module basic_1500_15000_2000_120_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_812,In_618);
xnor U1 (N_1,In_41,In_261);
xnor U2 (N_2,In_850,In_111);
nand U3 (N_3,In_143,In_668);
nand U4 (N_4,In_814,In_853);
nand U5 (N_5,In_862,In_1484);
xnor U6 (N_6,In_74,In_1000);
nor U7 (N_7,In_425,In_1248);
or U8 (N_8,In_1494,In_1451);
or U9 (N_9,In_108,In_1476);
nand U10 (N_10,In_212,In_1012);
or U11 (N_11,In_434,In_366);
and U12 (N_12,In_678,In_334);
nor U13 (N_13,In_153,In_441);
nor U14 (N_14,In_1060,In_1329);
xnor U15 (N_15,In_198,In_1445);
or U16 (N_16,In_134,In_624);
nor U17 (N_17,In_932,In_252);
xnor U18 (N_18,In_435,In_702);
nor U19 (N_19,In_698,In_682);
nand U20 (N_20,In_652,In_269);
xnor U21 (N_21,In_192,In_1303);
and U22 (N_22,In_625,In_1208);
or U23 (N_23,In_5,In_524);
nand U24 (N_24,In_283,In_273);
nor U25 (N_25,In_780,In_1374);
nor U26 (N_26,In_1061,In_1178);
nand U27 (N_27,In_681,In_117);
and U28 (N_28,In_1419,In_1467);
nor U29 (N_29,In_1073,In_1078);
nand U30 (N_30,In_555,In_1190);
nor U31 (N_31,In_287,In_34);
and U32 (N_32,In_1202,In_179);
xnor U33 (N_33,In_1225,In_878);
or U34 (N_34,In_952,In_1367);
nor U35 (N_35,In_552,In_772);
xor U36 (N_36,In_1007,In_68);
and U37 (N_37,In_712,In_1428);
xnor U38 (N_38,In_680,In_486);
and U39 (N_39,In_1294,In_172);
or U40 (N_40,In_962,In_351);
or U41 (N_41,In_1482,In_1145);
or U42 (N_42,In_1320,In_735);
xnor U43 (N_43,In_672,In_641);
and U44 (N_44,In_1010,In_245);
nor U45 (N_45,In_650,In_1097);
and U46 (N_46,In_859,In_1174);
and U47 (N_47,In_567,In_843);
and U48 (N_48,In_1126,In_515);
nor U49 (N_49,In_694,In_925);
xnor U50 (N_50,In_481,In_1412);
xor U51 (N_51,In_638,In_1459);
or U52 (N_52,In_185,In_1464);
or U53 (N_53,In_860,In_514);
xor U54 (N_54,In_464,In_232);
or U55 (N_55,In_1121,In_1328);
nor U56 (N_56,In_1474,In_1260);
nor U57 (N_57,In_1289,In_1159);
nand U58 (N_58,In_290,In_1353);
nand U59 (N_59,In_1239,In_762);
and U60 (N_60,In_851,In_332);
or U61 (N_61,In_297,In_568);
or U62 (N_62,In_1424,In_77);
nor U63 (N_63,In_765,In_258);
or U64 (N_64,In_1358,In_676);
nand U65 (N_65,In_651,In_1228);
xnor U66 (N_66,In_1258,In_661);
nand U67 (N_67,In_573,In_864);
and U68 (N_68,In_1259,In_386);
xor U69 (N_69,In_165,In_45);
or U70 (N_70,In_473,In_1483);
or U71 (N_71,In_353,In_855);
and U72 (N_72,In_385,In_1042);
xnor U73 (N_73,In_10,In_387);
nand U74 (N_74,In_873,In_622);
nand U75 (N_75,In_943,In_311);
xnor U76 (N_76,In_1344,In_240);
or U77 (N_77,In_299,In_688);
or U78 (N_78,In_1385,In_154);
and U79 (N_79,In_1296,In_1336);
or U80 (N_80,In_936,In_1216);
nand U81 (N_81,In_415,In_717);
xnor U82 (N_82,In_497,In_320);
or U83 (N_83,In_504,In_1172);
or U84 (N_84,In_1071,In_1312);
xnor U85 (N_85,In_1277,In_469);
or U86 (N_86,In_693,In_849);
nand U87 (N_87,In_699,In_1479);
nand U88 (N_88,In_583,In_163);
and U89 (N_89,In_1056,In_1346);
nand U90 (N_90,In_599,In_905);
or U91 (N_91,In_781,In_340);
xor U92 (N_92,In_912,In_1275);
nor U93 (N_93,In_364,In_1369);
nor U94 (N_94,In_646,In_1214);
xor U95 (N_95,In_49,In_725);
or U96 (N_96,In_23,In_731);
or U97 (N_97,In_136,In_1395);
nand U98 (N_98,In_35,In_671);
nand U99 (N_99,In_80,In_956);
and U100 (N_100,In_1351,In_1368);
nand U101 (N_101,In_1268,In_161);
and U102 (N_102,In_744,In_844);
nand U103 (N_103,In_257,In_1273);
or U104 (N_104,In_209,In_1106);
xor U105 (N_105,In_1249,In_101);
or U106 (N_106,In_0,In_1315);
and U107 (N_107,In_523,In_854);
and U108 (N_108,In_935,In_1408);
nor U109 (N_109,In_1447,In_1387);
nor U110 (N_110,In_1016,In_345);
nor U111 (N_111,In_1390,In_40);
or U112 (N_112,In_884,In_1107);
nor U113 (N_113,In_314,In_82);
nor U114 (N_114,In_1201,In_379);
xnor U115 (N_115,In_683,In_404);
nor U116 (N_116,In_405,In_592);
and U117 (N_117,In_895,In_748);
xor U118 (N_118,In_1188,In_1098);
and U119 (N_119,In_1195,In_992);
xnor U120 (N_120,In_217,In_1265);
xnor U121 (N_121,In_561,In_476);
and U122 (N_122,In_1077,In_141);
or U123 (N_123,In_708,In_424);
or U124 (N_124,In_381,In_426);
xnor U125 (N_125,In_871,In_915);
or U126 (N_126,In_380,N_120);
nand U127 (N_127,N_66,In_451);
and U128 (N_128,In_951,In_587);
and U129 (N_129,In_243,In_1182);
or U130 (N_130,N_10,In_317);
nand U131 (N_131,In_1354,N_62);
and U132 (N_132,In_1019,In_1095);
or U133 (N_133,N_94,In_1128);
nor U134 (N_134,In_689,In_1433);
nand U135 (N_135,In_253,N_27);
nor U136 (N_136,N_88,In_174);
nand U137 (N_137,N_57,In_1138);
and U138 (N_138,In_574,In_959);
and U139 (N_139,In_66,In_1438);
nand U140 (N_140,In_520,In_1123);
and U141 (N_141,In_178,In_1116);
nand U142 (N_142,In_1304,In_1376);
xnor U143 (N_143,In_865,In_1114);
xor U144 (N_144,In_103,In_1410);
nand U145 (N_145,In_737,In_1132);
xnor U146 (N_146,In_12,In_1119);
or U147 (N_147,In_743,In_642);
or U148 (N_148,In_118,In_532);
nor U149 (N_149,In_842,In_449);
or U150 (N_150,In_917,In_1231);
nor U151 (N_151,In_303,In_1161);
xor U152 (N_152,In_1052,In_350);
and U153 (N_153,In_83,In_966);
or U154 (N_154,In_1233,N_22);
nor U155 (N_155,In_116,In_1090);
nor U156 (N_156,In_1039,In_32);
and U157 (N_157,In_703,In_866);
nand U158 (N_158,In_1301,In_382);
xnor U159 (N_159,In_233,In_155);
nor U160 (N_160,In_439,In_110);
and U161 (N_161,In_633,In_869);
xor U162 (N_162,In_241,In_857);
nor U163 (N_163,In_392,In_191);
xor U164 (N_164,In_1244,In_1321);
and U165 (N_165,In_73,In_1285);
or U166 (N_166,In_1468,In_713);
xnor U167 (N_167,In_1238,In_896);
and U168 (N_168,In_1450,In_1025);
or U169 (N_169,In_1122,In_1261);
and U170 (N_170,In_626,In_766);
and U171 (N_171,In_8,In_1430);
xnor U172 (N_172,In_1490,In_824);
or U173 (N_173,In_557,In_1257);
and U174 (N_174,In_276,In_1462);
nand U175 (N_175,N_26,In_1453);
or U176 (N_176,In_13,In_503);
xor U177 (N_177,In_548,In_1488);
or U178 (N_178,In_230,In_655);
xor U179 (N_179,In_1324,In_937);
or U180 (N_180,In_540,In_911);
xnor U181 (N_181,In_1375,In_797);
nor U182 (N_182,In_675,In_1033);
xnor U183 (N_183,In_1271,In_304);
nand U184 (N_184,In_1302,In_341);
or U185 (N_185,In_816,In_827);
xor U186 (N_186,In_1082,In_354);
or U187 (N_187,In_1023,In_1064);
or U188 (N_188,In_1207,In_1074);
nor U189 (N_189,In_1256,In_938);
and U190 (N_190,In_121,In_443);
xnor U191 (N_191,In_1220,In_1309);
nor U192 (N_192,In_1327,In_156);
nor U193 (N_193,In_167,N_63);
xor U194 (N_194,In_128,In_531);
nor U195 (N_195,In_1036,In_1191);
nand U196 (N_196,N_76,In_833);
xnor U197 (N_197,In_566,In_742);
xnor U198 (N_198,In_750,N_7);
and U199 (N_199,N_90,In_280);
nand U200 (N_200,In_1196,In_899);
and U201 (N_201,In_1206,In_248);
or U202 (N_202,In_981,In_1499);
and U203 (N_203,In_1449,In_941);
and U204 (N_204,In_1030,In_611);
and U205 (N_205,In_1177,In_1135);
xor U206 (N_206,In_223,In_1396);
or U207 (N_207,In_919,In_769);
xor U208 (N_208,N_71,In_900);
nand U209 (N_209,In_547,In_886);
xnor U210 (N_210,In_856,In_57);
and U211 (N_211,In_31,In_1263);
xnor U212 (N_212,N_1,In_740);
or U213 (N_213,In_728,In_1144);
xor U214 (N_214,In_607,In_909);
or U215 (N_215,In_1429,N_100);
nor U216 (N_216,In_1293,In_1348);
or U217 (N_217,In_947,In_1165);
nand U218 (N_218,In_910,In_335);
nor U219 (N_219,In_1186,In_852);
nand U220 (N_220,In_997,In_228);
xor U221 (N_221,In_1209,In_333);
nand U222 (N_222,In_593,In_907);
nor U223 (N_223,In_898,In_272);
nand U224 (N_224,N_59,In_1470);
or U225 (N_225,In_640,In_199);
nor U226 (N_226,In_123,In_1330);
xor U227 (N_227,In_169,In_1218);
nand U228 (N_228,In_370,In_1065);
or U229 (N_229,N_8,In_104);
xnor U230 (N_230,In_554,In_724);
or U231 (N_231,In_205,In_1246);
nor U232 (N_232,In_183,In_994);
and U233 (N_233,In_489,In_444);
nor U234 (N_234,In_1437,In_1024);
nand U235 (N_235,In_914,In_1157);
nor U236 (N_236,In_648,In_792);
xnor U237 (N_237,In_1058,In_539);
nand U238 (N_238,N_17,N_43);
nor U239 (N_239,In_1146,N_97);
xnor U240 (N_240,In_202,In_391);
and U241 (N_241,In_85,In_926);
or U242 (N_242,In_358,In_100);
xnor U243 (N_243,In_578,N_30);
xor U244 (N_244,In_1099,N_92);
nand U245 (N_245,In_16,In_166);
and U246 (N_246,In_872,In_406);
nand U247 (N_247,In_928,In_470);
nor U248 (N_248,In_603,In_845);
nand U249 (N_249,In_7,In_1415);
or U250 (N_250,In_216,N_197);
nand U251 (N_251,In_1221,In_1264);
or U252 (N_252,In_563,In_1495);
or U253 (N_253,In_177,N_72);
or U254 (N_254,N_188,In_788);
xnor U255 (N_255,N_189,N_122);
or U256 (N_256,In_402,N_42);
or U257 (N_257,In_328,In_6);
nor U258 (N_258,In_53,In_58);
nand U259 (N_259,In_1487,In_1242);
and U260 (N_260,In_1362,N_109);
nand U261 (N_261,In_281,In_1020);
or U262 (N_262,N_127,In_56);
nand U263 (N_263,N_159,In_344);
or U264 (N_264,In_889,In_775);
nor U265 (N_265,N_231,In_1067);
or U266 (N_266,In_604,In_206);
nand U267 (N_267,In_374,N_37);
and U268 (N_268,In_739,N_244);
nor U269 (N_269,In_1226,In_600);
nor U270 (N_270,In_462,In_1401);
nor U271 (N_271,In_571,N_40);
or U272 (N_272,In_254,In_784);
xor U273 (N_273,In_1427,In_726);
xor U274 (N_274,N_241,In_870);
nand U275 (N_275,In_1109,In_802);
nor U276 (N_276,N_234,In_589);
nor U277 (N_277,N_143,In_946);
nand U278 (N_278,In_25,In_1147);
and U279 (N_279,N_207,In_764);
nand U280 (N_280,In_667,In_1291);
nand U281 (N_281,In_484,In_526);
and U282 (N_282,In_265,In_777);
xor U283 (N_283,N_85,In_1399);
or U284 (N_284,In_130,In_733);
nand U285 (N_285,In_623,In_767);
or U286 (N_286,In_1163,In_1469);
xnor U287 (N_287,In_863,In_1245);
xor U288 (N_288,In_591,In_1072);
nand U289 (N_289,N_131,In_21);
xor U290 (N_290,In_522,In_968);
and U291 (N_291,N_198,In_594);
and U292 (N_292,In_1381,In_270);
xor U293 (N_293,N_74,In_1267);
or U294 (N_294,In_569,In_1418);
nor U295 (N_295,In_643,In_1055);
xor U296 (N_296,In_90,In_953);
and U297 (N_297,In_54,In_830);
nand U298 (N_298,In_1241,In_882);
nand U299 (N_299,In_613,In_538);
nor U300 (N_300,In_975,N_78);
xor U301 (N_301,In_534,In_747);
and U302 (N_302,In_684,In_1115);
nand U303 (N_303,In_629,In_556);
xor U304 (N_304,In_420,In_1035);
and U305 (N_305,In_505,In_804);
nand U306 (N_306,In_499,In_806);
or U307 (N_307,In_431,N_21);
nand U308 (N_308,In_1306,In_355);
or U309 (N_309,In_239,In_348);
nand U310 (N_310,In_321,In_475);
xor U311 (N_311,In_1363,In_1085);
xor U312 (N_312,In_37,In_249);
xnor U313 (N_313,In_610,N_24);
or U314 (N_314,In_575,In_1466);
nand U315 (N_315,N_192,In_1);
or U316 (N_316,In_1409,In_368);
or U317 (N_317,In_89,N_205);
or U318 (N_318,In_418,N_248);
nor U319 (N_319,N_55,N_180);
and U320 (N_320,In_1153,In_969);
and U321 (N_321,N_69,In_175);
nand U322 (N_322,In_960,N_132);
nand U323 (N_323,In_398,In_729);
nor U324 (N_324,In_696,N_13);
and U325 (N_325,In_760,In_601);
nand U326 (N_326,In_933,In_581);
or U327 (N_327,In_1442,In_144);
or U328 (N_328,In_721,In_1425);
and U329 (N_329,In_986,In_536);
xnor U330 (N_330,In_944,In_302);
nor U331 (N_331,In_685,In_1211);
or U332 (N_332,In_263,N_181);
or U333 (N_333,In_989,N_106);
or U334 (N_334,In_1180,In_558);
or U335 (N_335,In_330,In_149);
nor U336 (N_336,In_244,In_300);
nand U337 (N_337,In_634,In_1370);
nor U338 (N_338,In_1287,In_663);
xor U339 (N_339,In_546,In_691);
or U340 (N_340,In_1156,In_468);
nor U341 (N_341,In_923,In_410);
and U342 (N_342,In_823,In_707);
nand U343 (N_343,In_1276,In_1152);
xor U344 (N_344,In_1102,In_140);
and U345 (N_345,N_151,In_1124);
xor U346 (N_346,In_709,In_33);
nor U347 (N_347,In_184,In_436);
xnor U348 (N_348,In_109,In_527);
nand U349 (N_349,In_614,In_700);
or U350 (N_350,In_1118,In_1377);
xnor U351 (N_351,In_1017,In_1011);
or U352 (N_352,In_876,In_590);
or U353 (N_353,In_1094,In_30);
nand U354 (N_354,N_134,In_846);
and U355 (N_355,N_163,In_112);
and U356 (N_356,In_1255,In_749);
and U357 (N_357,In_146,In_1334);
nor U358 (N_358,In_72,In_993);
nor U359 (N_359,N_39,In_1215);
or U360 (N_360,N_35,In_1444);
and U361 (N_361,In_649,In_437);
nand U362 (N_362,In_996,In_798);
and U363 (N_363,In_371,In_271);
and U364 (N_364,In_1021,In_606);
and U365 (N_365,In_1441,In_422);
or U366 (N_366,In_1359,In_978);
or U367 (N_367,In_832,N_28);
xnor U368 (N_368,In_1403,In_719);
and U369 (N_369,In_1254,N_200);
nor U370 (N_370,In_1069,In_372);
xnor U371 (N_371,In_602,In_450);
xor U372 (N_372,In_1050,In_231);
and U373 (N_373,In_1232,In_428);
nand U374 (N_374,In_949,In_1026);
nand U375 (N_375,In_879,In_483);
or U376 (N_376,In_746,N_211);
nand U377 (N_377,N_337,In_995);
and U378 (N_378,In_1179,N_36);
and U379 (N_379,N_339,In_461);
xnor U380 (N_380,In_1140,N_313);
nor U381 (N_381,In_782,In_874);
nor U382 (N_382,In_309,In_1197);
nand U383 (N_383,N_193,In_518);
xor U384 (N_384,In_357,In_401);
nand U385 (N_385,N_119,N_334);
xnor U386 (N_386,N_312,In_180);
nor U387 (N_387,N_270,In_1458);
nand U388 (N_388,In_1251,In_948);
or U389 (N_389,In_1333,In_562);
and U390 (N_390,In_38,In_736);
nor U391 (N_391,N_355,In_1372);
or U392 (N_392,In_757,N_250);
nor U393 (N_393,In_1461,N_343);
nor U394 (N_394,In_1100,In_564);
or U395 (N_395,In_1125,N_14);
and U396 (N_396,In_237,N_318);
or U397 (N_397,N_245,In_477);
and U398 (N_398,In_1027,In_324);
xnor U399 (N_399,N_147,N_70);
nor U400 (N_400,In_1093,N_52);
nor U401 (N_401,In_656,In_1292);
or U402 (N_402,In_1485,N_324);
nor U403 (N_403,In_129,In_247);
or U404 (N_404,N_172,N_82);
nand U405 (N_405,In_413,In_203);
or U406 (N_406,N_215,N_157);
nor U407 (N_407,N_38,N_144);
nand U408 (N_408,N_202,In_1166);
or U409 (N_409,In_1420,In_706);
nand U410 (N_410,In_1087,In_620);
xor U411 (N_411,In_868,N_262);
and U412 (N_412,In_412,In_1169);
and U413 (N_413,In_262,In_1005);
or U414 (N_414,In_1008,In_62);
nand U415 (N_415,N_110,In_268);
xnor U416 (N_416,N_148,In_1298);
nand U417 (N_417,In_388,N_206);
and U418 (N_418,In_984,In_1274);
and U419 (N_419,In_1373,N_289);
nand U420 (N_420,In_1394,In_463);
nor U421 (N_421,N_47,In_1253);
nand U422 (N_422,In_983,In_967);
nand U423 (N_423,In_697,In_195);
or U424 (N_424,N_259,In_342);
nand U425 (N_425,In_160,In_1240);
xnor U426 (N_426,In_1397,In_15);
or U427 (N_427,In_1084,In_487);
and U428 (N_428,In_1219,In_452);
and U429 (N_429,In_312,In_490);
xnor U430 (N_430,N_370,In_221);
nand U431 (N_431,N_116,In_791);
or U432 (N_432,N_102,In_403);
or U433 (N_433,N_89,In_211);
or U434 (N_434,In_881,In_1062);
or U435 (N_435,In_537,In_2);
nand U436 (N_436,N_208,N_167);
and U437 (N_437,In_1386,In_1319);
and U438 (N_438,N_301,In_138);
or U439 (N_439,In_295,In_1200);
nor U440 (N_440,N_166,N_284);
and U441 (N_441,In_1326,In_786);
and U442 (N_442,In_838,In_201);
nand U443 (N_443,N_347,In_1164);
nor U444 (N_444,In_27,In_1041);
nor U445 (N_445,In_194,In_349);
xor U446 (N_446,In_319,In_617);
nand U447 (N_447,N_306,In_474);
and U448 (N_448,N_235,In_596);
or U449 (N_449,N_133,In_1192);
xnor U450 (N_450,In_939,In_1391);
and U451 (N_451,N_277,N_117);
xor U452 (N_452,In_957,In_318);
or U453 (N_453,In_528,In_687);
and U454 (N_454,In_753,N_283);
nand U455 (N_455,N_209,In_60);
or U456 (N_456,N_137,In_819);
and U457 (N_457,N_366,In_550);
or U458 (N_458,In_847,In_510);
or U459 (N_459,In_1051,In_95);
and U460 (N_460,In_423,In_1371);
and U461 (N_461,In_390,In_972);
nor U462 (N_462,N_346,In_1141);
nand U463 (N_463,N_279,In_734);
nor U464 (N_464,In_584,N_152);
nand U465 (N_465,In_974,In_665);
or U466 (N_466,In_585,In_987);
nand U467 (N_467,In_456,In_1040);
nand U468 (N_468,In_18,In_480);
or U469 (N_469,N_265,In_1435);
nand U470 (N_470,In_1139,In_465);
or U471 (N_471,In_1431,In_376);
and U472 (N_472,In_107,In_517);
and U473 (N_473,In_466,In_24);
nor U474 (N_474,N_141,In_916);
nor U475 (N_475,In_378,In_255);
xor U476 (N_476,In_1343,N_150);
or U477 (N_477,In_97,In_647);
nand U478 (N_478,In_1160,N_121);
or U479 (N_479,In_1497,In_1443);
or U480 (N_480,In_285,N_365);
and U481 (N_481,N_276,In_331);
xnor U482 (N_482,In_1313,In_1400);
nor U483 (N_483,N_332,In_113);
nor U484 (N_484,In_1057,In_115);
or U485 (N_485,In_1383,In_52);
nand U486 (N_486,In_339,In_1170);
nor U487 (N_487,In_615,In_1493);
nand U488 (N_488,N_54,N_79);
nor U489 (N_489,In_1332,In_170);
and U490 (N_490,N_108,In_673);
or U491 (N_491,In_14,In_1158);
nor U492 (N_492,N_374,In_759);
and U493 (N_493,In_1411,N_367);
nor U494 (N_494,In_789,In_1189);
nor U495 (N_495,N_201,In_1352);
or U496 (N_496,N_83,In_861);
xor U497 (N_497,In_801,In_1213);
and U498 (N_498,In_137,In_87);
nand U499 (N_499,N_80,N_246);
xor U500 (N_500,N_380,In_1127);
nor U501 (N_501,N_187,In_39);
nand U502 (N_502,In_1492,In_373);
and U503 (N_503,In_512,N_194);
xnor U504 (N_504,N_56,In_472);
nand U505 (N_505,N_165,In_296);
nand U506 (N_506,In_1184,In_887);
nand U507 (N_507,In_940,In_807);
nand U508 (N_508,In_1338,In_529);
or U509 (N_509,In_674,In_1194);
and U510 (N_510,N_169,N_351);
or U511 (N_511,In_776,In_1181);
nor U512 (N_512,N_453,In_448);
nand U513 (N_513,N_302,In_1070);
nor U514 (N_514,In_400,N_352);
nand U515 (N_515,In_36,N_489);
nand U516 (N_516,In_1456,N_170);
and U517 (N_517,In_9,In_1108);
nand U518 (N_518,N_447,In_1001);
and U519 (N_519,In_1310,N_149);
and U520 (N_520,In_1129,In_551);
nand U521 (N_521,In_924,In_1053);
or U522 (N_522,N_432,N_232);
and U523 (N_523,In_1018,N_238);
and U524 (N_524,N_139,N_338);
xnor U525 (N_525,In_1288,N_140);
or U526 (N_526,In_1350,In_98);
nand U527 (N_527,In_65,In_1091);
nand U528 (N_528,In_930,In_1349);
nor U529 (N_529,N_423,In_901);
nand U530 (N_530,In_945,In_582);
xor U531 (N_531,In_1325,In_1342);
or U532 (N_532,In_1379,In_1171);
nand U533 (N_533,In_1227,In_579);
nand U534 (N_534,In_1199,In_365);
or U535 (N_535,In_577,N_376);
and U536 (N_536,N_326,In_695);
xnor U537 (N_537,N_178,In_720);
xor U538 (N_538,In_1299,N_60);
xor U539 (N_539,In_29,In_803);
nand U540 (N_540,In_525,In_1083);
or U541 (N_541,In_310,In_432);
xnor U542 (N_542,N_384,In_1339);
and U543 (N_543,In_1112,N_95);
nand U544 (N_544,In_215,N_493);
or U545 (N_545,N_462,In_608);
nor U546 (N_546,In_1079,In_1049);
and U547 (N_547,N_459,In_327);
nand U548 (N_548,In_825,In_1086);
nor U549 (N_549,N_34,In_394);
nand U550 (N_550,In_1407,In_159);
nor U551 (N_551,N_275,In_714);
xnor U552 (N_552,In_976,In_950);
nand U553 (N_553,In_1446,In_670);
nand U554 (N_554,In_1013,N_264);
xnor U555 (N_555,N_388,N_145);
or U556 (N_556,N_101,In_251);
nor U557 (N_557,In_1224,In_741);
or U558 (N_558,N_154,N_460);
and U559 (N_559,In_329,N_495);
xnor U560 (N_560,In_187,N_218);
xor U561 (N_561,In_369,In_1366);
xor U562 (N_562,In_999,In_811);
or U563 (N_563,N_426,In_190);
nand U564 (N_564,N_171,In_1281);
and U565 (N_565,In_471,In_131);
nand U566 (N_566,N_496,In_119);
nand U567 (N_567,In_289,In_307);
nor U568 (N_568,In_770,N_421);
nor U569 (N_569,N_411,In_210);
and U570 (N_570,In_507,In_222);
nor U571 (N_571,N_497,In_595);
xor U572 (N_572,N_320,In_457);
and U573 (N_573,N_282,In_384);
xnor U574 (N_574,In_1413,In_294);
nor U575 (N_575,N_229,In_1460);
and U576 (N_576,N_441,N_179);
xor U577 (N_577,In_1111,N_440);
nor U578 (N_578,In_71,N_473);
or U579 (N_579,In_875,N_399);
nand U580 (N_580,In_343,In_961);
or U581 (N_581,In_389,In_1496);
or U582 (N_582,In_888,In_704);
xnor U583 (N_583,In_1137,In_182);
nand U584 (N_584,In_1130,N_271);
xor U585 (N_585,In_1063,N_309);
nor U586 (N_586,In_396,N_240);
or U587 (N_587,In_570,N_216);
or U588 (N_588,In_157,In_1280);
and U589 (N_589,N_153,N_20);
nor U590 (N_590,N_331,In_745);
nand U591 (N_591,N_401,In_1162);
and U592 (N_592,N_297,N_203);
xor U593 (N_593,N_186,In_458);
xnor U594 (N_594,N_429,In_1038);
xnor U595 (N_595,In_282,In_841);
nand U596 (N_596,In_1471,In_1365);
nand U597 (N_597,In_632,In_47);
or U598 (N_598,In_877,N_373);
or U599 (N_599,N_44,In_277);
nor U600 (N_600,In_658,In_800);
nor U601 (N_601,In_653,In_1222);
xnor U602 (N_602,In_308,N_499);
xnor U603 (N_603,N_456,N_124);
or U604 (N_604,In_197,N_396);
and U605 (N_605,N_2,N_16);
or U606 (N_606,In_1175,In_1113);
xnor U607 (N_607,N_433,In_274);
xnor U608 (N_608,In_771,N_99);
and U609 (N_609,N_111,N_256);
and U610 (N_610,In_1034,In_235);
and U611 (N_611,N_257,In_1340);
and U612 (N_612,N_298,In_795);
or U613 (N_613,N_290,In_11);
and U614 (N_614,In_438,In_904);
or U615 (N_615,N_249,N_296);
nand U616 (N_616,N_303,In_158);
xnor U617 (N_617,N_104,In_453);
nor U618 (N_618,In_1266,In_1076);
xnor U619 (N_619,N_142,N_322);
xnor U620 (N_620,In_399,In_1167);
xor U621 (N_621,In_1131,In_1066);
or U622 (N_622,N_438,In_1089);
xnor U623 (N_623,In_1080,N_463);
nand U624 (N_624,N_41,N_458);
xnor U625 (N_625,N_443,N_603);
and U626 (N_626,N_305,In_836);
xnor U627 (N_627,In_774,N_417);
xnor U628 (N_628,N_457,N_602);
nand U629 (N_629,In_768,N_281);
nand U630 (N_630,N_316,In_1489);
nand U631 (N_631,N_442,In_711);
and U632 (N_632,In_1088,In_105);
and U633 (N_633,In_433,N_91);
or U634 (N_634,In_63,In_213);
or U635 (N_635,N_258,N_515);
or U636 (N_636,N_595,N_190);
nand U637 (N_637,N_222,In_67);
nand U638 (N_638,In_1388,In_1284);
or U639 (N_639,N_356,In_1380);
and U640 (N_640,N_474,N_414);
nand U641 (N_641,N_32,In_323);
nor U642 (N_642,N_540,In_1378);
xor U643 (N_643,In_894,N_183);
nor U644 (N_644,In_715,N_237);
nand U645 (N_645,In_164,In_662);
and U646 (N_646,In_70,In_26);
xnor U647 (N_647,In_171,In_727);
and U648 (N_648,In_635,In_1193);
or U649 (N_649,In_288,N_184);
and U650 (N_650,In_1002,N_6);
nand U651 (N_651,In_787,In_1250);
or U652 (N_652,In_597,In_834);
nand U653 (N_653,In_880,In_799);
or U654 (N_654,In_1203,In_560);
and U655 (N_655,In_619,In_1204);
xor U656 (N_656,In_442,N_562);
nand U657 (N_657,N_254,In_796);
xor U658 (N_658,In_250,In_502);
nand U659 (N_659,In_908,N_624);
or U660 (N_660,In_636,In_1475);
nand U661 (N_661,N_490,In_145);
and U662 (N_662,In_1237,N_113);
and U663 (N_663,In_347,N_379);
xnor U664 (N_664,N_561,In_1059);
xnor U665 (N_665,N_300,In_669);
or U666 (N_666,In_1223,In_409);
xnor U667 (N_667,In_511,N_185);
xnor U668 (N_668,N_476,In_1355);
nand U669 (N_669,In_207,N_393);
and U670 (N_670,N_466,In_586);
xnor U671 (N_671,In_1198,N_590);
nand U672 (N_672,In_1133,N_437);
or U673 (N_673,In_1295,In_723);
xor U674 (N_674,N_609,N_304);
nand U675 (N_675,In_1031,In_1455);
nor U676 (N_676,N_563,In_705);
and U677 (N_677,N_162,In_454);
or U678 (N_678,In_1143,In_751);
nor U679 (N_679,N_558,N_29);
xor U680 (N_680,N_576,In_659);
and U681 (N_681,In_848,In_565);
xnor U682 (N_682,In_92,N_9);
nor U683 (N_683,N_491,N_199);
nand U684 (N_684,In_132,In_1491);
xor U685 (N_685,In_1176,N_529);
and U686 (N_686,In_867,In_980);
nor U687 (N_687,In_42,In_1168);
and U688 (N_688,N_424,N_532);
nor U689 (N_689,N_330,N_543);
xor U690 (N_690,N_521,N_195);
xnor U691 (N_691,N_267,N_516);
nand U692 (N_692,In_660,In_1136);
nand U693 (N_693,In_1498,N_573);
xnor U694 (N_694,N_546,N_310);
nand U695 (N_695,In_542,In_1149);
or U696 (N_696,In_48,N_616);
nand U697 (N_697,N_416,N_418);
xnor U698 (N_698,In_716,In_1044);
nand U699 (N_699,N_556,N_353);
nand U700 (N_700,N_177,N_481);
and U701 (N_701,N_554,In_892);
or U702 (N_702,N_588,In_421);
nand U703 (N_703,N_219,In_971);
xnor U704 (N_704,In_1448,N_251);
nor U705 (N_705,N_511,N_571);
nand U706 (N_706,In_686,In_1457);
nor U707 (N_707,In_1361,In_1414);
nor U708 (N_708,In_785,N_239);
nand U709 (N_709,N_160,N_504);
and U710 (N_710,In_447,N_445);
or U711 (N_711,N_357,In_51);
nor U712 (N_712,N_314,In_1272);
nor U713 (N_713,N_484,N_98);
and U714 (N_714,N_175,N_549);
nor U715 (N_715,N_377,N_360);
and U716 (N_716,In_1434,In_1432);
nand U717 (N_717,N_252,N_514);
and U718 (N_718,In_730,N_286);
xor U719 (N_719,N_621,N_579);
nand U720 (N_720,In_1426,In_1117);
and U721 (N_721,In_1045,In_1205);
nand U722 (N_722,In_970,In_28);
and U723 (N_723,In_88,N_327);
and U724 (N_724,N_253,In_1230);
xnor U725 (N_725,In_1183,N_378);
and U726 (N_726,N_622,In_440);
and U727 (N_727,N_548,N_323);
nor U728 (N_728,In_267,In_91);
xnor U729 (N_729,N_526,In_152);
or U730 (N_730,In_543,N_299);
nor U731 (N_731,N_400,In_220);
or U732 (N_732,N_483,N_394);
and U733 (N_733,In_1290,In_305);
nor U734 (N_734,N_212,In_752);
and U735 (N_735,N_371,In_408);
nor U736 (N_736,In_122,N_115);
or U737 (N_737,N_553,N_492);
or U738 (N_738,N_451,N_449);
and U739 (N_739,In_831,N_507);
nor U740 (N_740,In_954,N_31);
xor U741 (N_741,In_106,N_584);
nand U742 (N_742,In_78,In_580);
or U743 (N_743,In_918,In_186);
xor U744 (N_744,In_363,N_512);
nand U745 (N_745,N_341,N_68);
nor U746 (N_746,N_412,In_494);
or U747 (N_747,N_223,N_176);
nand U748 (N_748,N_84,N_502);
and U749 (N_749,N_509,In_275);
xnor U750 (N_750,N_221,In_1006);
xnor U751 (N_751,In_459,In_151);
and U752 (N_752,N_4,In_559);
nor U753 (N_753,N_233,In_778);
nand U754 (N_754,In_236,In_417);
or U755 (N_755,In_1092,In_99);
nor U756 (N_756,In_509,In_1028);
nand U757 (N_757,In_313,N_53);
nor U758 (N_758,N_669,In_322);
nand U759 (N_759,N_674,In_1279);
or U760 (N_760,In_1402,In_55);
xnor U761 (N_761,In_1307,In_891);
xor U762 (N_762,N_670,In_20);
nor U763 (N_763,In_1212,In_1105);
nand U764 (N_764,N_648,N_475);
or U765 (N_765,N_720,N_395);
nand U766 (N_766,N_123,N_684);
or U767 (N_767,N_642,N_582);
or U768 (N_768,In_1142,N_263);
and U769 (N_769,N_643,N_217);
xnor U770 (N_770,N_587,In_1465);
nor U771 (N_771,In_1477,N_520);
and U772 (N_772,N_164,In_906);
nand U773 (N_773,In_1150,N_604);
nor U774 (N_774,N_628,N_130);
nor U775 (N_775,N_708,In_126);
and U776 (N_776,N_555,N_537);
xor U777 (N_777,N_358,In_902);
or U778 (N_778,In_316,N_640);
or U779 (N_779,N_717,N_311);
xnor U780 (N_780,In_84,In_718);
nor U781 (N_781,In_1269,N_699);
or U782 (N_782,N_444,N_636);
xnor U783 (N_783,N_420,N_652);
nor U784 (N_784,In_1185,In_616);
xor U785 (N_785,N_292,In_127);
xnor U786 (N_786,In_142,In_1236);
nor U787 (N_787,In_1405,N_125);
and U788 (N_788,N_614,N_733);
nand U789 (N_789,N_278,In_291);
nand U790 (N_790,N_431,N_634);
nand U791 (N_791,N_517,N_693);
nand U792 (N_792,N_606,In_1043);
nor U793 (N_793,In_260,In_1217);
and U794 (N_794,N_3,In_1104);
xor U795 (N_795,In_93,In_982);
and U796 (N_796,N_405,In_645);
xor U797 (N_797,N_578,N_738);
nor U798 (N_798,N_610,N_691);
or U799 (N_799,In_1037,In_1081);
nand U800 (N_800,N_452,In_493);
nand U801 (N_801,In_738,N_538);
and U802 (N_802,N_46,In_631);
nand U803 (N_803,N_227,N_138);
or U804 (N_804,In_988,N_630);
nor U805 (N_805,N_747,In_783);
nand U806 (N_806,In_1384,In_927);
nor U807 (N_807,N_719,In_664);
and U808 (N_808,N_505,In_521);
xnor U809 (N_809,N_0,N_385);
or U810 (N_810,In_120,N_247);
nor U811 (N_811,In_1341,In_858);
nand U812 (N_812,In_1393,In_478);
and U813 (N_813,N_406,In_114);
nand U814 (N_814,N_435,In_1439);
nand U815 (N_815,N_654,N_103);
or U816 (N_816,N_403,N_408);
and U817 (N_817,N_18,N_48);
and U818 (N_818,N_274,In_754);
or U819 (N_819,In_654,N_651);
nand U820 (N_820,In_506,In_407);
nand U821 (N_821,N_308,N_19);
nand U822 (N_822,N_173,In_377);
nand U823 (N_823,N_523,In_414);
nand U824 (N_824,N_748,N_409);
nor U825 (N_825,In_820,N_534);
or U826 (N_826,N_81,N_398);
nor U827 (N_827,N_629,N_354);
and U828 (N_828,N_687,N_392);
and U829 (N_829,In_979,In_773);
or U830 (N_830,N_464,N_557);
and U831 (N_831,N_702,In_793);
nor U832 (N_832,N_665,N_577);
nand U833 (N_833,N_655,N_689);
xnor U834 (N_834,N_469,In_965);
xnor U835 (N_835,In_1068,N_633);
nor U836 (N_836,In_492,N_448);
xnor U837 (N_837,In_533,N_740);
xnor U838 (N_838,In_1337,N_386);
nand U839 (N_839,In_495,N_461);
or U840 (N_840,In_942,N_93);
and U841 (N_841,In_627,N_524);
nand U842 (N_842,N_383,N_598);
nor U843 (N_843,In_498,In_813);
xor U844 (N_844,N_713,N_488);
and U845 (N_845,N_572,N_182);
nand U846 (N_846,In_485,In_284);
nand U847 (N_847,In_1360,N_696);
or U848 (N_848,N_112,In_1075);
nand U849 (N_849,N_204,In_612);
and U850 (N_850,N_430,In_1029);
nor U851 (N_851,N_23,N_480);
nand U852 (N_852,N_397,N_745);
or U853 (N_853,N_725,In_1382);
nor U854 (N_854,N_721,N_64);
nor U855 (N_855,In_214,N_653);
and U856 (N_856,N_333,In_826);
and U857 (N_857,In_508,In_790);
nor U858 (N_858,In_1323,In_359);
or U859 (N_859,N_638,N_319);
and U860 (N_860,In_1046,In_903);
nand U861 (N_861,In_541,N_716);
and U862 (N_862,N_731,N_618);
and U863 (N_863,In_779,N_710);
xnor U864 (N_864,N_294,N_735);
xnor U865 (N_865,N_506,In_278);
or U866 (N_866,N_11,In_416);
xnor U867 (N_867,N_498,N_711);
or U868 (N_868,In_991,In_19);
nand U869 (N_869,In_1436,In_929);
nor U870 (N_870,N_369,In_352);
xnor U871 (N_871,N_96,N_695);
nor U872 (N_872,N_288,N_706);
and U873 (N_873,In_488,N_161);
or U874 (N_874,N_340,In_1283);
nand U875 (N_875,N_734,N_800);
nand U876 (N_876,In_279,N_861);
and U877 (N_877,N_873,In_955);
nand U878 (N_878,N_685,N_847);
xor U879 (N_879,N_754,In_200);
nand U880 (N_880,In_446,In_383);
xnor U881 (N_881,N_865,N_677);
or U882 (N_882,N_839,N_678);
nor U883 (N_883,In_1480,In_79);
nand U884 (N_884,N_465,In_609);
or U885 (N_885,In_292,N_750);
xnor U886 (N_886,In_829,In_298);
xnor U887 (N_887,In_840,In_293);
nand U888 (N_888,In_922,N_782);
and U889 (N_889,N_761,In_460);
nand U890 (N_890,In_549,In_148);
or U891 (N_891,N_807,In_69);
nor U892 (N_892,N_454,N_228);
nand U893 (N_893,In_818,N_868);
nor U894 (N_894,N_671,In_1014);
nor U895 (N_895,In_1252,N_513);
xnor U896 (N_896,N_802,In_338);
nor U897 (N_897,N_649,N_501);
or U898 (N_898,N_518,N_773);
nor U899 (N_899,In_822,N_597);
and U900 (N_900,N_51,N_784);
nand U901 (N_901,N_820,In_1347);
xor U902 (N_902,N_382,N_389);
nand U903 (N_903,In_124,N_639);
or U904 (N_904,N_823,In_1154);
nor U905 (N_905,In_1416,N_220);
nand U906 (N_906,N_236,In_1357);
or U907 (N_907,N_762,In_931);
or U908 (N_908,N_841,N_350);
or U909 (N_909,N_805,In_1187);
xnor U910 (N_910,N_730,N_174);
nand U911 (N_911,N_830,In_1364);
nand U912 (N_912,In_1478,In_1243);
or U913 (N_913,N_856,N_478);
nor U914 (N_914,In_3,N_594);
and U915 (N_915,N_471,N_439);
or U916 (N_916,N_809,N_567);
nand U917 (N_917,N_790,In_920);
or U918 (N_918,In_692,N_568);
and U919 (N_919,N_566,N_419);
nand U920 (N_920,N_860,N_752);
and U921 (N_921,N_759,N_600);
nand U922 (N_922,N_105,N_844);
xor U923 (N_923,In_810,N_785);
nand U924 (N_924,In_1282,In_897);
and U925 (N_925,In_362,N_615);
or U926 (N_926,N_210,N_328);
nor U927 (N_927,In_1054,In_1210);
or U928 (N_928,In_218,In_817);
nand U929 (N_929,In_196,N_118);
nor U930 (N_930,N_834,In_375);
nor U931 (N_931,N_260,N_843);
and U932 (N_932,N_362,N_751);
nor U933 (N_933,N_852,N_704);
or U934 (N_934,N_547,N_683);
or U935 (N_935,N_833,In_1335);
or U936 (N_936,N_620,In_17);
xor U937 (N_937,In_598,In_535);
or U938 (N_938,In_679,In_1278);
and U939 (N_939,N_269,N_519);
nand U940 (N_940,N_701,In_605);
nor U941 (N_941,In_1314,N_857);
and U942 (N_942,In_1262,N_827);
and U943 (N_943,In_1322,In_1173);
and U944 (N_944,In_135,N_477);
or U945 (N_945,In_755,In_576);
nand U946 (N_946,N_77,N_372);
nand U947 (N_947,N_273,N_659);
xnor U948 (N_948,N_770,N_774);
xor U949 (N_949,In_1286,N_824);
xor U950 (N_950,In_337,N_5);
nand U951 (N_951,N_156,N_535);
nand U952 (N_952,In_809,In_963);
nand U953 (N_953,N_336,N_818);
nor U954 (N_954,N_552,In_1300);
nor U955 (N_955,In_139,N_436);
or U956 (N_956,N_560,N_612);
and U957 (N_957,N_613,N_317);
xnor U958 (N_958,N_635,N_344);
xnor U959 (N_959,N_407,N_832);
nor U960 (N_960,N_874,N_742);
nor U961 (N_961,N_87,N_255);
nor U962 (N_962,N_291,In_1317);
or U963 (N_963,N_863,In_637);
xor U964 (N_964,N_591,N_789);
and U965 (N_965,In_921,In_189);
or U966 (N_966,In_1009,N_842);
xor U967 (N_967,N_690,N_455);
nor U968 (N_968,In_1015,In_794);
nand U969 (N_969,In_1229,In_1234);
nand U970 (N_970,In_50,N_345);
nand U971 (N_971,In_973,In_1270);
and U972 (N_972,In_501,In_227);
and U973 (N_973,N_410,In_516);
nand U974 (N_974,In_1389,N_315);
xor U975 (N_975,In_934,N_242);
nor U976 (N_976,N_527,In_1101);
nor U977 (N_977,In_229,N_722);
or U978 (N_978,N_619,N_681);
xor U979 (N_979,N_530,N_726);
nor U980 (N_980,N_810,N_680);
nand U981 (N_981,N_812,In_958);
nor U982 (N_982,In_496,N_65);
or U983 (N_983,In_722,In_1148);
or U984 (N_984,N_335,N_467);
xor U985 (N_985,In_76,In_86);
or U986 (N_986,N_817,N_574);
xor U987 (N_987,In_1110,N_415);
and U988 (N_988,N_381,N_661);
xor U989 (N_989,In_208,N_826);
xnor U990 (N_990,N_698,N_829);
nor U991 (N_991,N_375,N_623);
or U992 (N_992,In_821,N_487);
and U993 (N_993,N_243,N_589);
nor U994 (N_994,In_883,N_136);
nor U995 (N_995,N_508,In_500);
xnor U996 (N_996,N_539,N_126);
and U997 (N_997,N_349,N_592);
xor U998 (N_998,In_168,N_570);
nand U999 (N_999,N_272,N_544);
and U1000 (N_1000,In_256,N_886);
and U1001 (N_1001,N_766,N_510);
nor U1002 (N_1002,N_956,In_701);
and U1003 (N_1003,In_411,N_872);
and U1004 (N_1004,N_895,N_268);
xor U1005 (N_1005,N_736,N_902);
or U1006 (N_1006,In_1331,N_927);
nor U1007 (N_1007,N_917,In_977);
nand U1008 (N_1008,N_811,N_884);
xnor U1009 (N_1009,N_565,N_676);
nand U1010 (N_1010,In_64,In_361);
or U1011 (N_1011,N_878,N_788);
nand U1012 (N_1012,N_828,N_960);
nor U1013 (N_1013,In_286,N_786);
nand U1014 (N_1014,In_427,N_976);
and U1015 (N_1015,N_743,N_993);
xor U1016 (N_1016,N_225,N_325);
or U1017 (N_1017,N_931,N_666);
nand U1018 (N_1018,In_1398,N_368);
or U1019 (N_1019,In_1481,In_828);
or U1020 (N_1020,N_67,N_937);
and U1021 (N_1021,N_107,N_816);
and U1022 (N_1022,N_894,N_718);
or U1023 (N_1023,N_694,N_775);
nor U1024 (N_1024,N_348,N_196);
and U1025 (N_1025,In_1454,In_1103);
nor U1026 (N_1026,N_470,In_1004);
nand U1027 (N_1027,In_758,N_391);
and U1028 (N_1028,In_1297,N_550);
nand U1029 (N_1029,N_974,In_188);
xnor U1030 (N_1030,N_575,In_360);
nor U1031 (N_1031,N_764,N_798);
nor U1032 (N_1032,N_660,In_44);
xor U1033 (N_1033,In_690,N_961);
nand U1034 (N_1034,In_419,N_755);
nand U1035 (N_1035,N_985,In_491);
nand U1036 (N_1036,In_346,N_646);
nand U1037 (N_1037,In_242,In_445);
xnor U1038 (N_1038,N_768,N_970);
or U1039 (N_1039,In_102,N_864);
or U1040 (N_1040,N_58,N_61);
nor U1041 (N_1041,In_393,N_915);
and U1042 (N_1042,N_923,In_479);
and U1043 (N_1043,In_234,N_907);
nand U1044 (N_1044,N_982,In_544);
nor U1045 (N_1045,N_583,N_942);
xnor U1046 (N_1046,N_213,In_985);
and U1047 (N_1047,N_968,In_224);
nand U1048 (N_1048,N_962,N_767);
or U1049 (N_1049,N_697,N_12);
nand U1050 (N_1050,N_758,In_1392);
nor U1051 (N_1051,In_588,N_975);
nor U1052 (N_1052,In_482,N_954);
nor U1053 (N_1053,N_819,N_724);
and U1054 (N_1054,N_607,N_536);
or U1055 (N_1055,N_771,N_932);
xor U1056 (N_1056,In_763,In_572);
nand U1057 (N_1057,N_280,In_395);
and U1058 (N_1058,In_181,In_1421);
and U1059 (N_1059,N_953,In_429);
xor U1060 (N_1060,N_808,N_542);
and U1061 (N_1061,N_869,N_285);
xor U1062 (N_1062,N_723,In_367);
nor U1063 (N_1063,N_984,N_627);
and U1064 (N_1064,In_553,In_204);
xnor U1065 (N_1065,In_226,In_325);
and U1066 (N_1066,N_796,N_73);
xor U1067 (N_1067,N_641,In_125);
nor U1068 (N_1068,N_364,N_679);
nand U1069 (N_1069,In_133,N_664);
and U1070 (N_1070,In_315,N_593);
nor U1071 (N_1071,N_925,N_715);
and U1072 (N_1072,N_129,N_760);
xor U1073 (N_1073,In_657,In_301);
xor U1074 (N_1074,N_230,In_639);
and U1075 (N_1075,N_293,N_935);
and U1076 (N_1076,N_605,N_50);
or U1077 (N_1077,N_893,N_998);
nand U1078 (N_1078,In_455,N_929);
or U1079 (N_1079,N_128,In_893);
xor U1080 (N_1080,N_995,N_662);
nand U1081 (N_1081,N_799,N_855);
xor U1082 (N_1082,N_737,N_657);
nand U1083 (N_1083,N_950,N_986);
and U1084 (N_1084,N_645,N_906);
nand U1085 (N_1085,N_783,N_892);
nand U1086 (N_1086,N_632,N_965);
and U1087 (N_1087,N_991,In_1345);
nor U1088 (N_1088,In_162,N_941);
xor U1089 (N_1089,N_155,N_806);
nor U1090 (N_1090,N_887,N_851);
nor U1091 (N_1091,N_647,In_513);
and U1092 (N_1092,N_971,N_821);
xnor U1093 (N_1093,In_964,N_191);
or U1094 (N_1094,N_390,N_531);
nor U1095 (N_1095,N_926,N_997);
nor U1096 (N_1096,N_434,N_479);
nor U1097 (N_1097,In_1463,N_825);
or U1098 (N_1098,N_911,N_940);
nand U1099 (N_1099,N_939,N_933);
or U1100 (N_1100,N_813,N_329);
nor U1101 (N_1101,N_972,N_703);
nand U1102 (N_1102,In_238,N_787);
nand U1103 (N_1103,N_224,In_1318);
or U1104 (N_1104,N_934,In_666);
and U1105 (N_1105,N_601,N_686);
nand U1106 (N_1106,In_306,N_528);
nand U1107 (N_1107,N_608,N_992);
xor U1108 (N_1108,N_503,N_904);
xor U1109 (N_1109,N_994,In_1311);
nand U1110 (N_1110,In_61,N_650);
or U1111 (N_1111,N_831,In_173);
nand U1112 (N_1112,N_114,N_321);
and U1113 (N_1113,N_919,In_264);
or U1114 (N_1114,N_541,In_890);
xnor U1115 (N_1115,N_778,N_744);
or U1116 (N_1116,N_891,N_692);
xor U1117 (N_1117,N_500,In_219);
or U1118 (N_1118,N_146,In_990);
nor U1119 (N_1119,N_900,N_672);
or U1120 (N_1120,N_885,N_836);
xnor U1121 (N_1121,N_880,N_402);
nand U1122 (N_1122,N_815,In_1096);
xor U1123 (N_1123,N_955,N_631);
xor U1124 (N_1124,N_947,N_978);
and U1125 (N_1125,N_525,N_1078);
nand U1126 (N_1126,N_472,In_1423);
xor U1127 (N_1127,N_1077,N_1003);
nand U1128 (N_1128,In_1452,In_1305);
or U1129 (N_1129,In_677,In_1247);
xor U1130 (N_1130,N_1072,N_753);
xnor U1131 (N_1131,N_996,N_1062);
nor U1132 (N_1132,N_795,N_1037);
or U1133 (N_1133,N_75,N_727);
or U1134 (N_1134,N_564,N_1036);
nand U1135 (N_1135,N_921,N_1073);
nand U1136 (N_1136,In_1308,N_1080);
xor U1137 (N_1137,N_875,N_404);
nor U1138 (N_1138,In_430,In_644);
and U1139 (N_1139,N_1123,In_1417);
or U1140 (N_1140,N_746,N_545);
xor U1141 (N_1141,N_876,N_909);
or U1142 (N_1142,N_700,N_903);
nand U1143 (N_1143,N_944,N_1020);
nand U1144 (N_1144,In_1155,N_1068);
and U1145 (N_1145,N_1093,N_990);
nor U1146 (N_1146,In_96,In_81);
xnor U1147 (N_1147,N_780,N_599);
xnor U1148 (N_1148,N_848,N_776);
nand U1149 (N_1149,N_980,N_1049);
xnor U1150 (N_1150,N_757,N_989);
and U1151 (N_1151,N_625,N_675);
or U1152 (N_1152,In_59,N_896);
xnor U1153 (N_1153,N_1015,In_4);
xnor U1154 (N_1154,N_1004,N_611);
or U1155 (N_1155,N_422,N_881);
or U1156 (N_1156,N_1007,N_261);
and U1157 (N_1157,N_1032,N_1091);
nor U1158 (N_1158,N_1075,N_1056);
xnor U1159 (N_1159,N_1070,N_1053);
nor U1160 (N_1160,N_1011,In_397);
or U1161 (N_1161,N_1101,N_226);
and U1162 (N_1162,In_1032,N_952);
nand U1163 (N_1163,N_801,N_1081);
nand U1164 (N_1164,N_1122,N_287);
nor U1165 (N_1165,N_663,N_916);
nand U1166 (N_1166,N_967,N_1117);
nand U1167 (N_1167,N_1017,N_494);
xnor U1168 (N_1168,N_918,N_1066);
or U1169 (N_1169,N_772,N_1047);
xnor U1170 (N_1170,N_951,In_1316);
nor U1171 (N_1171,N_1100,N_1031);
nor U1172 (N_1172,N_853,N_729);
or U1173 (N_1173,N_797,N_1046);
nor U1174 (N_1174,N_1110,In_22);
or U1175 (N_1175,N_596,N_763);
xnor U1176 (N_1176,N_977,In_326);
nor U1177 (N_1177,N_1088,N_854);
or U1178 (N_1178,In_519,N_946);
and U1179 (N_1179,In_530,In_1472);
nor U1180 (N_1180,N_33,N_359);
nor U1181 (N_1181,N_964,In_1134);
and U1182 (N_1182,In_815,N_1067);
nand U1183 (N_1183,N_769,N_866);
and U1184 (N_1184,In_150,N_1112);
xor U1185 (N_1185,N_658,N_551);
nor U1186 (N_1186,N_957,N_1090);
and U1187 (N_1187,N_1043,N_1098);
or U1188 (N_1188,N_1019,N_1113);
nor U1189 (N_1189,In_621,N_1039);
xor U1190 (N_1190,N_1001,N_981);
xnor U1191 (N_1191,In_1404,N_1065);
nand U1192 (N_1192,N_1054,N_883);
or U1193 (N_1193,N_1027,In_225);
nand U1194 (N_1194,In_1151,In_1440);
nor U1195 (N_1195,In_266,N_882);
or U1196 (N_1196,N_1087,N_682);
and U1197 (N_1197,N_846,N_850);
and U1198 (N_1198,N_1074,N_533);
or U1199 (N_1199,In_913,In_467);
nand U1200 (N_1200,N_342,N_862);
xor U1201 (N_1201,N_913,N_728);
or U1202 (N_1202,N_837,N_1086);
and U1203 (N_1203,N_936,In_1235);
nor U1204 (N_1204,N_1022,In_732);
xnor U1205 (N_1205,N_1096,N_45);
xnor U1206 (N_1206,N_1069,N_1044);
or U1207 (N_1207,N_793,In_710);
and U1208 (N_1208,In_75,N_1042);
nor U1209 (N_1209,N_1094,N_1120);
nor U1210 (N_1210,N_914,N_450);
nor U1211 (N_1211,N_1041,N_135);
xor U1212 (N_1212,N_1033,In_835);
nor U1213 (N_1213,N_1048,N_1005);
and U1214 (N_1214,N_814,N_673);
and U1215 (N_1215,N_581,N_899);
nand U1216 (N_1216,N_1103,N_973);
nor U1217 (N_1217,N_1124,N_963);
or U1218 (N_1218,N_1106,N_1063);
nor U1219 (N_1219,N_1089,N_979);
or U1220 (N_1220,N_1055,N_1104);
nand U1221 (N_1221,N_428,N_668);
nand U1222 (N_1222,N_688,N_867);
nor U1223 (N_1223,N_266,In_176);
xnor U1224 (N_1224,N_889,N_1012);
or U1225 (N_1225,N_949,N_1040);
nor U1226 (N_1226,N_779,N_1097);
or U1227 (N_1227,N_1076,N_765);
or U1228 (N_1228,In_805,N_413);
and U1229 (N_1229,N_707,N_361);
and U1230 (N_1230,N_749,N_667);
and U1231 (N_1231,N_930,N_791);
nand U1232 (N_1232,N_1116,N_468);
or U1233 (N_1233,N_1084,N_637);
or U1234 (N_1234,N_1008,N_656);
nand U1235 (N_1235,N_898,In_545);
or U1236 (N_1236,In_147,N_1108);
or U1237 (N_1237,N_1038,N_168);
nand U1238 (N_1238,N_1071,N_1114);
xor U1239 (N_1239,In_336,N_1009);
nor U1240 (N_1240,N_870,N_845);
and U1241 (N_1241,N_485,N_1035);
nand U1242 (N_1242,N_482,In_1003);
or U1243 (N_1243,N_905,In_94);
or U1244 (N_1244,N_969,N_25);
nor U1245 (N_1245,In_998,N_959);
xor U1246 (N_1246,N_943,N_1052);
xor U1247 (N_1247,N_569,N_1102);
nand U1248 (N_1248,In_756,N_948);
nand U1249 (N_1249,N_363,N_1000);
or U1250 (N_1250,N_987,N_486);
nor U1251 (N_1251,N_1230,N_1030);
nand U1252 (N_1252,N_1142,N_1132);
and U1253 (N_1253,In_837,N_1175);
and U1254 (N_1254,N_1216,N_1194);
xnor U1255 (N_1255,N_1095,N_158);
or U1256 (N_1256,N_1228,N_1184);
and U1257 (N_1257,N_803,N_859);
nor U1258 (N_1258,N_1179,N_1134);
nand U1259 (N_1259,N_999,N_1024);
xor U1260 (N_1260,N_425,N_1143);
and U1261 (N_1261,N_1025,N_644);
xor U1262 (N_1262,N_1236,In_630);
nor U1263 (N_1263,N_1183,N_804);
nor U1264 (N_1264,In_1120,N_1127);
xnor U1265 (N_1265,N_705,N_1204);
and U1266 (N_1266,N_1199,N_908);
nand U1267 (N_1267,N_1151,In_885);
nand U1268 (N_1268,N_781,N_945);
nand U1269 (N_1269,N_1176,N_1177);
or U1270 (N_1270,N_15,N_1131);
nand U1271 (N_1271,N_1152,N_1156);
nor U1272 (N_1272,N_617,N_1163);
and U1273 (N_1273,N_585,N_1150);
xor U1274 (N_1274,N_792,N_840);
nand U1275 (N_1275,N_714,N_1197);
and U1276 (N_1276,N_1168,N_1119);
nor U1277 (N_1277,N_1013,N_835);
nor U1278 (N_1278,In_1047,N_1018);
and U1279 (N_1279,N_928,N_1010);
nand U1280 (N_1280,N_1059,In_1048);
nand U1281 (N_1281,N_580,N_1164);
nor U1282 (N_1282,N_1219,N_1153);
or U1283 (N_1283,N_1006,In_1022);
xor U1284 (N_1284,N_1105,N_1173);
xnor U1285 (N_1285,N_1092,N_1185);
xnor U1286 (N_1286,N_1028,N_1130);
or U1287 (N_1287,N_924,N_888);
and U1288 (N_1288,N_1170,N_1212);
nor U1289 (N_1289,N_1058,N_1227);
nand U1290 (N_1290,N_1180,In_628);
and U1291 (N_1291,N_1158,N_1202);
and U1292 (N_1292,N_938,N_1211);
or U1293 (N_1293,N_877,N_1237);
or U1294 (N_1294,N_741,N_1026);
xor U1295 (N_1295,N_920,N_777);
nor U1296 (N_1296,N_1154,N_1169);
nand U1297 (N_1297,N_1162,N_1051);
or U1298 (N_1298,N_1165,N_1213);
xor U1299 (N_1299,N_1235,N_1160);
xor U1300 (N_1300,N_1016,N_1107);
xor U1301 (N_1301,N_1217,In_246);
xnor U1302 (N_1302,N_822,N_1246);
nor U1303 (N_1303,N_1083,N_1140);
xnor U1304 (N_1304,N_1243,N_1193);
or U1305 (N_1305,N_1157,N_1190);
nor U1306 (N_1306,N_1135,N_912);
xnor U1307 (N_1307,N_1182,N_1224);
xor U1308 (N_1308,N_1233,N_739);
xnor U1309 (N_1309,N_1146,N_1231);
nor U1310 (N_1310,N_1208,N_1002);
nor U1311 (N_1311,N_966,N_586);
nand U1312 (N_1312,N_49,N_1172);
nand U1313 (N_1313,N_1192,N_1247);
xor U1314 (N_1314,N_1045,N_732);
or U1315 (N_1315,N_1191,N_1206);
and U1316 (N_1316,N_1242,N_1220);
and U1317 (N_1317,N_1189,N_879);
nand U1318 (N_1318,In_1473,N_1136);
xor U1319 (N_1319,N_1126,N_1159);
xor U1320 (N_1320,N_1215,N_1244);
or U1321 (N_1321,N_709,In_1486);
xnor U1322 (N_1322,N_1171,N_712);
nor U1323 (N_1323,N_1121,N_1207);
nor U1324 (N_1324,N_1148,N_1249);
and U1325 (N_1325,N_1226,N_1205);
nor U1326 (N_1326,N_922,N_295);
nor U1327 (N_1327,N_1029,In_46);
and U1328 (N_1328,N_1223,N_756);
nor U1329 (N_1329,In_193,N_1210);
and U1330 (N_1330,N_958,N_1085);
or U1331 (N_1331,N_1050,N_1023);
xnor U1332 (N_1332,N_626,N_1060);
and U1333 (N_1333,In_43,N_1128);
xnor U1334 (N_1334,N_1167,N_1221);
and U1335 (N_1335,In_1422,N_86);
or U1336 (N_1336,N_1203,N_1225);
and U1337 (N_1337,N_1137,N_1238);
or U1338 (N_1338,N_1141,N_1155);
and U1339 (N_1339,N_1129,N_1109);
and U1340 (N_1340,In_1406,N_1166);
xnor U1341 (N_1341,N_1198,N_890);
xor U1342 (N_1342,N_1014,N_1232);
and U1343 (N_1343,N_1099,N_1222);
nand U1344 (N_1344,N_858,N_1187);
or U1345 (N_1345,N_1079,In_808);
nor U1346 (N_1346,N_214,N_1195);
xnor U1347 (N_1347,N_838,N_1082);
nand U1348 (N_1348,N_1144,N_1138);
or U1349 (N_1349,N_1161,N_988);
xnor U1350 (N_1350,N_1234,N_983);
nand U1351 (N_1351,N_871,N_1209);
and U1352 (N_1352,In_1356,N_1149);
xor U1353 (N_1353,N_1034,N_1188);
xnor U1354 (N_1354,N_427,N_1214);
xnor U1355 (N_1355,N_1061,N_522);
xnor U1356 (N_1356,N_897,N_1125);
nor U1357 (N_1357,N_1248,In_259);
nor U1358 (N_1358,N_1057,N_1200);
and U1359 (N_1359,In_356,N_1111);
nor U1360 (N_1360,N_1218,N_1241);
and U1361 (N_1361,In_761,N_1115);
nor U1362 (N_1362,N_559,N_1133);
xor U1363 (N_1363,N_910,N_1174);
xnor U1364 (N_1364,N_446,In_839);
and U1365 (N_1365,N_1178,N_1145);
and U1366 (N_1366,N_1139,N_1147);
nor U1367 (N_1367,N_1240,N_1245);
nand U1368 (N_1368,N_1181,N_387);
and U1369 (N_1369,N_1021,N_794);
nor U1370 (N_1370,N_901,N_1239);
xnor U1371 (N_1371,N_849,N_1064);
nor U1372 (N_1372,N_1118,N_1229);
and U1373 (N_1373,N_307,N_1186);
nand U1374 (N_1374,N_1196,N_1201);
nand U1375 (N_1375,N_1259,N_1294);
xnor U1376 (N_1376,N_1264,N_1355);
and U1377 (N_1377,N_1362,N_1344);
nand U1378 (N_1378,N_1267,N_1290);
or U1379 (N_1379,N_1351,N_1266);
and U1380 (N_1380,N_1357,N_1360);
xnor U1381 (N_1381,N_1313,N_1275);
xnor U1382 (N_1382,N_1345,N_1280);
and U1383 (N_1383,N_1302,N_1330);
or U1384 (N_1384,N_1347,N_1318);
nor U1385 (N_1385,N_1338,N_1333);
or U1386 (N_1386,N_1328,N_1308);
nand U1387 (N_1387,N_1321,N_1301);
or U1388 (N_1388,N_1281,N_1331);
xnor U1389 (N_1389,N_1370,N_1352);
nor U1390 (N_1390,N_1288,N_1285);
nor U1391 (N_1391,N_1373,N_1329);
nand U1392 (N_1392,N_1269,N_1295);
nand U1393 (N_1393,N_1340,N_1276);
and U1394 (N_1394,N_1303,N_1256);
xnor U1395 (N_1395,N_1282,N_1304);
or U1396 (N_1396,N_1271,N_1374);
nand U1397 (N_1397,N_1265,N_1358);
xnor U1398 (N_1398,N_1272,N_1372);
nand U1399 (N_1399,N_1332,N_1293);
nor U1400 (N_1400,N_1298,N_1371);
nand U1401 (N_1401,N_1268,N_1315);
nor U1402 (N_1402,N_1367,N_1322);
and U1403 (N_1403,N_1343,N_1310);
xnor U1404 (N_1404,N_1337,N_1324);
nor U1405 (N_1405,N_1314,N_1289);
or U1406 (N_1406,N_1291,N_1353);
nor U1407 (N_1407,N_1277,N_1356);
or U1408 (N_1408,N_1251,N_1260);
nor U1409 (N_1409,N_1258,N_1263);
and U1410 (N_1410,N_1316,N_1317);
xor U1411 (N_1411,N_1312,N_1300);
and U1412 (N_1412,N_1364,N_1336);
nor U1413 (N_1413,N_1366,N_1261);
and U1414 (N_1414,N_1346,N_1365);
or U1415 (N_1415,N_1309,N_1334);
and U1416 (N_1416,N_1319,N_1255);
and U1417 (N_1417,N_1305,N_1320);
and U1418 (N_1418,N_1297,N_1254);
and U1419 (N_1419,N_1286,N_1299);
nor U1420 (N_1420,N_1341,N_1363);
xnor U1421 (N_1421,N_1369,N_1349);
nor U1422 (N_1422,N_1274,N_1250);
or U1423 (N_1423,N_1287,N_1253);
xnor U1424 (N_1424,N_1279,N_1252);
and U1425 (N_1425,N_1311,N_1342);
or U1426 (N_1426,N_1283,N_1350);
nor U1427 (N_1427,N_1284,N_1307);
xnor U1428 (N_1428,N_1327,N_1323);
nand U1429 (N_1429,N_1359,N_1273);
nor U1430 (N_1430,N_1278,N_1348);
nand U1431 (N_1431,N_1368,N_1306);
nor U1432 (N_1432,N_1354,N_1325);
nand U1433 (N_1433,N_1257,N_1335);
nand U1434 (N_1434,N_1339,N_1361);
or U1435 (N_1435,N_1292,N_1326);
nor U1436 (N_1436,N_1270,N_1296);
nor U1437 (N_1437,N_1262,N_1313);
nor U1438 (N_1438,N_1282,N_1353);
nand U1439 (N_1439,N_1263,N_1272);
or U1440 (N_1440,N_1255,N_1258);
xor U1441 (N_1441,N_1279,N_1288);
nor U1442 (N_1442,N_1271,N_1351);
xor U1443 (N_1443,N_1304,N_1284);
nor U1444 (N_1444,N_1273,N_1269);
and U1445 (N_1445,N_1310,N_1362);
xnor U1446 (N_1446,N_1271,N_1310);
or U1447 (N_1447,N_1307,N_1306);
and U1448 (N_1448,N_1372,N_1276);
or U1449 (N_1449,N_1349,N_1328);
xnor U1450 (N_1450,N_1363,N_1331);
nor U1451 (N_1451,N_1355,N_1286);
or U1452 (N_1452,N_1255,N_1256);
nand U1453 (N_1453,N_1262,N_1285);
or U1454 (N_1454,N_1269,N_1293);
and U1455 (N_1455,N_1334,N_1326);
nand U1456 (N_1456,N_1339,N_1289);
xnor U1457 (N_1457,N_1269,N_1274);
or U1458 (N_1458,N_1362,N_1321);
nand U1459 (N_1459,N_1286,N_1268);
and U1460 (N_1460,N_1357,N_1372);
nor U1461 (N_1461,N_1332,N_1331);
and U1462 (N_1462,N_1280,N_1255);
or U1463 (N_1463,N_1265,N_1373);
or U1464 (N_1464,N_1308,N_1371);
and U1465 (N_1465,N_1339,N_1332);
or U1466 (N_1466,N_1344,N_1364);
or U1467 (N_1467,N_1342,N_1266);
xor U1468 (N_1468,N_1356,N_1350);
xor U1469 (N_1469,N_1261,N_1314);
or U1470 (N_1470,N_1320,N_1297);
and U1471 (N_1471,N_1319,N_1364);
or U1472 (N_1472,N_1307,N_1274);
xnor U1473 (N_1473,N_1350,N_1323);
or U1474 (N_1474,N_1332,N_1309);
or U1475 (N_1475,N_1334,N_1343);
xor U1476 (N_1476,N_1341,N_1267);
or U1477 (N_1477,N_1361,N_1321);
nor U1478 (N_1478,N_1347,N_1339);
xor U1479 (N_1479,N_1265,N_1352);
or U1480 (N_1480,N_1328,N_1323);
xor U1481 (N_1481,N_1348,N_1259);
and U1482 (N_1482,N_1278,N_1343);
xnor U1483 (N_1483,N_1269,N_1252);
nand U1484 (N_1484,N_1252,N_1328);
nand U1485 (N_1485,N_1340,N_1362);
or U1486 (N_1486,N_1259,N_1313);
or U1487 (N_1487,N_1351,N_1253);
and U1488 (N_1488,N_1326,N_1267);
nand U1489 (N_1489,N_1305,N_1323);
and U1490 (N_1490,N_1282,N_1256);
or U1491 (N_1491,N_1282,N_1306);
nand U1492 (N_1492,N_1278,N_1354);
and U1493 (N_1493,N_1287,N_1332);
and U1494 (N_1494,N_1327,N_1321);
and U1495 (N_1495,N_1293,N_1372);
xor U1496 (N_1496,N_1275,N_1342);
or U1497 (N_1497,N_1281,N_1362);
nand U1498 (N_1498,N_1325,N_1346);
or U1499 (N_1499,N_1311,N_1363);
xnor U1500 (N_1500,N_1491,N_1421);
xor U1501 (N_1501,N_1410,N_1489);
xor U1502 (N_1502,N_1446,N_1443);
nor U1503 (N_1503,N_1469,N_1401);
and U1504 (N_1504,N_1487,N_1404);
or U1505 (N_1505,N_1399,N_1479);
or U1506 (N_1506,N_1467,N_1492);
and U1507 (N_1507,N_1383,N_1495);
and U1508 (N_1508,N_1415,N_1440);
xor U1509 (N_1509,N_1429,N_1473);
xor U1510 (N_1510,N_1384,N_1456);
nor U1511 (N_1511,N_1454,N_1437);
nand U1512 (N_1512,N_1427,N_1442);
nor U1513 (N_1513,N_1388,N_1402);
or U1514 (N_1514,N_1475,N_1375);
nor U1515 (N_1515,N_1400,N_1478);
xor U1516 (N_1516,N_1379,N_1385);
or U1517 (N_1517,N_1482,N_1411);
nor U1518 (N_1518,N_1420,N_1460);
or U1519 (N_1519,N_1463,N_1445);
and U1520 (N_1520,N_1430,N_1409);
xor U1521 (N_1521,N_1441,N_1457);
or U1522 (N_1522,N_1408,N_1406);
and U1523 (N_1523,N_1398,N_1455);
xnor U1524 (N_1524,N_1439,N_1381);
nand U1525 (N_1525,N_1493,N_1432);
nor U1526 (N_1526,N_1458,N_1431);
nor U1527 (N_1527,N_1497,N_1481);
and U1528 (N_1528,N_1451,N_1403);
nor U1529 (N_1529,N_1419,N_1447);
nor U1530 (N_1530,N_1459,N_1477);
nor U1531 (N_1531,N_1396,N_1407);
and U1532 (N_1532,N_1393,N_1471);
xor U1533 (N_1533,N_1470,N_1425);
nor U1534 (N_1534,N_1412,N_1397);
nor U1535 (N_1535,N_1483,N_1428);
and U1536 (N_1536,N_1480,N_1418);
nor U1537 (N_1537,N_1448,N_1486);
xnor U1538 (N_1538,N_1394,N_1426);
xnor U1539 (N_1539,N_1474,N_1416);
and U1540 (N_1540,N_1387,N_1434);
nor U1541 (N_1541,N_1450,N_1449);
nand U1542 (N_1542,N_1378,N_1464);
or U1543 (N_1543,N_1436,N_1452);
and U1544 (N_1544,N_1466,N_1424);
or U1545 (N_1545,N_1391,N_1468);
nor U1546 (N_1546,N_1392,N_1433);
xor U1547 (N_1547,N_1476,N_1395);
xnor U1548 (N_1548,N_1438,N_1405);
nor U1549 (N_1549,N_1444,N_1417);
nand U1550 (N_1550,N_1496,N_1461);
or U1551 (N_1551,N_1422,N_1465);
or U1552 (N_1552,N_1462,N_1484);
xor U1553 (N_1553,N_1453,N_1413);
nand U1554 (N_1554,N_1376,N_1472);
nand U1555 (N_1555,N_1380,N_1435);
xor U1556 (N_1556,N_1488,N_1423);
or U1557 (N_1557,N_1498,N_1389);
and U1558 (N_1558,N_1485,N_1494);
nor U1559 (N_1559,N_1382,N_1377);
xnor U1560 (N_1560,N_1414,N_1499);
nor U1561 (N_1561,N_1386,N_1390);
or U1562 (N_1562,N_1490,N_1387);
nor U1563 (N_1563,N_1410,N_1449);
and U1564 (N_1564,N_1393,N_1406);
and U1565 (N_1565,N_1457,N_1485);
or U1566 (N_1566,N_1397,N_1464);
nand U1567 (N_1567,N_1398,N_1410);
nand U1568 (N_1568,N_1476,N_1473);
or U1569 (N_1569,N_1449,N_1483);
or U1570 (N_1570,N_1436,N_1433);
or U1571 (N_1571,N_1392,N_1455);
nor U1572 (N_1572,N_1411,N_1445);
nand U1573 (N_1573,N_1496,N_1441);
or U1574 (N_1574,N_1440,N_1389);
and U1575 (N_1575,N_1402,N_1417);
and U1576 (N_1576,N_1431,N_1463);
and U1577 (N_1577,N_1423,N_1418);
nand U1578 (N_1578,N_1480,N_1452);
and U1579 (N_1579,N_1434,N_1495);
and U1580 (N_1580,N_1412,N_1459);
or U1581 (N_1581,N_1446,N_1494);
xor U1582 (N_1582,N_1440,N_1437);
or U1583 (N_1583,N_1406,N_1454);
and U1584 (N_1584,N_1394,N_1437);
and U1585 (N_1585,N_1410,N_1379);
and U1586 (N_1586,N_1445,N_1443);
nor U1587 (N_1587,N_1394,N_1398);
nand U1588 (N_1588,N_1419,N_1388);
nor U1589 (N_1589,N_1483,N_1386);
xor U1590 (N_1590,N_1411,N_1497);
or U1591 (N_1591,N_1491,N_1470);
nor U1592 (N_1592,N_1416,N_1451);
or U1593 (N_1593,N_1434,N_1400);
and U1594 (N_1594,N_1450,N_1391);
nor U1595 (N_1595,N_1399,N_1411);
and U1596 (N_1596,N_1434,N_1446);
nor U1597 (N_1597,N_1490,N_1401);
and U1598 (N_1598,N_1392,N_1380);
nor U1599 (N_1599,N_1492,N_1440);
nor U1600 (N_1600,N_1499,N_1417);
xor U1601 (N_1601,N_1474,N_1475);
nor U1602 (N_1602,N_1482,N_1393);
nor U1603 (N_1603,N_1478,N_1453);
and U1604 (N_1604,N_1467,N_1406);
and U1605 (N_1605,N_1470,N_1434);
nand U1606 (N_1606,N_1475,N_1455);
nand U1607 (N_1607,N_1380,N_1385);
or U1608 (N_1608,N_1469,N_1383);
and U1609 (N_1609,N_1387,N_1421);
nand U1610 (N_1610,N_1409,N_1437);
and U1611 (N_1611,N_1459,N_1476);
nand U1612 (N_1612,N_1434,N_1432);
nand U1613 (N_1613,N_1462,N_1447);
nand U1614 (N_1614,N_1445,N_1419);
or U1615 (N_1615,N_1440,N_1412);
and U1616 (N_1616,N_1472,N_1466);
xor U1617 (N_1617,N_1487,N_1433);
xor U1618 (N_1618,N_1425,N_1381);
nor U1619 (N_1619,N_1378,N_1454);
nor U1620 (N_1620,N_1475,N_1477);
or U1621 (N_1621,N_1388,N_1394);
or U1622 (N_1622,N_1495,N_1419);
nand U1623 (N_1623,N_1496,N_1397);
xor U1624 (N_1624,N_1465,N_1404);
nand U1625 (N_1625,N_1554,N_1578);
and U1626 (N_1626,N_1504,N_1617);
xor U1627 (N_1627,N_1535,N_1547);
or U1628 (N_1628,N_1569,N_1591);
and U1629 (N_1629,N_1531,N_1581);
and U1630 (N_1630,N_1584,N_1603);
nand U1631 (N_1631,N_1563,N_1524);
or U1632 (N_1632,N_1506,N_1602);
nand U1633 (N_1633,N_1611,N_1608);
and U1634 (N_1634,N_1503,N_1588);
nor U1635 (N_1635,N_1577,N_1513);
nand U1636 (N_1636,N_1568,N_1533);
or U1637 (N_1637,N_1622,N_1509);
nor U1638 (N_1638,N_1559,N_1580);
nor U1639 (N_1639,N_1544,N_1539);
xnor U1640 (N_1640,N_1556,N_1623);
or U1641 (N_1641,N_1620,N_1530);
and U1642 (N_1642,N_1598,N_1564);
or U1643 (N_1643,N_1618,N_1561);
xnor U1644 (N_1644,N_1502,N_1565);
and U1645 (N_1645,N_1587,N_1605);
nor U1646 (N_1646,N_1551,N_1516);
xor U1647 (N_1647,N_1606,N_1546);
nand U1648 (N_1648,N_1548,N_1528);
and U1649 (N_1649,N_1553,N_1566);
or U1650 (N_1650,N_1610,N_1537);
nor U1651 (N_1651,N_1518,N_1596);
and U1652 (N_1652,N_1519,N_1555);
xnor U1653 (N_1653,N_1592,N_1624);
and U1654 (N_1654,N_1512,N_1576);
nand U1655 (N_1655,N_1579,N_1501);
or U1656 (N_1656,N_1514,N_1545);
or U1657 (N_1657,N_1607,N_1593);
xor U1658 (N_1658,N_1604,N_1590);
or U1659 (N_1659,N_1510,N_1525);
nor U1660 (N_1660,N_1599,N_1538);
or U1661 (N_1661,N_1595,N_1558);
or U1662 (N_1662,N_1574,N_1541);
nor U1663 (N_1663,N_1532,N_1562);
or U1664 (N_1664,N_1540,N_1619);
xnor U1665 (N_1665,N_1505,N_1621);
or U1666 (N_1666,N_1517,N_1575);
nand U1667 (N_1667,N_1614,N_1511);
xnor U1668 (N_1668,N_1589,N_1612);
nand U1669 (N_1669,N_1560,N_1582);
nor U1670 (N_1670,N_1542,N_1567);
nand U1671 (N_1671,N_1534,N_1583);
and U1672 (N_1672,N_1529,N_1520);
and U1673 (N_1673,N_1571,N_1601);
nand U1674 (N_1674,N_1616,N_1515);
xnor U1675 (N_1675,N_1549,N_1597);
and U1676 (N_1676,N_1500,N_1552);
xor U1677 (N_1677,N_1613,N_1573);
nand U1678 (N_1678,N_1523,N_1609);
xor U1679 (N_1679,N_1550,N_1615);
or U1680 (N_1680,N_1527,N_1572);
or U1681 (N_1681,N_1570,N_1508);
and U1682 (N_1682,N_1521,N_1585);
xor U1683 (N_1683,N_1522,N_1536);
nand U1684 (N_1684,N_1543,N_1557);
nor U1685 (N_1685,N_1600,N_1586);
xor U1686 (N_1686,N_1526,N_1594);
and U1687 (N_1687,N_1507,N_1599);
or U1688 (N_1688,N_1512,N_1579);
nand U1689 (N_1689,N_1552,N_1594);
nand U1690 (N_1690,N_1556,N_1512);
nor U1691 (N_1691,N_1545,N_1524);
or U1692 (N_1692,N_1538,N_1511);
xor U1693 (N_1693,N_1522,N_1582);
and U1694 (N_1694,N_1587,N_1532);
and U1695 (N_1695,N_1516,N_1589);
xor U1696 (N_1696,N_1526,N_1565);
nor U1697 (N_1697,N_1570,N_1597);
nand U1698 (N_1698,N_1530,N_1541);
and U1699 (N_1699,N_1504,N_1545);
xor U1700 (N_1700,N_1535,N_1587);
xor U1701 (N_1701,N_1528,N_1514);
nand U1702 (N_1702,N_1524,N_1579);
xnor U1703 (N_1703,N_1537,N_1528);
nand U1704 (N_1704,N_1501,N_1573);
xor U1705 (N_1705,N_1593,N_1547);
or U1706 (N_1706,N_1526,N_1570);
and U1707 (N_1707,N_1502,N_1563);
or U1708 (N_1708,N_1514,N_1589);
xor U1709 (N_1709,N_1575,N_1534);
nor U1710 (N_1710,N_1596,N_1505);
nand U1711 (N_1711,N_1572,N_1560);
xor U1712 (N_1712,N_1534,N_1558);
and U1713 (N_1713,N_1564,N_1568);
nor U1714 (N_1714,N_1600,N_1546);
nand U1715 (N_1715,N_1584,N_1545);
xor U1716 (N_1716,N_1617,N_1602);
xnor U1717 (N_1717,N_1539,N_1576);
nand U1718 (N_1718,N_1512,N_1594);
nand U1719 (N_1719,N_1543,N_1550);
nand U1720 (N_1720,N_1564,N_1541);
xor U1721 (N_1721,N_1617,N_1606);
nor U1722 (N_1722,N_1594,N_1569);
xor U1723 (N_1723,N_1624,N_1562);
nand U1724 (N_1724,N_1575,N_1617);
nor U1725 (N_1725,N_1601,N_1591);
nor U1726 (N_1726,N_1610,N_1535);
nor U1727 (N_1727,N_1518,N_1607);
and U1728 (N_1728,N_1566,N_1605);
or U1729 (N_1729,N_1505,N_1510);
nor U1730 (N_1730,N_1599,N_1580);
or U1731 (N_1731,N_1562,N_1525);
and U1732 (N_1732,N_1507,N_1601);
nand U1733 (N_1733,N_1564,N_1561);
and U1734 (N_1734,N_1533,N_1543);
nand U1735 (N_1735,N_1506,N_1509);
xnor U1736 (N_1736,N_1565,N_1539);
nand U1737 (N_1737,N_1542,N_1516);
and U1738 (N_1738,N_1562,N_1583);
nor U1739 (N_1739,N_1621,N_1532);
nand U1740 (N_1740,N_1559,N_1516);
xnor U1741 (N_1741,N_1593,N_1516);
and U1742 (N_1742,N_1540,N_1549);
xor U1743 (N_1743,N_1623,N_1564);
nor U1744 (N_1744,N_1539,N_1613);
nand U1745 (N_1745,N_1603,N_1541);
xnor U1746 (N_1746,N_1561,N_1560);
nand U1747 (N_1747,N_1590,N_1567);
nor U1748 (N_1748,N_1622,N_1596);
and U1749 (N_1749,N_1572,N_1564);
nand U1750 (N_1750,N_1712,N_1643);
nor U1751 (N_1751,N_1695,N_1665);
or U1752 (N_1752,N_1626,N_1700);
and U1753 (N_1753,N_1717,N_1719);
nor U1754 (N_1754,N_1732,N_1692);
nor U1755 (N_1755,N_1635,N_1646);
nor U1756 (N_1756,N_1741,N_1640);
xor U1757 (N_1757,N_1702,N_1682);
and U1758 (N_1758,N_1689,N_1644);
nor U1759 (N_1759,N_1658,N_1723);
and U1760 (N_1760,N_1722,N_1649);
xnor U1761 (N_1761,N_1735,N_1704);
and U1762 (N_1762,N_1709,N_1694);
nor U1763 (N_1763,N_1655,N_1663);
nor U1764 (N_1764,N_1730,N_1714);
nor U1765 (N_1765,N_1678,N_1742);
and U1766 (N_1766,N_1664,N_1639);
nor U1767 (N_1767,N_1657,N_1671);
nor U1768 (N_1768,N_1696,N_1638);
nand U1769 (N_1769,N_1660,N_1749);
or U1770 (N_1770,N_1744,N_1740);
nand U1771 (N_1771,N_1701,N_1691);
xor U1772 (N_1772,N_1641,N_1669);
nor U1773 (N_1773,N_1720,N_1668);
and U1774 (N_1774,N_1637,N_1666);
xnor U1775 (N_1775,N_1676,N_1710);
xnor U1776 (N_1776,N_1737,N_1650);
nand U1777 (N_1777,N_1630,N_1708);
nand U1778 (N_1778,N_1656,N_1667);
and U1779 (N_1779,N_1631,N_1721);
or U1780 (N_1780,N_1718,N_1738);
nor U1781 (N_1781,N_1705,N_1679);
nand U1782 (N_1782,N_1627,N_1725);
and U1783 (N_1783,N_1707,N_1745);
xor U1784 (N_1784,N_1683,N_1687);
nor U1785 (N_1785,N_1697,N_1636);
or U1786 (N_1786,N_1728,N_1659);
or U1787 (N_1787,N_1654,N_1681);
nor U1788 (N_1788,N_1706,N_1747);
or U1789 (N_1789,N_1634,N_1647);
xnor U1790 (N_1790,N_1688,N_1693);
nor U1791 (N_1791,N_1727,N_1739);
and U1792 (N_1792,N_1731,N_1715);
nor U1793 (N_1793,N_1677,N_1662);
or U1794 (N_1794,N_1686,N_1661);
and U1795 (N_1795,N_1633,N_1724);
and U1796 (N_1796,N_1698,N_1743);
nand U1797 (N_1797,N_1653,N_1680);
and U1798 (N_1798,N_1711,N_1748);
nor U1799 (N_1799,N_1699,N_1674);
or U1800 (N_1800,N_1628,N_1726);
xor U1801 (N_1801,N_1734,N_1713);
and U1802 (N_1802,N_1673,N_1716);
xnor U1803 (N_1803,N_1703,N_1690);
nand U1804 (N_1804,N_1651,N_1685);
xnor U1805 (N_1805,N_1675,N_1746);
nand U1806 (N_1806,N_1733,N_1632);
and U1807 (N_1807,N_1648,N_1670);
and U1808 (N_1808,N_1642,N_1684);
or U1809 (N_1809,N_1672,N_1629);
or U1810 (N_1810,N_1645,N_1736);
and U1811 (N_1811,N_1652,N_1625);
and U1812 (N_1812,N_1729,N_1639);
nor U1813 (N_1813,N_1701,N_1678);
and U1814 (N_1814,N_1628,N_1670);
nor U1815 (N_1815,N_1749,N_1646);
and U1816 (N_1816,N_1643,N_1656);
nand U1817 (N_1817,N_1666,N_1655);
nand U1818 (N_1818,N_1722,N_1642);
and U1819 (N_1819,N_1728,N_1747);
nand U1820 (N_1820,N_1655,N_1695);
xor U1821 (N_1821,N_1691,N_1747);
nand U1822 (N_1822,N_1667,N_1735);
nand U1823 (N_1823,N_1665,N_1700);
xor U1824 (N_1824,N_1726,N_1709);
nand U1825 (N_1825,N_1733,N_1730);
xnor U1826 (N_1826,N_1666,N_1745);
and U1827 (N_1827,N_1749,N_1642);
xnor U1828 (N_1828,N_1705,N_1739);
xor U1829 (N_1829,N_1744,N_1641);
or U1830 (N_1830,N_1629,N_1707);
nor U1831 (N_1831,N_1645,N_1701);
nand U1832 (N_1832,N_1655,N_1635);
and U1833 (N_1833,N_1713,N_1735);
nand U1834 (N_1834,N_1668,N_1739);
nand U1835 (N_1835,N_1680,N_1677);
nand U1836 (N_1836,N_1655,N_1722);
or U1837 (N_1837,N_1666,N_1747);
xor U1838 (N_1838,N_1647,N_1667);
nand U1839 (N_1839,N_1677,N_1748);
nand U1840 (N_1840,N_1729,N_1682);
nand U1841 (N_1841,N_1730,N_1647);
and U1842 (N_1842,N_1652,N_1649);
or U1843 (N_1843,N_1694,N_1665);
nand U1844 (N_1844,N_1627,N_1668);
nand U1845 (N_1845,N_1652,N_1731);
or U1846 (N_1846,N_1681,N_1685);
and U1847 (N_1847,N_1701,N_1685);
or U1848 (N_1848,N_1639,N_1703);
xor U1849 (N_1849,N_1667,N_1671);
nor U1850 (N_1850,N_1660,N_1695);
and U1851 (N_1851,N_1694,N_1669);
and U1852 (N_1852,N_1638,N_1652);
nor U1853 (N_1853,N_1727,N_1699);
and U1854 (N_1854,N_1744,N_1666);
or U1855 (N_1855,N_1708,N_1719);
and U1856 (N_1856,N_1647,N_1724);
or U1857 (N_1857,N_1679,N_1689);
xnor U1858 (N_1858,N_1722,N_1667);
xnor U1859 (N_1859,N_1719,N_1727);
nand U1860 (N_1860,N_1661,N_1650);
and U1861 (N_1861,N_1646,N_1702);
and U1862 (N_1862,N_1647,N_1686);
and U1863 (N_1863,N_1633,N_1653);
or U1864 (N_1864,N_1680,N_1648);
nor U1865 (N_1865,N_1721,N_1691);
nor U1866 (N_1866,N_1745,N_1677);
nor U1867 (N_1867,N_1692,N_1748);
or U1868 (N_1868,N_1643,N_1650);
or U1869 (N_1869,N_1724,N_1714);
or U1870 (N_1870,N_1743,N_1701);
nor U1871 (N_1871,N_1730,N_1685);
nor U1872 (N_1872,N_1654,N_1721);
or U1873 (N_1873,N_1737,N_1677);
nor U1874 (N_1874,N_1690,N_1746);
nand U1875 (N_1875,N_1787,N_1806);
and U1876 (N_1876,N_1757,N_1813);
nor U1877 (N_1877,N_1854,N_1873);
nand U1878 (N_1878,N_1839,N_1825);
xor U1879 (N_1879,N_1822,N_1869);
xnor U1880 (N_1880,N_1785,N_1815);
or U1881 (N_1881,N_1796,N_1857);
xor U1882 (N_1882,N_1820,N_1858);
or U1883 (N_1883,N_1819,N_1847);
or U1884 (N_1884,N_1760,N_1794);
nor U1885 (N_1885,N_1814,N_1784);
xnor U1886 (N_1886,N_1795,N_1752);
or U1887 (N_1887,N_1846,N_1792);
and U1888 (N_1888,N_1801,N_1810);
xnor U1889 (N_1889,N_1832,N_1790);
xnor U1890 (N_1890,N_1758,N_1824);
nor U1891 (N_1891,N_1826,N_1862);
or U1892 (N_1892,N_1840,N_1753);
nor U1893 (N_1893,N_1856,N_1834);
and U1894 (N_1894,N_1838,N_1770);
or U1895 (N_1895,N_1771,N_1833);
nor U1896 (N_1896,N_1804,N_1761);
or U1897 (N_1897,N_1831,N_1789);
nor U1898 (N_1898,N_1864,N_1837);
and U1899 (N_1899,N_1773,N_1871);
nor U1900 (N_1900,N_1821,N_1849);
or U1901 (N_1901,N_1860,N_1774);
xor U1902 (N_1902,N_1829,N_1827);
xnor U1903 (N_1903,N_1797,N_1768);
and U1904 (N_1904,N_1765,N_1764);
and U1905 (N_1905,N_1816,N_1872);
and U1906 (N_1906,N_1865,N_1798);
nor U1907 (N_1907,N_1852,N_1781);
and U1908 (N_1908,N_1800,N_1868);
or U1909 (N_1909,N_1867,N_1788);
nand U1910 (N_1910,N_1750,N_1786);
and U1911 (N_1911,N_1755,N_1807);
nor U1912 (N_1912,N_1855,N_1843);
or U1913 (N_1913,N_1778,N_1772);
xor U1914 (N_1914,N_1805,N_1802);
and U1915 (N_1915,N_1866,N_1841);
nor U1916 (N_1916,N_1776,N_1799);
or U1917 (N_1917,N_1793,N_1835);
nand U1918 (N_1918,N_1779,N_1751);
nand U1919 (N_1919,N_1769,N_1828);
xnor U1920 (N_1920,N_1818,N_1851);
or U1921 (N_1921,N_1874,N_1842);
nor U1922 (N_1922,N_1861,N_1782);
nand U1923 (N_1923,N_1766,N_1853);
xor U1924 (N_1924,N_1754,N_1777);
or U1925 (N_1925,N_1863,N_1850);
nor U1926 (N_1926,N_1791,N_1836);
or U1927 (N_1927,N_1830,N_1811);
or U1928 (N_1928,N_1763,N_1775);
and U1929 (N_1929,N_1817,N_1808);
nand U1930 (N_1930,N_1756,N_1848);
and U1931 (N_1931,N_1870,N_1759);
and U1932 (N_1932,N_1803,N_1812);
and U1933 (N_1933,N_1809,N_1767);
and U1934 (N_1934,N_1762,N_1780);
xor U1935 (N_1935,N_1859,N_1783);
nand U1936 (N_1936,N_1823,N_1845);
and U1937 (N_1937,N_1844,N_1810);
and U1938 (N_1938,N_1791,N_1855);
nand U1939 (N_1939,N_1814,N_1825);
nor U1940 (N_1940,N_1751,N_1778);
nor U1941 (N_1941,N_1852,N_1794);
nor U1942 (N_1942,N_1779,N_1770);
and U1943 (N_1943,N_1802,N_1781);
nand U1944 (N_1944,N_1855,N_1831);
or U1945 (N_1945,N_1820,N_1868);
xnor U1946 (N_1946,N_1816,N_1869);
nor U1947 (N_1947,N_1825,N_1841);
nor U1948 (N_1948,N_1812,N_1827);
or U1949 (N_1949,N_1843,N_1849);
or U1950 (N_1950,N_1839,N_1759);
nor U1951 (N_1951,N_1767,N_1754);
and U1952 (N_1952,N_1783,N_1845);
nand U1953 (N_1953,N_1820,N_1787);
or U1954 (N_1954,N_1782,N_1804);
xnor U1955 (N_1955,N_1822,N_1824);
xnor U1956 (N_1956,N_1810,N_1840);
nand U1957 (N_1957,N_1827,N_1861);
nand U1958 (N_1958,N_1782,N_1783);
xor U1959 (N_1959,N_1791,N_1832);
nor U1960 (N_1960,N_1830,N_1765);
or U1961 (N_1961,N_1853,N_1838);
nor U1962 (N_1962,N_1761,N_1862);
xnor U1963 (N_1963,N_1831,N_1788);
nand U1964 (N_1964,N_1789,N_1856);
xnor U1965 (N_1965,N_1826,N_1856);
xnor U1966 (N_1966,N_1750,N_1780);
nand U1967 (N_1967,N_1864,N_1846);
nand U1968 (N_1968,N_1817,N_1843);
nor U1969 (N_1969,N_1828,N_1801);
or U1970 (N_1970,N_1856,N_1765);
and U1971 (N_1971,N_1756,N_1801);
nand U1972 (N_1972,N_1814,N_1777);
and U1973 (N_1973,N_1831,N_1838);
xnor U1974 (N_1974,N_1856,N_1788);
or U1975 (N_1975,N_1789,N_1834);
and U1976 (N_1976,N_1790,N_1786);
or U1977 (N_1977,N_1780,N_1776);
and U1978 (N_1978,N_1838,N_1797);
nand U1979 (N_1979,N_1847,N_1868);
or U1980 (N_1980,N_1861,N_1821);
and U1981 (N_1981,N_1798,N_1824);
and U1982 (N_1982,N_1812,N_1799);
or U1983 (N_1983,N_1789,N_1771);
nor U1984 (N_1984,N_1819,N_1827);
or U1985 (N_1985,N_1797,N_1864);
nor U1986 (N_1986,N_1847,N_1778);
and U1987 (N_1987,N_1825,N_1794);
nand U1988 (N_1988,N_1863,N_1865);
and U1989 (N_1989,N_1761,N_1777);
or U1990 (N_1990,N_1758,N_1827);
nand U1991 (N_1991,N_1854,N_1784);
nand U1992 (N_1992,N_1838,N_1870);
or U1993 (N_1993,N_1804,N_1857);
or U1994 (N_1994,N_1801,N_1826);
nor U1995 (N_1995,N_1775,N_1858);
nor U1996 (N_1996,N_1835,N_1758);
nand U1997 (N_1997,N_1790,N_1848);
xor U1998 (N_1998,N_1808,N_1766);
nand U1999 (N_1999,N_1755,N_1810);
nand U2000 (N_2000,N_1875,N_1897);
nand U2001 (N_2001,N_1939,N_1941);
or U2002 (N_2002,N_1968,N_1986);
xor U2003 (N_2003,N_1972,N_1924);
nand U2004 (N_2004,N_1894,N_1971);
xnor U2005 (N_2005,N_1982,N_1948);
and U2006 (N_2006,N_1884,N_1906);
or U2007 (N_2007,N_1983,N_1947);
and U2008 (N_2008,N_1997,N_1996);
nor U2009 (N_2009,N_1902,N_1919);
and U2010 (N_2010,N_1891,N_1886);
and U2011 (N_2011,N_1967,N_1883);
and U2012 (N_2012,N_1989,N_1993);
nand U2013 (N_2013,N_1914,N_1908);
and U2014 (N_2014,N_1969,N_1879);
or U2015 (N_2015,N_1999,N_1928);
xor U2016 (N_2016,N_1961,N_1994);
xnor U2017 (N_2017,N_1905,N_1929);
nor U2018 (N_2018,N_1926,N_1974);
nand U2019 (N_2019,N_1899,N_1901);
and U2020 (N_2020,N_1950,N_1876);
and U2021 (N_2021,N_1937,N_1930);
xnor U2022 (N_2022,N_1903,N_1964);
nor U2023 (N_2023,N_1949,N_1935);
xor U2024 (N_2024,N_1957,N_1916);
nand U2025 (N_2025,N_1880,N_1960);
or U2026 (N_2026,N_1888,N_1915);
or U2027 (N_2027,N_1940,N_1920);
and U2028 (N_2028,N_1878,N_1885);
and U2029 (N_2029,N_1966,N_1979);
nor U2030 (N_2030,N_1944,N_1893);
and U2031 (N_2031,N_1907,N_1953);
nand U2032 (N_2032,N_1936,N_1896);
xor U2033 (N_2033,N_1921,N_1975);
or U2034 (N_2034,N_1912,N_1934);
or U2035 (N_2035,N_1922,N_1904);
xor U2036 (N_2036,N_1900,N_1887);
nor U2037 (N_2037,N_1987,N_1898);
or U2038 (N_2038,N_1933,N_1895);
nor U2039 (N_2039,N_1892,N_1956);
xnor U2040 (N_2040,N_1952,N_1951);
nand U2041 (N_2041,N_1977,N_1925);
nor U2042 (N_2042,N_1889,N_1965);
nand U2043 (N_2043,N_1909,N_1988);
xnor U2044 (N_2044,N_1973,N_1954);
or U2045 (N_2045,N_1984,N_1923);
xnor U2046 (N_2046,N_1946,N_1998);
or U2047 (N_2047,N_1942,N_1980);
nand U2048 (N_2048,N_1943,N_1945);
and U2049 (N_2049,N_1917,N_1976);
or U2050 (N_2050,N_1963,N_1981);
xor U2051 (N_2051,N_1995,N_1910);
nor U2052 (N_2052,N_1882,N_1992);
xor U2053 (N_2053,N_1970,N_1959);
or U2054 (N_2054,N_1918,N_1927);
nor U2055 (N_2055,N_1931,N_1890);
nand U2056 (N_2056,N_1932,N_1958);
nor U2057 (N_2057,N_1991,N_1962);
or U2058 (N_2058,N_1881,N_1877);
nand U2059 (N_2059,N_1990,N_1911);
nand U2060 (N_2060,N_1985,N_1978);
xor U2061 (N_2061,N_1938,N_1955);
nand U2062 (N_2062,N_1913,N_1952);
and U2063 (N_2063,N_1953,N_1946);
or U2064 (N_2064,N_1964,N_1995);
and U2065 (N_2065,N_1947,N_1877);
xnor U2066 (N_2066,N_1940,N_1954);
xor U2067 (N_2067,N_1916,N_1970);
nor U2068 (N_2068,N_1975,N_1956);
nor U2069 (N_2069,N_1938,N_1995);
nor U2070 (N_2070,N_1994,N_1954);
and U2071 (N_2071,N_1909,N_1912);
nand U2072 (N_2072,N_1955,N_1918);
and U2073 (N_2073,N_1991,N_1905);
nand U2074 (N_2074,N_1999,N_1899);
and U2075 (N_2075,N_1890,N_1976);
nor U2076 (N_2076,N_1974,N_1886);
nor U2077 (N_2077,N_1898,N_1917);
and U2078 (N_2078,N_1922,N_1983);
nand U2079 (N_2079,N_1930,N_1907);
or U2080 (N_2080,N_1978,N_1946);
nor U2081 (N_2081,N_1886,N_1986);
and U2082 (N_2082,N_1949,N_1997);
xnor U2083 (N_2083,N_1884,N_1943);
xnor U2084 (N_2084,N_1885,N_1940);
nand U2085 (N_2085,N_1919,N_1961);
or U2086 (N_2086,N_1996,N_1892);
or U2087 (N_2087,N_1884,N_1928);
nand U2088 (N_2088,N_1928,N_1898);
nor U2089 (N_2089,N_1877,N_1875);
nor U2090 (N_2090,N_1916,N_1950);
and U2091 (N_2091,N_1975,N_1906);
or U2092 (N_2092,N_1986,N_1983);
and U2093 (N_2093,N_1964,N_1943);
and U2094 (N_2094,N_1964,N_1875);
nand U2095 (N_2095,N_1891,N_1898);
xnor U2096 (N_2096,N_1938,N_1943);
nor U2097 (N_2097,N_1894,N_1997);
nand U2098 (N_2098,N_1931,N_1973);
or U2099 (N_2099,N_1892,N_1965);
nor U2100 (N_2100,N_1925,N_1983);
nand U2101 (N_2101,N_1998,N_1982);
and U2102 (N_2102,N_1920,N_1938);
and U2103 (N_2103,N_1895,N_1998);
xor U2104 (N_2104,N_1971,N_1893);
and U2105 (N_2105,N_1915,N_1896);
or U2106 (N_2106,N_1994,N_1908);
and U2107 (N_2107,N_1940,N_1883);
or U2108 (N_2108,N_1943,N_1926);
xnor U2109 (N_2109,N_1963,N_1901);
xnor U2110 (N_2110,N_1983,N_1896);
and U2111 (N_2111,N_1980,N_1924);
and U2112 (N_2112,N_1926,N_1981);
and U2113 (N_2113,N_1902,N_1937);
xor U2114 (N_2114,N_1954,N_1906);
and U2115 (N_2115,N_1882,N_1998);
or U2116 (N_2116,N_1982,N_1955);
or U2117 (N_2117,N_1987,N_1919);
or U2118 (N_2118,N_1901,N_1893);
or U2119 (N_2119,N_1907,N_1914);
xor U2120 (N_2120,N_1951,N_1894);
or U2121 (N_2121,N_1924,N_1888);
and U2122 (N_2122,N_1927,N_1920);
xnor U2123 (N_2123,N_1971,N_1902);
and U2124 (N_2124,N_1959,N_1887);
nand U2125 (N_2125,N_2095,N_2115);
nor U2126 (N_2126,N_2117,N_2004);
or U2127 (N_2127,N_2107,N_2055);
or U2128 (N_2128,N_2069,N_2005);
nand U2129 (N_2129,N_2018,N_2108);
nor U2130 (N_2130,N_2040,N_2087);
nand U2131 (N_2131,N_2081,N_2016);
or U2132 (N_2132,N_2027,N_2021);
nor U2133 (N_2133,N_2078,N_2092);
nor U2134 (N_2134,N_2116,N_2097);
nor U2135 (N_2135,N_2033,N_2028);
and U2136 (N_2136,N_2089,N_2048);
xor U2137 (N_2137,N_2013,N_2091);
nand U2138 (N_2138,N_2110,N_2062);
nand U2139 (N_2139,N_2067,N_2032);
nor U2140 (N_2140,N_2041,N_2059);
xor U2141 (N_2141,N_2010,N_2085);
nor U2142 (N_2142,N_2086,N_2096);
or U2143 (N_2143,N_2104,N_2052);
and U2144 (N_2144,N_2008,N_2009);
nor U2145 (N_2145,N_2049,N_2066);
and U2146 (N_2146,N_2063,N_2060);
or U2147 (N_2147,N_2068,N_2083);
or U2148 (N_2148,N_2042,N_2023);
nor U2149 (N_2149,N_2043,N_2030);
nor U2150 (N_2150,N_2029,N_2058);
xor U2151 (N_2151,N_2102,N_2099);
nor U2152 (N_2152,N_2056,N_2120);
nand U2153 (N_2153,N_2065,N_2047);
nand U2154 (N_2154,N_2017,N_2000);
nor U2155 (N_2155,N_2064,N_2019);
or U2156 (N_2156,N_2031,N_2012);
nor U2157 (N_2157,N_2100,N_2122);
or U2158 (N_2158,N_2118,N_2044);
or U2159 (N_2159,N_2082,N_2103);
xnor U2160 (N_2160,N_2112,N_2074);
xor U2161 (N_2161,N_2070,N_2114);
nor U2162 (N_2162,N_2075,N_2024);
nand U2163 (N_2163,N_2046,N_2079);
and U2164 (N_2164,N_2039,N_2098);
or U2165 (N_2165,N_2057,N_2035);
nor U2166 (N_2166,N_2045,N_2076);
or U2167 (N_2167,N_2088,N_2111);
nor U2168 (N_2168,N_2084,N_2051);
or U2169 (N_2169,N_2037,N_2007);
or U2170 (N_2170,N_2124,N_2123);
nor U2171 (N_2171,N_2080,N_2001);
or U2172 (N_2172,N_2053,N_2003);
nand U2173 (N_2173,N_2093,N_2050);
nand U2174 (N_2174,N_2026,N_2094);
or U2175 (N_2175,N_2101,N_2002);
nand U2176 (N_2176,N_2106,N_2121);
xor U2177 (N_2177,N_2038,N_2054);
nor U2178 (N_2178,N_2022,N_2077);
nor U2179 (N_2179,N_2011,N_2014);
or U2180 (N_2180,N_2015,N_2071);
nand U2181 (N_2181,N_2109,N_2061);
nand U2182 (N_2182,N_2025,N_2113);
nor U2183 (N_2183,N_2006,N_2020);
nor U2184 (N_2184,N_2090,N_2105);
and U2185 (N_2185,N_2034,N_2073);
nand U2186 (N_2186,N_2072,N_2036);
nand U2187 (N_2187,N_2119,N_2061);
nand U2188 (N_2188,N_2122,N_2095);
nor U2189 (N_2189,N_2052,N_2038);
xor U2190 (N_2190,N_2045,N_2017);
and U2191 (N_2191,N_2059,N_2069);
nand U2192 (N_2192,N_2123,N_2031);
xnor U2193 (N_2193,N_2094,N_2109);
and U2194 (N_2194,N_2109,N_2011);
xor U2195 (N_2195,N_2099,N_2053);
xnor U2196 (N_2196,N_2049,N_2074);
nor U2197 (N_2197,N_2034,N_2012);
nand U2198 (N_2198,N_2009,N_2117);
nor U2199 (N_2199,N_2101,N_2079);
nand U2200 (N_2200,N_2090,N_2014);
nor U2201 (N_2201,N_2056,N_2017);
and U2202 (N_2202,N_2032,N_2049);
or U2203 (N_2203,N_2047,N_2058);
nand U2204 (N_2204,N_2043,N_2098);
or U2205 (N_2205,N_2077,N_2083);
xnor U2206 (N_2206,N_2077,N_2102);
nand U2207 (N_2207,N_2122,N_2099);
nor U2208 (N_2208,N_2025,N_2118);
nand U2209 (N_2209,N_2028,N_2077);
and U2210 (N_2210,N_2093,N_2114);
xor U2211 (N_2211,N_2015,N_2085);
nor U2212 (N_2212,N_2079,N_2098);
nand U2213 (N_2213,N_2015,N_2075);
and U2214 (N_2214,N_2035,N_2083);
or U2215 (N_2215,N_2044,N_2019);
nand U2216 (N_2216,N_2043,N_2028);
or U2217 (N_2217,N_2013,N_2114);
nand U2218 (N_2218,N_2020,N_2101);
or U2219 (N_2219,N_2076,N_2058);
or U2220 (N_2220,N_2056,N_2011);
xnor U2221 (N_2221,N_2076,N_2027);
nor U2222 (N_2222,N_2047,N_2026);
xnor U2223 (N_2223,N_2032,N_2082);
or U2224 (N_2224,N_2010,N_2062);
nor U2225 (N_2225,N_2050,N_2015);
xor U2226 (N_2226,N_2074,N_2026);
nand U2227 (N_2227,N_2047,N_2043);
or U2228 (N_2228,N_2015,N_2081);
xor U2229 (N_2229,N_2108,N_2056);
nor U2230 (N_2230,N_2023,N_2049);
or U2231 (N_2231,N_2105,N_2072);
nand U2232 (N_2232,N_2087,N_2099);
or U2233 (N_2233,N_2076,N_2063);
or U2234 (N_2234,N_2072,N_2022);
nor U2235 (N_2235,N_2047,N_2067);
nor U2236 (N_2236,N_2092,N_2120);
nor U2237 (N_2237,N_2114,N_2025);
or U2238 (N_2238,N_2035,N_2040);
nand U2239 (N_2239,N_2023,N_2100);
nor U2240 (N_2240,N_2010,N_2019);
xnor U2241 (N_2241,N_2037,N_2103);
nor U2242 (N_2242,N_2067,N_2049);
nor U2243 (N_2243,N_2101,N_2083);
nand U2244 (N_2244,N_2071,N_2030);
and U2245 (N_2245,N_2124,N_2001);
or U2246 (N_2246,N_2047,N_2112);
nand U2247 (N_2247,N_2093,N_2082);
or U2248 (N_2248,N_2108,N_2020);
or U2249 (N_2249,N_2061,N_2072);
and U2250 (N_2250,N_2138,N_2143);
xnor U2251 (N_2251,N_2239,N_2189);
or U2252 (N_2252,N_2193,N_2235);
and U2253 (N_2253,N_2154,N_2157);
xor U2254 (N_2254,N_2139,N_2176);
nand U2255 (N_2255,N_2199,N_2246);
or U2256 (N_2256,N_2155,N_2172);
or U2257 (N_2257,N_2241,N_2227);
nand U2258 (N_2258,N_2133,N_2224);
nor U2259 (N_2259,N_2216,N_2188);
or U2260 (N_2260,N_2187,N_2228);
nand U2261 (N_2261,N_2226,N_2126);
nor U2262 (N_2262,N_2164,N_2184);
and U2263 (N_2263,N_2165,N_2147);
nand U2264 (N_2264,N_2173,N_2220);
and U2265 (N_2265,N_2207,N_2212);
and U2266 (N_2266,N_2217,N_2247);
nor U2267 (N_2267,N_2168,N_2135);
or U2268 (N_2268,N_2208,N_2209);
or U2269 (N_2269,N_2152,N_2240);
xnor U2270 (N_2270,N_2174,N_2236);
xnor U2271 (N_2271,N_2160,N_2128);
or U2272 (N_2272,N_2221,N_2134);
nor U2273 (N_2273,N_2202,N_2223);
xor U2274 (N_2274,N_2158,N_2183);
nand U2275 (N_2275,N_2162,N_2192);
nor U2276 (N_2276,N_2204,N_2175);
and U2277 (N_2277,N_2230,N_2177);
nor U2278 (N_2278,N_2132,N_2146);
and U2279 (N_2279,N_2218,N_2170);
xor U2280 (N_2280,N_2232,N_2182);
and U2281 (N_2281,N_2197,N_2245);
nor U2282 (N_2282,N_2150,N_2195);
and U2283 (N_2283,N_2178,N_2145);
or U2284 (N_2284,N_2169,N_2215);
xnor U2285 (N_2285,N_2234,N_2194);
or U2286 (N_2286,N_2243,N_2180);
nand U2287 (N_2287,N_2210,N_2242);
and U2288 (N_2288,N_2233,N_2151);
and U2289 (N_2289,N_2136,N_2156);
xor U2290 (N_2290,N_2213,N_2125);
nor U2291 (N_2291,N_2222,N_2130);
nand U2292 (N_2292,N_2237,N_2127);
nor U2293 (N_2293,N_2166,N_2198);
or U2294 (N_2294,N_2203,N_2185);
xnor U2295 (N_2295,N_2153,N_2191);
nor U2296 (N_2296,N_2141,N_2249);
and U2297 (N_2297,N_2161,N_2137);
xnor U2298 (N_2298,N_2196,N_2248);
and U2299 (N_2299,N_2238,N_2171);
xor U2300 (N_2300,N_2129,N_2225);
nor U2301 (N_2301,N_2200,N_2131);
or U2302 (N_2302,N_2206,N_2186);
and U2303 (N_2303,N_2179,N_2140);
nand U2304 (N_2304,N_2144,N_2159);
nor U2305 (N_2305,N_2211,N_2163);
nand U2306 (N_2306,N_2149,N_2214);
xor U2307 (N_2307,N_2167,N_2201);
nand U2308 (N_2308,N_2142,N_2205);
xor U2309 (N_2309,N_2231,N_2219);
nor U2310 (N_2310,N_2229,N_2190);
nor U2311 (N_2311,N_2181,N_2148);
nand U2312 (N_2312,N_2244,N_2129);
nand U2313 (N_2313,N_2148,N_2127);
and U2314 (N_2314,N_2248,N_2243);
nand U2315 (N_2315,N_2226,N_2137);
xnor U2316 (N_2316,N_2196,N_2164);
xor U2317 (N_2317,N_2131,N_2172);
and U2318 (N_2318,N_2233,N_2138);
nor U2319 (N_2319,N_2203,N_2183);
nor U2320 (N_2320,N_2214,N_2192);
and U2321 (N_2321,N_2127,N_2244);
or U2322 (N_2322,N_2135,N_2137);
xnor U2323 (N_2323,N_2129,N_2198);
or U2324 (N_2324,N_2171,N_2134);
nand U2325 (N_2325,N_2213,N_2134);
nor U2326 (N_2326,N_2134,N_2172);
xor U2327 (N_2327,N_2162,N_2212);
xor U2328 (N_2328,N_2149,N_2215);
nand U2329 (N_2329,N_2213,N_2215);
xnor U2330 (N_2330,N_2139,N_2201);
and U2331 (N_2331,N_2155,N_2186);
nand U2332 (N_2332,N_2163,N_2137);
and U2333 (N_2333,N_2156,N_2130);
and U2334 (N_2334,N_2223,N_2145);
nor U2335 (N_2335,N_2225,N_2147);
or U2336 (N_2336,N_2203,N_2209);
xor U2337 (N_2337,N_2227,N_2223);
nand U2338 (N_2338,N_2181,N_2184);
nand U2339 (N_2339,N_2221,N_2215);
nand U2340 (N_2340,N_2227,N_2173);
and U2341 (N_2341,N_2216,N_2182);
nand U2342 (N_2342,N_2174,N_2175);
nand U2343 (N_2343,N_2215,N_2204);
or U2344 (N_2344,N_2193,N_2241);
nand U2345 (N_2345,N_2185,N_2180);
nor U2346 (N_2346,N_2198,N_2203);
and U2347 (N_2347,N_2199,N_2224);
xnor U2348 (N_2348,N_2129,N_2138);
xnor U2349 (N_2349,N_2146,N_2176);
and U2350 (N_2350,N_2246,N_2160);
or U2351 (N_2351,N_2237,N_2149);
nor U2352 (N_2352,N_2171,N_2204);
nor U2353 (N_2353,N_2248,N_2217);
nor U2354 (N_2354,N_2175,N_2137);
nor U2355 (N_2355,N_2151,N_2185);
or U2356 (N_2356,N_2136,N_2188);
nand U2357 (N_2357,N_2137,N_2127);
and U2358 (N_2358,N_2210,N_2146);
nor U2359 (N_2359,N_2151,N_2152);
nor U2360 (N_2360,N_2219,N_2172);
or U2361 (N_2361,N_2177,N_2171);
nor U2362 (N_2362,N_2199,N_2147);
xnor U2363 (N_2363,N_2242,N_2240);
xnor U2364 (N_2364,N_2128,N_2179);
and U2365 (N_2365,N_2209,N_2154);
xnor U2366 (N_2366,N_2159,N_2225);
or U2367 (N_2367,N_2171,N_2219);
nor U2368 (N_2368,N_2225,N_2236);
xor U2369 (N_2369,N_2148,N_2217);
nand U2370 (N_2370,N_2146,N_2125);
or U2371 (N_2371,N_2208,N_2228);
nor U2372 (N_2372,N_2190,N_2202);
nor U2373 (N_2373,N_2140,N_2209);
nor U2374 (N_2374,N_2232,N_2160);
or U2375 (N_2375,N_2289,N_2351);
xnor U2376 (N_2376,N_2286,N_2319);
or U2377 (N_2377,N_2301,N_2264);
nand U2378 (N_2378,N_2348,N_2257);
nand U2379 (N_2379,N_2297,N_2345);
nand U2380 (N_2380,N_2312,N_2295);
and U2381 (N_2381,N_2284,N_2335);
nor U2382 (N_2382,N_2256,N_2262);
nor U2383 (N_2383,N_2261,N_2278);
nand U2384 (N_2384,N_2330,N_2300);
xnor U2385 (N_2385,N_2314,N_2294);
nor U2386 (N_2386,N_2373,N_2324);
or U2387 (N_2387,N_2267,N_2325);
xor U2388 (N_2388,N_2276,N_2367);
or U2389 (N_2389,N_2341,N_2309);
and U2390 (N_2390,N_2282,N_2350);
or U2391 (N_2391,N_2337,N_2327);
xor U2392 (N_2392,N_2349,N_2293);
and U2393 (N_2393,N_2359,N_2275);
nor U2394 (N_2394,N_2328,N_2272);
nand U2395 (N_2395,N_2281,N_2310);
and U2396 (N_2396,N_2279,N_2326);
nor U2397 (N_2397,N_2255,N_2342);
nor U2398 (N_2398,N_2265,N_2334);
nor U2399 (N_2399,N_2290,N_2344);
nand U2400 (N_2400,N_2303,N_2339);
nand U2401 (N_2401,N_2362,N_2365);
or U2402 (N_2402,N_2283,N_2298);
and U2403 (N_2403,N_2288,N_2277);
xnor U2404 (N_2404,N_2370,N_2331);
nor U2405 (N_2405,N_2258,N_2266);
and U2406 (N_2406,N_2299,N_2305);
nor U2407 (N_2407,N_2273,N_2287);
or U2408 (N_2408,N_2292,N_2346);
and U2409 (N_2409,N_2251,N_2311);
nand U2410 (N_2410,N_2374,N_2313);
nor U2411 (N_2411,N_2323,N_2316);
and U2412 (N_2412,N_2332,N_2271);
nand U2413 (N_2413,N_2304,N_2285);
or U2414 (N_2414,N_2357,N_2274);
nor U2415 (N_2415,N_2369,N_2354);
xor U2416 (N_2416,N_2296,N_2347);
nand U2417 (N_2417,N_2368,N_2356);
nand U2418 (N_2418,N_2372,N_2364);
and U2419 (N_2419,N_2338,N_2259);
nor U2420 (N_2420,N_2329,N_2308);
xor U2421 (N_2421,N_2253,N_2333);
xor U2422 (N_2422,N_2307,N_2353);
xnor U2423 (N_2423,N_2352,N_2315);
and U2424 (N_2424,N_2343,N_2321);
or U2425 (N_2425,N_2355,N_2252);
nor U2426 (N_2426,N_2371,N_2322);
and U2427 (N_2427,N_2366,N_2263);
or U2428 (N_2428,N_2361,N_2270);
or U2429 (N_2429,N_2302,N_2250);
or U2430 (N_2430,N_2291,N_2268);
and U2431 (N_2431,N_2306,N_2318);
xnor U2432 (N_2432,N_2317,N_2340);
and U2433 (N_2433,N_2254,N_2320);
and U2434 (N_2434,N_2336,N_2358);
nand U2435 (N_2435,N_2269,N_2363);
nand U2436 (N_2436,N_2360,N_2280);
nor U2437 (N_2437,N_2260,N_2323);
nand U2438 (N_2438,N_2258,N_2326);
and U2439 (N_2439,N_2296,N_2374);
and U2440 (N_2440,N_2261,N_2321);
or U2441 (N_2441,N_2323,N_2258);
or U2442 (N_2442,N_2318,N_2317);
nand U2443 (N_2443,N_2319,N_2325);
nand U2444 (N_2444,N_2306,N_2373);
nor U2445 (N_2445,N_2319,N_2254);
nand U2446 (N_2446,N_2291,N_2296);
or U2447 (N_2447,N_2301,N_2330);
nor U2448 (N_2448,N_2345,N_2272);
or U2449 (N_2449,N_2308,N_2314);
nand U2450 (N_2450,N_2256,N_2358);
and U2451 (N_2451,N_2371,N_2360);
nor U2452 (N_2452,N_2262,N_2352);
nor U2453 (N_2453,N_2365,N_2363);
and U2454 (N_2454,N_2371,N_2320);
nand U2455 (N_2455,N_2287,N_2308);
xnor U2456 (N_2456,N_2283,N_2348);
nor U2457 (N_2457,N_2368,N_2272);
nand U2458 (N_2458,N_2365,N_2374);
nor U2459 (N_2459,N_2329,N_2374);
or U2460 (N_2460,N_2273,N_2268);
and U2461 (N_2461,N_2324,N_2301);
and U2462 (N_2462,N_2366,N_2334);
xnor U2463 (N_2463,N_2366,N_2278);
or U2464 (N_2464,N_2257,N_2280);
and U2465 (N_2465,N_2305,N_2282);
nor U2466 (N_2466,N_2320,N_2368);
and U2467 (N_2467,N_2294,N_2281);
and U2468 (N_2468,N_2319,N_2253);
xnor U2469 (N_2469,N_2250,N_2354);
and U2470 (N_2470,N_2348,N_2282);
and U2471 (N_2471,N_2301,N_2303);
and U2472 (N_2472,N_2361,N_2268);
nor U2473 (N_2473,N_2320,N_2279);
and U2474 (N_2474,N_2332,N_2359);
nand U2475 (N_2475,N_2312,N_2260);
nor U2476 (N_2476,N_2345,N_2362);
and U2477 (N_2477,N_2295,N_2371);
or U2478 (N_2478,N_2319,N_2314);
nand U2479 (N_2479,N_2268,N_2289);
xnor U2480 (N_2480,N_2337,N_2254);
nand U2481 (N_2481,N_2272,N_2255);
and U2482 (N_2482,N_2267,N_2284);
xor U2483 (N_2483,N_2284,N_2301);
xor U2484 (N_2484,N_2318,N_2358);
or U2485 (N_2485,N_2332,N_2270);
or U2486 (N_2486,N_2346,N_2309);
nor U2487 (N_2487,N_2320,N_2253);
nand U2488 (N_2488,N_2271,N_2367);
xnor U2489 (N_2489,N_2360,N_2324);
nor U2490 (N_2490,N_2345,N_2336);
nor U2491 (N_2491,N_2286,N_2329);
and U2492 (N_2492,N_2280,N_2328);
or U2493 (N_2493,N_2354,N_2317);
or U2494 (N_2494,N_2277,N_2304);
and U2495 (N_2495,N_2270,N_2297);
or U2496 (N_2496,N_2308,N_2298);
xor U2497 (N_2497,N_2293,N_2343);
xor U2498 (N_2498,N_2272,N_2290);
and U2499 (N_2499,N_2339,N_2287);
nand U2500 (N_2500,N_2429,N_2452);
or U2501 (N_2501,N_2474,N_2457);
nor U2502 (N_2502,N_2490,N_2385);
or U2503 (N_2503,N_2497,N_2440);
xor U2504 (N_2504,N_2465,N_2383);
nand U2505 (N_2505,N_2389,N_2478);
xnor U2506 (N_2506,N_2477,N_2413);
xnor U2507 (N_2507,N_2476,N_2392);
xor U2508 (N_2508,N_2404,N_2405);
nor U2509 (N_2509,N_2393,N_2428);
or U2510 (N_2510,N_2398,N_2441);
or U2511 (N_2511,N_2412,N_2408);
nand U2512 (N_2512,N_2489,N_2459);
nand U2513 (N_2513,N_2400,N_2401);
and U2514 (N_2514,N_2443,N_2486);
nand U2515 (N_2515,N_2399,N_2484);
xnor U2516 (N_2516,N_2461,N_2480);
nand U2517 (N_2517,N_2499,N_2445);
nor U2518 (N_2518,N_2382,N_2379);
nor U2519 (N_2519,N_2384,N_2479);
and U2520 (N_2520,N_2475,N_2492);
and U2521 (N_2521,N_2495,N_2494);
xnor U2522 (N_2522,N_2431,N_2396);
nand U2523 (N_2523,N_2426,N_2435);
nand U2524 (N_2524,N_2462,N_2472);
nand U2525 (N_2525,N_2380,N_2451);
or U2526 (N_2526,N_2381,N_2436);
nor U2527 (N_2527,N_2427,N_2424);
or U2528 (N_2528,N_2432,N_2468);
nand U2529 (N_2529,N_2395,N_2444);
nor U2530 (N_2530,N_2425,N_2455);
nand U2531 (N_2531,N_2378,N_2488);
nand U2532 (N_2532,N_2447,N_2386);
or U2533 (N_2533,N_2482,N_2415);
or U2534 (N_2534,N_2407,N_2377);
or U2535 (N_2535,N_2390,N_2471);
or U2536 (N_2536,N_2421,N_2391);
and U2537 (N_2537,N_2460,N_2397);
nand U2538 (N_2538,N_2442,N_2469);
xnor U2539 (N_2539,N_2403,N_2473);
nor U2540 (N_2540,N_2439,N_2487);
nand U2541 (N_2541,N_2437,N_2456);
and U2542 (N_2542,N_2406,N_2483);
and U2543 (N_2543,N_2388,N_2375);
nand U2544 (N_2544,N_2423,N_2496);
and U2545 (N_2545,N_2438,N_2467);
nand U2546 (N_2546,N_2481,N_2464);
or U2547 (N_2547,N_2434,N_2409);
and U2548 (N_2548,N_2463,N_2458);
nand U2549 (N_2549,N_2420,N_2446);
xor U2550 (N_2550,N_2419,N_2410);
nor U2551 (N_2551,N_2498,N_2394);
and U2552 (N_2552,N_2418,N_2491);
xnor U2553 (N_2553,N_2453,N_2448);
or U2554 (N_2554,N_2485,N_2470);
nor U2555 (N_2555,N_2493,N_2430);
and U2556 (N_2556,N_2417,N_2376);
xnor U2557 (N_2557,N_2450,N_2414);
nor U2558 (N_2558,N_2411,N_2433);
and U2559 (N_2559,N_2454,N_2449);
nor U2560 (N_2560,N_2402,N_2416);
xor U2561 (N_2561,N_2422,N_2387);
nor U2562 (N_2562,N_2466,N_2391);
or U2563 (N_2563,N_2458,N_2410);
and U2564 (N_2564,N_2430,N_2401);
nor U2565 (N_2565,N_2420,N_2479);
or U2566 (N_2566,N_2397,N_2387);
and U2567 (N_2567,N_2498,N_2490);
nand U2568 (N_2568,N_2404,N_2473);
nor U2569 (N_2569,N_2473,N_2408);
nand U2570 (N_2570,N_2458,N_2440);
or U2571 (N_2571,N_2375,N_2448);
or U2572 (N_2572,N_2437,N_2469);
and U2573 (N_2573,N_2459,N_2456);
nor U2574 (N_2574,N_2376,N_2432);
or U2575 (N_2575,N_2384,N_2452);
nand U2576 (N_2576,N_2458,N_2379);
nand U2577 (N_2577,N_2435,N_2440);
or U2578 (N_2578,N_2493,N_2417);
nand U2579 (N_2579,N_2432,N_2445);
nand U2580 (N_2580,N_2432,N_2385);
xor U2581 (N_2581,N_2425,N_2416);
or U2582 (N_2582,N_2427,N_2486);
nor U2583 (N_2583,N_2399,N_2498);
nor U2584 (N_2584,N_2446,N_2380);
xor U2585 (N_2585,N_2405,N_2463);
xor U2586 (N_2586,N_2412,N_2396);
and U2587 (N_2587,N_2447,N_2438);
nand U2588 (N_2588,N_2379,N_2403);
nor U2589 (N_2589,N_2411,N_2432);
nand U2590 (N_2590,N_2499,N_2393);
xnor U2591 (N_2591,N_2456,N_2434);
and U2592 (N_2592,N_2450,N_2415);
xor U2593 (N_2593,N_2429,N_2455);
or U2594 (N_2594,N_2433,N_2487);
and U2595 (N_2595,N_2450,N_2449);
nor U2596 (N_2596,N_2447,N_2398);
xnor U2597 (N_2597,N_2492,N_2406);
xor U2598 (N_2598,N_2378,N_2422);
or U2599 (N_2599,N_2469,N_2383);
or U2600 (N_2600,N_2483,N_2421);
or U2601 (N_2601,N_2471,N_2397);
and U2602 (N_2602,N_2377,N_2494);
nor U2603 (N_2603,N_2383,N_2441);
xor U2604 (N_2604,N_2387,N_2391);
or U2605 (N_2605,N_2395,N_2430);
nand U2606 (N_2606,N_2498,N_2415);
nor U2607 (N_2607,N_2495,N_2497);
or U2608 (N_2608,N_2414,N_2425);
or U2609 (N_2609,N_2488,N_2496);
or U2610 (N_2610,N_2476,N_2430);
or U2611 (N_2611,N_2467,N_2405);
nor U2612 (N_2612,N_2483,N_2448);
or U2613 (N_2613,N_2494,N_2411);
nor U2614 (N_2614,N_2389,N_2396);
nor U2615 (N_2615,N_2483,N_2443);
nand U2616 (N_2616,N_2487,N_2413);
nand U2617 (N_2617,N_2486,N_2448);
nor U2618 (N_2618,N_2400,N_2458);
xor U2619 (N_2619,N_2426,N_2432);
or U2620 (N_2620,N_2388,N_2487);
nand U2621 (N_2621,N_2498,N_2429);
nor U2622 (N_2622,N_2422,N_2402);
nand U2623 (N_2623,N_2477,N_2388);
xnor U2624 (N_2624,N_2427,N_2476);
nand U2625 (N_2625,N_2546,N_2543);
nor U2626 (N_2626,N_2568,N_2529);
nand U2627 (N_2627,N_2502,N_2577);
nand U2628 (N_2628,N_2613,N_2616);
nand U2629 (N_2629,N_2586,N_2501);
xor U2630 (N_2630,N_2536,N_2575);
xor U2631 (N_2631,N_2560,N_2516);
nand U2632 (N_2632,N_2618,N_2510);
or U2633 (N_2633,N_2592,N_2549);
nand U2634 (N_2634,N_2559,N_2563);
nor U2635 (N_2635,N_2503,N_2500);
nor U2636 (N_2636,N_2544,N_2610);
and U2637 (N_2637,N_2581,N_2562);
nand U2638 (N_2638,N_2611,N_2506);
nor U2639 (N_2639,N_2558,N_2538);
nor U2640 (N_2640,N_2573,N_2583);
or U2641 (N_2641,N_2523,N_2580);
or U2642 (N_2642,N_2596,N_2569);
xor U2643 (N_2643,N_2572,N_2590);
or U2644 (N_2644,N_2621,N_2519);
nand U2645 (N_2645,N_2597,N_2508);
nand U2646 (N_2646,N_2540,N_2623);
and U2647 (N_2647,N_2522,N_2513);
nor U2648 (N_2648,N_2578,N_2620);
and U2649 (N_2649,N_2521,N_2601);
and U2650 (N_2650,N_2574,N_2619);
nor U2651 (N_2651,N_2589,N_2603);
nor U2652 (N_2652,N_2518,N_2554);
nor U2653 (N_2653,N_2552,N_2515);
or U2654 (N_2654,N_2524,N_2591);
xnor U2655 (N_2655,N_2588,N_2551);
or U2656 (N_2656,N_2605,N_2604);
xor U2657 (N_2657,N_2507,N_2566);
xnor U2658 (N_2658,N_2614,N_2557);
or U2659 (N_2659,N_2579,N_2509);
and U2660 (N_2660,N_2624,N_2533);
and U2661 (N_2661,N_2525,N_2520);
or U2662 (N_2662,N_2599,N_2505);
nor U2663 (N_2663,N_2587,N_2545);
or U2664 (N_2664,N_2528,N_2531);
nand U2665 (N_2665,N_2556,N_2537);
nor U2666 (N_2666,N_2530,N_2514);
or U2667 (N_2667,N_2582,N_2564);
or U2668 (N_2668,N_2593,N_2561);
and U2669 (N_2669,N_2585,N_2534);
xnor U2670 (N_2670,N_2532,N_2555);
nand U2671 (N_2671,N_2535,N_2541);
nand U2672 (N_2672,N_2606,N_2608);
xnor U2673 (N_2673,N_2576,N_2584);
nor U2674 (N_2674,N_2511,N_2550);
or U2675 (N_2675,N_2598,N_2547);
or U2676 (N_2676,N_2622,N_2565);
and U2677 (N_2677,N_2612,N_2548);
nor U2678 (N_2678,N_2595,N_2600);
nor U2679 (N_2679,N_2512,N_2567);
xor U2680 (N_2680,N_2594,N_2527);
or U2681 (N_2681,N_2517,N_2571);
or U2682 (N_2682,N_2504,N_2609);
xor U2683 (N_2683,N_2615,N_2526);
nor U2684 (N_2684,N_2617,N_2539);
xor U2685 (N_2685,N_2553,N_2570);
nand U2686 (N_2686,N_2607,N_2542);
and U2687 (N_2687,N_2602,N_2514);
xnor U2688 (N_2688,N_2530,N_2591);
nand U2689 (N_2689,N_2587,N_2617);
and U2690 (N_2690,N_2595,N_2617);
nand U2691 (N_2691,N_2562,N_2502);
and U2692 (N_2692,N_2551,N_2587);
and U2693 (N_2693,N_2608,N_2568);
nand U2694 (N_2694,N_2595,N_2528);
or U2695 (N_2695,N_2622,N_2572);
nand U2696 (N_2696,N_2607,N_2545);
nand U2697 (N_2697,N_2603,N_2531);
xnor U2698 (N_2698,N_2615,N_2514);
xor U2699 (N_2699,N_2573,N_2544);
or U2700 (N_2700,N_2538,N_2548);
nor U2701 (N_2701,N_2508,N_2556);
nand U2702 (N_2702,N_2528,N_2600);
and U2703 (N_2703,N_2538,N_2554);
and U2704 (N_2704,N_2602,N_2526);
and U2705 (N_2705,N_2500,N_2613);
xnor U2706 (N_2706,N_2502,N_2611);
xnor U2707 (N_2707,N_2516,N_2587);
or U2708 (N_2708,N_2510,N_2594);
or U2709 (N_2709,N_2574,N_2506);
nand U2710 (N_2710,N_2545,N_2532);
and U2711 (N_2711,N_2521,N_2538);
or U2712 (N_2712,N_2537,N_2622);
nand U2713 (N_2713,N_2534,N_2571);
nor U2714 (N_2714,N_2586,N_2509);
nor U2715 (N_2715,N_2603,N_2500);
or U2716 (N_2716,N_2605,N_2543);
nor U2717 (N_2717,N_2586,N_2575);
nor U2718 (N_2718,N_2523,N_2548);
nor U2719 (N_2719,N_2532,N_2610);
or U2720 (N_2720,N_2601,N_2509);
nor U2721 (N_2721,N_2501,N_2518);
and U2722 (N_2722,N_2607,N_2517);
nand U2723 (N_2723,N_2530,N_2506);
nand U2724 (N_2724,N_2585,N_2562);
nor U2725 (N_2725,N_2610,N_2546);
nor U2726 (N_2726,N_2534,N_2612);
and U2727 (N_2727,N_2511,N_2506);
nor U2728 (N_2728,N_2621,N_2534);
nor U2729 (N_2729,N_2527,N_2537);
and U2730 (N_2730,N_2517,N_2565);
nand U2731 (N_2731,N_2513,N_2558);
nor U2732 (N_2732,N_2583,N_2600);
and U2733 (N_2733,N_2621,N_2533);
and U2734 (N_2734,N_2532,N_2620);
or U2735 (N_2735,N_2510,N_2604);
nand U2736 (N_2736,N_2545,N_2557);
or U2737 (N_2737,N_2548,N_2524);
nor U2738 (N_2738,N_2522,N_2543);
and U2739 (N_2739,N_2581,N_2590);
or U2740 (N_2740,N_2510,N_2524);
or U2741 (N_2741,N_2620,N_2581);
xnor U2742 (N_2742,N_2560,N_2519);
and U2743 (N_2743,N_2558,N_2622);
and U2744 (N_2744,N_2504,N_2572);
and U2745 (N_2745,N_2561,N_2586);
xnor U2746 (N_2746,N_2611,N_2558);
xor U2747 (N_2747,N_2541,N_2553);
and U2748 (N_2748,N_2532,N_2548);
or U2749 (N_2749,N_2563,N_2622);
nand U2750 (N_2750,N_2658,N_2639);
xor U2751 (N_2751,N_2687,N_2653);
xor U2752 (N_2752,N_2690,N_2664);
and U2753 (N_2753,N_2627,N_2677);
xnor U2754 (N_2754,N_2652,N_2667);
or U2755 (N_2755,N_2713,N_2657);
nand U2756 (N_2756,N_2626,N_2715);
nand U2757 (N_2757,N_2697,N_2704);
and U2758 (N_2758,N_2685,N_2730);
and U2759 (N_2759,N_2702,N_2647);
nand U2760 (N_2760,N_2747,N_2719);
nor U2761 (N_2761,N_2726,N_2705);
xnor U2762 (N_2762,N_2633,N_2741);
xor U2763 (N_2763,N_2672,N_2695);
nand U2764 (N_2764,N_2640,N_2665);
xnor U2765 (N_2765,N_2717,N_2675);
nor U2766 (N_2766,N_2650,N_2708);
or U2767 (N_2767,N_2729,N_2628);
xor U2768 (N_2768,N_2720,N_2688);
nor U2769 (N_2769,N_2714,N_2638);
or U2770 (N_2770,N_2686,N_2651);
xnor U2771 (N_2771,N_2699,N_2625);
or U2772 (N_2772,N_2663,N_2703);
and U2773 (N_2773,N_2731,N_2746);
and U2774 (N_2774,N_2644,N_2724);
nor U2775 (N_2775,N_2678,N_2706);
xnor U2776 (N_2776,N_2740,N_2723);
nor U2777 (N_2777,N_2749,N_2721);
or U2778 (N_2778,N_2669,N_2737);
and U2779 (N_2779,N_2635,N_2679);
xnor U2780 (N_2780,N_2630,N_2693);
xor U2781 (N_2781,N_2738,N_2733);
nand U2782 (N_2782,N_2683,N_2691);
xor U2783 (N_2783,N_2722,N_2643);
nand U2784 (N_2784,N_2710,N_2646);
nor U2785 (N_2785,N_2641,N_2745);
nor U2786 (N_2786,N_2735,N_2707);
xor U2787 (N_2787,N_2734,N_2732);
xnor U2788 (N_2788,N_2742,N_2666);
nor U2789 (N_2789,N_2670,N_2682);
or U2790 (N_2790,N_2712,N_2739);
xor U2791 (N_2791,N_2673,N_2676);
nand U2792 (N_2792,N_2656,N_2637);
nand U2793 (N_2793,N_2727,N_2736);
or U2794 (N_2794,N_2684,N_2701);
xnor U2795 (N_2795,N_2654,N_2681);
nand U2796 (N_2796,N_2674,N_2700);
nand U2797 (N_2797,N_2725,N_2716);
nor U2798 (N_2798,N_2648,N_2661);
xor U2799 (N_2799,N_2748,N_2629);
and U2800 (N_2800,N_2631,N_2696);
or U2801 (N_2801,N_2645,N_2649);
nor U2802 (N_2802,N_2655,N_2711);
nor U2803 (N_2803,N_2634,N_2671);
and U2804 (N_2804,N_2659,N_2709);
xor U2805 (N_2805,N_2694,N_2642);
xor U2806 (N_2806,N_2660,N_2692);
nor U2807 (N_2807,N_2668,N_2689);
or U2808 (N_2808,N_2718,N_2632);
xor U2809 (N_2809,N_2743,N_2744);
nand U2810 (N_2810,N_2728,N_2680);
xor U2811 (N_2811,N_2662,N_2636);
xnor U2812 (N_2812,N_2698,N_2635);
nand U2813 (N_2813,N_2680,N_2638);
xor U2814 (N_2814,N_2648,N_2679);
nand U2815 (N_2815,N_2720,N_2693);
nor U2816 (N_2816,N_2715,N_2709);
nor U2817 (N_2817,N_2658,N_2663);
and U2818 (N_2818,N_2713,N_2725);
nor U2819 (N_2819,N_2631,N_2709);
nor U2820 (N_2820,N_2700,N_2733);
or U2821 (N_2821,N_2749,N_2675);
xnor U2822 (N_2822,N_2709,N_2628);
xor U2823 (N_2823,N_2707,N_2730);
xor U2824 (N_2824,N_2741,N_2714);
xnor U2825 (N_2825,N_2741,N_2718);
or U2826 (N_2826,N_2665,N_2678);
and U2827 (N_2827,N_2740,N_2726);
xnor U2828 (N_2828,N_2718,N_2634);
xnor U2829 (N_2829,N_2629,N_2701);
and U2830 (N_2830,N_2635,N_2722);
or U2831 (N_2831,N_2668,N_2639);
nand U2832 (N_2832,N_2682,N_2712);
nand U2833 (N_2833,N_2674,N_2749);
nor U2834 (N_2834,N_2733,N_2669);
xor U2835 (N_2835,N_2652,N_2720);
nor U2836 (N_2836,N_2720,N_2709);
nand U2837 (N_2837,N_2665,N_2725);
nand U2838 (N_2838,N_2666,N_2709);
and U2839 (N_2839,N_2706,N_2657);
nand U2840 (N_2840,N_2639,N_2654);
nor U2841 (N_2841,N_2711,N_2652);
nand U2842 (N_2842,N_2643,N_2673);
or U2843 (N_2843,N_2710,N_2677);
and U2844 (N_2844,N_2701,N_2677);
nor U2845 (N_2845,N_2651,N_2736);
and U2846 (N_2846,N_2680,N_2655);
nand U2847 (N_2847,N_2685,N_2692);
and U2848 (N_2848,N_2697,N_2730);
nor U2849 (N_2849,N_2634,N_2632);
nand U2850 (N_2850,N_2633,N_2715);
nand U2851 (N_2851,N_2663,N_2648);
or U2852 (N_2852,N_2690,N_2724);
xnor U2853 (N_2853,N_2745,N_2635);
nor U2854 (N_2854,N_2625,N_2731);
nand U2855 (N_2855,N_2694,N_2681);
or U2856 (N_2856,N_2675,N_2678);
xnor U2857 (N_2857,N_2644,N_2704);
nand U2858 (N_2858,N_2692,N_2701);
and U2859 (N_2859,N_2659,N_2679);
and U2860 (N_2860,N_2724,N_2675);
nand U2861 (N_2861,N_2668,N_2637);
or U2862 (N_2862,N_2698,N_2699);
and U2863 (N_2863,N_2745,N_2719);
nor U2864 (N_2864,N_2703,N_2749);
nand U2865 (N_2865,N_2654,N_2689);
nand U2866 (N_2866,N_2682,N_2740);
nor U2867 (N_2867,N_2638,N_2627);
xor U2868 (N_2868,N_2731,N_2669);
xnor U2869 (N_2869,N_2691,N_2669);
or U2870 (N_2870,N_2696,N_2664);
and U2871 (N_2871,N_2726,N_2663);
nor U2872 (N_2872,N_2730,N_2664);
xnor U2873 (N_2873,N_2666,N_2689);
and U2874 (N_2874,N_2635,N_2644);
nand U2875 (N_2875,N_2853,N_2774);
xnor U2876 (N_2876,N_2865,N_2779);
xor U2877 (N_2877,N_2790,N_2824);
and U2878 (N_2878,N_2791,N_2796);
or U2879 (N_2879,N_2834,N_2828);
nand U2880 (N_2880,N_2866,N_2783);
nor U2881 (N_2881,N_2789,N_2864);
xor U2882 (N_2882,N_2842,N_2802);
nand U2883 (N_2883,N_2849,N_2841);
xor U2884 (N_2884,N_2792,N_2831);
or U2885 (N_2885,N_2823,N_2773);
nor U2886 (N_2886,N_2797,N_2811);
and U2887 (N_2887,N_2847,N_2848);
nor U2888 (N_2888,N_2872,N_2817);
or U2889 (N_2889,N_2846,N_2758);
nand U2890 (N_2890,N_2835,N_2857);
or U2891 (N_2891,N_2754,N_2837);
nor U2892 (N_2892,N_2814,N_2839);
nand U2893 (N_2893,N_2852,N_2759);
nand U2894 (N_2894,N_2771,N_2810);
nand U2895 (N_2895,N_2809,N_2769);
xnor U2896 (N_2896,N_2840,N_2816);
and U2897 (N_2897,N_2766,N_2775);
or U2898 (N_2898,N_2788,N_2818);
nand U2899 (N_2899,N_2752,N_2757);
xor U2900 (N_2900,N_2761,N_2772);
nor U2901 (N_2901,N_2832,N_2874);
nor U2902 (N_2902,N_2830,N_2870);
or U2903 (N_2903,N_2803,N_2871);
nand U2904 (N_2904,N_2845,N_2873);
xnor U2905 (N_2905,N_2776,N_2860);
and U2906 (N_2906,N_2777,N_2787);
and U2907 (N_2907,N_2786,N_2856);
or U2908 (N_2908,N_2868,N_2760);
nand U2909 (N_2909,N_2855,N_2751);
or U2910 (N_2910,N_2782,N_2770);
nand U2911 (N_2911,N_2762,N_2812);
or U2912 (N_2912,N_2805,N_2780);
and U2913 (N_2913,N_2808,N_2784);
xnor U2914 (N_2914,N_2862,N_2843);
or U2915 (N_2915,N_2807,N_2756);
or U2916 (N_2916,N_2867,N_2795);
or U2917 (N_2917,N_2765,N_2815);
xor U2918 (N_2918,N_2763,N_2785);
nor U2919 (N_2919,N_2767,N_2768);
xor U2920 (N_2920,N_2820,N_2819);
and U2921 (N_2921,N_2753,N_2826);
or U2922 (N_2922,N_2822,N_2781);
xnor U2923 (N_2923,N_2858,N_2859);
nand U2924 (N_2924,N_2825,N_2750);
xor U2925 (N_2925,N_2861,N_2827);
and U2926 (N_2926,N_2844,N_2798);
nand U2927 (N_2927,N_2800,N_2829);
nor U2928 (N_2928,N_2863,N_2854);
nand U2929 (N_2929,N_2833,N_2850);
and U2930 (N_2930,N_2821,N_2799);
or U2931 (N_2931,N_2801,N_2851);
nor U2932 (N_2932,N_2793,N_2836);
or U2933 (N_2933,N_2764,N_2806);
nand U2934 (N_2934,N_2813,N_2778);
nand U2935 (N_2935,N_2794,N_2869);
nor U2936 (N_2936,N_2804,N_2755);
xnor U2937 (N_2937,N_2838,N_2852);
nand U2938 (N_2938,N_2796,N_2865);
nor U2939 (N_2939,N_2873,N_2793);
or U2940 (N_2940,N_2751,N_2830);
nand U2941 (N_2941,N_2844,N_2854);
nand U2942 (N_2942,N_2796,N_2837);
or U2943 (N_2943,N_2826,N_2839);
nand U2944 (N_2944,N_2844,N_2809);
nand U2945 (N_2945,N_2778,N_2754);
and U2946 (N_2946,N_2828,N_2870);
nand U2947 (N_2947,N_2817,N_2798);
nand U2948 (N_2948,N_2761,N_2768);
and U2949 (N_2949,N_2817,N_2764);
or U2950 (N_2950,N_2814,N_2781);
nor U2951 (N_2951,N_2769,N_2789);
nand U2952 (N_2952,N_2784,N_2834);
xnor U2953 (N_2953,N_2871,N_2808);
nand U2954 (N_2954,N_2789,N_2772);
and U2955 (N_2955,N_2789,N_2816);
nand U2956 (N_2956,N_2781,N_2872);
and U2957 (N_2957,N_2822,N_2867);
xnor U2958 (N_2958,N_2774,N_2757);
nor U2959 (N_2959,N_2790,N_2862);
or U2960 (N_2960,N_2802,N_2757);
nand U2961 (N_2961,N_2820,N_2753);
and U2962 (N_2962,N_2834,N_2816);
and U2963 (N_2963,N_2782,N_2868);
nand U2964 (N_2964,N_2757,N_2763);
nand U2965 (N_2965,N_2847,N_2764);
xor U2966 (N_2966,N_2854,N_2757);
and U2967 (N_2967,N_2843,N_2861);
nand U2968 (N_2968,N_2844,N_2788);
nand U2969 (N_2969,N_2857,N_2834);
xnor U2970 (N_2970,N_2860,N_2865);
xor U2971 (N_2971,N_2803,N_2821);
or U2972 (N_2972,N_2831,N_2803);
nor U2973 (N_2973,N_2859,N_2785);
nand U2974 (N_2974,N_2783,N_2777);
nor U2975 (N_2975,N_2858,N_2809);
and U2976 (N_2976,N_2799,N_2837);
xor U2977 (N_2977,N_2863,N_2774);
or U2978 (N_2978,N_2840,N_2859);
xor U2979 (N_2979,N_2775,N_2778);
or U2980 (N_2980,N_2792,N_2862);
nor U2981 (N_2981,N_2851,N_2853);
nand U2982 (N_2982,N_2764,N_2753);
xor U2983 (N_2983,N_2797,N_2810);
nand U2984 (N_2984,N_2830,N_2805);
or U2985 (N_2985,N_2779,N_2819);
nand U2986 (N_2986,N_2866,N_2841);
nand U2987 (N_2987,N_2759,N_2788);
xnor U2988 (N_2988,N_2789,N_2793);
or U2989 (N_2989,N_2851,N_2854);
nor U2990 (N_2990,N_2754,N_2786);
xor U2991 (N_2991,N_2780,N_2782);
xor U2992 (N_2992,N_2807,N_2837);
nor U2993 (N_2993,N_2827,N_2806);
and U2994 (N_2994,N_2838,N_2842);
nand U2995 (N_2995,N_2780,N_2767);
and U2996 (N_2996,N_2762,N_2846);
xor U2997 (N_2997,N_2832,N_2812);
nand U2998 (N_2998,N_2870,N_2780);
and U2999 (N_2999,N_2785,N_2822);
and U3000 (N_3000,N_2885,N_2970);
or U3001 (N_3001,N_2921,N_2933);
and U3002 (N_3002,N_2919,N_2883);
or U3003 (N_3003,N_2884,N_2988);
nor U3004 (N_3004,N_2879,N_2881);
xnor U3005 (N_3005,N_2907,N_2904);
nand U3006 (N_3006,N_2901,N_2940);
nor U3007 (N_3007,N_2877,N_2938);
and U3008 (N_3008,N_2913,N_2966);
xor U3009 (N_3009,N_2977,N_2914);
and U3010 (N_3010,N_2962,N_2953);
or U3011 (N_3011,N_2930,N_2915);
nor U3012 (N_3012,N_2982,N_2889);
nand U3013 (N_3013,N_2891,N_2939);
or U3014 (N_3014,N_2998,N_2945);
and U3015 (N_3015,N_2957,N_2990);
nor U3016 (N_3016,N_2886,N_2931);
xnor U3017 (N_3017,N_2952,N_2906);
xor U3018 (N_3018,N_2999,N_2965);
and U3019 (N_3019,N_2972,N_2934);
or U3020 (N_3020,N_2908,N_2880);
nor U3021 (N_3021,N_2887,N_2892);
nand U3022 (N_3022,N_2942,N_2897);
or U3023 (N_3023,N_2958,N_2959);
or U3024 (N_3024,N_2925,N_2956);
xnor U3025 (N_3025,N_2949,N_2987);
xnor U3026 (N_3026,N_2995,N_2882);
or U3027 (N_3027,N_2929,N_2893);
nand U3028 (N_3028,N_2968,N_2935);
and U3029 (N_3029,N_2916,N_2991);
and U3030 (N_3030,N_2961,N_2983);
or U3031 (N_3031,N_2946,N_2955);
xor U3032 (N_3032,N_2912,N_2928);
nand U3033 (N_3033,N_2924,N_2986);
xnor U3034 (N_3034,N_2993,N_2898);
or U3035 (N_3035,N_2964,N_2927);
xnor U3036 (N_3036,N_2932,N_2903);
or U3037 (N_3037,N_2979,N_2905);
and U3038 (N_3038,N_2917,N_2975);
nor U3039 (N_3039,N_2944,N_2948);
nand U3040 (N_3040,N_2947,N_2967);
xnor U3041 (N_3041,N_2876,N_2894);
xnor U3042 (N_3042,N_2984,N_2994);
and U3043 (N_3043,N_2910,N_2974);
nand U3044 (N_3044,N_2902,N_2985);
and U3045 (N_3045,N_2918,N_2937);
or U3046 (N_3046,N_2875,N_2896);
or U3047 (N_3047,N_2941,N_2943);
xor U3048 (N_3048,N_2900,N_2911);
and U3049 (N_3049,N_2963,N_2951);
and U3050 (N_3050,N_2878,N_2922);
and U3051 (N_3051,N_2895,N_2969);
xnor U3052 (N_3052,N_2936,N_2899);
or U3053 (N_3053,N_2888,N_2978);
xor U3054 (N_3054,N_2992,N_2997);
nand U3055 (N_3055,N_2971,N_2980);
and U3056 (N_3056,N_2973,N_2989);
nor U3057 (N_3057,N_2923,N_2954);
or U3058 (N_3058,N_2909,N_2960);
and U3059 (N_3059,N_2976,N_2950);
and U3060 (N_3060,N_2890,N_2996);
xnor U3061 (N_3061,N_2926,N_2920);
and U3062 (N_3062,N_2981,N_2967);
and U3063 (N_3063,N_2892,N_2878);
xor U3064 (N_3064,N_2939,N_2883);
nor U3065 (N_3065,N_2914,N_2978);
and U3066 (N_3066,N_2887,N_2993);
and U3067 (N_3067,N_2998,N_2925);
and U3068 (N_3068,N_2887,N_2952);
xnor U3069 (N_3069,N_2900,N_2934);
xor U3070 (N_3070,N_2983,N_2997);
nor U3071 (N_3071,N_2910,N_2899);
and U3072 (N_3072,N_2961,N_2877);
xor U3073 (N_3073,N_2893,N_2922);
xor U3074 (N_3074,N_2899,N_2996);
nor U3075 (N_3075,N_2949,N_2963);
and U3076 (N_3076,N_2918,N_2967);
nand U3077 (N_3077,N_2946,N_2908);
nor U3078 (N_3078,N_2969,N_2973);
and U3079 (N_3079,N_2902,N_2989);
xnor U3080 (N_3080,N_2958,N_2984);
nor U3081 (N_3081,N_2937,N_2906);
nand U3082 (N_3082,N_2977,N_2910);
and U3083 (N_3083,N_2943,N_2982);
or U3084 (N_3084,N_2910,N_2959);
nand U3085 (N_3085,N_2882,N_2955);
xnor U3086 (N_3086,N_2898,N_2949);
nand U3087 (N_3087,N_2958,N_2961);
nor U3088 (N_3088,N_2900,N_2991);
nand U3089 (N_3089,N_2930,N_2879);
or U3090 (N_3090,N_2962,N_2972);
and U3091 (N_3091,N_2945,N_2886);
xor U3092 (N_3092,N_2887,N_2955);
or U3093 (N_3093,N_2917,N_2878);
nor U3094 (N_3094,N_2886,N_2980);
nand U3095 (N_3095,N_2941,N_2903);
nor U3096 (N_3096,N_2992,N_2947);
xnor U3097 (N_3097,N_2963,N_2923);
nor U3098 (N_3098,N_2987,N_2938);
and U3099 (N_3099,N_2939,N_2926);
xor U3100 (N_3100,N_2894,N_2914);
xor U3101 (N_3101,N_2920,N_2912);
and U3102 (N_3102,N_2917,N_2896);
nor U3103 (N_3103,N_2879,N_2887);
nand U3104 (N_3104,N_2920,N_2879);
and U3105 (N_3105,N_2913,N_2881);
and U3106 (N_3106,N_2900,N_2913);
or U3107 (N_3107,N_2887,N_2973);
nor U3108 (N_3108,N_2987,N_2894);
nand U3109 (N_3109,N_2924,N_2954);
and U3110 (N_3110,N_2935,N_2996);
nand U3111 (N_3111,N_2977,N_2890);
xnor U3112 (N_3112,N_2998,N_2899);
or U3113 (N_3113,N_2901,N_2939);
nand U3114 (N_3114,N_2882,N_2960);
or U3115 (N_3115,N_2885,N_2948);
nor U3116 (N_3116,N_2939,N_2955);
xnor U3117 (N_3117,N_2894,N_2954);
nand U3118 (N_3118,N_2875,N_2912);
and U3119 (N_3119,N_2883,N_2969);
xor U3120 (N_3120,N_2880,N_2930);
nor U3121 (N_3121,N_2996,N_2897);
xor U3122 (N_3122,N_2901,N_2935);
nor U3123 (N_3123,N_2976,N_2879);
nor U3124 (N_3124,N_2919,N_2994);
and U3125 (N_3125,N_3063,N_3059);
or U3126 (N_3126,N_3010,N_3032);
or U3127 (N_3127,N_3114,N_3087);
xor U3128 (N_3128,N_3024,N_3043);
or U3129 (N_3129,N_3012,N_3061);
and U3130 (N_3130,N_3056,N_3099);
nand U3131 (N_3131,N_3121,N_3097);
or U3132 (N_3132,N_3111,N_3023);
or U3133 (N_3133,N_3051,N_3042);
nand U3134 (N_3134,N_3015,N_3106);
or U3135 (N_3135,N_3025,N_3048);
or U3136 (N_3136,N_3123,N_3054);
and U3137 (N_3137,N_3113,N_3039);
or U3138 (N_3138,N_3081,N_3008);
nor U3139 (N_3139,N_3004,N_3040);
or U3140 (N_3140,N_3072,N_3108);
and U3141 (N_3141,N_3078,N_3103);
xnor U3142 (N_3142,N_3090,N_3096);
and U3143 (N_3143,N_3016,N_3045);
nor U3144 (N_3144,N_3120,N_3058);
or U3145 (N_3145,N_3089,N_3036);
xnor U3146 (N_3146,N_3084,N_3031);
nand U3147 (N_3147,N_3022,N_3080);
or U3148 (N_3148,N_3071,N_3021);
xnor U3149 (N_3149,N_3104,N_3018);
nand U3150 (N_3150,N_3068,N_3076);
nor U3151 (N_3151,N_3067,N_3115);
nand U3152 (N_3152,N_3101,N_3073);
nand U3153 (N_3153,N_3013,N_3110);
xor U3154 (N_3154,N_3107,N_3003);
nand U3155 (N_3155,N_3086,N_3009);
or U3156 (N_3156,N_3029,N_3037);
nand U3157 (N_3157,N_3049,N_3044);
and U3158 (N_3158,N_3112,N_3124);
or U3159 (N_3159,N_3020,N_3070);
nor U3160 (N_3160,N_3069,N_3100);
and U3161 (N_3161,N_3119,N_3002);
or U3162 (N_3162,N_3006,N_3052);
or U3163 (N_3163,N_3028,N_3046);
and U3164 (N_3164,N_3053,N_3038);
or U3165 (N_3165,N_3026,N_3093);
xnor U3166 (N_3166,N_3118,N_3035);
nor U3167 (N_3167,N_3082,N_3030);
nand U3168 (N_3168,N_3083,N_3094);
and U3169 (N_3169,N_3019,N_3062);
nand U3170 (N_3170,N_3109,N_3055);
and U3171 (N_3171,N_3077,N_3095);
nand U3172 (N_3172,N_3005,N_3091);
nand U3173 (N_3173,N_3050,N_3065);
xor U3174 (N_3174,N_3057,N_3098);
or U3175 (N_3175,N_3092,N_3079);
nor U3176 (N_3176,N_3122,N_3116);
nor U3177 (N_3177,N_3047,N_3014);
nand U3178 (N_3178,N_3085,N_3001);
nand U3179 (N_3179,N_3007,N_3017);
nor U3180 (N_3180,N_3011,N_3060);
xor U3181 (N_3181,N_3102,N_3105);
or U3182 (N_3182,N_3000,N_3088);
and U3183 (N_3183,N_3117,N_3075);
nor U3184 (N_3184,N_3041,N_3066);
nor U3185 (N_3185,N_3033,N_3034);
or U3186 (N_3186,N_3064,N_3027);
xnor U3187 (N_3187,N_3074,N_3043);
xnor U3188 (N_3188,N_3017,N_3068);
or U3189 (N_3189,N_3100,N_3065);
nand U3190 (N_3190,N_3055,N_3025);
nand U3191 (N_3191,N_3013,N_3108);
nor U3192 (N_3192,N_3045,N_3047);
and U3193 (N_3193,N_3048,N_3090);
xor U3194 (N_3194,N_3010,N_3023);
nor U3195 (N_3195,N_3116,N_3028);
nand U3196 (N_3196,N_3005,N_3014);
nand U3197 (N_3197,N_3050,N_3107);
nor U3198 (N_3198,N_3065,N_3124);
xnor U3199 (N_3199,N_3045,N_3083);
xor U3200 (N_3200,N_3022,N_3010);
or U3201 (N_3201,N_3078,N_3081);
and U3202 (N_3202,N_3019,N_3021);
nand U3203 (N_3203,N_3053,N_3049);
xor U3204 (N_3204,N_3085,N_3083);
nand U3205 (N_3205,N_3119,N_3075);
nand U3206 (N_3206,N_3006,N_3095);
or U3207 (N_3207,N_3067,N_3029);
xnor U3208 (N_3208,N_3001,N_3116);
nor U3209 (N_3209,N_3068,N_3067);
or U3210 (N_3210,N_3113,N_3087);
xnor U3211 (N_3211,N_3070,N_3105);
or U3212 (N_3212,N_3032,N_3096);
xor U3213 (N_3213,N_3060,N_3036);
xor U3214 (N_3214,N_3091,N_3037);
or U3215 (N_3215,N_3086,N_3025);
nor U3216 (N_3216,N_3084,N_3019);
xnor U3217 (N_3217,N_3056,N_3047);
nand U3218 (N_3218,N_3045,N_3116);
nor U3219 (N_3219,N_3055,N_3010);
nor U3220 (N_3220,N_3091,N_3073);
and U3221 (N_3221,N_3073,N_3046);
nor U3222 (N_3222,N_3124,N_3049);
nor U3223 (N_3223,N_3007,N_3124);
xnor U3224 (N_3224,N_3061,N_3018);
xnor U3225 (N_3225,N_3111,N_3049);
nand U3226 (N_3226,N_3017,N_3122);
xor U3227 (N_3227,N_3080,N_3062);
or U3228 (N_3228,N_3108,N_3091);
nand U3229 (N_3229,N_3096,N_3046);
nor U3230 (N_3230,N_3071,N_3074);
nor U3231 (N_3231,N_3040,N_3088);
xor U3232 (N_3232,N_3119,N_3123);
nor U3233 (N_3233,N_3054,N_3056);
or U3234 (N_3234,N_3082,N_3095);
and U3235 (N_3235,N_3067,N_3100);
and U3236 (N_3236,N_3120,N_3048);
nor U3237 (N_3237,N_3083,N_3073);
xnor U3238 (N_3238,N_3073,N_3090);
xor U3239 (N_3239,N_3107,N_3055);
nor U3240 (N_3240,N_3047,N_3060);
nand U3241 (N_3241,N_3047,N_3096);
xnor U3242 (N_3242,N_3017,N_3008);
or U3243 (N_3243,N_3058,N_3051);
xor U3244 (N_3244,N_3113,N_3083);
xor U3245 (N_3245,N_3099,N_3031);
nand U3246 (N_3246,N_3115,N_3008);
or U3247 (N_3247,N_3079,N_3028);
or U3248 (N_3248,N_3046,N_3041);
xor U3249 (N_3249,N_3008,N_3070);
nor U3250 (N_3250,N_3204,N_3193);
xnor U3251 (N_3251,N_3183,N_3137);
nand U3252 (N_3252,N_3177,N_3169);
xnor U3253 (N_3253,N_3170,N_3232);
or U3254 (N_3254,N_3235,N_3218);
and U3255 (N_3255,N_3220,N_3156);
nand U3256 (N_3256,N_3141,N_3241);
or U3257 (N_3257,N_3219,N_3224);
nand U3258 (N_3258,N_3211,N_3188);
nand U3259 (N_3259,N_3228,N_3230);
nand U3260 (N_3260,N_3138,N_3209);
xnor U3261 (N_3261,N_3202,N_3179);
xor U3262 (N_3262,N_3195,N_3200);
xor U3263 (N_3263,N_3175,N_3160);
or U3264 (N_3264,N_3161,N_3237);
xor U3265 (N_3265,N_3231,N_3157);
xnor U3266 (N_3266,N_3142,N_3244);
or U3267 (N_3267,N_3171,N_3139);
nor U3268 (N_3268,N_3162,N_3143);
or U3269 (N_3269,N_3208,N_3165);
or U3270 (N_3270,N_3199,N_3242);
or U3271 (N_3271,N_3127,N_3243);
xnor U3272 (N_3272,N_3180,N_3216);
and U3273 (N_3273,N_3150,N_3197);
nand U3274 (N_3274,N_3125,N_3131);
nor U3275 (N_3275,N_3144,N_3129);
nand U3276 (N_3276,N_3155,N_3246);
xnor U3277 (N_3277,N_3163,N_3174);
and U3278 (N_3278,N_3132,N_3172);
or U3279 (N_3279,N_3210,N_3151);
and U3280 (N_3280,N_3198,N_3152);
and U3281 (N_3281,N_3203,N_3225);
nor U3282 (N_3282,N_3130,N_3215);
or U3283 (N_3283,N_3233,N_3166);
nor U3284 (N_3284,N_3217,N_3229);
or U3285 (N_3285,N_3207,N_3153);
nand U3286 (N_3286,N_3189,N_3154);
or U3287 (N_3287,N_3249,N_3159);
and U3288 (N_3288,N_3201,N_3133);
nand U3289 (N_3289,N_3181,N_3148);
xor U3290 (N_3290,N_3206,N_3136);
nor U3291 (N_3291,N_3145,N_3176);
or U3292 (N_3292,N_3158,N_3238);
xnor U3293 (N_3293,N_3146,N_3164);
xor U3294 (N_3294,N_3234,N_3227);
or U3295 (N_3295,N_3187,N_3221);
xnor U3296 (N_3296,N_3186,N_3240);
and U3297 (N_3297,N_3205,N_3167);
and U3298 (N_3298,N_3222,N_3192);
xor U3299 (N_3299,N_3213,N_3128);
and U3300 (N_3300,N_3184,N_3214);
nand U3301 (N_3301,N_3239,N_3194);
or U3302 (N_3302,N_3196,N_3212);
and U3303 (N_3303,N_3185,N_3134);
and U3304 (N_3304,N_3173,N_3140);
nand U3305 (N_3305,N_3191,N_3178);
or U3306 (N_3306,N_3226,N_3190);
or U3307 (N_3307,N_3248,N_3245);
and U3308 (N_3308,N_3147,N_3135);
nand U3309 (N_3309,N_3182,N_3126);
or U3310 (N_3310,N_3236,N_3168);
xor U3311 (N_3311,N_3149,N_3223);
xor U3312 (N_3312,N_3247,N_3240);
nor U3313 (N_3313,N_3228,N_3181);
nor U3314 (N_3314,N_3229,N_3153);
xnor U3315 (N_3315,N_3190,N_3197);
nor U3316 (N_3316,N_3199,N_3224);
and U3317 (N_3317,N_3247,N_3165);
or U3318 (N_3318,N_3196,N_3187);
nor U3319 (N_3319,N_3126,N_3234);
xnor U3320 (N_3320,N_3236,N_3176);
and U3321 (N_3321,N_3141,N_3127);
xor U3322 (N_3322,N_3159,N_3237);
and U3323 (N_3323,N_3174,N_3137);
or U3324 (N_3324,N_3229,N_3204);
nand U3325 (N_3325,N_3144,N_3184);
or U3326 (N_3326,N_3138,N_3161);
or U3327 (N_3327,N_3204,N_3178);
nand U3328 (N_3328,N_3163,N_3214);
and U3329 (N_3329,N_3248,N_3179);
xor U3330 (N_3330,N_3237,N_3178);
and U3331 (N_3331,N_3145,N_3224);
and U3332 (N_3332,N_3203,N_3142);
nand U3333 (N_3333,N_3163,N_3248);
nor U3334 (N_3334,N_3194,N_3204);
and U3335 (N_3335,N_3164,N_3196);
nand U3336 (N_3336,N_3143,N_3186);
or U3337 (N_3337,N_3194,N_3242);
nand U3338 (N_3338,N_3170,N_3129);
xor U3339 (N_3339,N_3185,N_3247);
nand U3340 (N_3340,N_3146,N_3149);
and U3341 (N_3341,N_3247,N_3141);
nor U3342 (N_3342,N_3204,N_3200);
and U3343 (N_3343,N_3227,N_3161);
or U3344 (N_3344,N_3159,N_3181);
nand U3345 (N_3345,N_3141,N_3245);
nand U3346 (N_3346,N_3208,N_3132);
nand U3347 (N_3347,N_3243,N_3141);
or U3348 (N_3348,N_3157,N_3239);
or U3349 (N_3349,N_3207,N_3166);
xor U3350 (N_3350,N_3199,N_3226);
xnor U3351 (N_3351,N_3153,N_3161);
and U3352 (N_3352,N_3130,N_3136);
and U3353 (N_3353,N_3158,N_3174);
xnor U3354 (N_3354,N_3158,N_3215);
nor U3355 (N_3355,N_3226,N_3234);
nand U3356 (N_3356,N_3153,N_3126);
nor U3357 (N_3357,N_3233,N_3182);
or U3358 (N_3358,N_3186,N_3153);
or U3359 (N_3359,N_3172,N_3208);
xnor U3360 (N_3360,N_3178,N_3242);
xor U3361 (N_3361,N_3178,N_3167);
and U3362 (N_3362,N_3138,N_3195);
xor U3363 (N_3363,N_3193,N_3224);
nand U3364 (N_3364,N_3204,N_3242);
or U3365 (N_3365,N_3162,N_3182);
and U3366 (N_3366,N_3197,N_3167);
or U3367 (N_3367,N_3231,N_3199);
nand U3368 (N_3368,N_3202,N_3130);
nand U3369 (N_3369,N_3136,N_3156);
nand U3370 (N_3370,N_3212,N_3235);
nand U3371 (N_3371,N_3204,N_3205);
or U3372 (N_3372,N_3237,N_3219);
nor U3373 (N_3373,N_3195,N_3183);
nor U3374 (N_3374,N_3228,N_3177);
and U3375 (N_3375,N_3319,N_3325);
nor U3376 (N_3376,N_3303,N_3306);
xnor U3377 (N_3377,N_3310,N_3370);
xor U3378 (N_3378,N_3294,N_3339);
xnor U3379 (N_3379,N_3374,N_3333);
and U3380 (N_3380,N_3309,N_3263);
nand U3381 (N_3381,N_3360,N_3365);
nand U3382 (N_3382,N_3335,N_3267);
xnor U3383 (N_3383,N_3350,N_3362);
and U3384 (N_3384,N_3254,N_3337);
nand U3385 (N_3385,N_3250,N_3285);
xnor U3386 (N_3386,N_3348,N_3264);
nand U3387 (N_3387,N_3274,N_3265);
and U3388 (N_3388,N_3327,N_3298);
or U3389 (N_3389,N_3353,N_3311);
xnor U3390 (N_3390,N_3367,N_3256);
and U3391 (N_3391,N_3363,N_3320);
and U3392 (N_3392,N_3347,N_3366);
or U3393 (N_3393,N_3364,N_3259);
nor U3394 (N_3394,N_3349,N_3282);
xnor U3395 (N_3395,N_3372,N_3251);
nand U3396 (N_3396,N_3359,N_3283);
or U3397 (N_3397,N_3345,N_3300);
xnor U3398 (N_3398,N_3358,N_3299);
nor U3399 (N_3399,N_3252,N_3288);
xor U3400 (N_3400,N_3290,N_3326);
nor U3401 (N_3401,N_3304,N_3322);
nand U3402 (N_3402,N_3280,N_3305);
nand U3403 (N_3403,N_3293,N_3281);
nor U3404 (N_3404,N_3271,N_3273);
and U3405 (N_3405,N_3352,N_3361);
and U3406 (N_3406,N_3276,N_3357);
nand U3407 (N_3407,N_3255,N_3344);
xor U3408 (N_3408,N_3278,N_3279);
xnor U3409 (N_3409,N_3307,N_3253);
nand U3410 (N_3410,N_3296,N_3346);
or U3411 (N_3411,N_3277,N_3284);
nand U3412 (N_3412,N_3341,N_3261);
nor U3413 (N_3413,N_3287,N_3330);
nor U3414 (N_3414,N_3340,N_3258);
nor U3415 (N_3415,N_3338,N_3371);
or U3416 (N_3416,N_3354,N_3272);
and U3417 (N_3417,N_3329,N_3356);
or U3418 (N_3418,N_3302,N_3291);
xnor U3419 (N_3419,N_3324,N_3336);
and U3420 (N_3420,N_3295,N_3343);
xor U3421 (N_3421,N_3316,N_3334);
or U3422 (N_3422,N_3257,N_3317);
xor U3423 (N_3423,N_3351,N_3313);
or U3424 (N_3424,N_3342,N_3260);
xor U3425 (N_3425,N_3301,N_3331);
nor U3426 (N_3426,N_3373,N_3355);
nand U3427 (N_3427,N_3289,N_3315);
nor U3428 (N_3428,N_3318,N_3308);
or U3429 (N_3429,N_3262,N_3312);
or U3430 (N_3430,N_3268,N_3328);
or U3431 (N_3431,N_3297,N_3314);
or U3432 (N_3432,N_3275,N_3292);
nand U3433 (N_3433,N_3323,N_3369);
nand U3434 (N_3434,N_3332,N_3270);
or U3435 (N_3435,N_3321,N_3269);
nor U3436 (N_3436,N_3266,N_3286);
nand U3437 (N_3437,N_3368,N_3361);
nor U3438 (N_3438,N_3325,N_3357);
xor U3439 (N_3439,N_3349,N_3295);
nor U3440 (N_3440,N_3265,N_3331);
xnor U3441 (N_3441,N_3315,N_3317);
nand U3442 (N_3442,N_3286,N_3264);
or U3443 (N_3443,N_3323,N_3373);
nand U3444 (N_3444,N_3302,N_3331);
nand U3445 (N_3445,N_3291,N_3333);
xor U3446 (N_3446,N_3339,N_3261);
or U3447 (N_3447,N_3260,N_3353);
nand U3448 (N_3448,N_3287,N_3338);
nand U3449 (N_3449,N_3349,N_3289);
nor U3450 (N_3450,N_3341,N_3265);
and U3451 (N_3451,N_3345,N_3325);
xnor U3452 (N_3452,N_3343,N_3319);
or U3453 (N_3453,N_3355,N_3344);
nor U3454 (N_3454,N_3358,N_3301);
nor U3455 (N_3455,N_3254,N_3280);
and U3456 (N_3456,N_3330,N_3374);
nand U3457 (N_3457,N_3261,N_3313);
nand U3458 (N_3458,N_3332,N_3307);
nand U3459 (N_3459,N_3288,N_3308);
or U3460 (N_3460,N_3277,N_3294);
nor U3461 (N_3461,N_3308,N_3333);
nor U3462 (N_3462,N_3332,N_3271);
nor U3463 (N_3463,N_3262,N_3365);
and U3464 (N_3464,N_3347,N_3294);
or U3465 (N_3465,N_3324,N_3279);
nand U3466 (N_3466,N_3354,N_3307);
xor U3467 (N_3467,N_3344,N_3341);
and U3468 (N_3468,N_3332,N_3315);
or U3469 (N_3469,N_3252,N_3316);
nor U3470 (N_3470,N_3308,N_3369);
xnor U3471 (N_3471,N_3355,N_3295);
and U3472 (N_3472,N_3254,N_3304);
and U3473 (N_3473,N_3355,N_3345);
xor U3474 (N_3474,N_3334,N_3290);
nor U3475 (N_3475,N_3343,N_3287);
nand U3476 (N_3476,N_3340,N_3311);
xor U3477 (N_3477,N_3276,N_3363);
or U3478 (N_3478,N_3264,N_3326);
nand U3479 (N_3479,N_3361,N_3274);
nor U3480 (N_3480,N_3252,N_3264);
or U3481 (N_3481,N_3275,N_3354);
nor U3482 (N_3482,N_3302,N_3325);
nand U3483 (N_3483,N_3368,N_3286);
or U3484 (N_3484,N_3264,N_3323);
nand U3485 (N_3485,N_3269,N_3275);
xor U3486 (N_3486,N_3319,N_3334);
nand U3487 (N_3487,N_3302,N_3369);
xor U3488 (N_3488,N_3278,N_3352);
nor U3489 (N_3489,N_3260,N_3320);
nor U3490 (N_3490,N_3338,N_3254);
nand U3491 (N_3491,N_3371,N_3265);
or U3492 (N_3492,N_3299,N_3286);
nor U3493 (N_3493,N_3319,N_3335);
xor U3494 (N_3494,N_3331,N_3342);
nor U3495 (N_3495,N_3295,N_3350);
and U3496 (N_3496,N_3353,N_3363);
or U3497 (N_3497,N_3326,N_3355);
xor U3498 (N_3498,N_3252,N_3258);
nand U3499 (N_3499,N_3355,N_3364);
or U3500 (N_3500,N_3382,N_3440);
and U3501 (N_3501,N_3402,N_3396);
nor U3502 (N_3502,N_3496,N_3410);
and U3503 (N_3503,N_3457,N_3376);
nand U3504 (N_3504,N_3487,N_3407);
nand U3505 (N_3505,N_3381,N_3392);
nor U3506 (N_3506,N_3375,N_3405);
xnor U3507 (N_3507,N_3425,N_3483);
or U3508 (N_3508,N_3434,N_3435);
or U3509 (N_3509,N_3436,N_3437);
nand U3510 (N_3510,N_3471,N_3426);
xor U3511 (N_3511,N_3445,N_3386);
or U3512 (N_3512,N_3474,N_3400);
or U3513 (N_3513,N_3384,N_3442);
or U3514 (N_3514,N_3422,N_3447);
nor U3515 (N_3515,N_3419,N_3395);
and U3516 (N_3516,N_3476,N_3462);
nor U3517 (N_3517,N_3473,N_3461);
xnor U3518 (N_3518,N_3497,N_3411);
nand U3519 (N_3519,N_3499,N_3421);
or U3520 (N_3520,N_3492,N_3469);
nand U3521 (N_3521,N_3482,N_3401);
xor U3522 (N_3522,N_3423,N_3478);
nor U3523 (N_3523,N_3387,N_3417);
xnor U3524 (N_3524,N_3488,N_3472);
nand U3525 (N_3525,N_3413,N_3439);
nand U3526 (N_3526,N_3416,N_3463);
nand U3527 (N_3527,N_3390,N_3491);
nand U3528 (N_3528,N_3451,N_3412);
nor U3529 (N_3529,N_3427,N_3409);
nand U3530 (N_3530,N_3383,N_3475);
or U3531 (N_3531,N_3430,N_3385);
or U3532 (N_3532,N_3438,N_3446);
or U3533 (N_3533,N_3399,N_3397);
xor U3534 (N_3534,N_3432,N_3398);
xnor U3535 (N_3535,N_3444,N_3467);
and U3536 (N_3536,N_3489,N_3403);
xnor U3537 (N_3537,N_3486,N_3393);
nand U3538 (N_3538,N_3480,N_3408);
and U3539 (N_3539,N_3441,N_3453);
or U3540 (N_3540,N_3428,N_3468);
and U3541 (N_3541,N_3443,N_3394);
nand U3542 (N_3542,N_3490,N_3459);
nand U3543 (N_3543,N_3378,N_3477);
xor U3544 (N_3544,N_3494,N_3388);
xor U3545 (N_3545,N_3498,N_3470);
or U3546 (N_3546,N_3433,N_3456);
nand U3547 (N_3547,N_3420,N_3404);
or U3548 (N_3548,N_3415,N_3418);
xnor U3549 (N_3549,N_3458,N_3485);
xnor U3550 (N_3550,N_3414,N_3380);
and U3551 (N_3551,N_3379,N_3484);
nor U3552 (N_3552,N_3460,N_3448);
or U3553 (N_3553,N_3406,N_3464);
nand U3554 (N_3554,N_3481,N_3454);
xor U3555 (N_3555,N_3424,N_3493);
and U3556 (N_3556,N_3452,N_3495);
or U3557 (N_3557,N_3431,N_3391);
xor U3558 (N_3558,N_3479,N_3465);
nor U3559 (N_3559,N_3377,N_3466);
xor U3560 (N_3560,N_3449,N_3429);
xor U3561 (N_3561,N_3450,N_3389);
or U3562 (N_3562,N_3455,N_3406);
or U3563 (N_3563,N_3394,N_3390);
nor U3564 (N_3564,N_3395,N_3464);
xnor U3565 (N_3565,N_3402,N_3413);
nor U3566 (N_3566,N_3441,N_3406);
nand U3567 (N_3567,N_3467,N_3494);
xor U3568 (N_3568,N_3378,N_3396);
xnor U3569 (N_3569,N_3433,N_3487);
nand U3570 (N_3570,N_3492,N_3437);
xor U3571 (N_3571,N_3376,N_3467);
and U3572 (N_3572,N_3465,N_3475);
nand U3573 (N_3573,N_3462,N_3432);
nand U3574 (N_3574,N_3383,N_3392);
xnor U3575 (N_3575,N_3452,N_3479);
and U3576 (N_3576,N_3482,N_3477);
or U3577 (N_3577,N_3493,N_3414);
and U3578 (N_3578,N_3405,N_3455);
and U3579 (N_3579,N_3469,N_3385);
xnor U3580 (N_3580,N_3491,N_3386);
nor U3581 (N_3581,N_3496,N_3444);
nand U3582 (N_3582,N_3406,N_3388);
nand U3583 (N_3583,N_3448,N_3440);
xor U3584 (N_3584,N_3463,N_3378);
and U3585 (N_3585,N_3397,N_3425);
and U3586 (N_3586,N_3399,N_3438);
and U3587 (N_3587,N_3422,N_3431);
and U3588 (N_3588,N_3473,N_3377);
or U3589 (N_3589,N_3487,N_3471);
xnor U3590 (N_3590,N_3456,N_3473);
nand U3591 (N_3591,N_3410,N_3453);
nand U3592 (N_3592,N_3402,N_3427);
nor U3593 (N_3593,N_3448,N_3489);
nand U3594 (N_3594,N_3441,N_3419);
and U3595 (N_3595,N_3426,N_3474);
xnor U3596 (N_3596,N_3375,N_3435);
nand U3597 (N_3597,N_3435,N_3462);
nand U3598 (N_3598,N_3390,N_3393);
or U3599 (N_3599,N_3473,N_3381);
xor U3600 (N_3600,N_3439,N_3442);
nand U3601 (N_3601,N_3398,N_3485);
or U3602 (N_3602,N_3467,N_3498);
nor U3603 (N_3603,N_3429,N_3416);
or U3604 (N_3604,N_3481,N_3399);
nand U3605 (N_3605,N_3494,N_3413);
nand U3606 (N_3606,N_3423,N_3421);
nor U3607 (N_3607,N_3494,N_3400);
nor U3608 (N_3608,N_3397,N_3454);
or U3609 (N_3609,N_3413,N_3422);
xnor U3610 (N_3610,N_3386,N_3468);
xor U3611 (N_3611,N_3471,N_3466);
nand U3612 (N_3612,N_3397,N_3474);
and U3613 (N_3613,N_3423,N_3496);
nor U3614 (N_3614,N_3417,N_3423);
nor U3615 (N_3615,N_3466,N_3434);
and U3616 (N_3616,N_3404,N_3391);
and U3617 (N_3617,N_3388,N_3391);
nand U3618 (N_3618,N_3484,N_3390);
nor U3619 (N_3619,N_3473,N_3380);
nand U3620 (N_3620,N_3485,N_3455);
nor U3621 (N_3621,N_3408,N_3432);
or U3622 (N_3622,N_3493,N_3492);
nor U3623 (N_3623,N_3481,N_3396);
and U3624 (N_3624,N_3452,N_3489);
nand U3625 (N_3625,N_3548,N_3571);
xnor U3626 (N_3626,N_3522,N_3608);
or U3627 (N_3627,N_3524,N_3540);
or U3628 (N_3628,N_3563,N_3566);
and U3629 (N_3629,N_3557,N_3618);
or U3630 (N_3630,N_3588,N_3550);
nand U3631 (N_3631,N_3546,N_3526);
nor U3632 (N_3632,N_3518,N_3619);
or U3633 (N_3633,N_3601,N_3511);
or U3634 (N_3634,N_3572,N_3542);
and U3635 (N_3635,N_3504,N_3575);
or U3636 (N_3636,N_3544,N_3529);
xnor U3637 (N_3637,N_3613,N_3609);
nand U3638 (N_3638,N_3584,N_3611);
nand U3639 (N_3639,N_3622,N_3545);
nor U3640 (N_3640,N_3620,N_3586);
xor U3641 (N_3641,N_3594,N_3505);
nand U3642 (N_3642,N_3587,N_3607);
and U3643 (N_3643,N_3585,N_3541);
and U3644 (N_3644,N_3614,N_3556);
xnor U3645 (N_3645,N_3503,N_3583);
xor U3646 (N_3646,N_3606,N_3502);
nand U3647 (N_3647,N_3532,N_3576);
or U3648 (N_3648,N_3543,N_3558);
nand U3649 (N_3649,N_3580,N_3577);
and U3650 (N_3650,N_3510,N_3514);
and U3651 (N_3651,N_3509,N_3617);
nor U3652 (N_3652,N_3501,N_3589);
and U3653 (N_3653,N_3554,N_3567);
xor U3654 (N_3654,N_3590,N_3570);
nor U3655 (N_3655,N_3561,N_3531);
nand U3656 (N_3656,N_3528,N_3621);
xor U3657 (N_3657,N_3506,N_3535);
nand U3658 (N_3658,N_3530,N_3592);
or U3659 (N_3659,N_3536,N_3515);
nand U3660 (N_3660,N_3539,N_3598);
xor U3661 (N_3661,N_3547,N_3565);
xor U3662 (N_3662,N_3600,N_3537);
nor U3663 (N_3663,N_3521,N_3624);
nand U3664 (N_3664,N_3562,N_3623);
or U3665 (N_3665,N_3605,N_3612);
nand U3666 (N_3666,N_3516,N_3602);
or U3667 (N_3667,N_3593,N_3596);
nand U3668 (N_3668,N_3552,N_3508);
or U3669 (N_3669,N_3500,N_3573);
nor U3670 (N_3670,N_3604,N_3538);
or U3671 (N_3671,N_3569,N_3581);
nand U3672 (N_3672,N_3603,N_3553);
xor U3673 (N_3673,N_3560,N_3512);
xnor U3674 (N_3674,N_3551,N_3610);
nor U3675 (N_3675,N_3579,N_3507);
nor U3676 (N_3676,N_3595,N_3527);
and U3677 (N_3677,N_3520,N_3615);
xnor U3678 (N_3678,N_3523,N_3568);
and U3679 (N_3679,N_3564,N_3533);
or U3680 (N_3680,N_3582,N_3559);
nand U3681 (N_3681,N_3616,N_3519);
or U3682 (N_3682,N_3513,N_3555);
nor U3683 (N_3683,N_3597,N_3525);
nor U3684 (N_3684,N_3591,N_3534);
and U3685 (N_3685,N_3574,N_3599);
nor U3686 (N_3686,N_3517,N_3578);
xnor U3687 (N_3687,N_3549,N_3514);
nand U3688 (N_3688,N_3516,N_3567);
xor U3689 (N_3689,N_3547,N_3557);
and U3690 (N_3690,N_3603,N_3584);
and U3691 (N_3691,N_3529,N_3535);
and U3692 (N_3692,N_3603,N_3581);
nand U3693 (N_3693,N_3551,N_3569);
nor U3694 (N_3694,N_3546,N_3613);
and U3695 (N_3695,N_3543,N_3540);
nor U3696 (N_3696,N_3512,N_3596);
xnor U3697 (N_3697,N_3528,N_3537);
xnor U3698 (N_3698,N_3545,N_3564);
and U3699 (N_3699,N_3595,N_3533);
or U3700 (N_3700,N_3573,N_3612);
nand U3701 (N_3701,N_3564,N_3539);
xor U3702 (N_3702,N_3513,N_3620);
and U3703 (N_3703,N_3522,N_3513);
or U3704 (N_3704,N_3543,N_3565);
nand U3705 (N_3705,N_3585,N_3595);
and U3706 (N_3706,N_3507,N_3557);
and U3707 (N_3707,N_3587,N_3535);
nand U3708 (N_3708,N_3578,N_3583);
and U3709 (N_3709,N_3554,N_3551);
and U3710 (N_3710,N_3501,N_3616);
xnor U3711 (N_3711,N_3564,N_3507);
xor U3712 (N_3712,N_3558,N_3555);
or U3713 (N_3713,N_3600,N_3615);
nand U3714 (N_3714,N_3570,N_3532);
nand U3715 (N_3715,N_3608,N_3599);
and U3716 (N_3716,N_3519,N_3591);
or U3717 (N_3717,N_3518,N_3555);
or U3718 (N_3718,N_3538,N_3533);
nor U3719 (N_3719,N_3564,N_3561);
or U3720 (N_3720,N_3600,N_3562);
or U3721 (N_3721,N_3502,N_3563);
and U3722 (N_3722,N_3592,N_3513);
or U3723 (N_3723,N_3541,N_3582);
and U3724 (N_3724,N_3604,N_3581);
or U3725 (N_3725,N_3600,N_3545);
nand U3726 (N_3726,N_3538,N_3558);
nand U3727 (N_3727,N_3591,N_3589);
and U3728 (N_3728,N_3502,N_3501);
or U3729 (N_3729,N_3512,N_3612);
nand U3730 (N_3730,N_3532,N_3609);
nor U3731 (N_3731,N_3546,N_3519);
nor U3732 (N_3732,N_3502,N_3623);
and U3733 (N_3733,N_3541,N_3505);
nand U3734 (N_3734,N_3572,N_3545);
and U3735 (N_3735,N_3605,N_3520);
xnor U3736 (N_3736,N_3594,N_3554);
or U3737 (N_3737,N_3580,N_3526);
nor U3738 (N_3738,N_3510,N_3554);
xnor U3739 (N_3739,N_3597,N_3510);
and U3740 (N_3740,N_3553,N_3532);
nand U3741 (N_3741,N_3565,N_3568);
and U3742 (N_3742,N_3557,N_3553);
and U3743 (N_3743,N_3577,N_3562);
nor U3744 (N_3744,N_3541,N_3522);
nand U3745 (N_3745,N_3504,N_3508);
nand U3746 (N_3746,N_3590,N_3562);
or U3747 (N_3747,N_3542,N_3552);
xnor U3748 (N_3748,N_3522,N_3606);
and U3749 (N_3749,N_3581,N_3545);
xnor U3750 (N_3750,N_3682,N_3680);
nand U3751 (N_3751,N_3709,N_3632);
nand U3752 (N_3752,N_3696,N_3693);
and U3753 (N_3753,N_3625,N_3719);
nand U3754 (N_3754,N_3729,N_3738);
nand U3755 (N_3755,N_3722,N_3698);
xor U3756 (N_3756,N_3646,N_3645);
nand U3757 (N_3757,N_3674,N_3748);
nand U3758 (N_3758,N_3715,N_3639);
nand U3759 (N_3759,N_3660,N_3666);
and U3760 (N_3760,N_3627,N_3692);
xnor U3761 (N_3761,N_3725,N_3676);
or U3762 (N_3762,N_3655,N_3626);
or U3763 (N_3763,N_3695,N_3665);
and U3764 (N_3764,N_3651,N_3683);
xnor U3765 (N_3765,N_3747,N_3737);
xor U3766 (N_3766,N_3721,N_3629);
nor U3767 (N_3767,N_3732,N_3647);
or U3768 (N_3768,N_3700,N_3642);
nand U3769 (N_3769,N_3749,N_3713);
nor U3770 (N_3770,N_3652,N_3689);
or U3771 (N_3771,N_3703,N_3649);
nor U3772 (N_3772,N_3728,N_3740);
nor U3773 (N_3773,N_3662,N_3672);
and U3774 (N_3774,N_3650,N_3681);
nand U3775 (N_3775,N_3744,N_3708);
nand U3776 (N_3776,N_3668,N_3677);
nand U3777 (N_3777,N_3685,N_3658);
nand U3778 (N_3778,N_3720,N_3630);
xnor U3779 (N_3779,N_3712,N_3741);
or U3780 (N_3780,N_3691,N_3697);
nand U3781 (N_3781,N_3684,N_3631);
nand U3782 (N_3782,N_3730,N_3717);
nor U3783 (N_3783,N_3669,N_3694);
and U3784 (N_3784,N_3742,N_3727);
nor U3785 (N_3785,N_3688,N_3637);
nand U3786 (N_3786,N_3648,N_3710);
or U3787 (N_3787,N_3745,N_3656);
nor U3788 (N_3788,N_3714,N_3699);
nor U3789 (N_3789,N_3739,N_3663);
or U3790 (N_3790,N_3657,N_3690);
xnor U3791 (N_3791,N_3736,N_3675);
and U3792 (N_3792,N_3653,N_3686);
nor U3793 (N_3793,N_3726,N_3743);
nand U3794 (N_3794,N_3679,N_3678);
xor U3795 (N_3795,N_3705,N_3733);
or U3796 (N_3796,N_3661,N_3635);
and U3797 (N_3797,N_3659,N_3735);
xor U3798 (N_3798,N_3724,N_3641);
nand U3799 (N_3799,N_3640,N_3654);
and U3800 (N_3800,N_3734,N_3638);
and U3801 (N_3801,N_3701,N_3664);
or U3802 (N_3802,N_3706,N_3687);
xnor U3803 (N_3803,N_3723,N_3702);
and U3804 (N_3804,N_3673,N_3746);
nor U3805 (N_3805,N_3636,N_3711);
xnor U3806 (N_3806,N_3716,N_3671);
nor U3807 (N_3807,N_3633,N_3731);
nor U3808 (N_3808,N_3644,N_3704);
and U3809 (N_3809,N_3707,N_3634);
nand U3810 (N_3810,N_3667,N_3718);
nand U3811 (N_3811,N_3670,N_3628);
and U3812 (N_3812,N_3643,N_3631);
or U3813 (N_3813,N_3660,N_3722);
nand U3814 (N_3814,N_3696,N_3747);
or U3815 (N_3815,N_3647,N_3748);
xnor U3816 (N_3816,N_3667,N_3699);
or U3817 (N_3817,N_3682,N_3695);
or U3818 (N_3818,N_3702,N_3716);
xnor U3819 (N_3819,N_3645,N_3652);
or U3820 (N_3820,N_3655,N_3651);
and U3821 (N_3821,N_3739,N_3705);
nand U3822 (N_3822,N_3707,N_3697);
xor U3823 (N_3823,N_3642,N_3691);
or U3824 (N_3824,N_3701,N_3681);
nand U3825 (N_3825,N_3628,N_3707);
xor U3826 (N_3826,N_3665,N_3659);
or U3827 (N_3827,N_3662,N_3637);
xnor U3828 (N_3828,N_3655,N_3705);
or U3829 (N_3829,N_3700,N_3693);
nor U3830 (N_3830,N_3687,N_3713);
nand U3831 (N_3831,N_3666,N_3725);
or U3832 (N_3832,N_3672,N_3689);
xnor U3833 (N_3833,N_3702,N_3674);
nand U3834 (N_3834,N_3653,N_3626);
nor U3835 (N_3835,N_3664,N_3725);
nand U3836 (N_3836,N_3668,N_3650);
nor U3837 (N_3837,N_3677,N_3699);
or U3838 (N_3838,N_3733,N_3708);
nand U3839 (N_3839,N_3638,N_3685);
or U3840 (N_3840,N_3626,N_3656);
nand U3841 (N_3841,N_3659,N_3655);
or U3842 (N_3842,N_3735,N_3683);
nand U3843 (N_3843,N_3638,N_3725);
nor U3844 (N_3844,N_3655,N_3665);
nor U3845 (N_3845,N_3657,N_3671);
and U3846 (N_3846,N_3650,N_3710);
nand U3847 (N_3847,N_3731,N_3737);
and U3848 (N_3848,N_3725,N_3660);
and U3849 (N_3849,N_3636,N_3680);
and U3850 (N_3850,N_3636,N_3709);
nor U3851 (N_3851,N_3652,N_3701);
or U3852 (N_3852,N_3659,N_3698);
and U3853 (N_3853,N_3653,N_3735);
xnor U3854 (N_3854,N_3656,N_3627);
nor U3855 (N_3855,N_3746,N_3667);
nor U3856 (N_3856,N_3655,N_3722);
xor U3857 (N_3857,N_3701,N_3684);
and U3858 (N_3858,N_3682,N_3697);
nand U3859 (N_3859,N_3703,N_3728);
nor U3860 (N_3860,N_3668,N_3715);
nor U3861 (N_3861,N_3630,N_3717);
xor U3862 (N_3862,N_3747,N_3713);
xor U3863 (N_3863,N_3723,N_3650);
nor U3864 (N_3864,N_3638,N_3626);
or U3865 (N_3865,N_3725,N_3702);
xnor U3866 (N_3866,N_3740,N_3627);
and U3867 (N_3867,N_3703,N_3654);
and U3868 (N_3868,N_3688,N_3747);
and U3869 (N_3869,N_3695,N_3701);
nor U3870 (N_3870,N_3649,N_3659);
xor U3871 (N_3871,N_3746,N_3664);
nand U3872 (N_3872,N_3644,N_3706);
nand U3873 (N_3873,N_3648,N_3652);
and U3874 (N_3874,N_3651,N_3668);
or U3875 (N_3875,N_3819,N_3848);
xor U3876 (N_3876,N_3761,N_3872);
xnor U3877 (N_3877,N_3844,N_3771);
nand U3878 (N_3878,N_3852,N_3816);
and U3879 (N_3879,N_3784,N_3799);
nor U3880 (N_3880,N_3811,N_3763);
xor U3881 (N_3881,N_3766,N_3830);
and U3882 (N_3882,N_3792,N_3756);
and U3883 (N_3883,N_3822,N_3793);
nor U3884 (N_3884,N_3812,N_3788);
nand U3885 (N_3885,N_3754,N_3873);
and U3886 (N_3886,N_3858,N_3828);
and U3887 (N_3887,N_3800,N_3791);
nand U3888 (N_3888,N_3757,N_3751);
nor U3889 (N_3889,N_3846,N_3772);
and U3890 (N_3890,N_3866,N_3758);
xnor U3891 (N_3891,N_3820,N_3854);
nand U3892 (N_3892,N_3836,N_3839);
and U3893 (N_3893,N_3868,N_3805);
nand U3894 (N_3894,N_3831,N_3871);
nor U3895 (N_3895,N_3856,N_3834);
nand U3896 (N_3896,N_3825,N_3759);
nand U3897 (N_3897,N_3808,N_3835);
nor U3898 (N_3898,N_3794,N_3752);
and U3899 (N_3899,N_3795,N_3774);
xor U3900 (N_3900,N_3797,N_3859);
nor U3901 (N_3901,N_3764,N_3860);
nor U3902 (N_3902,N_3760,N_3832);
and U3903 (N_3903,N_3787,N_3806);
and U3904 (N_3904,N_3777,N_3775);
nor U3905 (N_3905,N_3804,N_3865);
nor U3906 (N_3906,N_3807,N_3818);
and U3907 (N_3907,N_3769,N_3826);
and U3908 (N_3908,N_3801,N_3855);
nand U3909 (N_3909,N_3796,N_3850);
nand U3910 (N_3910,N_3845,N_3778);
nor U3911 (N_3911,N_3841,N_3861);
and U3912 (N_3912,N_3765,N_3780);
and U3913 (N_3913,N_3814,N_3842);
xnor U3914 (N_3914,N_3829,N_3862);
nand U3915 (N_3915,N_3767,N_3870);
xor U3916 (N_3916,N_3782,N_3867);
nor U3917 (N_3917,N_3790,N_3849);
xnor U3918 (N_3918,N_3810,N_3789);
or U3919 (N_3919,N_3770,N_3864);
nand U3920 (N_3920,N_3798,N_3750);
and U3921 (N_3921,N_3773,N_3874);
or U3922 (N_3922,N_3869,N_3853);
or U3923 (N_3923,N_3857,N_3813);
nor U3924 (N_3924,N_3753,N_3833);
nor U3925 (N_3925,N_3851,N_3815);
or U3926 (N_3926,N_3863,N_3768);
or U3927 (N_3927,N_3783,N_3824);
and U3928 (N_3928,N_3843,N_3817);
nor U3929 (N_3929,N_3762,N_3827);
or U3930 (N_3930,N_3776,N_3838);
and U3931 (N_3931,N_3785,N_3803);
nor U3932 (N_3932,N_3802,N_3821);
or U3933 (N_3933,N_3781,N_3840);
xnor U3934 (N_3934,N_3779,N_3823);
and U3935 (N_3935,N_3809,N_3847);
xor U3936 (N_3936,N_3786,N_3755);
nand U3937 (N_3937,N_3837,N_3813);
xnor U3938 (N_3938,N_3840,N_3792);
and U3939 (N_3939,N_3831,N_3759);
or U3940 (N_3940,N_3783,N_3804);
nand U3941 (N_3941,N_3848,N_3774);
and U3942 (N_3942,N_3868,N_3803);
nand U3943 (N_3943,N_3849,N_3760);
nor U3944 (N_3944,N_3801,N_3774);
nor U3945 (N_3945,N_3830,N_3761);
nand U3946 (N_3946,N_3871,N_3776);
xor U3947 (N_3947,N_3867,N_3854);
nor U3948 (N_3948,N_3839,N_3754);
xor U3949 (N_3949,N_3844,N_3799);
nand U3950 (N_3950,N_3858,N_3817);
or U3951 (N_3951,N_3837,N_3829);
and U3952 (N_3952,N_3820,N_3826);
nor U3953 (N_3953,N_3801,N_3836);
or U3954 (N_3954,N_3800,N_3823);
and U3955 (N_3955,N_3869,N_3864);
nor U3956 (N_3956,N_3770,N_3818);
nand U3957 (N_3957,N_3754,N_3838);
nor U3958 (N_3958,N_3774,N_3822);
nand U3959 (N_3959,N_3874,N_3786);
nand U3960 (N_3960,N_3806,N_3846);
nor U3961 (N_3961,N_3844,N_3770);
nor U3962 (N_3962,N_3798,N_3827);
xor U3963 (N_3963,N_3783,N_3851);
or U3964 (N_3964,N_3808,N_3821);
xor U3965 (N_3965,N_3800,N_3793);
nor U3966 (N_3966,N_3805,N_3814);
nor U3967 (N_3967,N_3840,N_3751);
or U3968 (N_3968,N_3824,N_3752);
nand U3969 (N_3969,N_3844,N_3793);
nor U3970 (N_3970,N_3857,N_3864);
and U3971 (N_3971,N_3840,N_3771);
nand U3972 (N_3972,N_3836,N_3855);
nand U3973 (N_3973,N_3827,N_3752);
nand U3974 (N_3974,N_3823,N_3788);
or U3975 (N_3975,N_3753,N_3809);
nand U3976 (N_3976,N_3771,N_3828);
nand U3977 (N_3977,N_3772,N_3850);
or U3978 (N_3978,N_3783,N_3753);
and U3979 (N_3979,N_3832,N_3802);
xnor U3980 (N_3980,N_3772,N_3812);
xor U3981 (N_3981,N_3793,N_3796);
nand U3982 (N_3982,N_3777,N_3860);
and U3983 (N_3983,N_3837,N_3842);
nand U3984 (N_3984,N_3770,N_3837);
xnor U3985 (N_3985,N_3755,N_3817);
and U3986 (N_3986,N_3827,N_3859);
nor U3987 (N_3987,N_3750,N_3820);
nor U3988 (N_3988,N_3808,N_3872);
and U3989 (N_3989,N_3829,N_3842);
or U3990 (N_3990,N_3847,N_3782);
or U3991 (N_3991,N_3802,N_3814);
and U3992 (N_3992,N_3822,N_3776);
xor U3993 (N_3993,N_3819,N_3843);
and U3994 (N_3994,N_3853,N_3757);
nand U3995 (N_3995,N_3874,N_3799);
and U3996 (N_3996,N_3804,N_3820);
or U3997 (N_3997,N_3756,N_3847);
xor U3998 (N_3998,N_3811,N_3770);
xor U3999 (N_3999,N_3835,N_3829);
nor U4000 (N_4000,N_3976,N_3983);
or U4001 (N_4001,N_3914,N_3919);
xor U4002 (N_4002,N_3964,N_3945);
nor U4003 (N_4003,N_3920,N_3879);
xor U4004 (N_4004,N_3877,N_3924);
nand U4005 (N_4005,N_3882,N_3990);
nor U4006 (N_4006,N_3997,N_3881);
or U4007 (N_4007,N_3939,N_3986);
nor U4008 (N_4008,N_3876,N_3937);
nand U4009 (N_4009,N_3903,N_3984);
nand U4010 (N_4010,N_3890,N_3940);
and U4011 (N_4011,N_3893,N_3958);
or U4012 (N_4012,N_3910,N_3948);
nor U4013 (N_4013,N_3951,N_3975);
nand U4014 (N_4014,N_3973,N_3956);
xor U4015 (N_4015,N_3918,N_3899);
nor U4016 (N_4016,N_3957,N_3929);
nand U4017 (N_4017,N_3921,N_3993);
nor U4018 (N_4018,N_3944,N_3901);
nor U4019 (N_4019,N_3988,N_3889);
xnor U4020 (N_4020,N_3972,N_3908);
nor U4021 (N_4021,N_3992,N_3917);
nor U4022 (N_4022,N_3911,N_3902);
xor U4023 (N_4023,N_3947,N_3935);
and U4024 (N_4024,N_3915,N_3966);
and U4025 (N_4025,N_3878,N_3894);
xnor U4026 (N_4026,N_3989,N_3967);
xor U4027 (N_4027,N_3965,N_3938);
nand U4028 (N_4028,N_3922,N_3886);
xnor U4029 (N_4029,N_3905,N_3960);
nor U4030 (N_4030,N_3934,N_3946);
xnor U4031 (N_4031,N_3981,N_3875);
and U4032 (N_4032,N_3994,N_3883);
or U4033 (N_4033,N_3880,N_3971);
or U4034 (N_4034,N_3931,N_3950);
nand U4035 (N_4035,N_3932,N_3979);
xnor U4036 (N_4036,N_3904,N_3927);
or U4037 (N_4037,N_3916,N_3985);
xor U4038 (N_4038,N_3978,N_3962);
and U4039 (N_4039,N_3952,N_3930);
nor U4040 (N_4040,N_3923,N_3996);
and U4041 (N_4041,N_3961,N_3888);
nor U4042 (N_4042,N_3898,N_3959);
and U4043 (N_4043,N_3926,N_3963);
or U4044 (N_4044,N_3955,N_3912);
nor U4045 (N_4045,N_3942,N_3900);
and U4046 (N_4046,N_3954,N_3887);
or U4047 (N_4047,N_3892,N_3896);
or U4048 (N_4048,N_3982,N_3977);
and U4049 (N_4049,N_3895,N_3925);
xnor U4050 (N_4050,N_3995,N_3891);
nand U4051 (N_4051,N_3991,N_3933);
nor U4052 (N_4052,N_3987,N_3906);
or U4053 (N_4053,N_3907,N_3897);
xnor U4054 (N_4054,N_3968,N_3998);
and U4055 (N_4055,N_3936,N_3974);
nor U4056 (N_4056,N_3999,N_3970);
or U4057 (N_4057,N_3909,N_3943);
nor U4058 (N_4058,N_3885,N_3949);
and U4059 (N_4059,N_3884,N_3980);
and U4060 (N_4060,N_3913,N_3969);
and U4061 (N_4061,N_3928,N_3953);
xor U4062 (N_4062,N_3941,N_3888);
and U4063 (N_4063,N_3922,N_3929);
xor U4064 (N_4064,N_3917,N_3881);
nor U4065 (N_4065,N_3927,N_3906);
xor U4066 (N_4066,N_3980,N_3885);
or U4067 (N_4067,N_3995,N_3973);
or U4068 (N_4068,N_3913,N_3925);
and U4069 (N_4069,N_3969,N_3945);
and U4070 (N_4070,N_3991,N_3880);
nand U4071 (N_4071,N_3896,N_3906);
nor U4072 (N_4072,N_3898,N_3974);
or U4073 (N_4073,N_3902,N_3949);
nand U4074 (N_4074,N_3992,N_3961);
nand U4075 (N_4075,N_3986,N_3922);
nand U4076 (N_4076,N_3911,N_3946);
nand U4077 (N_4077,N_3876,N_3961);
nor U4078 (N_4078,N_3925,N_3927);
nor U4079 (N_4079,N_3983,N_3881);
nor U4080 (N_4080,N_3962,N_3949);
xnor U4081 (N_4081,N_3967,N_3875);
nand U4082 (N_4082,N_3943,N_3972);
nor U4083 (N_4083,N_3988,N_3996);
xor U4084 (N_4084,N_3990,N_3903);
nor U4085 (N_4085,N_3962,N_3942);
nand U4086 (N_4086,N_3925,N_3948);
and U4087 (N_4087,N_3960,N_3982);
or U4088 (N_4088,N_3895,N_3879);
nand U4089 (N_4089,N_3980,N_3882);
nor U4090 (N_4090,N_3981,N_3954);
xor U4091 (N_4091,N_3956,N_3920);
nand U4092 (N_4092,N_3963,N_3929);
nand U4093 (N_4093,N_3993,N_3980);
nand U4094 (N_4094,N_3991,N_3890);
or U4095 (N_4095,N_3931,N_3910);
nand U4096 (N_4096,N_3909,N_3895);
and U4097 (N_4097,N_3960,N_3992);
or U4098 (N_4098,N_3974,N_3933);
xnor U4099 (N_4099,N_3877,N_3898);
nand U4100 (N_4100,N_3920,N_3999);
and U4101 (N_4101,N_3963,N_3888);
and U4102 (N_4102,N_3900,N_3948);
nor U4103 (N_4103,N_3912,N_3990);
xor U4104 (N_4104,N_3902,N_3958);
nand U4105 (N_4105,N_3984,N_3883);
nand U4106 (N_4106,N_3902,N_3986);
and U4107 (N_4107,N_3970,N_3955);
xnor U4108 (N_4108,N_3969,N_3984);
nor U4109 (N_4109,N_3918,N_3972);
nand U4110 (N_4110,N_3981,N_3970);
and U4111 (N_4111,N_3927,N_3929);
nand U4112 (N_4112,N_3923,N_3959);
nor U4113 (N_4113,N_3977,N_3971);
and U4114 (N_4114,N_3935,N_3924);
nand U4115 (N_4115,N_3887,N_3930);
and U4116 (N_4116,N_3906,N_3889);
nor U4117 (N_4117,N_3909,N_3899);
nor U4118 (N_4118,N_3878,N_3975);
and U4119 (N_4119,N_3970,N_3977);
nand U4120 (N_4120,N_3897,N_3969);
nand U4121 (N_4121,N_3967,N_3953);
or U4122 (N_4122,N_3902,N_3953);
and U4123 (N_4123,N_3880,N_3939);
nand U4124 (N_4124,N_3877,N_3955);
xnor U4125 (N_4125,N_4010,N_4092);
nor U4126 (N_4126,N_4088,N_4098);
xor U4127 (N_4127,N_4095,N_4004);
or U4128 (N_4128,N_4100,N_4072);
xor U4129 (N_4129,N_4053,N_4007);
or U4130 (N_4130,N_4060,N_4073);
nand U4131 (N_4131,N_4101,N_4091);
and U4132 (N_4132,N_4102,N_4103);
nand U4133 (N_4133,N_4124,N_4051);
nor U4134 (N_4134,N_4119,N_4071);
xnor U4135 (N_4135,N_4015,N_4087);
nor U4136 (N_4136,N_4027,N_4121);
nor U4137 (N_4137,N_4057,N_4038);
xor U4138 (N_4138,N_4041,N_4052);
nor U4139 (N_4139,N_4114,N_4040);
nor U4140 (N_4140,N_4120,N_4043);
or U4141 (N_4141,N_4078,N_4031);
nor U4142 (N_4142,N_4065,N_4122);
or U4143 (N_4143,N_4042,N_4047);
nor U4144 (N_4144,N_4014,N_4003);
or U4145 (N_4145,N_4044,N_4104);
nor U4146 (N_4146,N_4034,N_4096);
nor U4147 (N_4147,N_4116,N_4012);
or U4148 (N_4148,N_4062,N_4097);
nor U4149 (N_4149,N_4018,N_4056);
nor U4150 (N_4150,N_4061,N_4077);
nand U4151 (N_4151,N_4090,N_4108);
nand U4152 (N_4152,N_4111,N_4033);
xnor U4153 (N_4153,N_4115,N_4106);
and U4154 (N_4154,N_4109,N_4029);
or U4155 (N_4155,N_4084,N_4016);
nor U4156 (N_4156,N_4023,N_4093);
xor U4157 (N_4157,N_4080,N_4009);
xor U4158 (N_4158,N_4107,N_4067);
and U4159 (N_4159,N_4076,N_4112);
or U4160 (N_4160,N_4039,N_4035);
xor U4161 (N_4161,N_4070,N_4030);
nor U4162 (N_4162,N_4110,N_4036);
nand U4163 (N_4163,N_4045,N_4066);
xor U4164 (N_4164,N_4081,N_4026);
nor U4165 (N_4165,N_4024,N_4019);
and U4166 (N_4166,N_4082,N_4058);
xnor U4167 (N_4167,N_4074,N_4001);
or U4168 (N_4168,N_4075,N_4068);
nor U4169 (N_4169,N_4055,N_4105);
or U4170 (N_4170,N_4021,N_4046);
xnor U4171 (N_4171,N_4083,N_4017);
nand U4172 (N_4172,N_4118,N_4123);
and U4173 (N_4173,N_4054,N_4049);
or U4174 (N_4174,N_4099,N_4085);
nand U4175 (N_4175,N_4000,N_4059);
nor U4176 (N_4176,N_4028,N_4020);
and U4177 (N_4177,N_4069,N_4005);
xnor U4178 (N_4178,N_4094,N_4013);
or U4179 (N_4179,N_4079,N_4011);
nor U4180 (N_4180,N_4002,N_4064);
nor U4181 (N_4181,N_4089,N_4086);
nand U4182 (N_4182,N_4032,N_4006);
xor U4183 (N_4183,N_4037,N_4048);
and U4184 (N_4184,N_4113,N_4050);
nand U4185 (N_4185,N_4063,N_4117);
nor U4186 (N_4186,N_4008,N_4022);
xnor U4187 (N_4187,N_4025,N_4048);
nand U4188 (N_4188,N_4088,N_4013);
or U4189 (N_4189,N_4070,N_4067);
or U4190 (N_4190,N_4030,N_4052);
xnor U4191 (N_4191,N_4087,N_4024);
nand U4192 (N_4192,N_4087,N_4004);
nor U4193 (N_4193,N_4101,N_4059);
nor U4194 (N_4194,N_4085,N_4101);
nand U4195 (N_4195,N_4083,N_4027);
or U4196 (N_4196,N_4002,N_4082);
nand U4197 (N_4197,N_4068,N_4101);
and U4198 (N_4198,N_4116,N_4071);
or U4199 (N_4199,N_4112,N_4093);
nand U4200 (N_4200,N_4068,N_4072);
xnor U4201 (N_4201,N_4076,N_4078);
xnor U4202 (N_4202,N_4091,N_4095);
or U4203 (N_4203,N_4085,N_4049);
nor U4204 (N_4204,N_4123,N_4090);
nand U4205 (N_4205,N_4005,N_4067);
nor U4206 (N_4206,N_4093,N_4044);
nor U4207 (N_4207,N_4106,N_4020);
xnor U4208 (N_4208,N_4039,N_4034);
and U4209 (N_4209,N_4009,N_4074);
nor U4210 (N_4210,N_4050,N_4002);
and U4211 (N_4211,N_4071,N_4094);
nand U4212 (N_4212,N_4064,N_4027);
nor U4213 (N_4213,N_4040,N_4009);
nor U4214 (N_4214,N_4042,N_4005);
nor U4215 (N_4215,N_4087,N_4014);
nor U4216 (N_4216,N_4007,N_4120);
or U4217 (N_4217,N_4031,N_4070);
or U4218 (N_4218,N_4089,N_4087);
or U4219 (N_4219,N_4060,N_4006);
xor U4220 (N_4220,N_4115,N_4042);
xor U4221 (N_4221,N_4108,N_4119);
nor U4222 (N_4222,N_4070,N_4064);
nand U4223 (N_4223,N_4069,N_4092);
nor U4224 (N_4224,N_4112,N_4113);
nand U4225 (N_4225,N_4098,N_4063);
xor U4226 (N_4226,N_4112,N_4052);
nand U4227 (N_4227,N_4124,N_4032);
and U4228 (N_4228,N_4054,N_4001);
nor U4229 (N_4229,N_4045,N_4102);
xor U4230 (N_4230,N_4121,N_4045);
xnor U4231 (N_4231,N_4058,N_4069);
xnor U4232 (N_4232,N_4063,N_4004);
and U4233 (N_4233,N_4050,N_4070);
and U4234 (N_4234,N_4115,N_4084);
nand U4235 (N_4235,N_4082,N_4039);
nor U4236 (N_4236,N_4040,N_4036);
xor U4237 (N_4237,N_4030,N_4076);
and U4238 (N_4238,N_4054,N_4042);
nor U4239 (N_4239,N_4033,N_4096);
nand U4240 (N_4240,N_4042,N_4068);
nand U4241 (N_4241,N_4122,N_4058);
nor U4242 (N_4242,N_4113,N_4099);
nand U4243 (N_4243,N_4100,N_4019);
and U4244 (N_4244,N_4031,N_4112);
nand U4245 (N_4245,N_4004,N_4082);
xor U4246 (N_4246,N_4043,N_4124);
nand U4247 (N_4247,N_4118,N_4032);
nor U4248 (N_4248,N_4011,N_4087);
nor U4249 (N_4249,N_4065,N_4097);
nor U4250 (N_4250,N_4127,N_4151);
nor U4251 (N_4251,N_4198,N_4210);
or U4252 (N_4252,N_4147,N_4191);
or U4253 (N_4253,N_4248,N_4194);
or U4254 (N_4254,N_4163,N_4234);
and U4255 (N_4255,N_4197,N_4239);
nand U4256 (N_4256,N_4170,N_4203);
nand U4257 (N_4257,N_4189,N_4192);
or U4258 (N_4258,N_4230,N_4220);
and U4259 (N_4259,N_4219,N_4196);
nor U4260 (N_4260,N_4174,N_4222);
xnor U4261 (N_4261,N_4214,N_4178);
and U4262 (N_4262,N_4140,N_4217);
nand U4263 (N_4263,N_4158,N_4168);
or U4264 (N_4264,N_4136,N_4139);
xnor U4265 (N_4265,N_4167,N_4185);
nor U4266 (N_4266,N_4190,N_4244);
xor U4267 (N_4267,N_4157,N_4205);
or U4268 (N_4268,N_4200,N_4213);
or U4269 (N_4269,N_4129,N_4146);
or U4270 (N_4270,N_4161,N_4240);
nand U4271 (N_4271,N_4224,N_4226);
xor U4272 (N_4272,N_4128,N_4164);
or U4273 (N_4273,N_4169,N_4188);
nand U4274 (N_4274,N_4154,N_4232);
nand U4275 (N_4275,N_4159,N_4166);
xor U4276 (N_4276,N_4207,N_4186);
and U4277 (N_4277,N_4182,N_4181);
nand U4278 (N_4278,N_4135,N_4176);
or U4279 (N_4279,N_4247,N_4177);
nor U4280 (N_4280,N_4237,N_4141);
and U4281 (N_4281,N_4249,N_4236);
nor U4282 (N_4282,N_4195,N_4148);
xnor U4283 (N_4283,N_4216,N_4223);
and U4284 (N_4284,N_4153,N_4221);
and U4285 (N_4285,N_4199,N_4215);
or U4286 (N_4286,N_4201,N_4227);
nand U4287 (N_4287,N_4245,N_4160);
or U4288 (N_4288,N_4211,N_4132);
xor U4289 (N_4289,N_4171,N_4145);
or U4290 (N_4290,N_4246,N_4202);
xnor U4291 (N_4291,N_4152,N_4130);
or U4292 (N_4292,N_4243,N_4233);
or U4293 (N_4293,N_4179,N_4150);
nor U4294 (N_4294,N_4125,N_4162);
xnor U4295 (N_4295,N_4143,N_4165);
nor U4296 (N_4296,N_4138,N_4206);
or U4297 (N_4297,N_4208,N_4144);
or U4298 (N_4298,N_4133,N_4242);
and U4299 (N_4299,N_4212,N_4155);
nand U4300 (N_4300,N_4156,N_4137);
and U4301 (N_4301,N_4225,N_4231);
and U4302 (N_4302,N_4149,N_4187);
nand U4303 (N_4303,N_4126,N_4193);
nor U4304 (N_4304,N_4209,N_4180);
nand U4305 (N_4305,N_4183,N_4218);
and U4306 (N_4306,N_4204,N_4238);
and U4307 (N_4307,N_4241,N_4235);
nand U4308 (N_4308,N_4131,N_4134);
nand U4309 (N_4309,N_4142,N_4172);
xor U4310 (N_4310,N_4175,N_4184);
nor U4311 (N_4311,N_4173,N_4229);
and U4312 (N_4312,N_4228,N_4197);
nor U4313 (N_4313,N_4235,N_4156);
xor U4314 (N_4314,N_4144,N_4211);
nand U4315 (N_4315,N_4181,N_4221);
nor U4316 (N_4316,N_4141,N_4162);
and U4317 (N_4317,N_4140,N_4202);
xnor U4318 (N_4318,N_4139,N_4239);
and U4319 (N_4319,N_4145,N_4189);
or U4320 (N_4320,N_4203,N_4162);
or U4321 (N_4321,N_4217,N_4137);
and U4322 (N_4322,N_4200,N_4196);
and U4323 (N_4323,N_4179,N_4137);
nand U4324 (N_4324,N_4126,N_4185);
nand U4325 (N_4325,N_4175,N_4192);
nand U4326 (N_4326,N_4243,N_4152);
nand U4327 (N_4327,N_4180,N_4146);
nor U4328 (N_4328,N_4158,N_4201);
nand U4329 (N_4329,N_4195,N_4159);
and U4330 (N_4330,N_4195,N_4202);
nand U4331 (N_4331,N_4219,N_4241);
and U4332 (N_4332,N_4176,N_4143);
nand U4333 (N_4333,N_4199,N_4126);
and U4334 (N_4334,N_4161,N_4236);
or U4335 (N_4335,N_4152,N_4128);
or U4336 (N_4336,N_4130,N_4202);
xor U4337 (N_4337,N_4240,N_4229);
or U4338 (N_4338,N_4191,N_4168);
nand U4339 (N_4339,N_4135,N_4194);
or U4340 (N_4340,N_4164,N_4238);
or U4341 (N_4341,N_4132,N_4213);
xor U4342 (N_4342,N_4234,N_4197);
and U4343 (N_4343,N_4166,N_4209);
and U4344 (N_4344,N_4150,N_4138);
or U4345 (N_4345,N_4243,N_4192);
or U4346 (N_4346,N_4131,N_4162);
nor U4347 (N_4347,N_4213,N_4224);
nor U4348 (N_4348,N_4138,N_4180);
xor U4349 (N_4349,N_4248,N_4190);
nor U4350 (N_4350,N_4166,N_4236);
and U4351 (N_4351,N_4172,N_4201);
and U4352 (N_4352,N_4142,N_4134);
xnor U4353 (N_4353,N_4205,N_4246);
nand U4354 (N_4354,N_4220,N_4181);
or U4355 (N_4355,N_4125,N_4210);
xnor U4356 (N_4356,N_4127,N_4198);
nor U4357 (N_4357,N_4248,N_4199);
nand U4358 (N_4358,N_4221,N_4128);
nand U4359 (N_4359,N_4235,N_4128);
and U4360 (N_4360,N_4183,N_4191);
nor U4361 (N_4361,N_4187,N_4131);
or U4362 (N_4362,N_4243,N_4197);
and U4363 (N_4363,N_4226,N_4132);
and U4364 (N_4364,N_4194,N_4131);
or U4365 (N_4365,N_4128,N_4157);
and U4366 (N_4366,N_4144,N_4178);
nor U4367 (N_4367,N_4226,N_4189);
xnor U4368 (N_4368,N_4170,N_4205);
nor U4369 (N_4369,N_4151,N_4219);
nand U4370 (N_4370,N_4154,N_4142);
nand U4371 (N_4371,N_4234,N_4204);
and U4372 (N_4372,N_4177,N_4221);
or U4373 (N_4373,N_4148,N_4155);
nor U4374 (N_4374,N_4185,N_4204);
nand U4375 (N_4375,N_4348,N_4305);
xor U4376 (N_4376,N_4337,N_4298);
or U4377 (N_4377,N_4331,N_4262);
nand U4378 (N_4378,N_4372,N_4273);
nand U4379 (N_4379,N_4304,N_4277);
xor U4380 (N_4380,N_4322,N_4309);
nand U4381 (N_4381,N_4314,N_4317);
and U4382 (N_4382,N_4318,N_4371);
nand U4383 (N_4383,N_4306,N_4342);
nand U4384 (N_4384,N_4257,N_4275);
nand U4385 (N_4385,N_4296,N_4367);
nor U4386 (N_4386,N_4343,N_4285);
nand U4387 (N_4387,N_4347,N_4313);
and U4388 (N_4388,N_4350,N_4357);
or U4389 (N_4389,N_4312,N_4287);
nor U4390 (N_4390,N_4272,N_4292);
and U4391 (N_4391,N_4319,N_4316);
and U4392 (N_4392,N_4352,N_4320);
nand U4393 (N_4393,N_4370,N_4301);
nor U4394 (N_4394,N_4368,N_4267);
nor U4395 (N_4395,N_4253,N_4291);
nor U4396 (N_4396,N_4325,N_4258);
nor U4397 (N_4397,N_4271,N_4324);
nor U4398 (N_4398,N_4289,N_4270);
and U4399 (N_4399,N_4361,N_4280);
nand U4400 (N_4400,N_4264,N_4293);
nor U4401 (N_4401,N_4336,N_4329);
nand U4402 (N_4402,N_4295,N_4355);
nand U4403 (N_4403,N_4268,N_4328);
or U4404 (N_4404,N_4340,N_4300);
nand U4405 (N_4405,N_4374,N_4286);
and U4406 (N_4406,N_4333,N_4351);
and U4407 (N_4407,N_4327,N_4330);
and U4408 (N_4408,N_4335,N_4321);
xnor U4409 (N_4409,N_4297,N_4358);
nor U4410 (N_4410,N_4284,N_4344);
xnor U4411 (N_4411,N_4283,N_4261);
or U4412 (N_4412,N_4334,N_4363);
nand U4413 (N_4413,N_4302,N_4288);
or U4414 (N_4414,N_4269,N_4323);
nor U4415 (N_4415,N_4260,N_4266);
nand U4416 (N_4416,N_4373,N_4326);
or U4417 (N_4417,N_4346,N_4278);
and U4418 (N_4418,N_4369,N_4365);
and U4419 (N_4419,N_4339,N_4256);
or U4420 (N_4420,N_4307,N_4282);
nand U4421 (N_4421,N_4364,N_4290);
and U4422 (N_4422,N_4341,N_4349);
and U4423 (N_4423,N_4332,N_4263);
nor U4424 (N_4424,N_4255,N_4303);
or U4425 (N_4425,N_4299,N_4308);
and U4426 (N_4426,N_4356,N_4315);
or U4427 (N_4427,N_4252,N_4366);
or U4428 (N_4428,N_4281,N_4354);
nor U4429 (N_4429,N_4254,N_4259);
nand U4430 (N_4430,N_4279,N_4265);
nor U4431 (N_4431,N_4310,N_4345);
xnor U4432 (N_4432,N_4360,N_4294);
xnor U4433 (N_4433,N_4353,N_4338);
nor U4434 (N_4434,N_4362,N_4251);
xnor U4435 (N_4435,N_4250,N_4311);
or U4436 (N_4436,N_4276,N_4359);
xnor U4437 (N_4437,N_4274,N_4266);
nor U4438 (N_4438,N_4366,N_4292);
and U4439 (N_4439,N_4325,N_4278);
nor U4440 (N_4440,N_4297,N_4271);
nand U4441 (N_4441,N_4301,N_4283);
nor U4442 (N_4442,N_4278,N_4370);
and U4443 (N_4443,N_4370,N_4355);
nand U4444 (N_4444,N_4336,N_4278);
nand U4445 (N_4445,N_4346,N_4260);
and U4446 (N_4446,N_4317,N_4345);
and U4447 (N_4447,N_4281,N_4322);
and U4448 (N_4448,N_4307,N_4301);
xnor U4449 (N_4449,N_4268,N_4261);
and U4450 (N_4450,N_4312,N_4267);
xor U4451 (N_4451,N_4253,N_4369);
xor U4452 (N_4452,N_4330,N_4263);
nor U4453 (N_4453,N_4254,N_4358);
nor U4454 (N_4454,N_4329,N_4260);
nand U4455 (N_4455,N_4327,N_4290);
and U4456 (N_4456,N_4368,N_4372);
nand U4457 (N_4457,N_4369,N_4297);
and U4458 (N_4458,N_4289,N_4367);
xor U4459 (N_4459,N_4335,N_4364);
nor U4460 (N_4460,N_4304,N_4342);
nand U4461 (N_4461,N_4287,N_4361);
xnor U4462 (N_4462,N_4296,N_4353);
nor U4463 (N_4463,N_4349,N_4291);
nand U4464 (N_4464,N_4259,N_4343);
nand U4465 (N_4465,N_4327,N_4283);
nand U4466 (N_4466,N_4281,N_4286);
or U4467 (N_4467,N_4300,N_4290);
or U4468 (N_4468,N_4279,N_4355);
nor U4469 (N_4469,N_4302,N_4362);
and U4470 (N_4470,N_4280,N_4333);
or U4471 (N_4471,N_4266,N_4323);
and U4472 (N_4472,N_4323,N_4251);
nor U4473 (N_4473,N_4320,N_4332);
or U4474 (N_4474,N_4371,N_4314);
xor U4475 (N_4475,N_4326,N_4313);
nor U4476 (N_4476,N_4359,N_4324);
or U4477 (N_4477,N_4346,N_4306);
xnor U4478 (N_4478,N_4309,N_4261);
nor U4479 (N_4479,N_4281,N_4252);
or U4480 (N_4480,N_4280,N_4332);
nand U4481 (N_4481,N_4270,N_4359);
xor U4482 (N_4482,N_4326,N_4293);
and U4483 (N_4483,N_4336,N_4322);
xor U4484 (N_4484,N_4291,N_4354);
xnor U4485 (N_4485,N_4312,N_4300);
nand U4486 (N_4486,N_4314,N_4286);
xor U4487 (N_4487,N_4293,N_4325);
or U4488 (N_4488,N_4286,N_4293);
or U4489 (N_4489,N_4351,N_4318);
xor U4490 (N_4490,N_4360,N_4367);
xor U4491 (N_4491,N_4370,N_4312);
nand U4492 (N_4492,N_4335,N_4268);
nor U4493 (N_4493,N_4286,N_4334);
and U4494 (N_4494,N_4312,N_4310);
nor U4495 (N_4495,N_4371,N_4271);
and U4496 (N_4496,N_4334,N_4279);
nor U4497 (N_4497,N_4312,N_4328);
and U4498 (N_4498,N_4314,N_4361);
and U4499 (N_4499,N_4284,N_4318);
xor U4500 (N_4500,N_4478,N_4488);
nand U4501 (N_4501,N_4456,N_4445);
xor U4502 (N_4502,N_4435,N_4383);
xor U4503 (N_4503,N_4446,N_4391);
or U4504 (N_4504,N_4401,N_4461);
and U4505 (N_4505,N_4480,N_4432);
nand U4506 (N_4506,N_4386,N_4388);
or U4507 (N_4507,N_4466,N_4420);
nand U4508 (N_4508,N_4424,N_4455);
and U4509 (N_4509,N_4414,N_4473);
nor U4510 (N_4510,N_4458,N_4495);
and U4511 (N_4511,N_4477,N_4411);
nand U4512 (N_4512,N_4498,N_4467);
xor U4513 (N_4513,N_4393,N_4474);
xor U4514 (N_4514,N_4481,N_4492);
nand U4515 (N_4515,N_4475,N_4460);
nand U4516 (N_4516,N_4412,N_4403);
nand U4517 (N_4517,N_4448,N_4482);
nand U4518 (N_4518,N_4470,N_4394);
and U4519 (N_4519,N_4471,N_4485);
xor U4520 (N_4520,N_4493,N_4389);
and U4521 (N_4521,N_4465,N_4483);
or U4522 (N_4522,N_4399,N_4453);
or U4523 (N_4523,N_4380,N_4397);
nor U4524 (N_4524,N_4447,N_4489);
or U4525 (N_4525,N_4428,N_4384);
xor U4526 (N_4526,N_4407,N_4497);
and U4527 (N_4527,N_4499,N_4426);
or U4528 (N_4528,N_4395,N_4416);
and U4529 (N_4529,N_4417,N_4377);
nor U4530 (N_4530,N_4494,N_4443);
nand U4531 (N_4531,N_4487,N_4433);
nor U4532 (N_4532,N_4437,N_4436);
and U4533 (N_4533,N_4496,N_4408);
xnor U4534 (N_4534,N_4449,N_4486);
nand U4535 (N_4535,N_4419,N_4379);
nand U4536 (N_4536,N_4462,N_4457);
nor U4537 (N_4537,N_4469,N_4400);
and U4538 (N_4538,N_4450,N_4429);
nand U4539 (N_4539,N_4454,N_4398);
and U4540 (N_4540,N_4378,N_4413);
or U4541 (N_4541,N_4409,N_4376);
nor U4542 (N_4542,N_4434,N_4440);
or U4543 (N_4543,N_4410,N_4451);
xor U4544 (N_4544,N_4387,N_4441);
nand U4545 (N_4545,N_4479,N_4476);
and U4546 (N_4546,N_4390,N_4392);
nor U4547 (N_4547,N_4490,N_4402);
and U4548 (N_4548,N_4415,N_4404);
nand U4549 (N_4549,N_4431,N_4472);
nor U4550 (N_4550,N_4396,N_4381);
and U4551 (N_4551,N_4452,N_4439);
nor U4552 (N_4552,N_4459,N_4438);
nor U4553 (N_4553,N_4464,N_4430);
nor U4554 (N_4554,N_4418,N_4468);
or U4555 (N_4555,N_4444,N_4484);
nor U4556 (N_4556,N_4425,N_4422);
nor U4557 (N_4557,N_4442,N_4405);
or U4558 (N_4558,N_4406,N_4385);
nor U4559 (N_4559,N_4491,N_4421);
nand U4560 (N_4560,N_4463,N_4427);
xor U4561 (N_4561,N_4382,N_4423);
or U4562 (N_4562,N_4375,N_4471);
nor U4563 (N_4563,N_4421,N_4499);
xor U4564 (N_4564,N_4441,N_4388);
nor U4565 (N_4565,N_4383,N_4494);
xor U4566 (N_4566,N_4463,N_4464);
xnor U4567 (N_4567,N_4421,N_4484);
or U4568 (N_4568,N_4379,N_4378);
and U4569 (N_4569,N_4396,N_4427);
nor U4570 (N_4570,N_4413,N_4447);
nand U4571 (N_4571,N_4454,N_4429);
nand U4572 (N_4572,N_4422,N_4462);
xor U4573 (N_4573,N_4396,N_4412);
nand U4574 (N_4574,N_4451,N_4439);
nor U4575 (N_4575,N_4492,N_4460);
nor U4576 (N_4576,N_4407,N_4434);
and U4577 (N_4577,N_4388,N_4391);
xnor U4578 (N_4578,N_4429,N_4471);
or U4579 (N_4579,N_4444,N_4386);
or U4580 (N_4580,N_4457,N_4440);
nand U4581 (N_4581,N_4435,N_4493);
nand U4582 (N_4582,N_4450,N_4376);
nand U4583 (N_4583,N_4496,N_4476);
nor U4584 (N_4584,N_4449,N_4448);
nor U4585 (N_4585,N_4389,N_4460);
or U4586 (N_4586,N_4423,N_4457);
nor U4587 (N_4587,N_4498,N_4407);
or U4588 (N_4588,N_4417,N_4420);
and U4589 (N_4589,N_4398,N_4487);
and U4590 (N_4590,N_4390,N_4494);
or U4591 (N_4591,N_4415,N_4483);
xor U4592 (N_4592,N_4476,N_4403);
and U4593 (N_4593,N_4443,N_4398);
nand U4594 (N_4594,N_4452,N_4498);
xor U4595 (N_4595,N_4401,N_4387);
xor U4596 (N_4596,N_4401,N_4460);
and U4597 (N_4597,N_4397,N_4426);
or U4598 (N_4598,N_4404,N_4480);
or U4599 (N_4599,N_4378,N_4457);
nand U4600 (N_4600,N_4427,N_4431);
and U4601 (N_4601,N_4419,N_4425);
nand U4602 (N_4602,N_4406,N_4426);
nand U4603 (N_4603,N_4458,N_4488);
nor U4604 (N_4604,N_4421,N_4409);
nor U4605 (N_4605,N_4390,N_4407);
and U4606 (N_4606,N_4436,N_4483);
nand U4607 (N_4607,N_4390,N_4383);
nand U4608 (N_4608,N_4439,N_4404);
or U4609 (N_4609,N_4456,N_4471);
nor U4610 (N_4610,N_4398,N_4423);
nor U4611 (N_4611,N_4484,N_4483);
nor U4612 (N_4612,N_4421,N_4482);
xor U4613 (N_4613,N_4391,N_4444);
xor U4614 (N_4614,N_4379,N_4387);
nor U4615 (N_4615,N_4452,N_4442);
and U4616 (N_4616,N_4487,N_4456);
or U4617 (N_4617,N_4457,N_4450);
or U4618 (N_4618,N_4383,N_4396);
and U4619 (N_4619,N_4494,N_4384);
xnor U4620 (N_4620,N_4392,N_4482);
xor U4621 (N_4621,N_4465,N_4490);
nand U4622 (N_4622,N_4423,N_4471);
xnor U4623 (N_4623,N_4419,N_4452);
nand U4624 (N_4624,N_4461,N_4470);
and U4625 (N_4625,N_4547,N_4597);
nand U4626 (N_4626,N_4611,N_4580);
or U4627 (N_4627,N_4621,N_4528);
and U4628 (N_4628,N_4582,N_4616);
or U4629 (N_4629,N_4555,N_4619);
nor U4630 (N_4630,N_4512,N_4588);
or U4631 (N_4631,N_4561,N_4553);
or U4632 (N_4632,N_4583,N_4593);
nand U4633 (N_4633,N_4504,N_4569);
nand U4634 (N_4634,N_4530,N_4554);
nor U4635 (N_4635,N_4581,N_4538);
or U4636 (N_4636,N_4562,N_4510);
and U4637 (N_4637,N_4518,N_4624);
and U4638 (N_4638,N_4603,N_4513);
and U4639 (N_4639,N_4590,N_4594);
and U4640 (N_4640,N_4577,N_4601);
or U4641 (N_4641,N_4537,N_4516);
nand U4642 (N_4642,N_4568,N_4559);
and U4643 (N_4643,N_4578,N_4563);
nand U4644 (N_4644,N_4523,N_4526);
and U4645 (N_4645,N_4522,N_4543);
xor U4646 (N_4646,N_4505,N_4511);
nor U4647 (N_4647,N_4546,N_4531);
and U4648 (N_4648,N_4606,N_4520);
and U4649 (N_4649,N_4598,N_4571);
nor U4650 (N_4650,N_4587,N_4622);
or U4651 (N_4651,N_4532,N_4574);
xor U4652 (N_4652,N_4556,N_4623);
nand U4653 (N_4653,N_4552,N_4602);
or U4654 (N_4654,N_4525,N_4617);
xor U4655 (N_4655,N_4509,N_4605);
xnor U4656 (N_4656,N_4565,N_4506);
xor U4657 (N_4657,N_4533,N_4515);
xnor U4658 (N_4658,N_4540,N_4502);
or U4659 (N_4659,N_4592,N_4534);
or U4660 (N_4660,N_4508,N_4544);
and U4661 (N_4661,N_4613,N_4503);
nor U4662 (N_4662,N_4579,N_4591);
nand U4663 (N_4663,N_4567,N_4550);
nor U4664 (N_4664,N_4608,N_4557);
xnor U4665 (N_4665,N_4595,N_4558);
xor U4666 (N_4666,N_4620,N_4500);
nand U4667 (N_4667,N_4564,N_4519);
and U4668 (N_4668,N_4576,N_4507);
xnor U4669 (N_4669,N_4570,N_4539);
xnor U4670 (N_4670,N_4549,N_4514);
nand U4671 (N_4671,N_4575,N_4535);
xnor U4672 (N_4672,N_4560,N_4524);
nand U4673 (N_4673,N_4548,N_4584);
nand U4674 (N_4674,N_4589,N_4536);
nand U4675 (N_4675,N_4607,N_4542);
and U4676 (N_4676,N_4604,N_4573);
xor U4677 (N_4677,N_4529,N_4599);
or U4678 (N_4678,N_4551,N_4521);
nand U4679 (N_4679,N_4618,N_4596);
and U4680 (N_4680,N_4572,N_4527);
or U4681 (N_4681,N_4585,N_4501);
nor U4682 (N_4682,N_4517,N_4600);
and U4683 (N_4683,N_4615,N_4545);
and U4684 (N_4684,N_4609,N_4541);
and U4685 (N_4685,N_4586,N_4566);
nand U4686 (N_4686,N_4612,N_4614);
nor U4687 (N_4687,N_4610,N_4536);
xnor U4688 (N_4688,N_4545,N_4584);
nand U4689 (N_4689,N_4577,N_4622);
xnor U4690 (N_4690,N_4575,N_4562);
and U4691 (N_4691,N_4507,N_4605);
xnor U4692 (N_4692,N_4556,N_4619);
nor U4693 (N_4693,N_4583,N_4562);
nor U4694 (N_4694,N_4624,N_4527);
xor U4695 (N_4695,N_4616,N_4605);
xor U4696 (N_4696,N_4506,N_4523);
nand U4697 (N_4697,N_4542,N_4541);
nand U4698 (N_4698,N_4584,N_4514);
nor U4699 (N_4699,N_4617,N_4539);
nand U4700 (N_4700,N_4504,N_4597);
nor U4701 (N_4701,N_4564,N_4527);
or U4702 (N_4702,N_4580,N_4614);
xnor U4703 (N_4703,N_4609,N_4595);
and U4704 (N_4704,N_4507,N_4590);
xnor U4705 (N_4705,N_4597,N_4550);
nor U4706 (N_4706,N_4518,N_4596);
xnor U4707 (N_4707,N_4623,N_4595);
nand U4708 (N_4708,N_4605,N_4598);
nor U4709 (N_4709,N_4551,N_4505);
and U4710 (N_4710,N_4550,N_4590);
xor U4711 (N_4711,N_4603,N_4615);
nor U4712 (N_4712,N_4535,N_4528);
and U4713 (N_4713,N_4524,N_4578);
xor U4714 (N_4714,N_4598,N_4514);
nand U4715 (N_4715,N_4548,N_4539);
nor U4716 (N_4716,N_4584,N_4566);
nand U4717 (N_4717,N_4578,N_4599);
xor U4718 (N_4718,N_4551,N_4579);
or U4719 (N_4719,N_4579,N_4518);
and U4720 (N_4720,N_4624,N_4544);
or U4721 (N_4721,N_4558,N_4598);
nand U4722 (N_4722,N_4583,N_4617);
and U4723 (N_4723,N_4502,N_4595);
xor U4724 (N_4724,N_4504,N_4540);
nand U4725 (N_4725,N_4516,N_4506);
and U4726 (N_4726,N_4621,N_4619);
and U4727 (N_4727,N_4531,N_4533);
nand U4728 (N_4728,N_4527,N_4576);
or U4729 (N_4729,N_4508,N_4530);
or U4730 (N_4730,N_4583,N_4589);
xor U4731 (N_4731,N_4527,N_4571);
xor U4732 (N_4732,N_4545,N_4522);
xor U4733 (N_4733,N_4567,N_4524);
and U4734 (N_4734,N_4612,N_4592);
and U4735 (N_4735,N_4535,N_4584);
nand U4736 (N_4736,N_4604,N_4589);
nor U4737 (N_4737,N_4595,N_4533);
and U4738 (N_4738,N_4616,N_4568);
nand U4739 (N_4739,N_4616,N_4571);
nor U4740 (N_4740,N_4623,N_4532);
xor U4741 (N_4741,N_4539,N_4568);
or U4742 (N_4742,N_4579,N_4578);
nand U4743 (N_4743,N_4624,N_4553);
nor U4744 (N_4744,N_4539,N_4622);
nor U4745 (N_4745,N_4525,N_4615);
xnor U4746 (N_4746,N_4601,N_4622);
nor U4747 (N_4747,N_4562,N_4585);
xnor U4748 (N_4748,N_4571,N_4573);
or U4749 (N_4749,N_4599,N_4514);
or U4750 (N_4750,N_4649,N_4641);
nor U4751 (N_4751,N_4652,N_4703);
nor U4752 (N_4752,N_4735,N_4664);
and U4753 (N_4753,N_4686,N_4748);
xnor U4754 (N_4754,N_4696,N_4678);
nand U4755 (N_4755,N_4683,N_4702);
xnor U4756 (N_4756,N_4625,N_4638);
or U4757 (N_4757,N_4632,N_4650);
and U4758 (N_4758,N_4689,N_4634);
nor U4759 (N_4759,N_4692,N_4710);
nor U4760 (N_4760,N_4673,N_4745);
or U4761 (N_4761,N_4674,N_4714);
or U4762 (N_4762,N_4639,N_4690);
nor U4763 (N_4763,N_4712,N_4655);
xnor U4764 (N_4764,N_4734,N_4656);
nand U4765 (N_4765,N_4693,N_4661);
xor U4766 (N_4766,N_4726,N_4732);
and U4767 (N_4767,N_4642,N_4709);
xor U4768 (N_4768,N_4717,N_4628);
nor U4769 (N_4769,N_4665,N_4731);
nand U4770 (N_4770,N_4657,N_4727);
nor U4771 (N_4771,N_4699,N_4704);
nand U4772 (N_4772,N_4749,N_4654);
nor U4773 (N_4773,N_4708,N_4721);
nor U4774 (N_4774,N_4715,N_4705);
xnor U4775 (N_4775,N_4697,N_4694);
xnor U4776 (N_4776,N_4635,N_4725);
xnor U4777 (N_4777,N_4744,N_4640);
or U4778 (N_4778,N_4740,N_4722);
xor U4779 (N_4779,N_4716,N_4739);
nand U4780 (N_4780,N_4651,N_4698);
nor U4781 (N_4781,N_4733,N_4643);
xor U4782 (N_4782,N_4660,N_4645);
xnor U4783 (N_4783,N_4687,N_4743);
nor U4784 (N_4784,N_4653,N_4663);
and U4785 (N_4785,N_4679,N_4711);
nor U4786 (N_4786,N_4724,N_4747);
or U4787 (N_4787,N_4662,N_4701);
nor U4788 (N_4788,N_4626,N_4670);
or U4789 (N_4789,N_4682,N_4636);
nand U4790 (N_4790,N_4666,N_4680);
xor U4791 (N_4791,N_4720,N_4647);
nand U4792 (N_4792,N_4713,N_4742);
xor U4793 (N_4793,N_4671,N_4695);
or U4794 (N_4794,N_4675,N_4659);
nor U4795 (N_4795,N_4719,N_4738);
xor U4796 (N_4796,N_4637,N_4658);
nand U4797 (N_4797,N_4700,N_4631);
nor U4798 (N_4798,N_4672,N_4718);
xor U4799 (N_4799,N_4677,N_4667);
nor U4800 (N_4800,N_4684,N_4736);
xnor U4801 (N_4801,N_4627,N_4630);
xnor U4802 (N_4802,N_4633,N_4648);
xnor U4803 (N_4803,N_4723,N_4646);
nor U4804 (N_4804,N_4685,N_4669);
xor U4805 (N_4805,N_4681,N_4676);
xnor U4806 (N_4806,N_4741,N_4668);
nand U4807 (N_4807,N_4730,N_4737);
or U4808 (N_4808,N_4728,N_4729);
or U4809 (N_4809,N_4688,N_4706);
nand U4810 (N_4810,N_4707,N_4746);
xnor U4811 (N_4811,N_4644,N_4629);
or U4812 (N_4812,N_4691,N_4699);
or U4813 (N_4813,N_4626,N_4681);
nand U4814 (N_4814,N_4733,N_4705);
nor U4815 (N_4815,N_4732,N_4716);
nand U4816 (N_4816,N_4739,N_4662);
or U4817 (N_4817,N_4670,N_4705);
nand U4818 (N_4818,N_4693,N_4726);
nand U4819 (N_4819,N_4673,N_4658);
nor U4820 (N_4820,N_4698,N_4704);
nand U4821 (N_4821,N_4660,N_4726);
and U4822 (N_4822,N_4746,N_4721);
xnor U4823 (N_4823,N_4676,N_4670);
xnor U4824 (N_4824,N_4718,N_4748);
xor U4825 (N_4825,N_4684,N_4715);
or U4826 (N_4826,N_4642,N_4641);
nor U4827 (N_4827,N_4693,N_4655);
xor U4828 (N_4828,N_4718,N_4631);
nand U4829 (N_4829,N_4686,N_4698);
and U4830 (N_4830,N_4748,N_4641);
xnor U4831 (N_4831,N_4693,N_4692);
nand U4832 (N_4832,N_4634,N_4660);
xor U4833 (N_4833,N_4659,N_4708);
xor U4834 (N_4834,N_4704,N_4625);
nor U4835 (N_4835,N_4695,N_4647);
nand U4836 (N_4836,N_4631,N_4703);
nand U4837 (N_4837,N_4697,N_4717);
or U4838 (N_4838,N_4680,N_4704);
nand U4839 (N_4839,N_4677,N_4707);
and U4840 (N_4840,N_4655,N_4696);
nor U4841 (N_4841,N_4714,N_4742);
or U4842 (N_4842,N_4739,N_4737);
and U4843 (N_4843,N_4685,N_4716);
xnor U4844 (N_4844,N_4638,N_4709);
or U4845 (N_4845,N_4705,N_4735);
nand U4846 (N_4846,N_4734,N_4667);
nand U4847 (N_4847,N_4675,N_4726);
xor U4848 (N_4848,N_4695,N_4688);
and U4849 (N_4849,N_4742,N_4708);
or U4850 (N_4850,N_4720,N_4698);
nor U4851 (N_4851,N_4731,N_4739);
xnor U4852 (N_4852,N_4734,N_4708);
nor U4853 (N_4853,N_4688,N_4661);
xor U4854 (N_4854,N_4640,N_4715);
xnor U4855 (N_4855,N_4650,N_4704);
and U4856 (N_4856,N_4717,N_4724);
xnor U4857 (N_4857,N_4695,N_4728);
and U4858 (N_4858,N_4736,N_4630);
nor U4859 (N_4859,N_4742,N_4644);
xor U4860 (N_4860,N_4668,N_4657);
or U4861 (N_4861,N_4671,N_4670);
nor U4862 (N_4862,N_4679,N_4645);
nand U4863 (N_4863,N_4695,N_4721);
and U4864 (N_4864,N_4728,N_4652);
nand U4865 (N_4865,N_4745,N_4688);
or U4866 (N_4866,N_4630,N_4744);
nand U4867 (N_4867,N_4727,N_4675);
nand U4868 (N_4868,N_4699,N_4659);
and U4869 (N_4869,N_4717,N_4734);
or U4870 (N_4870,N_4646,N_4685);
nand U4871 (N_4871,N_4661,N_4728);
and U4872 (N_4872,N_4630,N_4682);
nand U4873 (N_4873,N_4641,N_4738);
and U4874 (N_4874,N_4714,N_4660);
nor U4875 (N_4875,N_4814,N_4827);
and U4876 (N_4876,N_4866,N_4775);
nand U4877 (N_4877,N_4753,N_4795);
nand U4878 (N_4878,N_4856,N_4777);
xnor U4879 (N_4879,N_4750,N_4847);
nand U4880 (N_4880,N_4767,N_4789);
xnor U4881 (N_4881,N_4836,N_4872);
xor U4882 (N_4882,N_4807,N_4774);
nand U4883 (N_4883,N_4843,N_4863);
and U4884 (N_4884,N_4758,N_4834);
nor U4885 (N_4885,N_4813,N_4845);
nor U4886 (N_4886,N_4848,N_4865);
nand U4887 (N_4887,N_4841,N_4844);
or U4888 (N_4888,N_4800,N_4802);
and U4889 (N_4889,N_4805,N_4756);
nand U4890 (N_4890,N_4793,N_4772);
nand U4891 (N_4891,N_4781,N_4852);
xnor U4892 (N_4892,N_4798,N_4842);
xor U4893 (N_4893,N_4780,N_4816);
and U4894 (N_4894,N_4768,N_4787);
xor U4895 (N_4895,N_4846,N_4764);
xnor U4896 (N_4896,N_4837,N_4851);
and U4897 (N_4897,N_4854,N_4796);
or U4898 (N_4898,N_4839,N_4760);
nand U4899 (N_4899,N_4861,N_4871);
or U4900 (N_4900,N_4754,N_4850);
and U4901 (N_4901,N_4765,N_4779);
nor U4902 (N_4902,N_4838,N_4868);
xnor U4903 (N_4903,N_4820,N_4828);
nor U4904 (N_4904,N_4812,N_4818);
nor U4905 (N_4905,N_4792,N_4809);
or U4906 (N_4906,N_4849,N_4794);
or U4907 (N_4907,N_4869,N_4858);
xnor U4908 (N_4908,N_4840,N_4755);
or U4909 (N_4909,N_4752,N_4867);
nor U4910 (N_4910,N_4819,N_4782);
nor U4911 (N_4911,N_4829,N_4776);
nor U4912 (N_4912,N_4810,N_4825);
and U4913 (N_4913,N_4808,N_4857);
or U4914 (N_4914,N_4801,N_4803);
xor U4915 (N_4915,N_4786,N_4799);
nand U4916 (N_4916,N_4831,N_4788);
and U4917 (N_4917,N_4806,N_4762);
or U4918 (N_4918,N_4830,N_4759);
and U4919 (N_4919,N_4853,N_4862);
nor U4920 (N_4920,N_4860,N_4821);
xnor U4921 (N_4921,N_4804,N_4835);
xor U4922 (N_4922,N_4864,N_4783);
and U4923 (N_4923,N_4784,N_4766);
or U4924 (N_4924,N_4763,N_4833);
and U4925 (N_4925,N_4771,N_4822);
xor U4926 (N_4926,N_4811,N_4770);
and U4927 (N_4927,N_4778,N_4874);
or U4928 (N_4928,N_4791,N_4826);
or U4929 (N_4929,N_4859,N_4773);
nor U4930 (N_4930,N_4815,N_4817);
or U4931 (N_4931,N_4757,N_4790);
nor U4932 (N_4932,N_4751,N_4855);
and U4933 (N_4933,N_4873,N_4823);
or U4934 (N_4934,N_4785,N_4824);
or U4935 (N_4935,N_4870,N_4797);
and U4936 (N_4936,N_4832,N_4761);
xor U4937 (N_4937,N_4769,N_4783);
or U4938 (N_4938,N_4852,N_4857);
xnor U4939 (N_4939,N_4782,N_4774);
or U4940 (N_4940,N_4829,N_4775);
xnor U4941 (N_4941,N_4807,N_4868);
nor U4942 (N_4942,N_4874,N_4769);
or U4943 (N_4943,N_4766,N_4787);
nor U4944 (N_4944,N_4761,N_4764);
and U4945 (N_4945,N_4786,N_4874);
or U4946 (N_4946,N_4764,N_4763);
nor U4947 (N_4947,N_4818,N_4847);
nand U4948 (N_4948,N_4763,N_4800);
nand U4949 (N_4949,N_4823,N_4794);
xnor U4950 (N_4950,N_4793,N_4816);
or U4951 (N_4951,N_4868,N_4805);
nor U4952 (N_4952,N_4770,N_4768);
or U4953 (N_4953,N_4790,N_4811);
xnor U4954 (N_4954,N_4766,N_4826);
nor U4955 (N_4955,N_4752,N_4873);
nor U4956 (N_4956,N_4833,N_4809);
xor U4957 (N_4957,N_4837,N_4793);
nor U4958 (N_4958,N_4868,N_4852);
nor U4959 (N_4959,N_4834,N_4835);
and U4960 (N_4960,N_4770,N_4861);
nor U4961 (N_4961,N_4847,N_4758);
xnor U4962 (N_4962,N_4800,N_4795);
nand U4963 (N_4963,N_4774,N_4825);
nor U4964 (N_4964,N_4779,N_4867);
xnor U4965 (N_4965,N_4835,N_4845);
or U4966 (N_4966,N_4861,N_4802);
and U4967 (N_4967,N_4783,N_4860);
and U4968 (N_4968,N_4790,N_4785);
xnor U4969 (N_4969,N_4863,N_4783);
or U4970 (N_4970,N_4863,N_4769);
or U4971 (N_4971,N_4866,N_4754);
xnor U4972 (N_4972,N_4865,N_4871);
xnor U4973 (N_4973,N_4815,N_4787);
and U4974 (N_4974,N_4834,N_4786);
nor U4975 (N_4975,N_4820,N_4849);
nor U4976 (N_4976,N_4870,N_4836);
nor U4977 (N_4977,N_4851,N_4824);
and U4978 (N_4978,N_4791,N_4753);
or U4979 (N_4979,N_4838,N_4865);
nand U4980 (N_4980,N_4780,N_4870);
nand U4981 (N_4981,N_4820,N_4807);
nor U4982 (N_4982,N_4867,N_4842);
xnor U4983 (N_4983,N_4821,N_4874);
nor U4984 (N_4984,N_4823,N_4797);
nand U4985 (N_4985,N_4813,N_4837);
or U4986 (N_4986,N_4796,N_4788);
or U4987 (N_4987,N_4813,N_4784);
nor U4988 (N_4988,N_4818,N_4794);
xor U4989 (N_4989,N_4863,N_4818);
nand U4990 (N_4990,N_4815,N_4843);
nand U4991 (N_4991,N_4783,N_4839);
or U4992 (N_4992,N_4869,N_4868);
or U4993 (N_4993,N_4860,N_4869);
or U4994 (N_4994,N_4778,N_4820);
nor U4995 (N_4995,N_4854,N_4848);
xnor U4996 (N_4996,N_4750,N_4828);
or U4997 (N_4997,N_4795,N_4778);
nor U4998 (N_4998,N_4858,N_4755);
and U4999 (N_4999,N_4824,N_4826);
and U5000 (N_5000,N_4886,N_4895);
nand U5001 (N_5001,N_4938,N_4997);
or U5002 (N_5002,N_4946,N_4904);
xnor U5003 (N_5003,N_4956,N_4881);
xor U5004 (N_5004,N_4897,N_4977);
and U5005 (N_5005,N_4990,N_4888);
nor U5006 (N_5006,N_4932,N_4890);
xor U5007 (N_5007,N_4905,N_4983);
nand U5008 (N_5008,N_4915,N_4995);
xor U5009 (N_5009,N_4978,N_4884);
xnor U5010 (N_5010,N_4943,N_4939);
xor U5011 (N_5011,N_4941,N_4914);
or U5012 (N_5012,N_4988,N_4962);
nand U5013 (N_5013,N_4976,N_4889);
and U5014 (N_5014,N_4937,N_4957);
and U5015 (N_5015,N_4921,N_4934);
nor U5016 (N_5016,N_4913,N_4925);
nor U5017 (N_5017,N_4930,N_4971);
nor U5018 (N_5018,N_4991,N_4961);
xnor U5019 (N_5019,N_4998,N_4892);
or U5020 (N_5020,N_4955,N_4965);
xnor U5021 (N_5021,N_4903,N_4918);
nand U5022 (N_5022,N_4894,N_4876);
or U5023 (N_5023,N_4901,N_4926);
xnor U5024 (N_5024,N_4935,N_4981);
xnor U5025 (N_5025,N_4909,N_4974);
nor U5026 (N_5026,N_4947,N_4911);
nor U5027 (N_5027,N_4979,N_4879);
nor U5028 (N_5028,N_4951,N_4899);
nor U5029 (N_5029,N_4880,N_4970);
nand U5030 (N_5030,N_4960,N_4906);
and U5031 (N_5031,N_4945,N_4982);
or U5032 (N_5032,N_4927,N_4968);
xnor U5033 (N_5033,N_4907,N_4989);
or U5034 (N_5034,N_4922,N_4958);
or U5035 (N_5035,N_4972,N_4973);
nand U5036 (N_5036,N_4987,N_4980);
nand U5037 (N_5037,N_4993,N_4984);
and U5038 (N_5038,N_4994,N_4942);
nor U5039 (N_5039,N_4966,N_4923);
or U5040 (N_5040,N_4940,N_4992);
nor U5041 (N_5041,N_4898,N_4964);
and U5042 (N_5042,N_4944,N_4875);
nor U5043 (N_5043,N_4896,N_4891);
nand U5044 (N_5044,N_4999,N_4948);
xor U5045 (N_5045,N_4910,N_4916);
or U5046 (N_5046,N_4936,N_4985);
nor U5047 (N_5047,N_4924,N_4928);
nor U5048 (N_5048,N_4931,N_4887);
nor U5049 (N_5049,N_4953,N_4996);
nor U5050 (N_5050,N_4929,N_4919);
nand U5051 (N_5051,N_4952,N_4883);
nand U5052 (N_5052,N_4912,N_4969);
or U5053 (N_5053,N_4949,N_4900);
and U5054 (N_5054,N_4967,N_4954);
and U5055 (N_5055,N_4950,N_4893);
nand U5056 (N_5056,N_4920,N_4933);
nand U5057 (N_5057,N_4975,N_4963);
and U5058 (N_5058,N_4917,N_4986);
and U5059 (N_5059,N_4877,N_4959);
and U5060 (N_5060,N_4902,N_4878);
or U5061 (N_5061,N_4885,N_4908);
xor U5062 (N_5062,N_4882,N_4988);
nor U5063 (N_5063,N_4892,N_4958);
and U5064 (N_5064,N_4886,N_4968);
and U5065 (N_5065,N_4884,N_4992);
nand U5066 (N_5066,N_4943,N_4991);
nor U5067 (N_5067,N_4951,N_4876);
and U5068 (N_5068,N_4984,N_4960);
and U5069 (N_5069,N_4905,N_4911);
and U5070 (N_5070,N_4955,N_4891);
or U5071 (N_5071,N_4907,N_4969);
nand U5072 (N_5072,N_4900,N_4992);
nand U5073 (N_5073,N_4921,N_4954);
xor U5074 (N_5074,N_4920,N_4989);
xor U5075 (N_5075,N_4958,N_4896);
and U5076 (N_5076,N_4946,N_4900);
xnor U5077 (N_5077,N_4959,N_4882);
or U5078 (N_5078,N_4964,N_4934);
or U5079 (N_5079,N_4999,N_4942);
xor U5080 (N_5080,N_4960,N_4965);
or U5081 (N_5081,N_4906,N_4908);
or U5082 (N_5082,N_4889,N_4974);
xnor U5083 (N_5083,N_4916,N_4957);
nand U5084 (N_5084,N_4912,N_4963);
and U5085 (N_5085,N_4882,N_4903);
nand U5086 (N_5086,N_4941,N_4882);
nand U5087 (N_5087,N_4906,N_4951);
nor U5088 (N_5088,N_4993,N_4931);
xnor U5089 (N_5089,N_4987,N_4924);
nor U5090 (N_5090,N_4960,N_4944);
and U5091 (N_5091,N_4987,N_4906);
and U5092 (N_5092,N_4979,N_4932);
xnor U5093 (N_5093,N_4923,N_4940);
or U5094 (N_5094,N_4974,N_4916);
nor U5095 (N_5095,N_4953,N_4886);
xor U5096 (N_5096,N_4902,N_4876);
and U5097 (N_5097,N_4927,N_4993);
or U5098 (N_5098,N_4887,N_4967);
xnor U5099 (N_5099,N_4982,N_4959);
xnor U5100 (N_5100,N_4981,N_4967);
xnor U5101 (N_5101,N_4997,N_4913);
nor U5102 (N_5102,N_4917,N_4924);
nor U5103 (N_5103,N_4918,N_4900);
or U5104 (N_5104,N_4987,N_4930);
nor U5105 (N_5105,N_4959,N_4947);
and U5106 (N_5106,N_4984,N_4967);
xnor U5107 (N_5107,N_4939,N_4895);
and U5108 (N_5108,N_4902,N_4949);
or U5109 (N_5109,N_4934,N_4890);
or U5110 (N_5110,N_4968,N_4890);
nand U5111 (N_5111,N_4881,N_4960);
or U5112 (N_5112,N_4914,N_4912);
nor U5113 (N_5113,N_4975,N_4875);
nor U5114 (N_5114,N_4953,N_4948);
or U5115 (N_5115,N_4963,N_4889);
and U5116 (N_5116,N_4903,N_4907);
nor U5117 (N_5117,N_4952,N_4910);
and U5118 (N_5118,N_4879,N_4961);
and U5119 (N_5119,N_4994,N_4939);
and U5120 (N_5120,N_4921,N_4953);
xor U5121 (N_5121,N_4921,N_4875);
or U5122 (N_5122,N_4963,N_4926);
xor U5123 (N_5123,N_4908,N_4932);
nand U5124 (N_5124,N_4876,N_4988);
xnor U5125 (N_5125,N_5100,N_5097);
xor U5126 (N_5126,N_5039,N_5075);
and U5127 (N_5127,N_5056,N_5035);
or U5128 (N_5128,N_5036,N_5019);
and U5129 (N_5129,N_5045,N_5041);
or U5130 (N_5130,N_5070,N_5093);
xnor U5131 (N_5131,N_5079,N_5105);
nor U5132 (N_5132,N_5037,N_5029);
nand U5133 (N_5133,N_5124,N_5121);
or U5134 (N_5134,N_5018,N_5102);
xnor U5135 (N_5135,N_5091,N_5011);
xnor U5136 (N_5136,N_5103,N_5088);
or U5137 (N_5137,N_5076,N_5024);
xnor U5138 (N_5138,N_5114,N_5020);
xor U5139 (N_5139,N_5013,N_5021);
nand U5140 (N_5140,N_5066,N_5002);
nor U5141 (N_5141,N_5050,N_5099);
xor U5142 (N_5142,N_5083,N_5030);
nor U5143 (N_5143,N_5109,N_5080);
and U5144 (N_5144,N_5110,N_5058);
nand U5145 (N_5145,N_5086,N_5003);
nand U5146 (N_5146,N_5046,N_5059);
and U5147 (N_5147,N_5032,N_5123);
nand U5148 (N_5148,N_5022,N_5023);
nand U5149 (N_5149,N_5062,N_5073);
and U5150 (N_5150,N_5064,N_5108);
and U5151 (N_5151,N_5087,N_5025);
and U5152 (N_5152,N_5112,N_5054);
nor U5153 (N_5153,N_5051,N_5063);
nand U5154 (N_5154,N_5004,N_5120);
and U5155 (N_5155,N_5052,N_5016);
nand U5156 (N_5156,N_5057,N_5082);
xor U5157 (N_5157,N_5034,N_5033);
nand U5158 (N_5158,N_5111,N_5010);
and U5159 (N_5159,N_5068,N_5027);
and U5160 (N_5160,N_5017,N_5014);
nand U5161 (N_5161,N_5106,N_5067);
and U5162 (N_5162,N_5101,N_5031);
nand U5163 (N_5163,N_5077,N_5049);
and U5164 (N_5164,N_5084,N_5090);
and U5165 (N_5165,N_5053,N_5107);
nand U5166 (N_5166,N_5038,N_5005);
xnor U5167 (N_5167,N_5078,N_5094);
or U5168 (N_5168,N_5000,N_5085);
or U5169 (N_5169,N_5072,N_5012);
and U5170 (N_5170,N_5071,N_5117);
and U5171 (N_5171,N_5113,N_5007);
nor U5172 (N_5172,N_5044,N_5042);
nor U5173 (N_5173,N_5069,N_5040);
or U5174 (N_5174,N_5104,N_5006);
xnor U5175 (N_5175,N_5098,N_5060);
or U5176 (N_5176,N_5009,N_5096);
or U5177 (N_5177,N_5122,N_5074);
nand U5178 (N_5178,N_5001,N_5095);
and U5179 (N_5179,N_5115,N_5028);
xnor U5180 (N_5180,N_5116,N_5119);
xor U5181 (N_5181,N_5092,N_5055);
and U5182 (N_5182,N_5048,N_5118);
nor U5183 (N_5183,N_5008,N_5015);
and U5184 (N_5184,N_5089,N_5026);
or U5185 (N_5185,N_5081,N_5061);
xnor U5186 (N_5186,N_5047,N_5065);
nand U5187 (N_5187,N_5043,N_5102);
xnor U5188 (N_5188,N_5049,N_5099);
xnor U5189 (N_5189,N_5074,N_5067);
nor U5190 (N_5190,N_5113,N_5044);
xor U5191 (N_5191,N_5065,N_5102);
or U5192 (N_5192,N_5047,N_5083);
or U5193 (N_5193,N_5085,N_5069);
nor U5194 (N_5194,N_5115,N_5043);
xnor U5195 (N_5195,N_5005,N_5080);
xor U5196 (N_5196,N_5061,N_5027);
xor U5197 (N_5197,N_5086,N_5087);
nand U5198 (N_5198,N_5116,N_5008);
nor U5199 (N_5199,N_5011,N_5052);
nand U5200 (N_5200,N_5112,N_5048);
or U5201 (N_5201,N_5081,N_5002);
xnor U5202 (N_5202,N_5035,N_5070);
nand U5203 (N_5203,N_5118,N_5109);
or U5204 (N_5204,N_5110,N_5056);
nand U5205 (N_5205,N_5087,N_5110);
or U5206 (N_5206,N_5083,N_5022);
nand U5207 (N_5207,N_5027,N_5118);
nand U5208 (N_5208,N_5098,N_5068);
nor U5209 (N_5209,N_5031,N_5073);
or U5210 (N_5210,N_5035,N_5037);
and U5211 (N_5211,N_5105,N_5066);
nor U5212 (N_5212,N_5051,N_5106);
xnor U5213 (N_5213,N_5109,N_5106);
nor U5214 (N_5214,N_5088,N_5085);
nand U5215 (N_5215,N_5076,N_5084);
xnor U5216 (N_5216,N_5065,N_5072);
and U5217 (N_5217,N_5089,N_5118);
or U5218 (N_5218,N_5052,N_5021);
nor U5219 (N_5219,N_5074,N_5002);
or U5220 (N_5220,N_5099,N_5005);
and U5221 (N_5221,N_5019,N_5115);
nor U5222 (N_5222,N_5043,N_5083);
and U5223 (N_5223,N_5049,N_5020);
nand U5224 (N_5224,N_5107,N_5077);
xor U5225 (N_5225,N_5000,N_5113);
or U5226 (N_5226,N_5105,N_5013);
nor U5227 (N_5227,N_5082,N_5069);
nand U5228 (N_5228,N_5079,N_5054);
and U5229 (N_5229,N_5013,N_5050);
or U5230 (N_5230,N_5086,N_5024);
or U5231 (N_5231,N_5115,N_5031);
or U5232 (N_5232,N_5035,N_5027);
and U5233 (N_5233,N_5096,N_5050);
xnor U5234 (N_5234,N_5070,N_5032);
or U5235 (N_5235,N_5075,N_5124);
nand U5236 (N_5236,N_5008,N_5042);
nor U5237 (N_5237,N_5101,N_5109);
xnor U5238 (N_5238,N_5056,N_5038);
nor U5239 (N_5239,N_5057,N_5007);
xor U5240 (N_5240,N_5034,N_5064);
or U5241 (N_5241,N_5078,N_5004);
or U5242 (N_5242,N_5046,N_5079);
xnor U5243 (N_5243,N_5077,N_5098);
nor U5244 (N_5244,N_5070,N_5033);
xnor U5245 (N_5245,N_5029,N_5043);
nor U5246 (N_5246,N_5120,N_5106);
xnor U5247 (N_5247,N_5067,N_5036);
nand U5248 (N_5248,N_5006,N_5015);
xnor U5249 (N_5249,N_5088,N_5119);
or U5250 (N_5250,N_5191,N_5165);
and U5251 (N_5251,N_5158,N_5149);
nand U5252 (N_5252,N_5198,N_5210);
xnor U5253 (N_5253,N_5173,N_5201);
or U5254 (N_5254,N_5197,N_5161);
xnor U5255 (N_5255,N_5204,N_5243);
or U5256 (N_5256,N_5238,N_5141);
nand U5257 (N_5257,N_5151,N_5240);
and U5258 (N_5258,N_5167,N_5164);
and U5259 (N_5259,N_5152,N_5246);
xor U5260 (N_5260,N_5144,N_5231);
xnor U5261 (N_5261,N_5142,N_5241);
and U5262 (N_5262,N_5216,N_5181);
nor U5263 (N_5263,N_5206,N_5163);
xor U5264 (N_5264,N_5217,N_5195);
or U5265 (N_5265,N_5226,N_5236);
or U5266 (N_5266,N_5242,N_5215);
and U5267 (N_5267,N_5160,N_5220);
or U5268 (N_5268,N_5187,N_5162);
nand U5269 (N_5269,N_5202,N_5219);
nor U5270 (N_5270,N_5147,N_5182);
and U5271 (N_5271,N_5138,N_5239);
and U5272 (N_5272,N_5245,N_5221);
nor U5273 (N_5273,N_5143,N_5218);
nand U5274 (N_5274,N_5211,N_5235);
xnor U5275 (N_5275,N_5159,N_5135);
xnor U5276 (N_5276,N_5196,N_5248);
nand U5277 (N_5277,N_5224,N_5190);
nand U5278 (N_5278,N_5131,N_5193);
nand U5279 (N_5279,N_5247,N_5130);
xnor U5280 (N_5280,N_5134,N_5174);
xor U5281 (N_5281,N_5213,N_5223);
xor U5282 (N_5282,N_5230,N_5183);
nor U5283 (N_5283,N_5146,N_5125);
nand U5284 (N_5284,N_5148,N_5171);
or U5285 (N_5285,N_5145,N_5234);
xor U5286 (N_5286,N_5132,N_5208);
nor U5287 (N_5287,N_5233,N_5176);
xor U5288 (N_5288,N_5168,N_5178);
or U5289 (N_5289,N_5212,N_5157);
nor U5290 (N_5290,N_5169,N_5170);
or U5291 (N_5291,N_5155,N_5189);
nor U5292 (N_5292,N_5156,N_5136);
or U5293 (N_5293,N_5140,N_5225);
nor U5294 (N_5294,N_5200,N_5222);
and U5295 (N_5295,N_5194,N_5229);
nor U5296 (N_5296,N_5129,N_5227);
or U5297 (N_5297,N_5137,N_5249);
nor U5298 (N_5298,N_5184,N_5205);
xor U5299 (N_5299,N_5214,N_5180);
nor U5300 (N_5300,N_5166,N_5133);
and U5301 (N_5301,N_5154,N_5150);
or U5302 (N_5302,N_5203,N_5185);
nor U5303 (N_5303,N_5172,N_5153);
and U5304 (N_5304,N_5209,N_5175);
nand U5305 (N_5305,N_5232,N_5139);
and U5306 (N_5306,N_5192,N_5126);
nor U5307 (N_5307,N_5207,N_5127);
nand U5308 (N_5308,N_5179,N_5199);
or U5309 (N_5309,N_5244,N_5128);
and U5310 (N_5310,N_5237,N_5186);
and U5311 (N_5311,N_5188,N_5228);
or U5312 (N_5312,N_5177,N_5182);
nor U5313 (N_5313,N_5164,N_5242);
and U5314 (N_5314,N_5196,N_5180);
nor U5315 (N_5315,N_5175,N_5219);
nor U5316 (N_5316,N_5213,N_5239);
and U5317 (N_5317,N_5212,N_5187);
or U5318 (N_5318,N_5222,N_5226);
or U5319 (N_5319,N_5147,N_5211);
nor U5320 (N_5320,N_5246,N_5216);
nand U5321 (N_5321,N_5141,N_5145);
nor U5322 (N_5322,N_5227,N_5208);
and U5323 (N_5323,N_5218,N_5189);
xor U5324 (N_5324,N_5178,N_5223);
or U5325 (N_5325,N_5232,N_5218);
and U5326 (N_5326,N_5237,N_5144);
and U5327 (N_5327,N_5224,N_5139);
and U5328 (N_5328,N_5210,N_5125);
xor U5329 (N_5329,N_5135,N_5143);
xnor U5330 (N_5330,N_5152,N_5144);
and U5331 (N_5331,N_5207,N_5238);
or U5332 (N_5332,N_5148,N_5158);
nor U5333 (N_5333,N_5241,N_5154);
and U5334 (N_5334,N_5212,N_5182);
and U5335 (N_5335,N_5249,N_5223);
and U5336 (N_5336,N_5131,N_5200);
xnor U5337 (N_5337,N_5248,N_5126);
or U5338 (N_5338,N_5202,N_5221);
nor U5339 (N_5339,N_5185,N_5137);
and U5340 (N_5340,N_5158,N_5160);
nor U5341 (N_5341,N_5203,N_5215);
nand U5342 (N_5342,N_5183,N_5218);
and U5343 (N_5343,N_5209,N_5164);
nand U5344 (N_5344,N_5162,N_5182);
or U5345 (N_5345,N_5178,N_5234);
or U5346 (N_5346,N_5179,N_5249);
or U5347 (N_5347,N_5133,N_5240);
nor U5348 (N_5348,N_5211,N_5227);
nand U5349 (N_5349,N_5125,N_5237);
nor U5350 (N_5350,N_5161,N_5215);
nor U5351 (N_5351,N_5134,N_5187);
or U5352 (N_5352,N_5159,N_5223);
xnor U5353 (N_5353,N_5142,N_5126);
xor U5354 (N_5354,N_5200,N_5185);
or U5355 (N_5355,N_5139,N_5131);
xnor U5356 (N_5356,N_5207,N_5220);
xnor U5357 (N_5357,N_5241,N_5180);
or U5358 (N_5358,N_5242,N_5224);
xor U5359 (N_5359,N_5236,N_5138);
and U5360 (N_5360,N_5243,N_5249);
or U5361 (N_5361,N_5158,N_5199);
xnor U5362 (N_5362,N_5186,N_5239);
and U5363 (N_5363,N_5228,N_5242);
or U5364 (N_5364,N_5220,N_5139);
or U5365 (N_5365,N_5216,N_5158);
and U5366 (N_5366,N_5127,N_5198);
and U5367 (N_5367,N_5184,N_5238);
and U5368 (N_5368,N_5245,N_5156);
xnor U5369 (N_5369,N_5177,N_5160);
and U5370 (N_5370,N_5125,N_5246);
or U5371 (N_5371,N_5143,N_5129);
nor U5372 (N_5372,N_5148,N_5130);
nor U5373 (N_5373,N_5167,N_5179);
or U5374 (N_5374,N_5201,N_5209);
or U5375 (N_5375,N_5283,N_5261);
xnor U5376 (N_5376,N_5374,N_5264);
xor U5377 (N_5377,N_5277,N_5347);
and U5378 (N_5378,N_5343,N_5367);
or U5379 (N_5379,N_5252,N_5269);
xor U5380 (N_5380,N_5327,N_5274);
nand U5381 (N_5381,N_5295,N_5253);
nor U5382 (N_5382,N_5302,N_5286);
and U5383 (N_5383,N_5263,N_5348);
nor U5384 (N_5384,N_5258,N_5271);
xor U5385 (N_5385,N_5312,N_5298);
xor U5386 (N_5386,N_5346,N_5337);
and U5387 (N_5387,N_5352,N_5294);
nand U5388 (N_5388,N_5338,N_5311);
xor U5389 (N_5389,N_5319,N_5344);
xor U5390 (N_5390,N_5308,N_5333);
or U5391 (N_5391,N_5361,N_5362);
nor U5392 (N_5392,N_5321,N_5260);
nand U5393 (N_5393,N_5280,N_5287);
nor U5394 (N_5394,N_5349,N_5254);
xor U5395 (N_5395,N_5325,N_5345);
or U5396 (N_5396,N_5341,N_5335);
nand U5397 (N_5397,N_5273,N_5285);
and U5398 (N_5398,N_5329,N_5296);
nand U5399 (N_5399,N_5315,N_5342);
nand U5400 (N_5400,N_5250,N_5265);
nand U5401 (N_5401,N_5282,N_5279);
nand U5402 (N_5402,N_5365,N_5320);
or U5403 (N_5403,N_5359,N_5370);
xor U5404 (N_5404,N_5363,N_5284);
or U5405 (N_5405,N_5313,N_5371);
nand U5406 (N_5406,N_5256,N_5290);
nor U5407 (N_5407,N_5306,N_5305);
xor U5408 (N_5408,N_5368,N_5336);
xor U5409 (N_5409,N_5353,N_5339);
nor U5410 (N_5410,N_5289,N_5364);
xnor U5411 (N_5411,N_5369,N_5357);
nor U5412 (N_5412,N_5324,N_5291);
nor U5413 (N_5413,N_5310,N_5372);
nand U5414 (N_5414,N_5328,N_5334);
or U5415 (N_5415,N_5251,N_5304);
and U5416 (N_5416,N_5373,N_5257);
and U5417 (N_5417,N_5266,N_5318);
or U5418 (N_5418,N_5314,N_5356);
or U5419 (N_5419,N_5322,N_5350);
xnor U5420 (N_5420,N_5303,N_5332);
xor U5421 (N_5421,N_5278,N_5267);
nand U5422 (N_5422,N_5323,N_5275);
nor U5423 (N_5423,N_5281,N_5262);
nor U5424 (N_5424,N_5292,N_5366);
xor U5425 (N_5425,N_5288,N_5259);
xnor U5426 (N_5426,N_5354,N_5358);
or U5427 (N_5427,N_5360,N_5330);
or U5428 (N_5428,N_5351,N_5326);
and U5429 (N_5429,N_5299,N_5316);
nand U5430 (N_5430,N_5270,N_5301);
xor U5431 (N_5431,N_5297,N_5272);
nand U5432 (N_5432,N_5355,N_5317);
nand U5433 (N_5433,N_5309,N_5307);
and U5434 (N_5434,N_5340,N_5268);
nand U5435 (N_5435,N_5300,N_5293);
xnor U5436 (N_5436,N_5276,N_5255);
xor U5437 (N_5437,N_5331,N_5305);
nand U5438 (N_5438,N_5287,N_5344);
nand U5439 (N_5439,N_5253,N_5300);
or U5440 (N_5440,N_5349,N_5337);
nand U5441 (N_5441,N_5279,N_5338);
nand U5442 (N_5442,N_5331,N_5357);
nor U5443 (N_5443,N_5270,N_5348);
xor U5444 (N_5444,N_5269,N_5340);
xor U5445 (N_5445,N_5282,N_5290);
or U5446 (N_5446,N_5370,N_5366);
or U5447 (N_5447,N_5361,N_5347);
or U5448 (N_5448,N_5285,N_5316);
nand U5449 (N_5449,N_5278,N_5293);
nand U5450 (N_5450,N_5283,N_5301);
or U5451 (N_5451,N_5291,N_5338);
xor U5452 (N_5452,N_5365,N_5340);
or U5453 (N_5453,N_5298,N_5284);
nor U5454 (N_5454,N_5344,N_5299);
xor U5455 (N_5455,N_5256,N_5267);
xnor U5456 (N_5456,N_5358,N_5329);
or U5457 (N_5457,N_5323,N_5346);
and U5458 (N_5458,N_5304,N_5336);
or U5459 (N_5459,N_5313,N_5305);
nand U5460 (N_5460,N_5287,N_5274);
nor U5461 (N_5461,N_5323,N_5308);
nand U5462 (N_5462,N_5347,N_5278);
nor U5463 (N_5463,N_5263,N_5356);
or U5464 (N_5464,N_5372,N_5303);
nand U5465 (N_5465,N_5349,N_5281);
or U5466 (N_5466,N_5350,N_5282);
or U5467 (N_5467,N_5310,N_5361);
nand U5468 (N_5468,N_5307,N_5282);
nand U5469 (N_5469,N_5267,N_5350);
nor U5470 (N_5470,N_5373,N_5271);
nand U5471 (N_5471,N_5361,N_5259);
nor U5472 (N_5472,N_5374,N_5346);
nor U5473 (N_5473,N_5255,N_5284);
nand U5474 (N_5474,N_5342,N_5373);
and U5475 (N_5475,N_5319,N_5284);
xor U5476 (N_5476,N_5323,N_5289);
nor U5477 (N_5477,N_5292,N_5346);
nand U5478 (N_5478,N_5302,N_5321);
xor U5479 (N_5479,N_5276,N_5287);
nand U5480 (N_5480,N_5365,N_5304);
nor U5481 (N_5481,N_5259,N_5336);
nand U5482 (N_5482,N_5373,N_5264);
xor U5483 (N_5483,N_5347,N_5282);
and U5484 (N_5484,N_5310,N_5328);
nand U5485 (N_5485,N_5374,N_5320);
nor U5486 (N_5486,N_5336,N_5323);
and U5487 (N_5487,N_5282,N_5364);
or U5488 (N_5488,N_5358,N_5319);
nand U5489 (N_5489,N_5338,N_5261);
nand U5490 (N_5490,N_5340,N_5271);
xnor U5491 (N_5491,N_5266,N_5278);
and U5492 (N_5492,N_5344,N_5367);
xnor U5493 (N_5493,N_5291,N_5278);
and U5494 (N_5494,N_5320,N_5334);
nor U5495 (N_5495,N_5274,N_5296);
and U5496 (N_5496,N_5352,N_5251);
xnor U5497 (N_5497,N_5365,N_5306);
or U5498 (N_5498,N_5360,N_5312);
nor U5499 (N_5499,N_5336,N_5355);
nand U5500 (N_5500,N_5383,N_5486);
nor U5501 (N_5501,N_5379,N_5398);
nor U5502 (N_5502,N_5431,N_5498);
xor U5503 (N_5503,N_5405,N_5467);
and U5504 (N_5504,N_5477,N_5404);
and U5505 (N_5505,N_5393,N_5392);
and U5506 (N_5506,N_5489,N_5471);
or U5507 (N_5507,N_5422,N_5481);
nand U5508 (N_5508,N_5375,N_5466);
nand U5509 (N_5509,N_5412,N_5480);
nand U5510 (N_5510,N_5494,N_5426);
and U5511 (N_5511,N_5464,N_5487);
xnor U5512 (N_5512,N_5483,N_5418);
nand U5513 (N_5513,N_5470,N_5419);
nand U5514 (N_5514,N_5459,N_5457);
and U5515 (N_5515,N_5473,N_5413);
nand U5516 (N_5516,N_5411,N_5462);
and U5517 (N_5517,N_5475,N_5440);
or U5518 (N_5518,N_5446,N_5414);
and U5519 (N_5519,N_5388,N_5380);
nand U5520 (N_5520,N_5463,N_5427);
nand U5521 (N_5521,N_5390,N_5485);
nor U5522 (N_5522,N_5402,N_5484);
xnor U5523 (N_5523,N_5469,N_5410);
nand U5524 (N_5524,N_5493,N_5434);
nand U5525 (N_5525,N_5472,N_5421);
and U5526 (N_5526,N_5381,N_5387);
nor U5527 (N_5527,N_5396,N_5382);
or U5528 (N_5528,N_5435,N_5445);
and U5529 (N_5529,N_5460,N_5443);
and U5530 (N_5530,N_5458,N_5451);
nand U5531 (N_5531,N_5496,N_5436);
or U5532 (N_5532,N_5461,N_5386);
or U5533 (N_5533,N_5497,N_5406);
or U5534 (N_5534,N_5384,N_5429);
nand U5535 (N_5535,N_5377,N_5409);
nor U5536 (N_5536,N_5447,N_5416);
xor U5537 (N_5537,N_5448,N_5389);
nor U5538 (N_5538,N_5400,N_5401);
xor U5539 (N_5539,N_5491,N_5482);
and U5540 (N_5540,N_5476,N_5391);
or U5541 (N_5541,N_5465,N_5442);
nor U5542 (N_5542,N_5453,N_5479);
nor U5543 (N_5543,N_5407,N_5433);
or U5544 (N_5544,N_5474,N_5378);
or U5545 (N_5545,N_5450,N_5438);
or U5546 (N_5546,N_5441,N_5399);
or U5547 (N_5547,N_5417,N_5452);
nand U5548 (N_5548,N_5376,N_5456);
xnor U5549 (N_5549,N_5468,N_5385);
nand U5550 (N_5550,N_5488,N_5428);
and U5551 (N_5551,N_5403,N_5395);
and U5552 (N_5552,N_5424,N_5397);
and U5553 (N_5553,N_5408,N_5420);
or U5554 (N_5554,N_5454,N_5437);
xnor U5555 (N_5555,N_5455,N_5430);
nand U5556 (N_5556,N_5478,N_5432);
or U5557 (N_5557,N_5492,N_5425);
nand U5558 (N_5558,N_5449,N_5439);
or U5559 (N_5559,N_5444,N_5490);
xnor U5560 (N_5560,N_5394,N_5499);
or U5561 (N_5561,N_5423,N_5495);
nor U5562 (N_5562,N_5415,N_5485);
nand U5563 (N_5563,N_5405,N_5443);
nand U5564 (N_5564,N_5438,N_5463);
nand U5565 (N_5565,N_5485,N_5398);
xor U5566 (N_5566,N_5398,N_5388);
and U5567 (N_5567,N_5494,N_5470);
or U5568 (N_5568,N_5480,N_5437);
or U5569 (N_5569,N_5413,N_5409);
nor U5570 (N_5570,N_5393,N_5487);
nor U5571 (N_5571,N_5408,N_5498);
xnor U5572 (N_5572,N_5459,N_5403);
and U5573 (N_5573,N_5440,N_5450);
nor U5574 (N_5574,N_5480,N_5380);
and U5575 (N_5575,N_5440,N_5406);
and U5576 (N_5576,N_5429,N_5446);
nand U5577 (N_5577,N_5384,N_5443);
xor U5578 (N_5578,N_5383,N_5433);
or U5579 (N_5579,N_5440,N_5483);
nor U5580 (N_5580,N_5404,N_5495);
nand U5581 (N_5581,N_5416,N_5451);
nor U5582 (N_5582,N_5489,N_5388);
or U5583 (N_5583,N_5400,N_5441);
nand U5584 (N_5584,N_5451,N_5494);
nand U5585 (N_5585,N_5468,N_5390);
or U5586 (N_5586,N_5391,N_5480);
nor U5587 (N_5587,N_5480,N_5462);
and U5588 (N_5588,N_5481,N_5458);
xor U5589 (N_5589,N_5453,N_5456);
or U5590 (N_5590,N_5488,N_5410);
xnor U5591 (N_5591,N_5464,N_5378);
and U5592 (N_5592,N_5402,N_5460);
and U5593 (N_5593,N_5448,N_5461);
or U5594 (N_5594,N_5394,N_5490);
and U5595 (N_5595,N_5494,N_5408);
and U5596 (N_5596,N_5446,N_5464);
and U5597 (N_5597,N_5466,N_5410);
nor U5598 (N_5598,N_5379,N_5463);
or U5599 (N_5599,N_5444,N_5397);
and U5600 (N_5600,N_5464,N_5428);
xor U5601 (N_5601,N_5494,N_5430);
or U5602 (N_5602,N_5499,N_5428);
xor U5603 (N_5603,N_5412,N_5426);
or U5604 (N_5604,N_5412,N_5415);
xor U5605 (N_5605,N_5412,N_5493);
xor U5606 (N_5606,N_5399,N_5394);
and U5607 (N_5607,N_5403,N_5462);
xnor U5608 (N_5608,N_5457,N_5427);
and U5609 (N_5609,N_5481,N_5482);
xnor U5610 (N_5610,N_5438,N_5418);
and U5611 (N_5611,N_5491,N_5383);
nand U5612 (N_5612,N_5413,N_5390);
and U5613 (N_5613,N_5397,N_5428);
or U5614 (N_5614,N_5417,N_5447);
nor U5615 (N_5615,N_5438,N_5412);
xnor U5616 (N_5616,N_5419,N_5462);
and U5617 (N_5617,N_5482,N_5456);
and U5618 (N_5618,N_5450,N_5451);
nor U5619 (N_5619,N_5440,N_5494);
and U5620 (N_5620,N_5490,N_5472);
nor U5621 (N_5621,N_5439,N_5483);
xnor U5622 (N_5622,N_5437,N_5479);
and U5623 (N_5623,N_5495,N_5385);
or U5624 (N_5624,N_5382,N_5376);
xnor U5625 (N_5625,N_5590,N_5613);
and U5626 (N_5626,N_5585,N_5600);
nor U5627 (N_5627,N_5609,N_5539);
nor U5628 (N_5628,N_5505,N_5531);
xnor U5629 (N_5629,N_5608,N_5564);
and U5630 (N_5630,N_5507,N_5533);
and U5631 (N_5631,N_5521,N_5549);
and U5632 (N_5632,N_5583,N_5602);
or U5633 (N_5633,N_5528,N_5553);
nand U5634 (N_5634,N_5614,N_5591);
nand U5635 (N_5635,N_5538,N_5510);
nand U5636 (N_5636,N_5569,N_5548);
nor U5637 (N_5637,N_5502,N_5573);
or U5638 (N_5638,N_5586,N_5612);
or U5639 (N_5639,N_5529,N_5558);
xor U5640 (N_5640,N_5588,N_5621);
or U5641 (N_5641,N_5576,N_5527);
xor U5642 (N_5642,N_5500,N_5554);
nand U5643 (N_5643,N_5530,N_5551);
or U5644 (N_5644,N_5525,N_5501);
xor U5645 (N_5645,N_5589,N_5598);
or U5646 (N_5646,N_5567,N_5603);
and U5647 (N_5647,N_5547,N_5575);
nor U5648 (N_5648,N_5556,N_5522);
nand U5649 (N_5649,N_5503,N_5519);
nand U5650 (N_5650,N_5592,N_5624);
xor U5651 (N_5651,N_5623,N_5601);
xor U5652 (N_5652,N_5618,N_5517);
and U5653 (N_5653,N_5559,N_5580);
or U5654 (N_5654,N_5615,N_5550);
nand U5655 (N_5655,N_5584,N_5563);
and U5656 (N_5656,N_5611,N_5574);
nand U5657 (N_5657,N_5596,N_5557);
nand U5658 (N_5658,N_5536,N_5523);
nor U5659 (N_5659,N_5509,N_5532);
nand U5660 (N_5660,N_5605,N_5599);
xor U5661 (N_5661,N_5593,N_5607);
xnor U5662 (N_5662,N_5565,N_5520);
nor U5663 (N_5663,N_5597,N_5508);
nand U5664 (N_5664,N_5577,N_5512);
nand U5665 (N_5665,N_5545,N_5604);
nor U5666 (N_5666,N_5537,N_5568);
nor U5667 (N_5667,N_5542,N_5540);
or U5668 (N_5668,N_5524,N_5606);
nor U5669 (N_5669,N_5587,N_5578);
and U5670 (N_5670,N_5513,N_5566);
xor U5671 (N_5671,N_5552,N_5582);
and U5672 (N_5672,N_5535,N_5534);
nor U5673 (N_5673,N_5516,N_5560);
nor U5674 (N_5674,N_5515,N_5572);
xor U5675 (N_5675,N_5595,N_5555);
or U5676 (N_5676,N_5581,N_5570);
and U5677 (N_5677,N_5546,N_5514);
and U5678 (N_5678,N_5504,N_5579);
and U5679 (N_5679,N_5619,N_5506);
xor U5680 (N_5680,N_5620,N_5541);
or U5681 (N_5681,N_5571,N_5616);
xor U5682 (N_5682,N_5511,N_5561);
and U5683 (N_5683,N_5594,N_5526);
nand U5684 (N_5684,N_5617,N_5518);
and U5685 (N_5685,N_5543,N_5562);
nand U5686 (N_5686,N_5622,N_5544);
and U5687 (N_5687,N_5610,N_5526);
xnor U5688 (N_5688,N_5541,N_5503);
nand U5689 (N_5689,N_5585,N_5546);
nand U5690 (N_5690,N_5546,N_5501);
or U5691 (N_5691,N_5505,N_5587);
or U5692 (N_5692,N_5523,N_5624);
nor U5693 (N_5693,N_5623,N_5556);
and U5694 (N_5694,N_5554,N_5589);
nor U5695 (N_5695,N_5583,N_5505);
or U5696 (N_5696,N_5574,N_5570);
nand U5697 (N_5697,N_5504,N_5611);
nor U5698 (N_5698,N_5579,N_5596);
or U5699 (N_5699,N_5536,N_5603);
or U5700 (N_5700,N_5582,N_5576);
nand U5701 (N_5701,N_5568,N_5517);
and U5702 (N_5702,N_5601,N_5562);
or U5703 (N_5703,N_5503,N_5608);
xnor U5704 (N_5704,N_5570,N_5598);
xnor U5705 (N_5705,N_5541,N_5527);
and U5706 (N_5706,N_5592,N_5564);
nor U5707 (N_5707,N_5600,N_5595);
xnor U5708 (N_5708,N_5595,N_5544);
or U5709 (N_5709,N_5566,N_5569);
or U5710 (N_5710,N_5617,N_5512);
nand U5711 (N_5711,N_5573,N_5558);
xor U5712 (N_5712,N_5577,N_5609);
and U5713 (N_5713,N_5552,N_5622);
and U5714 (N_5714,N_5577,N_5545);
or U5715 (N_5715,N_5558,N_5550);
nor U5716 (N_5716,N_5613,N_5597);
nand U5717 (N_5717,N_5621,N_5526);
and U5718 (N_5718,N_5607,N_5515);
nor U5719 (N_5719,N_5577,N_5546);
or U5720 (N_5720,N_5513,N_5572);
and U5721 (N_5721,N_5596,N_5504);
and U5722 (N_5722,N_5532,N_5537);
and U5723 (N_5723,N_5572,N_5583);
and U5724 (N_5724,N_5538,N_5617);
nor U5725 (N_5725,N_5545,N_5527);
xnor U5726 (N_5726,N_5587,N_5523);
and U5727 (N_5727,N_5560,N_5570);
and U5728 (N_5728,N_5555,N_5535);
or U5729 (N_5729,N_5540,N_5507);
or U5730 (N_5730,N_5584,N_5535);
xor U5731 (N_5731,N_5562,N_5610);
nor U5732 (N_5732,N_5579,N_5552);
nor U5733 (N_5733,N_5577,N_5602);
nor U5734 (N_5734,N_5529,N_5593);
and U5735 (N_5735,N_5575,N_5592);
nand U5736 (N_5736,N_5527,N_5535);
nand U5737 (N_5737,N_5525,N_5521);
or U5738 (N_5738,N_5548,N_5523);
xor U5739 (N_5739,N_5593,N_5509);
and U5740 (N_5740,N_5612,N_5509);
or U5741 (N_5741,N_5617,N_5587);
nand U5742 (N_5742,N_5526,N_5598);
nor U5743 (N_5743,N_5574,N_5610);
and U5744 (N_5744,N_5554,N_5542);
xor U5745 (N_5745,N_5507,N_5501);
or U5746 (N_5746,N_5563,N_5582);
or U5747 (N_5747,N_5556,N_5503);
and U5748 (N_5748,N_5505,N_5622);
nor U5749 (N_5749,N_5532,N_5559);
or U5750 (N_5750,N_5690,N_5696);
and U5751 (N_5751,N_5657,N_5705);
or U5752 (N_5752,N_5702,N_5729);
xor U5753 (N_5753,N_5714,N_5648);
nor U5754 (N_5754,N_5659,N_5736);
xnor U5755 (N_5755,N_5694,N_5720);
or U5756 (N_5756,N_5656,N_5725);
or U5757 (N_5757,N_5687,N_5661);
xor U5758 (N_5758,N_5654,N_5651);
xor U5759 (N_5759,N_5731,N_5633);
xnor U5760 (N_5760,N_5748,N_5710);
nand U5761 (N_5761,N_5677,N_5701);
xor U5762 (N_5762,N_5652,N_5745);
or U5763 (N_5763,N_5746,N_5674);
or U5764 (N_5764,N_5732,N_5653);
xor U5765 (N_5765,N_5704,N_5644);
nor U5766 (N_5766,N_5669,N_5639);
nand U5767 (N_5767,N_5715,N_5628);
and U5768 (N_5768,N_5672,N_5744);
or U5769 (N_5769,N_5703,N_5670);
xnor U5770 (N_5770,N_5636,N_5747);
and U5771 (N_5771,N_5655,N_5643);
xnor U5772 (N_5772,N_5634,N_5662);
xnor U5773 (N_5773,N_5660,N_5695);
or U5774 (N_5774,N_5666,N_5711);
nor U5775 (N_5775,N_5721,N_5685);
and U5776 (N_5776,N_5719,N_5734);
or U5777 (N_5777,N_5709,N_5650);
nor U5778 (N_5778,N_5675,N_5722);
nor U5779 (N_5779,N_5638,N_5649);
xor U5780 (N_5780,N_5686,N_5699);
nand U5781 (N_5781,N_5627,N_5642);
or U5782 (N_5782,N_5632,N_5724);
nand U5783 (N_5783,N_5716,N_5741);
or U5784 (N_5784,N_5663,N_5684);
or U5785 (N_5785,N_5645,N_5629);
xor U5786 (N_5786,N_5712,N_5692);
or U5787 (N_5787,N_5631,N_5665);
xnor U5788 (N_5788,N_5658,N_5738);
or U5789 (N_5789,N_5679,N_5689);
xor U5790 (N_5790,N_5707,N_5700);
nor U5791 (N_5791,N_5678,N_5733);
nor U5792 (N_5792,N_5718,N_5691);
or U5793 (N_5793,N_5676,N_5680);
nor U5794 (N_5794,N_5726,N_5646);
or U5795 (N_5795,N_5637,N_5693);
nor U5796 (N_5796,N_5697,N_5706);
xnor U5797 (N_5797,N_5739,N_5673);
or U5798 (N_5798,N_5742,N_5681);
and U5799 (N_5799,N_5708,N_5737);
nand U5800 (N_5800,N_5668,N_5682);
nand U5801 (N_5801,N_5626,N_5698);
nand U5802 (N_5802,N_5641,N_5730);
nor U5803 (N_5803,N_5723,N_5688);
xor U5804 (N_5804,N_5727,N_5717);
xor U5805 (N_5805,N_5667,N_5735);
xor U5806 (N_5806,N_5743,N_5640);
nor U5807 (N_5807,N_5683,N_5664);
xnor U5808 (N_5808,N_5625,N_5630);
nor U5809 (N_5809,N_5728,N_5749);
xor U5810 (N_5810,N_5713,N_5740);
nor U5811 (N_5811,N_5647,N_5671);
xor U5812 (N_5812,N_5635,N_5658);
or U5813 (N_5813,N_5661,N_5671);
or U5814 (N_5814,N_5669,N_5677);
xor U5815 (N_5815,N_5749,N_5640);
nand U5816 (N_5816,N_5745,N_5706);
xor U5817 (N_5817,N_5636,N_5625);
and U5818 (N_5818,N_5657,N_5707);
and U5819 (N_5819,N_5711,N_5649);
nand U5820 (N_5820,N_5658,N_5725);
or U5821 (N_5821,N_5693,N_5746);
or U5822 (N_5822,N_5654,N_5722);
nand U5823 (N_5823,N_5672,N_5649);
nor U5824 (N_5824,N_5729,N_5649);
or U5825 (N_5825,N_5628,N_5662);
xnor U5826 (N_5826,N_5707,N_5642);
nand U5827 (N_5827,N_5645,N_5746);
and U5828 (N_5828,N_5648,N_5627);
and U5829 (N_5829,N_5708,N_5669);
or U5830 (N_5830,N_5738,N_5718);
xor U5831 (N_5831,N_5636,N_5674);
or U5832 (N_5832,N_5661,N_5704);
or U5833 (N_5833,N_5668,N_5730);
or U5834 (N_5834,N_5654,N_5666);
xor U5835 (N_5835,N_5726,N_5625);
or U5836 (N_5836,N_5643,N_5725);
nor U5837 (N_5837,N_5721,N_5730);
nand U5838 (N_5838,N_5710,N_5747);
nor U5839 (N_5839,N_5693,N_5699);
or U5840 (N_5840,N_5698,N_5673);
xor U5841 (N_5841,N_5731,N_5655);
nor U5842 (N_5842,N_5723,N_5745);
and U5843 (N_5843,N_5734,N_5656);
and U5844 (N_5844,N_5728,N_5628);
nor U5845 (N_5845,N_5715,N_5724);
nand U5846 (N_5846,N_5711,N_5646);
nor U5847 (N_5847,N_5630,N_5715);
xnor U5848 (N_5848,N_5663,N_5689);
and U5849 (N_5849,N_5642,N_5644);
nand U5850 (N_5850,N_5660,N_5637);
xor U5851 (N_5851,N_5738,N_5698);
or U5852 (N_5852,N_5652,N_5747);
or U5853 (N_5853,N_5639,N_5733);
nand U5854 (N_5854,N_5711,N_5627);
nor U5855 (N_5855,N_5686,N_5740);
nand U5856 (N_5856,N_5691,N_5740);
nor U5857 (N_5857,N_5671,N_5640);
and U5858 (N_5858,N_5712,N_5631);
nor U5859 (N_5859,N_5647,N_5643);
nand U5860 (N_5860,N_5718,N_5736);
nor U5861 (N_5861,N_5664,N_5702);
xor U5862 (N_5862,N_5726,N_5660);
and U5863 (N_5863,N_5678,N_5692);
nor U5864 (N_5864,N_5630,N_5734);
and U5865 (N_5865,N_5694,N_5728);
and U5866 (N_5866,N_5650,N_5648);
nand U5867 (N_5867,N_5642,N_5652);
xor U5868 (N_5868,N_5659,N_5682);
or U5869 (N_5869,N_5679,N_5713);
nand U5870 (N_5870,N_5696,N_5670);
or U5871 (N_5871,N_5691,N_5699);
or U5872 (N_5872,N_5717,N_5714);
nor U5873 (N_5873,N_5718,N_5663);
nand U5874 (N_5874,N_5683,N_5740);
nand U5875 (N_5875,N_5780,N_5805);
xnor U5876 (N_5876,N_5856,N_5867);
nor U5877 (N_5877,N_5830,N_5802);
or U5878 (N_5878,N_5759,N_5874);
xor U5879 (N_5879,N_5848,N_5835);
and U5880 (N_5880,N_5871,N_5785);
nand U5881 (N_5881,N_5775,N_5790);
xor U5882 (N_5882,N_5819,N_5750);
or U5883 (N_5883,N_5752,N_5769);
xor U5884 (N_5884,N_5812,N_5852);
or U5885 (N_5885,N_5832,N_5807);
nor U5886 (N_5886,N_5806,N_5811);
or U5887 (N_5887,N_5808,N_5860);
nand U5888 (N_5888,N_5854,N_5777);
and U5889 (N_5889,N_5788,N_5774);
xnor U5890 (N_5890,N_5793,N_5839);
and U5891 (N_5891,N_5799,N_5761);
xor U5892 (N_5892,N_5797,N_5763);
nor U5893 (N_5893,N_5798,N_5764);
or U5894 (N_5894,N_5866,N_5762);
xnor U5895 (N_5895,N_5829,N_5840);
xor U5896 (N_5896,N_5861,N_5827);
xnor U5897 (N_5897,N_5841,N_5846);
nand U5898 (N_5898,N_5803,N_5809);
and U5899 (N_5899,N_5864,N_5784);
or U5900 (N_5900,N_5837,N_5767);
or U5901 (N_5901,N_5870,N_5825);
xor U5902 (N_5902,N_5789,N_5817);
nand U5903 (N_5903,N_5814,N_5843);
nor U5904 (N_5904,N_5765,N_5801);
nor U5905 (N_5905,N_5783,N_5773);
nand U5906 (N_5906,N_5804,N_5757);
and U5907 (N_5907,N_5868,N_5850);
or U5908 (N_5908,N_5824,N_5787);
nor U5909 (N_5909,N_5795,N_5820);
and U5910 (N_5910,N_5821,N_5778);
nand U5911 (N_5911,N_5863,N_5853);
nor U5912 (N_5912,N_5855,N_5770);
nand U5913 (N_5913,N_5776,N_5872);
nor U5914 (N_5914,N_5836,N_5838);
xnor U5915 (N_5915,N_5831,N_5849);
xor U5916 (N_5916,N_5766,N_5818);
and U5917 (N_5917,N_5858,N_5791);
nor U5918 (N_5918,N_5782,N_5873);
or U5919 (N_5919,N_5768,N_5815);
and U5920 (N_5920,N_5845,N_5834);
or U5921 (N_5921,N_5800,N_5859);
nor U5922 (N_5922,N_5862,N_5771);
nand U5923 (N_5923,N_5816,N_5779);
and U5924 (N_5924,N_5865,N_5826);
nand U5925 (N_5925,N_5781,N_5756);
or U5926 (N_5926,N_5842,N_5792);
xor U5927 (N_5927,N_5828,N_5794);
nor U5928 (N_5928,N_5755,N_5772);
and U5929 (N_5929,N_5751,N_5754);
xor U5930 (N_5930,N_5847,N_5869);
xnor U5931 (N_5931,N_5760,N_5822);
and U5932 (N_5932,N_5844,N_5753);
nand U5933 (N_5933,N_5796,N_5833);
or U5934 (N_5934,N_5813,N_5851);
nor U5935 (N_5935,N_5758,N_5786);
or U5936 (N_5936,N_5810,N_5857);
xnor U5937 (N_5937,N_5823,N_5821);
nand U5938 (N_5938,N_5782,N_5792);
or U5939 (N_5939,N_5785,N_5806);
or U5940 (N_5940,N_5772,N_5844);
nor U5941 (N_5941,N_5781,N_5851);
xor U5942 (N_5942,N_5824,N_5851);
nor U5943 (N_5943,N_5861,N_5817);
nand U5944 (N_5944,N_5855,N_5801);
xnor U5945 (N_5945,N_5859,N_5814);
nand U5946 (N_5946,N_5842,N_5840);
nor U5947 (N_5947,N_5848,N_5792);
or U5948 (N_5948,N_5780,N_5824);
or U5949 (N_5949,N_5770,N_5794);
nand U5950 (N_5950,N_5765,N_5854);
xor U5951 (N_5951,N_5789,N_5859);
nor U5952 (N_5952,N_5857,N_5779);
xor U5953 (N_5953,N_5759,N_5843);
nor U5954 (N_5954,N_5850,N_5793);
and U5955 (N_5955,N_5824,N_5806);
nor U5956 (N_5956,N_5837,N_5841);
and U5957 (N_5957,N_5764,N_5846);
nor U5958 (N_5958,N_5797,N_5771);
nand U5959 (N_5959,N_5752,N_5785);
nor U5960 (N_5960,N_5870,N_5817);
or U5961 (N_5961,N_5780,N_5870);
or U5962 (N_5962,N_5847,N_5765);
nand U5963 (N_5963,N_5816,N_5794);
or U5964 (N_5964,N_5755,N_5816);
nand U5965 (N_5965,N_5824,N_5841);
xor U5966 (N_5966,N_5831,N_5866);
or U5967 (N_5967,N_5861,N_5773);
and U5968 (N_5968,N_5771,N_5751);
and U5969 (N_5969,N_5804,N_5805);
nor U5970 (N_5970,N_5826,N_5810);
nand U5971 (N_5971,N_5807,N_5846);
and U5972 (N_5972,N_5765,N_5824);
nand U5973 (N_5973,N_5816,N_5808);
xor U5974 (N_5974,N_5758,N_5764);
and U5975 (N_5975,N_5777,N_5823);
or U5976 (N_5976,N_5857,N_5837);
or U5977 (N_5977,N_5868,N_5769);
nor U5978 (N_5978,N_5752,N_5767);
and U5979 (N_5979,N_5786,N_5834);
and U5980 (N_5980,N_5763,N_5835);
nand U5981 (N_5981,N_5801,N_5802);
nor U5982 (N_5982,N_5838,N_5841);
or U5983 (N_5983,N_5798,N_5783);
or U5984 (N_5984,N_5866,N_5796);
xnor U5985 (N_5985,N_5810,N_5759);
xnor U5986 (N_5986,N_5859,N_5824);
nor U5987 (N_5987,N_5855,N_5856);
nand U5988 (N_5988,N_5780,N_5871);
nor U5989 (N_5989,N_5817,N_5757);
xnor U5990 (N_5990,N_5786,N_5815);
xor U5991 (N_5991,N_5841,N_5794);
and U5992 (N_5992,N_5817,N_5845);
and U5993 (N_5993,N_5783,N_5753);
xor U5994 (N_5994,N_5867,N_5754);
xnor U5995 (N_5995,N_5854,N_5757);
or U5996 (N_5996,N_5811,N_5793);
nor U5997 (N_5997,N_5785,N_5775);
nand U5998 (N_5998,N_5838,N_5803);
nor U5999 (N_5999,N_5796,N_5804);
and U6000 (N_6000,N_5915,N_5985);
and U6001 (N_6001,N_5983,N_5893);
nor U6002 (N_6002,N_5965,N_5889);
or U6003 (N_6003,N_5999,N_5994);
nor U6004 (N_6004,N_5917,N_5878);
and U6005 (N_6005,N_5958,N_5953);
and U6006 (N_6006,N_5927,N_5892);
xor U6007 (N_6007,N_5976,N_5938);
nor U6008 (N_6008,N_5880,N_5903);
and U6009 (N_6009,N_5982,N_5951);
or U6010 (N_6010,N_5977,N_5905);
or U6011 (N_6011,N_5935,N_5993);
and U6012 (N_6012,N_5924,N_5901);
and U6013 (N_6013,N_5898,N_5995);
and U6014 (N_6014,N_5910,N_5939);
or U6015 (N_6015,N_5949,N_5975);
nand U6016 (N_6016,N_5877,N_5968);
and U6017 (N_6017,N_5998,N_5908);
and U6018 (N_6018,N_5967,N_5896);
nand U6019 (N_6019,N_5894,N_5974);
and U6020 (N_6020,N_5934,N_5990);
nor U6021 (N_6021,N_5984,N_5911);
nand U6022 (N_6022,N_5969,N_5971);
xnor U6023 (N_6023,N_5887,N_5921);
and U6024 (N_6024,N_5884,N_5972);
nor U6025 (N_6025,N_5897,N_5875);
or U6026 (N_6026,N_5970,N_5909);
nand U6027 (N_6027,N_5928,N_5964);
or U6028 (N_6028,N_5954,N_5918);
or U6029 (N_6029,N_5929,N_5950);
nor U6030 (N_6030,N_5992,N_5989);
or U6031 (N_6031,N_5952,N_5942);
nand U6032 (N_6032,N_5891,N_5900);
xor U6033 (N_6033,N_5945,N_5962);
and U6034 (N_6034,N_5933,N_5906);
or U6035 (N_6035,N_5926,N_5882);
nor U6036 (N_6036,N_5919,N_5980);
nand U6037 (N_6037,N_5943,N_5902);
nor U6038 (N_6038,N_5997,N_5899);
xor U6039 (N_6039,N_5883,N_5948);
or U6040 (N_6040,N_5940,N_5922);
nand U6041 (N_6041,N_5923,N_5876);
and U6042 (N_6042,N_5925,N_5946);
or U6043 (N_6043,N_5960,N_5895);
nor U6044 (N_6044,N_5955,N_5961);
nand U6045 (N_6045,N_5881,N_5904);
nor U6046 (N_6046,N_5963,N_5912);
nor U6047 (N_6047,N_5890,N_5941);
nor U6048 (N_6048,N_5956,N_5947);
nand U6049 (N_6049,N_5920,N_5936);
nor U6050 (N_6050,N_5885,N_5959);
and U6051 (N_6051,N_5957,N_5879);
xnor U6052 (N_6052,N_5930,N_5914);
or U6053 (N_6053,N_5973,N_5991);
xnor U6054 (N_6054,N_5981,N_5944);
nor U6055 (N_6055,N_5988,N_5986);
xnor U6056 (N_6056,N_5931,N_5978);
nand U6057 (N_6057,N_5937,N_5932);
nand U6058 (N_6058,N_5987,N_5966);
xor U6059 (N_6059,N_5979,N_5913);
xor U6060 (N_6060,N_5886,N_5888);
nor U6061 (N_6061,N_5907,N_5996);
nor U6062 (N_6062,N_5916,N_5938);
nand U6063 (N_6063,N_5890,N_5896);
xnor U6064 (N_6064,N_5911,N_5926);
or U6065 (N_6065,N_5916,N_5989);
xnor U6066 (N_6066,N_5962,N_5914);
and U6067 (N_6067,N_5964,N_5994);
xor U6068 (N_6068,N_5898,N_5899);
nand U6069 (N_6069,N_5965,N_5991);
nor U6070 (N_6070,N_5927,N_5942);
nor U6071 (N_6071,N_5913,N_5962);
and U6072 (N_6072,N_5889,N_5923);
nor U6073 (N_6073,N_5890,N_5882);
or U6074 (N_6074,N_5895,N_5963);
nor U6075 (N_6075,N_5943,N_5962);
or U6076 (N_6076,N_5988,N_5928);
nor U6077 (N_6077,N_5887,N_5939);
xor U6078 (N_6078,N_5997,N_5964);
nand U6079 (N_6079,N_5975,N_5925);
and U6080 (N_6080,N_5877,N_5878);
xor U6081 (N_6081,N_5900,N_5982);
xnor U6082 (N_6082,N_5909,N_5946);
and U6083 (N_6083,N_5925,N_5979);
nand U6084 (N_6084,N_5910,N_5938);
and U6085 (N_6085,N_5971,N_5953);
nand U6086 (N_6086,N_5966,N_5879);
nor U6087 (N_6087,N_5877,N_5937);
xnor U6088 (N_6088,N_5904,N_5977);
nand U6089 (N_6089,N_5893,N_5985);
xnor U6090 (N_6090,N_5987,N_5976);
nor U6091 (N_6091,N_5952,N_5997);
xor U6092 (N_6092,N_5912,N_5897);
nor U6093 (N_6093,N_5966,N_5899);
nor U6094 (N_6094,N_5882,N_5998);
nor U6095 (N_6095,N_5934,N_5883);
and U6096 (N_6096,N_5995,N_5895);
and U6097 (N_6097,N_5917,N_5906);
and U6098 (N_6098,N_5880,N_5972);
and U6099 (N_6099,N_5928,N_5906);
and U6100 (N_6100,N_5978,N_5981);
xnor U6101 (N_6101,N_5919,N_5987);
and U6102 (N_6102,N_5988,N_5995);
nor U6103 (N_6103,N_5925,N_5886);
nand U6104 (N_6104,N_5987,N_5968);
xor U6105 (N_6105,N_5928,N_5982);
and U6106 (N_6106,N_5965,N_5918);
nor U6107 (N_6107,N_5964,N_5945);
xor U6108 (N_6108,N_5976,N_5917);
and U6109 (N_6109,N_5919,N_5960);
xor U6110 (N_6110,N_5878,N_5975);
nor U6111 (N_6111,N_5970,N_5906);
nand U6112 (N_6112,N_5949,N_5879);
or U6113 (N_6113,N_5977,N_5921);
xnor U6114 (N_6114,N_5903,N_5982);
and U6115 (N_6115,N_5984,N_5905);
and U6116 (N_6116,N_5912,N_5955);
nor U6117 (N_6117,N_5987,N_5908);
and U6118 (N_6118,N_5960,N_5988);
xnor U6119 (N_6119,N_5954,N_5900);
nor U6120 (N_6120,N_5949,N_5963);
and U6121 (N_6121,N_5961,N_5881);
nor U6122 (N_6122,N_5972,N_5920);
nand U6123 (N_6123,N_5923,N_5925);
or U6124 (N_6124,N_5946,N_5975);
or U6125 (N_6125,N_6044,N_6051);
and U6126 (N_6126,N_6032,N_6041);
or U6127 (N_6127,N_6122,N_6031);
nand U6128 (N_6128,N_6116,N_6016);
or U6129 (N_6129,N_6118,N_6017);
nor U6130 (N_6130,N_6047,N_6106);
xnor U6131 (N_6131,N_6070,N_6124);
xor U6132 (N_6132,N_6095,N_6050);
nand U6133 (N_6133,N_6022,N_6102);
and U6134 (N_6134,N_6096,N_6072);
or U6135 (N_6135,N_6037,N_6113);
nand U6136 (N_6136,N_6093,N_6007);
nand U6137 (N_6137,N_6030,N_6056);
nor U6138 (N_6138,N_6052,N_6100);
nor U6139 (N_6139,N_6046,N_6002);
and U6140 (N_6140,N_6090,N_6006);
and U6141 (N_6141,N_6101,N_6001);
or U6142 (N_6142,N_6109,N_6099);
and U6143 (N_6143,N_6117,N_6059);
xnor U6144 (N_6144,N_6004,N_6062);
nor U6145 (N_6145,N_6103,N_6018);
xnor U6146 (N_6146,N_6073,N_6079);
nand U6147 (N_6147,N_6115,N_6028);
nand U6148 (N_6148,N_6107,N_6000);
xor U6149 (N_6149,N_6048,N_6038);
and U6150 (N_6150,N_6104,N_6091);
nor U6151 (N_6151,N_6045,N_6060);
nor U6152 (N_6152,N_6021,N_6008);
or U6153 (N_6153,N_6085,N_6058);
xor U6154 (N_6154,N_6066,N_6089);
and U6155 (N_6155,N_6123,N_6033);
xor U6156 (N_6156,N_6084,N_6092);
nor U6157 (N_6157,N_6086,N_6098);
or U6158 (N_6158,N_6081,N_6023);
nand U6159 (N_6159,N_6024,N_6035);
nand U6160 (N_6160,N_6043,N_6083);
xor U6161 (N_6161,N_6003,N_6121);
and U6162 (N_6162,N_6065,N_6039);
and U6163 (N_6163,N_6074,N_6049);
nand U6164 (N_6164,N_6080,N_6075);
or U6165 (N_6165,N_6071,N_6111);
nand U6166 (N_6166,N_6119,N_6042);
xnor U6167 (N_6167,N_6014,N_6015);
and U6168 (N_6168,N_6108,N_6114);
nand U6169 (N_6169,N_6069,N_6026);
and U6170 (N_6170,N_6067,N_6105);
and U6171 (N_6171,N_6076,N_6029);
and U6172 (N_6172,N_6011,N_6020);
nor U6173 (N_6173,N_6088,N_6013);
nor U6174 (N_6174,N_6057,N_6005);
or U6175 (N_6175,N_6012,N_6054);
xnor U6176 (N_6176,N_6068,N_6027);
and U6177 (N_6177,N_6061,N_6120);
nor U6178 (N_6178,N_6077,N_6082);
nand U6179 (N_6179,N_6064,N_6097);
or U6180 (N_6180,N_6025,N_6078);
xor U6181 (N_6181,N_6036,N_6019);
or U6182 (N_6182,N_6063,N_6110);
xnor U6183 (N_6183,N_6034,N_6087);
nor U6184 (N_6184,N_6094,N_6112);
nand U6185 (N_6185,N_6009,N_6053);
and U6186 (N_6186,N_6055,N_6040);
or U6187 (N_6187,N_6010,N_6086);
or U6188 (N_6188,N_6035,N_6114);
nand U6189 (N_6189,N_6123,N_6089);
nor U6190 (N_6190,N_6106,N_6014);
nor U6191 (N_6191,N_6053,N_6060);
and U6192 (N_6192,N_6027,N_6072);
nor U6193 (N_6193,N_6011,N_6058);
or U6194 (N_6194,N_6020,N_6121);
nor U6195 (N_6195,N_6015,N_6093);
nand U6196 (N_6196,N_6077,N_6003);
xnor U6197 (N_6197,N_6069,N_6091);
nand U6198 (N_6198,N_6110,N_6120);
nand U6199 (N_6199,N_6035,N_6111);
nor U6200 (N_6200,N_6082,N_6046);
xnor U6201 (N_6201,N_6107,N_6003);
or U6202 (N_6202,N_6084,N_6122);
nor U6203 (N_6203,N_6036,N_6006);
nand U6204 (N_6204,N_6028,N_6032);
nor U6205 (N_6205,N_6058,N_6003);
xnor U6206 (N_6206,N_6007,N_6009);
xor U6207 (N_6207,N_6037,N_6081);
and U6208 (N_6208,N_6007,N_6079);
nor U6209 (N_6209,N_6050,N_6119);
and U6210 (N_6210,N_6068,N_6120);
and U6211 (N_6211,N_6105,N_6036);
xnor U6212 (N_6212,N_6093,N_6043);
nor U6213 (N_6213,N_6038,N_6071);
and U6214 (N_6214,N_6045,N_6032);
nor U6215 (N_6215,N_6026,N_6019);
xor U6216 (N_6216,N_6023,N_6017);
xor U6217 (N_6217,N_6082,N_6102);
nor U6218 (N_6218,N_6073,N_6064);
xor U6219 (N_6219,N_6111,N_6106);
xor U6220 (N_6220,N_6096,N_6044);
nor U6221 (N_6221,N_6019,N_6081);
and U6222 (N_6222,N_6109,N_6028);
or U6223 (N_6223,N_6057,N_6000);
or U6224 (N_6224,N_6042,N_6100);
nand U6225 (N_6225,N_6102,N_6076);
xnor U6226 (N_6226,N_6043,N_6082);
or U6227 (N_6227,N_6119,N_6080);
or U6228 (N_6228,N_6109,N_6114);
nand U6229 (N_6229,N_6077,N_6096);
and U6230 (N_6230,N_6038,N_6069);
nand U6231 (N_6231,N_6012,N_6123);
and U6232 (N_6232,N_6011,N_6090);
and U6233 (N_6233,N_6033,N_6049);
or U6234 (N_6234,N_6093,N_6046);
and U6235 (N_6235,N_6051,N_6021);
nor U6236 (N_6236,N_6055,N_6025);
and U6237 (N_6237,N_6121,N_6060);
and U6238 (N_6238,N_6085,N_6008);
xor U6239 (N_6239,N_6110,N_6116);
nand U6240 (N_6240,N_6022,N_6008);
xor U6241 (N_6241,N_6081,N_6042);
nand U6242 (N_6242,N_6086,N_6054);
and U6243 (N_6243,N_6109,N_6021);
nand U6244 (N_6244,N_6092,N_6075);
xor U6245 (N_6245,N_6117,N_6110);
and U6246 (N_6246,N_6035,N_6000);
or U6247 (N_6247,N_6068,N_6023);
and U6248 (N_6248,N_6030,N_6063);
or U6249 (N_6249,N_6016,N_6040);
nand U6250 (N_6250,N_6237,N_6179);
and U6251 (N_6251,N_6204,N_6216);
xor U6252 (N_6252,N_6229,N_6202);
nand U6253 (N_6253,N_6157,N_6139);
nand U6254 (N_6254,N_6189,N_6165);
nand U6255 (N_6255,N_6129,N_6149);
nor U6256 (N_6256,N_6192,N_6242);
nor U6257 (N_6257,N_6147,N_6127);
xnor U6258 (N_6258,N_6188,N_6248);
or U6259 (N_6259,N_6158,N_6191);
and U6260 (N_6260,N_6238,N_6233);
or U6261 (N_6261,N_6214,N_6143);
or U6262 (N_6262,N_6225,N_6126);
or U6263 (N_6263,N_6141,N_6134);
and U6264 (N_6264,N_6222,N_6186);
nor U6265 (N_6265,N_6203,N_6249);
or U6266 (N_6266,N_6226,N_6136);
and U6267 (N_6267,N_6243,N_6241);
and U6268 (N_6268,N_6125,N_6180);
xnor U6269 (N_6269,N_6185,N_6239);
or U6270 (N_6270,N_6231,N_6151);
nand U6271 (N_6271,N_6246,N_6176);
nor U6272 (N_6272,N_6199,N_6144);
xor U6273 (N_6273,N_6245,N_6187);
nor U6274 (N_6274,N_6207,N_6206);
or U6275 (N_6275,N_6166,N_6142);
or U6276 (N_6276,N_6169,N_6168);
or U6277 (N_6277,N_6234,N_6128);
nor U6278 (N_6278,N_6181,N_6133);
nor U6279 (N_6279,N_6137,N_6212);
or U6280 (N_6280,N_6160,N_6244);
nor U6281 (N_6281,N_6175,N_6184);
nor U6282 (N_6282,N_6211,N_6172);
and U6283 (N_6283,N_6177,N_6193);
and U6284 (N_6284,N_6145,N_6223);
xor U6285 (N_6285,N_6135,N_6219);
nor U6286 (N_6286,N_6205,N_6235);
and U6287 (N_6287,N_6240,N_6218);
and U6288 (N_6288,N_6150,N_6162);
xnor U6289 (N_6289,N_6217,N_6155);
and U6290 (N_6290,N_6201,N_6228);
xnor U6291 (N_6291,N_6167,N_6153);
nand U6292 (N_6292,N_6190,N_6232);
nor U6293 (N_6293,N_6195,N_6163);
and U6294 (N_6294,N_6183,N_6224);
nand U6295 (N_6295,N_6140,N_6132);
xor U6296 (N_6296,N_6173,N_6148);
and U6297 (N_6297,N_6198,N_6159);
xnor U6298 (N_6298,N_6227,N_6220);
nand U6299 (N_6299,N_6174,N_6164);
or U6300 (N_6300,N_6152,N_6154);
and U6301 (N_6301,N_6208,N_6146);
nand U6302 (N_6302,N_6171,N_6196);
or U6303 (N_6303,N_6138,N_6182);
and U6304 (N_6304,N_6178,N_6221);
and U6305 (N_6305,N_6236,N_6213);
and U6306 (N_6306,N_6130,N_6131);
xor U6307 (N_6307,N_6170,N_6215);
nor U6308 (N_6308,N_6197,N_6161);
and U6309 (N_6309,N_6209,N_6194);
and U6310 (N_6310,N_6200,N_6210);
nand U6311 (N_6311,N_6230,N_6247);
or U6312 (N_6312,N_6156,N_6246);
nor U6313 (N_6313,N_6161,N_6206);
xnor U6314 (N_6314,N_6207,N_6228);
or U6315 (N_6315,N_6209,N_6162);
or U6316 (N_6316,N_6245,N_6205);
and U6317 (N_6317,N_6148,N_6224);
xnor U6318 (N_6318,N_6174,N_6188);
nor U6319 (N_6319,N_6213,N_6176);
or U6320 (N_6320,N_6211,N_6163);
or U6321 (N_6321,N_6158,N_6131);
or U6322 (N_6322,N_6222,N_6187);
xor U6323 (N_6323,N_6169,N_6193);
and U6324 (N_6324,N_6194,N_6171);
or U6325 (N_6325,N_6173,N_6131);
xor U6326 (N_6326,N_6212,N_6136);
nand U6327 (N_6327,N_6189,N_6186);
and U6328 (N_6328,N_6178,N_6152);
and U6329 (N_6329,N_6209,N_6217);
nand U6330 (N_6330,N_6141,N_6233);
or U6331 (N_6331,N_6206,N_6188);
xnor U6332 (N_6332,N_6163,N_6158);
or U6333 (N_6333,N_6226,N_6223);
or U6334 (N_6334,N_6232,N_6223);
xor U6335 (N_6335,N_6181,N_6190);
and U6336 (N_6336,N_6139,N_6198);
or U6337 (N_6337,N_6171,N_6170);
or U6338 (N_6338,N_6126,N_6222);
nor U6339 (N_6339,N_6242,N_6128);
nor U6340 (N_6340,N_6178,N_6164);
and U6341 (N_6341,N_6180,N_6140);
nor U6342 (N_6342,N_6162,N_6192);
or U6343 (N_6343,N_6165,N_6125);
nand U6344 (N_6344,N_6139,N_6203);
or U6345 (N_6345,N_6141,N_6208);
or U6346 (N_6346,N_6209,N_6195);
or U6347 (N_6347,N_6247,N_6176);
xor U6348 (N_6348,N_6218,N_6188);
and U6349 (N_6349,N_6237,N_6221);
or U6350 (N_6350,N_6133,N_6216);
xnor U6351 (N_6351,N_6234,N_6143);
and U6352 (N_6352,N_6157,N_6226);
or U6353 (N_6353,N_6150,N_6145);
or U6354 (N_6354,N_6242,N_6246);
and U6355 (N_6355,N_6172,N_6137);
xor U6356 (N_6356,N_6143,N_6197);
nor U6357 (N_6357,N_6233,N_6196);
nor U6358 (N_6358,N_6240,N_6196);
xnor U6359 (N_6359,N_6156,N_6174);
or U6360 (N_6360,N_6127,N_6243);
nor U6361 (N_6361,N_6141,N_6244);
or U6362 (N_6362,N_6234,N_6145);
or U6363 (N_6363,N_6203,N_6199);
nor U6364 (N_6364,N_6214,N_6246);
xor U6365 (N_6365,N_6225,N_6158);
nor U6366 (N_6366,N_6149,N_6152);
and U6367 (N_6367,N_6233,N_6201);
nor U6368 (N_6368,N_6196,N_6201);
xnor U6369 (N_6369,N_6222,N_6201);
xor U6370 (N_6370,N_6189,N_6143);
and U6371 (N_6371,N_6137,N_6153);
nand U6372 (N_6372,N_6157,N_6160);
xor U6373 (N_6373,N_6243,N_6168);
nand U6374 (N_6374,N_6199,N_6159);
or U6375 (N_6375,N_6348,N_6267);
nand U6376 (N_6376,N_6332,N_6261);
nor U6377 (N_6377,N_6263,N_6373);
or U6378 (N_6378,N_6346,N_6341);
and U6379 (N_6379,N_6277,N_6279);
or U6380 (N_6380,N_6276,N_6262);
nand U6381 (N_6381,N_6300,N_6347);
or U6382 (N_6382,N_6349,N_6252);
nor U6383 (N_6383,N_6318,N_6342);
nor U6384 (N_6384,N_6291,N_6359);
nor U6385 (N_6385,N_6372,N_6345);
nor U6386 (N_6386,N_6264,N_6284);
xnor U6387 (N_6387,N_6368,N_6288);
nor U6388 (N_6388,N_6358,N_6308);
or U6389 (N_6389,N_6369,N_6250);
nor U6390 (N_6390,N_6338,N_6370);
nor U6391 (N_6391,N_6272,N_6253);
xor U6392 (N_6392,N_6266,N_6283);
nand U6393 (N_6393,N_6336,N_6268);
nor U6394 (N_6394,N_6366,N_6323);
and U6395 (N_6395,N_6258,N_6357);
or U6396 (N_6396,N_6316,N_6313);
xor U6397 (N_6397,N_6304,N_6327);
and U6398 (N_6398,N_6321,N_6328);
and U6399 (N_6399,N_6367,N_6280);
and U6400 (N_6400,N_6364,N_6306);
xor U6401 (N_6401,N_6360,N_6324);
xor U6402 (N_6402,N_6312,N_6319);
nor U6403 (N_6403,N_6307,N_6297);
nand U6404 (N_6404,N_6270,N_6292);
nor U6405 (N_6405,N_6325,N_6285);
nand U6406 (N_6406,N_6309,N_6273);
nor U6407 (N_6407,N_6299,N_6329);
nand U6408 (N_6408,N_6260,N_6351);
xor U6409 (N_6409,N_6290,N_6289);
and U6410 (N_6410,N_6282,N_6259);
and U6411 (N_6411,N_6274,N_6343);
and U6412 (N_6412,N_6374,N_6340);
xnor U6413 (N_6413,N_6363,N_6337);
nor U6414 (N_6414,N_6256,N_6330);
and U6415 (N_6415,N_6305,N_6320);
nor U6416 (N_6416,N_6301,N_6296);
or U6417 (N_6417,N_6302,N_6371);
xor U6418 (N_6418,N_6317,N_6356);
nand U6419 (N_6419,N_6361,N_6335);
nand U6420 (N_6420,N_6278,N_6310);
nand U6421 (N_6421,N_6294,N_6293);
xnor U6422 (N_6422,N_6344,N_6315);
nor U6423 (N_6423,N_6286,N_6354);
nor U6424 (N_6424,N_6287,N_6311);
xnor U6425 (N_6425,N_6355,N_6251);
xnor U6426 (N_6426,N_6314,N_6269);
nand U6427 (N_6427,N_6322,N_6365);
or U6428 (N_6428,N_6257,N_6295);
nand U6429 (N_6429,N_6281,N_6271);
xnor U6430 (N_6430,N_6298,N_6303);
and U6431 (N_6431,N_6254,N_6326);
or U6432 (N_6432,N_6339,N_6275);
nor U6433 (N_6433,N_6334,N_6333);
and U6434 (N_6434,N_6362,N_6353);
xor U6435 (N_6435,N_6255,N_6350);
nor U6436 (N_6436,N_6352,N_6331);
or U6437 (N_6437,N_6265,N_6312);
or U6438 (N_6438,N_6288,N_6351);
nand U6439 (N_6439,N_6324,N_6262);
xor U6440 (N_6440,N_6332,N_6344);
xnor U6441 (N_6441,N_6286,N_6260);
nor U6442 (N_6442,N_6314,N_6283);
xor U6443 (N_6443,N_6313,N_6334);
nand U6444 (N_6444,N_6279,N_6264);
xor U6445 (N_6445,N_6331,N_6345);
nand U6446 (N_6446,N_6330,N_6309);
nand U6447 (N_6447,N_6305,N_6370);
nor U6448 (N_6448,N_6298,N_6325);
or U6449 (N_6449,N_6329,N_6333);
nor U6450 (N_6450,N_6365,N_6314);
nor U6451 (N_6451,N_6366,N_6269);
xor U6452 (N_6452,N_6322,N_6353);
and U6453 (N_6453,N_6368,N_6287);
nor U6454 (N_6454,N_6271,N_6299);
nor U6455 (N_6455,N_6310,N_6273);
and U6456 (N_6456,N_6360,N_6331);
or U6457 (N_6457,N_6351,N_6339);
or U6458 (N_6458,N_6313,N_6364);
nor U6459 (N_6459,N_6283,N_6273);
and U6460 (N_6460,N_6345,N_6361);
nand U6461 (N_6461,N_6275,N_6267);
xnor U6462 (N_6462,N_6373,N_6308);
xnor U6463 (N_6463,N_6280,N_6295);
nand U6464 (N_6464,N_6308,N_6320);
nor U6465 (N_6465,N_6358,N_6272);
xor U6466 (N_6466,N_6325,N_6296);
nand U6467 (N_6467,N_6373,N_6284);
nand U6468 (N_6468,N_6263,N_6345);
xor U6469 (N_6469,N_6332,N_6351);
nor U6470 (N_6470,N_6275,N_6373);
and U6471 (N_6471,N_6320,N_6283);
xor U6472 (N_6472,N_6303,N_6262);
nand U6473 (N_6473,N_6313,N_6278);
or U6474 (N_6474,N_6257,N_6270);
nand U6475 (N_6475,N_6323,N_6255);
and U6476 (N_6476,N_6263,N_6278);
nor U6477 (N_6477,N_6299,N_6366);
xor U6478 (N_6478,N_6339,N_6323);
or U6479 (N_6479,N_6370,N_6302);
xnor U6480 (N_6480,N_6360,N_6257);
or U6481 (N_6481,N_6295,N_6374);
xor U6482 (N_6482,N_6324,N_6288);
xnor U6483 (N_6483,N_6284,N_6268);
and U6484 (N_6484,N_6265,N_6332);
xnor U6485 (N_6485,N_6261,N_6283);
nand U6486 (N_6486,N_6288,N_6318);
xnor U6487 (N_6487,N_6328,N_6275);
or U6488 (N_6488,N_6328,N_6286);
or U6489 (N_6489,N_6360,N_6285);
nor U6490 (N_6490,N_6362,N_6266);
or U6491 (N_6491,N_6366,N_6254);
nand U6492 (N_6492,N_6369,N_6304);
nand U6493 (N_6493,N_6316,N_6264);
nand U6494 (N_6494,N_6271,N_6324);
nor U6495 (N_6495,N_6303,N_6353);
and U6496 (N_6496,N_6258,N_6268);
nand U6497 (N_6497,N_6293,N_6349);
or U6498 (N_6498,N_6327,N_6283);
nor U6499 (N_6499,N_6287,N_6371);
or U6500 (N_6500,N_6460,N_6458);
xor U6501 (N_6501,N_6435,N_6493);
xnor U6502 (N_6502,N_6413,N_6483);
xnor U6503 (N_6503,N_6439,N_6476);
or U6504 (N_6504,N_6433,N_6396);
or U6505 (N_6505,N_6417,N_6411);
nor U6506 (N_6506,N_6447,N_6495);
nand U6507 (N_6507,N_6418,N_6389);
and U6508 (N_6508,N_6406,N_6446);
xnor U6509 (N_6509,N_6395,N_6443);
or U6510 (N_6510,N_6393,N_6410);
or U6511 (N_6511,N_6390,N_6400);
nor U6512 (N_6512,N_6408,N_6422);
nand U6513 (N_6513,N_6394,N_6480);
and U6514 (N_6514,N_6398,N_6428);
and U6515 (N_6515,N_6386,N_6383);
or U6516 (N_6516,N_6401,N_6424);
xnor U6517 (N_6517,N_6463,N_6444);
or U6518 (N_6518,N_6440,N_6486);
xor U6519 (N_6519,N_6414,N_6430);
xor U6520 (N_6520,N_6482,N_6420);
and U6521 (N_6521,N_6454,N_6379);
xnor U6522 (N_6522,N_6416,N_6488);
and U6523 (N_6523,N_6481,N_6491);
nor U6524 (N_6524,N_6475,N_6478);
and U6525 (N_6525,N_6432,N_6442);
nor U6526 (N_6526,N_6489,N_6437);
and U6527 (N_6527,N_6397,N_6384);
nor U6528 (N_6528,N_6455,N_6497);
xnor U6529 (N_6529,N_6419,N_6388);
nor U6530 (N_6530,N_6387,N_6452);
xnor U6531 (N_6531,N_6376,N_6399);
xnor U6532 (N_6532,N_6474,N_6470);
xor U6533 (N_6533,N_6380,N_6453);
and U6534 (N_6534,N_6425,N_6464);
nor U6535 (N_6535,N_6448,N_6403);
nand U6536 (N_6536,N_6492,N_6467);
xnor U6537 (N_6537,N_6471,N_6485);
or U6538 (N_6538,N_6459,N_6404);
xnor U6539 (N_6539,N_6484,N_6494);
and U6540 (N_6540,N_6426,N_6407);
nand U6541 (N_6541,N_6465,N_6469);
nand U6542 (N_6542,N_6479,N_6423);
nand U6543 (N_6543,N_6441,N_6496);
or U6544 (N_6544,N_6449,N_6402);
nor U6545 (N_6545,N_6429,N_6436);
xor U6546 (N_6546,N_6462,N_6405);
nor U6547 (N_6547,N_6473,N_6392);
or U6548 (N_6548,N_6472,N_6438);
and U6549 (N_6549,N_6431,N_6498);
xnor U6550 (N_6550,N_6461,N_6499);
nand U6551 (N_6551,N_6466,N_6490);
nor U6552 (N_6552,N_6377,N_6385);
or U6553 (N_6553,N_6409,N_6445);
and U6554 (N_6554,N_6427,N_6457);
and U6555 (N_6555,N_6391,N_6451);
nor U6556 (N_6556,N_6412,N_6415);
xnor U6557 (N_6557,N_6375,N_6382);
nor U6558 (N_6558,N_6477,N_6456);
and U6559 (N_6559,N_6487,N_6434);
xor U6560 (N_6560,N_6450,N_6378);
xnor U6561 (N_6561,N_6381,N_6421);
nand U6562 (N_6562,N_6468,N_6396);
xor U6563 (N_6563,N_6431,N_6378);
or U6564 (N_6564,N_6449,N_6469);
xnor U6565 (N_6565,N_6421,N_6485);
and U6566 (N_6566,N_6480,N_6462);
or U6567 (N_6567,N_6487,N_6442);
nand U6568 (N_6568,N_6408,N_6486);
or U6569 (N_6569,N_6413,N_6451);
nand U6570 (N_6570,N_6437,N_6423);
and U6571 (N_6571,N_6466,N_6409);
nand U6572 (N_6572,N_6458,N_6482);
or U6573 (N_6573,N_6480,N_6423);
xor U6574 (N_6574,N_6488,N_6482);
xnor U6575 (N_6575,N_6377,N_6388);
and U6576 (N_6576,N_6462,N_6401);
nor U6577 (N_6577,N_6427,N_6496);
nor U6578 (N_6578,N_6452,N_6426);
xor U6579 (N_6579,N_6491,N_6446);
nand U6580 (N_6580,N_6452,N_6411);
or U6581 (N_6581,N_6375,N_6397);
or U6582 (N_6582,N_6409,N_6404);
nand U6583 (N_6583,N_6426,N_6495);
and U6584 (N_6584,N_6426,N_6490);
nor U6585 (N_6585,N_6485,N_6470);
or U6586 (N_6586,N_6481,N_6450);
and U6587 (N_6587,N_6456,N_6409);
and U6588 (N_6588,N_6450,N_6490);
and U6589 (N_6589,N_6495,N_6484);
nand U6590 (N_6590,N_6455,N_6444);
nor U6591 (N_6591,N_6462,N_6377);
or U6592 (N_6592,N_6488,N_6398);
and U6593 (N_6593,N_6454,N_6434);
xnor U6594 (N_6594,N_6423,N_6470);
or U6595 (N_6595,N_6414,N_6431);
or U6596 (N_6596,N_6384,N_6427);
or U6597 (N_6597,N_6483,N_6380);
nand U6598 (N_6598,N_6483,N_6444);
xnor U6599 (N_6599,N_6440,N_6477);
nand U6600 (N_6600,N_6410,N_6453);
or U6601 (N_6601,N_6486,N_6429);
nand U6602 (N_6602,N_6440,N_6384);
or U6603 (N_6603,N_6469,N_6402);
or U6604 (N_6604,N_6436,N_6380);
xor U6605 (N_6605,N_6443,N_6397);
nand U6606 (N_6606,N_6497,N_6403);
or U6607 (N_6607,N_6390,N_6462);
xnor U6608 (N_6608,N_6497,N_6496);
nor U6609 (N_6609,N_6494,N_6485);
nor U6610 (N_6610,N_6399,N_6432);
and U6611 (N_6611,N_6470,N_6439);
or U6612 (N_6612,N_6459,N_6474);
nand U6613 (N_6613,N_6384,N_6466);
or U6614 (N_6614,N_6470,N_6454);
or U6615 (N_6615,N_6433,N_6390);
nand U6616 (N_6616,N_6435,N_6394);
xor U6617 (N_6617,N_6441,N_6440);
and U6618 (N_6618,N_6420,N_6436);
or U6619 (N_6619,N_6415,N_6377);
xor U6620 (N_6620,N_6436,N_6408);
nor U6621 (N_6621,N_6396,N_6459);
xor U6622 (N_6622,N_6431,N_6493);
and U6623 (N_6623,N_6428,N_6474);
and U6624 (N_6624,N_6474,N_6421);
or U6625 (N_6625,N_6536,N_6501);
nor U6626 (N_6626,N_6577,N_6520);
and U6627 (N_6627,N_6567,N_6537);
or U6628 (N_6628,N_6571,N_6586);
xor U6629 (N_6629,N_6500,N_6556);
and U6630 (N_6630,N_6583,N_6508);
nand U6631 (N_6631,N_6522,N_6615);
xnor U6632 (N_6632,N_6527,N_6620);
xnor U6633 (N_6633,N_6598,N_6621);
xor U6634 (N_6634,N_6574,N_6516);
or U6635 (N_6635,N_6566,N_6543);
and U6636 (N_6636,N_6570,N_6582);
nand U6637 (N_6637,N_6563,N_6531);
and U6638 (N_6638,N_6575,N_6603);
and U6639 (N_6639,N_6573,N_6544);
and U6640 (N_6640,N_6529,N_6504);
nor U6641 (N_6641,N_6613,N_6513);
and U6642 (N_6642,N_6611,N_6589);
xnor U6643 (N_6643,N_6525,N_6509);
nor U6644 (N_6644,N_6532,N_6580);
nor U6645 (N_6645,N_6618,N_6600);
xnor U6646 (N_6646,N_6610,N_6534);
or U6647 (N_6647,N_6590,N_6503);
or U6648 (N_6648,N_6609,N_6594);
xnor U6649 (N_6649,N_6507,N_6550);
xnor U6650 (N_6650,N_6602,N_6521);
and U6651 (N_6651,N_6581,N_6555);
and U6652 (N_6652,N_6549,N_6542);
nand U6653 (N_6653,N_6524,N_6616);
xor U6654 (N_6654,N_6517,N_6514);
or U6655 (N_6655,N_6596,N_6540);
xor U6656 (N_6656,N_6576,N_6535);
xnor U6657 (N_6657,N_6617,N_6565);
nand U6658 (N_6658,N_6519,N_6623);
nand U6659 (N_6659,N_6606,N_6528);
or U6660 (N_6660,N_6558,N_6579);
nor U6661 (N_6661,N_6601,N_6551);
nand U6662 (N_6662,N_6530,N_6533);
nor U6663 (N_6663,N_6523,N_6548);
nand U6664 (N_6664,N_6541,N_6510);
nand U6665 (N_6665,N_6593,N_6624);
xor U6666 (N_6666,N_6614,N_6560);
nand U6667 (N_6667,N_6553,N_6506);
nor U6668 (N_6668,N_6545,N_6585);
xor U6669 (N_6669,N_6588,N_6568);
and U6670 (N_6670,N_6612,N_6538);
or U6671 (N_6671,N_6554,N_6512);
nand U6672 (N_6672,N_6546,N_6604);
and U6673 (N_6673,N_6599,N_6539);
and U6674 (N_6674,N_6595,N_6547);
nor U6675 (N_6675,N_6502,N_6557);
nor U6676 (N_6676,N_6597,N_6526);
nand U6677 (N_6677,N_6552,N_6578);
nor U6678 (N_6678,N_6608,N_6559);
xor U6679 (N_6679,N_6562,N_6518);
and U6680 (N_6680,N_6619,N_6515);
xnor U6681 (N_6681,N_6561,N_6591);
nand U6682 (N_6682,N_6584,N_6607);
nor U6683 (N_6683,N_6569,N_6592);
and U6684 (N_6684,N_6505,N_6605);
and U6685 (N_6685,N_6622,N_6511);
nor U6686 (N_6686,N_6572,N_6564);
or U6687 (N_6687,N_6587,N_6558);
and U6688 (N_6688,N_6609,N_6621);
and U6689 (N_6689,N_6575,N_6559);
nand U6690 (N_6690,N_6588,N_6532);
and U6691 (N_6691,N_6597,N_6525);
xor U6692 (N_6692,N_6527,N_6546);
and U6693 (N_6693,N_6574,N_6608);
and U6694 (N_6694,N_6581,N_6616);
xnor U6695 (N_6695,N_6618,N_6512);
or U6696 (N_6696,N_6540,N_6519);
xor U6697 (N_6697,N_6590,N_6541);
or U6698 (N_6698,N_6581,N_6614);
nand U6699 (N_6699,N_6540,N_6601);
and U6700 (N_6700,N_6592,N_6528);
xor U6701 (N_6701,N_6600,N_6568);
nand U6702 (N_6702,N_6516,N_6578);
xnor U6703 (N_6703,N_6592,N_6517);
or U6704 (N_6704,N_6615,N_6533);
or U6705 (N_6705,N_6515,N_6600);
nor U6706 (N_6706,N_6620,N_6579);
nor U6707 (N_6707,N_6601,N_6573);
nor U6708 (N_6708,N_6595,N_6604);
nor U6709 (N_6709,N_6613,N_6595);
and U6710 (N_6710,N_6549,N_6607);
nor U6711 (N_6711,N_6500,N_6534);
or U6712 (N_6712,N_6591,N_6602);
nor U6713 (N_6713,N_6593,N_6558);
xnor U6714 (N_6714,N_6539,N_6623);
xor U6715 (N_6715,N_6520,N_6513);
and U6716 (N_6716,N_6507,N_6524);
nor U6717 (N_6717,N_6612,N_6511);
and U6718 (N_6718,N_6520,N_6526);
and U6719 (N_6719,N_6544,N_6500);
nand U6720 (N_6720,N_6575,N_6530);
and U6721 (N_6721,N_6505,N_6517);
or U6722 (N_6722,N_6530,N_6501);
and U6723 (N_6723,N_6605,N_6544);
and U6724 (N_6724,N_6595,N_6523);
and U6725 (N_6725,N_6560,N_6553);
xor U6726 (N_6726,N_6542,N_6611);
nand U6727 (N_6727,N_6604,N_6544);
or U6728 (N_6728,N_6572,N_6563);
xnor U6729 (N_6729,N_6610,N_6502);
or U6730 (N_6730,N_6570,N_6511);
nand U6731 (N_6731,N_6607,N_6520);
or U6732 (N_6732,N_6567,N_6534);
xor U6733 (N_6733,N_6564,N_6596);
nor U6734 (N_6734,N_6525,N_6549);
xor U6735 (N_6735,N_6615,N_6573);
nor U6736 (N_6736,N_6555,N_6510);
nor U6737 (N_6737,N_6554,N_6558);
xor U6738 (N_6738,N_6572,N_6587);
and U6739 (N_6739,N_6530,N_6606);
or U6740 (N_6740,N_6580,N_6576);
nand U6741 (N_6741,N_6536,N_6549);
or U6742 (N_6742,N_6615,N_6568);
or U6743 (N_6743,N_6520,N_6564);
xnor U6744 (N_6744,N_6540,N_6604);
and U6745 (N_6745,N_6514,N_6576);
nand U6746 (N_6746,N_6542,N_6577);
and U6747 (N_6747,N_6591,N_6548);
nor U6748 (N_6748,N_6587,N_6575);
or U6749 (N_6749,N_6515,N_6584);
nor U6750 (N_6750,N_6684,N_6726);
and U6751 (N_6751,N_6695,N_6625);
xnor U6752 (N_6752,N_6730,N_6655);
or U6753 (N_6753,N_6643,N_6629);
nor U6754 (N_6754,N_6741,N_6649);
and U6755 (N_6755,N_6687,N_6708);
nand U6756 (N_6756,N_6636,N_6650);
and U6757 (N_6757,N_6642,N_6637);
nor U6758 (N_6758,N_6740,N_6644);
nor U6759 (N_6759,N_6679,N_6694);
xor U6760 (N_6760,N_6676,N_6685);
or U6761 (N_6761,N_6729,N_6725);
nor U6762 (N_6762,N_6723,N_6657);
nor U6763 (N_6763,N_6709,N_6630);
and U6764 (N_6764,N_6715,N_6666);
or U6765 (N_6765,N_6631,N_6732);
nand U6766 (N_6766,N_6711,N_6712);
and U6767 (N_6767,N_6646,N_6659);
or U6768 (N_6768,N_6633,N_6705);
and U6769 (N_6769,N_6736,N_6739);
xor U6770 (N_6770,N_6737,N_6647);
xnor U6771 (N_6771,N_6743,N_6640);
nor U6772 (N_6772,N_6742,N_6671);
nand U6773 (N_6773,N_6645,N_6721);
nand U6774 (N_6774,N_6717,N_6677);
nor U6775 (N_6775,N_6716,N_6674);
nor U6776 (N_6776,N_6697,N_6692);
nor U6777 (N_6777,N_6704,N_6735);
nor U6778 (N_6778,N_6749,N_6652);
and U6779 (N_6779,N_6673,N_6691);
and U6780 (N_6780,N_6648,N_6672);
nor U6781 (N_6781,N_6731,N_6638);
nand U6782 (N_6782,N_6722,N_6664);
or U6783 (N_6783,N_6706,N_6653);
xor U6784 (N_6784,N_6627,N_6703);
or U6785 (N_6785,N_6701,N_6665);
xor U6786 (N_6786,N_6713,N_6696);
nand U6787 (N_6787,N_6700,N_6693);
and U6788 (N_6788,N_6724,N_6675);
or U6789 (N_6789,N_6661,N_6682);
and U6790 (N_6790,N_6747,N_6688);
nand U6791 (N_6791,N_6718,N_6746);
nand U6792 (N_6792,N_6680,N_6707);
or U6793 (N_6793,N_6727,N_6670);
xnor U6794 (N_6794,N_6626,N_6719);
nor U6795 (N_6795,N_6641,N_6667);
or U6796 (N_6796,N_6698,N_6734);
nand U6797 (N_6797,N_6651,N_6635);
or U6798 (N_6798,N_6686,N_6710);
nor U6799 (N_6799,N_6720,N_6660);
and U6800 (N_6800,N_6690,N_6733);
nor U6801 (N_6801,N_6654,N_6662);
xor U6802 (N_6802,N_6668,N_6663);
nand U6803 (N_6803,N_6656,N_6689);
or U6804 (N_6804,N_6744,N_6632);
nand U6805 (N_6805,N_6745,N_6628);
nand U6806 (N_6806,N_6669,N_6658);
and U6807 (N_6807,N_6714,N_6678);
nand U6808 (N_6808,N_6681,N_6683);
or U6809 (N_6809,N_6634,N_6702);
xnor U6810 (N_6810,N_6699,N_6748);
or U6811 (N_6811,N_6728,N_6738);
xor U6812 (N_6812,N_6639,N_6705);
nand U6813 (N_6813,N_6711,N_6677);
xnor U6814 (N_6814,N_6641,N_6625);
nor U6815 (N_6815,N_6665,N_6690);
xnor U6816 (N_6816,N_6741,N_6648);
or U6817 (N_6817,N_6745,N_6746);
or U6818 (N_6818,N_6713,N_6732);
nor U6819 (N_6819,N_6735,N_6721);
nor U6820 (N_6820,N_6689,N_6730);
nand U6821 (N_6821,N_6671,N_6699);
or U6822 (N_6822,N_6642,N_6628);
xor U6823 (N_6823,N_6731,N_6660);
nand U6824 (N_6824,N_6725,N_6740);
nand U6825 (N_6825,N_6744,N_6686);
xnor U6826 (N_6826,N_6663,N_6625);
or U6827 (N_6827,N_6641,N_6729);
or U6828 (N_6828,N_6724,N_6740);
or U6829 (N_6829,N_6672,N_6662);
and U6830 (N_6830,N_6630,N_6723);
nand U6831 (N_6831,N_6707,N_6682);
and U6832 (N_6832,N_6718,N_6731);
or U6833 (N_6833,N_6651,N_6648);
or U6834 (N_6834,N_6722,N_6684);
nor U6835 (N_6835,N_6669,N_6645);
and U6836 (N_6836,N_6667,N_6723);
and U6837 (N_6837,N_6678,N_6748);
or U6838 (N_6838,N_6678,N_6643);
xnor U6839 (N_6839,N_6681,N_6652);
nand U6840 (N_6840,N_6700,N_6682);
nand U6841 (N_6841,N_6705,N_6718);
nor U6842 (N_6842,N_6743,N_6712);
or U6843 (N_6843,N_6634,N_6668);
nand U6844 (N_6844,N_6720,N_6727);
and U6845 (N_6845,N_6717,N_6699);
or U6846 (N_6846,N_6733,N_6639);
or U6847 (N_6847,N_6703,N_6673);
nand U6848 (N_6848,N_6738,N_6734);
nor U6849 (N_6849,N_6749,N_6668);
and U6850 (N_6850,N_6673,N_6726);
nand U6851 (N_6851,N_6704,N_6736);
and U6852 (N_6852,N_6735,N_6710);
xnor U6853 (N_6853,N_6664,N_6690);
nand U6854 (N_6854,N_6629,N_6670);
nor U6855 (N_6855,N_6640,N_6654);
xor U6856 (N_6856,N_6681,N_6688);
nor U6857 (N_6857,N_6640,N_6745);
nand U6858 (N_6858,N_6719,N_6722);
xnor U6859 (N_6859,N_6743,N_6665);
or U6860 (N_6860,N_6696,N_6691);
nand U6861 (N_6861,N_6637,N_6732);
xnor U6862 (N_6862,N_6707,N_6649);
nor U6863 (N_6863,N_6669,N_6726);
xnor U6864 (N_6864,N_6718,N_6674);
or U6865 (N_6865,N_6684,N_6701);
and U6866 (N_6866,N_6695,N_6745);
or U6867 (N_6867,N_6647,N_6727);
nand U6868 (N_6868,N_6744,N_6638);
nand U6869 (N_6869,N_6688,N_6635);
nor U6870 (N_6870,N_6639,N_6673);
and U6871 (N_6871,N_6723,N_6631);
or U6872 (N_6872,N_6687,N_6635);
nand U6873 (N_6873,N_6628,N_6721);
and U6874 (N_6874,N_6730,N_6649);
and U6875 (N_6875,N_6835,N_6823);
or U6876 (N_6876,N_6818,N_6755);
nor U6877 (N_6877,N_6766,N_6778);
or U6878 (N_6878,N_6845,N_6779);
or U6879 (N_6879,N_6750,N_6837);
xor U6880 (N_6880,N_6858,N_6792);
or U6881 (N_6881,N_6799,N_6828);
and U6882 (N_6882,N_6869,N_6795);
or U6883 (N_6883,N_6859,N_6809);
nand U6884 (N_6884,N_6788,N_6784);
or U6885 (N_6885,N_6759,N_6761);
nand U6886 (N_6886,N_6826,N_6827);
or U6887 (N_6887,N_6786,N_6820);
or U6888 (N_6888,N_6839,N_6781);
nor U6889 (N_6889,N_6861,N_6753);
or U6890 (N_6890,N_6851,N_6829);
and U6891 (N_6891,N_6842,N_6873);
xor U6892 (N_6892,N_6825,N_6773);
nand U6893 (N_6893,N_6782,N_6850);
or U6894 (N_6894,N_6760,N_6854);
nand U6895 (N_6895,N_6870,N_6814);
nor U6896 (N_6896,N_6840,N_6796);
nor U6897 (N_6897,N_6806,N_6774);
xnor U6898 (N_6898,N_6868,N_6758);
nor U6899 (N_6899,N_6821,N_6765);
and U6900 (N_6900,N_6871,N_6816);
and U6901 (N_6901,N_6857,N_6769);
nor U6902 (N_6902,N_6803,N_6756);
and U6903 (N_6903,N_6785,N_6810);
nand U6904 (N_6904,N_6844,N_6800);
nand U6905 (N_6905,N_6780,N_6768);
xnor U6906 (N_6906,N_6772,N_6824);
and U6907 (N_6907,N_6860,N_6808);
or U6908 (N_6908,N_6811,N_6831);
nand U6909 (N_6909,N_6754,N_6874);
xor U6910 (N_6910,N_6791,N_6863);
nor U6911 (N_6911,N_6752,N_6865);
and U6912 (N_6912,N_6776,N_6864);
or U6913 (N_6913,N_6775,N_6751);
and U6914 (N_6914,N_6853,N_6771);
or U6915 (N_6915,N_6841,N_6833);
xnor U6916 (N_6916,N_6856,N_6767);
nand U6917 (N_6917,N_6793,N_6802);
nand U6918 (N_6918,N_6855,N_6830);
nor U6919 (N_6919,N_6813,N_6801);
nand U6920 (N_6920,N_6797,N_6783);
nand U6921 (N_6921,N_6789,N_6867);
nand U6922 (N_6922,N_6838,N_6852);
or U6923 (N_6923,N_6798,N_6819);
or U6924 (N_6924,N_6817,N_6846);
and U6925 (N_6925,N_6843,N_6847);
nor U6926 (N_6926,N_6763,N_6815);
and U6927 (N_6927,N_6836,N_6787);
or U6928 (N_6928,N_6812,N_6794);
and U6929 (N_6929,N_6834,N_6790);
xor U6930 (N_6930,N_6805,N_6804);
nor U6931 (N_6931,N_6764,N_6807);
xnor U6932 (N_6932,N_6849,N_6762);
or U6933 (N_6933,N_6822,N_6757);
nand U6934 (N_6934,N_6848,N_6770);
nor U6935 (N_6935,N_6872,N_6862);
or U6936 (N_6936,N_6777,N_6832);
and U6937 (N_6937,N_6866,N_6830);
nand U6938 (N_6938,N_6803,N_6798);
xor U6939 (N_6939,N_6869,N_6825);
xnor U6940 (N_6940,N_6866,N_6865);
or U6941 (N_6941,N_6823,N_6813);
and U6942 (N_6942,N_6754,N_6851);
nor U6943 (N_6943,N_6801,N_6768);
nand U6944 (N_6944,N_6779,N_6782);
and U6945 (N_6945,N_6839,N_6829);
nand U6946 (N_6946,N_6788,N_6754);
nand U6947 (N_6947,N_6772,N_6840);
and U6948 (N_6948,N_6796,N_6802);
xnor U6949 (N_6949,N_6863,N_6850);
and U6950 (N_6950,N_6759,N_6836);
and U6951 (N_6951,N_6820,N_6808);
and U6952 (N_6952,N_6777,N_6789);
and U6953 (N_6953,N_6793,N_6800);
or U6954 (N_6954,N_6789,N_6874);
xor U6955 (N_6955,N_6859,N_6838);
and U6956 (N_6956,N_6868,N_6839);
nand U6957 (N_6957,N_6793,N_6856);
or U6958 (N_6958,N_6784,N_6830);
or U6959 (N_6959,N_6786,N_6793);
nor U6960 (N_6960,N_6819,N_6866);
xnor U6961 (N_6961,N_6853,N_6763);
nor U6962 (N_6962,N_6797,N_6766);
nand U6963 (N_6963,N_6761,N_6855);
xnor U6964 (N_6964,N_6838,N_6847);
xnor U6965 (N_6965,N_6826,N_6858);
nor U6966 (N_6966,N_6771,N_6809);
or U6967 (N_6967,N_6811,N_6849);
and U6968 (N_6968,N_6798,N_6765);
and U6969 (N_6969,N_6862,N_6849);
xor U6970 (N_6970,N_6866,N_6806);
xor U6971 (N_6971,N_6761,N_6863);
or U6972 (N_6972,N_6856,N_6872);
or U6973 (N_6973,N_6839,N_6837);
nand U6974 (N_6974,N_6856,N_6843);
and U6975 (N_6975,N_6873,N_6788);
nand U6976 (N_6976,N_6861,N_6779);
or U6977 (N_6977,N_6765,N_6757);
and U6978 (N_6978,N_6799,N_6759);
or U6979 (N_6979,N_6799,N_6791);
nor U6980 (N_6980,N_6870,N_6864);
nand U6981 (N_6981,N_6774,N_6812);
xor U6982 (N_6982,N_6835,N_6778);
or U6983 (N_6983,N_6837,N_6775);
nor U6984 (N_6984,N_6781,N_6759);
nor U6985 (N_6985,N_6823,N_6830);
nand U6986 (N_6986,N_6831,N_6764);
nand U6987 (N_6987,N_6763,N_6767);
or U6988 (N_6988,N_6830,N_6865);
and U6989 (N_6989,N_6816,N_6781);
xnor U6990 (N_6990,N_6814,N_6851);
nor U6991 (N_6991,N_6855,N_6842);
and U6992 (N_6992,N_6870,N_6773);
and U6993 (N_6993,N_6847,N_6768);
xnor U6994 (N_6994,N_6818,N_6793);
or U6995 (N_6995,N_6812,N_6845);
and U6996 (N_6996,N_6765,N_6861);
or U6997 (N_6997,N_6848,N_6862);
nor U6998 (N_6998,N_6798,N_6757);
or U6999 (N_6999,N_6784,N_6847);
nand U7000 (N_7000,N_6955,N_6887);
nor U7001 (N_7001,N_6928,N_6999);
nand U7002 (N_7002,N_6897,N_6882);
and U7003 (N_7003,N_6929,N_6995);
xor U7004 (N_7004,N_6964,N_6930);
nor U7005 (N_7005,N_6940,N_6919);
nand U7006 (N_7006,N_6987,N_6990);
nor U7007 (N_7007,N_6977,N_6970);
xnor U7008 (N_7008,N_6971,N_6960);
and U7009 (N_7009,N_6949,N_6993);
or U7010 (N_7010,N_6902,N_6876);
and U7011 (N_7011,N_6913,N_6989);
xor U7012 (N_7012,N_6886,N_6905);
and U7013 (N_7013,N_6956,N_6908);
xnor U7014 (N_7014,N_6877,N_6946);
or U7015 (N_7015,N_6957,N_6980);
nand U7016 (N_7016,N_6975,N_6927);
and U7017 (N_7017,N_6998,N_6951);
xnor U7018 (N_7018,N_6948,N_6896);
xor U7019 (N_7019,N_6910,N_6954);
xor U7020 (N_7020,N_6917,N_6879);
or U7021 (N_7021,N_6921,N_6965);
or U7022 (N_7022,N_6922,N_6944);
xnor U7023 (N_7023,N_6994,N_6932);
xor U7024 (N_7024,N_6972,N_6942);
nor U7025 (N_7025,N_6924,N_6996);
xor U7026 (N_7026,N_6939,N_6903);
xor U7027 (N_7027,N_6991,N_6976);
nand U7028 (N_7028,N_6935,N_6968);
nand U7029 (N_7029,N_6880,N_6883);
or U7030 (N_7030,N_6936,N_6969);
nand U7031 (N_7031,N_6881,N_6981);
xnor U7032 (N_7032,N_6901,N_6875);
and U7033 (N_7033,N_6904,N_6982);
xnor U7034 (N_7034,N_6938,N_6978);
and U7035 (N_7035,N_6952,N_6988);
xor U7036 (N_7036,N_6899,N_6985);
and U7037 (N_7037,N_6974,N_6885);
or U7038 (N_7038,N_6892,N_6888);
xor U7039 (N_7039,N_6966,N_6967);
and U7040 (N_7040,N_6884,N_6943);
and U7041 (N_7041,N_6933,N_6894);
and U7042 (N_7042,N_6926,N_6915);
xor U7043 (N_7043,N_6900,N_6898);
nand U7044 (N_7044,N_6914,N_6992);
and U7045 (N_7045,N_6893,N_6937);
nand U7046 (N_7046,N_6983,N_6906);
nand U7047 (N_7047,N_6920,N_6947);
or U7048 (N_7048,N_6895,N_6959);
nor U7049 (N_7049,N_6963,N_6912);
nand U7050 (N_7050,N_6950,N_6941);
nor U7051 (N_7051,N_6931,N_6918);
nor U7052 (N_7052,N_6958,N_6909);
nand U7053 (N_7053,N_6916,N_6891);
or U7054 (N_7054,N_6889,N_6979);
or U7055 (N_7055,N_6890,N_6984);
nor U7056 (N_7056,N_6997,N_6986);
and U7057 (N_7057,N_6973,N_6923);
nor U7058 (N_7058,N_6934,N_6907);
and U7059 (N_7059,N_6945,N_6925);
nor U7060 (N_7060,N_6911,N_6962);
xor U7061 (N_7061,N_6878,N_6953);
nor U7062 (N_7062,N_6961,N_6951);
nand U7063 (N_7063,N_6974,N_6880);
or U7064 (N_7064,N_6935,N_6983);
or U7065 (N_7065,N_6987,N_6963);
xnor U7066 (N_7066,N_6881,N_6933);
nor U7067 (N_7067,N_6982,N_6940);
xor U7068 (N_7068,N_6936,N_6957);
or U7069 (N_7069,N_6984,N_6975);
and U7070 (N_7070,N_6903,N_6919);
or U7071 (N_7071,N_6915,N_6894);
xor U7072 (N_7072,N_6986,N_6880);
nand U7073 (N_7073,N_6952,N_6927);
and U7074 (N_7074,N_6927,N_6885);
nand U7075 (N_7075,N_6896,N_6925);
xor U7076 (N_7076,N_6904,N_6887);
xnor U7077 (N_7077,N_6932,N_6880);
nand U7078 (N_7078,N_6995,N_6893);
nand U7079 (N_7079,N_6895,N_6998);
or U7080 (N_7080,N_6991,N_6903);
or U7081 (N_7081,N_6877,N_6998);
or U7082 (N_7082,N_6924,N_6948);
xnor U7083 (N_7083,N_6996,N_6971);
and U7084 (N_7084,N_6981,N_6948);
or U7085 (N_7085,N_6898,N_6956);
and U7086 (N_7086,N_6942,N_6879);
nor U7087 (N_7087,N_6878,N_6961);
or U7088 (N_7088,N_6987,N_6891);
xor U7089 (N_7089,N_6885,N_6986);
and U7090 (N_7090,N_6996,N_6972);
and U7091 (N_7091,N_6990,N_6894);
xor U7092 (N_7092,N_6886,N_6942);
or U7093 (N_7093,N_6940,N_6938);
xor U7094 (N_7094,N_6933,N_6968);
xor U7095 (N_7095,N_6906,N_6961);
or U7096 (N_7096,N_6948,N_6984);
nor U7097 (N_7097,N_6901,N_6919);
and U7098 (N_7098,N_6878,N_6947);
nor U7099 (N_7099,N_6957,N_6990);
xor U7100 (N_7100,N_6883,N_6942);
nor U7101 (N_7101,N_6895,N_6887);
or U7102 (N_7102,N_6922,N_6906);
and U7103 (N_7103,N_6996,N_6877);
nor U7104 (N_7104,N_6912,N_6981);
or U7105 (N_7105,N_6973,N_6884);
or U7106 (N_7106,N_6998,N_6922);
xor U7107 (N_7107,N_6949,N_6957);
nor U7108 (N_7108,N_6892,N_6882);
and U7109 (N_7109,N_6935,N_6986);
nand U7110 (N_7110,N_6997,N_6880);
nor U7111 (N_7111,N_6940,N_6929);
xnor U7112 (N_7112,N_6875,N_6963);
xnor U7113 (N_7113,N_6898,N_6923);
xor U7114 (N_7114,N_6880,N_6885);
nor U7115 (N_7115,N_6998,N_6975);
and U7116 (N_7116,N_6893,N_6891);
xnor U7117 (N_7117,N_6888,N_6997);
nor U7118 (N_7118,N_6893,N_6876);
and U7119 (N_7119,N_6921,N_6903);
nor U7120 (N_7120,N_6923,N_6893);
nor U7121 (N_7121,N_6948,N_6932);
xnor U7122 (N_7122,N_6897,N_6898);
or U7123 (N_7123,N_6920,N_6929);
nand U7124 (N_7124,N_6884,N_6923);
or U7125 (N_7125,N_7070,N_7063);
nand U7126 (N_7126,N_7002,N_7059);
or U7127 (N_7127,N_7055,N_7042);
nor U7128 (N_7128,N_7103,N_7102);
nor U7129 (N_7129,N_7081,N_7096);
xor U7130 (N_7130,N_7075,N_7046);
xnor U7131 (N_7131,N_7114,N_7011);
nand U7132 (N_7132,N_7093,N_7069);
nor U7133 (N_7133,N_7111,N_7026);
xnor U7134 (N_7134,N_7062,N_7020);
nor U7135 (N_7135,N_7057,N_7005);
xnor U7136 (N_7136,N_7048,N_7052);
xor U7137 (N_7137,N_7056,N_7033);
or U7138 (N_7138,N_7071,N_7060);
nand U7139 (N_7139,N_7051,N_7037);
and U7140 (N_7140,N_7123,N_7098);
nor U7141 (N_7141,N_7017,N_7110);
and U7142 (N_7142,N_7064,N_7004);
xor U7143 (N_7143,N_7074,N_7041);
nand U7144 (N_7144,N_7122,N_7032);
xnor U7145 (N_7145,N_7044,N_7007);
or U7146 (N_7146,N_7034,N_7080);
nor U7147 (N_7147,N_7010,N_7043);
and U7148 (N_7148,N_7104,N_7124);
xnor U7149 (N_7149,N_7118,N_7082);
xor U7150 (N_7150,N_7101,N_7066);
xnor U7151 (N_7151,N_7095,N_7106);
and U7152 (N_7152,N_7022,N_7009);
xnor U7153 (N_7153,N_7012,N_7077);
nand U7154 (N_7154,N_7094,N_7087);
or U7155 (N_7155,N_7039,N_7120);
nor U7156 (N_7156,N_7067,N_7105);
and U7157 (N_7157,N_7024,N_7092);
xnor U7158 (N_7158,N_7000,N_7083);
nor U7159 (N_7159,N_7016,N_7072);
or U7160 (N_7160,N_7021,N_7045);
xor U7161 (N_7161,N_7079,N_7030);
or U7162 (N_7162,N_7076,N_7008);
and U7163 (N_7163,N_7078,N_7113);
nand U7164 (N_7164,N_7121,N_7014);
nor U7165 (N_7165,N_7100,N_7003);
xnor U7166 (N_7166,N_7084,N_7031);
and U7167 (N_7167,N_7036,N_7090);
nor U7168 (N_7168,N_7091,N_7047);
nand U7169 (N_7169,N_7023,N_7025);
nor U7170 (N_7170,N_7116,N_7109);
or U7171 (N_7171,N_7053,N_7038);
xnor U7172 (N_7172,N_7097,N_7040);
nor U7173 (N_7173,N_7029,N_7088);
nor U7174 (N_7174,N_7107,N_7006);
and U7175 (N_7175,N_7001,N_7089);
and U7176 (N_7176,N_7085,N_7018);
nand U7177 (N_7177,N_7035,N_7049);
nor U7178 (N_7178,N_7068,N_7115);
nor U7179 (N_7179,N_7015,N_7108);
xnor U7180 (N_7180,N_7073,N_7061);
or U7181 (N_7181,N_7065,N_7058);
xnor U7182 (N_7182,N_7112,N_7119);
nand U7183 (N_7183,N_7099,N_7027);
and U7184 (N_7184,N_7054,N_7013);
and U7185 (N_7185,N_7050,N_7117);
and U7186 (N_7186,N_7028,N_7086);
nor U7187 (N_7187,N_7019,N_7007);
xnor U7188 (N_7188,N_7075,N_7088);
nor U7189 (N_7189,N_7116,N_7000);
nor U7190 (N_7190,N_7090,N_7114);
or U7191 (N_7191,N_7075,N_7077);
nor U7192 (N_7192,N_7058,N_7046);
nor U7193 (N_7193,N_7027,N_7094);
or U7194 (N_7194,N_7058,N_7119);
nor U7195 (N_7195,N_7094,N_7054);
and U7196 (N_7196,N_7099,N_7120);
nor U7197 (N_7197,N_7005,N_7009);
xnor U7198 (N_7198,N_7017,N_7119);
nor U7199 (N_7199,N_7052,N_7060);
nand U7200 (N_7200,N_7056,N_7032);
or U7201 (N_7201,N_7111,N_7004);
nand U7202 (N_7202,N_7111,N_7006);
nor U7203 (N_7203,N_7019,N_7117);
xnor U7204 (N_7204,N_7026,N_7045);
nand U7205 (N_7205,N_7013,N_7055);
nor U7206 (N_7206,N_7017,N_7025);
or U7207 (N_7207,N_7060,N_7120);
nand U7208 (N_7208,N_7072,N_7069);
or U7209 (N_7209,N_7069,N_7021);
nand U7210 (N_7210,N_7072,N_7055);
nand U7211 (N_7211,N_7069,N_7001);
nand U7212 (N_7212,N_7003,N_7101);
or U7213 (N_7213,N_7011,N_7082);
nand U7214 (N_7214,N_7068,N_7004);
xnor U7215 (N_7215,N_7007,N_7014);
nand U7216 (N_7216,N_7026,N_7005);
xnor U7217 (N_7217,N_7033,N_7120);
and U7218 (N_7218,N_7005,N_7067);
nor U7219 (N_7219,N_7065,N_7012);
and U7220 (N_7220,N_7087,N_7080);
or U7221 (N_7221,N_7025,N_7119);
or U7222 (N_7222,N_7082,N_7087);
xor U7223 (N_7223,N_7086,N_7097);
and U7224 (N_7224,N_7104,N_7000);
xor U7225 (N_7225,N_7032,N_7091);
or U7226 (N_7226,N_7115,N_7067);
or U7227 (N_7227,N_7030,N_7010);
nand U7228 (N_7228,N_7004,N_7036);
xnor U7229 (N_7229,N_7018,N_7116);
xnor U7230 (N_7230,N_7051,N_7052);
nand U7231 (N_7231,N_7102,N_7004);
and U7232 (N_7232,N_7114,N_7021);
xor U7233 (N_7233,N_7062,N_7069);
nor U7234 (N_7234,N_7096,N_7071);
nand U7235 (N_7235,N_7009,N_7069);
or U7236 (N_7236,N_7118,N_7043);
and U7237 (N_7237,N_7060,N_7039);
and U7238 (N_7238,N_7089,N_7084);
and U7239 (N_7239,N_7102,N_7041);
nand U7240 (N_7240,N_7030,N_7107);
nor U7241 (N_7241,N_7039,N_7119);
and U7242 (N_7242,N_7055,N_7039);
nand U7243 (N_7243,N_7083,N_7091);
nand U7244 (N_7244,N_7119,N_7084);
nor U7245 (N_7245,N_7012,N_7002);
nand U7246 (N_7246,N_7085,N_7097);
and U7247 (N_7247,N_7039,N_7068);
and U7248 (N_7248,N_7032,N_7106);
or U7249 (N_7249,N_7024,N_7025);
nand U7250 (N_7250,N_7183,N_7237);
xor U7251 (N_7251,N_7128,N_7146);
or U7252 (N_7252,N_7210,N_7209);
xnor U7253 (N_7253,N_7230,N_7196);
nor U7254 (N_7254,N_7136,N_7224);
nor U7255 (N_7255,N_7148,N_7150);
or U7256 (N_7256,N_7154,N_7248);
and U7257 (N_7257,N_7242,N_7149);
and U7258 (N_7258,N_7134,N_7163);
nand U7259 (N_7259,N_7144,N_7233);
nor U7260 (N_7260,N_7153,N_7177);
nor U7261 (N_7261,N_7140,N_7214);
nand U7262 (N_7262,N_7217,N_7221);
nand U7263 (N_7263,N_7231,N_7179);
nor U7264 (N_7264,N_7192,N_7145);
and U7265 (N_7265,N_7182,N_7194);
nand U7266 (N_7266,N_7185,N_7195);
and U7267 (N_7267,N_7173,N_7187);
nor U7268 (N_7268,N_7193,N_7171);
nand U7269 (N_7269,N_7151,N_7125);
or U7270 (N_7270,N_7168,N_7181);
and U7271 (N_7271,N_7226,N_7197);
and U7272 (N_7272,N_7169,N_7131);
nand U7273 (N_7273,N_7244,N_7202);
and U7274 (N_7274,N_7190,N_7238);
or U7275 (N_7275,N_7155,N_7229);
or U7276 (N_7276,N_7212,N_7158);
xnor U7277 (N_7277,N_7141,N_7160);
and U7278 (N_7278,N_7218,N_7137);
nand U7279 (N_7279,N_7204,N_7161);
nand U7280 (N_7280,N_7170,N_7199);
nand U7281 (N_7281,N_7191,N_7235);
or U7282 (N_7282,N_7164,N_7225);
nand U7283 (N_7283,N_7247,N_7147);
and U7284 (N_7284,N_7162,N_7184);
nand U7285 (N_7285,N_7220,N_7156);
and U7286 (N_7286,N_7246,N_7152);
nand U7287 (N_7287,N_7201,N_7206);
nor U7288 (N_7288,N_7186,N_7138);
or U7289 (N_7289,N_7211,N_7166);
nor U7290 (N_7290,N_7216,N_7143);
nor U7291 (N_7291,N_7245,N_7215);
xnor U7292 (N_7292,N_7205,N_7129);
or U7293 (N_7293,N_7198,N_7165);
nor U7294 (N_7294,N_7172,N_7178);
xor U7295 (N_7295,N_7167,N_7227);
and U7296 (N_7296,N_7176,N_7203);
nor U7297 (N_7297,N_7188,N_7126);
nand U7298 (N_7298,N_7200,N_7213);
xor U7299 (N_7299,N_7135,N_7232);
and U7300 (N_7300,N_7222,N_7132);
nand U7301 (N_7301,N_7180,N_7234);
nand U7302 (N_7302,N_7240,N_7174);
or U7303 (N_7303,N_7127,N_7175);
nor U7304 (N_7304,N_7189,N_7249);
xnor U7305 (N_7305,N_7228,N_7219);
nand U7306 (N_7306,N_7236,N_7243);
nand U7307 (N_7307,N_7142,N_7133);
nor U7308 (N_7308,N_7157,N_7159);
or U7309 (N_7309,N_7241,N_7130);
xor U7310 (N_7310,N_7239,N_7208);
or U7311 (N_7311,N_7207,N_7223);
and U7312 (N_7312,N_7139,N_7180);
or U7313 (N_7313,N_7170,N_7158);
or U7314 (N_7314,N_7172,N_7248);
nor U7315 (N_7315,N_7210,N_7241);
or U7316 (N_7316,N_7232,N_7217);
and U7317 (N_7317,N_7238,N_7149);
xnor U7318 (N_7318,N_7138,N_7144);
xnor U7319 (N_7319,N_7189,N_7153);
nand U7320 (N_7320,N_7212,N_7183);
nor U7321 (N_7321,N_7161,N_7248);
xnor U7322 (N_7322,N_7243,N_7221);
nor U7323 (N_7323,N_7134,N_7126);
and U7324 (N_7324,N_7227,N_7230);
and U7325 (N_7325,N_7245,N_7160);
or U7326 (N_7326,N_7248,N_7176);
nor U7327 (N_7327,N_7162,N_7163);
nand U7328 (N_7328,N_7191,N_7205);
nand U7329 (N_7329,N_7214,N_7239);
or U7330 (N_7330,N_7231,N_7142);
nor U7331 (N_7331,N_7227,N_7245);
or U7332 (N_7332,N_7162,N_7190);
nand U7333 (N_7333,N_7141,N_7240);
xor U7334 (N_7334,N_7170,N_7138);
nand U7335 (N_7335,N_7161,N_7211);
xnor U7336 (N_7336,N_7142,N_7195);
or U7337 (N_7337,N_7214,N_7147);
nand U7338 (N_7338,N_7168,N_7215);
xor U7339 (N_7339,N_7131,N_7148);
or U7340 (N_7340,N_7224,N_7232);
or U7341 (N_7341,N_7241,N_7195);
or U7342 (N_7342,N_7142,N_7134);
and U7343 (N_7343,N_7152,N_7142);
and U7344 (N_7344,N_7152,N_7198);
or U7345 (N_7345,N_7203,N_7159);
xor U7346 (N_7346,N_7179,N_7199);
nand U7347 (N_7347,N_7140,N_7243);
xnor U7348 (N_7348,N_7155,N_7208);
nor U7349 (N_7349,N_7181,N_7190);
xor U7350 (N_7350,N_7167,N_7192);
or U7351 (N_7351,N_7145,N_7209);
or U7352 (N_7352,N_7127,N_7226);
xor U7353 (N_7353,N_7158,N_7211);
nor U7354 (N_7354,N_7177,N_7138);
nor U7355 (N_7355,N_7205,N_7208);
and U7356 (N_7356,N_7171,N_7232);
nor U7357 (N_7357,N_7169,N_7141);
xnor U7358 (N_7358,N_7158,N_7242);
nor U7359 (N_7359,N_7192,N_7161);
and U7360 (N_7360,N_7196,N_7187);
nand U7361 (N_7361,N_7177,N_7136);
or U7362 (N_7362,N_7186,N_7183);
xor U7363 (N_7363,N_7142,N_7230);
nand U7364 (N_7364,N_7241,N_7181);
xnor U7365 (N_7365,N_7226,N_7183);
and U7366 (N_7366,N_7127,N_7179);
xnor U7367 (N_7367,N_7133,N_7201);
or U7368 (N_7368,N_7167,N_7139);
xnor U7369 (N_7369,N_7158,N_7230);
xor U7370 (N_7370,N_7181,N_7148);
and U7371 (N_7371,N_7178,N_7188);
and U7372 (N_7372,N_7234,N_7230);
or U7373 (N_7373,N_7245,N_7179);
and U7374 (N_7374,N_7196,N_7244);
xnor U7375 (N_7375,N_7347,N_7287);
nand U7376 (N_7376,N_7307,N_7275);
nor U7377 (N_7377,N_7318,N_7285);
nand U7378 (N_7378,N_7322,N_7283);
or U7379 (N_7379,N_7253,N_7368);
or U7380 (N_7380,N_7272,N_7327);
nor U7381 (N_7381,N_7273,N_7308);
xnor U7382 (N_7382,N_7313,N_7302);
xor U7383 (N_7383,N_7278,N_7331);
nand U7384 (N_7384,N_7303,N_7284);
or U7385 (N_7385,N_7265,N_7361);
nand U7386 (N_7386,N_7342,N_7326);
or U7387 (N_7387,N_7371,N_7356);
nand U7388 (N_7388,N_7362,N_7341);
nand U7389 (N_7389,N_7344,N_7261);
nor U7390 (N_7390,N_7255,N_7333);
nand U7391 (N_7391,N_7291,N_7281);
or U7392 (N_7392,N_7288,N_7369);
nor U7393 (N_7393,N_7359,N_7294);
nor U7394 (N_7394,N_7332,N_7364);
xor U7395 (N_7395,N_7329,N_7252);
and U7396 (N_7396,N_7292,N_7279);
xnor U7397 (N_7397,N_7337,N_7319);
nand U7398 (N_7398,N_7317,N_7309);
and U7399 (N_7399,N_7276,N_7311);
nor U7400 (N_7400,N_7340,N_7277);
nand U7401 (N_7401,N_7367,N_7343);
and U7402 (N_7402,N_7352,N_7260);
xnor U7403 (N_7403,N_7372,N_7325);
xor U7404 (N_7404,N_7274,N_7256);
xor U7405 (N_7405,N_7334,N_7301);
nand U7406 (N_7406,N_7315,N_7296);
nor U7407 (N_7407,N_7324,N_7365);
and U7408 (N_7408,N_7300,N_7355);
and U7409 (N_7409,N_7304,N_7289);
nand U7410 (N_7410,N_7251,N_7346);
xor U7411 (N_7411,N_7266,N_7349);
nand U7412 (N_7412,N_7312,N_7345);
and U7413 (N_7413,N_7267,N_7297);
nand U7414 (N_7414,N_7348,N_7290);
and U7415 (N_7415,N_7366,N_7295);
and U7416 (N_7416,N_7282,N_7286);
or U7417 (N_7417,N_7271,N_7298);
nand U7418 (N_7418,N_7323,N_7269);
or U7419 (N_7419,N_7336,N_7339);
nor U7420 (N_7420,N_7314,N_7280);
xnor U7421 (N_7421,N_7330,N_7363);
nor U7422 (N_7422,N_7257,N_7338);
or U7423 (N_7423,N_7350,N_7374);
and U7424 (N_7424,N_7310,N_7328);
xor U7425 (N_7425,N_7320,N_7268);
nor U7426 (N_7426,N_7258,N_7354);
nand U7427 (N_7427,N_7335,N_7353);
and U7428 (N_7428,N_7254,N_7270);
or U7429 (N_7429,N_7321,N_7250);
and U7430 (N_7430,N_7259,N_7263);
and U7431 (N_7431,N_7351,N_7370);
or U7432 (N_7432,N_7357,N_7306);
nand U7433 (N_7433,N_7293,N_7262);
nand U7434 (N_7434,N_7264,N_7373);
nand U7435 (N_7435,N_7360,N_7358);
and U7436 (N_7436,N_7316,N_7305);
and U7437 (N_7437,N_7299,N_7306);
and U7438 (N_7438,N_7254,N_7281);
nand U7439 (N_7439,N_7253,N_7305);
and U7440 (N_7440,N_7347,N_7300);
or U7441 (N_7441,N_7253,N_7313);
nor U7442 (N_7442,N_7331,N_7265);
and U7443 (N_7443,N_7307,N_7265);
and U7444 (N_7444,N_7281,N_7262);
and U7445 (N_7445,N_7323,N_7260);
or U7446 (N_7446,N_7332,N_7314);
and U7447 (N_7447,N_7346,N_7264);
nor U7448 (N_7448,N_7370,N_7294);
xor U7449 (N_7449,N_7283,N_7257);
nand U7450 (N_7450,N_7254,N_7264);
and U7451 (N_7451,N_7360,N_7303);
nand U7452 (N_7452,N_7306,N_7280);
and U7453 (N_7453,N_7330,N_7365);
xnor U7454 (N_7454,N_7295,N_7278);
or U7455 (N_7455,N_7268,N_7286);
xor U7456 (N_7456,N_7289,N_7335);
or U7457 (N_7457,N_7298,N_7289);
and U7458 (N_7458,N_7349,N_7338);
nand U7459 (N_7459,N_7324,N_7327);
nand U7460 (N_7460,N_7267,N_7362);
and U7461 (N_7461,N_7293,N_7317);
and U7462 (N_7462,N_7361,N_7350);
and U7463 (N_7463,N_7373,N_7293);
and U7464 (N_7464,N_7252,N_7296);
or U7465 (N_7465,N_7254,N_7273);
nor U7466 (N_7466,N_7357,N_7344);
xnor U7467 (N_7467,N_7266,N_7359);
or U7468 (N_7468,N_7264,N_7319);
or U7469 (N_7469,N_7312,N_7306);
nor U7470 (N_7470,N_7276,N_7251);
and U7471 (N_7471,N_7281,N_7294);
and U7472 (N_7472,N_7281,N_7252);
and U7473 (N_7473,N_7324,N_7337);
or U7474 (N_7474,N_7253,N_7258);
nor U7475 (N_7475,N_7326,N_7356);
or U7476 (N_7476,N_7346,N_7331);
nand U7477 (N_7477,N_7360,N_7329);
or U7478 (N_7478,N_7368,N_7372);
nor U7479 (N_7479,N_7344,N_7299);
nand U7480 (N_7480,N_7299,N_7343);
nand U7481 (N_7481,N_7353,N_7373);
nand U7482 (N_7482,N_7368,N_7316);
and U7483 (N_7483,N_7269,N_7331);
xor U7484 (N_7484,N_7334,N_7306);
or U7485 (N_7485,N_7276,N_7323);
and U7486 (N_7486,N_7261,N_7302);
nand U7487 (N_7487,N_7304,N_7294);
nand U7488 (N_7488,N_7320,N_7318);
nand U7489 (N_7489,N_7325,N_7306);
or U7490 (N_7490,N_7362,N_7278);
or U7491 (N_7491,N_7362,N_7292);
nor U7492 (N_7492,N_7314,N_7329);
and U7493 (N_7493,N_7354,N_7337);
nor U7494 (N_7494,N_7287,N_7353);
xnor U7495 (N_7495,N_7301,N_7260);
nand U7496 (N_7496,N_7293,N_7344);
and U7497 (N_7497,N_7313,N_7372);
nand U7498 (N_7498,N_7326,N_7309);
or U7499 (N_7499,N_7296,N_7353);
nand U7500 (N_7500,N_7383,N_7401);
or U7501 (N_7501,N_7408,N_7412);
or U7502 (N_7502,N_7434,N_7410);
and U7503 (N_7503,N_7440,N_7452);
nor U7504 (N_7504,N_7405,N_7486);
or U7505 (N_7505,N_7473,N_7441);
or U7506 (N_7506,N_7466,N_7482);
nand U7507 (N_7507,N_7445,N_7463);
and U7508 (N_7508,N_7485,N_7406);
and U7509 (N_7509,N_7380,N_7454);
and U7510 (N_7510,N_7492,N_7436);
xnor U7511 (N_7511,N_7424,N_7450);
nand U7512 (N_7512,N_7480,N_7460);
nor U7513 (N_7513,N_7430,N_7470);
nand U7514 (N_7514,N_7438,N_7404);
xor U7515 (N_7515,N_7421,N_7396);
xor U7516 (N_7516,N_7413,N_7475);
and U7517 (N_7517,N_7447,N_7455);
nor U7518 (N_7518,N_7435,N_7467);
and U7519 (N_7519,N_7431,N_7423);
and U7520 (N_7520,N_7493,N_7425);
xor U7521 (N_7521,N_7433,N_7394);
or U7522 (N_7522,N_7474,N_7476);
or U7523 (N_7523,N_7457,N_7489);
nand U7524 (N_7524,N_7465,N_7390);
xnor U7525 (N_7525,N_7449,N_7395);
xor U7526 (N_7526,N_7479,N_7439);
nand U7527 (N_7527,N_7414,N_7488);
and U7528 (N_7528,N_7400,N_7446);
or U7529 (N_7529,N_7464,N_7451);
xnor U7530 (N_7530,N_7416,N_7402);
xor U7531 (N_7531,N_7481,N_7429);
xnor U7532 (N_7532,N_7483,N_7382);
and U7533 (N_7533,N_7477,N_7377);
nand U7534 (N_7534,N_7444,N_7428);
and U7535 (N_7535,N_7391,N_7472);
nor U7536 (N_7536,N_7496,N_7427);
nand U7537 (N_7537,N_7462,N_7426);
nand U7538 (N_7538,N_7392,N_7393);
nor U7539 (N_7539,N_7376,N_7403);
xor U7540 (N_7540,N_7499,N_7422);
or U7541 (N_7541,N_7381,N_7399);
xnor U7542 (N_7542,N_7478,N_7442);
nand U7543 (N_7543,N_7389,N_7469);
or U7544 (N_7544,N_7484,N_7495);
xnor U7545 (N_7545,N_7388,N_7398);
nand U7546 (N_7546,N_7387,N_7384);
nor U7547 (N_7547,N_7471,N_7437);
nand U7548 (N_7548,N_7415,N_7411);
and U7549 (N_7549,N_7458,N_7494);
xnor U7550 (N_7550,N_7453,N_7417);
and U7551 (N_7551,N_7459,N_7487);
xor U7552 (N_7552,N_7490,N_7491);
or U7553 (N_7553,N_7432,N_7461);
nand U7554 (N_7554,N_7378,N_7418);
and U7555 (N_7555,N_7375,N_7385);
nor U7556 (N_7556,N_7497,N_7420);
nor U7557 (N_7557,N_7419,N_7386);
nor U7558 (N_7558,N_7456,N_7498);
and U7559 (N_7559,N_7443,N_7409);
and U7560 (N_7560,N_7379,N_7468);
or U7561 (N_7561,N_7397,N_7448);
and U7562 (N_7562,N_7407,N_7395);
nand U7563 (N_7563,N_7496,N_7380);
or U7564 (N_7564,N_7480,N_7403);
nor U7565 (N_7565,N_7404,N_7496);
and U7566 (N_7566,N_7497,N_7433);
nor U7567 (N_7567,N_7441,N_7406);
nor U7568 (N_7568,N_7447,N_7403);
or U7569 (N_7569,N_7451,N_7448);
and U7570 (N_7570,N_7487,N_7396);
nand U7571 (N_7571,N_7491,N_7409);
nor U7572 (N_7572,N_7452,N_7394);
nor U7573 (N_7573,N_7498,N_7417);
nand U7574 (N_7574,N_7435,N_7488);
xor U7575 (N_7575,N_7446,N_7442);
or U7576 (N_7576,N_7375,N_7464);
xor U7577 (N_7577,N_7483,N_7447);
nor U7578 (N_7578,N_7493,N_7416);
or U7579 (N_7579,N_7496,N_7401);
xor U7580 (N_7580,N_7378,N_7410);
xor U7581 (N_7581,N_7376,N_7400);
and U7582 (N_7582,N_7439,N_7494);
xor U7583 (N_7583,N_7448,N_7494);
nor U7584 (N_7584,N_7481,N_7468);
xnor U7585 (N_7585,N_7431,N_7449);
and U7586 (N_7586,N_7480,N_7379);
xnor U7587 (N_7587,N_7466,N_7434);
xnor U7588 (N_7588,N_7488,N_7439);
nor U7589 (N_7589,N_7416,N_7491);
and U7590 (N_7590,N_7378,N_7476);
nor U7591 (N_7591,N_7449,N_7420);
nand U7592 (N_7592,N_7434,N_7394);
nand U7593 (N_7593,N_7409,N_7407);
or U7594 (N_7594,N_7406,N_7448);
nor U7595 (N_7595,N_7439,N_7471);
nor U7596 (N_7596,N_7436,N_7431);
nand U7597 (N_7597,N_7452,N_7424);
and U7598 (N_7598,N_7422,N_7472);
nor U7599 (N_7599,N_7375,N_7411);
nand U7600 (N_7600,N_7439,N_7400);
and U7601 (N_7601,N_7457,N_7477);
or U7602 (N_7602,N_7486,N_7450);
nand U7603 (N_7603,N_7432,N_7389);
nand U7604 (N_7604,N_7497,N_7438);
or U7605 (N_7605,N_7398,N_7391);
xnor U7606 (N_7606,N_7476,N_7495);
nand U7607 (N_7607,N_7449,N_7384);
and U7608 (N_7608,N_7455,N_7432);
nand U7609 (N_7609,N_7388,N_7484);
nor U7610 (N_7610,N_7468,N_7498);
nand U7611 (N_7611,N_7402,N_7378);
nand U7612 (N_7612,N_7420,N_7405);
and U7613 (N_7613,N_7398,N_7406);
nor U7614 (N_7614,N_7427,N_7392);
nor U7615 (N_7615,N_7449,N_7428);
and U7616 (N_7616,N_7428,N_7395);
or U7617 (N_7617,N_7458,N_7453);
or U7618 (N_7618,N_7386,N_7395);
nand U7619 (N_7619,N_7421,N_7440);
nand U7620 (N_7620,N_7392,N_7390);
nor U7621 (N_7621,N_7375,N_7391);
nor U7622 (N_7622,N_7449,N_7476);
nor U7623 (N_7623,N_7413,N_7422);
nor U7624 (N_7624,N_7386,N_7412);
nand U7625 (N_7625,N_7580,N_7547);
or U7626 (N_7626,N_7502,N_7619);
or U7627 (N_7627,N_7526,N_7579);
nand U7628 (N_7628,N_7601,N_7512);
nand U7629 (N_7629,N_7510,N_7610);
or U7630 (N_7630,N_7527,N_7514);
or U7631 (N_7631,N_7548,N_7571);
and U7632 (N_7632,N_7563,N_7550);
or U7633 (N_7633,N_7613,N_7549);
nand U7634 (N_7634,N_7523,N_7582);
and U7635 (N_7635,N_7518,N_7539);
or U7636 (N_7636,N_7536,N_7504);
nand U7637 (N_7637,N_7577,N_7593);
or U7638 (N_7638,N_7501,N_7615);
nor U7639 (N_7639,N_7534,N_7519);
nand U7640 (N_7640,N_7543,N_7572);
and U7641 (N_7641,N_7612,N_7552);
and U7642 (N_7642,N_7594,N_7511);
or U7643 (N_7643,N_7516,N_7614);
and U7644 (N_7644,N_7569,N_7566);
nand U7645 (N_7645,N_7544,N_7595);
or U7646 (N_7646,N_7589,N_7576);
or U7647 (N_7647,N_7602,N_7624);
or U7648 (N_7648,N_7604,N_7554);
or U7649 (N_7649,N_7508,N_7620);
and U7650 (N_7650,N_7541,N_7591);
or U7651 (N_7651,N_7608,N_7513);
nand U7652 (N_7652,N_7521,N_7555);
nor U7653 (N_7653,N_7588,N_7598);
xnor U7654 (N_7654,N_7609,N_7611);
nor U7655 (N_7655,N_7605,N_7600);
nor U7656 (N_7656,N_7621,N_7533);
and U7657 (N_7657,N_7597,N_7574);
nand U7658 (N_7658,N_7568,N_7520);
xnor U7659 (N_7659,N_7535,N_7622);
and U7660 (N_7660,N_7606,N_7522);
and U7661 (N_7661,N_7596,N_7528);
or U7662 (N_7662,N_7532,N_7603);
or U7663 (N_7663,N_7575,N_7590);
or U7664 (N_7664,N_7560,N_7585);
nand U7665 (N_7665,N_7537,N_7570);
xnor U7666 (N_7666,N_7565,N_7553);
or U7667 (N_7667,N_7506,N_7586);
or U7668 (N_7668,N_7509,N_7542);
xor U7669 (N_7669,N_7573,N_7584);
xnor U7670 (N_7670,N_7581,N_7583);
or U7671 (N_7671,N_7540,N_7618);
nor U7672 (N_7672,N_7525,N_7558);
nand U7673 (N_7673,N_7524,N_7564);
nor U7674 (N_7674,N_7556,N_7503);
and U7675 (N_7675,N_7616,N_7500);
and U7676 (N_7676,N_7505,N_7587);
and U7677 (N_7677,N_7599,N_7529);
xor U7678 (N_7678,N_7561,N_7567);
or U7679 (N_7679,N_7515,N_7592);
nor U7680 (N_7680,N_7551,N_7538);
or U7681 (N_7681,N_7578,N_7545);
or U7682 (N_7682,N_7607,N_7623);
and U7683 (N_7683,N_7517,N_7562);
nor U7684 (N_7684,N_7617,N_7531);
nor U7685 (N_7685,N_7559,N_7546);
and U7686 (N_7686,N_7530,N_7507);
xor U7687 (N_7687,N_7557,N_7563);
nor U7688 (N_7688,N_7550,N_7601);
nor U7689 (N_7689,N_7513,N_7598);
nand U7690 (N_7690,N_7564,N_7584);
nor U7691 (N_7691,N_7557,N_7522);
and U7692 (N_7692,N_7553,N_7563);
and U7693 (N_7693,N_7599,N_7568);
or U7694 (N_7694,N_7551,N_7506);
xor U7695 (N_7695,N_7579,N_7547);
and U7696 (N_7696,N_7529,N_7601);
xnor U7697 (N_7697,N_7589,N_7529);
or U7698 (N_7698,N_7515,N_7529);
nor U7699 (N_7699,N_7550,N_7528);
or U7700 (N_7700,N_7616,N_7520);
xnor U7701 (N_7701,N_7615,N_7543);
xor U7702 (N_7702,N_7602,N_7525);
and U7703 (N_7703,N_7552,N_7589);
or U7704 (N_7704,N_7530,N_7620);
nor U7705 (N_7705,N_7524,N_7622);
or U7706 (N_7706,N_7619,N_7536);
nand U7707 (N_7707,N_7553,N_7509);
nor U7708 (N_7708,N_7539,N_7571);
and U7709 (N_7709,N_7613,N_7536);
nor U7710 (N_7710,N_7547,N_7517);
nor U7711 (N_7711,N_7597,N_7541);
nand U7712 (N_7712,N_7515,N_7561);
nand U7713 (N_7713,N_7596,N_7599);
nor U7714 (N_7714,N_7587,N_7549);
xor U7715 (N_7715,N_7514,N_7562);
nor U7716 (N_7716,N_7502,N_7588);
and U7717 (N_7717,N_7609,N_7503);
and U7718 (N_7718,N_7542,N_7595);
nand U7719 (N_7719,N_7557,N_7532);
xnor U7720 (N_7720,N_7589,N_7508);
or U7721 (N_7721,N_7527,N_7544);
nand U7722 (N_7722,N_7624,N_7547);
or U7723 (N_7723,N_7532,N_7518);
xor U7724 (N_7724,N_7624,N_7512);
and U7725 (N_7725,N_7532,N_7574);
or U7726 (N_7726,N_7551,N_7568);
and U7727 (N_7727,N_7559,N_7556);
and U7728 (N_7728,N_7504,N_7619);
xnor U7729 (N_7729,N_7612,N_7532);
nand U7730 (N_7730,N_7593,N_7584);
nand U7731 (N_7731,N_7561,N_7551);
nand U7732 (N_7732,N_7504,N_7583);
nand U7733 (N_7733,N_7578,N_7604);
nand U7734 (N_7734,N_7507,N_7555);
or U7735 (N_7735,N_7567,N_7605);
nand U7736 (N_7736,N_7568,N_7615);
nor U7737 (N_7737,N_7591,N_7617);
and U7738 (N_7738,N_7577,N_7612);
xor U7739 (N_7739,N_7594,N_7580);
or U7740 (N_7740,N_7617,N_7600);
nand U7741 (N_7741,N_7606,N_7575);
nor U7742 (N_7742,N_7579,N_7602);
xnor U7743 (N_7743,N_7557,N_7545);
xnor U7744 (N_7744,N_7522,N_7500);
and U7745 (N_7745,N_7504,N_7591);
nor U7746 (N_7746,N_7524,N_7540);
nand U7747 (N_7747,N_7580,N_7619);
xor U7748 (N_7748,N_7509,N_7511);
and U7749 (N_7749,N_7567,N_7615);
or U7750 (N_7750,N_7683,N_7681);
nor U7751 (N_7751,N_7665,N_7740);
xnor U7752 (N_7752,N_7706,N_7636);
nor U7753 (N_7753,N_7741,N_7649);
or U7754 (N_7754,N_7635,N_7701);
and U7755 (N_7755,N_7744,N_7644);
xor U7756 (N_7756,N_7721,N_7639);
nor U7757 (N_7757,N_7679,N_7697);
or U7758 (N_7758,N_7708,N_7715);
and U7759 (N_7759,N_7746,N_7733);
nor U7760 (N_7760,N_7749,N_7632);
nand U7761 (N_7761,N_7748,N_7707);
nor U7762 (N_7762,N_7734,N_7653);
xor U7763 (N_7763,N_7634,N_7717);
or U7764 (N_7764,N_7664,N_7705);
or U7765 (N_7765,N_7626,N_7641);
or U7766 (N_7766,N_7669,N_7720);
xnor U7767 (N_7767,N_7725,N_7637);
or U7768 (N_7768,N_7673,N_7731);
xnor U7769 (N_7769,N_7661,N_7689);
and U7770 (N_7770,N_7684,N_7703);
xor U7771 (N_7771,N_7685,N_7668);
nand U7772 (N_7772,N_7732,N_7698);
nor U7773 (N_7773,N_7724,N_7670);
and U7774 (N_7774,N_7682,N_7645);
nand U7775 (N_7775,N_7690,N_7691);
nand U7776 (N_7776,N_7659,N_7709);
nand U7777 (N_7777,N_7692,N_7738);
nor U7778 (N_7778,N_7745,N_7630);
nand U7779 (N_7779,N_7742,N_7657);
nand U7780 (N_7780,N_7662,N_7656);
or U7781 (N_7781,N_7693,N_7648);
xnor U7782 (N_7782,N_7688,N_7743);
nand U7783 (N_7783,N_7696,N_7640);
and U7784 (N_7784,N_7686,N_7722);
nor U7785 (N_7785,N_7633,N_7647);
nand U7786 (N_7786,N_7638,N_7710);
and U7787 (N_7787,N_7674,N_7672);
or U7788 (N_7788,N_7702,N_7727);
and U7789 (N_7789,N_7654,N_7719);
and U7790 (N_7790,N_7643,N_7729);
or U7791 (N_7791,N_7628,N_7675);
nand U7792 (N_7792,N_7642,N_7646);
and U7793 (N_7793,N_7737,N_7739);
xnor U7794 (N_7794,N_7714,N_7678);
nand U7795 (N_7795,N_7629,N_7677);
xor U7796 (N_7796,N_7700,N_7652);
or U7797 (N_7797,N_7663,N_7680);
and U7798 (N_7798,N_7736,N_7667);
or U7799 (N_7799,N_7713,N_7671);
xnor U7800 (N_7800,N_7676,N_7660);
nor U7801 (N_7801,N_7712,N_7627);
and U7802 (N_7802,N_7728,N_7658);
nand U7803 (N_7803,N_7694,N_7726);
or U7804 (N_7804,N_7747,N_7666);
nand U7805 (N_7805,N_7631,N_7723);
or U7806 (N_7806,N_7711,N_7718);
nor U7807 (N_7807,N_7655,N_7704);
and U7808 (N_7808,N_7651,N_7699);
xnor U7809 (N_7809,N_7687,N_7625);
and U7810 (N_7810,N_7650,N_7695);
and U7811 (N_7811,N_7735,N_7716);
or U7812 (N_7812,N_7730,N_7637);
nand U7813 (N_7813,N_7745,N_7639);
nor U7814 (N_7814,N_7642,N_7659);
or U7815 (N_7815,N_7676,N_7658);
or U7816 (N_7816,N_7663,N_7635);
xnor U7817 (N_7817,N_7667,N_7721);
or U7818 (N_7818,N_7681,N_7733);
or U7819 (N_7819,N_7650,N_7657);
or U7820 (N_7820,N_7684,N_7737);
xnor U7821 (N_7821,N_7642,N_7697);
or U7822 (N_7822,N_7680,N_7738);
nand U7823 (N_7823,N_7651,N_7722);
or U7824 (N_7824,N_7663,N_7702);
nand U7825 (N_7825,N_7716,N_7640);
nor U7826 (N_7826,N_7659,N_7648);
and U7827 (N_7827,N_7696,N_7630);
nand U7828 (N_7828,N_7712,N_7731);
and U7829 (N_7829,N_7675,N_7723);
and U7830 (N_7830,N_7640,N_7736);
and U7831 (N_7831,N_7631,N_7683);
nor U7832 (N_7832,N_7739,N_7677);
or U7833 (N_7833,N_7681,N_7649);
and U7834 (N_7834,N_7637,N_7710);
or U7835 (N_7835,N_7711,N_7640);
nand U7836 (N_7836,N_7726,N_7718);
xor U7837 (N_7837,N_7643,N_7692);
nand U7838 (N_7838,N_7722,N_7746);
and U7839 (N_7839,N_7630,N_7702);
xnor U7840 (N_7840,N_7728,N_7695);
nand U7841 (N_7841,N_7720,N_7715);
nand U7842 (N_7842,N_7661,N_7641);
nor U7843 (N_7843,N_7729,N_7703);
nor U7844 (N_7844,N_7688,N_7710);
or U7845 (N_7845,N_7702,N_7734);
nor U7846 (N_7846,N_7686,N_7709);
or U7847 (N_7847,N_7664,N_7655);
nand U7848 (N_7848,N_7678,N_7654);
nand U7849 (N_7849,N_7665,N_7651);
xnor U7850 (N_7850,N_7736,N_7707);
or U7851 (N_7851,N_7730,N_7690);
nand U7852 (N_7852,N_7695,N_7709);
or U7853 (N_7853,N_7707,N_7720);
or U7854 (N_7854,N_7681,N_7687);
nand U7855 (N_7855,N_7630,N_7653);
xnor U7856 (N_7856,N_7680,N_7669);
nand U7857 (N_7857,N_7746,N_7625);
nor U7858 (N_7858,N_7698,N_7746);
or U7859 (N_7859,N_7687,N_7649);
or U7860 (N_7860,N_7670,N_7678);
nor U7861 (N_7861,N_7669,N_7661);
xnor U7862 (N_7862,N_7646,N_7702);
nand U7863 (N_7863,N_7683,N_7739);
and U7864 (N_7864,N_7740,N_7671);
and U7865 (N_7865,N_7741,N_7650);
nor U7866 (N_7866,N_7651,N_7716);
nor U7867 (N_7867,N_7654,N_7639);
and U7868 (N_7868,N_7693,N_7728);
nor U7869 (N_7869,N_7641,N_7629);
xor U7870 (N_7870,N_7642,N_7705);
xor U7871 (N_7871,N_7684,N_7728);
or U7872 (N_7872,N_7727,N_7635);
nand U7873 (N_7873,N_7719,N_7705);
or U7874 (N_7874,N_7749,N_7634);
and U7875 (N_7875,N_7783,N_7820);
nor U7876 (N_7876,N_7757,N_7841);
and U7877 (N_7877,N_7770,N_7815);
nand U7878 (N_7878,N_7779,N_7781);
and U7879 (N_7879,N_7873,N_7805);
or U7880 (N_7880,N_7827,N_7818);
and U7881 (N_7881,N_7800,N_7808);
nor U7882 (N_7882,N_7769,N_7856);
nor U7883 (N_7883,N_7785,N_7858);
and U7884 (N_7884,N_7862,N_7838);
nor U7885 (N_7885,N_7792,N_7868);
or U7886 (N_7886,N_7831,N_7846);
nand U7887 (N_7887,N_7773,N_7834);
and U7888 (N_7888,N_7751,N_7829);
nand U7889 (N_7889,N_7810,N_7848);
nor U7890 (N_7890,N_7752,N_7819);
or U7891 (N_7891,N_7817,N_7850);
nand U7892 (N_7892,N_7797,N_7832);
and U7893 (N_7893,N_7772,N_7855);
and U7894 (N_7894,N_7758,N_7771);
or U7895 (N_7895,N_7830,N_7865);
nand U7896 (N_7896,N_7871,N_7837);
or U7897 (N_7897,N_7768,N_7777);
or U7898 (N_7898,N_7754,N_7816);
or U7899 (N_7899,N_7809,N_7863);
and U7900 (N_7900,N_7753,N_7767);
nor U7901 (N_7901,N_7755,N_7836);
nor U7902 (N_7902,N_7762,N_7766);
xor U7903 (N_7903,N_7852,N_7813);
nand U7904 (N_7904,N_7833,N_7782);
and U7905 (N_7905,N_7806,N_7823);
and U7906 (N_7906,N_7790,N_7821);
and U7907 (N_7907,N_7826,N_7799);
xor U7908 (N_7908,N_7750,N_7843);
or U7909 (N_7909,N_7857,N_7825);
or U7910 (N_7910,N_7794,N_7801);
and U7911 (N_7911,N_7842,N_7788);
xnor U7912 (N_7912,N_7824,N_7844);
or U7913 (N_7913,N_7845,N_7764);
nand U7914 (N_7914,N_7814,N_7787);
nor U7915 (N_7915,N_7803,N_7840);
and U7916 (N_7916,N_7869,N_7775);
nor U7917 (N_7917,N_7849,N_7786);
or U7918 (N_7918,N_7853,N_7864);
nand U7919 (N_7919,N_7859,N_7828);
nor U7920 (N_7920,N_7866,N_7791);
and U7921 (N_7921,N_7761,N_7756);
xnor U7922 (N_7922,N_7760,N_7835);
nand U7923 (N_7923,N_7774,N_7793);
nor U7924 (N_7924,N_7765,N_7763);
nor U7925 (N_7925,N_7870,N_7807);
xor U7926 (N_7926,N_7780,N_7839);
nand U7927 (N_7927,N_7847,N_7796);
xnor U7928 (N_7928,N_7759,N_7778);
nand U7929 (N_7929,N_7798,N_7776);
or U7930 (N_7930,N_7860,N_7851);
and U7931 (N_7931,N_7804,N_7874);
xor U7932 (N_7932,N_7789,N_7802);
nor U7933 (N_7933,N_7854,N_7812);
or U7934 (N_7934,N_7795,N_7822);
or U7935 (N_7935,N_7811,N_7872);
nand U7936 (N_7936,N_7861,N_7867);
nand U7937 (N_7937,N_7784,N_7821);
nand U7938 (N_7938,N_7874,N_7801);
nand U7939 (N_7939,N_7861,N_7801);
and U7940 (N_7940,N_7842,N_7844);
nand U7941 (N_7941,N_7847,N_7822);
or U7942 (N_7942,N_7796,N_7865);
and U7943 (N_7943,N_7818,N_7856);
and U7944 (N_7944,N_7854,N_7794);
xor U7945 (N_7945,N_7765,N_7834);
nor U7946 (N_7946,N_7862,N_7805);
or U7947 (N_7947,N_7832,N_7778);
or U7948 (N_7948,N_7814,N_7776);
nor U7949 (N_7949,N_7789,N_7774);
nand U7950 (N_7950,N_7751,N_7800);
xor U7951 (N_7951,N_7820,N_7827);
or U7952 (N_7952,N_7824,N_7758);
or U7953 (N_7953,N_7800,N_7782);
xnor U7954 (N_7954,N_7834,N_7811);
nand U7955 (N_7955,N_7760,N_7850);
xor U7956 (N_7956,N_7820,N_7781);
xor U7957 (N_7957,N_7751,N_7821);
and U7958 (N_7958,N_7835,N_7861);
or U7959 (N_7959,N_7850,N_7830);
or U7960 (N_7960,N_7830,N_7816);
xor U7961 (N_7961,N_7838,N_7870);
xor U7962 (N_7962,N_7764,N_7781);
nand U7963 (N_7963,N_7855,N_7786);
xor U7964 (N_7964,N_7769,N_7798);
or U7965 (N_7965,N_7859,N_7768);
nor U7966 (N_7966,N_7829,N_7781);
xor U7967 (N_7967,N_7800,N_7869);
or U7968 (N_7968,N_7816,N_7864);
or U7969 (N_7969,N_7817,N_7800);
xor U7970 (N_7970,N_7848,N_7788);
nand U7971 (N_7971,N_7785,N_7777);
nand U7972 (N_7972,N_7863,N_7873);
xnor U7973 (N_7973,N_7826,N_7860);
nand U7974 (N_7974,N_7808,N_7820);
nor U7975 (N_7975,N_7774,N_7838);
or U7976 (N_7976,N_7868,N_7822);
and U7977 (N_7977,N_7800,N_7835);
xor U7978 (N_7978,N_7783,N_7837);
nand U7979 (N_7979,N_7775,N_7789);
nor U7980 (N_7980,N_7843,N_7764);
nor U7981 (N_7981,N_7815,N_7778);
nand U7982 (N_7982,N_7859,N_7820);
nor U7983 (N_7983,N_7839,N_7859);
and U7984 (N_7984,N_7787,N_7791);
nand U7985 (N_7985,N_7839,N_7861);
nand U7986 (N_7986,N_7866,N_7822);
nor U7987 (N_7987,N_7796,N_7784);
or U7988 (N_7988,N_7809,N_7770);
nor U7989 (N_7989,N_7806,N_7757);
or U7990 (N_7990,N_7831,N_7871);
or U7991 (N_7991,N_7865,N_7822);
and U7992 (N_7992,N_7851,N_7801);
nand U7993 (N_7993,N_7874,N_7816);
and U7994 (N_7994,N_7850,N_7791);
and U7995 (N_7995,N_7782,N_7802);
nor U7996 (N_7996,N_7792,N_7874);
or U7997 (N_7997,N_7798,N_7832);
or U7998 (N_7998,N_7842,N_7846);
and U7999 (N_7999,N_7851,N_7799);
and U8000 (N_8000,N_7897,N_7948);
or U8001 (N_8001,N_7901,N_7938);
and U8002 (N_8002,N_7961,N_7962);
and U8003 (N_8003,N_7981,N_7896);
nor U8004 (N_8004,N_7886,N_7893);
and U8005 (N_8005,N_7918,N_7977);
or U8006 (N_8006,N_7944,N_7947);
and U8007 (N_8007,N_7959,N_7941);
and U8008 (N_8008,N_7928,N_7916);
or U8009 (N_8009,N_7914,N_7991);
xor U8010 (N_8010,N_7951,N_7910);
nor U8011 (N_8011,N_7898,N_7952);
nand U8012 (N_8012,N_7880,N_7957);
or U8013 (N_8013,N_7934,N_7882);
nand U8014 (N_8014,N_7956,N_7906);
nor U8015 (N_8015,N_7905,N_7930);
nor U8016 (N_8016,N_7958,N_7993);
and U8017 (N_8017,N_7963,N_7936);
nand U8018 (N_8018,N_7978,N_7877);
or U8019 (N_8019,N_7979,N_7965);
and U8020 (N_8020,N_7982,N_7904);
nand U8021 (N_8021,N_7945,N_7975);
and U8022 (N_8022,N_7922,N_7881);
nor U8023 (N_8023,N_7935,N_7964);
or U8024 (N_8024,N_7968,N_7926);
nand U8025 (N_8025,N_7908,N_7949);
or U8026 (N_8026,N_7996,N_7889);
or U8027 (N_8027,N_7899,N_7876);
nor U8028 (N_8028,N_7997,N_7915);
and U8029 (N_8029,N_7900,N_7920);
nand U8030 (N_8030,N_7967,N_7943);
and U8031 (N_8031,N_7925,N_7984);
xor U8032 (N_8032,N_7890,N_7972);
xor U8033 (N_8033,N_7891,N_7970);
or U8034 (N_8034,N_7911,N_7955);
nor U8035 (N_8035,N_7885,N_7913);
xnor U8036 (N_8036,N_7879,N_7888);
nor U8037 (N_8037,N_7960,N_7929);
xor U8038 (N_8038,N_7995,N_7989);
nand U8039 (N_8039,N_7998,N_7912);
nand U8040 (N_8040,N_7903,N_7969);
or U8041 (N_8041,N_7902,N_7980);
nand U8042 (N_8042,N_7953,N_7924);
xor U8043 (N_8043,N_7990,N_7992);
nand U8044 (N_8044,N_7909,N_7942);
nor U8045 (N_8045,N_7931,N_7907);
and U8046 (N_8046,N_7940,N_7999);
nand U8047 (N_8047,N_7973,N_7974);
xnor U8048 (N_8048,N_7917,N_7976);
nand U8049 (N_8049,N_7932,N_7987);
or U8050 (N_8050,N_7875,N_7950);
nand U8051 (N_8051,N_7919,N_7971);
nand U8052 (N_8052,N_7985,N_7946);
or U8053 (N_8053,N_7986,N_7923);
or U8054 (N_8054,N_7892,N_7983);
xor U8055 (N_8055,N_7927,N_7933);
nand U8056 (N_8056,N_7894,N_7895);
nand U8057 (N_8057,N_7921,N_7939);
or U8058 (N_8058,N_7878,N_7994);
xor U8059 (N_8059,N_7954,N_7887);
and U8060 (N_8060,N_7937,N_7966);
nor U8061 (N_8061,N_7883,N_7884);
or U8062 (N_8062,N_7988,N_7982);
nor U8063 (N_8063,N_7896,N_7911);
and U8064 (N_8064,N_7951,N_7878);
nor U8065 (N_8065,N_7962,N_7901);
and U8066 (N_8066,N_7899,N_7973);
xor U8067 (N_8067,N_7936,N_7923);
and U8068 (N_8068,N_7976,N_7900);
nand U8069 (N_8069,N_7946,N_7990);
xnor U8070 (N_8070,N_7956,N_7939);
nor U8071 (N_8071,N_7991,N_7886);
or U8072 (N_8072,N_7974,N_7950);
or U8073 (N_8073,N_7987,N_7881);
and U8074 (N_8074,N_7946,N_7923);
xnor U8075 (N_8075,N_7994,N_7896);
and U8076 (N_8076,N_7933,N_7882);
or U8077 (N_8077,N_7894,N_7936);
or U8078 (N_8078,N_7938,N_7890);
or U8079 (N_8079,N_7889,N_7921);
nand U8080 (N_8080,N_7918,N_7972);
xor U8081 (N_8081,N_7954,N_7933);
xnor U8082 (N_8082,N_7997,N_7982);
or U8083 (N_8083,N_7989,N_7974);
xnor U8084 (N_8084,N_7930,N_7900);
or U8085 (N_8085,N_7888,N_7976);
nand U8086 (N_8086,N_7952,N_7938);
nand U8087 (N_8087,N_7984,N_7917);
xor U8088 (N_8088,N_7984,N_7914);
or U8089 (N_8089,N_7936,N_7943);
nor U8090 (N_8090,N_7920,N_7990);
nand U8091 (N_8091,N_7987,N_7904);
or U8092 (N_8092,N_7956,N_7951);
xor U8093 (N_8093,N_7983,N_7888);
nor U8094 (N_8094,N_7937,N_7942);
nor U8095 (N_8095,N_7980,N_7952);
and U8096 (N_8096,N_7955,N_7918);
xnor U8097 (N_8097,N_7976,N_7912);
nor U8098 (N_8098,N_7916,N_7924);
nand U8099 (N_8099,N_7905,N_7899);
xnor U8100 (N_8100,N_7955,N_7995);
xor U8101 (N_8101,N_7940,N_7944);
or U8102 (N_8102,N_7970,N_7907);
nand U8103 (N_8103,N_7975,N_7950);
or U8104 (N_8104,N_7904,N_7877);
nor U8105 (N_8105,N_7922,N_7890);
nand U8106 (N_8106,N_7909,N_7920);
nor U8107 (N_8107,N_7924,N_7966);
nand U8108 (N_8108,N_7875,N_7948);
and U8109 (N_8109,N_7993,N_7939);
or U8110 (N_8110,N_7970,N_7964);
nand U8111 (N_8111,N_7951,N_7965);
nor U8112 (N_8112,N_7913,N_7956);
nor U8113 (N_8113,N_7963,N_7950);
or U8114 (N_8114,N_7937,N_7913);
nand U8115 (N_8115,N_7931,N_7893);
or U8116 (N_8116,N_7896,N_7954);
nand U8117 (N_8117,N_7916,N_7879);
xnor U8118 (N_8118,N_7879,N_7983);
nand U8119 (N_8119,N_7899,N_7981);
or U8120 (N_8120,N_7987,N_7954);
xor U8121 (N_8121,N_7952,N_7897);
nand U8122 (N_8122,N_7952,N_7927);
nand U8123 (N_8123,N_7926,N_7974);
nor U8124 (N_8124,N_7947,N_7996);
nand U8125 (N_8125,N_8020,N_8043);
nand U8126 (N_8126,N_8116,N_8015);
or U8127 (N_8127,N_8117,N_8056);
and U8128 (N_8128,N_8014,N_8098);
xnor U8129 (N_8129,N_8067,N_8088);
xnor U8130 (N_8130,N_8105,N_8031);
xnor U8131 (N_8131,N_8061,N_8107);
or U8132 (N_8132,N_8090,N_8121);
and U8133 (N_8133,N_8097,N_8096);
and U8134 (N_8134,N_8082,N_8085);
or U8135 (N_8135,N_8072,N_8080);
nor U8136 (N_8136,N_8075,N_8028);
and U8137 (N_8137,N_8039,N_8035);
and U8138 (N_8138,N_8106,N_8062);
xnor U8139 (N_8139,N_8027,N_8063);
or U8140 (N_8140,N_8110,N_8000);
xnor U8141 (N_8141,N_8047,N_8005);
nor U8142 (N_8142,N_8040,N_8114);
nor U8143 (N_8143,N_8089,N_8004);
nand U8144 (N_8144,N_8123,N_8030);
xor U8145 (N_8145,N_8095,N_8001);
and U8146 (N_8146,N_8073,N_8059);
or U8147 (N_8147,N_8050,N_8071);
nand U8148 (N_8148,N_8037,N_8083);
or U8149 (N_8149,N_8011,N_8058);
or U8150 (N_8150,N_8112,N_8124);
or U8151 (N_8151,N_8021,N_8016);
and U8152 (N_8152,N_8079,N_8091);
nand U8153 (N_8153,N_8102,N_8086);
nor U8154 (N_8154,N_8038,N_8053);
nand U8155 (N_8155,N_8013,N_8007);
nor U8156 (N_8156,N_8034,N_8094);
nand U8157 (N_8157,N_8100,N_8066);
xnor U8158 (N_8158,N_8024,N_8010);
nor U8159 (N_8159,N_8002,N_8101);
nor U8160 (N_8160,N_8006,N_8041);
xnor U8161 (N_8161,N_8008,N_8051);
nor U8162 (N_8162,N_8057,N_8019);
xor U8163 (N_8163,N_8064,N_8084);
and U8164 (N_8164,N_8070,N_8122);
xnor U8165 (N_8165,N_8099,N_8054);
or U8166 (N_8166,N_8046,N_8009);
or U8167 (N_8167,N_8092,N_8081);
or U8168 (N_8168,N_8049,N_8033);
or U8169 (N_8169,N_8042,N_8025);
or U8170 (N_8170,N_8078,N_8104);
nand U8171 (N_8171,N_8044,N_8113);
and U8172 (N_8172,N_8048,N_8029);
and U8173 (N_8173,N_8108,N_8118);
and U8174 (N_8174,N_8077,N_8120);
nand U8175 (N_8175,N_8018,N_8103);
nor U8176 (N_8176,N_8060,N_8003);
or U8177 (N_8177,N_8119,N_8074);
xnor U8178 (N_8178,N_8109,N_8065);
or U8179 (N_8179,N_8069,N_8026);
xnor U8180 (N_8180,N_8076,N_8055);
and U8181 (N_8181,N_8022,N_8017);
nand U8182 (N_8182,N_8087,N_8045);
xnor U8183 (N_8183,N_8036,N_8052);
or U8184 (N_8184,N_8032,N_8068);
nand U8185 (N_8185,N_8093,N_8111);
nand U8186 (N_8186,N_8115,N_8012);
nor U8187 (N_8187,N_8023,N_8000);
nor U8188 (N_8188,N_8019,N_8047);
nor U8189 (N_8189,N_8063,N_8086);
nand U8190 (N_8190,N_8119,N_8077);
or U8191 (N_8191,N_8105,N_8015);
or U8192 (N_8192,N_8020,N_8105);
or U8193 (N_8193,N_8001,N_8076);
nand U8194 (N_8194,N_8034,N_8023);
nor U8195 (N_8195,N_8071,N_8002);
and U8196 (N_8196,N_8003,N_8063);
nor U8197 (N_8197,N_8088,N_8059);
or U8198 (N_8198,N_8036,N_8060);
nand U8199 (N_8199,N_8066,N_8118);
nor U8200 (N_8200,N_8065,N_8022);
nor U8201 (N_8201,N_8115,N_8001);
and U8202 (N_8202,N_8019,N_8063);
or U8203 (N_8203,N_8000,N_8064);
nand U8204 (N_8204,N_8117,N_8058);
nand U8205 (N_8205,N_8095,N_8078);
nand U8206 (N_8206,N_8112,N_8025);
nor U8207 (N_8207,N_8087,N_8071);
and U8208 (N_8208,N_8119,N_8105);
and U8209 (N_8209,N_8080,N_8034);
or U8210 (N_8210,N_8114,N_8094);
nand U8211 (N_8211,N_8093,N_8016);
xnor U8212 (N_8212,N_8043,N_8012);
xnor U8213 (N_8213,N_8053,N_8122);
nand U8214 (N_8214,N_8075,N_8100);
or U8215 (N_8215,N_8079,N_8107);
nand U8216 (N_8216,N_8033,N_8058);
or U8217 (N_8217,N_8014,N_8104);
or U8218 (N_8218,N_8080,N_8098);
or U8219 (N_8219,N_8037,N_8095);
xor U8220 (N_8220,N_8057,N_8028);
and U8221 (N_8221,N_8089,N_8074);
xor U8222 (N_8222,N_8085,N_8099);
xnor U8223 (N_8223,N_8020,N_8051);
xor U8224 (N_8224,N_8001,N_8048);
and U8225 (N_8225,N_8063,N_8022);
and U8226 (N_8226,N_8107,N_8094);
nand U8227 (N_8227,N_8040,N_8121);
and U8228 (N_8228,N_8063,N_8112);
or U8229 (N_8229,N_8055,N_8011);
and U8230 (N_8230,N_8043,N_8057);
or U8231 (N_8231,N_8025,N_8066);
nand U8232 (N_8232,N_8124,N_8120);
xor U8233 (N_8233,N_8078,N_8023);
xor U8234 (N_8234,N_8073,N_8003);
nor U8235 (N_8235,N_8103,N_8067);
or U8236 (N_8236,N_8101,N_8016);
nor U8237 (N_8237,N_8123,N_8042);
xor U8238 (N_8238,N_8088,N_8073);
or U8239 (N_8239,N_8087,N_8088);
or U8240 (N_8240,N_8058,N_8021);
nand U8241 (N_8241,N_8010,N_8050);
and U8242 (N_8242,N_8096,N_8067);
and U8243 (N_8243,N_8061,N_8070);
xnor U8244 (N_8244,N_8119,N_8063);
or U8245 (N_8245,N_8097,N_8064);
xnor U8246 (N_8246,N_8012,N_8114);
xor U8247 (N_8247,N_8042,N_8106);
and U8248 (N_8248,N_8033,N_8113);
nand U8249 (N_8249,N_8123,N_8073);
xor U8250 (N_8250,N_8132,N_8240);
nor U8251 (N_8251,N_8236,N_8208);
and U8252 (N_8252,N_8195,N_8223);
xnor U8253 (N_8253,N_8235,N_8207);
xnor U8254 (N_8254,N_8148,N_8174);
nand U8255 (N_8255,N_8149,N_8230);
nor U8256 (N_8256,N_8152,N_8245);
and U8257 (N_8257,N_8151,N_8238);
nor U8258 (N_8258,N_8204,N_8177);
and U8259 (N_8259,N_8170,N_8164);
nand U8260 (N_8260,N_8167,N_8214);
or U8261 (N_8261,N_8218,N_8157);
and U8262 (N_8262,N_8165,N_8139);
and U8263 (N_8263,N_8231,N_8183);
and U8264 (N_8264,N_8196,N_8187);
nor U8265 (N_8265,N_8166,N_8127);
and U8266 (N_8266,N_8125,N_8192);
nand U8267 (N_8267,N_8241,N_8138);
or U8268 (N_8268,N_8205,N_8202);
nand U8269 (N_8269,N_8175,N_8225);
nor U8270 (N_8270,N_8147,N_8140);
xnor U8271 (N_8271,N_8133,N_8201);
and U8272 (N_8272,N_8190,N_8173);
and U8273 (N_8273,N_8243,N_8155);
xnor U8274 (N_8274,N_8134,N_8163);
and U8275 (N_8275,N_8178,N_8217);
nand U8276 (N_8276,N_8179,N_8181);
nor U8277 (N_8277,N_8249,N_8129);
or U8278 (N_8278,N_8219,N_8213);
nor U8279 (N_8279,N_8221,N_8211);
and U8280 (N_8280,N_8189,N_8161);
nor U8281 (N_8281,N_8180,N_8212);
xnor U8282 (N_8282,N_8169,N_8171);
or U8283 (N_8283,N_8153,N_8244);
nor U8284 (N_8284,N_8156,N_8186);
nand U8285 (N_8285,N_8232,N_8198);
nand U8286 (N_8286,N_8228,N_8220);
or U8287 (N_8287,N_8160,N_8247);
xnor U8288 (N_8288,N_8209,N_8199);
nand U8289 (N_8289,N_8203,N_8242);
xor U8290 (N_8290,N_8158,N_8206);
or U8291 (N_8291,N_8136,N_8210);
nand U8292 (N_8292,N_8191,N_8131);
or U8293 (N_8293,N_8248,N_8246);
nand U8294 (N_8294,N_8188,N_8197);
nor U8295 (N_8295,N_8145,N_8239);
nand U8296 (N_8296,N_8185,N_8154);
and U8297 (N_8297,N_8168,N_8234);
xor U8298 (N_8298,N_8222,N_8229);
and U8299 (N_8299,N_8130,N_8200);
nand U8300 (N_8300,N_8159,N_8128);
nand U8301 (N_8301,N_8216,N_8237);
nand U8302 (N_8302,N_8162,N_8150);
and U8303 (N_8303,N_8142,N_8224);
or U8304 (N_8304,N_8226,N_8176);
and U8305 (N_8305,N_8184,N_8233);
nand U8306 (N_8306,N_8227,N_8146);
or U8307 (N_8307,N_8182,N_8144);
and U8308 (N_8308,N_8193,N_8172);
and U8309 (N_8309,N_8215,N_8135);
or U8310 (N_8310,N_8141,N_8137);
nor U8311 (N_8311,N_8194,N_8143);
and U8312 (N_8312,N_8126,N_8143);
xnor U8313 (N_8313,N_8199,N_8136);
nor U8314 (N_8314,N_8133,N_8180);
xor U8315 (N_8315,N_8199,N_8187);
and U8316 (N_8316,N_8213,N_8207);
xor U8317 (N_8317,N_8140,N_8214);
and U8318 (N_8318,N_8171,N_8196);
nor U8319 (N_8319,N_8162,N_8215);
or U8320 (N_8320,N_8195,N_8245);
xnor U8321 (N_8321,N_8190,N_8242);
nand U8322 (N_8322,N_8161,N_8228);
xnor U8323 (N_8323,N_8180,N_8231);
nor U8324 (N_8324,N_8185,N_8125);
xnor U8325 (N_8325,N_8154,N_8181);
or U8326 (N_8326,N_8230,N_8160);
nand U8327 (N_8327,N_8150,N_8227);
and U8328 (N_8328,N_8131,N_8188);
or U8329 (N_8329,N_8218,N_8217);
nand U8330 (N_8330,N_8148,N_8236);
nand U8331 (N_8331,N_8216,N_8167);
or U8332 (N_8332,N_8229,N_8131);
nand U8333 (N_8333,N_8141,N_8155);
xnor U8334 (N_8334,N_8235,N_8198);
nand U8335 (N_8335,N_8209,N_8212);
and U8336 (N_8336,N_8214,N_8239);
or U8337 (N_8337,N_8206,N_8208);
or U8338 (N_8338,N_8148,N_8206);
nand U8339 (N_8339,N_8163,N_8246);
and U8340 (N_8340,N_8155,N_8143);
or U8341 (N_8341,N_8175,N_8244);
xor U8342 (N_8342,N_8209,N_8204);
nor U8343 (N_8343,N_8182,N_8176);
nor U8344 (N_8344,N_8228,N_8137);
and U8345 (N_8345,N_8211,N_8151);
xnor U8346 (N_8346,N_8160,N_8224);
and U8347 (N_8347,N_8212,N_8159);
xor U8348 (N_8348,N_8144,N_8215);
or U8349 (N_8349,N_8157,N_8247);
or U8350 (N_8350,N_8136,N_8245);
and U8351 (N_8351,N_8241,N_8202);
or U8352 (N_8352,N_8138,N_8202);
xor U8353 (N_8353,N_8195,N_8247);
nand U8354 (N_8354,N_8143,N_8133);
nand U8355 (N_8355,N_8175,N_8136);
nand U8356 (N_8356,N_8150,N_8167);
and U8357 (N_8357,N_8222,N_8166);
or U8358 (N_8358,N_8152,N_8239);
nand U8359 (N_8359,N_8169,N_8217);
nand U8360 (N_8360,N_8243,N_8163);
or U8361 (N_8361,N_8156,N_8160);
nor U8362 (N_8362,N_8227,N_8136);
nor U8363 (N_8363,N_8127,N_8128);
and U8364 (N_8364,N_8171,N_8133);
nand U8365 (N_8365,N_8128,N_8186);
and U8366 (N_8366,N_8240,N_8170);
nor U8367 (N_8367,N_8141,N_8170);
xor U8368 (N_8368,N_8236,N_8186);
nor U8369 (N_8369,N_8159,N_8239);
and U8370 (N_8370,N_8217,N_8162);
nor U8371 (N_8371,N_8153,N_8133);
nand U8372 (N_8372,N_8146,N_8172);
nand U8373 (N_8373,N_8158,N_8164);
or U8374 (N_8374,N_8198,N_8177);
or U8375 (N_8375,N_8286,N_8304);
nand U8376 (N_8376,N_8258,N_8292);
nand U8377 (N_8377,N_8264,N_8297);
nand U8378 (N_8378,N_8300,N_8333);
and U8379 (N_8379,N_8347,N_8335);
nand U8380 (N_8380,N_8260,N_8352);
and U8381 (N_8381,N_8315,N_8322);
xor U8382 (N_8382,N_8362,N_8349);
xnor U8383 (N_8383,N_8350,N_8290);
and U8384 (N_8384,N_8281,N_8351);
nor U8385 (N_8385,N_8283,N_8318);
and U8386 (N_8386,N_8293,N_8294);
nand U8387 (N_8387,N_8269,N_8275);
and U8388 (N_8388,N_8251,N_8346);
or U8389 (N_8389,N_8274,N_8278);
or U8390 (N_8390,N_8366,N_8262);
nor U8391 (N_8391,N_8344,N_8372);
nand U8392 (N_8392,N_8280,N_8267);
nor U8393 (N_8393,N_8287,N_8268);
or U8394 (N_8394,N_8250,N_8310);
nor U8395 (N_8395,N_8325,N_8299);
nor U8396 (N_8396,N_8259,N_8265);
xor U8397 (N_8397,N_8309,N_8308);
or U8398 (N_8398,N_8374,N_8354);
xor U8399 (N_8399,N_8261,N_8343);
and U8400 (N_8400,N_8279,N_8364);
xor U8401 (N_8401,N_8340,N_8370);
xor U8402 (N_8402,N_8306,N_8311);
xnor U8403 (N_8403,N_8302,N_8342);
xor U8404 (N_8404,N_8336,N_8252);
nor U8405 (N_8405,N_8338,N_8288);
and U8406 (N_8406,N_8345,N_8359);
and U8407 (N_8407,N_8341,N_8326);
nor U8408 (N_8408,N_8356,N_8313);
nor U8409 (N_8409,N_8276,N_8266);
xor U8410 (N_8410,N_8348,N_8360);
nand U8411 (N_8411,N_8337,N_8289);
nor U8412 (N_8412,N_8256,N_8319);
xor U8413 (N_8413,N_8368,N_8331);
xnor U8414 (N_8414,N_8291,N_8303);
and U8415 (N_8415,N_8263,N_8301);
nor U8416 (N_8416,N_8357,N_8353);
or U8417 (N_8417,N_8312,N_8255);
and U8418 (N_8418,N_8323,N_8254);
nand U8419 (N_8419,N_8332,N_8334);
or U8420 (N_8420,N_8282,N_8314);
nand U8421 (N_8421,N_8329,N_8373);
nand U8422 (N_8422,N_8363,N_8272);
xnor U8423 (N_8423,N_8298,N_8327);
nand U8424 (N_8424,N_8321,N_8369);
nor U8425 (N_8425,N_8367,N_8253);
nand U8426 (N_8426,N_8358,N_8271);
xor U8427 (N_8427,N_8330,N_8295);
xnor U8428 (N_8428,N_8317,N_8361);
nand U8429 (N_8429,N_8371,N_8328);
xnor U8430 (N_8430,N_8257,N_8324);
or U8431 (N_8431,N_8316,N_8355);
xnor U8432 (N_8432,N_8284,N_8365);
xnor U8433 (N_8433,N_8307,N_8296);
or U8434 (N_8434,N_8285,N_8339);
nand U8435 (N_8435,N_8320,N_8305);
nor U8436 (N_8436,N_8270,N_8277);
nor U8437 (N_8437,N_8273,N_8289);
xor U8438 (N_8438,N_8348,N_8303);
and U8439 (N_8439,N_8294,N_8296);
nor U8440 (N_8440,N_8272,N_8356);
nand U8441 (N_8441,N_8323,N_8337);
nor U8442 (N_8442,N_8342,N_8281);
nand U8443 (N_8443,N_8278,N_8363);
xor U8444 (N_8444,N_8307,N_8287);
xor U8445 (N_8445,N_8346,N_8317);
nor U8446 (N_8446,N_8279,N_8272);
nor U8447 (N_8447,N_8298,N_8350);
nor U8448 (N_8448,N_8250,N_8341);
or U8449 (N_8449,N_8250,N_8350);
and U8450 (N_8450,N_8276,N_8258);
nand U8451 (N_8451,N_8334,N_8290);
and U8452 (N_8452,N_8260,N_8342);
xnor U8453 (N_8453,N_8353,N_8316);
and U8454 (N_8454,N_8282,N_8258);
nor U8455 (N_8455,N_8307,N_8323);
nor U8456 (N_8456,N_8281,N_8330);
and U8457 (N_8457,N_8293,N_8276);
nor U8458 (N_8458,N_8372,N_8357);
nand U8459 (N_8459,N_8324,N_8352);
or U8460 (N_8460,N_8358,N_8333);
xor U8461 (N_8461,N_8321,N_8307);
nand U8462 (N_8462,N_8270,N_8361);
or U8463 (N_8463,N_8255,N_8352);
nand U8464 (N_8464,N_8324,N_8293);
nor U8465 (N_8465,N_8358,N_8354);
xor U8466 (N_8466,N_8372,N_8280);
nor U8467 (N_8467,N_8312,N_8371);
or U8468 (N_8468,N_8283,N_8314);
or U8469 (N_8469,N_8312,N_8273);
or U8470 (N_8470,N_8347,N_8317);
or U8471 (N_8471,N_8326,N_8269);
nor U8472 (N_8472,N_8296,N_8313);
xor U8473 (N_8473,N_8296,N_8300);
xnor U8474 (N_8474,N_8269,N_8251);
xor U8475 (N_8475,N_8253,N_8271);
or U8476 (N_8476,N_8256,N_8325);
nand U8477 (N_8477,N_8330,N_8364);
nor U8478 (N_8478,N_8368,N_8304);
or U8479 (N_8479,N_8303,N_8329);
and U8480 (N_8480,N_8283,N_8326);
or U8481 (N_8481,N_8367,N_8261);
or U8482 (N_8482,N_8366,N_8356);
nor U8483 (N_8483,N_8366,N_8263);
or U8484 (N_8484,N_8344,N_8328);
nand U8485 (N_8485,N_8369,N_8367);
nor U8486 (N_8486,N_8276,N_8321);
and U8487 (N_8487,N_8322,N_8360);
and U8488 (N_8488,N_8319,N_8265);
nor U8489 (N_8489,N_8337,N_8314);
or U8490 (N_8490,N_8321,N_8338);
or U8491 (N_8491,N_8341,N_8265);
nor U8492 (N_8492,N_8279,N_8275);
xnor U8493 (N_8493,N_8374,N_8280);
nand U8494 (N_8494,N_8328,N_8299);
nor U8495 (N_8495,N_8370,N_8312);
and U8496 (N_8496,N_8267,N_8283);
xnor U8497 (N_8497,N_8252,N_8330);
nand U8498 (N_8498,N_8257,N_8353);
or U8499 (N_8499,N_8277,N_8321);
xor U8500 (N_8500,N_8414,N_8408);
nor U8501 (N_8501,N_8426,N_8385);
or U8502 (N_8502,N_8379,N_8390);
and U8503 (N_8503,N_8480,N_8423);
and U8504 (N_8504,N_8416,N_8384);
nand U8505 (N_8505,N_8495,N_8466);
and U8506 (N_8506,N_8393,N_8420);
xor U8507 (N_8507,N_8473,N_8491);
nand U8508 (N_8508,N_8386,N_8482);
or U8509 (N_8509,N_8484,N_8411);
and U8510 (N_8510,N_8391,N_8492);
nor U8511 (N_8511,N_8382,N_8424);
nor U8512 (N_8512,N_8446,N_8410);
xnor U8513 (N_8513,N_8433,N_8375);
nand U8514 (N_8514,N_8459,N_8440);
and U8515 (N_8515,N_8475,N_8432);
and U8516 (N_8516,N_8464,N_8401);
or U8517 (N_8517,N_8447,N_8377);
nor U8518 (N_8518,N_8395,N_8450);
xnor U8519 (N_8519,N_8387,N_8438);
nor U8520 (N_8520,N_8430,N_8409);
and U8521 (N_8521,N_8389,N_8462);
or U8522 (N_8522,N_8429,N_8476);
or U8523 (N_8523,N_8439,N_8442);
xor U8524 (N_8524,N_8403,N_8376);
and U8525 (N_8525,N_8481,N_8471);
nor U8526 (N_8526,N_8406,N_8456);
or U8527 (N_8527,N_8415,N_8469);
xnor U8528 (N_8528,N_8496,N_8457);
nor U8529 (N_8529,N_8499,N_8397);
nand U8530 (N_8530,N_8418,N_8402);
xnor U8531 (N_8531,N_8497,N_8434);
or U8532 (N_8532,N_8460,N_8488);
nand U8533 (N_8533,N_8441,N_8392);
and U8534 (N_8534,N_8463,N_8483);
nor U8535 (N_8535,N_8428,N_8461);
and U8536 (N_8536,N_8479,N_8436);
nand U8537 (N_8537,N_8468,N_8467);
nor U8538 (N_8538,N_8425,N_8485);
nor U8539 (N_8539,N_8443,N_8431);
or U8540 (N_8540,N_8421,N_8380);
and U8541 (N_8541,N_8486,N_8396);
nand U8542 (N_8542,N_8452,N_8444);
nor U8543 (N_8543,N_8477,N_8413);
and U8544 (N_8544,N_8470,N_8381);
or U8545 (N_8545,N_8445,N_8422);
nor U8546 (N_8546,N_8494,N_8388);
nand U8547 (N_8547,N_8465,N_8399);
xnor U8548 (N_8548,N_8417,N_8474);
and U8549 (N_8549,N_8435,N_8448);
xnor U8550 (N_8550,N_8394,N_8490);
nor U8551 (N_8551,N_8412,N_8419);
and U8552 (N_8552,N_8454,N_8449);
nor U8553 (N_8553,N_8455,N_8498);
xor U8554 (N_8554,N_8400,N_8487);
or U8555 (N_8555,N_8478,N_8453);
or U8556 (N_8556,N_8383,N_8398);
nand U8557 (N_8557,N_8493,N_8405);
nor U8558 (N_8558,N_8427,N_8472);
nor U8559 (N_8559,N_8407,N_8458);
and U8560 (N_8560,N_8451,N_8378);
xor U8561 (N_8561,N_8489,N_8404);
nor U8562 (N_8562,N_8437,N_8385);
xor U8563 (N_8563,N_8454,N_8453);
xor U8564 (N_8564,N_8392,N_8488);
nand U8565 (N_8565,N_8429,N_8484);
nand U8566 (N_8566,N_8490,N_8398);
xnor U8567 (N_8567,N_8438,N_8420);
or U8568 (N_8568,N_8387,N_8435);
or U8569 (N_8569,N_8376,N_8388);
or U8570 (N_8570,N_8481,N_8408);
and U8571 (N_8571,N_8422,N_8382);
xor U8572 (N_8572,N_8385,N_8442);
and U8573 (N_8573,N_8485,N_8489);
or U8574 (N_8574,N_8421,N_8401);
nand U8575 (N_8575,N_8454,N_8425);
nand U8576 (N_8576,N_8420,N_8400);
or U8577 (N_8577,N_8499,N_8489);
nor U8578 (N_8578,N_8480,N_8395);
and U8579 (N_8579,N_8491,N_8388);
and U8580 (N_8580,N_8476,N_8416);
and U8581 (N_8581,N_8389,N_8454);
nand U8582 (N_8582,N_8424,N_8391);
or U8583 (N_8583,N_8380,N_8463);
xnor U8584 (N_8584,N_8377,N_8396);
and U8585 (N_8585,N_8377,N_8440);
and U8586 (N_8586,N_8495,N_8429);
nand U8587 (N_8587,N_8449,N_8433);
and U8588 (N_8588,N_8492,N_8438);
and U8589 (N_8589,N_8467,N_8420);
and U8590 (N_8590,N_8443,N_8388);
nand U8591 (N_8591,N_8422,N_8402);
or U8592 (N_8592,N_8406,N_8457);
or U8593 (N_8593,N_8382,N_8460);
and U8594 (N_8594,N_8430,N_8493);
nand U8595 (N_8595,N_8432,N_8495);
or U8596 (N_8596,N_8436,N_8380);
and U8597 (N_8597,N_8486,N_8394);
xnor U8598 (N_8598,N_8454,N_8474);
nor U8599 (N_8599,N_8422,N_8400);
or U8600 (N_8600,N_8485,N_8381);
or U8601 (N_8601,N_8413,N_8492);
xnor U8602 (N_8602,N_8479,N_8426);
nor U8603 (N_8603,N_8380,N_8466);
or U8604 (N_8604,N_8463,N_8473);
nor U8605 (N_8605,N_8475,N_8454);
nand U8606 (N_8606,N_8420,N_8402);
nand U8607 (N_8607,N_8400,N_8477);
xor U8608 (N_8608,N_8416,N_8402);
nor U8609 (N_8609,N_8469,N_8404);
nor U8610 (N_8610,N_8438,N_8418);
xnor U8611 (N_8611,N_8484,N_8432);
and U8612 (N_8612,N_8457,N_8415);
nor U8613 (N_8613,N_8406,N_8422);
or U8614 (N_8614,N_8421,N_8499);
and U8615 (N_8615,N_8403,N_8398);
or U8616 (N_8616,N_8483,N_8391);
xnor U8617 (N_8617,N_8455,N_8431);
nand U8618 (N_8618,N_8430,N_8484);
or U8619 (N_8619,N_8429,N_8395);
xnor U8620 (N_8620,N_8432,N_8452);
nor U8621 (N_8621,N_8389,N_8424);
and U8622 (N_8622,N_8474,N_8497);
nand U8623 (N_8623,N_8391,N_8385);
and U8624 (N_8624,N_8441,N_8425);
nor U8625 (N_8625,N_8536,N_8503);
nor U8626 (N_8626,N_8569,N_8530);
nor U8627 (N_8627,N_8525,N_8508);
nor U8628 (N_8628,N_8572,N_8615);
or U8629 (N_8629,N_8551,N_8548);
xor U8630 (N_8630,N_8506,N_8592);
xnor U8631 (N_8631,N_8518,N_8554);
xor U8632 (N_8632,N_8558,N_8521);
nand U8633 (N_8633,N_8623,N_8564);
or U8634 (N_8634,N_8579,N_8581);
or U8635 (N_8635,N_8616,N_8586);
xnor U8636 (N_8636,N_8561,N_8513);
nor U8637 (N_8637,N_8500,N_8526);
nor U8638 (N_8638,N_8620,N_8597);
nor U8639 (N_8639,N_8618,N_8598);
xnor U8640 (N_8640,N_8585,N_8556);
and U8641 (N_8641,N_8529,N_8613);
and U8642 (N_8642,N_8540,N_8543);
and U8643 (N_8643,N_8574,N_8505);
and U8644 (N_8644,N_8565,N_8568);
nor U8645 (N_8645,N_8578,N_8571);
and U8646 (N_8646,N_8504,N_8609);
xor U8647 (N_8647,N_8527,N_8624);
or U8648 (N_8648,N_8570,N_8555);
nand U8649 (N_8649,N_8612,N_8514);
nor U8650 (N_8650,N_8537,N_8582);
nor U8651 (N_8651,N_8534,N_8516);
and U8652 (N_8652,N_8535,N_8509);
nand U8653 (N_8653,N_8602,N_8619);
and U8654 (N_8654,N_8550,N_8559);
or U8655 (N_8655,N_8575,N_8560);
and U8656 (N_8656,N_8608,N_8595);
or U8657 (N_8657,N_8567,N_8607);
and U8658 (N_8658,N_8528,N_8593);
xnor U8659 (N_8659,N_8510,N_8541);
nand U8660 (N_8660,N_8591,N_8600);
xor U8661 (N_8661,N_8524,N_8515);
and U8662 (N_8662,N_8617,N_8566);
nand U8663 (N_8663,N_8614,N_8532);
xor U8664 (N_8664,N_8587,N_8522);
nor U8665 (N_8665,N_8577,N_8610);
and U8666 (N_8666,N_8611,N_8544);
or U8667 (N_8667,N_8501,N_8512);
or U8668 (N_8668,N_8596,N_8563);
nand U8669 (N_8669,N_8604,N_8622);
xnor U8670 (N_8670,N_8517,N_8599);
and U8671 (N_8671,N_8502,N_8601);
and U8672 (N_8672,N_8523,N_8549);
and U8673 (N_8673,N_8605,N_8603);
nor U8674 (N_8674,N_8546,N_8533);
or U8675 (N_8675,N_8594,N_8519);
nand U8676 (N_8676,N_8553,N_8588);
nand U8677 (N_8677,N_8552,N_8580);
or U8678 (N_8678,N_8583,N_8562);
or U8679 (N_8679,N_8520,N_8545);
nor U8680 (N_8680,N_8542,N_8576);
and U8681 (N_8681,N_8511,N_8538);
and U8682 (N_8682,N_8531,N_8621);
or U8683 (N_8683,N_8590,N_8606);
or U8684 (N_8684,N_8557,N_8539);
xor U8685 (N_8685,N_8547,N_8584);
nand U8686 (N_8686,N_8507,N_8573);
nand U8687 (N_8687,N_8589,N_8508);
and U8688 (N_8688,N_8559,N_8621);
xor U8689 (N_8689,N_8589,N_8518);
and U8690 (N_8690,N_8585,N_8521);
xor U8691 (N_8691,N_8555,N_8622);
nor U8692 (N_8692,N_8612,N_8598);
xor U8693 (N_8693,N_8560,N_8566);
xnor U8694 (N_8694,N_8500,N_8583);
and U8695 (N_8695,N_8613,N_8592);
and U8696 (N_8696,N_8555,N_8504);
or U8697 (N_8697,N_8567,N_8604);
nand U8698 (N_8698,N_8574,N_8582);
nor U8699 (N_8699,N_8581,N_8615);
or U8700 (N_8700,N_8592,N_8558);
nand U8701 (N_8701,N_8570,N_8590);
or U8702 (N_8702,N_8590,N_8602);
xnor U8703 (N_8703,N_8506,N_8616);
and U8704 (N_8704,N_8604,N_8502);
or U8705 (N_8705,N_8506,N_8530);
nand U8706 (N_8706,N_8560,N_8592);
nand U8707 (N_8707,N_8605,N_8514);
xor U8708 (N_8708,N_8576,N_8588);
or U8709 (N_8709,N_8616,N_8611);
and U8710 (N_8710,N_8508,N_8564);
or U8711 (N_8711,N_8510,N_8567);
nand U8712 (N_8712,N_8502,N_8526);
xor U8713 (N_8713,N_8531,N_8586);
nand U8714 (N_8714,N_8582,N_8515);
xor U8715 (N_8715,N_8523,N_8577);
or U8716 (N_8716,N_8501,N_8544);
xnor U8717 (N_8717,N_8526,N_8587);
nand U8718 (N_8718,N_8501,N_8603);
or U8719 (N_8719,N_8543,N_8615);
nor U8720 (N_8720,N_8588,N_8589);
or U8721 (N_8721,N_8533,N_8515);
nand U8722 (N_8722,N_8540,N_8621);
nand U8723 (N_8723,N_8543,N_8619);
nor U8724 (N_8724,N_8591,N_8536);
or U8725 (N_8725,N_8543,N_8531);
xnor U8726 (N_8726,N_8511,N_8585);
nor U8727 (N_8727,N_8604,N_8562);
nand U8728 (N_8728,N_8618,N_8550);
xor U8729 (N_8729,N_8573,N_8546);
nand U8730 (N_8730,N_8622,N_8539);
nand U8731 (N_8731,N_8617,N_8622);
nand U8732 (N_8732,N_8603,N_8617);
nor U8733 (N_8733,N_8565,N_8523);
and U8734 (N_8734,N_8511,N_8551);
nand U8735 (N_8735,N_8584,N_8561);
nor U8736 (N_8736,N_8602,N_8573);
and U8737 (N_8737,N_8516,N_8519);
nand U8738 (N_8738,N_8613,N_8501);
nand U8739 (N_8739,N_8569,N_8559);
xor U8740 (N_8740,N_8515,N_8558);
and U8741 (N_8741,N_8603,N_8548);
nand U8742 (N_8742,N_8601,N_8524);
nor U8743 (N_8743,N_8525,N_8514);
xnor U8744 (N_8744,N_8592,N_8579);
and U8745 (N_8745,N_8502,N_8519);
or U8746 (N_8746,N_8577,N_8624);
or U8747 (N_8747,N_8584,N_8522);
and U8748 (N_8748,N_8534,N_8506);
xnor U8749 (N_8749,N_8592,N_8549);
nor U8750 (N_8750,N_8680,N_8730);
xor U8751 (N_8751,N_8699,N_8686);
xnor U8752 (N_8752,N_8650,N_8716);
nor U8753 (N_8753,N_8648,N_8745);
and U8754 (N_8754,N_8693,N_8689);
nor U8755 (N_8755,N_8640,N_8690);
nand U8756 (N_8756,N_8664,N_8704);
nand U8757 (N_8757,N_8637,N_8630);
xnor U8758 (N_8758,N_8719,N_8721);
nand U8759 (N_8759,N_8696,N_8705);
or U8760 (N_8760,N_8700,N_8677);
xnor U8761 (N_8761,N_8729,N_8651);
nand U8762 (N_8762,N_8702,N_8748);
xor U8763 (N_8763,N_8654,N_8692);
or U8764 (N_8764,N_8731,N_8652);
and U8765 (N_8765,N_8691,N_8679);
nand U8766 (N_8766,N_8649,N_8634);
nor U8767 (N_8767,N_8625,N_8744);
xor U8768 (N_8768,N_8697,N_8739);
or U8769 (N_8769,N_8627,N_8667);
and U8770 (N_8770,N_8707,N_8645);
nand U8771 (N_8771,N_8687,N_8647);
or U8772 (N_8772,N_8671,N_8646);
xnor U8773 (N_8773,N_8643,N_8669);
nand U8774 (N_8774,N_8714,N_8656);
xor U8775 (N_8775,N_8711,N_8694);
nor U8776 (N_8776,N_8712,N_8747);
xnor U8777 (N_8777,N_8715,N_8629);
xor U8778 (N_8778,N_8674,N_8628);
nand U8779 (N_8779,N_8746,N_8658);
nand U8780 (N_8780,N_8703,N_8743);
nor U8781 (N_8781,N_8661,N_8723);
and U8782 (N_8782,N_8720,N_8631);
and U8783 (N_8783,N_8636,N_8668);
nor U8784 (N_8784,N_8742,N_8688);
or U8785 (N_8785,N_8635,N_8732);
xor U8786 (N_8786,N_8659,N_8670);
and U8787 (N_8787,N_8725,N_8626);
nand U8788 (N_8788,N_8638,N_8655);
nand U8789 (N_8789,N_8713,N_8698);
or U8790 (N_8790,N_8737,N_8633);
nand U8791 (N_8791,N_8672,N_8644);
or U8792 (N_8792,N_8710,N_8632);
or U8793 (N_8793,N_8657,N_8665);
and U8794 (N_8794,N_8701,N_8736);
and U8795 (N_8795,N_8734,N_8662);
xor U8796 (N_8796,N_8663,N_8683);
nor U8797 (N_8797,N_8676,N_8728);
xnor U8798 (N_8798,N_8722,N_8653);
nand U8799 (N_8799,N_8685,N_8708);
nor U8800 (N_8800,N_8724,N_8749);
and U8801 (N_8801,N_8718,N_8641);
nor U8802 (N_8802,N_8681,N_8695);
or U8803 (N_8803,N_8733,N_8660);
or U8804 (N_8804,N_8639,N_8709);
nor U8805 (N_8805,N_8678,N_8684);
and U8806 (N_8806,N_8673,N_8735);
or U8807 (N_8807,N_8675,N_8642);
nand U8808 (N_8808,N_8727,N_8740);
nor U8809 (N_8809,N_8717,N_8741);
and U8810 (N_8810,N_8706,N_8682);
nor U8811 (N_8811,N_8666,N_8738);
xnor U8812 (N_8812,N_8726,N_8723);
or U8813 (N_8813,N_8672,N_8650);
nor U8814 (N_8814,N_8709,N_8748);
and U8815 (N_8815,N_8684,N_8746);
nand U8816 (N_8816,N_8728,N_8656);
nor U8817 (N_8817,N_8702,N_8714);
nand U8818 (N_8818,N_8707,N_8668);
xor U8819 (N_8819,N_8628,N_8725);
nor U8820 (N_8820,N_8627,N_8655);
and U8821 (N_8821,N_8746,N_8654);
nor U8822 (N_8822,N_8743,N_8652);
nor U8823 (N_8823,N_8704,N_8685);
or U8824 (N_8824,N_8682,N_8654);
nand U8825 (N_8825,N_8735,N_8723);
xor U8826 (N_8826,N_8744,N_8712);
or U8827 (N_8827,N_8634,N_8626);
nand U8828 (N_8828,N_8658,N_8722);
or U8829 (N_8829,N_8749,N_8672);
nor U8830 (N_8830,N_8736,N_8741);
nand U8831 (N_8831,N_8629,N_8737);
and U8832 (N_8832,N_8684,N_8648);
and U8833 (N_8833,N_8740,N_8743);
and U8834 (N_8834,N_8734,N_8681);
and U8835 (N_8835,N_8715,N_8628);
nor U8836 (N_8836,N_8637,N_8712);
and U8837 (N_8837,N_8722,N_8734);
xor U8838 (N_8838,N_8739,N_8689);
xnor U8839 (N_8839,N_8707,N_8739);
and U8840 (N_8840,N_8745,N_8657);
xnor U8841 (N_8841,N_8743,N_8738);
and U8842 (N_8842,N_8708,N_8669);
and U8843 (N_8843,N_8635,N_8659);
xnor U8844 (N_8844,N_8739,N_8734);
xnor U8845 (N_8845,N_8630,N_8676);
or U8846 (N_8846,N_8660,N_8674);
nor U8847 (N_8847,N_8637,N_8727);
or U8848 (N_8848,N_8663,N_8682);
or U8849 (N_8849,N_8742,N_8647);
xor U8850 (N_8850,N_8633,N_8638);
nor U8851 (N_8851,N_8719,N_8626);
nor U8852 (N_8852,N_8695,N_8706);
or U8853 (N_8853,N_8729,N_8646);
or U8854 (N_8854,N_8690,N_8663);
nand U8855 (N_8855,N_8640,N_8748);
nand U8856 (N_8856,N_8684,N_8730);
nand U8857 (N_8857,N_8728,N_8647);
xor U8858 (N_8858,N_8738,N_8740);
xnor U8859 (N_8859,N_8745,N_8743);
xor U8860 (N_8860,N_8743,N_8699);
or U8861 (N_8861,N_8647,N_8747);
and U8862 (N_8862,N_8657,N_8731);
nand U8863 (N_8863,N_8648,N_8748);
nor U8864 (N_8864,N_8670,N_8671);
xnor U8865 (N_8865,N_8698,N_8695);
nor U8866 (N_8866,N_8693,N_8711);
xor U8867 (N_8867,N_8707,N_8650);
and U8868 (N_8868,N_8626,N_8658);
nand U8869 (N_8869,N_8638,N_8730);
and U8870 (N_8870,N_8747,N_8737);
nand U8871 (N_8871,N_8660,N_8713);
nor U8872 (N_8872,N_8726,N_8738);
nand U8873 (N_8873,N_8687,N_8738);
xnor U8874 (N_8874,N_8714,N_8635);
or U8875 (N_8875,N_8796,N_8793);
and U8876 (N_8876,N_8810,N_8855);
nand U8877 (N_8877,N_8785,N_8841);
xnor U8878 (N_8878,N_8777,N_8853);
and U8879 (N_8879,N_8820,N_8756);
or U8880 (N_8880,N_8839,N_8856);
nor U8881 (N_8881,N_8773,N_8852);
xnor U8882 (N_8882,N_8857,N_8761);
xor U8883 (N_8883,N_8800,N_8817);
and U8884 (N_8884,N_8873,N_8847);
or U8885 (N_8885,N_8818,N_8845);
and U8886 (N_8886,N_8754,N_8781);
and U8887 (N_8887,N_8782,N_8752);
and U8888 (N_8888,N_8794,N_8836);
xnor U8889 (N_8889,N_8823,N_8751);
nand U8890 (N_8890,N_8872,N_8860);
and U8891 (N_8891,N_8757,N_8868);
and U8892 (N_8892,N_8828,N_8806);
or U8893 (N_8893,N_8816,N_8833);
and U8894 (N_8894,N_8774,N_8813);
xnor U8895 (N_8895,N_8861,N_8768);
nand U8896 (N_8896,N_8797,N_8770);
or U8897 (N_8897,N_8831,N_8815);
or U8898 (N_8898,N_8775,N_8863);
nor U8899 (N_8899,N_8829,N_8783);
and U8900 (N_8900,N_8870,N_8753);
nor U8901 (N_8901,N_8784,N_8843);
or U8902 (N_8902,N_8865,N_8838);
xnor U8903 (N_8903,N_8786,N_8776);
or U8904 (N_8904,N_8814,N_8851);
nand U8905 (N_8905,N_8826,N_8805);
xnor U8906 (N_8906,N_8825,N_8801);
nor U8907 (N_8907,N_8772,N_8755);
nor U8908 (N_8908,N_8779,N_8811);
nor U8909 (N_8909,N_8802,N_8798);
nand U8910 (N_8910,N_8763,N_8791);
or U8911 (N_8911,N_8799,N_8807);
nand U8912 (N_8912,N_8780,N_8862);
or U8913 (N_8913,N_8758,N_8869);
nor U8914 (N_8914,N_8771,N_8790);
and U8915 (N_8915,N_8767,N_8859);
xor U8916 (N_8916,N_8778,N_8789);
xnor U8917 (N_8917,N_8835,N_8858);
xnor U8918 (N_8918,N_8760,N_8822);
xnor U8919 (N_8919,N_8824,N_8795);
or U8920 (N_8920,N_8809,N_8866);
nand U8921 (N_8921,N_8766,N_8834);
and U8922 (N_8922,N_8871,N_8792);
xnor U8923 (N_8923,N_8850,N_8804);
xnor U8924 (N_8924,N_8819,N_8837);
and U8925 (N_8925,N_8788,N_8750);
xnor U8926 (N_8926,N_8867,N_8759);
nor U8927 (N_8927,N_8874,N_8827);
and U8928 (N_8928,N_8844,N_8830);
xnor U8929 (N_8929,N_8840,N_8812);
nor U8930 (N_8930,N_8842,N_8769);
nor U8931 (N_8931,N_8764,N_8808);
nand U8932 (N_8932,N_8821,N_8848);
nor U8933 (N_8933,N_8765,N_8854);
xnor U8934 (N_8934,N_8849,N_8832);
and U8935 (N_8935,N_8846,N_8864);
and U8936 (N_8936,N_8787,N_8762);
xor U8937 (N_8937,N_8803,N_8775);
nor U8938 (N_8938,N_8860,N_8815);
nand U8939 (N_8939,N_8873,N_8843);
nand U8940 (N_8940,N_8852,N_8798);
xnor U8941 (N_8941,N_8858,N_8799);
or U8942 (N_8942,N_8803,N_8770);
xor U8943 (N_8943,N_8826,N_8868);
or U8944 (N_8944,N_8841,N_8791);
and U8945 (N_8945,N_8850,N_8769);
nor U8946 (N_8946,N_8833,N_8766);
nand U8947 (N_8947,N_8870,N_8817);
xnor U8948 (N_8948,N_8755,N_8780);
nand U8949 (N_8949,N_8834,N_8836);
and U8950 (N_8950,N_8769,N_8757);
nor U8951 (N_8951,N_8793,N_8797);
and U8952 (N_8952,N_8799,N_8868);
nor U8953 (N_8953,N_8868,N_8758);
or U8954 (N_8954,N_8873,N_8794);
and U8955 (N_8955,N_8788,N_8755);
and U8956 (N_8956,N_8764,N_8851);
xnor U8957 (N_8957,N_8800,N_8873);
or U8958 (N_8958,N_8844,N_8794);
or U8959 (N_8959,N_8782,N_8869);
and U8960 (N_8960,N_8873,N_8830);
xnor U8961 (N_8961,N_8819,N_8760);
nor U8962 (N_8962,N_8802,N_8786);
or U8963 (N_8963,N_8873,N_8805);
or U8964 (N_8964,N_8831,N_8791);
and U8965 (N_8965,N_8761,N_8806);
xor U8966 (N_8966,N_8829,N_8818);
nand U8967 (N_8967,N_8870,N_8825);
nor U8968 (N_8968,N_8820,N_8805);
nand U8969 (N_8969,N_8768,N_8837);
nand U8970 (N_8970,N_8827,N_8825);
nand U8971 (N_8971,N_8787,N_8815);
and U8972 (N_8972,N_8827,N_8823);
and U8973 (N_8973,N_8810,N_8833);
nand U8974 (N_8974,N_8793,N_8801);
xnor U8975 (N_8975,N_8763,N_8848);
nand U8976 (N_8976,N_8873,N_8758);
and U8977 (N_8977,N_8837,N_8772);
or U8978 (N_8978,N_8841,N_8774);
or U8979 (N_8979,N_8841,N_8840);
and U8980 (N_8980,N_8836,N_8774);
and U8981 (N_8981,N_8767,N_8799);
nor U8982 (N_8982,N_8775,N_8750);
nand U8983 (N_8983,N_8830,N_8839);
or U8984 (N_8984,N_8808,N_8799);
nand U8985 (N_8985,N_8804,N_8776);
and U8986 (N_8986,N_8871,N_8854);
nor U8987 (N_8987,N_8824,N_8862);
xor U8988 (N_8988,N_8797,N_8816);
or U8989 (N_8989,N_8865,N_8825);
xnor U8990 (N_8990,N_8794,N_8862);
and U8991 (N_8991,N_8751,N_8862);
or U8992 (N_8992,N_8808,N_8812);
nand U8993 (N_8993,N_8752,N_8836);
and U8994 (N_8994,N_8796,N_8843);
and U8995 (N_8995,N_8829,N_8787);
nor U8996 (N_8996,N_8793,N_8843);
and U8997 (N_8997,N_8759,N_8792);
nor U8998 (N_8998,N_8785,N_8794);
nand U8999 (N_8999,N_8807,N_8795);
nor U9000 (N_9000,N_8896,N_8885);
and U9001 (N_9001,N_8916,N_8887);
nand U9002 (N_9002,N_8927,N_8883);
nand U9003 (N_9003,N_8950,N_8905);
or U9004 (N_9004,N_8965,N_8930);
or U9005 (N_9005,N_8918,N_8989);
xnor U9006 (N_9006,N_8877,N_8907);
nand U9007 (N_9007,N_8892,N_8881);
nand U9008 (N_9008,N_8937,N_8976);
and U9009 (N_9009,N_8948,N_8924);
xnor U9010 (N_9010,N_8914,N_8879);
xor U9011 (N_9011,N_8941,N_8934);
or U9012 (N_9012,N_8998,N_8991);
nand U9013 (N_9013,N_8899,N_8895);
or U9014 (N_9014,N_8897,N_8969);
nor U9015 (N_9015,N_8977,N_8982);
or U9016 (N_9016,N_8954,N_8943);
and U9017 (N_9017,N_8888,N_8964);
nor U9018 (N_9018,N_8882,N_8952);
xor U9019 (N_9019,N_8901,N_8900);
and U9020 (N_9020,N_8909,N_8960);
nor U9021 (N_9021,N_8995,N_8876);
nand U9022 (N_9022,N_8957,N_8935);
and U9023 (N_9023,N_8922,N_8939);
nor U9024 (N_9024,N_8926,N_8908);
and U9025 (N_9025,N_8903,N_8981);
and U9026 (N_9026,N_8893,N_8985);
nor U9027 (N_9027,N_8915,N_8999);
xor U9028 (N_9028,N_8972,N_8945);
or U9029 (N_9029,N_8890,N_8955);
or U9030 (N_9030,N_8938,N_8912);
xor U9031 (N_9031,N_8980,N_8884);
nand U9032 (N_9032,N_8913,N_8936);
xor U9033 (N_9033,N_8933,N_8917);
nand U9034 (N_9034,N_8947,N_8928);
or U9035 (N_9035,N_8974,N_8946);
or U9036 (N_9036,N_8894,N_8971);
nor U9037 (N_9037,N_8973,N_8932);
or U9038 (N_9038,N_8940,N_8949);
nand U9039 (N_9039,N_8959,N_8910);
xor U9040 (N_9040,N_8923,N_8986);
or U9041 (N_9041,N_8962,N_8956);
and U9042 (N_9042,N_8994,N_8920);
nand U9043 (N_9043,N_8966,N_8875);
and U9044 (N_9044,N_8889,N_8979);
nand U9045 (N_9045,N_8951,N_8987);
xnor U9046 (N_9046,N_8961,N_8978);
nand U9047 (N_9047,N_8911,N_8898);
and U9048 (N_9048,N_8942,N_8953);
xnor U9049 (N_9049,N_8988,N_8958);
or U9050 (N_9050,N_8925,N_8963);
nand U9051 (N_9051,N_8996,N_8891);
or U9052 (N_9052,N_8904,N_8983);
and U9053 (N_9053,N_8880,N_8902);
and U9054 (N_9054,N_8984,N_8997);
nor U9055 (N_9055,N_8993,N_8929);
and U9056 (N_9056,N_8975,N_8970);
nand U9057 (N_9057,N_8921,N_8878);
nand U9058 (N_9058,N_8968,N_8990);
nor U9059 (N_9059,N_8931,N_8906);
nor U9060 (N_9060,N_8967,N_8992);
nor U9061 (N_9061,N_8919,N_8886);
nand U9062 (N_9062,N_8944,N_8949);
xnor U9063 (N_9063,N_8990,N_8953);
nand U9064 (N_9064,N_8966,N_8942);
nor U9065 (N_9065,N_8885,N_8906);
or U9066 (N_9066,N_8953,N_8975);
nor U9067 (N_9067,N_8909,N_8990);
xor U9068 (N_9068,N_8977,N_8876);
xnor U9069 (N_9069,N_8967,N_8991);
nand U9070 (N_9070,N_8906,N_8903);
or U9071 (N_9071,N_8981,N_8945);
and U9072 (N_9072,N_8988,N_8888);
xor U9073 (N_9073,N_8932,N_8898);
and U9074 (N_9074,N_8905,N_8890);
nand U9075 (N_9075,N_8905,N_8911);
xnor U9076 (N_9076,N_8995,N_8878);
or U9077 (N_9077,N_8911,N_8978);
nand U9078 (N_9078,N_8993,N_8988);
nand U9079 (N_9079,N_8919,N_8918);
or U9080 (N_9080,N_8973,N_8880);
xor U9081 (N_9081,N_8989,N_8881);
or U9082 (N_9082,N_8966,N_8969);
nand U9083 (N_9083,N_8877,N_8930);
nand U9084 (N_9084,N_8887,N_8932);
nand U9085 (N_9085,N_8912,N_8878);
xor U9086 (N_9086,N_8892,N_8954);
or U9087 (N_9087,N_8979,N_8930);
and U9088 (N_9088,N_8890,N_8896);
xor U9089 (N_9089,N_8906,N_8965);
nor U9090 (N_9090,N_8895,N_8935);
xnor U9091 (N_9091,N_8961,N_8965);
and U9092 (N_9092,N_8914,N_8948);
xor U9093 (N_9093,N_8962,N_8954);
xnor U9094 (N_9094,N_8916,N_8937);
nor U9095 (N_9095,N_8910,N_8888);
and U9096 (N_9096,N_8920,N_8914);
xor U9097 (N_9097,N_8894,N_8956);
or U9098 (N_9098,N_8936,N_8931);
xor U9099 (N_9099,N_8993,N_8878);
nand U9100 (N_9100,N_8945,N_8950);
and U9101 (N_9101,N_8884,N_8894);
nand U9102 (N_9102,N_8978,N_8951);
nand U9103 (N_9103,N_8907,N_8925);
nand U9104 (N_9104,N_8995,N_8984);
and U9105 (N_9105,N_8947,N_8896);
nand U9106 (N_9106,N_8989,N_8900);
xor U9107 (N_9107,N_8879,N_8902);
nor U9108 (N_9108,N_8943,N_8917);
nor U9109 (N_9109,N_8897,N_8906);
xnor U9110 (N_9110,N_8931,N_8881);
or U9111 (N_9111,N_8884,N_8939);
nor U9112 (N_9112,N_8985,N_8977);
or U9113 (N_9113,N_8947,N_8998);
nor U9114 (N_9114,N_8881,N_8952);
xnor U9115 (N_9115,N_8938,N_8973);
nand U9116 (N_9116,N_8924,N_8967);
nor U9117 (N_9117,N_8991,N_8981);
and U9118 (N_9118,N_8892,N_8943);
and U9119 (N_9119,N_8980,N_8958);
nand U9120 (N_9120,N_8987,N_8956);
or U9121 (N_9121,N_8981,N_8890);
or U9122 (N_9122,N_8997,N_8935);
nor U9123 (N_9123,N_8916,N_8917);
nor U9124 (N_9124,N_8877,N_8976);
xor U9125 (N_9125,N_9077,N_9021);
or U9126 (N_9126,N_9062,N_9094);
or U9127 (N_9127,N_9096,N_9113);
xor U9128 (N_9128,N_9080,N_9058);
and U9129 (N_9129,N_9007,N_9029);
nand U9130 (N_9130,N_9117,N_9037);
nand U9131 (N_9131,N_9067,N_9009);
nand U9132 (N_9132,N_9033,N_9044);
xnor U9133 (N_9133,N_9065,N_9024);
nand U9134 (N_9134,N_9122,N_9098);
and U9135 (N_9135,N_9015,N_9063);
or U9136 (N_9136,N_9038,N_9006);
nor U9137 (N_9137,N_9057,N_9073);
xor U9138 (N_9138,N_9023,N_9056);
or U9139 (N_9139,N_9012,N_9079);
nor U9140 (N_9140,N_9074,N_9008);
and U9141 (N_9141,N_9114,N_9035);
and U9142 (N_9142,N_9052,N_9048);
or U9143 (N_9143,N_9103,N_9032);
xnor U9144 (N_9144,N_9076,N_9014);
and U9145 (N_9145,N_9016,N_9115);
or U9146 (N_9146,N_9053,N_9100);
and U9147 (N_9147,N_9121,N_9059);
or U9148 (N_9148,N_9020,N_9085);
xnor U9149 (N_9149,N_9105,N_9041);
nor U9150 (N_9150,N_9064,N_9099);
nor U9151 (N_9151,N_9072,N_9089);
xor U9152 (N_9152,N_9054,N_9061);
or U9153 (N_9153,N_9026,N_9019);
nand U9154 (N_9154,N_9111,N_9066);
or U9155 (N_9155,N_9071,N_9083);
nor U9156 (N_9156,N_9092,N_9123);
nand U9157 (N_9157,N_9060,N_9082);
and U9158 (N_9158,N_9018,N_9107);
xor U9159 (N_9159,N_9124,N_9116);
xor U9160 (N_9160,N_9010,N_9091);
and U9161 (N_9161,N_9034,N_9011);
nor U9162 (N_9162,N_9027,N_9078);
or U9163 (N_9163,N_9050,N_9005);
or U9164 (N_9164,N_9097,N_9087);
and U9165 (N_9165,N_9051,N_9104);
xnor U9166 (N_9166,N_9075,N_9109);
nor U9167 (N_9167,N_9046,N_9022);
and U9168 (N_9168,N_9000,N_9040);
nor U9169 (N_9169,N_9028,N_9081);
xnor U9170 (N_9170,N_9049,N_9047);
or U9171 (N_9171,N_9045,N_9070);
xor U9172 (N_9172,N_9110,N_9042);
and U9173 (N_9173,N_9036,N_9013);
or U9174 (N_9174,N_9108,N_9088);
or U9175 (N_9175,N_9101,N_9017);
or U9176 (N_9176,N_9095,N_9068);
nand U9177 (N_9177,N_9039,N_9106);
or U9178 (N_9178,N_9025,N_9031);
xnor U9179 (N_9179,N_9112,N_9102);
xnor U9180 (N_9180,N_9086,N_9003);
and U9181 (N_9181,N_9090,N_9120);
and U9182 (N_9182,N_9119,N_9004);
or U9183 (N_9183,N_9030,N_9069);
nand U9184 (N_9184,N_9055,N_9043);
or U9185 (N_9185,N_9084,N_9118);
nor U9186 (N_9186,N_9001,N_9002);
nand U9187 (N_9187,N_9093,N_9049);
xor U9188 (N_9188,N_9002,N_9067);
xor U9189 (N_9189,N_9116,N_9033);
xnor U9190 (N_9190,N_9006,N_9107);
and U9191 (N_9191,N_9073,N_9080);
and U9192 (N_9192,N_9076,N_9124);
nor U9193 (N_9193,N_9038,N_9031);
nor U9194 (N_9194,N_9049,N_9069);
or U9195 (N_9195,N_9116,N_9105);
xnor U9196 (N_9196,N_9031,N_9056);
nor U9197 (N_9197,N_9037,N_9011);
or U9198 (N_9198,N_9073,N_9072);
nor U9199 (N_9199,N_9099,N_9066);
and U9200 (N_9200,N_9091,N_9012);
or U9201 (N_9201,N_9117,N_9073);
and U9202 (N_9202,N_9071,N_9010);
nor U9203 (N_9203,N_9021,N_9033);
and U9204 (N_9204,N_9044,N_9106);
xnor U9205 (N_9205,N_9109,N_9124);
nor U9206 (N_9206,N_9070,N_9003);
nor U9207 (N_9207,N_9102,N_9072);
nor U9208 (N_9208,N_9073,N_9071);
nor U9209 (N_9209,N_9091,N_9101);
xor U9210 (N_9210,N_9110,N_9043);
xnor U9211 (N_9211,N_9017,N_9060);
or U9212 (N_9212,N_9117,N_9095);
and U9213 (N_9213,N_9110,N_9001);
nor U9214 (N_9214,N_9015,N_9036);
and U9215 (N_9215,N_9037,N_9077);
nand U9216 (N_9216,N_9028,N_9091);
or U9217 (N_9217,N_9089,N_9018);
nand U9218 (N_9218,N_9077,N_9080);
and U9219 (N_9219,N_9098,N_9017);
nor U9220 (N_9220,N_9072,N_9045);
or U9221 (N_9221,N_9031,N_9100);
and U9222 (N_9222,N_9093,N_9112);
and U9223 (N_9223,N_9028,N_9089);
nor U9224 (N_9224,N_9013,N_9025);
or U9225 (N_9225,N_9088,N_9004);
and U9226 (N_9226,N_9062,N_9028);
or U9227 (N_9227,N_9104,N_9065);
and U9228 (N_9228,N_9024,N_9092);
and U9229 (N_9229,N_9042,N_9085);
xor U9230 (N_9230,N_9088,N_9027);
nor U9231 (N_9231,N_9058,N_9049);
xor U9232 (N_9232,N_9096,N_9022);
xor U9233 (N_9233,N_9047,N_9004);
and U9234 (N_9234,N_9073,N_9090);
xnor U9235 (N_9235,N_9110,N_9123);
xor U9236 (N_9236,N_9084,N_9029);
xor U9237 (N_9237,N_9032,N_9067);
nand U9238 (N_9238,N_9013,N_9123);
or U9239 (N_9239,N_9002,N_9096);
or U9240 (N_9240,N_9056,N_9012);
nand U9241 (N_9241,N_9065,N_9111);
or U9242 (N_9242,N_9060,N_9058);
nand U9243 (N_9243,N_9030,N_9102);
nor U9244 (N_9244,N_9049,N_9096);
or U9245 (N_9245,N_9026,N_9054);
nor U9246 (N_9246,N_9117,N_9008);
and U9247 (N_9247,N_9048,N_9091);
or U9248 (N_9248,N_9014,N_9005);
or U9249 (N_9249,N_9084,N_9019);
or U9250 (N_9250,N_9158,N_9153);
nor U9251 (N_9251,N_9185,N_9169);
and U9252 (N_9252,N_9188,N_9160);
nand U9253 (N_9253,N_9203,N_9176);
xor U9254 (N_9254,N_9215,N_9181);
or U9255 (N_9255,N_9128,N_9211);
xnor U9256 (N_9256,N_9177,N_9205);
and U9257 (N_9257,N_9240,N_9237);
nor U9258 (N_9258,N_9156,N_9207);
or U9259 (N_9259,N_9150,N_9179);
or U9260 (N_9260,N_9129,N_9209);
xor U9261 (N_9261,N_9152,N_9242);
nand U9262 (N_9262,N_9157,N_9196);
nand U9263 (N_9263,N_9241,N_9218);
nand U9264 (N_9264,N_9151,N_9194);
nand U9265 (N_9265,N_9161,N_9217);
nand U9266 (N_9266,N_9133,N_9140);
nor U9267 (N_9267,N_9142,N_9171);
nand U9268 (N_9268,N_9130,N_9132);
nand U9269 (N_9269,N_9219,N_9225);
nor U9270 (N_9270,N_9146,N_9214);
and U9271 (N_9271,N_9248,N_9197);
nand U9272 (N_9272,N_9235,N_9172);
nand U9273 (N_9273,N_9147,N_9144);
or U9274 (N_9274,N_9206,N_9247);
xnor U9275 (N_9275,N_9210,N_9127);
nand U9276 (N_9276,N_9134,N_9208);
nand U9277 (N_9277,N_9154,N_9192);
nor U9278 (N_9278,N_9180,N_9249);
and U9279 (N_9279,N_9182,N_9229);
nand U9280 (N_9280,N_9200,N_9245);
and U9281 (N_9281,N_9126,N_9226);
xor U9282 (N_9282,N_9239,N_9216);
or U9283 (N_9283,N_9187,N_9204);
xnor U9284 (N_9284,N_9148,N_9174);
or U9285 (N_9285,N_9201,N_9143);
xor U9286 (N_9286,N_9212,N_9168);
xor U9287 (N_9287,N_9183,N_9141);
xnor U9288 (N_9288,N_9145,N_9167);
xor U9289 (N_9289,N_9131,N_9202);
nor U9290 (N_9290,N_9213,N_9155);
nor U9291 (N_9291,N_9223,N_9138);
xnor U9292 (N_9292,N_9166,N_9222);
nor U9293 (N_9293,N_9224,N_9186);
or U9294 (N_9294,N_9135,N_9191);
nand U9295 (N_9295,N_9230,N_9159);
xnor U9296 (N_9296,N_9163,N_9233);
nor U9297 (N_9297,N_9165,N_9244);
nand U9298 (N_9298,N_9162,N_9231);
xor U9299 (N_9299,N_9189,N_9243);
nand U9300 (N_9300,N_9173,N_9193);
or U9301 (N_9301,N_9227,N_9236);
and U9302 (N_9302,N_9190,N_9221);
xnor U9303 (N_9303,N_9136,N_9246);
nand U9304 (N_9304,N_9164,N_9137);
nand U9305 (N_9305,N_9178,N_9184);
or U9306 (N_9306,N_9232,N_9234);
and U9307 (N_9307,N_9199,N_9228);
nor U9308 (N_9308,N_9149,N_9139);
and U9309 (N_9309,N_9220,N_9170);
nor U9310 (N_9310,N_9198,N_9175);
xor U9311 (N_9311,N_9238,N_9195);
xor U9312 (N_9312,N_9125,N_9239);
or U9313 (N_9313,N_9154,N_9130);
nand U9314 (N_9314,N_9142,N_9235);
nand U9315 (N_9315,N_9178,N_9126);
or U9316 (N_9316,N_9183,N_9128);
or U9317 (N_9317,N_9202,N_9152);
nand U9318 (N_9318,N_9133,N_9228);
xor U9319 (N_9319,N_9248,N_9169);
or U9320 (N_9320,N_9175,N_9206);
xnor U9321 (N_9321,N_9245,N_9204);
nor U9322 (N_9322,N_9225,N_9246);
nor U9323 (N_9323,N_9125,N_9128);
and U9324 (N_9324,N_9183,N_9197);
or U9325 (N_9325,N_9133,N_9214);
nand U9326 (N_9326,N_9161,N_9230);
or U9327 (N_9327,N_9212,N_9246);
nand U9328 (N_9328,N_9241,N_9194);
xnor U9329 (N_9329,N_9157,N_9183);
xnor U9330 (N_9330,N_9158,N_9227);
or U9331 (N_9331,N_9182,N_9159);
nand U9332 (N_9332,N_9174,N_9154);
and U9333 (N_9333,N_9233,N_9207);
nand U9334 (N_9334,N_9238,N_9151);
nor U9335 (N_9335,N_9225,N_9130);
or U9336 (N_9336,N_9133,N_9224);
and U9337 (N_9337,N_9235,N_9137);
xnor U9338 (N_9338,N_9202,N_9132);
or U9339 (N_9339,N_9224,N_9196);
or U9340 (N_9340,N_9245,N_9237);
or U9341 (N_9341,N_9248,N_9183);
and U9342 (N_9342,N_9179,N_9242);
or U9343 (N_9343,N_9241,N_9208);
nand U9344 (N_9344,N_9183,N_9196);
xor U9345 (N_9345,N_9165,N_9247);
and U9346 (N_9346,N_9155,N_9174);
xor U9347 (N_9347,N_9239,N_9153);
or U9348 (N_9348,N_9171,N_9168);
or U9349 (N_9349,N_9149,N_9220);
nor U9350 (N_9350,N_9173,N_9202);
xnor U9351 (N_9351,N_9220,N_9204);
and U9352 (N_9352,N_9225,N_9141);
nand U9353 (N_9353,N_9199,N_9187);
and U9354 (N_9354,N_9195,N_9240);
nand U9355 (N_9355,N_9217,N_9148);
or U9356 (N_9356,N_9185,N_9196);
or U9357 (N_9357,N_9220,N_9167);
nor U9358 (N_9358,N_9199,N_9147);
nor U9359 (N_9359,N_9179,N_9229);
xnor U9360 (N_9360,N_9213,N_9143);
and U9361 (N_9361,N_9125,N_9245);
and U9362 (N_9362,N_9236,N_9166);
nor U9363 (N_9363,N_9226,N_9165);
nor U9364 (N_9364,N_9174,N_9161);
or U9365 (N_9365,N_9214,N_9242);
or U9366 (N_9366,N_9147,N_9134);
and U9367 (N_9367,N_9228,N_9195);
nor U9368 (N_9368,N_9222,N_9245);
xnor U9369 (N_9369,N_9150,N_9186);
nor U9370 (N_9370,N_9228,N_9146);
nand U9371 (N_9371,N_9168,N_9248);
nand U9372 (N_9372,N_9220,N_9199);
or U9373 (N_9373,N_9234,N_9148);
xor U9374 (N_9374,N_9200,N_9134);
nor U9375 (N_9375,N_9265,N_9304);
and U9376 (N_9376,N_9367,N_9319);
or U9377 (N_9377,N_9271,N_9284);
xor U9378 (N_9378,N_9326,N_9252);
nand U9379 (N_9379,N_9341,N_9358);
nor U9380 (N_9380,N_9331,N_9307);
and U9381 (N_9381,N_9321,N_9296);
nor U9382 (N_9382,N_9350,N_9337);
xnor U9383 (N_9383,N_9298,N_9324);
and U9384 (N_9384,N_9270,N_9274);
xnor U9385 (N_9385,N_9363,N_9255);
or U9386 (N_9386,N_9339,N_9365);
or U9387 (N_9387,N_9335,N_9366);
or U9388 (N_9388,N_9287,N_9317);
xor U9389 (N_9389,N_9286,N_9300);
xnor U9390 (N_9390,N_9344,N_9254);
nand U9391 (N_9391,N_9374,N_9313);
and U9392 (N_9392,N_9261,N_9311);
xnor U9393 (N_9393,N_9281,N_9276);
nand U9394 (N_9394,N_9314,N_9299);
nand U9395 (N_9395,N_9273,N_9347);
xor U9396 (N_9396,N_9332,N_9318);
or U9397 (N_9397,N_9343,N_9302);
xnor U9398 (N_9398,N_9334,N_9301);
and U9399 (N_9399,N_9278,N_9362);
or U9400 (N_9400,N_9258,N_9269);
xor U9401 (N_9401,N_9306,N_9303);
nand U9402 (N_9402,N_9309,N_9312);
nor U9403 (N_9403,N_9355,N_9369);
nor U9404 (N_9404,N_9280,N_9293);
nand U9405 (N_9405,N_9360,N_9354);
nor U9406 (N_9406,N_9330,N_9349);
and U9407 (N_9407,N_9289,N_9325);
xnor U9408 (N_9408,N_9372,N_9257);
xor U9409 (N_9409,N_9268,N_9338);
xor U9410 (N_9410,N_9297,N_9294);
nand U9411 (N_9411,N_9345,N_9322);
and U9412 (N_9412,N_9327,N_9251);
nand U9413 (N_9413,N_9277,N_9279);
nor U9414 (N_9414,N_9368,N_9259);
and U9415 (N_9415,N_9260,N_9266);
and U9416 (N_9416,N_9373,N_9310);
xor U9417 (N_9417,N_9357,N_9250);
nor U9418 (N_9418,N_9256,N_9364);
or U9419 (N_9419,N_9267,N_9264);
xor U9420 (N_9420,N_9361,N_9305);
nand U9421 (N_9421,N_9371,N_9353);
nor U9422 (N_9422,N_9333,N_9351);
and U9423 (N_9423,N_9282,N_9323);
and U9424 (N_9424,N_9340,N_9329);
xor U9425 (N_9425,N_9292,N_9346);
and U9426 (N_9426,N_9285,N_9342);
nor U9427 (N_9427,N_9308,N_9263);
nand U9428 (N_9428,N_9272,N_9316);
or U9429 (N_9429,N_9352,N_9356);
nor U9430 (N_9430,N_9328,N_9253);
nand U9431 (N_9431,N_9283,N_9336);
nand U9432 (N_9432,N_9315,N_9290);
nand U9433 (N_9433,N_9320,N_9291);
and U9434 (N_9434,N_9295,N_9370);
or U9435 (N_9435,N_9288,N_9359);
or U9436 (N_9436,N_9348,N_9275);
xnor U9437 (N_9437,N_9262,N_9315);
xnor U9438 (N_9438,N_9265,N_9362);
nor U9439 (N_9439,N_9266,N_9309);
and U9440 (N_9440,N_9346,N_9260);
and U9441 (N_9441,N_9362,N_9285);
nor U9442 (N_9442,N_9374,N_9353);
or U9443 (N_9443,N_9270,N_9347);
xor U9444 (N_9444,N_9324,N_9274);
xor U9445 (N_9445,N_9328,N_9250);
nand U9446 (N_9446,N_9322,N_9273);
xor U9447 (N_9447,N_9325,N_9348);
nor U9448 (N_9448,N_9301,N_9295);
nand U9449 (N_9449,N_9329,N_9268);
and U9450 (N_9450,N_9295,N_9333);
xor U9451 (N_9451,N_9326,N_9268);
or U9452 (N_9452,N_9305,N_9300);
and U9453 (N_9453,N_9300,N_9370);
nand U9454 (N_9454,N_9250,N_9294);
nand U9455 (N_9455,N_9344,N_9354);
nor U9456 (N_9456,N_9370,N_9341);
nor U9457 (N_9457,N_9338,N_9367);
and U9458 (N_9458,N_9356,N_9336);
and U9459 (N_9459,N_9347,N_9295);
nor U9460 (N_9460,N_9369,N_9278);
and U9461 (N_9461,N_9280,N_9291);
and U9462 (N_9462,N_9331,N_9347);
or U9463 (N_9463,N_9291,N_9301);
xor U9464 (N_9464,N_9336,N_9331);
and U9465 (N_9465,N_9254,N_9315);
and U9466 (N_9466,N_9288,N_9258);
nor U9467 (N_9467,N_9284,N_9373);
and U9468 (N_9468,N_9322,N_9268);
nor U9469 (N_9469,N_9281,N_9351);
xor U9470 (N_9470,N_9297,N_9342);
and U9471 (N_9471,N_9355,N_9331);
nand U9472 (N_9472,N_9262,N_9261);
or U9473 (N_9473,N_9279,N_9265);
nand U9474 (N_9474,N_9272,N_9366);
nor U9475 (N_9475,N_9266,N_9354);
nor U9476 (N_9476,N_9353,N_9308);
nor U9477 (N_9477,N_9371,N_9365);
xor U9478 (N_9478,N_9331,N_9257);
nand U9479 (N_9479,N_9293,N_9373);
nand U9480 (N_9480,N_9368,N_9295);
nor U9481 (N_9481,N_9274,N_9317);
nand U9482 (N_9482,N_9272,N_9336);
nor U9483 (N_9483,N_9295,N_9332);
xnor U9484 (N_9484,N_9322,N_9357);
xor U9485 (N_9485,N_9287,N_9330);
or U9486 (N_9486,N_9345,N_9254);
nand U9487 (N_9487,N_9366,N_9374);
nor U9488 (N_9488,N_9362,N_9252);
and U9489 (N_9489,N_9319,N_9300);
nand U9490 (N_9490,N_9288,N_9362);
and U9491 (N_9491,N_9315,N_9282);
xor U9492 (N_9492,N_9295,N_9350);
nand U9493 (N_9493,N_9354,N_9334);
nor U9494 (N_9494,N_9337,N_9302);
and U9495 (N_9495,N_9361,N_9268);
xor U9496 (N_9496,N_9337,N_9317);
and U9497 (N_9497,N_9276,N_9325);
or U9498 (N_9498,N_9350,N_9294);
nor U9499 (N_9499,N_9315,N_9343);
nand U9500 (N_9500,N_9450,N_9377);
and U9501 (N_9501,N_9478,N_9405);
nand U9502 (N_9502,N_9491,N_9398);
or U9503 (N_9503,N_9479,N_9426);
nand U9504 (N_9504,N_9411,N_9482);
or U9505 (N_9505,N_9419,N_9401);
or U9506 (N_9506,N_9464,N_9446);
and U9507 (N_9507,N_9433,N_9461);
or U9508 (N_9508,N_9448,N_9386);
nand U9509 (N_9509,N_9463,N_9472);
nor U9510 (N_9510,N_9412,N_9495);
nand U9511 (N_9511,N_9499,N_9438);
nor U9512 (N_9512,N_9470,N_9467);
or U9513 (N_9513,N_9441,N_9395);
or U9514 (N_9514,N_9408,N_9418);
nor U9515 (N_9515,N_9428,N_9442);
or U9516 (N_9516,N_9403,N_9431);
nand U9517 (N_9517,N_9407,N_9417);
or U9518 (N_9518,N_9415,N_9493);
xnor U9519 (N_9519,N_9390,N_9484);
nand U9520 (N_9520,N_9459,N_9424);
and U9521 (N_9521,N_9432,N_9468);
and U9522 (N_9522,N_9447,N_9382);
or U9523 (N_9523,N_9496,N_9489);
or U9524 (N_9524,N_9425,N_9399);
xor U9525 (N_9525,N_9477,N_9492);
nor U9526 (N_9526,N_9423,N_9490);
and U9527 (N_9527,N_9466,N_9420);
or U9528 (N_9528,N_9487,N_9400);
xor U9529 (N_9529,N_9465,N_9460);
or U9530 (N_9530,N_9430,N_9485);
and U9531 (N_9531,N_9391,N_9437);
and U9532 (N_9532,N_9486,N_9427);
xor U9533 (N_9533,N_9384,N_9440);
nand U9534 (N_9534,N_9422,N_9443);
xor U9535 (N_9535,N_9421,N_9483);
nand U9536 (N_9536,N_9455,N_9436);
xnor U9537 (N_9537,N_9381,N_9388);
nand U9538 (N_9538,N_9473,N_9454);
or U9539 (N_9539,N_9383,N_9409);
or U9540 (N_9540,N_9457,N_9379);
nand U9541 (N_9541,N_9396,N_9378);
or U9542 (N_9542,N_9474,N_9476);
or U9543 (N_9543,N_9416,N_9404);
nand U9544 (N_9544,N_9402,N_9380);
xnor U9545 (N_9545,N_9445,N_9456);
or U9546 (N_9546,N_9452,N_9451);
or U9547 (N_9547,N_9449,N_9385);
xnor U9548 (N_9548,N_9429,N_9444);
and U9549 (N_9549,N_9406,N_9387);
nand U9550 (N_9550,N_9462,N_9494);
nand U9551 (N_9551,N_9453,N_9439);
xor U9552 (N_9552,N_9393,N_9414);
or U9553 (N_9553,N_9389,N_9413);
or U9554 (N_9554,N_9394,N_9481);
nor U9555 (N_9555,N_9498,N_9376);
and U9556 (N_9556,N_9488,N_9471);
or U9557 (N_9557,N_9410,N_9375);
nor U9558 (N_9558,N_9497,N_9397);
nor U9559 (N_9559,N_9469,N_9434);
or U9560 (N_9560,N_9435,N_9458);
xor U9561 (N_9561,N_9475,N_9480);
or U9562 (N_9562,N_9392,N_9432);
xor U9563 (N_9563,N_9418,N_9462);
xor U9564 (N_9564,N_9438,N_9426);
or U9565 (N_9565,N_9402,N_9475);
nor U9566 (N_9566,N_9493,N_9382);
and U9567 (N_9567,N_9384,N_9472);
xnor U9568 (N_9568,N_9404,N_9405);
nand U9569 (N_9569,N_9477,N_9425);
xnor U9570 (N_9570,N_9445,N_9479);
nor U9571 (N_9571,N_9412,N_9463);
nand U9572 (N_9572,N_9409,N_9431);
nand U9573 (N_9573,N_9472,N_9446);
nor U9574 (N_9574,N_9394,N_9430);
or U9575 (N_9575,N_9447,N_9490);
and U9576 (N_9576,N_9484,N_9465);
nor U9577 (N_9577,N_9494,N_9386);
xnor U9578 (N_9578,N_9438,N_9481);
nor U9579 (N_9579,N_9412,N_9413);
nor U9580 (N_9580,N_9430,N_9467);
nand U9581 (N_9581,N_9428,N_9380);
xor U9582 (N_9582,N_9407,N_9379);
and U9583 (N_9583,N_9409,N_9435);
or U9584 (N_9584,N_9461,N_9411);
nand U9585 (N_9585,N_9451,N_9405);
or U9586 (N_9586,N_9438,N_9455);
xor U9587 (N_9587,N_9464,N_9499);
nor U9588 (N_9588,N_9462,N_9391);
and U9589 (N_9589,N_9438,N_9474);
xor U9590 (N_9590,N_9473,N_9394);
or U9591 (N_9591,N_9478,N_9464);
xor U9592 (N_9592,N_9424,N_9422);
nor U9593 (N_9593,N_9409,N_9487);
nor U9594 (N_9594,N_9475,N_9464);
nand U9595 (N_9595,N_9433,N_9420);
and U9596 (N_9596,N_9375,N_9398);
or U9597 (N_9597,N_9485,N_9476);
nand U9598 (N_9598,N_9442,N_9449);
xnor U9599 (N_9599,N_9485,N_9394);
and U9600 (N_9600,N_9485,N_9416);
xor U9601 (N_9601,N_9439,N_9476);
xnor U9602 (N_9602,N_9389,N_9416);
and U9603 (N_9603,N_9426,N_9436);
or U9604 (N_9604,N_9385,N_9390);
and U9605 (N_9605,N_9454,N_9436);
nor U9606 (N_9606,N_9470,N_9428);
xor U9607 (N_9607,N_9439,N_9407);
and U9608 (N_9608,N_9427,N_9399);
or U9609 (N_9609,N_9462,N_9463);
or U9610 (N_9610,N_9495,N_9442);
nand U9611 (N_9611,N_9441,N_9381);
or U9612 (N_9612,N_9430,N_9483);
and U9613 (N_9613,N_9426,N_9396);
or U9614 (N_9614,N_9490,N_9415);
or U9615 (N_9615,N_9403,N_9392);
nand U9616 (N_9616,N_9418,N_9441);
xnor U9617 (N_9617,N_9435,N_9433);
nand U9618 (N_9618,N_9496,N_9484);
nand U9619 (N_9619,N_9385,N_9497);
xor U9620 (N_9620,N_9376,N_9431);
nand U9621 (N_9621,N_9439,N_9464);
and U9622 (N_9622,N_9441,N_9430);
and U9623 (N_9623,N_9416,N_9480);
or U9624 (N_9624,N_9395,N_9387);
nand U9625 (N_9625,N_9602,N_9554);
and U9626 (N_9626,N_9607,N_9574);
nor U9627 (N_9627,N_9611,N_9564);
xor U9628 (N_9628,N_9541,N_9514);
nor U9629 (N_9629,N_9519,N_9580);
or U9630 (N_9630,N_9586,N_9539);
xnor U9631 (N_9631,N_9615,N_9588);
and U9632 (N_9632,N_9618,N_9579);
nor U9633 (N_9633,N_9523,N_9590);
nand U9634 (N_9634,N_9597,N_9581);
nand U9635 (N_9635,N_9507,N_9617);
nand U9636 (N_9636,N_9526,N_9546);
and U9637 (N_9637,N_9533,N_9545);
nor U9638 (N_9638,N_9605,N_9560);
nor U9639 (N_9639,N_9616,N_9622);
nor U9640 (N_9640,N_9510,N_9513);
nor U9641 (N_9641,N_9559,N_9515);
nor U9642 (N_9642,N_9516,N_9522);
xor U9643 (N_9643,N_9595,N_9535);
or U9644 (N_9644,N_9551,N_9601);
or U9645 (N_9645,N_9540,N_9511);
xor U9646 (N_9646,N_9583,N_9571);
nand U9647 (N_9647,N_9585,N_9538);
and U9648 (N_9648,N_9500,N_9592);
or U9649 (N_9649,N_9509,N_9600);
nor U9650 (N_9650,N_9529,N_9548);
nand U9651 (N_9651,N_9598,N_9512);
nor U9652 (N_9652,N_9565,N_9505);
nand U9653 (N_9653,N_9620,N_9502);
or U9654 (N_9654,N_9543,N_9593);
nand U9655 (N_9655,N_9562,N_9596);
and U9656 (N_9656,N_9524,N_9604);
and U9657 (N_9657,N_9623,N_9549);
xnor U9658 (N_9658,N_9504,N_9503);
and U9659 (N_9659,N_9528,N_9619);
and U9660 (N_9660,N_9573,N_9589);
nand U9661 (N_9661,N_9575,N_9603);
nand U9662 (N_9662,N_9578,N_9550);
and U9663 (N_9663,N_9566,N_9558);
nand U9664 (N_9664,N_9572,N_9520);
xnor U9665 (N_9665,N_9576,N_9584);
xor U9666 (N_9666,N_9547,N_9518);
xnor U9667 (N_9667,N_9561,N_9555);
xor U9668 (N_9668,N_9612,N_9501);
nor U9669 (N_9669,N_9613,N_9567);
nand U9670 (N_9670,N_9525,N_9537);
and U9671 (N_9671,N_9563,N_9556);
nor U9672 (N_9672,N_9577,N_9624);
xnor U9673 (N_9673,N_9506,N_9582);
or U9674 (N_9674,N_9599,N_9614);
xnor U9675 (N_9675,N_9536,N_9534);
or U9676 (N_9676,N_9517,N_9591);
xnor U9677 (N_9677,N_9530,N_9557);
xor U9678 (N_9678,N_9569,N_9621);
and U9679 (N_9679,N_9606,N_9570);
nor U9680 (N_9680,N_9544,N_9610);
nand U9681 (N_9681,N_9531,N_9568);
and U9682 (N_9682,N_9532,N_9609);
xor U9683 (N_9683,N_9594,N_9508);
and U9684 (N_9684,N_9542,N_9521);
and U9685 (N_9685,N_9587,N_9608);
or U9686 (N_9686,N_9527,N_9553);
and U9687 (N_9687,N_9552,N_9603);
and U9688 (N_9688,N_9581,N_9554);
xnor U9689 (N_9689,N_9617,N_9545);
xor U9690 (N_9690,N_9607,N_9564);
and U9691 (N_9691,N_9501,N_9594);
xnor U9692 (N_9692,N_9561,N_9529);
nand U9693 (N_9693,N_9604,N_9572);
nor U9694 (N_9694,N_9609,N_9607);
or U9695 (N_9695,N_9504,N_9508);
xnor U9696 (N_9696,N_9587,N_9598);
or U9697 (N_9697,N_9591,N_9624);
nand U9698 (N_9698,N_9544,N_9586);
nor U9699 (N_9699,N_9591,N_9581);
nor U9700 (N_9700,N_9607,N_9514);
and U9701 (N_9701,N_9515,N_9516);
or U9702 (N_9702,N_9603,N_9556);
and U9703 (N_9703,N_9519,N_9583);
xor U9704 (N_9704,N_9544,N_9546);
or U9705 (N_9705,N_9584,N_9561);
or U9706 (N_9706,N_9620,N_9515);
and U9707 (N_9707,N_9593,N_9548);
or U9708 (N_9708,N_9585,N_9542);
or U9709 (N_9709,N_9543,N_9562);
and U9710 (N_9710,N_9533,N_9618);
xnor U9711 (N_9711,N_9608,N_9526);
and U9712 (N_9712,N_9524,N_9575);
or U9713 (N_9713,N_9622,N_9619);
nor U9714 (N_9714,N_9508,N_9550);
nand U9715 (N_9715,N_9559,N_9563);
xnor U9716 (N_9716,N_9542,N_9537);
and U9717 (N_9717,N_9601,N_9573);
nor U9718 (N_9718,N_9540,N_9567);
xnor U9719 (N_9719,N_9567,N_9578);
or U9720 (N_9720,N_9589,N_9539);
and U9721 (N_9721,N_9577,N_9508);
or U9722 (N_9722,N_9512,N_9571);
nor U9723 (N_9723,N_9608,N_9565);
nor U9724 (N_9724,N_9606,N_9562);
nand U9725 (N_9725,N_9612,N_9601);
nor U9726 (N_9726,N_9522,N_9608);
nor U9727 (N_9727,N_9512,N_9595);
and U9728 (N_9728,N_9606,N_9547);
nor U9729 (N_9729,N_9518,N_9525);
and U9730 (N_9730,N_9586,N_9501);
nor U9731 (N_9731,N_9530,N_9542);
xnor U9732 (N_9732,N_9569,N_9584);
nand U9733 (N_9733,N_9563,N_9504);
or U9734 (N_9734,N_9590,N_9510);
xnor U9735 (N_9735,N_9561,N_9607);
or U9736 (N_9736,N_9603,N_9501);
nand U9737 (N_9737,N_9615,N_9550);
nand U9738 (N_9738,N_9602,N_9514);
xor U9739 (N_9739,N_9570,N_9522);
and U9740 (N_9740,N_9542,N_9574);
nand U9741 (N_9741,N_9618,N_9611);
nand U9742 (N_9742,N_9526,N_9564);
nand U9743 (N_9743,N_9580,N_9539);
nor U9744 (N_9744,N_9537,N_9505);
xor U9745 (N_9745,N_9532,N_9578);
nand U9746 (N_9746,N_9531,N_9536);
xor U9747 (N_9747,N_9504,N_9566);
or U9748 (N_9748,N_9560,N_9592);
or U9749 (N_9749,N_9615,N_9612);
or U9750 (N_9750,N_9670,N_9719);
nand U9751 (N_9751,N_9711,N_9728);
xor U9752 (N_9752,N_9646,N_9700);
xnor U9753 (N_9753,N_9674,N_9691);
or U9754 (N_9754,N_9729,N_9673);
nand U9755 (N_9755,N_9648,N_9745);
xor U9756 (N_9756,N_9725,N_9749);
nor U9757 (N_9757,N_9685,N_9692);
and U9758 (N_9758,N_9637,N_9626);
nor U9759 (N_9759,N_9655,N_9718);
xor U9760 (N_9760,N_9676,N_9723);
or U9761 (N_9761,N_9748,N_9667);
xnor U9762 (N_9762,N_9682,N_9690);
and U9763 (N_9763,N_9644,N_9726);
xnor U9764 (N_9764,N_9689,N_9703);
or U9765 (N_9765,N_9661,N_9641);
xnor U9766 (N_9766,N_9686,N_9742);
nor U9767 (N_9767,N_9628,N_9656);
or U9768 (N_9768,N_9734,N_9629);
nand U9769 (N_9769,N_9645,N_9634);
xor U9770 (N_9770,N_9654,N_9638);
or U9771 (N_9771,N_9647,N_9735);
and U9772 (N_9772,N_9704,N_9677);
nand U9773 (N_9773,N_9712,N_9705);
xor U9774 (N_9774,N_9747,N_9732);
xnor U9775 (N_9775,N_9636,N_9649);
or U9776 (N_9776,N_9695,N_9630);
and U9777 (N_9777,N_9720,N_9631);
xnor U9778 (N_9778,N_9662,N_9721);
nand U9779 (N_9779,N_9639,N_9651);
nor U9780 (N_9780,N_9668,N_9696);
and U9781 (N_9781,N_9743,N_9632);
nor U9782 (N_9782,N_9627,N_9730);
and U9783 (N_9783,N_9675,N_9643);
or U9784 (N_9784,N_9706,N_9678);
or U9785 (N_9785,N_9681,N_9642);
nand U9786 (N_9786,N_9664,N_9625);
and U9787 (N_9787,N_9741,N_9698);
nor U9788 (N_9788,N_9640,N_9717);
nand U9789 (N_9789,N_9727,N_9633);
nand U9790 (N_9790,N_9739,N_9709);
and U9791 (N_9791,N_9650,N_9671);
nand U9792 (N_9792,N_9659,N_9669);
nand U9793 (N_9793,N_9710,N_9744);
xor U9794 (N_9794,N_9724,N_9679);
nand U9795 (N_9795,N_9699,N_9716);
or U9796 (N_9796,N_9666,N_9713);
and U9797 (N_9797,N_9684,N_9714);
xnor U9798 (N_9798,N_9702,N_9693);
and U9799 (N_9799,N_9708,N_9733);
xor U9800 (N_9800,N_9731,N_9660);
nand U9801 (N_9801,N_9683,N_9736);
and U9802 (N_9802,N_9657,N_9665);
nand U9803 (N_9803,N_9697,N_9694);
nor U9804 (N_9804,N_9738,N_9707);
xor U9805 (N_9805,N_9635,N_9715);
nor U9806 (N_9806,N_9653,N_9672);
xor U9807 (N_9807,N_9722,N_9687);
xor U9808 (N_9808,N_9663,N_9688);
and U9809 (N_9809,N_9680,N_9701);
and U9810 (N_9810,N_9740,N_9737);
nor U9811 (N_9811,N_9746,N_9658);
nand U9812 (N_9812,N_9652,N_9705);
nor U9813 (N_9813,N_9630,N_9694);
nand U9814 (N_9814,N_9741,N_9694);
xnor U9815 (N_9815,N_9715,N_9744);
nor U9816 (N_9816,N_9706,N_9681);
nand U9817 (N_9817,N_9701,N_9632);
xor U9818 (N_9818,N_9632,N_9716);
or U9819 (N_9819,N_9661,N_9657);
or U9820 (N_9820,N_9649,N_9645);
nand U9821 (N_9821,N_9722,N_9720);
xnor U9822 (N_9822,N_9625,N_9739);
or U9823 (N_9823,N_9681,N_9669);
and U9824 (N_9824,N_9698,N_9715);
xor U9825 (N_9825,N_9699,N_9698);
and U9826 (N_9826,N_9633,N_9656);
xor U9827 (N_9827,N_9691,N_9646);
nor U9828 (N_9828,N_9632,N_9731);
and U9829 (N_9829,N_9638,N_9728);
xor U9830 (N_9830,N_9637,N_9715);
nand U9831 (N_9831,N_9678,N_9743);
or U9832 (N_9832,N_9709,N_9701);
or U9833 (N_9833,N_9742,N_9741);
xnor U9834 (N_9834,N_9678,N_9659);
and U9835 (N_9835,N_9719,N_9675);
nand U9836 (N_9836,N_9700,N_9668);
nand U9837 (N_9837,N_9661,N_9745);
and U9838 (N_9838,N_9639,N_9734);
or U9839 (N_9839,N_9659,N_9689);
xor U9840 (N_9840,N_9746,N_9650);
and U9841 (N_9841,N_9724,N_9714);
or U9842 (N_9842,N_9693,N_9747);
xnor U9843 (N_9843,N_9701,N_9691);
nand U9844 (N_9844,N_9687,N_9649);
and U9845 (N_9845,N_9688,N_9668);
nor U9846 (N_9846,N_9672,N_9633);
or U9847 (N_9847,N_9688,N_9666);
nor U9848 (N_9848,N_9709,N_9717);
and U9849 (N_9849,N_9665,N_9628);
xor U9850 (N_9850,N_9700,N_9661);
xor U9851 (N_9851,N_9699,N_9710);
nand U9852 (N_9852,N_9724,N_9633);
nand U9853 (N_9853,N_9707,N_9665);
nor U9854 (N_9854,N_9723,N_9719);
nor U9855 (N_9855,N_9691,N_9707);
nor U9856 (N_9856,N_9649,N_9700);
xnor U9857 (N_9857,N_9646,N_9631);
nand U9858 (N_9858,N_9705,N_9673);
and U9859 (N_9859,N_9703,N_9677);
nor U9860 (N_9860,N_9685,N_9743);
or U9861 (N_9861,N_9711,N_9651);
or U9862 (N_9862,N_9647,N_9679);
and U9863 (N_9863,N_9697,N_9687);
xnor U9864 (N_9864,N_9740,N_9689);
nand U9865 (N_9865,N_9673,N_9663);
and U9866 (N_9866,N_9721,N_9726);
and U9867 (N_9867,N_9734,N_9679);
or U9868 (N_9868,N_9727,N_9724);
xnor U9869 (N_9869,N_9671,N_9708);
nand U9870 (N_9870,N_9681,N_9639);
and U9871 (N_9871,N_9658,N_9685);
nand U9872 (N_9872,N_9698,N_9710);
and U9873 (N_9873,N_9672,N_9701);
or U9874 (N_9874,N_9661,N_9645);
nor U9875 (N_9875,N_9778,N_9855);
nand U9876 (N_9876,N_9753,N_9808);
or U9877 (N_9877,N_9870,N_9787);
and U9878 (N_9878,N_9827,N_9843);
xnor U9879 (N_9879,N_9750,N_9846);
nor U9880 (N_9880,N_9790,N_9780);
or U9881 (N_9881,N_9776,N_9854);
nand U9882 (N_9882,N_9819,N_9844);
nor U9883 (N_9883,N_9794,N_9793);
nand U9884 (N_9884,N_9848,N_9766);
or U9885 (N_9885,N_9828,N_9812);
nand U9886 (N_9886,N_9871,N_9770);
nor U9887 (N_9887,N_9864,N_9850);
xor U9888 (N_9888,N_9851,N_9837);
or U9889 (N_9889,N_9803,N_9752);
xor U9890 (N_9890,N_9802,N_9866);
nor U9891 (N_9891,N_9810,N_9796);
or U9892 (N_9892,N_9811,N_9852);
or U9893 (N_9893,N_9774,N_9777);
or U9894 (N_9894,N_9772,N_9860);
and U9895 (N_9895,N_9757,N_9818);
or U9896 (N_9896,N_9761,N_9861);
nand U9897 (N_9897,N_9763,N_9813);
or U9898 (N_9898,N_9862,N_9849);
xor U9899 (N_9899,N_9824,N_9820);
nand U9900 (N_9900,N_9775,N_9853);
xor U9901 (N_9901,N_9773,N_9797);
and U9902 (N_9902,N_9756,N_9814);
or U9903 (N_9903,N_9807,N_9779);
and U9904 (N_9904,N_9798,N_9825);
or U9905 (N_9905,N_9783,N_9832);
nand U9906 (N_9906,N_9792,N_9865);
and U9907 (N_9907,N_9841,N_9872);
and U9908 (N_9908,N_9838,N_9868);
nand U9909 (N_9909,N_9815,N_9826);
nor U9910 (N_9910,N_9816,N_9830);
or U9911 (N_9911,N_9833,N_9799);
nor U9912 (N_9912,N_9869,N_9823);
and U9913 (N_9913,N_9831,N_9835);
xor U9914 (N_9914,N_9769,N_9751);
xnor U9915 (N_9915,N_9804,N_9767);
nor U9916 (N_9916,N_9806,N_9755);
and U9917 (N_9917,N_9847,N_9805);
nor U9918 (N_9918,N_9782,N_9836);
nor U9919 (N_9919,N_9781,N_9834);
and U9920 (N_9920,N_9840,N_9842);
and U9921 (N_9921,N_9859,N_9829);
xnor U9922 (N_9922,N_9768,N_9801);
xor U9923 (N_9923,N_9765,N_9759);
and U9924 (N_9924,N_9788,N_9786);
and U9925 (N_9925,N_9856,N_9817);
and U9926 (N_9926,N_9845,N_9785);
nor U9927 (N_9927,N_9789,N_9867);
xor U9928 (N_9928,N_9873,N_9874);
nor U9929 (N_9929,N_9762,N_9858);
nor U9930 (N_9930,N_9800,N_9771);
or U9931 (N_9931,N_9839,N_9784);
and U9932 (N_9932,N_9760,N_9795);
nor U9933 (N_9933,N_9754,N_9791);
xnor U9934 (N_9934,N_9863,N_9821);
and U9935 (N_9935,N_9764,N_9857);
nor U9936 (N_9936,N_9809,N_9822);
xor U9937 (N_9937,N_9758,N_9862);
xor U9938 (N_9938,N_9850,N_9787);
nand U9939 (N_9939,N_9758,N_9751);
nand U9940 (N_9940,N_9761,N_9858);
nand U9941 (N_9941,N_9845,N_9752);
xor U9942 (N_9942,N_9780,N_9796);
nor U9943 (N_9943,N_9798,N_9807);
nand U9944 (N_9944,N_9829,N_9797);
nand U9945 (N_9945,N_9846,N_9796);
and U9946 (N_9946,N_9810,N_9753);
xnor U9947 (N_9947,N_9823,N_9790);
nand U9948 (N_9948,N_9840,N_9760);
xor U9949 (N_9949,N_9871,N_9846);
nand U9950 (N_9950,N_9836,N_9803);
or U9951 (N_9951,N_9765,N_9818);
nand U9952 (N_9952,N_9862,N_9848);
nor U9953 (N_9953,N_9789,N_9791);
nand U9954 (N_9954,N_9863,N_9837);
or U9955 (N_9955,N_9860,N_9804);
and U9956 (N_9956,N_9863,N_9826);
or U9957 (N_9957,N_9793,N_9800);
and U9958 (N_9958,N_9788,N_9794);
or U9959 (N_9959,N_9868,N_9798);
nor U9960 (N_9960,N_9823,N_9762);
and U9961 (N_9961,N_9774,N_9808);
and U9962 (N_9962,N_9862,N_9763);
or U9963 (N_9963,N_9803,N_9773);
or U9964 (N_9964,N_9841,N_9796);
nand U9965 (N_9965,N_9763,N_9833);
nand U9966 (N_9966,N_9874,N_9839);
nand U9967 (N_9967,N_9791,N_9837);
nor U9968 (N_9968,N_9816,N_9801);
xnor U9969 (N_9969,N_9835,N_9759);
nor U9970 (N_9970,N_9788,N_9813);
xor U9971 (N_9971,N_9871,N_9840);
and U9972 (N_9972,N_9866,N_9779);
or U9973 (N_9973,N_9815,N_9824);
and U9974 (N_9974,N_9771,N_9797);
and U9975 (N_9975,N_9770,N_9799);
or U9976 (N_9976,N_9821,N_9837);
nand U9977 (N_9977,N_9815,N_9850);
nand U9978 (N_9978,N_9802,N_9783);
and U9979 (N_9979,N_9782,N_9844);
xnor U9980 (N_9980,N_9798,N_9821);
and U9981 (N_9981,N_9809,N_9873);
nor U9982 (N_9982,N_9819,N_9870);
and U9983 (N_9983,N_9872,N_9859);
and U9984 (N_9984,N_9829,N_9870);
xor U9985 (N_9985,N_9859,N_9849);
and U9986 (N_9986,N_9756,N_9791);
or U9987 (N_9987,N_9854,N_9837);
and U9988 (N_9988,N_9800,N_9769);
xor U9989 (N_9989,N_9751,N_9849);
and U9990 (N_9990,N_9867,N_9857);
nor U9991 (N_9991,N_9793,N_9855);
xor U9992 (N_9992,N_9856,N_9827);
or U9993 (N_9993,N_9826,N_9795);
and U9994 (N_9994,N_9827,N_9755);
nor U9995 (N_9995,N_9770,N_9794);
nand U9996 (N_9996,N_9759,N_9840);
xor U9997 (N_9997,N_9794,N_9858);
nor U9998 (N_9998,N_9755,N_9844);
nand U9999 (N_9999,N_9776,N_9833);
nor U10000 (N_10000,N_9903,N_9901);
and U10001 (N_10001,N_9985,N_9922);
nor U10002 (N_10002,N_9937,N_9958);
and U10003 (N_10003,N_9947,N_9989);
or U10004 (N_10004,N_9991,N_9929);
nand U10005 (N_10005,N_9880,N_9876);
xor U10006 (N_10006,N_9900,N_9939);
and U10007 (N_10007,N_9983,N_9952);
or U10008 (N_10008,N_9894,N_9918);
nor U10009 (N_10009,N_9964,N_9980);
xor U10010 (N_10010,N_9878,N_9954);
xor U10011 (N_10011,N_9884,N_9956);
xnor U10012 (N_10012,N_9938,N_9946);
xnor U10013 (N_10013,N_9959,N_9877);
xor U10014 (N_10014,N_9967,N_9889);
nand U10015 (N_10015,N_9935,N_9982);
nor U10016 (N_10016,N_9988,N_9925);
xor U10017 (N_10017,N_9999,N_9986);
nor U10018 (N_10018,N_9914,N_9905);
or U10019 (N_10019,N_9981,N_9969);
nand U10020 (N_10020,N_9893,N_9879);
or U10021 (N_10021,N_9927,N_9971);
or U10022 (N_10022,N_9906,N_9926);
and U10023 (N_10023,N_9984,N_9978);
nand U10024 (N_10024,N_9992,N_9943);
or U10025 (N_10025,N_9966,N_9902);
or U10026 (N_10026,N_9963,N_9979);
and U10027 (N_10027,N_9931,N_9998);
xor U10028 (N_10028,N_9883,N_9917);
xor U10029 (N_10029,N_9949,N_9933);
and U10030 (N_10030,N_9936,N_9891);
or U10031 (N_10031,N_9923,N_9888);
xor U10032 (N_10032,N_9934,N_9951);
xor U10033 (N_10033,N_9990,N_9895);
and U10034 (N_10034,N_9928,N_9910);
or U10035 (N_10035,N_9955,N_9962);
or U10036 (N_10036,N_9950,N_9975);
xor U10037 (N_10037,N_9898,N_9875);
xor U10038 (N_10038,N_9976,N_9973);
or U10039 (N_10039,N_9913,N_9945);
and U10040 (N_10040,N_9886,N_9960);
nand U10041 (N_10041,N_9920,N_9953);
or U10042 (N_10042,N_9961,N_9899);
or U10043 (N_10043,N_9941,N_9882);
xnor U10044 (N_10044,N_9885,N_9957);
nor U10045 (N_10045,N_9994,N_9965);
and U10046 (N_10046,N_9897,N_9993);
xor U10047 (N_10047,N_9909,N_9904);
xnor U10048 (N_10048,N_9921,N_9974);
nor U10049 (N_10049,N_9997,N_9907);
nand U10050 (N_10050,N_9987,N_9996);
and U10051 (N_10051,N_9919,N_9944);
and U10052 (N_10052,N_9887,N_9970);
and U10053 (N_10053,N_9890,N_9916);
nor U10054 (N_10054,N_9915,N_9972);
or U10055 (N_10055,N_9942,N_9892);
or U10056 (N_10056,N_9912,N_9896);
nor U10057 (N_10057,N_9911,N_9924);
nand U10058 (N_10058,N_9968,N_9995);
and U10059 (N_10059,N_9908,N_9948);
or U10060 (N_10060,N_9977,N_9932);
and U10061 (N_10061,N_9930,N_9881);
xnor U10062 (N_10062,N_9940,N_9909);
or U10063 (N_10063,N_9999,N_9943);
nand U10064 (N_10064,N_9997,N_9989);
nand U10065 (N_10065,N_9926,N_9999);
and U10066 (N_10066,N_9951,N_9947);
and U10067 (N_10067,N_9894,N_9916);
and U10068 (N_10068,N_9945,N_9978);
xnor U10069 (N_10069,N_9910,N_9907);
nand U10070 (N_10070,N_9968,N_9942);
or U10071 (N_10071,N_9882,N_9923);
or U10072 (N_10072,N_9950,N_9934);
and U10073 (N_10073,N_9953,N_9966);
nand U10074 (N_10074,N_9944,N_9974);
or U10075 (N_10075,N_9942,N_9954);
or U10076 (N_10076,N_9974,N_9879);
nand U10077 (N_10077,N_9978,N_9897);
nand U10078 (N_10078,N_9902,N_9988);
nand U10079 (N_10079,N_9931,N_9962);
nand U10080 (N_10080,N_9939,N_9998);
nand U10081 (N_10081,N_9899,N_9932);
xor U10082 (N_10082,N_9879,N_9942);
or U10083 (N_10083,N_9990,N_9890);
xnor U10084 (N_10084,N_9950,N_9994);
and U10085 (N_10085,N_9996,N_9906);
and U10086 (N_10086,N_9972,N_9987);
nand U10087 (N_10087,N_9931,N_9984);
nor U10088 (N_10088,N_9907,N_9995);
and U10089 (N_10089,N_9987,N_9974);
nand U10090 (N_10090,N_9960,N_9923);
or U10091 (N_10091,N_9922,N_9951);
nor U10092 (N_10092,N_9976,N_9926);
nor U10093 (N_10093,N_9980,N_9968);
nor U10094 (N_10094,N_9966,N_9884);
nand U10095 (N_10095,N_9965,N_9931);
nor U10096 (N_10096,N_9882,N_9970);
and U10097 (N_10097,N_9991,N_9878);
nor U10098 (N_10098,N_9922,N_9971);
nand U10099 (N_10099,N_9960,N_9978);
nand U10100 (N_10100,N_9991,N_9903);
or U10101 (N_10101,N_9925,N_9956);
xnor U10102 (N_10102,N_9918,N_9980);
nand U10103 (N_10103,N_9951,N_9929);
nor U10104 (N_10104,N_9990,N_9903);
xnor U10105 (N_10105,N_9920,N_9963);
nand U10106 (N_10106,N_9882,N_9920);
nand U10107 (N_10107,N_9905,N_9884);
and U10108 (N_10108,N_9903,N_9913);
and U10109 (N_10109,N_9962,N_9894);
nand U10110 (N_10110,N_9900,N_9960);
nand U10111 (N_10111,N_9977,N_9968);
xor U10112 (N_10112,N_9956,N_9900);
nor U10113 (N_10113,N_9952,N_9937);
or U10114 (N_10114,N_9900,N_9935);
nor U10115 (N_10115,N_9973,N_9930);
xnor U10116 (N_10116,N_9944,N_9895);
xnor U10117 (N_10117,N_9924,N_9934);
and U10118 (N_10118,N_9895,N_9902);
nand U10119 (N_10119,N_9963,N_9913);
and U10120 (N_10120,N_9997,N_9903);
or U10121 (N_10121,N_9971,N_9880);
nand U10122 (N_10122,N_9892,N_9895);
xnor U10123 (N_10123,N_9943,N_9903);
nor U10124 (N_10124,N_9887,N_9879);
and U10125 (N_10125,N_10102,N_10109);
and U10126 (N_10126,N_10092,N_10089);
xnor U10127 (N_10127,N_10017,N_10020);
nor U10128 (N_10128,N_10121,N_10096);
nand U10129 (N_10129,N_10064,N_10103);
and U10130 (N_10130,N_10083,N_10033);
xor U10131 (N_10131,N_10050,N_10044);
or U10132 (N_10132,N_10015,N_10122);
xor U10133 (N_10133,N_10008,N_10084);
and U10134 (N_10134,N_10081,N_10013);
nor U10135 (N_10135,N_10032,N_10000);
and U10136 (N_10136,N_10009,N_10024);
xor U10137 (N_10137,N_10088,N_10077);
xnor U10138 (N_10138,N_10075,N_10073);
xor U10139 (N_10139,N_10060,N_10021);
xor U10140 (N_10140,N_10004,N_10112);
xnor U10141 (N_10141,N_10001,N_10057);
nand U10142 (N_10142,N_10104,N_10022);
or U10143 (N_10143,N_10026,N_10115);
or U10144 (N_10144,N_10035,N_10068);
nor U10145 (N_10145,N_10038,N_10119);
or U10146 (N_10146,N_10124,N_10019);
xor U10147 (N_10147,N_10036,N_10074);
nor U10148 (N_10148,N_10100,N_10037);
nor U10149 (N_10149,N_10046,N_10094);
or U10150 (N_10150,N_10011,N_10051);
and U10151 (N_10151,N_10018,N_10114);
or U10152 (N_10152,N_10093,N_10101);
or U10153 (N_10153,N_10085,N_10106);
or U10154 (N_10154,N_10113,N_10117);
nor U10155 (N_10155,N_10052,N_10025);
or U10156 (N_10156,N_10120,N_10002);
or U10157 (N_10157,N_10076,N_10043);
or U10158 (N_10158,N_10058,N_10039);
or U10159 (N_10159,N_10099,N_10080);
and U10160 (N_10160,N_10056,N_10082);
nor U10161 (N_10161,N_10027,N_10069);
or U10162 (N_10162,N_10014,N_10123);
and U10163 (N_10163,N_10086,N_10111);
xor U10164 (N_10164,N_10007,N_10067);
and U10165 (N_10165,N_10097,N_10091);
and U10166 (N_10166,N_10010,N_10053);
nor U10167 (N_10167,N_10062,N_10107);
nand U10168 (N_10168,N_10116,N_10048);
nor U10169 (N_10169,N_10079,N_10071);
nand U10170 (N_10170,N_10059,N_10005);
nor U10171 (N_10171,N_10090,N_10098);
nor U10172 (N_10172,N_10047,N_10108);
or U10173 (N_10173,N_10054,N_10012);
nor U10174 (N_10174,N_10028,N_10061);
or U10175 (N_10175,N_10066,N_10105);
and U10176 (N_10176,N_10003,N_10029);
nor U10177 (N_10177,N_10070,N_10023);
nor U10178 (N_10178,N_10110,N_10078);
nand U10179 (N_10179,N_10031,N_10030);
or U10180 (N_10180,N_10042,N_10072);
and U10181 (N_10181,N_10055,N_10034);
nor U10182 (N_10182,N_10045,N_10118);
nor U10183 (N_10183,N_10006,N_10065);
or U10184 (N_10184,N_10040,N_10063);
xor U10185 (N_10185,N_10016,N_10041);
and U10186 (N_10186,N_10095,N_10087);
and U10187 (N_10187,N_10049,N_10044);
xnor U10188 (N_10188,N_10086,N_10041);
or U10189 (N_10189,N_10104,N_10082);
nor U10190 (N_10190,N_10095,N_10122);
or U10191 (N_10191,N_10011,N_10042);
xor U10192 (N_10192,N_10093,N_10008);
nand U10193 (N_10193,N_10082,N_10018);
and U10194 (N_10194,N_10077,N_10100);
or U10195 (N_10195,N_10107,N_10111);
and U10196 (N_10196,N_10086,N_10099);
nor U10197 (N_10197,N_10009,N_10036);
or U10198 (N_10198,N_10063,N_10046);
and U10199 (N_10199,N_10045,N_10076);
or U10200 (N_10200,N_10085,N_10077);
nor U10201 (N_10201,N_10007,N_10075);
xnor U10202 (N_10202,N_10112,N_10099);
or U10203 (N_10203,N_10027,N_10113);
or U10204 (N_10204,N_10049,N_10081);
xnor U10205 (N_10205,N_10049,N_10104);
xor U10206 (N_10206,N_10073,N_10010);
nand U10207 (N_10207,N_10031,N_10057);
and U10208 (N_10208,N_10026,N_10030);
nor U10209 (N_10209,N_10101,N_10104);
or U10210 (N_10210,N_10082,N_10118);
or U10211 (N_10211,N_10049,N_10023);
and U10212 (N_10212,N_10014,N_10075);
and U10213 (N_10213,N_10111,N_10092);
xnor U10214 (N_10214,N_10022,N_10106);
and U10215 (N_10215,N_10086,N_10014);
xnor U10216 (N_10216,N_10027,N_10117);
nand U10217 (N_10217,N_10005,N_10083);
xnor U10218 (N_10218,N_10108,N_10040);
and U10219 (N_10219,N_10019,N_10020);
or U10220 (N_10220,N_10101,N_10088);
or U10221 (N_10221,N_10022,N_10070);
nor U10222 (N_10222,N_10117,N_10102);
and U10223 (N_10223,N_10004,N_10025);
or U10224 (N_10224,N_10099,N_10076);
or U10225 (N_10225,N_10055,N_10098);
and U10226 (N_10226,N_10027,N_10006);
or U10227 (N_10227,N_10035,N_10071);
and U10228 (N_10228,N_10117,N_10119);
or U10229 (N_10229,N_10123,N_10066);
and U10230 (N_10230,N_10104,N_10083);
and U10231 (N_10231,N_10058,N_10022);
or U10232 (N_10232,N_10104,N_10053);
or U10233 (N_10233,N_10070,N_10074);
or U10234 (N_10234,N_10093,N_10099);
or U10235 (N_10235,N_10051,N_10082);
xor U10236 (N_10236,N_10123,N_10012);
nand U10237 (N_10237,N_10065,N_10108);
nand U10238 (N_10238,N_10118,N_10074);
xor U10239 (N_10239,N_10013,N_10049);
or U10240 (N_10240,N_10019,N_10082);
and U10241 (N_10241,N_10087,N_10061);
nor U10242 (N_10242,N_10061,N_10085);
and U10243 (N_10243,N_10079,N_10074);
and U10244 (N_10244,N_10050,N_10114);
nor U10245 (N_10245,N_10068,N_10019);
xor U10246 (N_10246,N_10001,N_10086);
xor U10247 (N_10247,N_10115,N_10054);
xor U10248 (N_10248,N_10001,N_10112);
nand U10249 (N_10249,N_10066,N_10015);
xnor U10250 (N_10250,N_10171,N_10149);
and U10251 (N_10251,N_10207,N_10221);
and U10252 (N_10252,N_10215,N_10218);
and U10253 (N_10253,N_10142,N_10174);
and U10254 (N_10254,N_10182,N_10212);
xnor U10255 (N_10255,N_10223,N_10187);
nand U10256 (N_10256,N_10128,N_10132);
and U10257 (N_10257,N_10194,N_10137);
xnor U10258 (N_10258,N_10166,N_10247);
nand U10259 (N_10259,N_10170,N_10211);
xnor U10260 (N_10260,N_10203,N_10147);
xor U10261 (N_10261,N_10244,N_10206);
and U10262 (N_10262,N_10176,N_10130);
xnor U10263 (N_10263,N_10185,N_10159);
or U10264 (N_10264,N_10191,N_10144);
nand U10265 (N_10265,N_10175,N_10129);
nor U10266 (N_10266,N_10200,N_10158);
nand U10267 (N_10267,N_10131,N_10180);
or U10268 (N_10268,N_10145,N_10195);
nand U10269 (N_10269,N_10240,N_10161);
and U10270 (N_10270,N_10225,N_10140);
nand U10271 (N_10271,N_10226,N_10165);
and U10272 (N_10272,N_10192,N_10245);
nand U10273 (N_10273,N_10246,N_10242);
and U10274 (N_10274,N_10167,N_10169);
xor U10275 (N_10275,N_10133,N_10188);
nor U10276 (N_10276,N_10154,N_10143);
and U10277 (N_10277,N_10249,N_10205);
or U10278 (N_10278,N_10155,N_10236);
nor U10279 (N_10279,N_10231,N_10190);
and U10280 (N_10280,N_10216,N_10135);
nor U10281 (N_10281,N_10217,N_10163);
nor U10282 (N_10282,N_10184,N_10141);
xor U10283 (N_10283,N_10224,N_10153);
nor U10284 (N_10284,N_10199,N_10173);
nand U10285 (N_10285,N_10222,N_10196);
xnor U10286 (N_10286,N_10151,N_10220);
xnor U10287 (N_10287,N_10235,N_10152);
and U10288 (N_10288,N_10227,N_10148);
xnor U10289 (N_10289,N_10134,N_10229);
nand U10290 (N_10290,N_10214,N_10127);
xor U10291 (N_10291,N_10183,N_10150);
nand U10292 (N_10292,N_10208,N_10233);
and U10293 (N_10293,N_10179,N_10138);
and U10294 (N_10294,N_10202,N_10238);
or U10295 (N_10295,N_10232,N_10160);
nand U10296 (N_10296,N_10228,N_10139);
nor U10297 (N_10297,N_10146,N_10209);
and U10298 (N_10298,N_10198,N_10237);
nand U10299 (N_10299,N_10243,N_10125);
nor U10300 (N_10300,N_10234,N_10201);
and U10301 (N_10301,N_10186,N_10157);
nor U10302 (N_10302,N_10239,N_10197);
and U10303 (N_10303,N_10136,N_10248);
or U10304 (N_10304,N_10230,N_10181);
xnor U10305 (N_10305,N_10189,N_10168);
and U10306 (N_10306,N_10241,N_10162);
and U10307 (N_10307,N_10210,N_10178);
and U10308 (N_10308,N_10204,N_10177);
and U10309 (N_10309,N_10213,N_10219);
and U10310 (N_10310,N_10164,N_10193);
nor U10311 (N_10311,N_10156,N_10126);
nand U10312 (N_10312,N_10172,N_10236);
nor U10313 (N_10313,N_10158,N_10184);
or U10314 (N_10314,N_10157,N_10242);
nand U10315 (N_10315,N_10244,N_10136);
and U10316 (N_10316,N_10143,N_10150);
nand U10317 (N_10317,N_10126,N_10177);
and U10318 (N_10318,N_10183,N_10223);
or U10319 (N_10319,N_10185,N_10182);
xnor U10320 (N_10320,N_10239,N_10190);
xor U10321 (N_10321,N_10207,N_10194);
xor U10322 (N_10322,N_10171,N_10146);
xnor U10323 (N_10323,N_10172,N_10221);
xor U10324 (N_10324,N_10239,N_10138);
nand U10325 (N_10325,N_10235,N_10139);
nor U10326 (N_10326,N_10234,N_10196);
and U10327 (N_10327,N_10219,N_10186);
xnor U10328 (N_10328,N_10135,N_10201);
xnor U10329 (N_10329,N_10182,N_10220);
xnor U10330 (N_10330,N_10210,N_10163);
nor U10331 (N_10331,N_10223,N_10201);
or U10332 (N_10332,N_10225,N_10239);
nor U10333 (N_10333,N_10236,N_10186);
nand U10334 (N_10334,N_10209,N_10184);
nand U10335 (N_10335,N_10199,N_10236);
nor U10336 (N_10336,N_10151,N_10246);
or U10337 (N_10337,N_10184,N_10165);
and U10338 (N_10338,N_10234,N_10185);
and U10339 (N_10339,N_10224,N_10206);
and U10340 (N_10340,N_10180,N_10177);
and U10341 (N_10341,N_10202,N_10242);
nor U10342 (N_10342,N_10189,N_10191);
and U10343 (N_10343,N_10246,N_10191);
nor U10344 (N_10344,N_10158,N_10211);
nand U10345 (N_10345,N_10186,N_10187);
and U10346 (N_10346,N_10232,N_10222);
and U10347 (N_10347,N_10190,N_10220);
nor U10348 (N_10348,N_10216,N_10213);
and U10349 (N_10349,N_10197,N_10151);
nor U10350 (N_10350,N_10229,N_10182);
xor U10351 (N_10351,N_10234,N_10131);
nand U10352 (N_10352,N_10137,N_10229);
nand U10353 (N_10353,N_10205,N_10203);
nor U10354 (N_10354,N_10153,N_10184);
or U10355 (N_10355,N_10125,N_10128);
and U10356 (N_10356,N_10128,N_10159);
or U10357 (N_10357,N_10241,N_10220);
or U10358 (N_10358,N_10150,N_10152);
and U10359 (N_10359,N_10170,N_10155);
xnor U10360 (N_10360,N_10171,N_10136);
or U10361 (N_10361,N_10187,N_10234);
nand U10362 (N_10362,N_10184,N_10227);
and U10363 (N_10363,N_10214,N_10155);
nand U10364 (N_10364,N_10154,N_10195);
nand U10365 (N_10365,N_10174,N_10248);
or U10366 (N_10366,N_10237,N_10206);
and U10367 (N_10367,N_10235,N_10241);
or U10368 (N_10368,N_10170,N_10152);
xnor U10369 (N_10369,N_10195,N_10156);
or U10370 (N_10370,N_10142,N_10195);
nand U10371 (N_10371,N_10197,N_10193);
nand U10372 (N_10372,N_10150,N_10227);
xor U10373 (N_10373,N_10196,N_10141);
nor U10374 (N_10374,N_10236,N_10218);
and U10375 (N_10375,N_10280,N_10272);
or U10376 (N_10376,N_10261,N_10309);
and U10377 (N_10377,N_10301,N_10372);
nand U10378 (N_10378,N_10279,N_10360);
or U10379 (N_10379,N_10357,N_10342);
or U10380 (N_10380,N_10356,N_10255);
nand U10381 (N_10381,N_10374,N_10288);
and U10382 (N_10382,N_10278,N_10369);
nor U10383 (N_10383,N_10330,N_10274);
and U10384 (N_10384,N_10318,N_10322);
nand U10385 (N_10385,N_10269,N_10340);
xnor U10386 (N_10386,N_10328,N_10316);
or U10387 (N_10387,N_10329,N_10286);
or U10388 (N_10388,N_10271,N_10292);
or U10389 (N_10389,N_10315,N_10281);
nor U10390 (N_10390,N_10289,N_10268);
nor U10391 (N_10391,N_10327,N_10366);
xor U10392 (N_10392,N_10339,N_10338);
or U10393 (N_10393,N_10256,N_10298);
and U10394 (N_10394,N_10364,N_10323);
or U10395 (N_10395,N_10347,N_10262);
xor U10396 (N_10396,N_10326,N_10258);
nor U10397 (N_10397,N_10314,N_10355);
xnor U10398 (N_10398,N_10308,N_10311);
xor U10399 (N_10399,N_10341,N_10295);
xor U10400 (N_10400,N_10349,N_10253);
and U10401 (N_10401,N_10254,N_10276);
nor U10402 (N_10402,N_10319,N_10303);
xnor U10403 (N_10403,N_10275,N_10359);
nor U10404 (N_10404,N_10265,N_10305);
or U10405 (N_10405,N_10307,N_10336);
nand U10406 (N_10406,N_10285,N_10284);
nand U10407 (N_10407,N_10348,N_10373);
or U10408 (N_10408,N_10259,N_10358);
or U10409 (N_10409,N_10310,N_10267);
and U10410 (N_10410,N_10368,N_10252);
xor U10411 (N_10411,N_10335,N_10304);
and U10412 (N_10412,N_10264,N_10331);
or U10413 (N_10413,N_10367,N_10296);
or U10414 (N_10414,N_10302,N_10290);
and U10415 (N_10415,N_10333,N_10334);
nor U10416 (N_10416,N_10352,N_10287);
and U10417 (N_10417,N_10299,N_10365);
nand U10418 (N_10418,N_10282,N_10343);
nand U10419 (N_10419,N_10350,N_10344);
and U10420 (N_10420,N_10371,N_10257);
or U10421 (N_10421,N_10332,N_10263);
and U10422 (N_10422,N_10277,N_10345);
nor U10423 (N_10423,N_10260,N_10251);
nor U10424 (N_10424,N_10351,N_10300);
nor U10425 (N_10425,N_10362,N_10266);
nor U10426 (N_10426,N_10337,N_10306);
and U10427 (N_10427,N_10324,N_10361);
nand U10428 (N_10428,N_10325,N_10317);
and U10429 (N_10429,N_10293,N_10313);
or U10430 (N_10430,N_10354,N_10283);
and U10431 (N_10431,N_10297,N_10312);
nor U10432 (N_10432,N_10353,N_10346);
xor U10433 (N_10433,N_10294,N_10250);
nand U10434 (N_10434,N_10321,N_10370);
or U10435 (N_10435,N_10320,N_10291);
or U10436 (N_10436,N_10273,N_10270);
or U10437 (N_10437,N_10363,N_10367);
nor U10438 (N_10438,N_10287,N_10254);
nand U10439 (N_10439,N_10368,N_10305);
nor U10440 (N_10440,N_10250,N_10298);
or U10441 (N_10441,N_10297,N_10344);
nor U10442 (N_10442,N_10308,N_10293);
or U10443 (N_10443,N_10253,N_10350);
or U10444 (N_10444,N_10261,N_10319);
nor U10445 (N_10445,N_10343,N_10256);
or U10446 (N_10446,N_10287,N_10316);
xnor U10447 (N_10447,N_10335,N_10265);
xnor U10448 (N_10448,N_10281,N_10336);
xnor U10449 (N_10449,N_10300,N_10315);
and U10450 (N_10450,N_10351,N_10321);
and U10451 (N_10451,N_10347,N_10260);
xnor U10452 (N_10452,N_10366,N_10371);
nand U10453 (N_10453,N_10268,N_10321);
or U10454 (N_10454,N_10336,N_10323);
nand U10455 (N_10455,N_10254,N_10373);
nand U10456 (N_10456,N_10282,N_10253);
xnor U10457 (N_10457,N_10347,N_10270);
nor U10458 (N_10458,N_10314,N_10371);
xnor U10459 (N_10459,N_10324,N_10287);
and U10460 (N_10460,N_10336,N_10318);
and U10461 (N_10461,N_10363,N_10259);
or U10462 (N_10462,N_10279,N_10300);
nor U10463 (N_10463,N_10274,N_10360);
nor U10464 (N_10464,N_10289,N_10311);
nand U10465 (N_10465,N_10278,N_10359);
nand U10466 (N_10466,N_10258,N_10310);
or U10467 (N_10467,N_10340,N_10257);
nand U10468 (N_10468,N_10320,N_10289);
and U10469 (N_10469,N_10295,N_10288);
nor U10470 (N_10470,N_10261,N_10294);
xnor U10471 (N_10471,N_10350,N_10356);
or U10472 (N_10472,N_10312,N_10258);
xor U10473 (N_10473,N_10366,N_10311);
and U10474 (N_10474,N_10270,N_10365);
nor U10475 (N_10475,N_10276,N_10347);
nand U10476 (N_10476,N_10290,N_10367);
xnor U10477 (N_10477,N_10353,N_10273);
nor U10478 (N_10478,N_10371,N_10323);
nor U10479 (N_10479,N_10349,N_10304);
xor U10480 (N_10480,N_10273,N_10365);
nand U10481 (N_10481,N_10263,N_10317);
xnor U10482 (N_10482,N_10328,N_10300);
xnor U10483 (N_10483,N_10350,N_10289);
nor U10484 (N_10484,N_10358,N_10260);
nand U10485 (N_10485,N_10263,N_10278);
xor U10486 (N_10486,N_10274,N_10288);
xor U10487 (N_10487,N_10303,N_10329);
nor U10488 (N_10488,N_10361,N_10299);
nand U10489 (N_10489,N_10255,N_10281);
nand U10490 (N_10490,N_10264,N_10288);
or U10491 (N_10491,N_10329,N_10284);
nand U10492 (N_10492,N_10359,N_10311);
xor U10493 (N_10493,N_10277,N_10270);
nand U10494 (N_10494,N_10278,N_10297);
and U10495 (N_10495,N_10301,N_10323);
nor U10496 (N_10496,N_10297,N_10292);
nand U10497 (N_10497,N_10253,N_10326);
xnor U10498 (N_10498,N_10260,N_10313);
and U10499 (N_10499,N_10277,N_10336);
and U10500 (N_10500,N_10479,N_10453);
nand U10501 (N_10501,N_10456,N_10435);
or U10502 (N_10502,N_10396,N_10381);
or U10503 (N_10503,N_10442,N_10491);
xor U10504 (N_10504,N_10473,N_10388);
or U10505 (N_10505,N_10413,N_10380);
or U10506 (N_10506,N_10402,N_10411);
and U10507 (N_10507,N_10400,N_10450);
and U10508 (N_10508,N_10393,N_10457);
nor U10509 (N_10509,N_10446,N_10461);
and U10510 (N_10510,N_10385,N_10485);
nand U10511 (N_10511,N_10391,N_10474);
nand U10512 (N_10512,N_10459,N_10403);
nor U10513 (N_10513,N_10395,N_10497);
or U10514 (N_10514,N_10472,N_10437);
nand U10515 (N_10515,N_10423,N_10431);
xnor U10516 (N_10516,N_10392,N_10495);
xor U10517 (N_10517,N_10469,N_10428);
and U10518 (N_10518,N_10464,N_10488);
and U10519 (N_10519,N_10451,N_10484);
xor U10520 (N_10520,N_10470,N_10487);
nand U10521 (N_10521,N_10376,N_10440);
xnor U10522 (N_10522,N_10489,N_10438);
nor U10523 (N_10523,N_10415,N_10468);
nand U10524 (N_10524,N_10441,N_10454);
or U10525 (N_10525,N_10421,N_10406);
or U10526 (N_10526,N_10445,N_10434);
and U10527 (N_10527,N_10409,N_10412);
and U10528 (N_10528,N_10444,N_10462);
xnor U10529 (N_10529,N_10493,N_10455);
and U10530 (N_10530,N_10420,N_10443);
nor U10531 (N_10531,N_10398,N_10378);
and U10532 (N_10532,N_10448,N_10382);
xor U10533 (N_10533,N_10426,N_10430);
nand U10534 (N_10534,N_10481,N_10399);
nor U10535 (N_10535,N_10404,N_10418);
nor U10536 (N_10536,N_10486,N_10383);
nand U10537 (N_10537,N_10460,N_10436);
nand U10538 (N_10538,N_10414,N_10439);
nor U10539 (N_10539,N_10490,N_10408);
and U10540 (N_10540,N_10390,N_10427);
nor U10541 (N_10541,N_10480,N_10496);
or U10542 (N_10542,N_10384,N_10416);
and U10543 (N_10543,N_10458,N_10432);
nand U10544 (N_10544,N_10466,N_10463);
nand U10545 (N_10545,N_10483,N_10375);
or U10546 (N_10546,N_10477,N_10498);
or U10547 (N_10547,N_10405,N_10379);
nand U10548 (N_10548,N_10419,N_10482);
xor U10549 (N_10549,N_10452,N_10447);
xnor U10550 (N_10550,N_10377,N_10475);
and U10551 (N_10551,N_10389,N_10465);
nand U10552 (N_10552,N_10494,N_10492);
and U10553 (N_10553,N_10422,N_10425);
xor U10554 (N_10554,N_10449,N_10499);
xnor U10555 (N_10555,N_10476,N_10386);
xor U10556 (N_10556,N_10433,N_10478);
and U10557 (N_10557,N_10471,N_10429);
xor U10558 (N_10558,N_10467,N_10401);
xor U10559 (N_10559,N_10410,N_10407);
or U10560 (N_10560,N_10387,N_10424);
and U10561 (N_10561,N_10397,N_10417);
and U10562 (N_10562,N_10394,N_10380);
xor U10563 (N_10563,N_10384,N_10477);
nand U10564 (N_10564,N_10441,N_10381);
nand U10565 (N_10565,N_10424,N_10457);
nand U10566 (N_10566,N_10390,N_10440);
nand U10567 (N_10567,N_10488,N_10490);
nand U10568 (N_10568,N_10415,N_10489);
nor U10569 (N_10569,N_10394,N_10403);
nor U10570 (N_10570,N_10382,N_10472);
nand U10571 (N_10571,N_10488,N_10474);
or U10572 (N_10572,N_10475,N_10484);
and U10573 (N_10573,N_10477,N_10454);
xnor U10574 (N_10574,N_10388,N_10499);
or U10575 (N_10575,N_10389,N_10458);
or U10576 (N_10576,N_10455,N_10459);
or U10577 (N_10577,N_10449,N_10391);
and U10578 (N_10578,N_10393,N_10419);
xor U10579 (N_10579,N_10486,N_10456);
and U10580 (N_10580,N_10488,N_10478);
nand U10581 (N_10581,N_10447,N_10492);
and U10582 (N_10582,N_10477,N_10471);
nor U10583 (N_10583,N_10485,N_10463);
nor U10584 (N_10584,N_10381,N_10480);
nand U10585 (N_10585,N_10427,N_10447);
or U10586 (N_10586,N_10428,N_10451);
or U10587 (N_10587,N_10441,N_10485);
and U10588 (N_10588,N_10486,N_10492);
and U10589 (N_10589,N_10404,N_10452);
xnor U10590 (N_10590,N_10398,N_10477);
nand U10591 (N_10591,N_10418,N_10478);
or U10592 (N_10592,N_10449,N_10424);
nor U10593 (N_10593,N_10467,N_10455);
xor U10594 (N_10594,N_10491,N_10459);
nor U10595 (N_10595,N_10375,N_10484);
nor U10596 (N_10596,N_10437,N_10452);
and U10597 (N_10597,N_10433,N_10444);
or U10598 (N_10598,N_10387,N_10388);
nor U10599 (N_10599,N_10459,N_10480);
or U10600 (N_10600,N_10429,N_10414);
xor U10601 (N_10601,N_10493,N_10470);
and U10602 (N_10602,N_10420,N_10484);
and U10603 (N_10603,N_10429,N_10492);
and U10604 (N_10604,N_10471,N_10425);
or U10605 (N_10605,N_10396,N_10427);
or U10606 (N_10606,N_10477,N_10417);
xor U10607 (N_10607,N_10422,N_10443);
nor U10608 (N_10608,N_10476,N_10478);
nand U10609 (N_10609,N_10444,N_10424);
nand U10610 (N_10610,N_10433,N_10422);
or U10611 (N_10611,N_10399,N_10468);
or U10612 (N_10612,N_10474,N_10384);
nor U10613 (N_10613,N_10486,N_10488);
or U10614 (N_10614,N_10480,N_10477);
nor U10615 (N_10615,N_10387,N_10426);
xnor U10616 (N_10616,N_10493,N_10381);
nand U10617 (N_10617,N_10428,N_10377);
nand U10618 (N_10618,N_10497,N_10381);
nor U10619 (N_10619,N_10419,N_10473);
or U10620 (N_10620,N_10490,N_10401);
or U10621 (N_10621,N_10425,N_10450);
or U10622 (N_10622,N_10422,N_10429);
or U10623 (N_10623,N_10495,N_10448);
xor U10624 (N_10624,N_10463,N_10435);
and U10625 (N_10625,N_10592,N_10563);
nand U10626 (N_10626,N_10589,N_10500);
nand U10627 (N_10627,N_10523,N_10618);
or U10628 (N_10628,N_10516,N_10606);
xor U10629 (N_10629,N_10614,N_10507);
nor U10630 (N_10630,N_10531,N_10543);
xor U10631 (N_10631,N_10577,N_10527);
and U10632 (N_10632,N_10539,N_10542);
xor U10633 (N_10633,N_10508,N_10587);
nor U10634 (N_10634,N_10502,N_10530);
and U10635 (N_10635,N_10571,N_10550);
nor U10636 (N_10636,N_10552,N_10521);
nor U10637 (N_10637,N_10533,N_10566);
nand U10638 (N_10638,N_10528,N_10522);
nand U10639 (N_10639,N_10600,N_10611);
and U10640 (N_10640,N_10619,N_10610);
nor U10641 (N_10641,N_10593,N_10561);
and U10642 (N_10642,N_10613,N_10564);
and U10643 (N_10643,N_10590,N_10517);
and U10644 (N_10644,N_10540,N_10513);
and U10645 (N_10645,N_10570,N_10535);
xnor U10646 (N_10646,N_10558,N_10608);
xnor U10647 (N_10647,N_10576,N_10588);
xnor U10648 (N_10648,N_10504,N_10605);
or U10649 (N_10649,N_10572,N_10599);
nand U10650 (N_10650,N_10519,N_10612);
and U10651 (N_10651,N_10551,N_10574);
nor U10652 (N_10652,N_10556,N_10511);
nand U10653 (N_10653,N_10586,N_10622);
xor U10654 (N_10654,N_10615,N_10545);
nand U10655 (N_10655,N_10529,N_10503);
nor U10656 (N_10656,N_10510,N_10601);
nand U10657 (N_10657,N_10617,N_10621);
nand U10658 (N_10658,N_10569,N_10505);
and U10659 (N_10659,N_10526,N_10562);
nor U10660 (N_10660,N_10509,N_10581);
xnor U10661 (N_10661,N_10538,N_10541);
and U10662 (N_10662,N_10501,N_10568);
nor U10663 (N_10663,N_10537,N_10560);
nor U10664 (N_10664,N_10514,N_10554);
xor U10665 (N_10665,N_10575,N_10515);
nand U10666 (N_10666,N_10547,N_10524);
or U10667 (N_10667,N_10609,N_10525);
nor U10668 (N_10668,N_10506,N_10520);
xor U10669 (N_10669,N_10548,N_10578);
nor U10670 (N_10670,N_10534,N_10532);
nor U10671 (N_10671,N_10596,N_10546);
and U10672 (N_10672,N_10555,N_10580);
and U10673 (N_10673,N_10518,N_10557);
nor U10674 (N_10674,N_10579,N_10602);
xor U10675 (N_10675,N_10544,N_10598);
or U10676 (N_10676,N_10597,N_10603);
xor U10677 (N_10677,N_10607,N_10583);
nor U10678 (N_10678,N_10567,N_10512);
nand U10679 (N_10679,N_10559,N_10553);
or U10680 (N_10680,N_10624,N_10594);
nand U10681 (N_10681,N_10549,N_10623);
xnor U10682 (N_10682,N_10604,N_10582);
nand U10683 (N_10683,N_10591,N_10595);
or U10684 (N_10684,N_10616,N_10565);
or U10685 (N_10685,N_10585,N_10536);
xnor U10686 (N_10686,N_10573,N_10620);
nor U10687 (N_10687,N_10584,N_10548);
or U10688 (N_10688,N_10548,N_10603);
nor U10689 (N_10689,N_10547,N_10598);
nor U10690 (N_10690,N_10583,N_10580);
xor U10691 (N_10691,N_10605,N_10623);
nor U10692 (N_10692,N_10607,N_10527);
xnor U10693 (N_10693,N_10520,N_10579);
or U10694 (N_10694,N_10518,N_10541);
and U10695 (N_10695,N_10591,N_10613);
nor U10696 (N_10696,N_10557,N_10574);
nand U10697 (N_10697,N_10557,N_10617);
or U10698 (N_10698,N_10539,N_10584);
or U10699 (N_10699,N_10551,N_10523);
xor U10700 (N_10700,N_10501,N_10516);
and U10701 (N_10701,N_10579,N_10555);
or U10702 (N_10702,N_10591,N_10506);
and U10703 (N_10703,N_10514,N_10592);
nor U10704 (N_10704,N_10543,N_10519);
nand U10705 (N_10705,N_10528,N_10624);
nand U10706 (N_10706,N_10593,N_10566);
or U10707 (N_10707,N_10579,N_10593);
nor U10708 (N_10708,N_10531,N_10566);
and U10709 (N_10709,N_10554,N_10577);
nand U10710 (N_10710,N_10581,N_10576);
or U10711 (N_10711,N_10598,N_10581);
nor U10712 (N_10712,N_10529,N_10620);
or U10713 (N_10713,N_10508,N_10560);
or U10714 (N_10714,N_10604,N_10596);
xnor U10715 (N_10715,N_10502,N_10596);
and U10716 (N_10716,N_10524,N_10616);
or U10717 (N_10717,N_10567,N_10514);
or U10718 (N_10718,N_10568,N_10543);
nor U10719 (N_10719,N_10585,N_10550);
and U10720 (N_10720,N_10513,N_10530);
xor U10721 (N_10721,N_10620,N_10512);
and U10722 (N_10722,N_10568,N_10589);
or U10723 (N_10723,N_10590,N_10551);
xnor U10724 (N_10724,N_10532,N_10517);
nand U10725 (N_10725,N_10613,N_10503);
xor U10726 (N_10726,N_10527,N_10616);
nand U10727 (N_10727,N_10523,N_10545);
nand U10728 (N_10728,N_10501,N_10561);
xor U10729 (N_10729,N_10619,N_10518);
and U10730 (N_10730,N_10610,N_10566);
nand U10731 (N_10731,N_10545,N_10501);
nand U10732 (N_10732,N_10515,N_10505);
or U10733 (N_10733,N_10558,N_10533);
or U10734 (N_10734,N_10507,N_10558);
or U10735 (N_10735,N_10529,N_10527);
xor U10736 (N_10736,N_10531,N_10578);
nor U10737 (N_10737,N_10549,N_10521);
nor U10738 (N_10738,N_10508,N_10539);
nand U10739 (N_10739,N_10574,N_10547);
xnor U10740 (N_10740,N_10575,N_10552);
nand U10741 (N_10741,N_10599,N_10554);
nor U10742 (N_10742,N_10582,N_10562);
xor U10743 (N_10743,N_10591,N_10582);
nand U10744 (N_10744,N_10593,N_10508);
nand U10745 (N_10745,N_10609,N_10621);
and U10746 (N_10746,N_10503,N_10554);
xnor U10747 (N_10747,N_10555,N_10523);
xnor U10748 (N_10748,N_10526,N_10553);
nand U10749 (N_10749,N_10591,N_10611);
nand U10750 (N_10750,N_10715,N_10651);
nor U10751 (N_10751,N_10648,N_10644);
xor U10752 (N_10752,N_10718,N_10713);
and U10753 (N_10753,N_10627,N_10642);
nor U10754 (N_10754,N_10668,N_10685);
or U10755 (N_10755,N_10664,N_10730);
and U10756 (N_10756,N_10725,N_10721);
nor U10757 (N_10757,N_10655,N_10714);
xor U10758 (N_10758,N_10739,N_10654);
nor U10759 (N_10759,N_10649,N_10704);
or U10760 (N_10760,N_10724,N_10632);
nor U10761 (N_10761,N_10639,N_10660);
and U10762 (N_10762,N_10650,N_10638);
nor U10763 (N_10763,N_10706,N_10677);
nand U10764 (N_10764,N_10705,N_10686);
and U10765 (N_10765,N_10740,N_10747);
nand U10766 (N_10766,N_10625,N_10667);
and U10767 (N_10767,N_10736,N_10675);
xor U10768 (N_10768,N_10733,N_10681);
and U10769 (N_10769,N_10701,N_10643);
xor U10770 (N_10770,N_10663,N_10645);
and U10771 (N_10771,N_10676,N_10631);
and U10772 (N_10772,N_10687,N_10628);
nand U10773 (N_10773,N_10744,N_10629);
xnor U10774 (N_10774,N_10743,N_10732);
xnor U10775 (N_10775,N_10712,N_10722);
and U10776 (N_10776,N_10646,N_10696);
nand U10777 (N_10777,N_10693,N_10683);
nand U10778 (N_10778,N_10689,N_10717);
and U10779 (N_10779,N_10734,N_10727);
and U10780 (N_10780,N_10695,N_10690);
or U10781 (N_10781,N_10708,N_10694);
nand U10782 (N_10782,N_10640,N_10634);
xor U10783 (N_10783,N_10659,N_10636);
nor U10784 (N_10784,N_10728,N_10633);
and U10785 (N_10785,N_10657,N_10662);
or U10786 (N_10786,N_10720,N_10680);
or U10787 (N_10787,N_10674,N_10738);
xor U10788 (N_10788,N_10691,N_10656);
xor U10789 (N_10789,N_10710,N_10742);
xnor U10790 (N_10790,N_10658,N_10684);
xnor U10791 (N_10791,N_10726,N_10711);
xor U10792 (N_10792,N_10748,N_10678);
or U10793 (N_10793,N_10653,N_10647);
or U10794 (N_10794,N_10703,N_10707);
xnor U10795 (N_10795,N_10635,N_10749);
nand U10796 (N_10796,N_10637,N_10692);
nand U10797 (N_10797,N_10731,N_10745);
xnor U10798 (N_10798,N_10702,N_10716);
and U10799 (N_10799,N_10666,N_10729);
or U10800 (N_10800,N_10688,N_10709);
nand U10801 (N_10801,N_10741,N_10626);
nand U10802 (N_10802,N_10671,N_10641);
xor U10803 (N_10803,N_10665,N_10700);
nor U10804 (N_10804,N_10698,N_10661);
xnor U10805 (N_10805,N_10682,N_10652);
nor U10806 (N_10806,N_10699,N_10679);
or U10807 (N_10807,N_10697,N_10719);
or U10808 (N_10808,N_10669,N_10630);
xnor U10809 (N_10809,N_10735,N_10672);
xnor U10810 (N_10810,N_10737,N_10670);
nor U10811 (N_10811,N_10746,N_10723);
and U10812 (N_10812,N_10673,N_10674);
nor U10813 (N_10813,N_10685,N_10701);
xor U10814 (N_10814,N_10666,N_10737);
or U10815 (N_10815,N_10717,N_10632);
xor U10816 (N_10816,N_10707,N_10743);
nand U10817 (N_10817,N_10733,N_10729);
or U10818 (N_10818,N_10704,N_10673);
xnor U10819 (N_10819,N_10661,N_10749);
and U10820 (N_10820,N_10731,N_10672);
xor U10821 (N_10821,N_10703,N_10654);
xor U10822 (N_10822,N_10641,N_10731);
nand U10823 (N_10823,N_10639,N_10668);
xor U10824 (N_10824,N_10630,N_10702);
xnor U10825 (N_10825,N_10663,N_10635);
xor U10826 (N_10826,N_10713,N_10734);
xnor U10827 (N_10827,N_10689,N_10626);
or U10828 (N_10828,N_10697,N_10671);
nand U10829 (N_10829,N_10744,N_10749);
nor U10830 (N_10830,N_10712,N_10654);
nand U10831 (N_10831,N_10710,N_10708);
nand U10832 (N_10832,N_10666,N_10639);
or U10833 (N_10833,N_10731,N_10634);
or U10834 (N_10834,N_10636,N_10638);
nand U10835 (N_10835,N_10635,N_10691);
nand U10836 (N_10836,N_10651,N_10625);
and U10837 (N_10837,N_10642,N_10651);
xnor U10838 (N_10838,N_10703,N_10659);
nor U10839 (N_10839,N_10695,N_10650);
or U10840 (N_10840,N_10685,N_10728);
or U10841 (N_10841,N_10632,N_10723);
nand U10842 (N_10842,N_10658,N_10641);
and U10843 (N_10843,N_10638,N_10714);
or U10844 (N_10844,N_10664,N_10646);
xor U10845 (N_10845,N_10660,N_10678);
or U10846 (N_10846,N_10657,N_10738);
nand U10847 (N_10847,N_10666,N_10711);
or U10848 (N_10848,N_10660,N_10710);
xnor U10849 (N_10849,N_10683,N_10732);
or U10850 (N_10850,N_10655,N_10717);
and U10851 (N_10851,N_10677,N_10739);
or U10852 (N_10852,N_10728,N_10631);
nand U10853 (N_10853,N_10728,N_10738);
or U10854 (N_10854,N_10670,N_10648);
and U10855 (N_10855,N_10655,N_10749);
and U10856 (N_10856,N_10655,N_10634);
or U10857 (N_10857,N_10633,N_10725);
nand U10858 (N_10858,N_10731,N_10679);
or U10859 (N_10859,N_10711,N_10671);
and U10860 (N_10860,N_10734,N_10739);
and U10861 (N_10861,N_10690,N_10680);
nor U10862 (N_10862,N_10666,N_10637);
xor U10863 (N_10863,N_10740,N_10710);
xor U10864 (N_10864,N_10644,N_10679);
nand U10865 (N_10865,N_10713,N_10656);
nor U10866 (N_10866,N_10675,N_10646);
nor U10867 (N_10867,N_10704,N_10718);
and U10868 (N_10868,N_10699,N_10711);
nand U10869 (N_10869,N_10649,N_10645);
or U10870 (N_10870,N_10714,N_10637);
or U10871 (N_10871,N_10696,N_10630);
xor U10872 (N_10872,N_10702,N_10658);
nor U10873 (N_10873,N_10687,N_10655);
nor U10874 (N_10874,N_10647,N_10729);
nor U10875 (N_10875,N_10825,N_10848);
nor U10876 (N_10876,N_10857,N_10776);
nand U10877 (N_10877,N_10775,N_10774);
nand U10878 (N_10878,N_10792,N_10765);
nor U10879 (N_10879,N_10771,N_10809);
nand U10880 (N_10880,N_10789,N_10832);
or U10881 (N_10881,N_10852,N_10863);
xnor U10882 (N_10882,N_10833,N_10760);
nor U10883 (N_10883,N_10821,N_10847);
nand U10884 (N_10884,N_10758,N_10800);
nor U10885 (N_10885,N_10845,N_10777);
nand U10886 (N_10886,N_10864,N_10838);
xor U10887 (N_10887,N_10868,N_10843);
nand U10888 (N_10888,N_10766,N_10813);
xnor U10889 (N_10889,N_10824,N_10820);
and U10890 (N_10890,N_10778,N_10869);
or U10891 (N_10891,N_10815,N_10768);
nand U10892 (N_10892,N_10779,N_10803);
nor U10893 (N_10893,N_10783,N_10859);
or U10894 (N_10894,N_10811,N_10871);
and U10895 (N_10895,N_10804,N_10819);
nand U10896 (N_10896,N_10769,N_10849);
nor U10897 (N_10897,N_10851,N_10806);
and U10898 (N_10898,N_10814,N_10796);
or U10899 (N_10899,N_10782,N_10830);
or U10900 (N_10900,N_10767,N_10764);
or U10901 (N_10901,N_10754,N_10785);
or U10902 (N_10902,N_10798,N_10750);
xnor U10903 (N_10903,N_10772,N_10829);
and U10904 (N_10904,N_10795,N_10874);
or U10905 (N_10905,N_10816,N_10836);
nand U10906 (N_10906,N_10788,N_10794);
nor U10907 (N_10907,N_10841,N_10834);
nor U10908 (N_10908,N_10801,N_10812);
nor U10909 (N_10909,N_10827,N_10831);
and U10910 (N_10910,N_10751,N_10786);
nor U10911 (N_10911,N_10773,N_10854);
nor U10912 (N_10912,N_10844,N_10850);
and U10913 (N_10913,N_10872,N_10837);
nor U10914 (N_10914,N_10793,N_10808);
nand U10915 (N_10915,N_10826,N_10858);
xor U10916 (N_10916,N_10762,N_10805);
xor U10917 (N_10917,N_10790,N_10752);
xnor U10918 (N_10918,N_10853,N_10761);
and U10919 (N_10919,N_10861,N_10781);
or U10920 (N_10920,N_10770,N_10870);
or U10921 (N_10921,N_10784,N_10763);
and U10922 (N_10922,N_10865,N_10818);
nor U10923 (N_10923,N_10835,N_10856);
and U10924 (N_10924,N_10757,N_10822);
nor U10925 (N_10925,N_10787,N_10873);
nand U10926 (N_10926,N_10802,N_10860);
nor U10927 (N_10927,N_10817,N_10755);
and U10928 (N_10928,N_10840,N_10866);
or U10929 (N_10929,N_10753,N_10797);
or U10930 (N_10930,N_10759,N_10846);
or U10931 (N_10931,N_10842,N_10756);
xnor U10932 (N_10932,N_10810,N_10828);
or U10933 (N_10933,N_10780,N_10791);
nand U10934 (N_10934,N_10807,N_10799);
nor U10935 (N_10935,N_10823,N_10855);
nand U10936 (N_10936,N_10839,N_10867);
nand U10937 (N_10937,N_10862,N_10856);
xnor U10938 (N_10938,N_10859,N_10781);
or U10939 (N_10939,N_10870,N_10778);
xnor U10940 (N_10940,N_10852,N_10815);
and U10941 (N_10941,N_10826,N_10811);
xnor U10942 (N_10942,N_10771,N_10836);
or U10943 (N_10943,N_10865,N_10823);
xor U10944 (N_10944,N_10803,N_10847);
nand U10945 (N_10945,N_10799,N_10874);
nor U10946 (N_10946,N_10774,N_10785);
or U10947 (N_10947,N_10860,N_10751);
or U10948 (N_10948,N_10761,N_10768);
nor U10949 (N_10949,N_10788,N_10824);
nor U10950 (N_10950,N_10856,N_10823);
nor U10951 (N_10951,N_10807,N_10832);
and U10952 (N_10952,N_10832,N_10796);
nor U10953 (N_10953,N_10849,N_10756);
and U10954 (N_10954,N_10869,N_10751);
nor U10955 (N_10955,N_10815,N_10760);
nor U10956 (N_10956,N_10792,N_10840);
or U10957 (N_10957,N_10858,N_10841);
or U10958 (N_10958,N_10852,N_10798);
and U10959 (N_10959,N_10823,N_10799);
nand U10960 (N_10960,N_10835,N_10834);
nand U10961 (N_10961,N_10788,N_10810);
nand U10962 (N_10962,N_10753,N_10848);
xnor U10963 (N_10963,N_10865,N_10769);
and U10964 (N_10964,N_10827,N_10865);
xnor U10965 (N_10965,N_10779,N_10822);
and U10966 (N_10966,N_10764,N_10873);
and U10967 (N_10967,N_10819,N_10799);
xnor U10968 (N_10968,N_10806,N_10844);
and U10969 (N_10969,N_10838,N_10859);
or U10970 (N_10970,N_10826,N_10787);
or U10971 (N_10971,N_10824,N_10828);
or U10972 (N_10972,N_10794,N_10792);
nor U10973 (N_10973,N_10809,N_10760);
nand U10974 (N_10974,N_10839,N_10874);
xor U10975 (N_10975,N_10765,N_10842);
nand U10976 (N_10976,N_10759,N_10817);
xnor U10977 (N_10977,N_10839,N_10756);
xor U10978 (N_10978,N_10869,N_10844);
nand U10979 (N_10979,N_10848,N_10766);
and U10980 (N_10980,N_10796,N_10807);
nor U10981 (N_10981,N_10874,N_10824);
nand U10982 (N_10982,N_10874,N_10869);
or U10983 (N_10983,N_10800,N_10783);
nor U10984 (N_10984,N_10823,N_10789);
and U10985 (N_10985,N_10784,N_10834);
or U10986 (N_10986,N_10822,N_10869);
nor U10987 (N_10987,N_10805,N_10826);
xor U10988 (N_10988,N_10820,N_10867);
nor U10989 (N_10989,N_10854,N_10819);
or U10990 (N_10990,N_10851,N_10797);
and U10991 (N_10991,N_10852,N_10842);
nand U10992 (N_10992,N_10783,N_10848);
xor U10993 (N_10993,N_10792,N_10788);
xor U10994 (N_10994,N_10770,N_10844);
xor U10995 (N_10995,N_10869,N_10849);
and U10996 (N_10996,N_10817,N_10761);
xnor U10997 (N_10997,N_10869,N_10813);
nor U10998 (N_10998,N_10869,N_10850);
and U10999 (N_10999,N_10786,N_10835);
nand U11000 (N_11000,N_10929,N_10997);
nor U11001 (N_11001,N_10915,N_10923);
and U11002 (N_11002,N_10937,N_10916);
and U11003 (N_11003,N_10903,N_10947);
or U11004 (N_11004,N_10967,N_10930);
and U11005 (N_11005,N_10880,N_10894);
and U11006 (N_11006,N_10898,N_10983);
nand U11007 (N_11007,N_10910,N_10987);
or U11008 (N_11008,N_10912,N_10934);
nand U11009 (N_11009,N_10900,N_10984);
or U11010 (N_11010,N_10927,N_10952);
nand U11011 (N_11011,N_10981,N_10978);
xnor U11012 (N_11012,N_10932,N_10877);
nand U11013 (N_11013,N_10922,N_10897);
xor U11014 (N_11014,N_10973,N_10999);
nand U11015 (N_11015,N_10969,N_10881);
and U11016 (N_11016,N_10919,N_10931);
and U11017 (N_11017,N_10892,N_10977);
nand U11018 (N_11018,N_10926,N_10996);
nor U11019 (N_11019,N_10879,N_10909);
and U11020 (N_11020,N_10875,N_10976);
nor U11021 (N_11021,N_10908,N_10913);
nand U11022 (N_11022,N_10960,N_10975);
nand U11023 (N_11023,N_10959,N_10914);
and U11024 (N_11024,N_10985,N_10886);
and U11025 (N_11025,N_10882,N_10933);
nand U11026 (N_11026,N_10962,N_10995);
xnor U11027 (N_11027,N_10949,N_10951);
and U11028 (N_11028,N_10940,N_10905);
or U11029 (N_11029,N_10893,N_10889);
and U11030 (N_11030,N_10925,N_10979);
nand U11031 (N_11031,N_10918,N_10911);
and U11032 (N_11032,N_10974,N_10986);
or U11033 (N_11033,N_10955,N_10921);
xor U11034 (N_11034,N_10891,N_10964);
or U11035 (N_11035,N_10943,N_10991);
nor U11036 (N_11036,N_10904,N_10878);
xor U11037 (N_11037,N_10953,N_10902);
or U11038 (N_11038,N_10939,N_10998);
and U11039 (N_11039,N_10907,N_10982);
nor U11040 (N_11040,N_10938,N_10970);
or U11041 (N_11041,N_10945,N_10989);
nor U11042 (N_11042,N_10946,N_10906);
nand U11043 (N_11043,N_10888,N_10884);
or U11044 (N_11044,N_10990,N_10885);
nand U11045 (N_11045,N_10883,N_10971);
nand U11046 (N_11046,N_10890,N_10965);
nor U11047 (N_11047,N_10917,N_10896);
xnor U11048 (N_11048,N_10901,N_10972);
xor U11049 (N_11049,N_10956,N_10948);
nand U11050 (N_11050,N_10876,N_10950);
and U11051 (N_11051,N_10994,N_10935);
and U11052 (N_11052,N_10992,N_10941);
nor U11053 (N_11053,N_10957,N_10899);
nand U11054 (N_11054,N_10961,N_10928);
and U11055 (N_11055,N_10920,N_10895);
xnor U11056 (N_11056,N_10944,N_10966);
and U11057 (N_11057,N_10942,N_10980);
or U11058 (N_11058,N_10968,N_10936);
nor U11059 (N_11059,N_10887,N_10963);
nor U11060 (N_11060,N_10988,N_10954);
or U11061 (N_11061,N_10958,N_10924);
nand U11062 (N_11062,N_10993,N_10926);
xnor U11063 (N_11063,N_10950,N_10960);
nand U11064 (N_11064,N_10884,N_10889);
and U11065 (N_11065,N_10885,N_10894);
nand U11066 (N_11066,N_10907,N_10997);
or U11067 (N_11067,N_10892,N_10910);
or U11068 (N_11068,N_10931,N_10938);
nand U11069 (N_11069,N_10884,N_10972);
nand U11070 (N_11070,N_10920,N_10964);
xnor U11071 (N_11071,N_10940,N_10934);
nand U11072 (N_11072,N_10948,N_10906);
nand U11073 (N_11073,N_10955,N_10987);
and U11074 (N_11074,N_10926,N_10897);
xnor U11075 (N_11075,N_10919,N_10936);
xnor U11076 (N_11076,N_10949,N_10971);
and U11077 (N_11077,N_10969,N_10891);
nand U11078 (N_11078,N_10908,N_10878);
nand U11079 (N_11079,N_10900,N_10968);
xnor U11080 (N_11080,N_10916,N_10972);
and U11081 (N_11081,N_10986,N_10879);
xnor U11082 (N_11082,N_10938,N_10911);
and U11083 (N_11083,N_10910,N_10935);
or U11084 (N_11084,N_10922,N_10977);
nor U11085 (N_11085,N_10923,N_10899);
nand U11086 (N_11086,N_10969,N_10900);
xnor U11087 (N_11087,N_10893,N_10969);
xor U11088 (N_11088,N_10966,N_10940);
nand U11089 (N_11089,N_10959,N_10967);
or U11090 (N_11090,N_10957,N_10965);
and U11091 (N_11091,N_10952,N_10973);
or U11092 (N_11092,N_10949,N_10969);
nor U11093 (N_11093,N_10972,N_10991);
xor U11094 (N_11094,N_10897,N_10913);
or U11095 (N_11095,N_10918,N_10976);
xnor U11096 (N_11096,N_10940,N_10981);
or U11097 (N_11097,N_10970,N_10971);
or U11098 (N_11098,N_10995,N_10957);
or U11099 (N_11099,N_10896,N_10901);
nand U11100 (N_11100,N_10941,N_10934);
xor U11101 (N_11101,N_10883,N_10978);
nor U11102 (N_11102,N_10987,N_10887);
and U11103 (N_11103,N_10962,N_10932);
nand U11104 (N_11104,N_10968,N_10945);
nand U11105 (N_11105,N_10939,N_10936);
or U11106 (N_11106,N_10888,N_10972);
or U11107 (N_11107,N_10925,N_10880);
xor U11108 (N_11108,N_10962,N_10989);
or U11109 (N_11109,N_10957,N_10890);
nor U11110 (N_11110,N_10975,N_10884);
xnor U11111 (N_11111,N_10947,N_10986);
or U11112 (N_11112,N_10965,N_10915);
or U11113 (N_11113,N_10888,N_10877);
nand U11114 (N_11114,N_10876,N_10907);
xor U11115 (N_11115,N_10925,N_10945);
or U11116 (N_11116,N_10905,N_10908);
and U11117 (N_11117,N_10933,N_10958);
xor U11118 (N_11118,N_10945,N_10914);
xor U11119 (N_11119,N_10949,N_10975);
xor U11120 (N_11120,N_10890,N_10989);
xnor U11121 (N_11121,N_10985,N_10941);
or U11122 (N_11122,N_10919,N_10978);
or U11123 (N_11123,N_10940,N_10889);
nand U11124 (N_11124,N_10946,N_10979);
and U11125 (N_11125,N_11076,N_11105);
or U11126 (N_11126,N_11087,N_11046);
and U11127 (N_11127,N_11038,N_11118);
or U11128 (N_11128,N_11096,N_11034);
or U11129 (N_11129,N_11006,N_11120);
nor U11130 (N_11130,N_11123,N_11112);
nand U11131 (N_11131,N_11021,N_11012);
and U11132 (N_11132,N_11124,N_11094);
nor U11133 (N_11133,N_11022,N_11019);
xor U11134 (N_11134,N_11071,N_11050);
and U11135 (N_11135,N_11007,N_11063);
nand U11136 (N_11136,N_11069,N_11113);
and U11137 (N_11137,N_11080,N_11001);
xor U11138 (N_11138,N_11008,N_11093);
nand U11139 (N_11139,N_11117,N_11029);
xnor U11140 (N_11140,N_11033,N_11020);
and U11141 (N_11141,N_11106,N_11043);
and U11142 (N_11142,N_11010,N_11041);
and U11143 (N_11143,N_11100,N_11060);
nor U11144 (N_11144,N_11055,N_11122);
nand U11145 (N_11145,N_11099,N_11025);
nand U11146 (N_11146,N_11049,N_11109);
and U11147 (N_11147,N_11115,N_11078);
xnor U11148 (N_11148,N_11037,N_11042);
or U11149 (N_11149,N_11104,N_11013);
nand U11150 (N_11150,N_11075,N_11040);
xor U11151 (N_11151,N_11086,N_11068);
nor U11152 (N_11152,N_11107,N_11039);
nor U11153 (N_11153,N_11091,N_11079);
nor U11154 (N_11154,N_11000,N_11056);
nor U11155 (N_11155,N_11002,N_11088);
nor U11156 (N_11156,N_11030,N_11121);
or U11157 (N_11157,N_11072,N_11083);
nor U11158 (N_11158,N_11015,N_11102);
nor U11159 (N_11159,N_11057,N_11048);
nand U11160 (N_11160,N_11066,N_11101);
and U11161 (N_11161,N_11045,N_11116);
and U11162 (N_11162,N_11077,N_11110);
xor U11163 (N_11163,N_11061,N_11114);
and U11164 (N_11164,N_11005,N_11097);
nand U11165 (N_11165,N_11017,N_11082);
nand U11166 (N_11166,N_11058,N_11044);
xnor U11167 (N_11167,N_11062,N_11073);
nand U11168 (N_11168,N_11089,N_11014);
nor U11169 (N_11169,N_11064,N_11092);
or U11170 (N_11170,N_11051,N_11095);
xnor U11171 (N_11171,N_11052,N_11081);
nand U11172 (N_11172,N_11024,N_11074);
and U11173 (N_11173,N_11084,N_11111);
nand U11174 (N_11174,N_11009,N_11018);
nand U11175 (N_11175,N_11090,N_11054);
nand U11176 (N_11176,N_11098,N_11053);
nor U11177 (N_11177,N_11026,N_11028);
and U11178 (N_11178,N_11027,N_11023);
nor U11179 (N_11179,N_11036,N_11103);
nor U11180 (N_11180,N_11016,N_11047);
nand U11181 (N_11181,N_11108,N_11004);
or U11182 (N_11182,N_11067,N_11070);
nor U11183 (N_11183,N_11032,N_11003);
xor U11184 (N_11184,N_11031,N_11035);
nand U11185 (N_11185,N_11065,N_11011);
xnor U11186 (N_11186,N_11085,N_11119);
nand U11187 (N_11187,N_11059,N_11063);
and U11188 (N_11188,N_11030,N_11065);
or U11189 (N_11189,N_11089,N_11081);
xnor U11190 (N_11190,N_11001,N_11072);
xnor U11191 (N_11191,N_11066,N_11123);
nor U11192 (N_11192,N_11012,N_11044);
and U11193 (N_11193,N_11038,N_11040);
xnor U11194 (N_11194,N_11015,N_11049);
xor U11195 (N_11195,N_11075,N_11041);
xor U11196 (N_11196,N_11002,N_11090);
nor U11197 (N_11197,N_11119,N_11026);
or U11198 (N_11198,N_11054,N_11043);
and U11199 (N_11199,N_11095,N_11015);
nor U11200 (N_11200,N_11070,N_11082);
or U11201 (N_11201,N_11100,N_11052);
xor U11202 (N_11202,N_11010,N_11033);
nor U11203 (N_11203,N_11082,N_11069);
nor U11204 (N_11204,N_11102,N_11066);
or U11205 (N_11205,N_11099,N_11055);
or U11206 (N_11206,N_11070,N_11105);
nor U11207 (N_11207,N_11074,N_11122);
nor U11208 (N_11208,N_11017,N_11081);
nor U11209 (N_11209,N_11120,N_11013);
nand U11210 (N_11210,N_11071,N_11111);
xor U11211 (N_11211,N_11090,N_11013);
or U11212 (N_11212,N_11050,N_11112);
and U11213 (N_11213,N_11036,N_11051);
xnor U11214 (N_11214,N_11044,N_11014);
xnor U11215 (N_11215,N_11058,N_11120);
nor U11216 (N_11216,N_11091,N_11065);
nand U11217 (N_11217,N_11069,N_11004);
and U11218 (N_11218,N_11029,N_11073);
nor U11219 (N_11219,N_11093,N_11085);
or U11220 (N_11220,N_11056,N_11033);
and U11221 (N_11221,N_11105,N_11060);
and U11222 (N_11222,N_11094,N_11061);
xnor U11223 (N_11223,N_11037,N_11074);
and U11224 (N_11224,N_11105,N_11082);
xor U11225 (N_11225,N_11069,N_11050);
xor U11226 (N_11226,N_11036,N_11118);
or U11227 (N_11227,N_11070,N_11004);
or U11228 (N_11228,N_11056,N_11043);
nand U11229 (N_11229,N_11097,N_11085);
xnor U11230 (N_11230,N_11025,N_11091);
or U11231 (N_11231,N_11079,N_11064);
or U11232 (N_11232,N_11026,N_11049);
or U11233 (N_11233,N_11033,N_11120);
and U11234 (N_11234,N_11025,N_11018);
nor U11235 (N_11235,N_11099,N_11006);
and U11236 (N_11236,N_11007,N_11098);
xnor U11237 (N_11237,N_11118,N_11015);
and U11238 (N_11238,N_11089,N_11096);
nor U11239 (N_11239,N_11022,N_11007);
nor U11240 (N_11240,N_11004,N_11013);
nor U11241 (N_11241,N_11048,N_11039);
nor U11242 (N_11242,N_11053,N_11059);
nand U11243 (N_11243,N_11050,N_11039);
or U11244 (N_11244,N_11082,N_11121);
or U11245 (N_11245,N_11020,N_11056);
nand U11246 (N_11246,N_11098,N_11063);
nor U11247 (N_11247,N_11104,N_11084);
and U11248 (N_11248,N_11066,N_11054);
and U11249 (N_11249,N_11017,N_11120);
nor U11250 (N_11250,N_11173,N_11242);
and U11251 (N_11251,N_11176,N_11142);
or U11252 (N_11252,N_11161,N_11240);
and U11253 (N_11253,N_11199,N_11196);
nor U11254 (N_11254,N_11146,N_11165);
nor U11255 (N_11255,N_11222,N_11206);
xor U11256 (N_11256,N_11220,N_11200);
or U11257 (N_11257,N_11227,N_11137);
and U11258 (N_11258,N_11214,N_11166);
or U11259 (N_11259,N_11186,N_11145);
and U11260 (N_11260,N_11225,N_11177);
nand U11261 (N_11261,N_11231,N_11131);
or U11262 (N_11262,N_11157,N_11204);
nand U11263 (N_11263,N_11128,N_11156);
nor U11264 (N_11264,N_11239,N_11217);
xnor U11265 (N_11265,N_11215,N_11153);
or U11266 (N_11266,N_11182,N_11144);
and U11267 (N_11267,N_11167,N_11202);
xor U11268 (N_11268,N_11174,N_11171);
xnor U11269 (N_11269,N_11183,N_11129);
or U11270 (N_11270,N_11152,N_11169);
and U11271 (N_11271,N_11226,N_11234);
or U11272 (N_11272,N_11224,N_11133);
and U11273 (N_11273,N_11198,N_11245);
xor U11274 (N_11274,N_11158,N_11243);
nor U11275 (N_11275,N_11249,N_11172);
nand U11276 (N_11276,N_11143,N_11185);
and U11277 (N_11277,N_11189,N_11135);
nor U11278 (N_11278,N_11208,N_11228);
and U11279 (N_11279,N_11162,N_11187);
or U11280 (N_11280,N_11188,N_11238);
and U11281 (N_11281,N_11211,N_11181);
xor U11282 (N_11282,N_11197,N_11125);
nor U11283 (N_11283,N_11221,N_11179);
nand U11284 (N_11284,N_11149,N_11164);
and U11285 (N_11285,N_11141,N_11194);
xor U11286 (N_11286,N_11232,N_11127);
nand U11287 (N_11287,N_11159,N_11233);
xor U11288 (N_11288,N_11190,N_11223);
or U11289 (N_11289,N_11184,N_11154);
xnor U11290 (N_11290,N_11136,N_11147);
and U11291 (N_11291,N_11175,N_11193);
xnor U11292 (N_11292,N_11140,N_11168);
xor U11293 (N_11293,N_11148,N_11218);
nor U11294 (N_11294,N_11241,N_11212);
and U11295 (N_11295,N_11195,N_11138);
or U11296 (N_11296,N_11229,N_11192);
xor U11297 (N_11297,N_11151,N_11237);
nor U11298 (N_11298,N_11247,N_11248);
or U11299 (N_11299,N_11244,N_11210);
nor U11300 (N_11300,N_11180,N_11139);
nor U11301 (N_11301,N_11201,N_11205);
xor U11302 (N_11302,N_11126,N_11203);
nand U11303 (N_11303,N_11130,N_11246);
or U11304 (N_11304,N_11219,N_11209);
and U11305 (N_11305,N_11170,N_11150);
or U11306 (N_11306,N_11132,N_11236);
nand U11307 (N_11307,N_11230,N_11134);
nand U11308 (N_11308,N_11178,N_11160);
nor U11309 (N_11309,N_11207,N_11155);
and U11310 (N_11310,N_11216,N_11235);
or U11311 (N_11311,N_11163,N_11213);
xnor U11312 (N_11312,N_11191,N_11176);
or U11313 (N_11313,N_11247,N_11234);
nor U11314 (N_11314,N_11125,N_11173);
or U11315 (N_11315,N_11211,N_11130);
xor U11316 (N_11316,N_11195,N_11143);
nand U11317 (N_11317,N_11125,N_11151);
nor U11318 (N_11318,N_11217,N_11169);
xnor U11319 (N_11319,N_11138,N_11140);
and U11320 (N_11320,N_11154,N_11221);
xor U11321 (N_11321,N_11148,N_11151);
nand U11322 (N_11322,N_11132,N_11189);
nor U11323 (N_11323,N_11167,N_11162);
xor U11324 (N_11324,N_11176,N_11217);
or U11325 (N_11325,N_11193,N_11170);
xor U11326 (N_11326,N_11181,N_11127);
nand U11327 (N_11327,N_11221,N_11208);
nor U11328 (N_11328,N_11243,N_11163);
nand U11329 (N_11329,N_11159,N_11200);
xnor U11330 (N_11330,N_11237,N_11172);
and U11331 (N_11331,N_11187,N_11248);
and U11332 (N_11332,N_11245,N_11247);
or U11333 (N_11333,N_11219,N_11176);
xor U11334 (N_11334,N_11176,N_11229);
or U11335 (N_11335,N_11188,N_11183);
and U11336 (N_11336,N_11164,N_11202);
nor U11337 (N_11337,N_11153,N_11136);
xnor U11338 (N_11338,N_11230,N_11209);
and U11339 (N_11339,N_11148,N_11128);
nor U11340 (N_11340,N_11171,N_11137);
nand U11341 (N_11341,N_11221,N_11240);
nor U11342 (N_11342,N_11139,N_11202);
or U11343 (N_11343,N_11176,N_11137);
nand U11344 (N_11344,N_11193,N_11249);
nor U11345 (N_11345,N_11179,N_11249);
or U11346 (N_11346,N_11142,N_11136);
or U11347 (N_11347,N_11152,N_11165);
or U11348 (N_11348,N_11188,N_11218);
and U11349 (N_11349,N_11243,N_11145);
or U11350 (N_11350,N_11210,N_11145);
xor U11351 (N_11351,N_11162,N_11211);
nand U11352 (N_11352,N_11246,N_11146);
or U11353 (N_11353,N_11221,N_11239);
and U11354 (N_11354,N_11127,N_11221);
xor U11355 (N_11355,N_11150,N_11198);
nor U11356 (N_11356,N_11174,N_11240);
nand U11357 (N_11357,N_11233,N_11171);
nor U11358 (N_11358,N_11181,N_11247);
nor U11359 (N_11359,N_11161,N_11204);
nand U11360 (N_11360,N_11209,N_11142);
and U11361 (N_11361,N_11220,N_11163);
or U11362 (N_11362,N_11144,N_11151);
or U11363 (N_11363,N_11227,N_11165);
or U11364 (N_11364,N_11249,N_11145);
nor U11365 (N_11365,N_11146,N_11173);
nor U11366 (N_11366,N_11174,N_11128);
and U11367 (N_11367,N_11133,N_11195);
nor U11368 (N_11368,N_11164,N_11179);
nand U11369 (N_11369,N_11149,N_11180);
nand U11370 (N_11370,N_11159,N_11190);
or U11371 (N_11371,N_11137,N_11177);
nor U11372 (N_11372,N_11215,N_11192);
nand U11373 (N_11373,N_11201,N_11181);
xnor U11374 (N_11374,N_11209,N_11196);
nor U11375 (N_11375,N_11346,N_11326);
nor U11376 (N_11376,N_11337,N_11350);
xnor U11377 (N_11377,N_11256,N_11266);
xor U11378 (N_11378,N_11289,N_11345);
or U11379 (N_11379,N_11349,N_11300);
nand U11380 (N_11380,N_11364,N_11282);
nor U11381 (N_11381,N_11374,N_11369);
xor U11382 (N_11382,N_11361,N_11293);
nor U11383 (N_11383,N_11268,N_11275);
xnor U11384 (N_11384,N_11331,N_11270);
nor U11385 (N_11385,N_11355,N_11291);
and U11386 (N_11386,N_11296,N_11366);
and U11387 (N_11387,N_11318,N_11323);
and U11388 (N_11388,N_11278,N_11359);
xnor U11389 (N_11389,N_11299,N_11258);
nand U11390 (N_11390,N_11303,N_11322);
or U11391 (N_11391,N_11252,N_11265);
and U11392 (N_11392,N_11339,N_11314);
nand U11393 (N_11393,N_11288,N_11274);
nand U11394 (N_11394,N_11301,N_11295);
xnor U11395 (N_11395,N_11363,N_11372);
or U11396 (N_11396,N_11332,N_11281);
or U11397 (N_11397,N_11351,N_11271);
nor U11398 (N_11398,N_11340,N_11316);
or U11399 (N_11399,N_11327,N_11294);
nor U11400 (N_11400,N_11264,N_11255);
or U11401 (N_11401,N_11324,N_11259);
nand U11402 (N_11402,N_11360,N_11309);
and U11403 (N_11403,N_11261,N_11357);
nand U11404 (N_11404,N_11283,N_11253);
nand U11405 (N_11405,N_11335,N_11329);
and U11406 (N_11406,N_11352,N_11371);
nand U11407 (N_11407,N_11305,N_11373);
xor U11408 (N_11408,N_11347,N_11312);
or U11409 (N_11409,N_11260,N_11272);
and U11410 (N_11410,N_11358,N_11273);
and U11411 (N_11411,N_11353,N_11280);
xor U11412 (N_11412,N_11298,N_11263);
or U11413 (N_11413,N_11356,N_11365);
and U11414 (N_11414,N_11284,N_11267);
and U11415 (N_11415,N_11367,N_11308);
and U11416 (N_11416,N_11251,N_11343);
and U11417 (N_11417,N_11320,N_11315);
or U11418 (N_11418,N_11286,N_11342);
nor U11419 (N_11419,N_11344,N_11341);
nand U11420 (N_11420,N_11317,N_11338);
or U11421 (N_11421,N_11333,N_11262);
or U11422 (N_11422,N_11348,N_11370);
and U11423 (N_11423,N_11257,N_11354);
or U11424 (N_11424,N_11330,N_11310);
and U11425 (N_11425,N_11368,N_11292);
and U11426 (N_11426,N_11313,N_11325);
xor U11427 (N_11427,N_11287,N_11306);
xnor U11428 (N_11428,N_11307,N_11254);
and U11429 (N_11429,N_11279,N_11269);
and U11430 (N_11430,N_11334,N_11321);
nand U11431 (N_11431,N_11250,N_11311);
nand U11432 (N_11432,N_11362,N_11290);
nor U11433 (N_11433,N_11285,N_11302);
nor U11434 (N_11434,N_11276,N_11336);
and U11435 (N_11435,N_11328,N_11319);
and U11436 (N_11436,N_11277,N_11304);
or U11437 (N_11437,N_11297,N_11360);
nor U11438 (N_11438,N_11317,N_11277);
nand U11439 (N_11439,N_11344,N_11342);
xor U11440 (N_11440,N_11257,N_11373);
xnor U11441 (N_11441,N_11341,N_11323);
and U11442 (N_11442,N_11275,N_11307);
and U11443 (N_11443,N_11351,N_11363);
and U11444 (N_11444,N_11337,N_11324);
or U11445 (N_11445,N_11260,N_11318);
nand U11446 (N_11446,N_11315,N_11362);
xor U11447 (N_11447,N_11304,N_11351);
xor U11448 (N_11448,N_11321,N_11347);
nand U11449 (N_11449,N_11271,N_11302);
or U11450 (N_11450,N_11364,N_11346);
nand U11451 (N_11451,N_11288,N_11280);
and U11452 (N_11452,N_11341,N_11307);
nand U11453 (N_11453,N_11345,N_11352);
and U11454 (N_11454,N_11319,N_11371);
or U11455 (N_11455,N_11345,N_11306);
nor U11456 (N_11456,N_11327,N_11356);
nand U11457 (N_11457,N_11314,N_11328);
or U11458 (N_11458,N_11348,N_11343);
xor U11459 (N_11459,N_11353,N_11261);
or U11460 (N_11460,N_11254,N_11333);
or U11461 (N_11461,N_11255,N_11334);
nor U11462 (N_11462,N_11281,N_11306);
nand U11463 (N_11463,N_11355,N_11251);
and U11464 (N_11464,N_11369,N_11332);
nor U11465 (N_11465,N_11318,N_11370);
xnor U11466 (N_11466,N_11250,N_11296);
xnor U11467 (N_11467,N_11280,N_11373);
xor U11468 (N_11468,N_11262,N_11307);
or U11469 (N_11469,N_11251,N_11331);
xor U11470 (N_11470,N_11357,N_11373);
nand U11471 (N_11471,N_11259,N_11250);
xor U11472 (N_11472,N_11319,N_11348);
or U11473 (N_11473,N_11266,N_11296);
and U11474 (N_11474,N_11339,N_11313);
xor U11475 (N_11475,N_11293,N_11349);
nor U11476 (N_11476,N_11329,N_11365);
and U11477 (N_11477,N_11255,N_11369);
or U11478 (N_11478,N_11293,N_11276);
xnor U11479 (N_11479,N_11272,N_11309);
nand U11480 (N_11480,N_11252,N_11259);
or U11481 (N_11481,N_11300,N_11273);
nor U11482 (N_11482,N_11312,N_11309);
or U11483 (N_11483,N_11371,N_11264);
or U11484 (N_11484,N_11260,N_11363);
nor U11485 (N_11485,N_11371,N_11344);
xor U11486 (N_11486,N_11273,N_11363);
or U11487 (N_11487,N_11347,N_11262);
nor U11488 (N_11488,N_11323,N_11369);
and U11489 (N_11489,N_11358,N_11270);
xor U11490 (N_11490,N_11291,N_11362);
or U11491 (N_11491,N_11268,N_11286);
nand U11492 (N_11492,N_11315,N_11371);
xnor U11493 (N_11493,N_11306,N_11324);
and U11494 (N_11494,N_11273,N_11357);
nor U11495 (N_11495,N_11259,N_11374);
nand U11496 (N_11496,N_11349,N_11259);
nand U11497 (N_11497,N_11347,N_11287);
and U11498 (N_11498,N_11267,N_11256);
nor U11499 (N_11499,N_11261,N_11254);
and U11500 (N_11500,N_11489,N_11478);
nand U11501 (N_11501,N_11438,N_11417);
and U11502 (N_11502,N_11496,N_11389);
nor U11503 (N_11503,N_11451,N_11492);
nor U11504 (N_11504,N_11416,N_11409);
xor U11505 (N_11505,N_11406,N_11441);
xnor U11506 (N_11506,N_11493,N_11475);
or U11507 (N_11507,N_11399,N_11485);
nand U11508 (N_11508,N_11402,N_11379);
nor U11509 (N_11509,N_11463,N_11425);
nand U11510 (N_11510,N_11408,N_11488);
xor U11511 (N_11511,N_11486,N_11386);
or U11512 (N_11512,N_11384,N_11445);
or U11513 (N_11513,N_11482,N_11419);
nand U11514 (N_11514,N_11387,N_11413);
nor U11515 (N_11515,N_11397,N_11465);
xor U11516 (N_11516,N_11472,N_11467);
or U11517 (N_11517,N_11455,N_11381);
nand U11518 (N_11518,N_11490,N_11412);
or U11519 (N_11519,N_11498,N_11460);
xor U11520 (N_11520,N_11418,N_11375);
and U11521 (N_11521,N_11423,N_11434);
or U11522 (N_11522,N_11380,N_11414);
nand U11523 (N_11523,N_11483,N_11477);
and U11524 (N_11524,N_11470,N_11440);
nor U11525 (N_11525,N_11476,N_11428);
and U11526 (N_11526,N_11433,N_11429);
and U11527 (N_11527,N_11459,N_11466);
nand U11528 (N_11528,N_11405,N_11401);
nor U11529 (N_11529,N_11422,N_11450);
and U11530 (N_11530,N_11411,N_11396);
nor U11531 (N_11531,N_11437,N_11468);
and U11532 (N_11532,N_11446,N_11439);
nand U11533 (N_11533,N_11407,N_11479);
and U11534 (N_11534,N_11473,N_11453);
xor U11535 (N_11535,N_11448,N_11432);
nand U11536 (N_11536,N_11435,N_11400);
and U11537 (N_11537,N_11377,N_11457);
nand U11538 (N_11538,N_11464,N_11388);
and U11539 (N_11539,N_11447,N_11394);
and U11540 (N_11540,N_11452,N_11499);
or U11541 (N_11541,N_11383,N_11491);
xnor U11542 (N_11542,N_11436,N_11385);
nand U11543 (N_11543,N_11481,N_11430);
nand U11544 (N_11544,N_11420,N_11426);
or U11545 (N_11545,N_11393,N_11462);
nor U11546 (N_11546,N_11487,N_11398);
and U11547 (N_11547,N_11495,N_11442);
xor U11548 (N_11548,N_11421,N_11390);
or U11549 (N_11549,N_11403,N_11449);
nand U11550 (N_11550,N_11484,N_11461);
nand U11551 (N_11551,N_11469,N_11454);
and U11552 (N_11552,N_11474,N_11376);
or U11553 (N_11553,N_11391,N_11410);
nor U11554 (N_11554,N_11392,N_11480);
or U11555 (N_11555,N_11424,N_11471);
and U11556 (N_11556,N_11444,N_11404);
xor U11557 (N_11557,N_11458,N_11415);
or U11558 (N_11558,N_11456,N_11427);
nor U11559 (N_11559,N_11382,N_11378);
nor U11560 (N_11560,N_11431,N_11395);
and U11561 (N_11561,N_11494,N_11497);
nor U11562 (N_11562,N_11443,N_11422);
or U11563 (N_11563,N_11425,N_11478);
and U11564 (N_11564,N_11449,N_11457);
nand U11565 (N_11565,N_11386,N_11452);
and U11566 (N_11566,N_11492,N_11486);
nor U11567 (N_11567,N_11440,N_11424);
nor U11568 (N_11568,N_11423,N_11435);
nor U11569 (N_11569,N_11492,N_11376);
or U11570 (N_11570,N_11377,N_11496);
or U11571 (N_11571,N_11423,N_11432);
nand U11572 (N_11572,N_11447,N_11468);
nor U11573 (N_11573,N_11379,N_11496);
nor U11574 (N_11574,N_11396,N_11444);
nand U11575 (N_11575,N_11461,N_11439);
xor U11576 (N_11576,N_11393,N_11440);
and U11577 (N_11577,N_11428,N_11483);
nand U11578 (N_11578,N_11433,N_11389);
nand U11579 (N_11579,N_11400,N_11467);
and U11580 (N_11580,N_11462,N_11407);
nand U11581 (N_11581,N_11480,N_11442);
xor U11582 (N_11582,N_11393,N_11411);
nor U11583 (N_11583,N_11413,N_11442);
xor U11584 (N_11584,N_11441,N_11382);
xor U11585 (N_11585,N_11475,N_11376);
or U11586 (N_11586,N_11453,N_11399);
or U11587 (N_11587,N_11383,N_11415);
nand U11588 (N_11588,N_11467,N_11431);
and U11589 (N_11589,N_11430,N_11393);
or U11590 (N_11590,N_11404,N_11470);
and U11591 (N_11591,N_11460,N_11401);
xnor U11592 (N_11592,N_11440,N_11467);
or U11593 (N_11593,N_11474,N_11408);
nor U11594 (N_11594,N_11495,N_11466);
and U11595 (N_11595,N_11404,N_11423);
xor U11596 (N_11596,N_11392,N_11494);
or U11597 (N_11597,N_11498,N_11447);
and U11598 (N_11598,N_11451,N_11488);
and U11599 (N_11599,N_11489,N_11426);
or U11600 (N_11600,N_11424,N_11378);
or U11601 (N_11601,N_11382,N_11495);
nor U11602 (N_11602,N_11393,N_11410);
and U11603 (N_11603,N_11379,N_11457);
or U11604 (N_11604,N_11418,N_11435);
nor U11605 (N_11605,N_11430,N_11405);
xnor U11606 (N_11606,N_11460,N_11461);
and U11607 (N_11607,N_11403,N_11467);
nand U11608 (N_11608,N_11382,N_11435);
nor U11609 (N_11609,N_11402,N_11381);
and U11610 (N_11610,N_11389,N_11455);
xor U11611 (N_11611,N_11416,N_11402);
xnor U11612 (N_11612,N_11432,N_11445);
nand U11613 (N_11613,N_11438,N_11497);
nand U11614 (N_11614,N_11419,N_11472);
nor U11615 (N_11615,N_11484,N_11402);
or U11616 (N_11616,N_11488,N_11498);
nor U11617 (N_11617,N_11453,N_11380);
or U11618 (N_11618,N_11471,N_11394);
nand U11619 (N_11619,N_11450,N_11377);
nand U11620 (N_11620,N_11480,N_11395);
and U11621 (N_11621,N_11383,N_11419);
nor U11622 (N_11622,N_11390,N_11467);
and U11623 (N_11623,N_11442,N_11468);
xnor U11624 (N_11624,N_11382,N_11496);
and U11625 (N_11625,N_11622,N_11567);
nand U11626 (N_11626,N_11624,N_11511);
and U11627 (N_11627,N_11584,N_11514);
nor U11628 (N_11628,N_11534,N_11519);
or U11629 (N_11629,N_11556,N_11557);
or U11630 (N_11630,N_11616,N_11528);
nand U11631 (N_11631,N_11621,N_11599);
and U11632 (N_11632,N_11532,N_11503);
and U11633 (N_11633,N_11571,N_11613);
xor U11634 (N_11634,N_11538,N_11588);
or U11635 (N_11635,N_11541,N_11506);
and U11636 (N_11636,N_11510,N_11573);
and U11637 (N_11637,N_11515,N_11546);
nand U11638 (N_11638,N_11596,N_11590);
nand U11639 (N_11639,N_11531,N_11592);
nor U11640 (N_11640,N_11582,N_11605);
or U11641 (N_11641,N_11524,N_11566);
or U11642 (N_11642,N_11558,N_11600);
and U11643 (N_11643,N_11518,N_11550);
or U11644 (N_11644,N_11521,N_11562);
and U11645 (N_11645,N_11620,N_11598);
xor U11646 (N_11646,N_11509,N_11607);
and U11647 (N_11647,N_11522,N_11569);
nand U11648 (N_11648,N_11504,N_11568);
and U11649 (N_11649,N_11505,N_11577);
or U11650 (N_11650,N_11500,N_11610);
or U11651 (N_11651,N_11554,N_11570);
nand U11652 (N_11652,N_11594,N_11580);
nand U11653 (N_11653,N_11533,N_11561);
or U11654 (N_11654,N_11555,N_11537);
xnor U11655 (N_11655,N_11603,N_11508);
or U11656 (N_11656,N_11530,N_11543);
or U11657 (N_11657,N_11606,N_11576);
nand U11658 (N_11658,N_11560,N_11523);
nand U11659 (N_11659,N_11617,N_11611);
nor U11660 (N_11660,N_11585,N_11615);
xnor U11661 (N_11661,N_11589,N_11597);
nor U11662 (N_11662,N_11618,N_11608);
nor U11663 (N_11663,N_11525,N_11540);
nand U11664 (N_11664,N_11512,N_11623);
or U11665 (N_11665,N_11578,N_11549);
xnor U11666 (N_11666,N_11583,N_11553);
or U11667 (N_11667,N_11551,N_11609);
or U11668 (N_11668,N_11574,N_11536);
and U11669 (N_11669,N_11563,N_11595);
xor U11670 (N_11670,N_11565,N_11507);
and U11671 (N_11671,N_11591,N_11619);
nor U11672 (N_11672,N_11593,N_11564);
nand U11673 (N_11673,N_11513,N_11545);
nor U11674 (N_11674,N_11516,N_11601);
and U11675 (N_11675,N_11575,N_11602);
xnor U11676 (N_11676,N_11527,N_11502);
and U11677 (N_11677,N_11526,N_11559);
or U11678 (N_11678,N_11501,N_11520);
nor U11679 (N_11679,N_11529,N_11548);
and U11680 (N_11680,N_11604,N_11586);
nand U11681 (N_11681,N_11552,N_11572);
xor U11682 (N_11682,N_11614,N_11547);
and U11683 (N_11683,N_11544,N_11579);
or U11684 (N_11684,N_11517,N_11535);
and U11685 (N_11685,N_11539,N_11581);
nor U11686 (N_11686,N_11612,N_11542);
and U11687 (N_11687,N_11587,N_11526);
or U11688 (N_11688,N_11563,N_11503);
nand U11689 (N_11689,N_11571,N_11504);
or U11690 (N_11690,N_11529,N_11593);
and U11691 (N_11691,N_11619,N_11579);
xnor U11692 (N_11692,N_11601,N_11567);
or U11693 (N_11693,N_11617,N_11526);
or U11694 (N_11694,N_11517,N_11556);
nor U11695 (N_11695,N_11534,N_11597);
nand U11696 (N_11696,N_11616,N_11534);
or U11697 (N_11697,N_11516,N_11517);
and U11698 (N_11698,N_11612,N_11508);
and U11699 (N_11699,N_11544,N_11554);
nand U11700 (N_11700,N_11578,N_11506);
and U11701 (N_11701,N_11545,N_11598);
xnor U11702 (N_11702,N_11586,N_11591);
and U11703 (N_11703,N_11511,N_11532);
nor U11704 (N_11704,N_11595,N_11593);
nand U11705 (N_11705,N_11598,N_11581);
or U11706 (N_11706,N_11526,N_11607);
nand U11707 (N_11707,N_11537,N_11543);
and U11708 (N_11708,N_11560,N_11598);
xor U11709 (N_11709,N_11511,N_11573);
nand U11710 (N_11710,N_11555,N_11609);
nor U11711 (N_11711,N_11578,N_11624);
or U11712 (N_11712,N_11506,N_11607);
or U11713 (N_11713,N_11531,N_11527);
or U11714 (N_11714,N_11546,N_11557);
nand U11715 (N_11715,N_11589,N_11514);
xor U11716 (N_11716,N_11597,N_11554);
or U11717 (N_11717,N_11617,N_11536);
xor U11718 (N_11718,N_11512,N_11542);
and U11719 (N_11719,N_11612,N_11557);
xnor U11720 (N_11720,N_11514,N_11577);
xor U11721 (N_11721,N_11593,N_11555);
nand U11722 (N_11722,N_11503,N_11500);
nor U11723 (N_11723,N_11533,N_11538);
nor U11724 (N_11724,N_11622,N_11605);
and U11725 (N_11725,N_11510,N_11602);
or U11726 (N_11726,N_11615,N_11588);
and U11727 (N_11727,N_11596,N_11526);
nor U11728 (N_11728,N_11595,N_11509);
nand U11729 (N_11729,N_11618,N_11539);
nor U11730 (N_11730,N_11547,N_11506);
nor U11731 (N_11731,N_11528,N_11561);
or U11732 (N_11732,N_11615,N_11597);
or U11733 (N_11733,N_11520,N_11549);
nor U11734 (N_11734,N_11595,N_11562);
and U11735 (N_11735,N_11610,N_11609);
nand U11736 (N_11736,N_11530,N_11560);
nor U11737 (N_11737,N_11612,N_11528);
and U11738 (N_11738,N_11624,N_11569);
or U11739 (N_11739,N_11611,N_11524);
nand U11740 (N_11740,N_11582,N_11530);
nor U11741 (N_11741,N_11514,N_11527);
nand U11742 (N_11742,N_11515,N_11519);
xor U11743 (N_11743,N_11623,N_11588);
xnor U11744 (N_11744,N_11612,N_11554);
nor U11745 (N_11745,N_11526,N_11528);
or U11746 (N_11746,N_11541,N_11510);
or U11747 (N_11747,N_11524,N_11519);
nand U11748 (N_11748,N_11596,N_11530);
and U11749 (N_11749,N_11612,N_11539);
nand U11750 (N_11750,N_11693,N_11648);
or U11751 (N_11751,N_11656,N_11729);
nor U11752 (N_11752,N_11631,N_11639);
nand U11753 (N_11753,N_11646,N_11735);
and U11754 (N_11754,N_11625,N_11722);
or U11755 (N_11755,N_11691,N_11653);
nor U11756 (N_11756,N_11685,N_11634);
nand U11757 (N_11757,N_11642,N_11740);
nand U11758 (N_11758,N_11700,N_11724);
and U11759 (N_11759,N_11738,N_11660);
nor U11760 (N_11760,N_11629,N_11661);
or U11761 (N_11761,N_11652,N_11665);
xor U11762 (N_11762,N_11657,N_11718);
and U11763 (N_11763,N_11702,N_11650);
nand U11764 (N_11764,N_11737,N_11694);
nor U11765 (N_11765,N_11635,N_11739);
nor U11766 (N_11766,N_11743,N_11644);
nor U11767 (N_11767,N_11711,N_11721);
nor U11768 (N_11768,N_11728,N_11730);
nor U11769 (N_11769,N_11626,N_11632);
and U11770 (N_11770,N_11734,N_11697);
or U11771 (N_11771,N_11704,N_11643);
or U11772 (N_11772,N_11637,N_11667);
xor U11773 (N_11773,N_11719,N_11720);
or U11774 (N_11774,N_11723,N_11659);
xor U11775 (N_11775,N_11678,N_11692);
nand U11776 (N_11776,N_11688,N_11628);
or U11777 (N_11777,N_11682,N_11749);
and U11778 (N_11778,N_11669,N_11705);
xnor U11779 (N_11779,N_11649,N_11706);
nand U11780 (N_11780,N_11636,N_11683);
nor U11781 (N_11781,N_11741,N_11714);
nand U11782 (N_11782,N_11630,N_11673);
nor U11783 (N_11783,N_11712,N_11675);
nor U11784 (N_11784,N_11703,N_11726);
and U11785 (N_11785,N_11654,N_11696);
xor U11786 (N_11786,N_11658,N_11745);
nor U11787 (N_11787,N_11717,N_11736);
or U11788 (N_11788,N_11746,N_11641);
nand U11789 (N_11789,N_11684,N_11689);
nand U11790 (N_11790,N_11679,N_11645);
or U11791 (N_11791,N_11742,N_11701);
nand U11792 (N_11792,N_11677,N_11709);
nand U11793 (N_11793,N_11690,N_11671);
xnor U11794 (N_11794,N_11664,N_11686);
xor U11795 (N_11795,N_11699,N_11713);
xor U11796 (N_11796,N_11708,N_11676);
xnor U11797 (N_11797,N_11662,N_11674);
or U11798 (N_11798,N_11668,N_11651);
or U11799 (N_11799,N_11627,N_11716);
and U11800 (N_11800,N_11698,N_11681);
xor U11801 (N_11801,N_11672,N_11666);
and U11802 (N_11802,N_11695,N_11732);
and U11803 (N_11803,N_11663,N_11655);
nand U11804 (N_11804,N_11733,N_11731);
nor U11805 (N_11805,N_11727,N_11748);
or U11806 (N_11806,N_11680,N_11715);
xnor U11807 (N_11807,N_11638,N_11633);
nor U11808 (N_11808,N_11710,N_11744);
xor U11809 (N_11809,N_11725,N_11640);
xor U11810 (N_11810,N_11687,N_11747);
or U11811 (N_11811,N_11670,N_11707);
and U11812 (N_11812,N_11647,N_11738);
or U11813 (N_11813,N_11704,N_11731);
and U11814 (N_11814,N_11704,N_11721);
and U11815 (N_11815,N_11628,N_11705);
and U11816 (N_11816,N_11674,N_11638);
nor U11817 (N_11817,N_11663,N_11708);
or U11818 (N_11818,N_11647,N_11675);
nand U11819 (N_11819,N_11654,N_11672);
nor U11820 (N_11820,N_11734,N_11684);
nor U11821 (N_11821,N_11709,N_11726);
nor U11822 (N_11822,N_11677,N_11640);
or U11823 (N_11823,N_11712,N_11651);
nor U11824 (N_11824,N_11727,N_11655);
or U11825 (N_11825,N_11730,N_11690);
and U11826 (N_11826,N_11739,N_11661);
and U11827 (N_11827,N_11742,N_11645);
and U11828 (N_11828,N_11747,N_11742);
or U11829 (N_11829,N_11665,N_11668);
or U11830 (N_11830,N_11704,N_11709);
nor U11831 (N_11831,N_11628,N_11749);
and U11832 (N_11832,N_11696,N_11722);
and U11833 (N_11833,N_11695,N_11726);
nor U11834 (N_11834,N_11633,N_11697);
or U11835 (N_11835,N_11693,N_11729);
or U11836 (N_11836,N_11674,N_11627);
nand U11837 (N_11837,N_11737,N_11687);
xnor U11838 (N_11838,N_11634,N_11645);
nand U11839 (N_11839,N_11651,N_11721);
xnor U11840 (N_11840,N_11740,N_11720);
nand U11841 (N_11841,N_11705,N_11666);
and U11842 (N_11842,N_11669,N_11702);
nor U11843 (N_11843,N_11660,N_11730);
and U11844 (N_11844,N_11711,N_11733);
and U11845 (N_11845,N_11698,N_11737);
nand U11846 (N_11846,N_11742,N_11697);
nand U11847 (N_11847,N_11633,N_11635);
nand U11848 (N_11848,N_11684,N_11741);
nand U11849 (N_11849,N_11703,N_11638);
nand U11850 (N_11850,N_11657,N_11685);
xor U11851 (N_11851,N_11702,N_11654);
nor U11852 (N_11852,N_11633,N_11708);
nand U11853 (N_11853,N_11632,N_11636);
nor U11854 (N_11854,N_11672,N_11690);
nand U11855 (N_11855,N_11688,N_11708);
xnor U11856 (N_11856,N_11739,N_11667);
xnor U11857 (N_11857,N_11713,N_11660);
nand U11858 (N_11858,N_11645,N_11662);
nand U11859 (N_11859,N_11692,N_11705);
and U11860 (N_11860,N_11718,N_11665);
xnor U11861 (N_11861,N_11629,N_11651);
nand U11862 (N_11862,N_11629,N_11736);
or U11863 (N_11863,N_11695,N_11640);
nor U11864 (N_11864,N_11712,N_11738);
xnor U11865 (N_11865,N_11741,N_11721);
and U11866 (N_11866,N_11669,N_11714);
nand U11867 (N_11867,N_11732,N_11728);
nor U11868 (N_11868,N_11631,N_11727);
xnor U11869 (N_11869,N_11748,N_11632);
nor U11870 (N_11870,N_11689,N_11683);
or U11871 (N_11871,N_11638,N_11715);
xnor U11872 (N_11872,N_11715,N_11667);
or U11873 (N_11873,N_11638,N_11650);
nor U11874 (N_11874,N_11697,N_11646);
or U11875 (N_11875,N_11750,N_11753);
nor U11876 (N_11876,N_11777,N_11751);
nor U11877 (N_11877,N_11773,N_11785);
and U11878 (N_11878,N_11841,N_11772);
nand U11879 (N_11879,N_11808,N_11783);
or U11880 (N_11880,N_11782,N_11761);
or U11881 (N_11881,N_11813,N_11788);
nor U11882 (N_11882,N_11752,N_11871);
xor U11883 (N_11883,N_11860,N_11812);
and U11884 (N_11884,N_11818,N_11817);
or U11885 (N_11885,N_11865,N_11791);
and U11886 (N_11886,N_11795,N_11846);
and U11887 (N_11887,N_11819,N_11854);
xor U11888 (N_11888,N_11779,N_11815);
xor U11889 (N_11889,N_11873,N_11814);
nand U11890 (N_11890,N_11840,N_11835);
nor U11891 (N_11891,N_11760,N_11759);
and U11892 (N_11892,N_11831,N_11862);
and U11893 (N_11893,N_11857,N_11825);
or U11894 (N_11894,N_11863,N_11789);
or U11895 (N_11895,N_11836,N_11799);
or U11896 (N_11896,N_11855,N_11784);
and U11897 (N_11897,N_11832,N_11816);
and U11898 (N_11898,N_11792,N_11866);
or U11899 (N_11899,N_11858,N_11872);
and U11900 (N_11900,N_11771,N_11765);
and U11901 (N_11901,N_11847,N_11829);
nor U11902 (N_11902,N_11770,N_11806);
or U11903 (N_11903,N_11793,N_11804);
or U11904 (N_11904,N_11767,N_11837);
and U11905 (N_11905,N_11868,N_11798);
or U11906 (N_11906,N_11820,N_11762);
and U11907 (N_11907,N_11787,N_11823);
nor U11908 (N_11908,N_11833,N_11756);
nor U11909 (N_11909,N_11850,N_11822);
and U11910 (N_11910,N_11828,N_11802);
and U11911 (N_11911,N_11859,N_11811);
or U11912 (N_11912,N_11797,N_11800);
nor U11913 (N_11913,N_11769,N_11834);
and U11914 (N_11914,N_11775,N_11774);
and U11915 (N_11915,N_11830,N_11839);
nor U11916 (N_11916,N_11870,N_11807);
nand U11917 (N_11917,N_11826,N_11848);
and U11918 (N_11918,N_11796,N_11764);
and U11919 (N_11919,N_11809,N_11778);
or U11920 (N_11920,N_11845,N_11824);
and U11921 (N_11921,N_11786,N_11766);
nand U11922 (N_11922,N_11852,N_11763);
xnor U11923 (N_11923,N_11849,N_11758);
or U11924 (N_11924,N_11851,N_11821);
nand U11925 (N_11925,N_11781,N_11803);
nand U11926 (N_11926,N_11864,N_11776);
and U11927 (N_11927,N_11827,N_11843);
and U11928 (N_11928,N_11754,N_11853);
and U11929 (N_11929,N_11874,N_11861);
and U11930 (N_11930,N_11869,N_11842);
and U11931 (N_11931,N_11790,N_11780);
nor U11932 (N_11932,N_11810,N_11801);
nand U11933 (N_11933,N_11838,N_11805);
and U11934 (N_11934,N_11768,N_11856);
nor U11935 (N_11935,N_11755,N_11867);
and U11936 (N_11936,N_11794,N_11844);
and U11937 (N_11937,N_11757,N_11805);
or U11938 (N_11938,N_11792,N_11805);
xor U11939 (N_11939,N_11857,N_11759);
and U11940 (N_11940,N_11764,N_11777);
and U11941 (N_11941,N_11787,N_11806);
and U11942 (N_11942,N_11868,N_11767);
and U11943 (N_11943,N_11865,N_11867);
nand U11944 (N_11944,N_11860,N_11849);
nor U11945 (N_11945,N_11776,N_11764);
xor U11946 (N_11946,N_11851,N_11847);
or U11947 (N_11947,N_11823,N_11764);
xor U11948 (N_11948,N_11794,N_11857);
xor U11949 (N_11949,N_11780,N_11758);
nor U11950 (N_11950,N_11776,N_11837);
and U11951 (N_11951,N_11824,N_11865);
nor U11952 (N_11952,N_11830,N_11859);
xor U11953 (N_11953,N_11857,N_11784);
and U11954 (N_11954,N_11802,N_11766);
nor U11955 (N_11955,N_11787,N_11834);
nor U11956 (N_11956,N_11797,N_11815);
nand U11957 (N_11957,N_11822,N_11849);
nor U11958 (N_11958,N_11801,N_11857);
xor U11959 (N_11959,N_11832,N_11865);
nand U11960 (N_11960,N_11860,N_11764);
nor U11961 (N_11961,N_11857,N_11803);
xor U11962 (N_11962,N_11769,N_11812);
nor U11963 (N_11963,N_11846,N_11806);
and U11964 (N_11964,N_11848,N_11847);
nand U11965 (N_11965,N_11763,N_11813);
and U11966 (N_11966,N_11831,N_11797);
nor U11967 (N_11967,N_11781,N_11824);
nand U11968 (N_11968,N_11847,N_11806);
or U11969 (N_11969,N_11862,N_11772);
or U11970 (N_11970,N_11839,N_11766);
nand U11971 (N_11971,N_11835,N_11845);
or U11972 (N_11972,N_11798,N_11810);
nor U11973 (N_11973,N_11799,N_11869);
xnor U11974 (N_11974,N_11764,N_11766);
nand U11975 (N_11975,N_11757,N_11833);
xor U11976 (N_11976,N_11788,N_11771);
and U11977 (N_11977,N_11792,N_11809);
xnor U11978 (N_11978,N_11834,N_11843);
nand U11979 (N_11979,N_11779,N_11794);
or U11980 (N_11980,N_11780,N_11769);
nor U11981 (N_11981,N_11840,N_11830);
xnor U11982 (N_11982,N_11832,N_11796);
nand U11983 (N_11983,N_11861,N_11782);
nor U11984 (N_11984,N_11850,N_11858);
or U11985 (N_11985,N_11805,N_11839);
nand U11986 (N_11986,N_11769,N_11781);
nand U11987 (N_11987,N_11764,N_11835);
xnor U11988 (N_11988,N_11797,N_11770);
nor U11989 (N_11989,N_11828,N_11753);
nor U11990 (N_11990,N_11797,N_11750);
xnor U11991 (N_11991,N_11868,N_11787);
and U11992 (N_11992,N_11768,N_11824);
or U11993 (N_11993,N_11761,N_11777);
and U11994 (N_11994,N_11784,N_11824);
or U11995 (N_11995,N_11761,N_11860);
nand U11996 (N_11996,N_11828,N_11873);
and U11997 (N_11997,N_11777,N_11781);
nor U11998 (N_11998,N_11849,N_11864);
and U11999 (N_11999,N_11760,N_11790);
or U12000 (N_12000,N_11909,N_11888);
xor U12001 (N_12001,N_11962,N_11933);
nand U12002 (N_12002,N_11999,N_11904);
and U12003 (N_12003,N_11928,N_11976);
nand U12004 (N_12004,N_11935,N_11988);
nor U12005 (N_12005,N_11954,N_11993);
nor U12006 (N_12006,N_11914,N_11939);
nor U12007 (N_12007,N_11911,N_11883);
nand U12008 (N_12008,N_11951,N_11921);
nand U12009 (N_12009,N_11961,N_11968);
or U12010 (N_12010,N_11896,N_11912);
or U12011 (N_12011,N_11932,N_11978);
and U12012 (N_12012,N_11929,N_11897);
xor U12013 (N_12013,N_11877,N_11958);
or U12014 (N_12014,N_11894,N_11992);
xor U12015 (N_12015,N_11947,N_11881);
nor U12016 (N_12016,N_11891,N_11908);
or U12017 (N_12017,N_11991,N_11945);
or U12018 (N_12018,N_11882,N_11998);
nor U12019 (N_12019,N_11952,N_11918);
and U12020 (N_12020,N_11920,N_11900);
nand U12021 (N_12021,N_11878,N_11949);
nand U12022 (N_12022,N_11892,N_11938);
or U12023 (N_12023,N_11995,N_11983);
xnor U12024 (N_12024,N_11927,N_11989);
nor U12025 (N_12025,N_11971,N_11946);
or U12026 (N_12026,N_11981,N_11955);
or U12027 (N_12027,N_11922,N_11887);
or U12028 (N_12028,N_11899,N_11996);
or U12029 (N_12029,N_11943,N_11957);
and U12030 (N_12030,N_11948,N_11987);
and U12031 (N_12031,N_11984,N_11919);
or U12032 (N_12032,N_11880,N_11953);
nand U12033 (N_12033,N_11926,N_11916);
nor U12034 (N_12034,N_11964,N_11893);
xor U12035 (N_12035,N_11885,N_11905);
and U12036 (N_12036,N_11972,N_11985);
nand U12037 (N_12037,N_11963,N_11941);
nor U12038 (N_12038,N_11977,N_11910);
and U12039 (N_12039,N_11944,N_11931);
nor U12040 (N_12040,N_11913,N_11902);
nor U12041 (N_12041,N_11979,N_11901);
and U12042 (N_12042,N_11986,N_11940);
xnor U12043 (N_12043,N_11959,N_11970);
or U12044 (N_12044,N_11967,N_11982);
and U12045 (N_12045,N_11934,N_11965);
or U12046 (N_12046,N_11889,N_11936);
nor U12047 (N_12047,N_11975,N_11942);
and U12048 (N_12048,N_11875,N_11960);
or U12049 (N_12049,N_11923,N_11930);
nor U12050 (N_12050,N_11903,N_11994);
xnor U12051 (N_12051,N_11980,N_11884);
or U12052 (N_12052,N_11966,N_11990);
and U12053 (N_12053,N_11969,N_11917);
and U12054 (N_12054,N_11915,N_11950);
nand U12055 (N_12055,N_11895,N_11886);
or U12056 (N_12056,N_11898,N_11876);
and U12057 (N_12057,N_11879,N_11997);
nor U12058 (N_12058,N_11890,N_11925);
nand U12059 (N_12059,N_11973,N_11937);
or U12060 (N_12060,N_11956,N_11907);
and U12061 (N_12061,N_11906,N_11924);
and U12062 (N_12062,N_11974,N_11907);
xor U12063 (N_12063,N_11901,N_11893);
xor U12064 (N_12064,N_11880,N_11998);
and U12065 (N_12065,N_11955,N_11906);
nor U12066 (N_12066,N_11895,N_11937);
nand U12067 (N_12067,N_11959,N_11885);
or U12068 (N_12068,N_11886,N_11880);
and U12069 (N_12069,N_11921,N_11991);
or U12070 (N_12070,N_11901,N_11930);
or U12071 (N_12071,N_11972,N_11882);
nor U12072 (N_12072,N_11960,N_11929);
nor U12073 (N_12073,N_11977,N_11958);
xor U12074 (N_12074,N_11892,N_11884);
xnor U12075 (N_12075,N_11979,N_11919);
or U12076 (N_12076,N_11926,N_11929);
and U12077 (N_12077,N_11973,N_11915);
nand U12078 (N_12078,N_11895,N_11955);
xor U12079 (N_12079,N_11928,N_11960);
nand U12080 (N_12080,N_11970,N_11909);
nand U12081 (N_12081,N_11915,N_11977);
and U12082 (N_12082,N_11984,N_11913);
or U12083 (N_12083,N_11883,N_11875);
nand U12084 (N_12084,N_11921,N_11962);
xnor U12085 (N_12085,N_11878,N_11900);
nor U12086 (N_12086,N_11895,N_11952);
and U12087 (N_12087,N_11973,N_11994);
or U12088 (N_12088,N_11911,N_11961);
or U12089 (N_12089,N_11979,N_11923);
nor U12090 (N_12090,N_11990,N_11880);
nor U12091 (N_12091,N_11988,N_11899);
and U12092 (N_12092,N_11898,N_11875);
xnor U12093 (N_12093,N_11926,N_11895);
nor U12094 (N_12094,N_11941,N_11905);
nand U12095 (N_12095,N_11910,N_11995);
and U12096 (N_12096,N_11957,N_11931);
xor U12097 (N_12097,N_11998,N_11875);
nor U12098 (N_12098,N_11901,N_11880);
nor U12099 (N_12099,N_11999,N_11978);
or U12100 (N_12100,N_11888,N_11892);
and U12101 (N_12101,N_11956,N_11915);
or U12102 (N_12102,N_11921,N_11889);
nand U12103 (N_12103,N_11989,N_11951);
and U12104 (N_12104,N_11903,N_11904);
xor U12105 (N_12105,N_11875,N_11953);
nor U12106 (N_12106,N_11931,N_11932);
xnor U12107 (N_12107,N_11889,N_11995);
or U12108 (N_12108,N_11919,N_11938);
and U12109 (N_12109,N_11906,N_11901);
nor U12110 (N_12110,N_11903,N_11891);
or U12111 (N_12111,N_11889,N_11930);
or U12112 (N_12112,N_11974,N_11908);
xor U12113 (N_12113,N_11970,N_11989);
nor U12114 (N_12114,N_11892,N_11966);
and U12115 (N_12115,N_11925,N_11907);
or U12116 (N_12116,N_11907,N_11918);
nor U12117 (N_12117,N_11904,N_11915);
or U12118 (N_12118,N_11930,N_11997);
or U12119 (N_12119,N_11964,N_11890);
and U12120 (N_12120,N_11961,N_11980);
nand U12121 (N_12121,N_11990,N_11879);
and U12122 (N_12122,N_11945,N_11885);
nand U12123 (N_12123,N_11923,N_11924);
xnor U12124 (N_12124,N_11919,N_11944);
nand U12125 (N_12125,N_12002,N_12006);
or U12126 (N_12126,N_12056,N_12045);
and U12127 (N_12127,N_12023,N_12099);
and U12128 (N_12128,N_12104,N_12120);
nor U12129 (N_12129,N_12097,N_12122);
or U12130 (N_12130,N_12007,N_12054);
xor U12131 (N_12131,N_12014,N_12030);
nand U12132 (N_12132,N_12085,N_12049);
or U12133 (N_12133,N_12088,N_12087);
nand U12134 (N_12134,N_12025,N_12073);
or U12135 (N_12135,N_12036,N_12121);
nor U12136 (N_12136,N_12101,N_12020);
or U12137 (N_12137,N_12011,N_12110);
or U12138 (N_12138,N_12062,N_12096);
nor U12139 (N_12139,N_12076,N_12052);
nand U12140 (N_12140,N_12041,N_12053);
xor U12141 (N_12141,N_12103,N_12080);
or U12142 (N_12142,N_12005,N_12024);
and U12143 (N_12143,N_12015,N_12113);
nand U12144 (N_12144,N_12107,N_12070);
nor U12145 (N_12145,N_12013,N_12100);
and U12146 (N_12146,N_12065,N_12086);
xor U12147 (N_12147,N_12075,N_12078);
and U12148 (N_12148,N_12040,N_12072);
xor U12149 (N_12149,N_12067,N_12057);
and U12150 (N_12150,N_12061,N_12089);
and U12151 (N_12151,N_12047,N_12026);
or U12152 (N_12152,N_12032,N_12090);
or U12153 (N_12153,N_12034,N_12031);
xor U12154 (N_12154,N_12050,N_12000);
nor U12155 (N_12155,N_12009,N_12051);
nand U12156 (N_12156,N_12058,N_12111);
or U12157 (N_12157,N_12106,N_12092);
xnor U12158 (N_12158,N_12029,N_12119);
nand U12159 (N_12159,N_12066,N_12083);
nand U12160 (N_12160,N_12069,N_12004);
xnor U12161 (N_12161,N_12064,N_12102);
or U12162 (N_12162,N_12012,N_12035);
and U12163 (N_12163,N_12019,N_12117);
or U12164 (N_12164,N_12094,N_12098);
nor U12165 (N_12165,N_12071,N_12044);
or U12166 (N_12166,N_12068,N_12115);
and U12167 (N_12167,N_12039,N_12124);
xor U12168 (N_12168,N_12081,N_12043);
and U12169 (N_12169,N_12008,N_12060);
xor U12170 (N_12170,N_12027,N_12116);
and U12171 (N_12171,N_12028,N_12118);
nor U12172 (N_12172,N_12037,N_12112);
nor U12173 (N_12173,N_12109,N_12114);
or U12174 (N_12174,N_12063,N_12021);
nor U12175 (N_12175,N_12079,N_12091);
xnor U12176 (N_12176,N_12123,N_12093);
nand U12177 (N_12177,N_12082,N_12003);
nand U12178 (N_12178,N_12001,N_12059);
nor U12179 (N_12179,N_12018,N_12022);
xnor U12180 (N_12180,N_12074,N_12055);
and U12181 (N_12181,N_12095,N_12010);
nand U12182 (N_12182,N_12048,N_12077);
xor U12183 (N_12183,N_12038,N_12033);
nor U12184 (N_12184,N_12016,N_12046);
nor U12185 (N_12185,N_12108,N_12042);
nand U12186 (N_12186,N_12017,N_12084);
or U12187 (N_12187,N_12105,N_12011);
nor U12188 (N_12188,N_12004,N_12058);
xnor U12189 (N_12189,N_12103,N_12061);
and U12190 (N_12190,N_12113,N_12049);
or U12191 (N_12191,N_12113,N_12070);
or U12192 (N_12192,N_12038,N_12083);
nor U12193 (N_12193,N_12080,N_12108);
or U12194 (N_12194,N_12007,N_12057);
and U12195 (N_12195,N_12110,N_12001);
nand U12196 (N_12196,N_12069,N_12029);
or U12197 (N_12197,N_12112,N_12046);
xnor U12198 (N_12198,N_12094,N_12076);
and U12199 (N_12199,N_12119,N_12074);
nor U12200 (N_12200,N_12071,N_12094);
nand U12201 (N_12201,N_12042,N_12036);
nand U12202 (N_12202,N_12063,N_12016);
xor U12203 (N_12203,N_12043,N_12006);
xnor U12204 (N_12204,N_12066,N_12121);
and U12205 (N_12205,N_12101,N_12008);
or U12206 (N_12206,N_12124,N_12056);
and U12207 (N_12207,N_12034,N_12041);
xor U12208 (N_12208,N_12109,N_12108);
and U12209 (N_12209,N_12066,N_12123);
or U12210 (N_12210,N_12118,N_12006);
and U12211 (N_12211,N_12025,N_12049);
nor U12212 (N_12212,N_12107,N_12043);
or U12213 (N_12213,N_12024,N_12088);
xor U12214 (N_12214,N_12001,N_12032);
xor U12215 (N_12215,N_12053,N_12003);
and U12216 (N_12216,N_12098,N_12067);
nand U12217 (N_12217,N_12030,N_12040);
xnor U12218 (N_12218,N_12080,N_12098);
nor U12219 (N_12219,N_12021,N_12030);
or U12220 (N_12220,N_12110,N_12017);
xnor U12221 (N_12221,N_12031,N_12121);
nor U12222 (N_12222,N_12123,N_12091);
nor U12223 (N_12223,N_12013,N_12044);
and U12224 (N_12224,N_12094,N_12084);
or U12225 (N_12225,N_12114,N_12108);
xnor U12226 (N_12226,N_12011,N_12032);
xnor U12227 (N_12227,N_12045,N_12032);
and U12228 (N_12228,N_12118,N_12032);
and U12229 (N_12229,N_12045,N_12122);
and U12230 (N_12230,N_12027,N_12010);
or U12231 (N_12231,N_12071,N_12019);
or U12232 (N_12232,N_12106,N_12060);
nor U12233 (N_12233,N_12071,N_12028);
xor U12234 (N_12234,N_12041,N_12090);
nand U12235 (N_12235,N_12058,N_12019);
nor U12236 (N_12236,N_12008,N_12098);
xnor U12237 (N_12237,N_12111,N_12035);
and U12238 (N_12238,N_12013,N_12113);
nor U12239 (N_12239,N_12009,N_12058);
nor U12240 (N_12240,N_12012,N_12091);
nor U12241 (N_12241,N_12063,N_12014);
nand U12242 (N_12242,N_12124,N_12099);
nor U12243 (N_12243,N_12110,N_12085);
and U12244 (N_12244,N_12095,N_12054);
or U12245 (N_12245,N_12116,N_12023);
nor U12246 (N_12246,N_12037,N_12001);
or U12247 (N_12247,N_12066,N_12019);
and U12248 (N_12248,N_12059,N_12007);
xor U12249 (N_12249,N_12052,N_12035);
and U12250 (N_12250,N_12204,N_12135);
or U12251 (N_12251,N_12184,N_12174);
xnor U12252 (N_12252,N_12216,N_12159);
nor U12253 (N_12253,N_12169,N_12232);
nor U12254 (N_12254,N_12185,N_12214);
nor U12255 (N_12255,N_12209,N_12243);
xor U12256 (N_12256,N_12161,N_12242);
and U12257 (N_12257,N_12234,N_12141);
nand U12258 (N_12258,N_12136,N_12188);
nor U12259 (N_12259,N_12177,N_12194);
nand U12260 (N_12260,N_12142,N_12158);
xnor U12261 (N_12261,N_12150,N_12165);
nand U12262 (N_12262,N_12182,N_12171);
nor U12263 (N_12263,N_12130,N_12144);
nand U12264 (N_12264,N_12132,N_12152);
nand U12265 (N_12265,N_12133,N_12183);
and U12266 (N_12266,N_12192,N_12248);
and U12267 (N_12267,N_12128,N_12186);
or U12268 (N_12268,N_12200,N_12149);
and U12269 (N_12269,N_12160,N_12138);
nand U12270 (N_12270,N_12131,N_12202);
xnor U12271 (N_12271,N_12235,N_12168);
nor U12272 (N_12272,N_12226,N_12230);
nand U12273 (N_12273,N_12198,N_12220);
xor U12274 (N_12274,N_12127,N_12175);
nor U12275 (N_12275,N_12180,N_12176);
and U12276 (N_12276,N_12239,N_12241);
nand U12277 (N_12277,N_12181,N_12140);
or U12278 (N_12278,N_12195,N_12231);
nand U12279 (N_12279,N_12219,N_12148);
nor U12280 (N_12280,N_12143,N_12237);
nand U12281 (N_12281,N_12153,N_12172);
nor U12282 (N_12282,N_12203,N_12146);
nor U12283 (N_12283,N_12217,N_12166);
and U12284 (N_12284,N_12126,N_12238);
nor U12285 (N_12285,N_12240,N_12212);
or U12286 (N_12286,N_12137,N_12173);
nand U12287 (N_12287,N_12207,N_12208);
nand U12288 (N_12288,N_12139,N_12245);
nand U12289 (N_12289,N_12134,N_12129);
nor U12290 (N_12290,N_12223,N_12179);
or U12291 (N_12291,N_12224,N_12199);
xor U12292 (N_12292,N_12170,N_12162);
nand U12293 (N_12293,N_12246,N_12178);
xor U12294 (N_12294,N_12156,N_12225);
xnor U12295 (N_12295,N_12218,N_12157);
nor U12296 (N_12296,N_12215,N_12227);
xor U12297 (N_12297,N_12164,N_12190);
nand U12298 (N_12298,N_12210,N_12145);
xnor U12299 (N_12299,N_12187,N_12197);
xor U12300 (N_12300,N_12247,N_12233);
nand U12301 (N_12301,N_12213,N_12249);
nand U12302 (N_12302,N_12193,N_12167);
nand U12303 (N_12303,N_12191,N_12201);
and U12304 (N_12304,N_12229,N_12221);
nand U12305 (N_12305,N_12244,N_12125);
nand U12306 (N_12306,N_12189,N_12228);
or U12307 (N_12307,N_12154,N_12205);
or U12308 (N_12308,N_12211,N_12155);
and U12309 (N_12309,N_12151,N_12206);
and U12310 (N_12310,N_12196,N_12163);
or U12311 (N_12311,N_12236,N_12222);
and U12312 (N_12312,N_12147,N_12132);
nand U12313 (N_12313,N_12249,N_12207);
xnor U12314 (N_12314,N_12206,N_12240);
xor U12315 (N_12315,N_12204,N_12162);
and U12316 (N_12316,N_12231,N_12204);
nor U12317 (N_12317,N_12213,N_12234);
nand U12318 (N_12318,N_12225,N_12136);
nor U12319 (N_12319,N_12147,N_12234);
or U12320 (N_12320,N_12211,N_12210);
nand U12321 (N_12321,N_12160,N_12245);
and U12322 (N_12322,N_12153,N_12235);
nand U12323 (N_12323,N_12125,N_12150);
nand U12324 (N_12324,N_12213,N_12136);
nand U12325 (N_12325,N_12150,N_12239);
nor U12326 (N_12326,N_12171,N_12245);
nand U12327 (N_12327,N_12172,N_12177);
nor U12328 (N_12328,N_12205,N_12136);
nand U12329 (N_12329,N_12161,N_12126);
and U12330 (N_12330,N_12191,N_12167);
nand U12331 (N_12331,N_12200,N_12167);
nor U12332 (N_12332,N_12133,N_12151);
nand U12333 (N_12333,N_12157,N_12190);
and U12334 (N_12334,N_12192,N_12171);
nand U12335 (N_12335,N_12220,N_12148);
and U12336 (N_12336,N_12247,N_12219);
xor U12337 (N_12337,N_12236,N_12144);
nor U12338 (N_12338,N_12146,N_12148);
and U12339 (N_12339,N_12128,N_12208);
and U12340 (N_12340,N_12240,N_12127);
nor U12341 (N_12341,N_12235,N_12203);
xor U12342 (N_12342,N_12197,N_12231);
or U12343 (N_12343,N_12221,N_12178);
nor U12344 (N_12344,N_12128,N_12198);
nand U12345 (N_12345,N_12133,N_12221);
xnor U12346 (N_12346,N_12202,N_12214);
and U12347 (N_12347,N_12224,N_12156);
or U12348 (N_12348,N_12163,N_12174);
nor U12349 (N_12349,N_12183,N_12144);
or U12350 (N_12350,N_12155,N_12157);
and U12351 (N_12351,N_12154,N_12198);
xnor U12352 (N_12352,N_12188,N_12154);
xnor U12353 (N_12353,N_12189,N_12147);
nand U12354 (N_12354,N_12137,N_12126);
nor U12355 (N_12355,N_12193,N_12166);
xnor U12356 (N_12356,N_12219,N_12206);
or U12357 (N_12357,N_12188,N_12221);
nand U12358 (N_12358,N_12220,N_12229);
nand U12359 (N_12359,N_12162,N_12209);
nand U12360 (N_12360,N_12247,N_12199);
nor U12361 (N_12361,N_12219,N_12203);
nand U12362 (N_12362,N_12221,N_12129);
xor U12363 (N_12363,N_12223,N_12237);
or U12364 (N_12364,N_12243,N_12229);
and U12365 (N_12365,N_12125,N_12191);
nor U12366 (N_12366,N_12152,N_12166);
nand U12367 (N_12367,N_12141,N_12208);
nand U12368 (N_12368,N_12248,N_12198);
or U12369 (N_12369,N_12193,N_12151);
and U12370 (N_12370,N_12145,N_12163);
nand U12371 (N_12371,N_12244,N_12142);
xor U12372 (N_12372,N_12147,N_12140);
and U12373 (N_12373,N_12153,N_12165);
nor U12374 (N_12374,N_12209,N_12135);
nor U12375 (N_12375,N_12260,N_12293);
xor U12376 (N_12376,N_12309,N_12334);
xor U12377 (N_12377,N_12325,N_12305);
nor U12378 (N_12378,N_12291,N_12333);
and U12379 (N_12379,N_12290,N_12351);
or U12380 (N_12380,N_12259,N_12313);
or U12381 (N_12381,N_12274,N_12354);
and U12382 (N_12382,N_12303,N_12292);
nand U12383 (N_12383,N_12367,N_12271);
xnor U12384 (N_12384,N_12364,N_12299);
nand U12385 (N_12385,N_12308,N_12263);
xnor U12386 (N_12386,N_12282,N_12342);
nor U12387 (N_12387,N_12353,N_12345);
nor U12388 (N_12388,N_12337,N_12300);
nand U12389 (N_12389,N_12258,N_12338);
nand U12390 (N_12390,N_12301,N_12286);
xor U12391 (N_12391,N_12350,N_12283);
nor U12392 (N_12392,N_12356,N_12358);
and U12393 (N_12393,N_12341,N_12253);
or U12394 (N_12394,N_12317,N_12369);
nand U12395 (N_12395,N_12298,N_12347);
xor U12396 (N_12396,N_12294,N_12297);
nor U12397 (N_12397,N_12262,N_12315);
and U12398 (N_12398,N_12321,N_12251);
and U12399 (N_12399,N_12273,N_12267);
xor U12400 (N_12400,N_12370,N_12343);
or U12401 (N_12401,N_12327,N_12296);
and U12402 (N_12402,N_12302,N_12371);
xnor U12403 (N_12403,N_12363,N_12348);
nor U12404 (N_12404,N_12307,N_12320);
xnor U12405 (N_12405,N_12322,N_12314);
and U12406 (N_12406,N_12326,N_12355);
or U12407 (N_12407,N_12323,N_12295);
nor U12408 (N_12408,N_12346,N_12266);
nand U12409 (N_12409,N_12340,N_12310);
nand U12410 (N_12410,N_12319,N_12287);
nand U12411 (N_12411,N_12250,N_12276);
or U12412 (N_12412,N_12336,N_12280);
or U12413 (N_12413,N_12285,N_12349);
or U12414 (N_12414,N_12257,N_12264);
nor U12415 (N_12415,N_12255,N_12284);
nor U12416 (N_12416,N_12366,N_12311);
nor U12417 (N_12417,N_12331,N_12359);
nor U12418 (N_12418,N_12365,N_12281);
nand U12419 (N_12419,N_12328,N_12277);
nor U12420 (N_12420,N_12357,N_12335);
or U12421 (N_12421,N_12352,N_12278);
nor U12422 (N_12422,N_12344,N_12360);
nand U12423 (N_12423,N_12269,N_12275);
or U12424 (N_12424,N_12268,N_12304);
and U12425 (N_12425,N_12372,N_12252);
and U12426 (N_12426,N_12318,N_12368);
nor U12427 (N_12427,N_12373,N_12279);
xor U12428 (N_12428,N_12339,N_12361);
or U12429 (N_12429,N_12329,N_12374);
nor U12430 (N_12430,N_12324,N_12332);
nand U12431 (N_12431,N_12330,N_12270);
and U12432 (N_12432,N_12316,N_12288);
nand U12433 (N_12433,N_12312,N_12272);
nand U12434 (N_12434,N_12289,N_12362);
nand U12435 (N_12435,N_12261,N_12254);
and U12436 (N_12436,N_12256,N_12265);
xnor U12437 (N_12437,N_12306,N_12291);
nor U12438 (N_12438,N_12338,N_12372);
or U12439 (N_12439,N_12316,N_12356);
or U12440 (N_12440,N_12281,N_12269);
and U12441 (N_12441,N_12358,N_12366);
nor U12442 (N_12442,N_12290,N_12314);
nor U12443 (N_12443,N_12369,N_12292);
xor U12444 (N_12444,N_12277,N_12309);
nor U12445 (N_12445,N_12309,N_12282);
nor U12446 (N_12446,N_12330,N_12255);
nand U12447 (N_12447,N_12279,N_12260);
and U12448 (N_12448,N_12299,N_12312);
nand U12449 (N_12449,N_12343,N_12371);
nor U12450 (N_12450,N_12288,N_12299);
and U12451 (N_12451,N_12261,N_12317);
nor U12452 (N_12452,N_12270,N_12360);
and U12453 (N_12453,N_12340,N_12316);
or U12454 (N_12454,N_12266,N_12352);
and U12455 (N_12455,N_12374,N_12318);
and U12456 (N_12456,N_12356,N_12353);
xnor U12457 (N_12457,N_12330,N_12252);
nand U12458 (N_12458,N_12279,N_12334);
xor U12459 (N_12459,N_12291,N_12288);
or U12460 (N_12460,N_12257,N_12301);
and U12461 (N_12461,N_12349,N_12337);
nor U12462 (N_12462,N_12319,N_12336);
xor U12463 (N_12463,N_12289,N_12298);
nand U12464 (N_12464,N_12335,N_12345);
nand U12465 (N_12465,N_12340,N_12270);
and U12466 (N_12466,N_12254,N_12301);
nor U12467 (N_12467,N_12283,N_12307);
or U12468 (N_12468,N_12278,N_12286);
or U12469 (N_12469,N_12339,N_12260);
nor U12470 (N_12470,N_12262,N_12293);
nand U12471 (N_12471,N_12279,N_12372);
nor U12472 (N_12472,N_12272,N_12325);
nand U12473 (N_12473,N_12283,N_12358);
nand U12474 (N_12474,N_12260,N_12333);
nor U12475 (N_12475,N_12324,N_12310);
or U12476 (N_12476,N_12374,N_12342);
nor U12477 (N_12477,N_12318,N_12285);
or U12478 (N_12478,N_12265,N_12322);
xor U12479 (N_12479,N_12251,N_12333);
xnor U12480 (N_12480,N_12315,N_12346);
and U12481 (N_12481,N_12346,N_12347);
or U12482 (N_12482,N_12354,N_12363);
xnor U12483 (N_12483,N_12318,N_12286);
nor U12484 (N_12484,N_12371,N_12276);
xnor U12485 (N_12485,N_12355,N_12321);
nand U12486 (N_12486,N_12340,N_12304);
nor U12487 (N_12487,N_12369,N_12312);
nand U12488 (N_12488,N_12263,N_12369);
nand U12489 (N_12489,N_12305,N_12330);
or U12490 (N_12490,N_12335,N_12263);
or U12491 (N_12491,N_12356,N_12363);
nor U12492 (N_12492,N_12360,N_12261);
and U12493 (N_12493,N_12274,N_12357);
or U12494 (N_12494,N_12309,N_12349);
and U12495 (N_12495,N_12273,N_12330);
nor U12496 (N_12496,N_12279,N_12359);
and U12497 (N_12497,N_12287,N_12338);
or U12498 (N_12498,N_12301,N_12318);
nor U12499 (N_12499,N_12363,N_12340);
nand U12500 (N_12500,N_12498,N_12492);
and U12501 (N_12501,N_12497,N_12423);
nor U12502 (N_12502,N_12397,N_12484);
nand U12503 (N_12503,N_12449,N_12380);
nor U12504 (N_12504,N_12388,N_12424);
and U12505 (N_12505,N_12473,N_12448);
or U12506 (N_12506,N_12447,N_12462);
nor U12507 (N_12507,N_12436,N_12443);
and U12508 (N_12508,N_12435,N_12469);
nand U12509 (N_12509,N_12421,N_12412);
xnor U12510 (N_12510,N_12394,N_12417);
nor U12511 (N_12511,N_12483,N_12482);
and U12512 (N_12512,N_12476,N_12496);
nor U12513 (N_12513,N_12437,N_12486);
nor U12514 (N_12514,N_12493,N_12403);
or U12515 (N_12515,N_12419,N_12416);
or U12516 (N_12516,N_12392,N_12460);
or U12517 (N_12517,N_12451,N_12471);
nor U12518 (N_12518,N_12405,N_12415);
nor U12519 (N_12519,N_12444,N_12377);
nor U12520 (N_12520,N_12453,N_12465);
or U12521 (N_12521,N_12378,N_12464);
or U12522 (N_12522,N_12446,N_12408);
or U12523 (N_12523,N_12432,N_12426);
xnor U12524 (N_12524,N_12458,N_12379);
or U12525 (N_12525,N_12457,N_12428);
and U12526 (N_12526,N_12450,N_12390);
nand U12527 (N_12527,N_12488,N_12459);
nor U12528 (N_12528,N_12396,N_12406);
xnor U12529 (N_12529,N_12409,N_12441);
and U12530 (N_12530,N_12434,N_12485);
and U12531 (N_12531,N_12439,N_12431);
xor U12532 (N_12532,N_12386,N_12491);
nand U12533 (N_12533,N_12395,N_12499);
nor U12534 (N_12534,N_12399,N_12381);
and U12535 (N_12535,N_12393,N_12385);
or U12536 (N_12536,N_12433,N_12384);
or U12537 (N_12537,N_12454,N_12414);
xnor U12538 (N_12538,N_12425,N_12398);
nand U12539 (N_12539,N_12376,N_12461);
and U12540 (N_12540,N_12404,N_12418);
nand U12541 (N_12541,N_12413,N_12442);
or U12542 (N_12542,N_12375,N_12479);
nand U12543 (N_12543,N_12389,N_12445);
nor U12544 (N_12544,N_12440,N_12452);
nor U12545 (N_12545,N_12470,N_12427);
nor U12546 (N_12546,N_12494,N_12382);
xnor U12547 (N_12547,N_12468,N_12472);
xor U12548 (N_12548,N_12391,N_12387);
nor U12549 (N_12549,N_12466,N_12487);
or U12550 (N_12550,N_12495,N_12420);
xor U12551 (N_12551,N_12400,N_12463);
nor U12552 (N_12552,N_12467,N_12490);
or U12553 (N_12553,N_12430,N_12407);
and U12554 (N_12554,N_12478,N_12477);
xnor U12555 (N_12555,N_12475,N_12422);
nand U12556 (N_12556,N_12480,N_12489);
nand U12557 (N_12557,N_12402,N_12481);
xor U12558 (N_12558,N_12383,N_12429);
or U12559 (N_12559,N_12474,N_12410);
nor U12560 (N_12560,N_12438,N_12455);
nand U12561 (N_12561,N_12456,N_12411);
nor U12562 (N_12562,N_12401,N_12409);
or U12563 (N_12563,N_12440,N_12403);
nor U12564 (N_12564,N_12475,N_12431);
nand U12565 (N_12565,N_12419,N_12445);
nor U12566 (N_12566,N_12476,N_12482);
nor U12567 (N_12567,N_12377,N_12404);
nor U12568 (N_12568,N_12488,N_12409);
and U12569 (N_12569,N_12455,N_12474);
nor U12570 (N_12570,N_12467,N_12411);
nand U12571 (N_12571,N_12440,N_12433);
or U12572 (N_12572,N_12435,N_12480);
nor U12573 (N_12573,N_12436,N_12464);
and U12574 (N_12574,N_12440,N_12488);
nand U12575 (N_12575,N_12455,N_12422);
and U12576 (N_12576,N_12495,N_12411);
nand U12577 (N_12577,N_12496,N_12438);
and U12578 (N_12578,N_12456,N_12397);
or U12579 (N_12579,N_12390,N_12465);
and U12580 (N_12580,N_12431,N_12433);
and U12581 (N_12581,N_12489,N_12424);
nand U12582 (N_12582,N_12458,N_12430);
and U12583 (N_12583,N_12381,N_12497);
xor U12584 (N_12584,N_12439,N_12405);
nand U12585 (N_12585,N_12434,N_12397);
and U12586 (N_12586,N_12417,N_12434);
and U12587 (N_12587,N_12493,N_12487);
xor U12588 (N_12588,N_12452,N_12400);
and U12589 (N_12589,N_12395,N_12455);
or U12590 (N_12590,N_12388,N_12418);
nand U12591 (N_12591,N_12433,N_12400);
nor U12592 (N_12592,N_12495,N_12467);
and U12593 (N_12593,N_12487,N_12441);
and U12594 (N_12594,N_12475,N_12493);
nand U12595 (N_12595,N_12418,N_12469);
nor U12596 (N_12596,N_12411,N_12426);
or U12597 (N_12597,N_12407,N_12434);
xor U12598 (N_12598,N_12406,N_12383);
and U12599 (N_12599,N_12408,N_12411);
nor U12600 (N_12600,N_12390,N_12474);
nor U12601 (N_12601,N_12428,N_12455);
and U12602 (N_12602,N_12380,N_12438);
or U12603 (N_12603,N_12499,N_12484);
nand U12604 (N_12604,N_12496,N_12383);
nand U12605 (N_12605,N_12497,N_12444);
xnor U12606 (N_12606,N_12471,N_12436);
nand U12607 (N_12607,N_12484,N_12441);
nand U12608 (N_12608,N_12417,N_12466);
nor U12609 (N_12609,N_12430,N_12490);
nand U12610 (N_12610,N_12458,N_12492);
and U12611 (N_12611,N_12491,N_12391);
and U12612 (N_12612,N_12478,N_12382);
nor U12613 (N_12613,N_12402,N_12429);
xnor U12614 (N_12614,N_12436,N_12461);
or U12615 (N_12615,N_12494,N_12442);
nand U12616 (N_12616,N_12438,N_12453);
nor U12617 (N_12617,N_12485,N_12424);
nor U12618 (N_12618,N_12471,N_12446);
and U12619 (N_12619,N_12412,N_12400);
nor U12620 (N_12620,N_12484,N_12385);
xnor U12621 (N_12621,N_12475,N_12494);
or U12622 (N_12622,N_12483,N_12417);
or U12623 (N_12623,N_12377,N_12408);
and U12624 (N_12624,N_12407,N_12490);
nor U12625 (N_12625,N_12501,N_12527);
nor U12626 (N_12626,N_12607,N_12596);
and U12627 (N_12627,N_12591,N_12585);
or U12628 (N_12628,N_12595,N_12581);
nor U12629 (N_12629,N_12547,N_12579);
or U12630 (N_12630,N_12523,N_12587);
or U12631 (N_12631,N_12537,N_12571);
xnor U12632 (N_12632,N_12609,N_12602);
xor U12633 (N_12633,N_12541,N_12614);
nor U12634 (N_12634,N_12540,N_12560);
xor U12635 (N_12635,N_12530,N_12573);
and U12636 (N_12636,N_12512,N_12549);
or U12637 (N_12637,N_12603,N_12576);
nor U12638 (N_12638,N_12566,N_12505);
and U12639 (N_12639,N_12506,N_12557);
nand U12640 (N_12640,N_12522,N_12601);
or U12641 (N_12641,N_12551,N_12533);
or U12642 (N_12642,N_12565,N_12508);
and U12643 (N_12643,N_12546,N_12590);
nand U12644 (N_12644,N_12572,N_12562);
and U12645 (N_12645,N_12619,N_12531);
nand U12646 (N_12646,N_12509,N_12611);
nand U12647 (N_12647,N_12582,N_12574);
and U12648 (N_12648,N_12553,N_12520);
nand U12649 (N_12649,N_12616,N_12516);
and U12650 (N_12650,N_12564,N_12623);
or U12651 (N_12651,N_12511,N_12594);
nand U12652 (N_12652,N_12598,N_12612);
and U12653 (N_12653,N_12525,N_12532);
nand U12654 (N_12654,N_12577,N_12575);
nand U12655 (N_12655,N_12500,N_12567);
or U12656 (N_12656,N_12524,N_12615);
and U12657 (N_12657,N_12586,N_12518);
or U12658 (N_12658,N_12561,N_12513);
nor U12659 (N_12659,N_12605,N_12510);
or U12660 (N_12660,N_12502,N_12592);
nor U12661 (N_12661,N_12504,N_12556);
nor U12662 (N_12662,N_12608,N_12618);
nand U12663 (N_12663,N_12593,N_12521);
nand U12664 (N_12664,N_12554,N_12600);
xnor U12665 (N_12665,N_12599,N_12578);
nand U12666 (N_12666,N_12528,N_12559);
nor U12667 (N_12667,N_12545,N_12570);
or U12668 (N_12668,N_12534,N_12622);
or U12669 (N_12669,N_12624,N_12569);
nand U12670 (N_12670,N_12515,N_12588);
and U12671 (N_12671,N_12604,N_12542);
xnor U12672 (N_12672,N_12563,N_12620);
xor U12673 (N_12673,N_12610,N_12568);
or U12674 (N_12674,N_12583,N_12597);
nand U12675 (N_12675,N_12535,N_12543);
nor U12676 (N_12676,N_12538,N_12544);
nand U12677 (N_12677,N_12552,N_12503);
and U12678 (N_12678,N_12539,N_12529);
xnor U12679 (N_12679,N_12558,N_12613);
xnor U12680 (N_12680,N_12550,N_12526);
nand U12681 (N_12681,N_12617,N_12584);
nor U12682 (N_12682,N_12514,N_12589);
nand U12683 (N_12683,N_12621,N_12517);
xor U12684 (N_12684,N_12606,N_12555);
xor U12685 (N_12685,N_12507,N_12580);
nor U12686 (N_12686,N_12548,N_12519);
nand U12687 (N_12687,N_12536,N_12531);
and U12688 (N_12688,N_12565,N_12507);
nor U12689 (N_12689,N_12503,N_12519);
or U12690 (N_12690,N_12550,N_12609);
or U12691 (N_12691,N_12502,N_12595);
xnor U12692 (N_12692,N_12544,N_12569);
and U12693 (N_12693,N_12522,N_12517);
nand U12694 (N_12694,N_12537,N_12525);
nand U12695 (N_12695,N_12533,N_12531);
or U12696 (N_12696,N_12580,N_12589);
or U12697 (N_12697,N_12507,N_12568);
and U12698 (N_12698,N_12588,N_12603);
and U12699 (N_12699,N_12612,N_12528);
nor U12700 (N_12700,N_12545,N_12532);
or U12701 (N_12701,N_12543,N_12592);
nor U12702 (N_12702,N_12540,N_12503);
or U12703 (N_12703,N_12505,N_12567);
and U12704 (N_12704,N_12620,N_12553);
nand U12705 (N_12705,N_12582,N_12581);
xor U12706 (N_12706,N_12526,N_12598);
nor U12707 (N_12707,N_12558,N_12584);
xor U12708 (N_12708,N_12537,N_12603);
xor U12709 (N_12709,N_12519,N_12604);
xor U12710 (N_12710,N_12598,N_12605);
xnor U12711 (N_12711,N_12556,N_12590);
nor U12712 (N_12712,N_12585,N_12519);
or U12713 (N_12713,N_12534,N_12602);
nor U12714 (N_12714,N_12602,N_12595);
and U12715 (N_12715,N_12568,N_12541);
nand U12716 (N_12716,N_12542,N_12500);
xor U12717 (N_12717,N_12616,N_12512);
nand U12718 (N_12718,N_12587,N_12518);
nor U12719 (N_12719,N_12542,N_12509);
and U12720 (N_12720,N_12548,N_12571);
xor U12721 (N_12721,N_12559,N_12562);
xnor U12722 (N_12722,N_12618,N_12535);
nor U12723 (N_12723,N_12619,N_12590);
xnor U12724 (N_12724,N_12615,N_12580);
xnor U12725 (N_12725,N_12535,N_12571);
xor U12726 (N_12726,N_12599,N_12518);
nor U12727 (N_12727,N_12547,N_12534);
xor U12728 (N_12728,N_12561,N_12506);
or U12729 (N_12729,N_12576,N_12556);
and U12730 (N_12730,N_12532,N_12551);
or U12731 (N_12731,N_12624,N_12571);
and U12732 (N_12732,N_12573,N_12586);
or U12733 (N_12733,N_12588,N_12557);
nand U12734 (N_12734,N_12553,N_12570);
or U12735 (N_12735,N_12563,N_12597);
and U12736 (N_12736,N_12541,N_12575);
and U12737 (N_12737,N_12602,N_12517);
xnor U12738 (N_12738,N_12573,N_12504);
or U12739 (N_12739,N_12560,N_12512);
and U12740 (N_12740,N_12584,N_12614);
xor U12741 (N_12741,N_12524,N_12561);
and U12742 (N_12742,N_12581,N_12614);
nor U12743 (N_12743,N_12574,N_12519);
and U12744 (N_12744,N_12546,N_12536);
xnor U12745 (N_12745,N_12599,N_12529);
and U12746 (N_12746,N_12623,N_12560);
nor U12747 (N_12747,N_12558,N_12545);
nor U12748 (N_12748,N_12556,N_12591);
nand U12749 (N_12749,N_12528,N_12553);
and U12750 (N_12750,N_12644,N_12696);
xnor U12751 (N_12751,N_12749,N_12735);
nand U12752 (N_12752,N_12640,N_12663);
xnor U12753 (N_12753,N_12686,N_12737);
xor U12754 (N_12754,N_12685,N_12648);
xor U12755 (N_12755,N_12664,N_12680);
and U12756 (N_12756,N_12661,N_12647);
nor U12757 (N_12757,N_12746,N_12638);
nor U12758 (N_12758,N_12651,N_12697);
or U12759 (N_12759,N_12710,N_12712);
or U12760 (N_12760,N_12673,N_12694);
and U12761 (N_12761,N_12630,N_12650);
nor U12762 (N_12762,N_12718,N_12695);
or U12763 (N_12763,N_12649,N_12681);
or U12764 (N_12764,N_12625,N_12721);
or U12765 (N_12765,N_12748,N_12662);
nor U12766 (N_12766,N_12688,N_12634);
nand U12767 (N_12767,N_12679,N_12646);
nor U12768 (N_12768,N_12631,N_12671);
nand U12769 (N_12769,N_12667,N_12684);
xor U12770 (N_12770,N_12675,N_12730);
or U12771 (N_12771,N_12692,N_12629);
and U12772 (N_12772,N_12668,N_12690);
or U12773 (N_12773,N_12722,N_12732);
or U12774 (N_12774,N_12659,N_12636);
and U12775 (N_12775,N_12645,N_12708);
and U12776 (N_12776,N_12683,N_12677);
nand U12777 (N_12777,N_12652,N_12698);
xnor U12778 (N_12778,N_12632,N_12719);
or U12779 (N_12779,N_12744,N_12728);
nor U12780 (N_12780,N_12736,N_12742);
and U12781 (N_12781,N_12738,N_12637);
nor U12782 (N_12782,N_12672,N_12653);
or U12783 (N_12783,N_12727,N_12733);
nor U12784 (N_12784,N_12703,N_12639);
xnor U12785 (N_12785,N_12635,N_12725);
or U12786 (N_12786,N_12726,N_12702);
xor U12787 (N_12787,N_12655,N_12704);
nor U12788 (N_12788,N_12691,N_12657);
or U12789 (N_12789,N_12699,N_12747);
xnor U12790 (N_12790,N_12676,N_12670);
nor U12791 (N_12791,N_12740,N_12628);
xor U12792 (N_12792,N_12723,N_12693);
xnor U12793 (N_12793,N_12656,N_12720);
or U12794 (N_12794,N_12739,N_12714);
nor U12795 (N_12795,N_12658,N_12705);
and U12796 (N_12796,N_12716,N_12689);
nor U12797 (N_12797,N_12724,N_12715);
or U12798 (N_12798,N_12678,N_12707);
or U12799 (N_12799,N_12731,N_12701);
or U12800 (N_12800,N_12654,N_12706);
and U12801 (N_12801,N_12641,N_12682);
xor U12802 (N_12802,N_12669,N_12666);
xor U12803 (N_12803,N_12717,N_12627);
nand U12804 (N_12804,N_12665,N_12660);
nand U12805 (N_12805,N_12713,N_12643);
and U12806 (N_12806,N_12626,N_12687);
xor U12807 (N_12807,N_12642,N_12633);
nor U12808 (N_12808,N_12729,N_12674);
nor U12809 (N_12809,N_12734,N_12743);
nand U12810 (N_12810,N_12709,N_12700);
and U12811 (N_12811,N_12741,N_12711);
xor U12812 (N_12812,N_12745,N_12693);
and U12813 (N_12813,N_12673,N_12686);
nor U12814 (N_12814,N_12684,N_12632);
nand U12815 (N_12815,N_12725,N_12677);
or U12816 (N_12816,N_12640,N_12673);
or U12817 (N_12817,N_12635,N_12636);
xor U12818 (N_12818,N_12654,N_12695);
nor U12819 (N_12819,N_12630,N_12668);
xor U12820 (N_12820,N_12656,N_12672);
and U12821 (N_12821,N_12710,N_12631);
or U12822 (N_12822,N_12714,N_12705);
nor U12823 (N_12823,N_12646,N_12703);
xor U12824 (N_12824,N_12647,N_12689);
or U12825 (N_12825,N_12715,N_12711);
nor U12826 (N_12826,N_12626,N_12659);
nor U12827 (N_12827,N_12736,N_12659);
nand U12828 (N_12828,N_12645,N_12635);
nor U12829 (N_12829,N_12635,N_12698);
nand U12830 (N_12830,N_12689,N_12676);
nand U12831 (N_12831,N_12629,N_12741);
and U12832 (N_12832,N_12707,N_12648);
xnor U12833 (N_12833,N_12640,N_12674);
xnor U12834 (N_12834,N_12681,N_12705);
nor U12835 (N_12835,N_12745,N_12675);
and U12836 (N_12836,N_12710,N_12688);
nand U12837 (N_12837,N_12711,N_12625);
and U12838 (N_12838,N_12640,N_12664);
nand U12839 (N_12839,N_12678,N_12701);
nor U12840 (N_12840,N_12640,N_12700);
nor U12841 (N_12841,N_12748,N_12731);
nand U12842 (N_12842,N_12718,N_12700);
nor U12843 (N_12843,N_12718,N_12699);
and U12844 (N_12844,N_12628,N_12729);
nand U12845 (N_12845,N_12717,N_12708);
or U12846 (N_12846,N_12712,N_12629);
xor U12847 (N_12847,N_12661,N_12720);
nand U12848 (N_12848,N_12703,N_12657);
and U12849 (N_12849,N_12699,N_12626);
nand U12850 (N_12850,N_12642,N_12647);
nand U12851 (N_12851,N_12724,N_12735);
or U12852 (N_12852,N_12661,N_12690);
or U12853 (N_12853,N_12626,N_12682);
xnor U12854 (N_12854,N_12721,N_12681);
or U12855 (N_12855,N_12675,N_12722);
xnor U12856 (N_12856,N_12715,N_12694);
and U12857 (N_12857,N_12680,N_12628);
or U12858 (N_12858,N_12717,N_12672);
and U12859 (N_12859,N_12693,N_12677);
and U12860 (N_12860,N_12674,N_12728);
or U12861 (N_12861,N_12641,N_12655);
xor U12862 (N_12862,N_12689,N_12705);
xor U12863 (N_12863,N_12700,N_12719);
or U12864 (N_12864,N_12685,N_12679);
nor U12865 (N_12865,N_12704,N_12707);
nor U12866 (N_12866,N_12667,N_12626);
nand U12867 (N_12867,N_12687,N_12713);
nor U12868 (N_12868,N_12655,N_12666);
and U12869 (N_12869,N_12628,N_12743);
nor U12870 (N_12870,N_12628,N_12661);
nor U12871 (N_12871,N_12649,N_12682);
or U12872 (N_12872,N_12660,N_12643);
nand U12873 (N_12873,N_12651,N_12667);
nand U12874 (N_12874,N_12669,N_12699);
and U12875 (N_12875,N_12760,N_12780);
nand U12876 (N_12876,N_12822,N_12754);
and U12877 (N_12877,N_12830,N_12862);
nor U12878 (N_12878,N_12861,N_12824);
or U12879 (N_12879,N_12870,N_12874);
nand U12880 (N_12880,N_12779,N_12794);
xnor U12881 (N_12881,N_12752,N_12840);
or U12882 (N_12882,N_12781,N_12852);
and U12883 (N_12883,N_12848,N_12823);
nor U12884 (N_12884,N_12806,N_12792);
nand U12885 (N_12885,N_12765,N_12783);
and U12886 (N_12886,N_12801,N_12759);
xnor U12887 (N_12887,N_12827,N_12856);
nand U12888 (N_12888,N_12858,N_12787);
nor U12889 (N_12889,N_12771,N_12857);
xor U12890 (N_12890,N_12797,N_12812);
or U12891 (N_12891,N_12853,N_12756);
or U12892 (N_12892,N_12831,N_12834);
or U12893 (N_12893,N_12762,N_12820);
xor U12894 (N_12894,N_12753,N_12828);
nor U12895 (N_12895,N_12776,N_12800);
nor U12896 (N_12896,N_12810,N_12850);
nand U12897 (N_12897,N_12763,N_12821);
nor U12898 (N_12898,N_12805,N_12757);
nand U12899 (N_12899,N_12844,N_12802);
nor U12900 (N_12900,N_12795,N_12838);
nand U12901 (N_12901,N_12767,N_12761);
nor U12902 (N_12902,N_12864,N_12817);
xor U12903 (N_12903,N_12793,N_12815);
xnor U12904 (N_12904,N_12841,N_12769);
or U12905 (N_12905,N_12829,N_12766);
nor U12906 (N_12906,N_12842,N_12835);
nor U12907 (N_12907,N_12774,N_12784);
nor U12908 (N_12908,N_12871,N_12775);
xor U12909 (N_12909,N_12837,N_12778);
xor U12910 (N_12910,N_12782,N_12814);
nand U12911 (N_12911,N_12789,N_12818);
or U12912 (N_12912,N_12799,N_12855);
or U12913 (N_12913,N_12796,N_12854);
or U12914 (N_12914,N_12859,N_12758);
and U12915 (N_12915,N_12873,N_12839);
xor U12916 (N_12916,N_12770,N_12813);
xnor U12917 (N_12917,N_12809,N_12790);
nand U12918 (N_12918,N_12811,N_12863);
or U12919 (N_12919,N_12836,N_12849);
and U12920 (N_12920,N_12785,N_12833);
nor U12921 (N_12921,N_12777,N_12865);
or U12922 (N_12922,N_12768,N_12826);
and U12923 (N_12923,N_12867,N_12750);
nor U12924 (N_12924,N_12803,N_12791);
nor U12925 (N_12925,N_12860,N_12866);
nand U12926 (N_12926,N_12788,N_12816);
or U12927 (N_12927,N_12832,N_12764);
nand U12928 (N_12928,N_12872,N_12807);
and U12929 (N_12929,N_12846,N_12825);
nand U12930 (N_12930,N_12843,N_12772);
xor U12931 (N_12931,N_12786,N_12808);
or U12932 (N_12932,N_12868,N_12751);
xor U12933 (N_12933,N_12847,N_12851);
xnor U12934 (N_12934,N_12804,N_12845);
and U12935 (N_12935,N_12773,N_12755);
xor U12936 (N_12936,N_12819,N_12798);
and U12937 (N_12937,N_12869,N_12824);
or U12938 (N_12938,N_12812,N_12805);
or U12939 (N_12939,N_12763,N_12751);
or U12940 (N_12940,N_12753,N_12789);
xnor U12941 (N_12941,N_12852,N_12799);
or U12942 (N_12942,N_12827,N_12831);
nand U12943 (N_12943,N_12773,N_12836);
or U12944 (N_12944,N_12779,N_12760);
or U12945 (N_12945,N_12822,N_12872);
xor U12946 (N_12946,N_12823,N_12792);
xnor U12947 (N_12947,N_12808,N_12784);
nor U12948 (N_12948,N_12751,N_12843);
or U12949 (N_12949,N_12794,N_12772);
xor U12950 (N_12950,N_12835,N_12757);
nand U12951 (N_12951,N_12851,N_12750);
nor U12952 (N_12952,N_12865,N_12782);
nor U12953 (N_12953,N_12808,N_12810);
nand U12954 (N_12954,N_12851,N_12816);
nand U12955 (N_12955,N_12835,N_12866);
nand U12956 (N_12956,N_12865,N_12811);
xnor U12957 (N_12957,N_12865,N_12870);
or U12958 (N_12958,N_12761,N_12813);
or U12959 (N_12959,N_12806,N_12872);
or U12960 (N_12960,N_12787,N_12758);
nor U12961 (N_12961,N_12840,N_12792);
nor U12962 (N_12962,N_12794,N_12813);
and U12963 (N_12963,N_12782,N_12858);
or U12964 (N_12964,N_12837,N_12769);
xnor U12965 (N_12965,N_12848,N_12825);
nor U12966 (N_12966,N_12866,N_12837);
nand U12967 (N_12967,N_12830,N_12783);
nor U12968 (N_12968,N_12867,N_12752);
and U12969 (N_12969,N_12859,N_12826);
and U12970 (N_12970,N_12820,N_12833);
and U12971 (N_12971,N_12870,N_12817);
nor U12972 (N_12972,N_12819,N_12822);
or U12973 (N_12973,N_12858,N_12870);
nor U12974 (N_12974,N_12785,N_12865);
nor U12975 (N_12975,N_12816,N_12766);
or U12976 (N_12976,N_12771,N_12770);
nor U12977 (N_12977,N_12834,N_12792);
nand U12978 (N_12978,N_12751,N_12873);
or U12979 (N_12979,N_12863,N_12815);
xnor U12980 (N_12980,N_12836,N_12868);
nor U12981 (N_12981,N_12768,N_12806);
xnor U12982 (N_12982,N_12795,N_12798);
and U12983 (N_12983,N_12778,N_12769);
xor U12984 (N_12984,N_12809,N_12808);
and U12985 (N_12985,N_12862,N_12813);
or U12986 (N_12986,N_12752,N_12754);
nor U12987 (N_12987,N_12779,N_12751);
nand U12988 (N_12988,N_12829,N_12801);
nand U12989 (N_12989,N_12773,N_12765);
and U12990 (N_12990,N_12861,N_12783);
nor U12991 (N_12991,N_12822,N_12786);
nand U12992 (N_12992,N_12807,N_12763);
and U12993 (N_12993,N_12825,N_12780);
and U12994 (N_12994,N_12792,N_12790);
xor U12995 (N_12995,N_12757,N_12867);
nand U12996 (N_12996,N_12754,N_12808);
nor U12997 (N_12997,N_12817,N_12825);
or U12998 (N_12998,N_12874,N_12866);
and U12999 (N_12999,N_12758,N_12856);
nor U13000 (N_13000,N_12967,N_12970);
or U13001 (N_13001,N_12987,N_12916);
nor U13002 (N_13002,N_12921,N_12878);
xor U13003 (N_13003,N_12966,N_12890);
nand U13004 (N_13004,N_12897,N_12904);
xor U13005 (N_13005,N_12953,N_12886);
nand U13006 (N_13006,N_12946,N_12943);
or U13007 (N_13007,N_12876,N_12982);
xnor U13008 (N_13008,N_12894,N_12998);
and U13009 (N_13009,N_12910,N_12920);
xnor U13010 (N_13010,N_12952,N_12900);
xnor U13011 (N_13011,N_12983,N_12934);
nand U13012 (N_13012,N_12999,N_12907);
nand U13013 (N_13013,N_12914,N_12981);
nand U13014 (N_13014,N_12989,N_12902);
nand U13015 (N_13015,N_12942,N_12911);
and U13016 (N_13016,N_12961,N_12891);
and U13017 (N_13017,N_12888,N_12925);
or U13018 (N_13018,N_12947,N_12991);
and U13019 (N_13019,N_12924,N_12978);
xor U13020 (N_13020,N_12937,N_12899);
xnor U13021 (N_13021,N_12918,N_12906);
nand U13022 (N_13022,N_12923,N_12949);
or U13023 (N_13023,N_12927,N_12940);
or U13024 (N_13024,N_12905,N_12931);
and U13025 (N_13025,N_12932,N_12915);
nor U13026 (N_13026,N_12955,N_12964);
nor U13027 (N_13027,N_12901,N_12877);
nand U13028 (N_13028,N_12880,N_12893);
and U13029 (N_13029,N_12945,N_12883);
or U13030 (N_13030,N_12960,N_12971);
xnor U13031 (N_13031,N_12988,N_12917);
nor U13032 (N_13032,N_12980,N_12939);
xor U13033 (N_13033,N_12979,N_12875);
xor U13034 (N_13034,N_12990,N_12889);
and U13035 (N_13035,N_12976,N_12993);
nor U13036 (N_13036,N_12969,N_12957);
and U13037 (N_13037,N_12985,N_12950);
and U13038 (N_13038,N_12965,N_12912);
nand U13039 (N_13039,N_12958,N_12887);
nor U13040 (N_13040,N_12936,N_12928);
nand U13041 (N_13041,N_12974,N_12977);
nand U13042 (N_13042,N_12885,N_12909);
nand U13043 (N_13043,N_12973,N_12929);
nand U13044 (N_13044,N_12992,N_12919);
xnor U13045 (N_13045,N_12908,N_12951);
xnor U13046 (N_13046,N_12933,N_12935);
or U13047 (N_13047,N_12968,N_12895);
and U13048 (N_13048,N_12984,N_12975);
or U13049 (N_13049,N_12995,N_12884);
nand U13050 (N_13050,N_12892,N_12954);
and U13051 (N_13051,N_12896,N_12972);
or U13052 (N_13052,N_12944,N_12882);
nand U13053 (N_13053,N_12938,N_12930);
nand U13054 (N_13054,N_12922,N_12997);
nor U13055 (N_13055,N_12903,N_12948);
nand U13056 (N_13056,N_12963,N_12881);
nand U13057 (N_13057,N_12994,N_12913);
or U13058 (N_13058,N_12962,N_12941);
xnor U13059 (N_13059,N_12879,N_12956);
nand U13060 (N_13060,N_12898,N_12996);
and U13061 (N_13061,N_12926,N_12986);
xnor U13062 (N_13062,N_12959,N_12962);
xnor U13063 (N_13063,N_12975,N_12900);
nand U13064 (N_13064,N_12953,N_12981);
nor U13065 (N_13065,N_12922,N_12893);
and U13066 (N_13066,N_12949,N_12958);
nand U13067 (N_13067,N_12911,N_12895);
nand U13068 (N_13068,N_12887,N_12980);
or U13069 (N_13069,N_12957,N_12931);
nand U13070 (N_13070,N_12977,N_12895);
nor U13071 (N_13071,N_12956,N_12970);
nand U13072 (N_13072,N_12890,N_12993);
and U13073 (N_13073,N_12998,N_12899);
and U13074 (N_13074,N_12972,N_12969);
and U13075 (N_13075,N_12901,N_12986);
nor U13076 (N_13076,N_12886,N_12941);
nand U13077 (N_13077,N_12915,N_12880);
nand U13078 (N_13078,N_12995,N_12916);
nand U13079 (N_13079,N_12980,N_12944);
nand U13080 (N_13080,N_12989,N_12892);
or U13081 (N_13081,N_12945,N_12936);
nor U13082 (N_13082,N_12973,N_12927);
or U13083 (N_13083,N_12980,N_12882);
xor U13084 (N_13084,N_12882,N_12906);
nand U13085 (N_13085,N_12950,N_12984);
and U13086 (N_13086,N_12885,N_12939);
xnor U13087 (N_13087,N_12970,N_12999);
xnor U13088 (N_13088,N_12963,N_12988);
or U13089 (N_13089,N_12947,N_12875);
nand U13090 (N_13090,N_12928,N_12992);
and U13091 (N_13091,N_12932,N_12962);
or U13092 (N_13092,N_12944,N_12945);
nand U13093 (N_13093,N_12985,N_12948);
nor U13094 (N_13094,N_12880,N_12875);
nand U13095 (N_13095,N_12970,N_12952);
nor U13096 (N_13096,N_12925,N_12949);
and U13097 (N_13097,N_12891,N_12982);
or U13098 (N_13098,N_12883,N_12882);
or U13099 (N_13099,N_12887,N_12905);
or U13100 (N_13100,N_12995,N_12909);
nand U13101 (N_13101,N_12899,N_12975);
nand U13102 (N_13102,N_12941,N_12909);
xnor U13103 (N_13103,N_12877,N_12935);
nand U13104 (N_13104,N_12881,N_12936);
or U13105 (N_13105,N_12977,N_12887);
nor U13106 (N_13106,N_12902,N_12999);
and U13107 (N_13107,N_12995,N_12964);
and U13108 (N_13108,N_12905,N_12879);
or U13109 (N_13109,N_12900,N_12979);
xor U13110 (N_13110,N_12896,N_12885);
nand U13111 (N_13111,N_12958,N_12954);
nor U13112 (N_13112,N_12878,N_12929);
xnor U13113 (N_13113,N_12910,N_12949);
xor U13114 (N_13114,N_12910,N_12995);
nor U13115 (N_13115,N_12901,N_12990);
nand U13116 (N_13116,N_12948,N_12889);
nand U13117 (N_13117,N_12896,N_12905);
and U13118 (N_13118,N_12877,N_12934);
nand U13119 (N_13119,N_12984,N_12919);
nand U13120 (N_13120,N_12928,N_12912);
or U13121 (N_13121,N_12989,N_12968);
nor U13122 (N_13122,N_12904,N_12935);
or U13123 (N_13123,N_12924,N_12883);
xor U13124 (N_13124,N_12943,N_12918);
and U13125 (N_13125,N_13042,N_13012);
xor U13126 (N_13126,N_13051,N_13026);
and U13127 (N_13127,N_13107,N_13028);
nand U13128 (N_13128,N_13022,N_13027);
or U13129 (N_13129,N_13071,N_13076);
xnor U13130 (N_13130,N_13038,N_13121);
nand U13131 (N_13131,N_13078,N_13083);
nor U13132 (N_13132,N_13105,N_13090);
nand U13133 (N_13133,N_13109,N_13056);
nor U13134 (N_13134,N_13014,N_13117);
or U13135 (N_13135,N_13072,N_13032);
and U13136 (N_13136,N_13112,N_13104);
nor U13137 (N_13137,N_13123,N_13098);
or U13138 (N_13138,N_13031,N_13011);
and U13139 (N_13139,N_13095,N_13053);
nand U13140 (N_13140,N_13059,N_13120);
nor U13141 (N_13141,N_13005,N_13067);
nand U13142 (N_13142,N_13110,N_13054);
nand U13143 (N_13143,N_13077,N_13087);
xor U13144 (N_13144,N_13004,N_13007);
nor U13145 (N_13145,N_13111,N_13115);
nor U13146 (N_13146,N_13015,N_13050);
or U13147 (N_13147,N_13033,N_13093);
or U13148 (N_13148,N_13037,N_13000);
xnor U13149 (N_13149,N_13069,N_13039);
or U13150 (N_13150,N_13021,N_13114);
or U13151 (N_13151,N_13013,N_13096);
nand U13152 (N_13152,N_13119,N_13019);
or U13153 (N_13153,N_13043,N_13001);
or U13154 (N_13154,N_13081,N_13089);
nor U13155 (N_13155,N_13020,N_13044);
xnor U13156 (N_13156,N_13075,N_13025);
xnor U13157 (N_13157,N_13108,N_13084);
or U13158 (N_13158,N_13003,N_13055);
nand U13159 (N_13159,N_13073,N_13046);
and U13160 (N_13160,N_13023,N_13029);
nor U13161 (N_13161,N_13035,N_13092);
nor U13162 (N_13162,N_13030,N_13079);
and U13163 (N_13163,N_13099,N_13116);
xnor U13164 (N_13164,N_13009,N_13062);
nand U13165 (N_13165,N_13058,N_13048);
nor U13166 (N_13166,N_13118,N_13088);
or U13167 (N_13167,N_13106,N_13024);
xnor U13168 (N_13168,N_13008,N_13097);
nor U13169 (N_13169,N_13018,N_13036);
and U13170 (N_13170,N_13061,N_13066);
xor U13171 (N_13171,N_13086,N_13102);
xor U13172 (N_13172,N_13034,N_13124);
nand U13173 (N_13173,N_13057,N_13082);
or U13174 (N_13174,N_13101,N_13006);
nor U13175 (N_13175,N_13002,N_13065);
and U13176 (N_13176,N_13094,N_13010);
and U13177 (N_13177,N_13045,N_13040);
nor U13178 (N_13178,N_13041,N_13060);
nand U13179 (N_13179,N_13063,N_13122);
or U13180 (N_13180,N_13080,N_13100);
and U13181 (N_13181,N_13074,N_13091);
xor U13182 (N_13182,N_13070,N_13017);
xnor U13183 (N_13183,N_13113,N_13016);
xnor U13184 (N_13184,N_13052,N_13103);
nand U13185 (N_13185,N_13064,N_13068);
xnor U13186 (N_13186,N_13085,N_13047);
nand U13187 (N_13187,N_13049,N_13108);
nor U13188 (N_13188,N_13040,N_13013);
xnor U13189 (N_13189,N_13081,N_13036);
nand U13190 (N_13190,N_13076,N_13031);
xnor U13191 (N_13191,N_13054,N_13009);
nand U13192 (N_13192,N_13043,N_13011);
and U13193 (N_13193,N_13014,N_13118);
xor U13194 (N_13194,N_13010,N_13043);
nand U13195 (N_13195,N_13118,N_13099);
xor U13196 (N_13196,N_13115,N_13062);
nand U13197 (N_13197,N_13101,N_13033);
or U13198 (N_13198,N_13101,N_13018);
nor U13199 (N_13199,N_13048,N_13025);
and U13200 (N_13200,N_13003,N_13019);
xor U13201 (N_13201,N_13024,N_13064);
nand U13202 (N_13202,N_13041,N_13047);
xor U13203 (N_13203,N_13078,N_13053);
and U13204 (N_13204,N_13102,N_13051);
xnor U13205 (N_13205,N_13073,N_13100);
xor U13206 (N_13206,N_13093,N_13066);
nand U13207 (N_13207,N_13099,N_13051);
and U13208 (N_13208,N_13087,N_13089);
and U13209 (N_13209,N_13078,N_13027);
and U13210 (N_13210,N_13124,N_13067);
or U13211 (N_13211,N_13098,N_13086);
xnor U13212 (N_13212,N_13017,N_13116);
nor U13213 (N_13213,N_13008,N_13077);
and U13214 (N_13214,N_13080,N_13014);
nor U13215 (N_13215,N_13030,N_13001);
nand U13216 (N_13216,N_13115,N_13104);
nor U13217 (N_13217,N_13047,N_13057);
nor U13218 (N_13218,N_13116,N_13060);
or U13219 (N_13219,N_13092,N_13083);
nand U13220 (N_13220,N_13017,N_13023);
or U13221 (N_13221,N_13084,N_13114);
nand U13222 (N_13222,N_13007,N_13102);
and U13223 (N_13223,N_13066,N_13087);
nor U13224 (N_13224,N_13113,N_13103);
and U13225 (N_13225,N_13071,N_13010);
and U13226 (N_13226,N_13072,N_13121);
and U13227 (N_13227,N_13091,N_13108);
and U13228 (N_13228,N_13072,N_13081);
nand U13229 (N_13229,N_13031,N_13002);
or U13230 (N_13230,N_13021,N_13054);
nor U13231 (N_13231,N_13029,N_13123);
nor U13232 (N_13232,N_13065,N_13090);
nand U13233 (N_13233,N_13058,N_13111);
nand U13234 (N_13234,N_13044,N_13052);
and U13235 (N_13235,N_13073,N_13051);
nor U13236 (N_13236,N_13095,N_13024);
or U13237 (N_13237,N_13019,N_13016);
or U13238 (N_13238,N_13005,N_13083);
nor U13239 (N_13239,N_13100,N_13007);
nor U13240 (N_13240,N_13115,N_13013);
nor U13241 (N_13241,N_13118,N_13006);
and U13242 (N_13242,N_13046,N_13038);
and U13243 (N_13243,N_13004,N_13070);
or U13244 (N_13244,N_13015,N_13059);
nor U13245 (N_13245,N_13005,N_13089);
nor U13246 (N_13246,N_13076,N_13059);
nor U13247 (N_13247,N_13069,N_13031);
or U13248 (N_13248,N_13118,N_13020);
xnor U13249 (N_13249,N_13113,N_13085);
xnor U13250 (N_13250,N_13164,N_13149);
nor U13251 (N_13251,N_13220,N_13204);
nand U13252 (N_13252,N_13208,N_13225);
xnor U13253 (N_13253,N_13229,N_13163);
and U13254 (N_13254,N_13244,N_13240);
and U13255 (N_13255,N_13178,N_13172);
or U13256 (N_13256,N_13239,N_13223);
nand U13257 (N_13257,N_13155,N_13158);
xnor U13258 (N_13258,N_13199,N_13186);
nand U13259 (N_13259,N_13167,N_13219);
nand U13260 (N_13260,N_13152,N_13227);
xnor U13261 (N_13261,N_13210,N_13195);
nand U13262 (N_13262,N_13194,N_13129);
or U13263 (N_13263,N_13185,N_13198);
or U13264 (N_13264,N_13126,N_13211);
nand U13265 (N_13265,N_13206,N_13197);
nor U13266 (N_13266,N_13212,N_13173);
nor U13267 (N_13267,N_13188,N_13131);
xnor U13268 (N_13268,N_13168,N_13159);
nand U13269 (N_13269,N_13189,N_13241);
xnor U13270 (N_13270,N_13145,N_13169);
and U13271 (N_13271,N_13228,N_13151);
nand U13272 (N_13272,N_13184,N_13127);
nor U13273 (N_13273,N_13214,N_13153);
or U13274 (N_13274,N_13237,N_13200);
or U13275 (N_13275,N_13134,N_13138);
or U13276 (N_13276,N_13130,N_13190);
or U13277 (N_13277,N_13157,N_13148);
nor U13278 (N_13278,N_13135,N_13232);
or U13279 (N_13279,N_13183,N_13176);
xor U13280 (N_13280,N_13162,N_13202);
or U13281 (N_13281,N_13141,N_13221);
nand U13282 (N_13282,N_13142,N_13222);
xnor U13283 (N_13283,N_13125,N_13224);
xnor U13284 (N_13284,N_13215,N_13249);
or U13285 (N_13285,N_13166,N_13205);
or U13286 (N_13286,N_13180,N_13245);
or U13287 (N_13287,N_13132,N_13179);
nand U13288 (N_13288,N_13143,N_13191);
xor U13289 (N_13289,N_13174,N_13217);
and U13290 (N_13290,N_13147,N_13144);
nand U13291 (N_13291,N_13160,N_13170);
nand U13292 (N_13292,N_13230,N_13146);
or U13293 (N_13293,N_13156,N_13196);
xor U13294 (N_13294,N_13218,N_13246);
nand U13295 (N_13295,N_13247,N_13154);
xor U13296 (N_13296,N_13234,N_13238);
nand U13297 (N_13297,N_13233,N_13187);
and U13298 (N_13298,N_13140,N_13128);
nor U13299 (N_13299,N_13165,N_13231);
nor U13300 (N_13300,N_13193,N_13182);
nand U13301 (N_13301,N_13248,N_13236);
and U13302 (N_13302,N_13207,N_13201);
nand U13303 (N_13303,N_13203,N_13150);
or U13304 (N_13304,N_13139,N_13213);
nor U13305 (N_13305,N_13209,N_13133);
xnor U13306 (N_13306,N_13243,N_13216);
or U13307 (N_13307,N_13161,N_13242);
nor U13308 (N_13308,N_13192,N_13137);
xnor U13309 (N_13309,N_13171,N_13235);
nand U13310 (N_13310,N_13226,N_13181);
and U13311 (N_13311,N_13177,N_13175);
or U13312 (N_13312,N_13136,N_13191);
nand U13313 (N_13313,N_13231,N_13175);
and U13314 (N_13314,N_13205,N_13183);
nand U13315 (N_13315,N_13217,N_13153);
xnor U13316 (N_13316,N_13195,N_13149);
nor U13317 (N_13317,N_13203,N_13245);
and U13318 (N_13318,N_13145,N_13130);
nand U13319 (N_13319,N_13145,N_13227);
nor U13320 (N_13320,N_13172,N_13151);
nand U13321 (N_13321,N_13202,N_13198);
or U13322 (N_13322,N_13186,N_13128);
and U13323 (N_13323,N_13238,N_13146);
xnor U13324 (N_13324,N_13216,N_13234);
and U13325 (N_13325,N_13162,N_13237);
xor U13326 (N_13326,N_13221,N_13222);
xnor U13327 (N_13327,N_13191,N_13141);
and U13328 (N_13328,N_13210,N_13161);
nand U13329 (N_13329,N_13157,N_13217);
nor U13330 (N_13330,N_13246,N_13170);
and U13331 (N_13331,N_13147,N_13180);
xnor U13332 (N_13332,N_13226,N_13159);
xnor U13333 (N_13333,N_13147,N_13237);
or U13334 (N_13334,N_13157,N_13215);
or U13335 (N_13335,N_13232,N_13156);
and U13336 (N_13336,N_13249,N_13176);
and U13337 (N_13337,N_13238,N_13213);
or U13338 (N_13338,N_13187,N_13152);
and U13339 (N_13339,N_13135,N_13193);
xnor U13340 (N_13340,N_13139,N_13155);
xor U13341 (N_13341,N_13157,N_13128);
or U13342 (N_13342,N_13140,N_13174);
and U13343 (N_13343,N_13163,N_13145);
or U13344 (N_13344,N_13189,N_13183);
and U13345 (N_13345,N_13239,N_13178);
xnor U13346 (N_13346,N_13172,N_13180);
nor U13347 (N_13347,N_13239,N_13213);
nand U13348 (N_13348,N_13134,N_13132);
and U13349 (N_13349,N_13227,N_13197);
xnor U13350 (N_13350,N_13212,N_13151);
nor U13351 (N_13351,N_13218,N_13223);
nand U13352 (N_13352,N_13177,N_13242);
and U13353 (N_13353,N_13243,N_13245);
nor U13354 (N_13354,N_13173,N_13230);
or U13355 (N_13355,N_13228,N_13173);
nor U13356 (N_13356,N_13176,N_13181);
or U13357 (N_13357,N_13206,N_13200);
nand U13358 (N_13358,N_13126,N_13215);
nor U13359 (N_13359,N_13169,N_13125);
nand U13360 (N_13360,N_13182,N_13184);
xnor U13361 (N_13361,N_13199,N_13215);
nor U13362 (N_13362,N_13169,N_13196);
nor U13363 (N_13363,N_13137,N_13225);
or U13364 (N_13364,N_13231,N_13163);
and U13365 (N_13365,N_13168,N_13218);
or U13366 (N_13366,N_13221,N_13208);
or U13367 (N_13367,N_13204,N_13168);
and U13368 (N_13368,N_13226,N_13201);
and U13369 (N_13369,N_13140,N_13222);
xor U13370 (N_13370,N_13128,N_13223);
xnor U13371 (N_13371,N_13143,N_13199);
nand U13372 (N_13372,N_13231,N_13162);
xnor U13373 (N_13373,N_13141,N_13219);
or U13374 (N_13374,N_13203,N_13207);
nand U13375 (N_13375,N_13337,N_13288);
or U13376 (N_13376,N_13315,N_13335);
xor U13377 (N_13377,N_13306,N_13291);
xnor U13378 (N_13378,N_13271,N_13327);
nand U13379 (N_13379,N_13343,N_13256);
nor U13380 (N_13380,N_13319,N_13345);
and U13381 (N_13381,N_13290,N_13325);
and U13382 (N_13382,N_13294,N_13340);
or U13383 (N_13383,N_13264,N_13365);
nand U13384 (N_13384,N_13313,N_13359);
nand U13385 (N_13385,N_13351,N_13322);
nor U13386 (N_13386,N_13366,N_13277);
nand U13387 (N_13387,N_13250,N_13317);
and U13388 (N_13388,N_13292,N_13316);
or U13389 (N_13389,N_13265,N_13275);
and U13390 (N_13390,N_13303,N_13344);
or U13391 (N_13391,N_13301,N_13364);
and U13392 (N_13392,N_13312,N_13353);
and U13393 (N_13393,N_13311,N_13360);
and U13394 (N_13394,N_13320,N_13296);
and U13395 (N_13395,N_13302,N_13286);
xor U13396 (N_13396,N_13355,N_13289);
xor U13397 (N_13397,N_13347,N_13338);
nor U13398 (N_13398,N_13333,N_13371);
nor U13399 (N_13399,N_13300,N_13280);
xnor U13400 (N_13400,N_13263,N_13299);
xor U13401 (N_13401,N_13314,N_13334);
nand U13402 (N_13402,N_13267,N_13252);
and U13403 (N_13403,N_13339,N_13284);
nor U13404 (N_13404,N_13323,N_13251);
and U13405 (N_13405,N_13281,N_13309);
and U13406 (N_13406,N_13282,N_13370);
nor U13407 (N_13407,N_13356,N_13349);
nand U13408 (N_13408,N_13326,N_13260);
xor U13409 (N_13409,N_13266,N_13278);
xor U13410 (N_13410,N_13258,N_13310);
nand U13411 (N_13411,N_13363,N_13321);
nand U13412 (N_13412,N_13352,N_13253);
and U13413 (N_13413,N_13298,N_13318);
xor U13414 (N_13414,N_13269,N_13279);
and U13415 (N_13415,N_13330,N_13262);
nor U13416 (N_13416,N_13297,N_13348);
nor U13417 (N_13417,N_13367,N_13255);
nor U13418 (N_13418,N_13354,N_13358);
or U13419 (N_13419,N_13261,N_13293);
or U13420 (N_13420,N_13331,N_13372);
and U13421 (N_13421,N_13308,N_13368);
nor U13422 (N_13422,N_13273,N_13305);
and U13423 (N_13423,N_13307,N_13259);
nor U13424 (N_13424,N_13350,N_13287);
or U13425 (N_13425,N_13328,N_13270);
xnor U13426 (N_13426,N_13257,N_13357);
or U13427 (N_13427,N_13295,N_13329);
xor U13428 (N_13428,N_13304,N_13373);
xnor U13429 (N_13429,N_13324,N_13369);
or U13430 (N_13430,N_13361,N_13362);
and U13431 (N_13431,N_13285,N_13341);
xnor U13432 (N_13432,N_13274,N_13374);
xnor U13433 (N_13433,N_13283,N_13332);
xnor U13434 (N_13434,N_13346,N_13254);
xor U13435 (N_13435,N_13276,N_13268);
and U13436 (N_13436,N_13336,N_13272);
xnor U13437 (N_13437,N_13342,N_13349);
nor U13438 (N_13438,N_13288,N_13294);
nand U13439 (N_13439,N_13363,N_13318);
and U13440 (N_13440,N_13340,N_13374);
xnor U13441 (N_13441,N_13348,N_13291);
and U13442 (N_13442,N_13366,N_13324);
xnor U13443 (N_13443,N_13316,N_13295);
nand U13444 (N_13444,N_13315,N_13304);
nand U13445 (N_13445,N_13273,N_13339);
nor U13446 (N_13446,N_13295,N_13346);
nand U13447 (N_13447,N_13281,N_13273);
nor U13448 (N_13448,N_13271,N_13331);
xor U13449 (N_13449,N_13272,N_13319);
and U13450 (N_13450,N_13277,N_13302);
and U13451 (N_13451,N_13292,N_13266);
nand U13452 (N_13452,N_13343,N_13274);
xor U13453 (N_13453,N_13344,N_13268);
xnor U13454 (N_13454,N_13364,N_13251);
and U13455 (N_13455,N_13331,N_13346);
nor U13456 (N_13456,N_13326,N_13297);
or U13457 (N_13457,N_13326,N_13308);
nand U13458 (N_13458,N_13323,N_13292);
and U13459 (N_13459,N_13366,N_13348);
xnor U13460 (N_13460,N_13358,N_13327);
and U13461 (N_13461,N_13270,N_13322);
or U13462 (N_13462,N_13261,N_13265);
xnor U13463 (N_13463,N_13371,N_13330);
or U13464 (N_13464,N_13310,N_13297);
nor U13465 (N_13465,N_13332,N_13351);
xnor U13466 (N_13466,N_13284,N_13356);
nor U13467 (N_13467,N_13355,N_13254);
nor U13468 (N_13468,N_13337,N_13338);
nor U13469 (N_13469,N_13274,N_13310);
or U13470 (N_13470,N_13301,N_13371);
xor U13471 (N_13471,N_13340,N_13261);
nand U13472 (N_13472,N_13262,N_13255);
xor U13473 (N_13473,N_13362,N_13269);
nand U13474 (N_13474,N_13299,N_13290);
xnor U13475 (N_13475,N_13345,N_13281);
xnor U13476 (N_13476,N_13337,N_13310);
or U13477 (N_13477,N_13278,N_13256);
and U13478 (N_13478,N_13318,N_13258);
nand U13479 (N_13479,N_13276,N_13334);
nor U13480 (N_13480,N_13335,N_13253);
nor U13481 (N_13481,N_13344,N_13271);
or U13482 (N_13482,N_13285,N_13289);
xor U13483 (N_13483,N_13296,N_13289);
xnor U13484 (N_13484,N_13321,N_13359);
nor U13485 (N_13485,N_13307,N_13331);
xnor U13486 (N_13486,N_13369,N_13350);
nor U13487 (N_13487,N_13361,N_13350);
and U13488 (N_13488,N_13321,N_13322);
and U13489 (N_13489,N_13297,N_13340);
nor U13490 (N_13490,N_13264,N_13318);
and U13491 (N_13491,N_13342,N_13326);
and U13492 (N_13492,N_13273,N_13307);
nor U13493 (N_13493,N_13298,N_13366);
or U13494 (N_13494,N_13338,N_13251);
or U13495 (N_13495,N_13371,N_13271);
nand U13496 (N_13496,N_13251,N_13269);
and U13497 (N_13497,N_13321,N_13272);
nor U13498 (N_13498,N_13256,N_13276);
and U13499 (N_13499,N_13353,N_13372);
xor U13500 (N_13500,N_13418,N_13386);
or U13501 (N_13501,N_13429,N_13471);
or U13502 (N_13502,N_13425,N_13492);
nor U13503 (N_13503,N_13484,N_13467);
or U13504 (N_13504,N_13480,N_13411);
nand U13505 (N_13505,N_13476,N_13451);
nor U13506 (N_13506,N_13376,N_13420);
and U13507 (N_13507,N_13479,N_13375);
xor U13508 (N_13508,N_13426,N_13460);
or U13509 (N_13509,N_13409,N_13398);
and U13510 (N_13510,N_13384,N_13434);
and U13511 (N_13511,N_13413,N_13452);
and U13512 (N_13512,N_13412,N_13483);
nor U13513 (N_13513,N_13441,N_13459);
nand U13514 (N_13514,N_13447,N_13446);
xnor U13515 (N_13515,N_13407,N_13481);
nor U13516 (N_13516,N_13475,N_13383);
nand U13517 (N_13517,N_13406,N_13472);
xor U13518 (N_13518,N_13443,N_13482);
xor U13519 (N_13519,N_13489,N_13419);
and U13520 (N_13520,N_13495,N_13458);
xor U13521 (N_13521,N_13401,N_13391);
and U13522 (N_13522,N_13448,N_13416);
nand U13523 (N_13523,N_13424,N_13485);
nand U13524 (N_13524,N_13498,N_13402);
and U13525 (N_13525,N_13437,N_13463);
or U13526 (N_13526,N_13497,N_13493);
nor U13527 (N_13527,N_13445,N_13450);
and U13528 (N_13528,N_13440,N_13410);
nor U13529 (N_13529,N_13496,N_13377);
nand U13530 (N_13530,N_13432,N_13455);
or U13531 (N_13531,N_13442,N_13408);
nor U13532 (N_13532,N_13385,N_13444);
and U13533 (N_13533,N_13393,N_13449);
xnor U13534 (N_13534,N_13387,N_13468);
or U13535 (N_13535,N_13473,N_13422);
nor U13536 (N_13536,N_13433,N_13474);
nand U13537 (N_13537,N_13453,N_13478);
or U13538 (N_13538,N_13494,N_13397);
nand U13539 (N_13539,N_13392,N_13469);
nand U13540 (N_13540,N_13487,N_13428);
xor U13541 (N_13541,N_13414,N_13404);
xor U13542 (N_13542,N_13415,N_13381);
nand U13543 (N_13543,N_13394,N_13390);
nor U13544 (N_13544,N_13396,N_13465);
nor U13545 (N_13545,N_13400,N_13430);
nor U13546 (N_13546,N_13499,N_13405);
nor U13547 (N_13547,N_13399,N_13403);
or U13548 (N_13548,N_13427,N_13438);
xnor U13549 (N_13549,N_13466,N_13380);
or U13550 (N_13550,N_13388,N_13477);
nand U13551 (N_13551,N_13423,N_13378);
or U13552 (N_13552,N_13382,N_13389);
xnor U13553 (N_13553,N_13486,N_13457);
or U13554 (N_13554,N_13431,N_13435);
or U13555 (N_13555,N_13436,N_13491);
nand U13556 (N_13556,N_13488,N_13470);
nor U13557 (N_13557,N_13454,N_13395);
and U13558 (N_13558,N_13379,N_13490);
xnor U13559 (N_13559,N_13464,N_13462);
and U13560 (N_13560,N_13439,N_13421);
nand U13561 (N_13561,N_13417,N_13461);
xor U13562 (N_13562,N_13456,N_13448);
nand U13563 (N_13563,N_13432,N_13435);
or U13564 (N_13564,N_13393,N_13485);
or U13565 (N_13565,N_13406,N_13466);
xnor U13566 (N_13566,N_13405,N_13396);
xnor U13567 (N_13567,N_13495,N_13499);
or U13568 (N_13568,N_13420,N_13446);
and U13569 (N_13569,N_13495,N_13417);
xnor U13570 (N_13570,N_13416,N_13462);
xor U13571 (N_13571,N_13450,N_13499);
xnor U13572 (N_13572,N_13382,N_13478);
xnor U13573 (N_13573,N_13401,N_13402);
nand U13574 (N_13574,N_13377,N_13493);
or U13575 (N_13575,N_13499,N_13407);
or U13576 (N_13576,N_13458,N_13437);
nand U13577 (N_13577,N_13424,N_13451);
nand U13578 (N_13578,N_13449,N_13429);
or U13579 (N_13579,N_13498,N_13405);
or U13580 (N_13580,N_13449,N_13459);
xnor U13581 (N_13581,N_13393,N_13389);
or U13582 (N_13582,N_13445,N_13449);
nand U13583 (N_13583,N_13404,N_13375);
and U13584 (N_13584,N_13434,N_13382);
and U13585 (N_13585,N_13479,N_13412);
or U13586 (N_13586,N_13383,N_13451);
or U13587 (N_13587,N_13435,N_13403);
xor U13588 (N_13588,N_13451,N_13459);
nand U13589 (N_13589,N_13461,N_13412);
and U13590 (N_13590,N_13423,N_13485);
or U13591 (N_13591,N_13432,N_13482);
nand U13592 (N_13592,N_13438,N_13494);
nor U13593 (N_13593,N_13474,N_13476);
or U13594 (N_13594,N_13442,N_13410);
or U13595 (N_13595,N_13419,N_13468);
or U13596 (N_13596,N_13442,N_13381);
or U13597 (N_13597,N_13452,N_13398);
nand U13598 (N_13598,N_13443,N_13429);
nor U13599 (N_13599,N_13493,N_13472);
or U13600 (N_13600,N_13401,N_13471);
nand U13601 (N_13601,N_13454,N_13467);
nor U13602 (N_13602,N_13376,N_13434);
and U13603 (N_13603,N_13385,N_13478);
nor U13604 (N_13604,N_13380,N_13445);
or U13605 (N_13605,N_13378,N_13485);
or U13606 (N_13606,N_13435,N_13472);
and U13607 (N_13607,N_13412,N_13471);
and U13608 (N_13608,N_13412,N_13423);
xor U13609 (N_13609,N_13488,N_13462);
or U13610 (N_13610,N_13460,N_13429);
xor U13611 (N_13611,N_13486,N_13378);
and U13612 (N_13612,N_13438,N_13416);
xnor U13613 (N_13613,N_13498,N_13399);
nor U13614 (N_13614,N_13381,N_13486);
xnor U13615 (N_13615,N_13454,N_13498);
nor U13616 (N_13616,N_13383,N_13457);
xnor U13617 (N_13617,N_13474,N_13402);
nor U13618 (N_13618,N_13461,N_13433);
nand U13619 (N_13619,N_13464,N_13414);
nand U13620 (N_13620,N_13494,N_13466);
nor U13621 (N_13621,N_13490,N_13403);
and U13622 (N_13622,N_13394,N_13467);
nor U13623 (N_13623,N_13399,N_13474);
and U13624 (N_13624,N_13423,N_13431);
nand U13625 (N_13625,N_13620,N_13604);
and U13626 (N_13626,N_13595,N_13569);
nand U13627 (N_13627,N_13599,N_13552);
or U13628 (N_13628,N_13566,N_13586);
nand U13629 (N_13629,N_13531,N_13536);
and U13630 (N_13630,N_13544,N_13590);
xnor U13631 (N_13631,N_13539,N_13543);
or U13632 (N_13632,N_13504,N_13613);
and U13633 (N_13633,N_13614,N_13572);
nor U13634 (N_13634,N_13580,N_13592);
and U13635 (N_13635,N_13502,N_13550);
nand U13636 (N_13636,N_13567,N_13583);
nor U13637 (N_13637,N_13579,N_13512);
nand U13638 (N_13638,N_13549,N_13616);
nand U13639 (N_13639,N_13621,N_13622);
nand U13640 (N_13640,N_13594,N_13582);
and U13641 (N_13641,N_13540,N_13612);
nand U13642 (N_13642,N_13603,N_13548);
and U13643 (N_13643,N_13578,N_13519);
and U13644 (N_13644,N_13522,N_13591);
nor U13645 (N_13645,N_13562,N_13505);
nand U13646 (N_13646,N_13551,N_13523);
nand U13647 (N_13647,N_13598,N_13568);
or U13648 (N_13648,N_13597,N_13518);
xor U13649 (N_13649,N_13556,N_13611);
and U13650 (N_13650,N_13596,N_13609);
and U13651 (N_13651,N_13624,N_13547);
nand U13652 (N_13652,N_13619,N_13601);
xnor U13653 (N_13653,N_13546,N_13506);
or U13654 (N_13654,N_13608,N_13517);
and U13655 (N_13655,N_13514,N_13513);
nand U13656 (N_13656,N_13585,N_13533);
nand U13657 (N_13657,N_13554,N_13529);
xnor U13658 (N_13658,N_13508,N_13526);
or U13659 (N_13659,N_13576,N_13617);
or U13660 (N_13660,N_13500,N_13538);
nor U13661 (N_13661,N_13535,N_13537);
or U13662 (N_13662,N_13593,N_13555);
or U13663 (N_13663,N_13581,N_13605);
and U13664 (N_13664,N_13516,N_13571);
xnor U13665 (N_13665,N_13524,N_13558);
nor U13666 (N_13666,N_13541,N_13557);
nor U13667 (N_13667,N_13606,N_13559);
nor U13668 (N_13668,N_13530,N_13563);
xor U13669 (N_13669,N_13525,N_13528);
or U13670 (N_13670,N_13618,N_13588);
nor U13671 (N_13671,N_13511,N_13509);
and U13672 (N_13672,N_13553,N_13573);
and U13673 (N_13673,N_13623,N_13534);
or U13674 (N_13674,N_13575,N_13542);
nand U13675 (N_13675,N_13600,N_13610);
and U13676 (N_13676,N_13565,N_13607);
xnor U13677 (N_13677,N_13532,N_13615);
nor U13678 (N_13678,N_13570,N_13507);
nor U13679 (N_13679,N_13602,N_13501);
and U13680 (N_13680,N_13510,N_13584);
nor U13681 (N_13681,N_13577,N_13527);
nor U13682 (N_13682,N_13503,N_13589);
nand U13683 (N_13683,N_13587,N_13520);
nand U13684 (N_13684,N_13515,N_13545);
nand U13685 (N_13685,N_13561,N_13564);
or U13686 (N_13686,N_13560,N_13521);
nand U13687 (N_13687,N_13574,N_13547);
nand U13688 (N_13688,N_13504,N_13523);
and U13689 (N_13689,N_13618,N_13579);
nand U13690 (N_13690,N_13584,N_13561);
nor U13691 (N_13691,N_13569,N_13602);
nand U13692 (N_13692,N_13617,N_13505);
nand U13693 (N_13693,N_13571,N_13535);
and U13694 (N_13694,N_13547,N_13535);
nor U13695 (N_13695,N_13518,N_13544);
and U13696 (N_13696,N_13559,N_13567);
or U13697 (N_13697,N_13521,N_13525);
xor U13698 (N_13698,N_13534,N_13561);
and U13699 (N_13699,N_13518,N_13615);
nor U13700 (N_13700,N_13521,N_13541);
and U13701 (N_13701,N_13531,N_13565);
or U13702 (N_13702,N_13537,N_13602);
nor U13703 (N_13703,N_13580,N_13550);
and U13704 (N_13704,N_13518,N_13582);
or U13705 (N_13705,N_13579,N_13511);
or U13706 (N_13706,N_13615,N_13561);
nand U13707 (N_13707,N_13585,N_13584);
nand U13708 (N_13708,N_13512,N_13551);
and U13709 (N_13709,N_13586,N_13591);
nand U13710 (N_13710,N_13541,N_13572);
or U13711 (N_13711,N_13524,N_13560);
nor U13712 (N_13712,N_13599,N_13601);
nor U13713 (N_13713,N_13553,N_13500);
nor U13714 (N_13714,N_13504,N_13542);
nand U13715 (N_13715,N_13619,N_13593);
xnor U13716 (N_13716,N_13525,N_13602);
or U13717 (N_13717,N_13559,N_13618);
nand U13718 (N_13718,N_13567,N_13618);
nand U13719 (N_13719,N_13505,N_13552);
nand U13720 (N_13720,N_13609,N_13605);
xor U13721 (N_13721,N_13577,N_13565);
nor U13722 (N_13722,N_13548,N_13611);
and U13723 (N_13723,N_13543,N_13544);
nor U13724 (N_13724,N_13526,N_13528);
and U13725 (N_13725,N_13513,N_13622);
or U13726 (N_13726,N_13531,N_13540);
nand U13727 (N_13727,N_13504,N_13531);
or U13728 (N_13728,N_13612,N_13613);
or U13729 (N_13729,N_13534,N_13565);
and U13730 (N_13730,N_13526,N_13572);
or U13731 (N_13731,N_13604,N_13611);
nor U13732 (N_13732,N_13507,N_13613);
and U13733 (N_13733,N_13610,N_13582);
and U13734 (N_13734,N_13619,N_13617);
and U13735 (N_13735,N_13598,N_13511);
and U13736 (N_13736,N_13518,N_13585);
or U13737 (N_13737,N_13515,N_13535);
nand U13738 (N_13738,N_13601,N_13501);
nand U13739 (N_13739,N_13507,N_13552);
or U13740 (N_13740,N_13508,N_13550);
xor U13741 (N_13741,N_13565,N_13519);
and U13742 (N_13742,N_13567,N_13551);
or U13743 (N_13743,N_13597,N_13552);
nand U13744 (N_13744,N_13585,N_13558);
and U13745 (N_13745,N_13540,N_13586);
xor U13746 (N_13746,N_13563,N_13579);
nand U13747 (N_13747,N_13524,N_13574);
nand U13748 (N_13748,N_13620,N_13619);
nor U13749 (N_13749,N_13522,N_13517);
or U13750 (N_13750,N_13741,N_13649);
nand U13751 (N_13751,N_13692,N_13643);
nand U13752 (N_13752,N_13689,N_13734);
xor U13753 (N_13753,N_13668,N_13642);
xnor U13754 (N_13754,N_13717,N_13666);
nor U13755 (N_13755,N_13742,N_13701);
and U13756 (N_13756,N_13627,N_13662);
and U13757 (N_13757,N_13735,N_13683);
nor U13758 (N_13758,N_13715,N_13625);
nand U13759 (N_13759,N_13638,N_13723);
or U13760 (N_13760,N_13675,N_13637);
nand U13761 (N_13761,N_13738,N_13660);
or U13762 (N_13762,N_13711,N_13646);
or U13763 (N_13763,N_13703,N_13740);
or U13764 (N_13764,N_13700,N_13631);
or U13765 (N_13765,N_13647,N_13640);
xnor U13766 (N_13766,N_13749,N_13710);
or U13767 (N_13767,N_13634,N_13746);
nor U13768 (N_13768,N_13733,N_13648);
xnor U13769 (N_13769,N_13714,N_13678);
nor U13770 (N_13770,N_13669,N_13665);
or U13771 (N_13771,N_13684,N_13667);
and U13772 (N_13772,N_13676,N_13626);
xor U13773 (N_13773,N_13636,N_13663);
nor U13774 (N_13774,N_13744,N_13645);
xor U13775 (N_13775,N_13629,N_13721);
nand U13776 (N_13776,N_13695,N_13687);
nor U13777 (N_13777,N_13658,N_13661);
xor U13778 (N_13778,N_13677,N_13718);
or U13779 (N_13779,N_13641,N_13664);
and U13780 (N_13780,N_13674,N_13747);
nand U13781 (N_13781,N_13697,N_13651);
nor U13782 (N_13782,N_13659,N_13730);
nand U13783 (N_13783,N_13632,N_13716);
xnor U13784 (N_13784,N_13727,N_13644);
nand U13785 (N_13785,N_13708,N_13705);
xnor U13786 (N_13786,N_13685,N_13639);
and U13787 (N_13787,N_13707,N_13709);
or U13788 (N_13788,N_13635,N_13737);
or U13789 (N_13789,N_13680,N_13686);
xor U13790 (N_13790,N_13688,N_13706);
nor U13791 (N_13791,N_13630,N_13691);
or U13792 (N_13792,N_13698,N_13724);
nand U13793 (N_13793,N_13743,N_13722);
and U13794 (N_13794,N_13650,N_13719);
xnor U13795 (N_13795,N_13671,N_13748);
or U13796 (N_13796,N_13693,N_13731);
or U13797 (N_13797,N_13628,N_13702);
nor U13798 (N_13798,N_13745,N_13657);
or U13799 (N_13799,N_13712,N_13655);
nand U13800 (N_13800,N_13725,N_13654);
and U13801 (N_13801,N_13652,N_13633);
xnor U13802 (N_13802,N_13726,N_13699);
and U13803 (N_13803,N_13728,N_13694);
nor U13804 (N_13804,N_13704,N_13653);
nor U13805 (N_13805,N_13682,N_13690);
or U13806 (N_13806,N_13679,N_13736);
nand U13807 (N_13807,N_13656,N_13681);
or U13808 (N_13808,N_13732,N_13739);
nand U13809 (N_13809,N_13729,N_13673);
xor U13810 (N_13810,N_13720,N_13670);
or U13811 (N_13811,N_13713,N_13696);
or U13812 (N_13812,N_13672,N_13679);
nor U13813 (N_13813,N_13646,N_13625);
and U13814 (N_13814,N_13713,N_13709);
xor U13815 (N_13815,N_13683,N_13704);
nand U13816 (N_13816,N_13682,N_13748);
and U13817 (N_13817,N_13681,N_13662);
nand U13818 (N_13818,N_13655,N_13703);
xor U13819 (N_13819,N_13736,N_13640);
and U13820 (N_13820,N_13633,N_13661);
or U13821 (N_13821,N_13711,N_13692);
or U13822 (N_13822,N_13723,N_13661);
and U13823 (N_13823,N_13710,N_13697);
nor U13824 (N_13824,N_13667,N_13666);
xnor U13825 (N_13825,N_13719,N_13734);
xor U13826 (N_13826,N_13658,N_13678);
or U13827 (N_13827,N_13670,N_13717);
nand U13828 (N_13828,N_13657,N_13669);
xnor U13829 (N_13829,N_13675,N_13693);
nor U13830 (N_13830,N_13648,N_13626);
xnor U13831 (N_13831,N_13696,N_13706);
or U13832 (N_13832,N_13708,N_13676);
or U13833 (N_13833,N_13747,N_13709);
xor U13834 (N_13834,N_13716,N_13663);
and U13835 (N_13835,N_13713,N_13653);
xor U13836 (N_13836,N_13678,N_13639);
nor U13837 (N_13837,N_13686,N_13718);
or U13838 (N_13838,N_13638,N_13733);
or U13839 (N_13839,N_13665,N_13675);
or U13840 (N_13840,N_13686,N_13681);
xnor U13841 (N_13841,N_13688,N_13744);
xnor U13842 (N_13842,N_13656,N_13648);
nor U13843 (N_13843,N_13676,N_13638);
or U13844 (N_13844,N_13680,N_13707);
xor U13845 (N_13845,N_13734,N_13646);
or U13846 (N_13846,N_13731,N_13697);
nand U13847 (N_13847,N_13674,N_13740);
xnor U13848 (N_13848,N_13687,N_13651);
nand U13849 (N_13849,N_13719,N_13630);
xnor U13850 (N_13850,N_13628,N_13714);
xor U13851 (N_13851,N_13691,N_13693);
nor U13852 (N_13852,N_13682,N_13683);
nand U13853 (N_13853,N_13743,N_13706);
nor U13854 (N_13854,N_13743,N_13638);
or U13855 (N_13855,N_13673,N_13629);
and U13856 (N_13856,N_13747,N_13705);
or U13857 (N_13857,N_13661,N_13645);
nand U13858 (N_13858,N_13645,N_13637);
and U13859 (N_13859,N_13657,N_13687);
nand U13860 (N_13860,N_13657,N_13731);
nor U13861 (N_13861,N_13665,N_13680);
and U13862 (N_13862,N_13654,N_13710);
and U13863 (N_13863,N_13716,N_13711);
xor U13864 (N_13864,N_13666,N_13748);
nand U13865 (N_13865,N_13636,N_13691);
nand U13866 (N_13866,N_13728,N_13640);
xnor U13867 (N_13867,N_13659,N_13706);
xor U13868 (N_13868,N_13678,N_13632);
or U13869 (N_13869,N_13648,N_13676);
nor U13870 (N_13870,N_13671,N_13731);
nor U13871 (N_13871,N_13630,N_13693);
or U13872 (N_13872,N_13665,N_13635);
xor U13873 (N_13873,N_13681,N_13701);
xor U13874 (N_13874,N_13746,N_13701);
xnor U13875 (N_13875,N_13756,N_13771);
xnor U13876 (N_13876,N_13755,N_13782);
nand U13877 (N_13877,N_13846,N_13809);
xor U13878 (N_13878,N_13830,N_13753);
nor U13879 (N_13879,N_13844,N_13777);
nand U13880 (N_13880,N_13867,N_13869);
nand U13881 (N_13881,N_13849,N_13852);
nand U13882 (N_13882,N_13770,N_13870);
nand U13883 (N_13883,N_13833,N_13776);
xor U13884 (N_13884,N_13750,N_13874);
xnor U13885 (N_13885,N_13807,N_13847);
nor U13886 (N_13886,N_13765,N_13864);
nor U13887 (N_13887,N_13805,N_13797);
and U13888 (N_13888,N_13783,N_13803);
nor U13889 (N_13889,N_13779,N_13780);
or U13890 (N_13890,N_13822,N_13812);
nor U13891 (N_13891,N_13793,N_13813);
and U13892 (N_13892,N_13834,N_13860);
or U13893 (N_13893,N_13856,N_13866);
nand U13894 (N_13894,N_13759,N_13837);
nand U13895 (N_13895,N_13775,N_13804);
xnor U13896 (N_13896,N_13766,N_13819);
xor U13897 (N_13897,N_13845,N_13840);
xnor U13898 (N_13898,N_13778,N_13773);
or U13899 (N_13899,N_13788,N_13752);
and U13900 (N_13900,N_13761,N_13832);
nor U13901 (N_13901,N_13763,N_13826);
nor U13902 (N_13902,N_13854,N_13810);
xor U13903 (N_13903,N_13787,N_13814);
or U13904 (N_13904,N_13858,N_13796);
xnor U13905 (N_13905,N_13769,N_13784);
or U13906 (N_13906,N_13789,N_13873);
xor U13907 (N_13907,N_13872,N_13808);
and U13908 (N_13908,N_13758,N_13800);
or U13909 (N_13909,N_13848,N_13859);
nand U13910 (N_13910,N_13855,N_13839);
nand U13911 (N_13911,N_13843,N_13825);
xor U13912 (N_13912,N_13863,N_13768);
and U13913 (N_13913,N_13801,N_13790);
or U13914 (N_13914,N_13853,N_13836);
xor U13915 (N_13915,N_13827,N_13831);
nand U13916 (N_13916,N_13751,N_13786);
nor U13917 (N_13917,N_13767,N_13850);
nor U13918 (N_13918,N_13861,N_13760);
nand U13919 (N_13919,N_13757,N_13841);
nand U13920 (N_13920,N_13871,N_13811);
nand U13921 (N_13921,N_13838,N_13785);
nand U13922 (N_13922,N_13806,N_13815);
nand U13923 (N_13923,N_13791,N_13823);
or U13924 (N_13924,N_13798,N_13802);
or U13925 (N_13925,N_13817,N_13818);
nor U13926 (N_13926,N_13835,N_13865);
and U13927 (N_13927,N_13799,N_13820);
nor U13928 (N_13928,N_13821,N_13868);
xor U13929 (N_13929,N_13764,N_13774);
nand U13930 (N_13930,N_13772,N_13816);
xnor U13931 (N_13931,N_13842,N_13851);
nand U13932 (N_13932,N_13781,N_13754);
nand U13933 (N_13933,N_13795,N_13762);
or U13934 (N_13934,N_13824,N_13862);
or U13935 (N_13935,N_13829,N_13792);
or U13936 (N_13936,N_13857,N_13828);
nand U13937 (N_13937,N_13794,N_13831);
and U13938 (N_13938,N_13769,N_13821);
or U13939 (N_13939,N_13783,N_13851);
nor U13940 (N_13940,N_13755,N_13812);
nand U13941 (N_13941,N_13849,N_13810);
nor U13942 (N_13942,N_13853,N_13869);
and U13943 (N_13943,N_13797,N_13861);
nor U13944 (N_13944,N_13874,N_13857);
and U13945 (N_13945,N_13860,N_13807);
xor U13946 (N_13946,N_13846,N_13768);
nor U13947 (N_13947,N_13792,N_13844);
nor U13948 (N_13948,N_13784,N_13873);
or U13949 (N_13949,N_13810,N_13758);
and U13950 (N_13950,N_13806,N_13866);
nand U13951 (N_13951,N_13795,N_13791);
or U13952 (N_13952,N_13786,N_13752);
and U13953 (N_13953,N_13785,N_13861);
or U13954 (N_13954,N_13778,N_13770);
nand U13955 (N_13955,N_13863,N_13776);
and U13956 (N_13956,N_13839,N_13810);
and U13957 (N_13957,N_13871,N_13859);
or U13958 (N_13958,N_13801,N_13775);
nand U13959 (N_13959,N_13857,N_13794);
nor U13960 (N_13960,N_13839,N_13847);
nand U13961 (N_13961,N_13774,N_13755);
nand U13962 (N_13962,N_13816,N_13855);
nand U13963 (N_13963,N_13845,N_13837);
nor U13964 (N_13964,N_13755,N_13868);
and U13965 (N_13965,N_13844,N_13842);
xor U13966 (N_13966,N_13807,N_13804);
xor U13967 (N_13967,N_13821,N_13777);
or U13968 (N_13968,N_13823,N_13846);
or U13969 (N_13969,N_13763,N_13866);
nor U13970 (N_13970,N_13841,N_13772);
nand U13971 (N_13971,N_13751,N_13846);
and U13972 (N_13972,N_13752,N_13857);
nand U13973 (N_13973,N_13792,N_13780);
and U13974 (N_13974,N_13847,N_13818);
and U13975 (N_13975,N_13754,N_13871);
nor U13976 (N_13976,N_13793,N_13799);
nand U13977 (N_13977,N_13751,N_13810);
or U13978 (N_13978,N_13767,N_13771);
nand U13979 (N_13979,N_13871,N_13807);
or U13980 (N_13980,N_13862,N_13859);
or U13981 (N_13981,N_13846,N_13787);
or U13982 (N_13982,N_13841,N_13794);
nand U13983 (N_13983,N_13825,N_13829);
xnor U13984 (N_13984,N_13859,N_13752);
xor U13985 (N_13985,N_13828,N_13767);
nor U13986 (N_13986,N_13863,N_13855);
or U13987 (N_13987,N_13837,N_13816);
nor U13988 (N_13988,N_13776,N_13810);
nor U13989 (N_13989,N_13774,N_13870);
or U13990 (N_13990,N_13780,N_13773);
nand U13991 (N_13991,N_13851,N_13814);
or U13992 (N_13992,N_13792,N_13872);
nand U13993 (N_13993,N_13859,N_13844);
xnor U13994 (N_13994,N_13756,N_13753);
or U13995 (N_13995,N_13782,N_13786);
nand U13996 (N_13996,N_13864,N_13848);
nand U13997 (N_13997,N_13798,N_13760);
nor U13998 (N_13998,N_13837,N_13861);
nand U13999 (N_13999,N_13791,N_13754);
xnor U14000 (N_14000,N_13902,N_13909);
nor U14001 (N_14001,N_13968,N_13895);
and U14002 (N_14002,N_13990,N_13992);
and U14003 (N_14003,N_13999,N_13965);
nor U14004 (N_14004,N_13919,N_13914);
xnor U14005 (N_14005,N_13967,N_13916);
nand U14006 (N_14006,N_13945,N_13917);
nand U14007 (N_14007,N_13948,N_13882);
nand U14008 (N_14008,N_13982,N_13986);
nor U14009 (N_14009,N_13994,N_13924);
nand U14010 (N_14010,N_13877,N_13953);
nand U14011 (N_14011,N_13946,N_13906);
xnor U14012 (N_14012,N_13957,N_13960);
or U14013 (N_14013,N_13971,N_13905);
xor U14014 (N_14014,N_13884,N_13941);
nor U14015 (N_14015,N_13911,N_13883);
or U14016 (N_14016,N_13937,N_13981);
xor U14017 (N_14017,N_13983,N_13977);
and U14018 (N_14018,N_13897,N_13880);
xnor U14019 (N_14019,N_13942,N_13975);
or U14020 (N_14020,N_13940,N_13943);
or U14021 (N_14021,N_13993,N_13956);
or U14022 (N_14022,N_13961,N_13875);
nand U14023 (N_14023,N_13972,N_13913);
or U14024 (N_14024,N_13889,N_13944);
or U14025 (N_14025,N_13952,N_13927);
nor U14026 (N_14026,N_13932,N_13947);
and U14027 (N_14027,N_13885,N_13959);
and U14028 (N_14028,N_13915,N_13984);
xor U14029 (N_14029,N_13939,N_13923);
or U14030 (N_14030,N_13996,N_13962);
nand U14031 (N_14031,N_13963,N_13966);
or U14032 (N_14032,N_13998,N_13886);
nor U14033 (N_14033,N_13893,N_13876);
xnor U14034 (N_14034,N_13938,N_13979);
or U14035 (N_14035,N_13991,N_13925);
xnor U14036 (N_14036,N_13955,N_13910);
and U14037 (N_14037,N_13907,N_13903);
nand U14038 (N_14038,N_13951,N_13989);
nand U14039 (N_14039,N_13890,N_13934);
nand U14040 (N_14040,N_13929,N_13958);
or U14041 (N_14041,N_13995,N_13949);
nand U14042 (N_14042,N_13980,N_13888);
xor U14043 (N_14043,N_13904,N_13988);
or U14044 (N_14044,N_13930,N_13928);
xnor U14045 (N_14045,N_13922,N_13918);
nand U14046 (N_14046,N_13936,N_13900);
xor U14047 (N_14047,N_13935,N_13964);
or U14048 (N_14048,N_13978,N_13954);
nand U14049 (N_14049,N_13921,N_13896);
nand U14050 (N_14050,N_13892,N_13879);
xor U14051 (N_14051,N_13912,N_13976);
xnor U14052 (N_14052,N_13985,N_13881);
nor U14053 (N_14053,N_13920,N_13926);
nand U14054 (N_14054,N_13894,N_13987);
nand U14055 (N_14055,N_13901,N_13899);
xnor U14056 (N_14056,N_13950,N_13970);
or U14057 (N_14057,N_13973,N_13878);
xnor U14058 (N_14058,N_13908,N_13933);
xor U14059 (N_14059,N_13931,N_13997);
xnor U14060 (N_14060,N_13887,N_13974);
xnor U14061 (N_14061,N_13898,N_13969);
xor U14062 (N_14062,N_13891,N_13893);
and U14063 (N_14063,N_13898,N_13888);
nand U14064 (N_14064,N_13880,N_13982);
nand U14065 (N_14065,N_13987,N_13970);
or U14066 (N_14066,N_13877,N_13898);
nand U14067 (N_14067,N_13927,N_13986);
and U14068 (N_14068,N_13965,N_13986);
or U14069 (N_14069,N_13876,N_13894);
xnor U14070 (N_14070,N_13941,N_13929);
xnor U14071 (N_14071,N_13954,N_13983);
nor U14072 (N_14072,N_13953,N_13898);
nand U14073 (N_14073,N_13929,N_13928);
and U14074 (N_14074,N_13879,N_13949);
nor U14075 (N_14075,N_13939,N_13950);
xor U14076 (N_14076,N_13979,N_13990);
nor U14077 (N_14077,N_13905,N_13940);
nand U14078 (N_14078,N_13886,N_13935);
nand U14079 (N_14079,N_13969,N_13954);
and U14080 (N_14080,N_13896,N_13910);
nand U14081 (N_14081,N_13963,N_13984);
nor U14082 (N_14082,N_13904,N_13892);
nor U14083 (N_14083,N_13954,N_13893);
or U14084 (N_14084,N_13936,N_13925);
nand U14085 (N_14085,N_13967,N_13891);
nor U14086 (N_14086,N_13928,N_13972);
and U14087 (N_14087,N_13918,N_13953);
or U14088 (N_14088,N_13931,N_13976);
and U14089 (N_14089,N_13934,N_13896);
and U14090 (N_14090,N_13926,N_13915);
or U14091 (N_14091,N_13909,N_13986);
and U14092 (N_14092,N_13941,N_13947);
nand U14093 (N_14093,N_13938,N_13966);
or U14094 (N_14094,N_13996,N_13926);
xnor U14095 (N_14095,N_13917,N_13978);
and U14096 (N_14096,N_13959,N_13966);
nand U14097 (N_14097,N_13923,N_13943);
xor U14098 (N_14098,N_13890,N_13882);
and U14099 (N_14099,N_13972,N_13877);
nand U14100 (N_14100,N_13927,N_13946);
nand U14101 (N_14101,N_13991,N_13957);
xnor U14102 (N_14102,N_13984,N_13979);
nand U14103 (N_14103,N_13908,N_13991);
or U14104 (N_14104,N_13966,N_13945);
xor U14105 (N_14105,N_13913,N_13968);
or U14106 (N_14106,N_13990,N_13936);
nor U14107 (N_14107,N_13943,N_13934);
or U14108 (N_14108,N_13927,N_13963);
or U14109 (N_14109,N_13875,N_13996);
xor U14110 (N_14110,N_13969,N_13891);
and U14111 (N_14111,N_13952,N_13945);
or U14112 (N_14112,N_13980,N_13909);
and U14113 (N_14113,N_13955,N_13887);
nand U14114 (N_14114,N_13989,N_13877);
and U14115 (N_14115,N_13899,N_13927);
xor U14116 (N_14116,N_13906,N_13947);
nor U14117 (N_14117,N_13878,N_13917);
nor U14118 (N_14118,N_13919,N_13881);
nand U14119 (N_14119,N_13897,N_13926);
xnor U14120 (N_14120,N_13922,N_13967);
and U14121 (N_14121,N_13963,N_13883);
nand U14122 (N_14122,N_13937,N_13964);
nor U14123 (N_14123,N_13886,N_13946);
or U14124 (N_14124,N_13905,N_13908);
nor U14125 (N_14125,N_14024,N_14095);
nor U14126 (N_14126,N_14080,N_14113);
and U14127 (N_14127,N_14104,N_14012);
nand U14128 (N_14128,N_14021,N_14056);
or U14129 (N_14129,N_14034,N_14057);
and U14130 (N_14130,N_14002,N_14118);
and U14131 (N_14131,N_14026,N_14058);
and U14132 (N_14132,N_14003,N_14008);
xor U14133 (N_14133,N_14000,N_14105);
or U14134 (N_14134,N_14007,N_14018);
or U14135 (N_14135,N_14098,N_14040);
nand U14136 (N_14136,N_14072,N_14088);
and U14137 (N_14137,N_14044,N_14090);
or U14138 (N_14138,N_14038,N_14089);
nor U14139 (N_14139,N_14049,N_14087);
xnor U14140 (N_14140,N_14081,N_14096);
and U14141 (N_14141,N_14083,N_14102);
or U14142 (N_14142,N_14063,N_14020);
and U14143 (N_14143,N_14070,N_14108);
xnor U14144 (N_14144,N_14116,N_14101);
or U14145 (N_14145,N_14065,N_14027);
nand U14146 (N_14146,N_14062,N_14009);
and U14147 (N_14147,N_14100,N_14053);
xor U14148 (N_14148,N_14015,N_14120);
or U14149 (N_14149,N_14112,N_14097);
nor U14150 (N_14150,N_14050,N_14029);
nor U14151 (N_14151,N_14051,N_14022);
or U14152 (N_14152,N_14006,N_14066);
nor U14153 (N_14153,N_14041,N_14093);
or U14154 (N_14154,N_14061,N_14091);
and U14155 (N_14155,N_14059,N_14075);
nand U14156 (N_14156,N_14025,N_14117);
xor U14157 (N_14157,N_14030,N_14111);
nand U14158 (N_14158,N_14033,N_14019);
xnor U14159 (N_14159,N_14010,N_14121);
or U14160 (N_14160,N_14067,N_14122);
or U14161 (N_14161,N_14043,N_14076);
or U14162 (N_14162,N_14068,N_14013);
or U14163 (N_14163,N_14077,N_14109);
and U14164 (N_14164,N_14047,N_14103);
and U14165 (N_14165,N_14124,N_14079);
xnor U14166 (N_14166,N_14054,N_14036);
nand U14167 (N_14167,N_14052,N_14085);
nand U14168 (N_14168,N_14046,N_14069);
xor U14169 (N_14169,N_14055,N_14028);
nor U14170 (N_14170,N_14073,N_14074);
and U14171 (N_14171,N_14016,N_14119);
nand U14172 (N_14172,N_14064,N_14107);
nor U14173 (N_14173,N_14115,N_14123);
nor U14174 (N_14174,N_14110,N_14078);
nor U14175 (N_14175,N_14060,N_14042);
nor U14176 (N_14176,N_14039,N_14084);
xor U14177 (N_14177,N_14071,N_14023);
xor U14178 (N_14178,N_14106,N_14114);
nor U14179 (N_14179,N_14014,N_14099);
xor U14180 (N_14180,N_14032,N_14005);
xor U14181 (N_14181,N_14092,N_14035);
nand U14182 (N_14182,N_14031,N_14082);
and U14183 (N_14183,N_14017,N_14001);
and U14184 (N_14184,N_14004,N_14037);
nor U14185 (N_14185,N_14094,N_14086);
nor U14186 (N_14186,N_14045,N_14048);
nand U14187 (N_14187,N_14011,N_14048);
nand U14188 (N_14188,N_14091,N_14059);
and U14189 (N_14189,N_14082,N_14007);
nand U14190 (N_14190,N_14016,N_14066);
and U14191 (N_14191,N_14074,N_14032);
and U14192 (N_14192,N_14049,N_14068);
nor U14193 (N_14193,N_14048,N_14070);
or U14194 (N_14194,N_14040,N_14074);
nor U14195 (N_14195,N_14007,N_14113);
or U14196 (N_14196,N_14044,N_14038);
or U14197 (N_14197,N_14005,N_14057);
or U14198 (N_14198,N_14026,N_14079);
nor U14199 (N_14199,N_14051,N_14120);
or U14200 (N_14200,N_14026,N_14033);
nor U14201 (N_14201,N_14026,N_14076);
xor U14202 (N_14202,N_14049,N_14013);
and U14203 (N_14203,N_14041,N_14105);
xnor U14204 (N_14204,N_14088,N_14010);
xor U14205 (N_14205,N_14056,N_14075);
or U14206 (N_14206,N_14103,N_14010);
nor U14207 (N_14207,N_14078,N_14091);
xnor U14208 (N_14208,N_14012,N_14065);
xnor U14209 (N_14209,N_14013,N_14035);
nand U14210 (N_14210,N_14121,N_14114);
and U14211 (N_14211,N_14061,N_14090);
nand U14212 (N_14212,N_14124,N_14109);
xor U14213 (N_14213,N_14070,N_14004);
nand U14214 (N_14214,N_14058,N_14053);
xor U14215 (N_14215,N_14040,N_14035);
and U14216 (N_14216,N_14100,N_14076);
nand U14217 (N_14217,N_14002,N_14041);
nand U14218 (N_14218,N_14082,N_14061);
xor U14219 (N_14219,N_14075,N_14112);
and U14220 (N_14220,N_14079,N_14110);
xnor U14221 (N_14221,N_14048,N_14030);
or U14222 (N_14222,N_14077,N_14124);
nand U14223 (N_14223,N_14114,N_14064);
nor U14224 (N_14224,N_14048,N_14021);
xor U14225 (N_14225,N_14120,N_14036);
nor U14226 (N_14226,N_14070,N_14059);
and U14227 (N_14227,N_14039,N_14023);
or U14228 (N_14228,N_14000,N_14017);
and U14229 (N_14229,N_14078,N_14117);
and U14230 (N_14230,N_14067,N_14042);
nor U14231 (N_14231,N_14073,N_14004);
nand U14232 (N_14232,N_14002,N_14054);
or U14233 (N_14233,N_14106,N_14034);
nand U14234 (N_14234,N_14051,N_14121);
nor U14235 (N_14235,N_14108,N_14067);
nand U14236 (N_14236,N_14015,N_14011);
or U14237 (N_14237,N_14015,N_14067);
xnor U14238 (N_14238,N_14044,N_14020);
nand U14239 (N_14239,N_14001,N_14028);
and U14240 (N_14240,N_14120,N_14039);
and U14241 (N_14241,N_14051,N_14100);
nor U14242 (N_14242,N_14059,N_14049);
and U14243 (N_14243,N_14100,N_14059);
or U14244 (N_14244,N_14100,N_14044);
nand U14245 (N_14245,N_14016,N_14099);
or U14246 (N_14246,N_14010,N_14033);
and U14247 (N_14247,N_14000,N_14107);
xnor U14248 (N_14248,N_14080,N_14069);
and U14249 (N_14249,N_14121,N_14064);
nor U14250 (N_14250,N_14192,N_14229);
and U14251 (N_14251,N_14226,N_14210);
and U14252 (N_14252,N_14184,N_14198);
and U14253 (N_14253,N_14154,N_14178);
xor U14254 (N_14254,N_14130,N_14180);
nor U14255 (N_14255,N_14141,N_14225);
nand U14256 (N_14256,N_14245,N_14230);
and U14257 (N_14257,N_14214,N_14126);
or U14258 (N_14258,N_14211,N_14191);
or U14259 (N_14259,N_14157,N_14162);
and U14260 (N_14260,N_14139,N_14216);
nor U14261 (N_14261,N_14167,N_14146);
nor U14262 (N_14262,N_14238,N_14196);
nand U14263 (N_14263,N_14248,N_14143);
nor U14264 (N_14264,N_14161,N_14246);
and U14265 (N_14265,N_14175,N_14235);
or U14266 (N_14266,N_14159,N_14204);
and U14267 (N_14267,N_14125,N_14170);
nor U14268 (N_14268,N_14131,N_14165);
xor U14269 (N_14269,N_14205,N_14247);
nor U14270 (N_14270,N_14183,N_14249);
nor U14271 (N_14271,N_14176,N_14222);
and U14272 (N_14272,N_14213,N_14138);
and U14273 (N_14273,N_14231,N_14243);
xnor U14274 (N_14274,N_14197,N_14151);
nor U14275 (N_14275,N_14163,N_14177);
nor U14276 (N_14276,N_14145,N_14134);
and U14277 (N_14277,N_14187,N_14241);
nor U14278 (N_14278,N_14158,N_14148);
nor U14279 (N_14279,N_14228,N_14149);
and U14280 (N_14280,N_14215,N_14206);
and U14281 (N_14281,N_14239,N_14224);
nor U14282 (N_14282,N_14174,N_14142);
nor U14283 (N_14283,N_14227,N_14144);
nor U14284 (N_14284,N_14153,N_14212);
and U14285 (N_14285,N_14240,N_14169);
xor U14286 (N_14286,N_14242,N_14171);
nor U14287 (N_14287,N_14166,N_14218);
xnor U14288 (N_14288,N_14193,N_14127);
nand U14289 (N_14289,N_14137,N_14190);
nor U14290 (N_14290,N_14173,N_14182);
xnor U14291 (N_14291,N_14164,N_14133);
and U14292 (N_14292,N_14244,N_14155);
xor U14293 (N_14293,N_14150,N_14189);
nor U14294 (N_14294,N_14203,N_14207);
or U14295 (N_14295,N_14129,N_14199);
and U14296 (N_14296,N_14140,N_14217);
or U14297 (N_14297,N_14219,N_14136);
xnor U14298 (N_14298,N_14128,N_14208);
xor U14299 (N_14299,N_14234,N_14201);
xor U14300 (N_14300,N_14172,N_14233);
and U14301 (N_14301,N_14186,N_14168);
and U14302 (N_14302,N_14147,N_14188);
and U14303 (N_14303,N_14209,N_14232);
xnor U14304 (N_14304,N_14221,N_14132);
nor U14305 (N_14305,N_14185,N_14220);
or U14306 (N_14306,N_14152,N_14195);
nor U14307 (N_14307,N_14237,N_14179);
nor U14308 (N_14308,N_14202,N_14160);
nor U14309 (N_14309,N_14194,N_14156);
nand U14310 (N_14310,N_14135,N_14236);
nand U14311 (N_14311,N_14200,N_14223);
nand U14312 (N_14312,N_14181,N_14221);
or U14313 (N_14313,N_14166,N_14192);
and U14314 (N_14314,N_14173,N_14131);
or U14315 (N_14315,N_14214,N_14174);
or U14316 (N_14316,N_14248,N_14184);
or U14317 (N_14317,N_14170,N_14180);
xnor U14318 (N_14318,N_14206,N_14216);
nor U14319 (N_14319,N_14219,N_14235);
xor U14320 (N_14320,N_14125,N_14246);
nand U14321 (N_14321,N_14162,N_14206);
nor U14322 (N_14322,N_14222,N_14193);
nand U14323 (N_14323,N_14209,N_14230);
and U14324 (N_14324,N_14207,N_14135);
or U14325 (N_14325,N_14166,N_14238);
nand U14326 (N_14326,N_14175,N_14246);
and U14327 (N_14327,N_14224,N_14191);
xnor U14328 (N_14328,N_14216,N_14237);
and U14329 (N_14329,N_14136,N_14196);
xor U14330 (N_14330,N_14180,N_14193);
or U14331 (N_14331,N_14169,N_14185);
nor U14332 (N_14332,N_14138,N_14201);
or U14333 (N_14333,N_14202,N_14178);
and U14334 (N_14334,N_14160,N_14243);
xnor U14335 (N_14335,N_14125,N_14141);
or U14336 (N_14336,N_14197,N_14248);
nand U14337 (N_14337,N_14229,N_14249);
and U14338 (N_14338,N_14191,N_14139);
xnor U14339 (N_14339,N_14131,N_14194);
nor U14340 (N_14340,N_14233,N_14147);
xor U14341 (N_14341,N_14204,N_14165);
xor U14342 (N_14342,N_14181,N_14148);
nor U14343 (N_14343,N_14139,N_14208);
or U14344 (N_14344,N_14236,N_14204);
nand U14345 (N_14345,N_14134,N_14235);
and U14346 (N_14346,N_14236,N_14158);
or U14347 (N_14347,N_14221,N_14186);
and U14348 (N_14348,N_14149,N_14227);
or U14349 (N_14349,N_14187,N_14196);
xnor U14350 (N_14350,N_14135,N_14169);
xnor U14351 (N_14351,N_14139,N_14200);
or U14352 (N_14352,N_14213,N_14197);
nand U14353 (N_14353,N_14173,N_14197);
xor U14354 (N_14354,N_14156,N_14165);
or U14355 (N_14355,N_14128,N_14228);
xor U14356 (N_14356,N_14232,N_14154);
nand U14357 (N_14357,N_14134,N_14180);
nand U14358 (N_14358,N_14126,N_14234);
nor U14359 (N_14359,N_14225,N_14232);
xor U14360 (N_14360,N_14217,N_14243);
nand U14361 (N_14361,N_14151,N_14127);
nand U14362 (N_14362,N_14221,N_14173);
nand U14363 (N_14363,N_14236,N_14217);
or U14364 (N_14364,N_14234,N_14182);
and U14365 (N_14365,N_14132,N_14191);
xnor U14366 (N_14366,N_14210,N_14237);
nor U14367 (N_14367,N_14159,N_14229);
xor U14368 (N_14368,N_14151,N_14205);
or U14369 (N_14369,N_14187,N_14227);
nand U14370 (N_14370,N_14127,N_14237);
nor U14371 (N_14371,N_14195,N_14223);
nand U14372 (N_14372,N_14174,N_14134);
or U14373 (N_14373,N_14248,N_14198);
nand U14374 (N_14374,N_14242,N_14198);
nor U14375 (N_14375,N_14324,N_14360);
nor U14376 (N_14376,N_14297,N_14358);
or U14377 (N_14377,N_14274,N_14333);
nand U14378 (N_14378,N_14361,N_14321);
or U14379 (N_14379,N_14289,N_14264);
and U14380 (N_14380,N_14294,N_14349);
nand U14381 (N_14381,N_14364,N_14296);
and U14382 (N_14382,N_14266,N_14320);
or U14383 (N_14383,N_14263,N_14254);
nor U14384 (N_14384,N_14312,N_14292);
xnor U14385 (N_14385,N_14268,N_14287);
xor U14386 (N_14386,N_14257,N_14332);
and U14387 (N_14387,N_14348,N_14314);
or U14388 (N_14388,N_14347,N_14340);
or U14389 (N_14389,N_14372,N_14305);
nand U14390 (N_14390,N_14295,N_14369);
nand U14391 (N_14391,N_14354,N_14319);
and U14392 (N_14392,N_14350,N_14288);
nor U14393 (N_14393,N_14346,N_14286);
xor U14394 (N_14394,N_14273,N_14325);
xnor U14395 (N_14395,N_14276,N_14265);
or U14396 (N_14396,N_14258,N_14281);
nor U14397 (N_14397,N_14278,N_14302);
nand U14398 (N_14398,N_14303,N_14251);
xor U14399 (N_14399,N_14341,N_14363);
or U14400 (N_14400,N_14367,N_14301);
and U14401 (N_14401,N_14366,N_14271);
xor U14402 (N_14402,N_14374,N_14262);
and U14403 (N_14403,N_14343,N_14261);
and U14404 (N_14404,N_14315,N_14269);
or U14405 (N_14405,N_14282,N_14309);
or U14406 (N_14406,N_14352,N_14290);
or U14407 (N_14407,N_14368,N_14357);
or U14408 (N_14408,N_14291,N_14250);
nand U14409 (N_14409,N_14318,N_14356);
nor U14410 (N_14410,N_14284,N_14370);
and U14411 (N_14411,N_14277,N_14344);
or U14412 (N_14412,N_14300,N_14353);
xor U14413 (N_14413,N_14283,N_14373);
or U14414 (N_14414,N_14280,N_14316);
xor U14415 (N_14415,N_14342,N_14362);
or U14416 (N_14416,N_14256,N_14253);
xnor U14417 (N_14417,N_14313,N_14336);
or U14418 (N_14418,N_14308,N_14328);
nand U14419 (N_14419,N_14311,N_14267);
xor U14420 (N_14420,N_14326,N_14331);
and U14421 (N_14421,N_14310,N_14260);
and U14422 (N_14422,N_14323,N_14293);
nand U14423 (N_14423,N_14272,N_14327);
xor U14424 (N_14424,N_14307,N_14351);
xnor U14425 (N_14425,N_14359,N_14285);
or U14426 (N_14426,N_14329,N_14306);
xor U14427 (N_14427,N_14279,N_14317);
nand U14428 (N_14428,N_14330,N_14299);
or U14429 (N_14429,N_14339,N_14275);
nand U14430 (N_14430,N_14334,N_14270);
and U14431 (N_14431,N_14371,N_14355);
xnor U14432 (N_14432,N_14337,N_14252);
xnor U14433 (N_14433,N_14304,N_14335);
or U14434 (N_14434,N_14338,N_14365);
xor U14435 (N_14435,N_14345,N_14259);
nand U14436 (N_14436,N_14322,N_14298);
or U14437 (N_14437,N_14255,N_14262);
or U14438 (N_14438,N_14327,N_14356);
nand U14439 (N_14439,N_14308,N_14294);
nor U14440 (N_14440,N_14252,N_14251);
nor U14441 (N_14441,N_14330,N_14293);
xor U14442 (N_14442,N_14362,N_14300);
nor U14443 (N_14443,N_14295,N_14320);
and U14444 (N_14444,N_14290,N_14331);
xor U14445 (N_14445,N_14327,N_14349);
or U14446 (N_14446,N_14298,N_14290);
nand U14447 (N_14447,N_14276,N_14277);
xor U14448 (N_14448,N_14335,N_14313);
xor U14449 (N_14449,N_14369,N_14254);
and U14450 (N_14450,N_14316,N_14300);
nand U14451 (N_14451,N_14273,N_14336);
or U14452 (N_14452,N_14336,N_14253);
and U14453 (N_14453,N_14259,N_14268);
xor U14454 (N_14454,N_14291,N_14360);
nand U14455 (N_14455,N_14308,N_14275);
or U14456 (N_14456,N_14345,N_14289);
nand U14457 (N_14457,N_14281,N_14324);
nand U14458 (N_14458,N_14289,N_14298);
or U14459 (N_14459,N_14312,N_14296);
xor U14460 (N_14460,N_14269,N_14292);
xor U14461 (N_14461,N_14317,N_14326);
and U14462 (N_14462,N_14296,N_14367);
nor U14463 (N_14463,N_14320,N_14278);
nor U14464 (N_14464,N_14277,N_14259);
or U14465 (N_14465,N_14372,N_14294);
xnor U14466 (N_14466,N_14344,N_14286);
xor U14467 (N_14467,N_14316,N_14365);
nor U14468 (N_14468,N_14250,N_14351);
nor U14469 (N_14469,N_14341,N_14310);
nor U14470 (N_14470,N_14309,N_14258);
xor U14471 (N_14471,N_14261,N_14270);
nand U14472 (N_14472,N_14289,N_14341);
xor U14473 (N_14473,N_14305,N_14253);
nand U14474 (N_14474,N_14305,N_14274);
and U14475 (N_14475,N_14372,N_14369);
and U14476 (N_14476,N_14370,N_14307);
xor U14477 (N_14477,N_14368,N_14361);
nand U14478 (N_14478,N_14274,N_14357);
nor U14479 (N_14479,N_14344,N_14334);
nor U14480 (N_14480,N_14355,N_14278);
and U14481 (N_14481,N_14336,N_14298);
and U14482 (N_14482,N_14344,N_14262);
nand U14483 (N_14483,N_14359,N_14330);
nor U14484 (N_14484,N_14271,N_14332);
nand U14485 (N_14485,N_14310,N_14256);
or U14486 (N_14486,N_14303,N_14278);
nor U14487 (N_14487,N_14326,N_14294);
or U14488 (N_14488,N_14319,N_14347);
or U14489 (N_14489,N_14319,N_14274);
or U14490 (N_14490,N_14274,N_14292);
xor U14491 (N_14491,N_14278,N_14342);
and U14492 (N_14492,N_14270,N_14346);
xnor U14493 (N_14493,N_14281,N_14337);
nor U14494 (N_14494,N_14283,N_14324);
or U14495 (N_14495,N_14314,N_14344);
xnor U14496 (N_14496,N_14372,N_14276);
or U14497 (N_14497,N_14284,N_14295);
nor U14498 (N_14498,N_14272,N_14366);
nor U14499 (N_14499,N_14332,N_14305);
nor U14500 (N_14500,N_14499,N_14417);
nand U14501 (N_14501,N_14446,N_14426);
or U14502 (N_14502,N_14424,N_14403);
and U14503 (N_14503,N_14421,N_14404);
xor U14504 (N_14504,N_14447,N_14420);
nor U14505 (N_14505,N_14431,N_14414);
nand U14506 (N_14506,N_14493,N_14449);
nand U14507 (N_14507,N_14472,N_14380);
nand U14508 (N_14508,N_14445,N_14425);
xnor U14509 (N_14509,N_14413,N_14397);
nand U14510 (N_14510,N_14456,N_14443);
or U14511 (N_14511,N_14415,N_14455);
xor U14512 (N_14512,N_14393,N_14379);
or U14513 (N_14513,N_14440,N_14383);
or U14514 (N_14514,N_14468,N_14460);
or U14515 (N_14515,N_14432,N_14450);
or U14516 (N_14516,N_14395,N_14427);
nand U14517 (N_14517,N_14444,N_14390);
xor U14518 (N_14518,N_14489,N_14469);
nor U14519 (N_14519,N_14448,N_14490);
xor U14520 (N_14520,N_14485,N_14461);
nor U14521 (N_14521,N_14465,N_14408);
xor U14522 (N_14522,N_14452,N_14451);
or U14523 (N_14523,N_14410,N_14478);
xor U14524 (N_14524,N_14406,N_14480);
and U14525 (N_14525,N_14459,N_14392);
or U14526 (N_14526,N_14387,N_14418);
nand U14527 (N_14527,N_14439,N_14492);
or U14528 (N_14528,N_14384,N_14441);
nand U14529 (N_14529,N_14385,N_14442);
nor U14530 (N_14530,N_14496,N_14399);
and U14531 (N_14531,N_14400,N_14389);
or U14532 (N_14532,N_14388,N_14474);
or U14533 (N_14533,N_14467,N_14470);
or U14534 (N_14534,N_14476,N_14454);
nand U14535 (N_14535,N_14464,N_14463);
and U14536 (N_14536,N_14436,N_14433);
and U14537 (N_14537,N_14428,N_14473);
nand U14538 (N_14538,N_14484,N_14405);
or U14539 (N_14539,N_14401,N_14494);
nor U14540 (N_14540,N_14495,N_14416);
nor U14541 (N_14541,N_14423,N_14412);
and U14542 (N_14542,N_14377,N_14497);
or U14543 (N_14543,N_14477,N_14458);
or U14544 (N_14544,N_14419,N_14375);
xor U14545 (N_14545,N_14483,N_14498);
xnor U14546 (N_14546,N_14491,N_14471);
xnor U14547 (N_14547,N_14429,N_14396);
nor U14548 (N_14548,N_14486,N_14453);
xor U14549 (N_14549,N_14430,N_14434);
or U14550 (N_14550,N_14457,N_14407);
and U14551 (N_14551,N_14411,N_14402);
or U14552 (N_14552,N_14386,N_14378);
xnor U14553 (N_14553,N_14437,N_14479);
or U14554 (N_14554,N_14409,N_14462);
nand U14555 (N_14555,N_14466,N_14438);
or U14556 (N_14556,N_14488,N_14398);
or U14557 (N_14557,N_14475,N_14422);
nand U14558 (N_14558,N_14394,N_14381);
nand U14559 (N_14559,N_14482,N_14391);
nor U14560 (N_14560,N_14382,N_14487);
and U14561 (N_14561,N_14376,N_14481);
xnor U14562 (N_14562,N_14435,N_14449);
or U14563 (N_14563,N_14463,N_14376);
xor U14564 (N_14564,N_14404,N_14486);
nand U14565 (N_14565,N_14474,N_14386);
or U14566 (N_14566,N_14411,N_14401);
nor U14567 (N_14567,N_14381,N_14412);
and U14568 (N_14568,N_14483,N_14460);
xnor U14569 (N_14569,N_14430,N_14445);
xnor U14570 (N_14570,N_14461,N_14382);
or U14571 (N_14571,N_14451,N_14495);
nand U14572 (N_14572,N_14473,N_14425);
xnor U14573 (N_14573,N_14392,N_14475);
and U14574 (N_14574,N_14454,N_14385);
or U14575 (N_14575,N_14428,N_14444);
nand U14576 (N_14576,N_14395,N_14440);
nor U14577 (N_14577,N_14486,N_14489);
or U14578 (N_14578,N_14468,N_14444);
nand U14579 (N_14579,N_14474,N_14447);
and U14580 (N_14580,N_14485,N_14465);
xnor U14581 (N_14581,N_14434,N_14493);
xor U14582 (N_14582,N_14491,N_14465);
xnor U14583 (N_14583,N_14472,N_14435);
nor U14584 (N_14584,N_14493,N_14452);
and U14585 (N_14585,N_14423,N_14456);
or U14586 (N_14586,N_14497,N_14418);
and U14587 (N_14587,N_14474,N_14487);
nor U14588 (N_14588,N_14387,N_14467);
nand U14589 (N_14589,N_14436,N_14418);
or U14590 (N_14590,N_14441,N_14430);
nand U14591 (N_14591,N_14440,N_14463);
nor U14592 (N_14592,N_14451,N_14423);
nor U14593 (N_14593,N_14479,N_14491);
nor U14594 (N_14594,N_14432,N_14491);
nor U14595 (N_14595,N_14456,N_14388);
and U14596 (N_14596,N_14394,N_14398);
or U14597 (N_14597,N_14397,N_14375);
or U14598 (N_14598,N_14412,N_14414);
nor U14599 (N_14599,N_14412,N_14446);
nor U14600 (N_14600,N_14422,N_14446);
xor U14601 (N_14601,N_14468,N_14410);
nor U14602 (N_14602,N_14439,N_14408);
nand U14603 (N_14603,N_14454,N_14487);
xor U14604 (N_14604,N_14419,N_14385);
xor U14605 (N_14605,N_14420,N_14495);
xnor U14606 (N_14606,N_14490,N_14441);
or U14607 (N_14607,N_14435,N_14484);
nand U14608 (N_14608,N_14424,N_14484);
xor U14609 (N_14609,N_14407,N_14432);
or U14610 (N_14610,N_14415,N_14425);
nand U14611 (N_14611,N_14411,N_14428);
nor U14612 (N_14612,N_14425,N_14404);
xnor U14613 (N_14613,N_14499,N_14493);
nor U14614 (N_14614,N_14472,N_14400);
nand U14615 (N_14615,N_14460,N_14390);
and U14616 (N_14616,N_14463,N_14442);
nor U14617 (N_14617,N_14381,N_14388);
xor U14618 (N_14618,N_14406,N_14388);
or U14619 (N_14619,N_14417,N_14388);
nand U14620 (N_14620,N_14463,N_14490);
and U14621 (N_14621,N_14376,N_14416);
xor U14622 (N_14622,N_14383,N_14385);
and U14623 (N_14623,N_14384,N_14426);
xnor U14624 (N_14624,N_14481,N_14408);
nand U14625 (N_14625,N_14570,N_14569);
and U14626 (N_14626,N_14541,N_14522);
or U14627 (N_14627,N_14562,N_14539);
xor U14628 (N_14628,N_14502,N_14533);
or U14629 (N_14629,N_14538,N_14587);
and U14630 (N_14630,N_14528,N_14503);
xor U14631 (N_14631,N_14555,N_14515);
xor U14632 (N_14632,N_14506,N_14607);
xnor U14633 (N_14633,N_14512,N_14610);
and U14634 (N_14634,N_14589,N_14558);
nand U14635 (N_14635,N_14606,N_14573);
nor U14636 (N_14636,N_14575,N_14580);
nor U14637 (N_14637,N_14585,N_14521);
nor U14638 (N_14638,N_14596,N_14611);
and U14639 (N_14639,N_14553,N_14540);
and U14640 (N_14640,N_14513,N_14508);
nor U14641 (N_14641,N_14561,N_14590);
nand U14642 (N_14642,N_14586,N_14516);
nand U14643 (N_14643,N_14615,N_14602);
nand U14644 (N_14644,N_14604,N_14603);
and U14645 (N_14645,N_14544,N_14517);
nand U14646 (N_14646,N_14621,N_14595);
xor U14647 (N_14647,N_14614,N_14574);
nand U14648 (N_14648,N_14601,N_14529);
or U14649 (N_14649,N_14549,N_14520);
xnor U14650 (N_14650,N_14609,N_14592);
nor U14651 (N_14651,N_14619,N_14551);
nor U14652 (N_14652,N_14598,N_14524);
or U14653 (N_14653,N_14500,N_14552);
or U14654 (N_14654,N_14501,N_14545);
and U14655 (N_14655,N_14554,N_14616);
nor U14656 (N_14656,N_14568,N_14618);
and U14657 (N_14657,N_14523,N_14608);
xor U14658 (N_14658,N_14526,N_14566);
and U14659 (N_14659,N_14505,N_14594);
and U14660 (N_14660,N_14559,N_14563);
nand U14661 (N_14661,N_14557,N_14530);
nor U14662 (N_14662,N_14532,N_14507);
nand U14663 (N_14663,N_14593,N_14536);
and U14664 (N_14664,N_14600,N_14542);
or U14665 (N_14665,N_14620,N_14577);
xor U14666 (N_14666,N_14583,N_14556);
nor U14667 (N_14667,N_14548,N_14504);
or U14668 (N_14668,N_14576,N_14612);
nor U14669 (N_14669,N_14514,N_14582);
and U14670 (N_14670,N_14546,N_14550);
or U14671 (N_14671,N_14560,N_14518);
or U14672 (N_14672,N_14547,N_14509);
nor U14673 (N_14673,N_14591,N_14537);
or U14674 (N_14674,N_14565,N_14613);
nand U14675 (N_14675,N_14605,N_14564);
xor U14676 (N_14676,N_14510,N_14623);
or U14677 (N_14677,N_14579,N_14617);
nor U14678 (N_14678,N_14578,N_14535);
nand U14679 (N_14679,N_14599,N_14622);
or U14680 (N_14680,N_14588,N_14567);
and U14681 (N_14681,N_14525,N_14584);
xor U14682 (N_14682,N_14511,N_14581);
nor U14683 (N_14683,N_14543,N_14519);
and U14684 (N_14684,N_14534,N_14571);
or U14685 (N_14685,N_14597,N_14527);
nand U14686 (N_14686,N_14531,N_14624);
and U14687 (N_14687,N_14572,N_14609);
or U14688 (N_14688,N_14573,N_14610);
or U14689 (N_14689,N_14578,N_14597);
xor U14690 (N_14690,N_14537,N_14595);
xor U14691 (N_14691,N_14541,N_14581);
nor U14692 (N_14692,N_14543,N_14605);
and U14693 (N_14693,N_14511,N_14509);
nor U14694 (N_14694,N_14510,N_14527);
nand U14695 (N_14695,N_14569,N_14560);
or U14696 (N_14696,N_14518,N_14519);
or U14697 (N_14697,N_14622,N_14558);
xor U14698 (N_14698,N_14525,N_14621);
nor U14699 (N_14699,N_14610,N_14500);
nand U14700 (N_14700,N_14597,N_14541);
and U14701 (N_14701,N_14560,N_14607);
xnor U14702 (N_14702,N_14542,N_14553);
and U14703 (N_14703,N_14575,N_14591);
and U14704 (N_14704,N_14529,N_14532);
nor U14705 (N_14705,N_14597,N_14570);
and U14706 (N_14706,N_14528,N_14606);
nor U14707 (N_14707,N_14520,N_14603);
nand U14708 (N_14708,N_14502,N_14582);
nor U14709 (N_14709,N_14603,N_14581);
and U14710 (N_14710,N_14535,N_14547);
and U14711 (N_14711,N_14508,N_14574);
nand U14712 (N_14712,N_14519,N_14560);
and U14713 (N_14713,N_14561,N_14610);
or U14714 (N_14714,N_14536,N_14586);
nor U14715 (N_14715,N_14504,N_14542);
nor U14716 (N_14716,N_14571,N_14547);
and U14717 (N_14717,N_14551,N_14527);
xnor U14718 (N_14718,N_14559,N_14565);
xor U14719 (N_14719,N_14574,N_14607);
nor U14720 (N_14720,N_14621,N_14601);
nand U14721 (N_14721,N_14616,N_14531);
nor U14722 (N_14722,N_14578,N_14575);
and U14723 (N_14723,N_14568,N_14563);
and U14724 (N_14724,N_14623,N_14567);
xor U14725 (N_14725,N_14530,N_14600);
xor U14726 (N_14726,N_14526,N_14591);
and U14727 (N_14727,N_14537,N_14511);
nor U14728 (N_14728,N_14554,N_14511);
xor U14729 (N_14729,N_14587,N_14606);
xnor U14730 (N_14730,N_14506,N_14612);
or U14731 (N_14731,N_14536,N_14508);
nand U14732 (N_14732,N_14520,N_14510);
and U14733 (N_14733,N_14589,N_14586);
or U14734 (N_14734,N_14509,N_14587);
xnor U14735 (N_14735,N_14526,N_14505);
and U14736 (N_14736,N_14526,N_14550);
and U14737 (N_14737,N_14558,N_14531);
nand U14738 (N_14738,N_14505,N_14536);
and U14739 (N_14739,N_14566,N_14537);
nor U14740 (N_14740,N_14560,N_14621);
nor U14741 (N_14741,N_14503,N_14586);
and U14742 (N_14742,N_14535,N_14501);
or U14743 (N_14743,N_14524,N_14538);
nor U14744 (N_14744,N_14555,N_14593);
nand U14745 (N_14745,N_14531,N_14537);
nor U14746 (N_14746,N_14539,N_14578);
and U14747 (N_14747,N_14523,N_14551);
and U14748 (N_14748,N_14601,N_14566);
or U14749 (N_14749,N_14553,N_14557);
nand U14750 (N_14750,N_14651,N_14688);
nor U14751 (N_14751,N_14662,N_14635);
nand U14752 (N_14752,N_14681,N_14630);
xnor U14753 (N_14753,N_14728,N_14653);
or U14754 (N_14754,N_14671,N_14652);
nand U14755 (N_14755,N_14697,N_14737);
xnor U14756 (N_14756,N_14684,N_14740);
nand U14757 (N_14757,N_14720,N_14736);
and U14758 (N_14758,N_14704,N_14699);
and U14759 (N_14759,N_14747,N_14655);
xor U14760 (N_14760,N_14717,N_14746);
nand U14761 (N_14761,N_14649,N_14659);
xnor U14762 (N_14762,N_14660,N_14705);
and U14763 (N_14763,N_14647,N_14643);
nor U14764 (N_14764,N_14644,N_14679);
nand U14765 (N_14765,N_14636,N_14708);
nand U14766 (N_14766,N_14666,N_14725);
or U14767 (N_14767,N_14709,N_14631);
xor U14768 (N_14768,N_14689,N_14673);
nand U14769 (N_14769,N_14661,N_14626);
and U14770 (N_14770,N_14743,N_14748);
xnor U14771 (N_14771,N_14641,N_14744);
xor U14772 (N_14772,N_14718,N_14731);
or U14773 (N_14773,N_14658,N_14739);
or U14774 (N_14774,N_14698,N_14675);
nor U14775 (N_14775,N_14721,N_14634);
or U14776 (N_14776,N_14654,N_14707);
xor U14777 (N_14777,N_14719,N_14686);
nor U14778 (N_14778,N_14713,N_14642);
or U14779 (N_14779,N_14678,N_14742);
nand U14780 (N_14780,N_14669,N_14648);
or U14781 (N_14781,N_14700,N_14638);
xor U14782 (N_14782,N_14667,N_14637);
or U14783 (N_14783,N_14745,N_14682);
nor U14784 (N_14784,N_14702,N_14665);
nand U14785 (N_14785,N_14646,N_14711);
xor U14786 (N_14786,N_14732,N_14628);
and U14787 (N_14787,N_14735,N_14625);
nand U14788 (N_14788,N_14693,N_14695);
nor U14789 (N_14789,N_14672,N_14677);
nor U14790 (N_14790,N_14687,N_14656);
or U14791 (N_14791,N_14724,N_14680);
or U14792 (N_14792,N_14632,N_14629);
and U14793 (N_14793,N_14710,N_14650);
or U14794 (N_14794,N_14727,N_14701);
or U14795 (N_14795,N_14674,N_14639);
xor U14796 (N_14796,N_14726,N_14664);
xnor U14797 (N_14797,N_14722,N_14714);
and U14798 (N_14798,N_14663,N_14668);
nand U14799 (N_14799,N_14676,N_14691);
or U14800 (N_14800,N_14670,N_14696);
and U14801 (N_14801,N_14692,N_14627);
nand U14802 (N_14802,N_14633,N_14729);
nand U14803 (N_14803,N_14734,N_14706);
nand U14804 (N_14804,N_14645,N_14694);
nand U14805 (N_14805,N_14741,N_14690);
nor U14806 (N_14806,N_14723,N_14685);
xnor U14807 (N_14807,N_14715,N_14712);
nor U14808 (N_14808,N_14738,N_14657);
or U14809 (N_14809,N_14733,N_14640);
xor U14810 (N_14810,N_14730,N_14716);
xnor U14811 (N_14811,N_14749,N_14703);
or U14812 (N_14812,N_14683,N_14715);
or U14813 (N_14813,N_14683,N_14719);
nor U14814 (N_14814,N_14734,N_14732);
or U14815 (N_14815,N_14627,N_14635);
xnor U14816 (N_14816,N_14712,N_14742);
and U14817 (N_14817,N_14675,N_14721);
nand U14818 (N_14818,N_14643,N_14668);
or U14819 (N_14819,N_14688,N_14743);
nor U14820 (N_14820,N_14714,N_14744);
nor U14821 (N_14821,N_14636,N_14740);
and U14822 (N_14822,N_14675,N_14690);
nor U14823 (N_14823,N_14679,N_14664);
or U14824 (N_14824,N_14688,N_14734);
and U14825 (N_14825,N_14625,N_14668);
nand U14826 (N_14826,N_14729,N_14631);
and U14827 (N_14827,N_14654,N_14635);
nand U14828 (N_14828,N_14718,N_14719);
and U14829 (N_14829,N_14701,N_14732);
or U14830 (N_14830,N_14648,N_14732);
nor U14831 (N_14831,N_14637,N_14695);
nand U14832 (N_14832,N_14661,N_14628);
xnor U14833 (N_14833,N_14683,N_14664);
and U14834 (N_14834,N_14714,N_14716);
nor U14835 (N_14835,N_14687,N_14642);
nor U14836 (N_14836,N_14715,N_14716);
xnor U14837 (N_14837,N_14722,N_14680);
and U14838 (N_14838,N_14714,N_14733);
nand U14839 (N_14839,N_14636,N_14635);
nand U14840 (N_14840,N_14679,N_14637);
nand U14841 (N_14841,N_14649,N_14666);
xor U14842 (N_14842,N_14706,N_14639);
nor U14843 (N_14843,N_14703,N_14739);
nor U14844 (N_14844,N_14745,N_14675);
and U14845 (N_14845,N_14698,N_14656);
nor U14846 (N_14846,N_14657,N_14667);
nor U14847 (N_14847,N_14625,N_14677);
and U14848 (N_14848,N_14730,N_14696);
nand U14849 (N_14849,N_14739,N_14713);
or U14850 (N_14850,N_14640,N_14697);
nand U14851 (N_14851,N_14659,N_14648);
or U14852 (N_14852,N_14670,N_14649);
or U14853 (N_14853,N_14652,N_14738);
nand U14854 (N_14854,N_14648,N_14689);
nand U14855 (N_14855,N_14630,N_14653);
or U14856 (N_14856,N_14727,N_14692);
xor U14857 (N_14857,N_14626,N_14639);
xor U14858 (N_14858,N_14719,N_14680);
nor U14859 (N_14859,N_14639,N_14676);
nand U14860 (N_14860,N_14647,N_14665);
or U14861 (N_14861,N_14647,N_14646);
and U14862 (N_14862,N_14729,N_14663);
and U14863 (N_14863,N_14731,N_14632);
xor U14864 (N_14864,N_14628,N_14686);
or U14865 (N_14865,N_14630,N_14675);
or U14866 (N_14866,N_14671,N_14676);
nor U14867 (N_14867,N_14706,N_14705);
xnor U14868 (N_14868,N_14646,N_14717);
and U14869 (N_14869,N_14677,N_14745);
and U14870 (N_14870,N_14684,N_14728);
and U14871 (N_14871,N_14634,N_14678);
and U14872 (N_14872,N_14720,N_14632);
or U14873 (N_14873,N_14669,N_14687);
or U14874 (N_14874,N_14682,N_14629);
nor U14875 (N_14875,N_14758,N_14835);
nor U14876 (N_14876,N_14803,N_14836);
and U14877 (N_14877,N_14869,N_14857);
nor U14878 (N_14878,N_14839,N_14785);
nand U14879 (N_14879,N_14787,N_14872);
xnor U14880 (N_14880,N_14853,N_14778);
or U14881 (N_14881,N_14865,N_14811);
nand U14882 (N_14882,N_14783,N_14757);
nand U14883 (N_14883,N_14826,N_14855);
or U14884 (N_14884,N_14780,N_14838);
and U14885 (N_14885,N_14786,N_14792);
and U14886 (N_14886,N_14847,N_14788);
xnor U14887 (N_14887,N_14799,N_14795);
and U14888 (N_14888,N_14751,N_14790);
nor U14889 (N_14889,N_14779,N_14831);
or U14890 (N_14890,N_14837,N_14784);
xor U14891 (N_14891,N_14762,N_14764);
nand U14892 (N_14892,N_14770,N_14761);
or U14893 (N_14893,N_14775,N_14793);
nor U14894 (N_14894,N_14796,N_14767);
and U14895 (N_14895,N_14804,N_14871);
or U14896 (N_14896,N_14794,N_14812);
or U14897 (N_14897,N_14813,N_14829);
nand U14898 (N_14898,N_14858,N_14769);
and U14899 (N_14899,N_14854,N_14830);
nor U14900 (N_14900,N_14773,N_14861);
xor U14901 (N_14901,N_14859,N_14874);
and U14902 (N_14902,N_14798,N_14810);
nand U14903 (N_14903,N_14862,N_14846);
and U14904 (N_14904,N_14800,N_14821);
nor U14905 (N_14905,N_14819,N_14772);
xor U14906 (N_14906,N_14833,N_14817);
nand U14907 (N_14907,N_14848,N_14873);
or U14908 (N_14908,N_14852,N_14844);
xor U14909 (N_14909,N_14755,N_14791);
xor U14910 (N_14910,N_14774,N_14809);
xor U14911 (N_14911,N_14824,N_14849);
nand U14912 (N_14912,N_14822,N_14864);
xor U14913 (N_14913,N_14860,N_14805);
nand U14914 (N_14914,N_14856,N_14789);
nor U14915 (N_14915,N_14814,N_14782);
xnor U14916 (N_14916,N_14806,N_14818);
nor U14917 (N_14917,N_14827,N_14825);
and U14918 (N_14918,N_14820,N_14766);
or U14919 (N_14919,N_14808,N_14834);
nand U14920 (N_14920,N_14867,N_14753);
or U14921 (N_14921,N_14828,N_14850);
nor U14922 (N_14922,N_14750,N_14756);
nand U14923 (N_14923,N_14807,N_14752);
nand U14924 (N_14924,N_14781,N_14866);
xnor U14925 (N_14925,N_14801,N_14765);
nor U14926 (N_14926,N_14768,N_14863);
nand U14927 (N_14927,N_14754,N_14760);
xor U14928 (N_14928,N_14841,N_14840);
and U14929 (N_14929,N_14851,N_14776);
or U14930 (N_14930,N_14823,N_14816);
xor U14931 (N_14931,N_14777,N_14868);
nand U14932 (N_14932,N_14763,N_14842);
and U14933 (N_14933,N_14870,N_14845);
nand U14934 (N_14934,N_14843,N_14759);
xnor U14935 (N_14935,N_14832,N_14797);
or U14936 (N_14936,N_14802,N_14771);
xnor U14937 (N_14937,N_14815,N_14828);
and U14938 (N_14938,N_14757,N_14838);
nor U14939 (N_14939,N_14855,N_14850);
or U14940 (N_14940,N_14785,N_14813);
nand U14941 (N_14941,N_14843,N_14856);
nand U14942 (N_14942,N_14821,N_14757);
xor U14943 (N_14943,N_14854,N_14763);
nand U14944 (N_14944,N_14859,N_14772);
nor U14945 (N_14945,N_14868,N_14810);
nor U14946 (N_14946,N_14806,N_14809);
xor U14947 (N_14947,N_14865,N_14814);
nand U14948 (N_14948,N_14860,N_14775);
or U14949 (N_14949,N_14842,N_14861);
xor U14950 (N_14950,N_14843,N_14858);
and U14951 (N_14951,N_14782,N_14840);
nand U14952 (N_14952,N_14833,N_14784);
xor U14953 (N_14953,N_14797,N_14751);
xnor U14954 (N_14954,N_14865,N_14782);
or U14955 (N_14955,N_14752,N_14872);
nand U14956 (N_14956,N_14864,N_14765);
nor U14957 (N_14957,N_14796,N_14869);
or U14958 (N_14958,N_14763,N_14864);
and U14959 (N_14959,N_14832,N_14849);
xnor U14960 (N_14960,N_14852,N_14838);
nand U14961 (N_14961,N_14841,N_14837);
xor U14962 (N_14962,N_14855,N_14810);
nor U14963 (N_14963,N_14859,N_14770);
and U14964 (N_14964,N_14818,N_14827);
nor U14965 (N_14965,N_14833,N_14846);
or U14966 (N_14966,N_14764,N_14867);
and U14967 (N_14967,N_14819,N_14804);
nor U14968 (N_14968,N_14780,N_14870);
nand U14969 (N_14969,N_14800,N_14802);
or U14970 (N_14970,N_14769,N_14838);
and U14971 (N_14971,N_14751,N_14795);
nor U14972 (N_14972,N_14821,N_14750);
nor U14973 (N_14973,N_14790,N_14854);
and U14974 (N_14974,N_14772,N_14789);
nor U14975 (N_14975,N_14802,N_14837);
or U14976 (N_14976,N_14751,N_14826);
xor U14977 (N_14977,N_14846,N_14796);
or U14978 (N_14978,N_14801,N_14824);
nand U14979 (N_14979,N_14865,N_14847);
or U14980 (N_14980,N_14865,N_14830);
nor U14981 (N_14981,N_14804,N_14859);
or U14982 (N_14982,N_14856,N_14865);
or U14983 (N_14983,N_14847,N_14772);
nor U14984 (N_14984,N_14842,N_14857);
xor U14985 (N_14985,N_14774,N_14832);
or U14986 (N_14986,N_14831,N_14813);
or U14987 (N_14987,N_14761,N_14753);
nor U14988 (N_14988,N_14813,N_14778);
xnor U14989 (N_14989,N_14858,N_14820);
nand U14990 (N_14990,N_14819,N_14870);
or U14991 (N_14991,N_14805,N_14775);
nand U14992 (N_14992,N_14806,N_14785);
nor U14993 (N_14993,N_14817,N_14769);
and U14994 (N_14994,N_14839,N_14794);
nor U14995 (N_14995,N_14776,N_14852);
nand U14996 (N_14996,N_14811,N_14854);
xor U14997 (N_14997,N_14785,N_14807);
nand U14998 (N_14998,N_14785,N_14768);
nand U14999 (N_14999,N_14802,N_14868);
nand UO_0 (O_0,N_14950,N_14905);
nand UO_1 (O_1,N_14932,N_14890);
and UO_2 (O_2,N_14981,N_14955);
xnor UO_3 (O_3,N_14945,N_14893);
nand UO_4 (O_4,N_14991,N_14973);
xnor UO_5 (O_5,N_14883,N_14988);
or UO_6 (O_6,N_14938,N_14910);
or UO_7 (O_7,N_14923,N_14976);
nor UO_8 (O_8,N_14913,N_14954);
or UO_9 (O_9,N_14901,N_14990);
nor UO_10 (O_10,N_14898,N_14989);
xnor UO_11 (O_11,N_14939,N_14980);
and UO_12 (O_12,N_14878,N_14982);
nor UO_13 (O_13,N_14891,N_14907);
or UO_14 (O_14,N_14902,N_14953);
and UO_15 (O_15,N_14975,N_14935);
and UO_16 (O_16,N_14969,N_14904);
or UO_17 (O_17,N_14962,N_14992);
nand UO_18 (O_18,N_14925,N_14900);
and UO_19 (O_19,N_14963,N_14978);
and UO_20 (O_20,N_14877,N_14952);
xor UO_21 (O_21,N_14931,N_14959);
and UO_22 (O_22,N_14972,N_14944);
nand UO_23 (O_23,N_14940,N_14974);
nand UO_24 (O_24,N_14934,N_14886);
xnor UO_25 (O_25,N_14911,N_14968);
nor UO_26 (O_26,N_14929,N_14876);
nand UO_27 (O_27,N_14996,N_14983);
and UO_28 (O_28,N_14998,N_14994);
and UO_29 (O_29,N_14958,N_14930);
xor UO_30 (O_30,N_14894,N_14916);
nor UO_31 (O_31,N_14896,N_14951);
nand UO_32 (O_32,N_14933,N_14920);
nand UO_33 (O_33,N_14906,N_14879);
nand UO_34 (O_34,N_14888,N_14899);
xor UO_35 (O_35,N_14915,N_14942);
nor UO_36 (O_36,N_14947,N_14943);
nor UO_37 (O_37,N_14971,N_14964);
nor UO_38 (O_38,N_14927,N_14922);
nand UO_39 (O_39,N_14882,N_14887);
nand UO_40 (O_40,N_14914,N_14997);
xor UO_41 (O_41,N_14961,N_14881);
nor UO_42 (O_42,N_14875,N_14924);
nand UO_43 (O_43,N_14895,N_14937);
xnor UO_44 (O_44,N_14912,N_14987);
nor UO_45 (O_45,N_14949,N_14948);
or UO_46 (O_46,N_14909,N_14880);
and UO_47 (O_47,N_14903,N_14941);
or UO_48 (O_48,N_14921,N_14885);
xnor UO_49 (O_49,N_14884,N_14889);
nand UO_50 (O_50,N_14936,N_14977);
nand UO_51 (O_51,N_14966,N_14979);
nor UO_52 (O_52,N_14919,N_14999);
and UO_53 (O_53,N_14897,N_14984);
xnor UO_54 (O_54,N_14970,N_14917);
and UO_55 (O_55,N_14908,N_14960);
or UO_56 (O_56,N_14946,N_14993);
and UO_57 (O_57,N_14985,N_14967);
and UO_58 (O_58,N_14986,N_14956);
or UO_59 (O_59,N_14995,N_14965);
xnor UO_60 (O_60,N_14918,N_14926);
xnor UO_61 (O_61,N_14928,N_14892);
or UO_62 (O_62,N_14957,N_14983);
nand UO_63 (O_63,N_14923,N_14891);
or UO_64 (O_64,N_14903,N_14898);
or UO_65 (O_65,N_14961,N_14953);
and UO_66 (O_66,N_14916,N_14914);
nand UO_67 (O_67,N_14931,N_14920);
nor UO_68 (O_68,N_14907,N_14938);
nand UO_69 (O_69,N_14935,N_14989);
or UO_70 (O_70,N_14999,N_14895);
or UO_71 (O_71,N_14938,N_14926);
or UO_72 (O_72,N_14896,N_14997);
xnor UO_73 (O_73,N_14982,N_14908);
or UO_74 (O_74,N_14902,N_14982);
xnor UO_75 (O_75,N_14925,N_14927);
or UO_76 (O_76,N_14960,N_14901);
nand UO_77 (O_77,N_14954,N_14947);
or UO_78 (O_78,N_14977,N_14927);
or UO_79 (O_79,N_14931,N_14906);
nand UO_80 (O_80,N_14973,N_14908);
and UO_81 (O_81,N_14958,N_14960);
nor UO_82 (O_82,N_14905,N_14900);
nand UO_83 (O_83,N_14935,N_14882);
nand UO_84 (O_84,N_14998,N_14876);
xnor UO_85 (O_85,N_14939,N_14998);
and UO_86 (O_86,N_14919,N_14987);
and UO_87 (O_87,N_14876,N_14982);
nand UO_88 (O_88,N_14983,N_14959);
or UO_89 (O_89,N_14889,N_14971);
nand UO_90 (O_90,N_14907,N_14992);
and UO_91 (O_91,N_14983,N_14987);
and UO_92 (O_92,N_14933,N_14911);
nor UO_93 (O_93,N_14922,N_14954);
or UO_94 (O_94,N_14910,N_14907);
nand UO_95 (O_95,N_14914,N_14956);
nand UO_96 (O_96,N_14973,N_14983);
and UO_97 (O_97,N_14926,N_14892);
nand UO_98 (O_98,N_14914,N_14946);
and UO_99 (O_99,N_14953,N_14888);
and UO_100 (O_100,N_14919,N_14962);
nand UO_101 (O_101,N_14961,N_14938);
and UO_102 (O_102,N_14884,N_14985);
or UO_103 (O_103,N_14973,N_14876);
or UO_104 (O_104,N_14911,N_14998);
and UO_105 (O_105,N_14950,N_14919);
nand UO_106 (O_106,N_14909,N_14900);
and UO_107 (O_107,N_14939,N_14991);
or UO_108 (O_108,N_14876,N_14927);
nor UO_109 (O_109,N_14981,N_14929);
or UO_110 (O_110,N_14899,N_14944);
xnor UO_111 (O_111,N_14922,N_14997);
or UO_112 (O_112,N_14889,N_14887);
and UO_113 (O_113,N_14966,N_14999);
xor UO_114 (O_114,N_14924,N_14914);
and UO_115 (O_115,N_14963,N_14908);
xnor UO_116 (O_116,N_14904,N_14883);
and UO_117 (O_117,N_14941,N_14920);
and UO_118 (O_118,N_14960,N_14955);
nor UO_119 (O_119,N_14880,N_14917);
nand UO_120 (O_120,N_14904,N_14961);
xor UO_121 (O_121,N_14997,N_14891);
and UO_122 (O_122,N_14915,N_14935);
xor UO_123 (O_123,N_14939,N_14964);
nor UO_124 (O_124,N_14941,N_14985);
or UO_125 (O_125,N_14988,N_14922);
nand UO_126 (O_126,N_14906,N_14981);
or UO_127 (O_127,N_14983,N_14942);
nand UO_128 (O_128,N_14938,N_14915);
and UO_129 (O_129,N_14898,N_14884);
xnor UO_130 (O_130,N_14929,N_14998);
or UO_131 (O_131,N_14908,N_14899);
and UO_132 (O_132,N_14942,N_14890);
and UO_133 (O_133,N_14962,N_14947);
nor UO_134 (O_134,N_14953,N_14965);
nand UO_135 (O_135,N_14897,N_14902);
nor UO_136 (O_136,N_14879,N_14968);
nand UO_137 (O_137,N_14876,N_14937);
nand UO_138 (O_138,N_14929,N_14928);
nor UO_139 (O_139,N_14879,N_14993);
nand UO_140 (O_140,N_14986,N_14979);
nand UO_141 (O_141,N_14953,N_14898);
nor UO_142 (O_142,N_14988,N_14921);
nor UO_143 (O_143,N_14994,N_14979);
nand UO_144 (O_144,N_14909,N_14913);
nand UO_145 (O_145,N_14979,N_14960);
and UO_146 (O_146,N_14876,N_14978);
nor UO_147 (O_147,N_14911,N_14956);
nor UO_148 (O_148,N_14903,N_14957);
xnor UO_149 (O_149,N_14979,N_14947);
nand UO_150 (O_150,N_14893,N_14911);
xnor UO_151 (O_151,N_14962,N_14883);
nor UO_152 (O_152,N_14938,N_14923);
nand UO_153 (O_153,N_14943,N_14900);
or UO_154 (O_154,N_14961,N_14923);
nand UO_155 (O_155,N_14899,N_14937);
nand UO_156 (O_156,N_14881,N_14951);
or UO_157 (O_157,N_14943,N_14890);
nand UO_158 (O_158,N_14878,N_14992);
xor UO_159 (O_159,N_14992,N_14973);
or UO_160 (O_160,N_14888,N_14890);
nor UO_161 (O_161,N_14878,N_14888);
xnor UO_162 (O_162,N_14897,N_14992);
or UO_163 (O_163,N_14879,N_14877);
nand UO_164 (O_164,N_14931,N_14973);
or UO_165 (O_165,N_14881,N_14981);
or UO_166 (O_166,N_14903,N_14938);
nand UO_167 (O_167,N_14942,N_14911);
nand UO_168 (O_168,N_14876,N_14895);
xor UO_169 (O_169,N_14913,N_14914);
nor UO_170 (O_170,N_14884,N_14977);
or UO_171 (O_171,N_14978,N_14900);
or UO_172 (O_172,N_14939,N_14883);
nor UO_173 (O_173,N_14920,N_14898);
and UO_174 (O_174,N_14904,N_14896);
xnor UO_175 (O_175,N_14998,N_14916);
and UO_176 (O_176,N_14996,N_14957);
nand UO_177 (O_177,N_14944,N_14968);
nor UO_178 (O_178,N_14978,N_14985);
nor UO_179 (O_179,N_14927,N_14998);
and UO_180 (O_180,N_14956,N_14943);
nand UO_181 (O_181,N_14894,N_14985);
nor UO_182 (O_182,N_14885,N_14982);
nand UO_183 (O_183,N_14946,N_14913);
nand UO_184 (O_184,N_14949,N_14914);
nand UO_185 (O_185,N_14951,N_14962);
xnor UO_186 (O_186,N_14912,N_14948);
and UO_187 (O_187,N_14974,N_14902);
or UO_188 (O_188,N_14989,N_14937);
or UO_189 (O_189,N_14904,N_14999);
xor UO_190 (O_190,N_14887,N_14997);
nor UO_191 (O_191,N_14913,N_14926);
or UO_192 (O_192,N_14894,N_14980);
nand UO_193 (O_193,N_14995,N_14875);
or UO_194 (O_194,N_14883,N_14919);
or UO_195 (O_195,N_14885,N_14883);
or UO_196 (O_196,N_14974,N_14979);
nand UO_197 (O_197,N_14906,N_14946);
nor UO_198 (O_198,N_14936,N_14901);
nor UO_199 (O_199,N_14928,N_14980);
and UO_200 (O_200,N_14973,N_14922);
nor UO_201 (O_201,N_14942,N_14943);
or UO_202 (O_202,N_14949,N_14912);
nor UO_203 (O_203,N_14959,N_14996);
nand UO_204 (O_204,N_14950,N_14999);
and UO_205 (O_205,N_14957,N_14889);
nor UO_206 (O_206,N_14875,N_14893);
and UO_207 (O_207,N_14933,N_14980);
nor UO_208 (O_208,N_14902,N_14951);
and UO_209 (O_209,N_14920,N_14970);
nand UO_210 (O_210,N_14894,N_14909);
and UO_211 (O_211,N_14951,N_14917);
and UO_212 (O_212,N_14934,N_14901);
and UO_213 (O_213,N_14935,N_14939);
xor UO_214 (O_214,N_14945,N_14920);
nand UO_215 (O_215,N_14968,N_14939);
nand UO_216 (O_216,N_14906,N_14939);
and UO_217 (O_217,N_14978,N_14933);
or UO_218 (O_218,N_14948,N_14937);
nor UO_219 (O_219,N_14983,N_14941);
or UO_220 (O_220,N_14927,N_14920);
nor UO_221 (O_221,N_14879,N_14978);
xor UO_222 (O_222,N_14898,N_14998);
or UO_223 (O_223,N_14952,N_14906);
xnor UO_224 (O_224,N_14895,N_14978);
xor UO_225 (O_225,N_14969,N_14912);
xnor UO_226 (O_226,N_14883,N_14944);
xor UO_227 (O_227,N_14916,N_14939);
or UO_228 (O_228,N_14882,N_14943);
or UO_229 (O_229,N_14960,N_14998);
xor UO_230 (O_230,N_14878,N_14887);
nand UO_231 (O_231,N_14955,N_14888);
xor UO_232 (O_232,N_14928,N_14887);
and UO_233 (O_233,N_14914,N_14888);
xnor UO_234 (O_234,N_14931,N_14878);
xnor UO_235 (O_235,N_14891,N_14915);
or UO_236 (O_236,N_14895,N_14915);
nor UO_237 (O_237,N_14884,N_14948);
nor UO_238 (O_238,N_14994,N_14913);
nand UO_239 (O_239,N_14935,N_14937);
xnor UO_240 (O_240,N_14987,N_14896);
xnor UO_241 (O_241,N_14931,N_14893);
or UO_242 (O_242,N_14948,N_14935);
or UO_243 (O_243,N_14892,N_14883);
or UO_244 (O_244,N_14992,N_14940);
xor UO_245 (O_245,N_14893,N_14942);
or UO_246 (O_246,N_14888,N_14892);
and UO_247 (O_247,N_14993,N_14883);
and UO_248 (O_248,N_14879,N_14935);
nor UO_249 (O_249,N_14960,N_14963);
and UO_250 (O_250,N_14985,N_14937);
nand UO_251 (O_251,N_14967,N_14943);
or UO_252 (O_252,N_14963,N_14888);
xor UO_253 (O_253,N_14906,N_14924);
nor UO_254 (O_254,N_14950,N_14993);
nor UO_255 (O_255,N_14982,N_14920);
nand UO_256 (O_256,N_14909,N_14885);
xor UO_257 (O_257,N_14990,N_14970);
xnor UO_258 (O_258,N_14939,N_14977);
nand UO_259 (O_259,N_14906,N_14878);
and UO_260 (O_260,N_14925,N_14959);
nand UO_261 (O_261,N_14969,N_14909);
xnor UO_262 (O_262,N_14894,N_14939);
xor UO_263 (O_263,N_14895,N_14922);
xnor UO_264 (O_264,N_14985,N_14990);
nor UO_265 (O_265,N_14927,N_14986);
nor UO_266 (O_266,N_14989,N_14985);
nand UO_267 (O_267,N_14973,N_14950);
nor UO_268 (O_268,N_14953,N_14940);
nor UO_269 (O_269,N_14895,N_14883);
and UO_270 (O_270,N_14975,N_14991);
and UO_271 (O_271,N_14903,N_14920);
nor UO_272 (O_272,N_14917,N_14879);
xnor UO_273 (O_273,N_14952,N_14989);
xnor UO_274 (O_274,N_14908,N_14877);
xnor UO_275 (O_275,N_14982,N_14979);
nand UO_276 (O_276,N_14953,N_14993);
or UO_277 (O_277,N_14995,N_14958);
xnor UO_278 (O_278,N_14883,N_14913);
or UO_279 (O_279,N_14991,N_14897);
and UO_280 (O_280,N_14960,N_14882);
nor UO_281 (O_281,N_14986,N_14967);
nand UO_282 (O_282,N_14914,N_14926);
or UO_283 (O_283,N_14915,N_14961);
or UO_284 (O_284,N_14945,N_14953);
or UO_285 (O_285,N_14880,N_14995);
or UO_286 (O_286,N_14876,N_14940);
nand UO_287 (O_287,N_14931,N_14919);
and UO_288 (O_288,N_14999,N_14963);
or UO_289 (O_289,N_14898,N_14990);
nor UO_290 (O_290,N_14966,N_14895);
or UO_291 (O_291,N_14952,N_14899);
nor UO_292 (O_292,N_14954,N_14975);
or UO_293 (O_293,N_14948,N_14883);
and UO_294 (O_294,N_14876,N_14886);
xnor UO_295 (O_295,N_14879,N_14912);
nand UO_296 (O_296,N_14949,N_14977);
xnor UO_297 (O_297,N_14974,N_14997);
and UO_298 (O_298,N_14876,N_14904);
nor UO_299 (O_299,N_14886,N_14940);
nor UO_300 (O_300,N_14976,N_14903);
or UO_301 (O_301,N_14883,N_14933);
and UO_302 (O_302,N_14973,N_14929);
or UO_303 (O_303,N_14989,N_14913);
or UO_304 (O_304,N_14918,N_14887);
xnor UO_305 (O_305,N_14882,N_14924);
xnor UO_306 (O_306,N_14967,N_14915);
and UO_307 (O_307,N_14890,N_14909);
nor UO_308 (O_308,N_14876,N_14875);
xor UO_309 (O_309,N_14882,N_14900);
xor UO_310 (O_310,N_14946,N_14922);
and UO_311 (O_311,N_14935,N_14914);
nand UO_312 (O_312,N_14915,N_14920);
xnor UO_313 (O_313,N_14994,N_14933);
nand UO_314 (O_314,N_14877,N_14878);
nand UO_315 (O_315,N_14941,N_14962);
and UO_316 (O_316,N_14981,N_14913);
xor UO_317 (O_317,N_14918,N_14910);
nand UO_318 (O_318,N_14974,N_14939);
and UO_319 (O_319,N_14996,N_14984);
or UO_320 (O_320,N_14998,N_14955);
or UO_321 (O_321,N_14976,N_14888);
or UO_322 (O_322,N_14999,N_14967);
nor UO_323 (O_323,N_14962,N_14902);
and UO_324 (O_324,N_14891,N_14935);
nor UO_325 (O_325,N_14910,N_14998);
xnor UO_326 (O_326,N_14977,N_14901);
nor UO_327 (O_327,N_14936,N_14880);
nor UO_328 (O_328,N_14878,N_14934);
or UO_329 (O_329,N_14942,N_14898);
xnor UO_330 (O_330,N_14917,N_14875);
xor UO_331 (O_331,N_14978,N_14890);
nor UO_332 (O_332,N_14883,N_14877);
and UO_333 (O_333,N_14887,N_14992);
xor UO_334 (O_334,N_14876,N_14905);
nor UO_335 (O_335,N_14902,N_14885);
nor UO_336 (O_336,N_14948,N_14879);
or UO_337 (O_337,N_14913,N_14904);
nor UO_338 (O_338,N_14979,N_14944);
and UO_339 (O_339,N_14974,N_14991);
and UO_340 (O_340,N_14898,N_14976);
nand UO_341 (O_341,N_14911,N_14926);
xor UO_342 (O_342,N_14951,N_14910);
nand UO_343 (O_343,N_14952,N_14883);
and UO_344 (O_344,N_14940,N_14946);
nand UO_345 (O_345,N_14918,N_14971);
and UO_346 (O_346,N_14959,N_14888);
nand UO_347 (O_347,N_14958,N_14878);
nor UO_348 (O_348,N_14885,N_14907);
nor UO_349 (O_349,N_14876,N_14999);
and UO_350 (O_350,N_14972,N_14984);
xnor UO_351 (O_351,N_14918,N_14880);
or UO_352 (O_352,N_14926,N_14928);
xor UO_353 (O_353,N_14879,N_14950);
nand UO_354 (O_354,N_14992,N_14875);
and UO_355 (O_355,N_14998,N_14976);
nor UO_356 (O_356,N_14952,N_14950);
nand UO_357 (O_357,N_14988,N_14981);
xnor UO_358 (O_358,N_14956,N_14912);
and UO_359 (O_359,N_14994,N_14991);
or UO_360 (O_360,N_14895,N_14952);
and UO_361 (O_361,N_14966,N_14933);
nand UO_362 (O_362,N_14908,N_14940);
xor UO_363 (O_363,N_14954,N_14974);
nor UO_364 (O_364,N_14997,N_14885);
or UO_365 (O_365,N_14899,N_14991);
and UO_366 (O_366,N_14986,N_14947);
nand UO_367 (O_367,N_14983,N_14995);
nor UO_368 (O_368,N_14967,N_14954);
nor UO_369 (O_369,N_14948,N_14886);
nand UO_370 (O_370,N_14969,N_14950);
xor UO_371 (O_371,N_14995,N_14899);
and UO_372 (O_372,N_14891,N_14917);
xnor UO_373 (O_373,N_14914,N_14970);
xor UO_374 (O_374,N_14881,N_14885);
or UO_375 (O_375,N_14983,N_14965);
nor UO_376 (O_376,N_14949,N_14880);
nand UO_377 (O_377,N_14910,N_14906);
nand UO_378 (O_378,N_14973,N_14911);
xnor UO_379 (O_379,N_14911,N_14997);
nor UO_380 (O_380,N_14928,N_14906);
or UO_381 (O_381,N_14930,N_14903);
nand UO_382 (O_382,N_14987,N_14922);
and UO_383 (O_383,N_14919,N_14921);
nand UO_384 (O_384,N_14930,N_14934);
and UO_385 (O_385,N_14994,N_14894);
nor UO_386 (O_386,N_14997,N_14926);
nand UO_387 (O_387,N_14907,N_14941);
nand UO_388 (O_388,N_14917,N_14979);
and UO_389 (O_389,N_14930,N_14932);
xnor UO_390 (O_390,N_14988,N_14877);
and UO_391 (O_391,N_14877,N_14944);
xnor UO_392 (O_392,N_14975,N_14891);
xor UO_393 (O_393,N_14982,N_14953);
xor UO_394 (O_394,N_14943,N_14928);
and UO_395 (O_395,N_14884,N_14999);
and UO_396 (O_396,N_14906,N_14923);
xor UO_397 (O_397,N_14976,N_14987);
xor UO_398 (O_398,N_14932,N_14985);
or UO_399 (O_399,N_14893,N_14948);
xnor UO_400 (O_400,N_14889,N_14882);
nor UO_401 (O_401,N_14920,N_14889);
or UO_402 (O_402,N_14898,N_14971);
nand UO_403 (O_403,N_14978,N_14980);
xor UO_404 (O_404,N_14896,N_14927);
or UO_405 (O_405,N_14996,N_14905);
or UO_406 (O_406,N_14950,N_14923);
nor UO_407 (O_407,N_14911,N_14943);
nor UO_408 (O_408,N_14960,N_14981);
nand UO_409 (O_409,N_14884,N_14993);
and UO_410 (O_410,N_14995,N_14968);
and UO_411 (O_411,N_14940,N_14973);
or UO_412 (O_412,N_14995,N_14966);
and UO_413 (O_413,N_14883,N_14886);
nor UO_414 (O_414,N_14957,N_14905);
nand UO_415 (O_415,N_14910,N_14923);
or UO_416 (O_416,N_14929,N_14984);
xor UO_417 (O_417,N_14924,N_14892);
or UO_418 (O_418,N_14913,N_14877);
or UO_419 (O_419,N_14934,N_14915);
nor UO_420 (O_420,N_14996,N_14958);
nand UO_421 (O_421,N_14954,N_14976);
and UO_422 (O_422,N_14906,N_14938);
nand UO_423 (O_423,N_14894,N_14920);
and UO_424 (O_424,N_14945,N_14895);
and UO_425 (O_425,N_14894,N_14885);
nand UO_426 (O_426,N_14987,N_14979);
and UO_427 (O_427,N_14899,N_14986);
or UO_428 (O_428,N_14941,N_14967);
or UO_429 (O_429,N_14911,N_14892);
xor UO_430 (O_430,N_14971,N_14995);
nand UO_431 (O_431,N_14901,N_14963);
or UO_432 (O_432,N_14997,N_14912);
xnor UO_433 (O_433,N_14877,N_14971);
nand UO_434 (O_434,N_14883,N_14956);
or UO_435 (O_435,N_14926,N_14934);
or UO_436 (O_436,N_14963,N_14983);
and UO_437 (O_437,N_14975,N_14882);
or UO_438 (O_438,N_14886,N_14916);
or UO_439 (O_439,N_14899,N_14975);
nor UO_440 (O_440,N_14925,N_14953);
nand UO_441 (O_441,N_14985,N_14902);
nand UO_442 (O_442,N_14964,N_14996);
nand UO_443 (O_443,N_14921,N_14900);
xor UO_444 (O_444,N_14972,N_14959);
nand UO_445 (O_445,N_14918,N_14972);
or UO_446 (O_446,N_14954,N_14935);
xnor UO_447 (O_447,N_14914,N_14991);
and UO_448 (O_448,N_14914,N_14904);
and UO_449 (O_449,N_14882,N_14951);
nor UO_450 (O_450,N_14936,N_14906);
and UO_451 (O_451,N_14956,N_14959);
nand UO_452 (O_452,N_14951,N_14894);
nand UO_453 (O_453,N_14879,N_14982);
or UO_454 (O_454,N_14892,N_14938);
and UO_455 (O_455,N_14903,N_14978);
nand UO_456 (O_456,N_14902,N_14924);
or UO_457 (O_457,N_14977,N_14889);
nor UO_458 (O_458,N_14961,N_14887);
nor UO_459 (O_459,N_14925,N_14913);
or UO_460 (O_460,N_14960,N_14903);
nor UO_461 (O_461,N_14926,N_14875);
nor UO_462 (O_462,N_14984,N_14952);
nand UO_463 (O_463,N_14917,N_14923);
nor UO_464 (O_464,N_14876,N_14950);
or UO_465 (O_465,N_14987,N_14994);
nand UO_466 (O_466,N_14959,N_14884);
and UO_467 (O_467,N_14966,N_14936);
and UO_468 (O_468,N_14959,N_14921);
xnor UO_469 (O_469,N_14887,N_14901);
xnor UO_470 (O_470,N_14939,N_14971);
nand UO_471 (O_471,N_14936,N_14917);
xnor UO_472 (O_472,N_14876,N_14883);
nor UO_473 (O_473,N_14975,N_14939);
xnor UO_474 (O_474,N_14986,N_14961);
xor UO_475 (O_475,N_14902,N_14893);
or UO_476 (O_476,N_14923,N_14998);
nor UO_477 (O_477,N_14927,N_14936);
nor UO_478 (O_478,N_14996,N_14920);
nor UO_479 (O_479,N_14968,N_14949);
nand UO_480 (O_480,N_14923,N_14972);
xnor UO_481 (O_481,N_14948,N_14905);
xnor UO_482 (O_482,N_14952,N_14919);
nor UO_483 (O_483,N_14903,N_14906);
nor UO_484 (O_484,N_14955,N_14958);
or UO_485 (O_485,N_14885,N_14915);
and UO_486 (O_486,N_14918,N_14900);
and UO_487 (O_487,N_14992,N_14891);
nand UO_488 (O_488,N_14888,N_14937);
xnor UO_489 (O_489,N_14924,N_14893);
nor UO_490 (O_490,N_14922,N_14892);
and UO_491 (O_491,N_14915,N_14933);
nand UO_492 (O_492,N_14898,N_14890);
and UO_493 (O_493,N_14997,N_14935);
xnor UO_494 (O_494,N_14983,N_14916);
or UO_495 (O_495,N_14907,N_14917);
nand UO_496 (O_496,N_14902,N_14892);
and UO_497 (O_497,N_14893,N_14935);
nand UO_498 (O_498,N_14933,N_14990);
or UO_499 (O_499,N_14924,N_14897);
or UO_500 (O_500,N_14944,N_14935);
nor UO_501 (O_501,N_14945,N_14938);
xor UO_502 (O_502,N_14938,N_14881);
xnor UO_503 (O_503,N_14985,N_14996);
or UO_504 (O_504,N_14939,N_14920);
xor UO_505 (O_505,N_14942,N_14912);
and UO_506 (O_506,N_14965,N_14941);
or UO_507 (O_507,N_14977,N_14903);
nor UO_508 (O_508,N_14898,N_14916);
nor UO_509 (O_509,N_14949,N_14924);
xor UO_510 (O_510,N_14878,N_14950);
nor UO_511 (O_511,N_14953,N_14978);
nor UO_512 (O_512,N_14958,N_14988);
and UO_513 (O_513,N_14953,N_14948);
nand UO_514 (O_514,N_14959,N_14964);
nand UO_515 (O_515,N_14957,N_14911);
nand UO_516 (O_516,N_14982,N_14969);
and UO_517 (O_517,N_14992,N_14933);
xor UO_518 (O_518,N_14924,N_14999);
or UO_519 (O_519,N_14887,N_14933);
or UO_520 (O_520,N_14973,N_14928);
xor UO_521 (O_521,N_14981,N_14978);
and UO_522 (O_522,N_14977,N_14928);
nor UO_523 (O_523,N_14927,N_14989);
nand UO_524 (O_524,N_14887,N_14989);
nand UO_525 (O_525,N_14991,N_14907);
nand UO_526 (O_526,N_14915,N_14890);
xnor UO_527 (O_527,N_14886,N_14878);
or UO_528 (O_528,N_14957,N_14907);
nand UO_529 (O_529,N_14966,N_14875);
and UO_530 (O_530,N_14895,N_14974);
nand UO_531 (O_531,N_14947,N_14937);
xor UO_532 (O_532,N_14909,N_14881);
nand UO_533 (O_533,N_14960,N_14948);
and UO_534 (O_534,N_14886,N_14978);
nor UO_535 (O_535,N_14958,N_14990);
and UO_536 (O_536,N_14878,N_14996);
nand UO_537 (O_537,N_14990,N_14955);
nor UO_538 (O_538,N_14928,N_14878);
or UO_539 (O_539,N_14917,N_14953);
nor UO_540 (O_540,N_14961,N_14990);
or UO_541 (O_541,N_14966,N_14952);
nand UO_542 (O_542,N_14966,N_14892);
or UO_543 (O_543,N_14925,N_14997);
xnor UO_544 (O_544,N_14956,N_14881);
nor UO_545 (O_545,N_14910,N_14898);
nor UO_546 (O_546,N_14933,N_14885);
or UO_547 (O_547,N_14990,N_14879);
nor UO_548 (O_548,N_14971,N_14981);
nand UO_549 (O_549,N_14900,N_14965);
or UO_550 (O_550,N_14957,N_14902);
xor UO_551 (O_551,N_14917,N_14904);
xnor UO_552 (O_552,N_14906,N_14943);
nand UO_553 (O_553,N_14884,N_14957);
nor UO_554 (O_554,N_14879,N_14972);
nor UO_555 (O_555,N_14929,N_14941);
xor UO_556 (O_556,N_14931,N_14974);
or UO_557 (O_557,N_14876,N_14932);
and UO_558 (O_558,N_14911,N_14963);
nor UO_559 (O_559,N_14906,N_14940);
and UO_560 (O_560,N_14935,N_14919);
xor UO_561 (O_561,N_14997,N_14879);
nand UO_562 (O_562,N_14947,N_14950);
xor UO_563 (O_563,N_14922,N_14962);
xnor UO_564 (O_564,N_14983,N_14954);
nor UO_565 (O_565,N_14891,N_14952);
and UO_566 (O_566,N_14952,N_14996);
nand UO_567 (O_567,N_14977,N_14879);
and UO_568 (O_568,N_14973,N_14901);
xor UO_569 (O_569,N_14928,N_14879);
xnor UO_570 (O_570,N_14956,N_14880);
xor UO_571 (O_571,N_14925,N_14940);
nor UO_572 (O_572,N_14888,N_14991);
and UO_573 (O_573,N_14925,N_14919);
or UO_574 (O_574,N_14885,N_14953);
and UO_575 (O_575,N_14989,N_14955);
or UO_576 (O_576,N_14948,N_14990);
or UO_577 (O_577,N_14885,N_14914);
nor UO_578 (O_578,N_14875,N_14878);
nand UO_579 (O_579,N_14948,N_14890);
and UO_580 (O_580,N_14963,N_14958);
nor UO_581 (O_581,N_14927,N_14934);
and UO_582 (O_582,N_14895,N_14918);
nand UO_583 (O_583,N_14973,N_14889);
nand UO_584 (O_584,N_14893,N_14884);
nor UO_585 (O_585,N_14932,N_14934);
and UO_586 (O_586,N_14945,N_14878);
xnor UO_587 (O_587,N_14929,N_14937);
and UO_588 (O_588,N_14950,N_14911);
or UO_589 (O_589,N_14993,N_14934);
and UO_590 (O_590,N_14940,N_14963);
nand UO_591 (O_591,N_14909,N_14928);
or UO_592 (O_592,N_14978,N_14971);
nand UO_593 (O_593,N_14934,N_14893);
or UO_594 (O_594,N_14990,N_14957);
or UO_595 (O_595,N_14882,N_14916);
nor UO_596 (O_596,N_14909,N_14896);
nor UO_597 (O_597,N_14986,N_14925);
nand UO_598 (O_598,N_14970,N_14989);
or UO_599 (O_599,N_14881,N_14949);
and UO_600 (O_600,N_14948,N_14945);
nand UO_601 (O_601,N_14894,N_14962);
xnor UO_602 (O_602,N_14997,N_14953);
and UO_603 (O_603,N_14954,N_14962);
nand UO_604 (O_604,N_14881,N_14898);
or UO_605 (O_605,N_14993,N_14992);
nor UO_606 (O_606,N_14971,N_14954);
xor UO_607 (O_607,N_14929,N_14968);
and UO_608 (O_608,N_14924,N_14890);
and UO_609 (O_609,N_14957,N_14963);
nand UO_610 (O_610,N_14956,N_14935);
nor UO_611 (O_611,N_14974,N_14919);
nor UO_612 (O_612,N_14886,N_14938);
xnor UO_613 (O_613,N_14988,N_14937);
nand UO_614 (O_614,N_14961,N_14929);
nor UO_615 (O_615,N_14979,N_14984);
nor UO_616 (O_616,N_14973,N_14894);
and UO_617 (O_617,N_14989,N_14923);
nor UO_618 (O_618,N_14937,N_14960);
and UO_619 (O_619,N_14971,N_14941);
nand UO_620 (O_620,N_14897,N_14898);
nor UO_621 (O_621,N_14905,N_14992);
and UO_622 (O_622,N_14952,N_14979);
nand UO_623 (O_623,N_14927,N_14951);
nor UO_624 (O_624,N_14971,N_14993);
nor UO_625 (O_625,N_14962,N_14999);
or UO_626 (O_626,N_14875,N_14956);
nor UO_627 (O_627,N_14976,N_14946);
xnor UO_628 (O_628,N_14921,N_14980);
nor UO_629 (O_629,N_14895,N_14887);
nand UO_630 (O_630,N_14913,N_14950);
and UO_631 (O_631,N_14890,N_14913);
xor UO_632 (O_632,N_14993,N_14931);
nand UO_633 (O_633,N_14936,N_14960);
nor UO_634 (O_634,N_14935,N_14923);
nor UO_635 (O_635,N_14906,N_14882);
nand UO_636 (O_636,N_14901,N_14893);
nor UO_637 (O_637,N_14884,N_14918);
and UO_638 (O_638,N_14901,N_14953);
nor UO_639 (O_639,N_14942,N_14946);
xor UO_640 (O_640,N_14955,N_14903);
nor UO_641 (O_641,N_14933,N_14947);
nor UO_642 (O_642,N_14977,N_14952);
or UO_643 (O_643,N_14955,N_14985);
xor UO_644 (O_644,N_14991,N_14989);
or UO_645 (O_645,N_14920,N_14881);
nor UO_646 (O_646,N_14922,N_14975);
xnor UO_647 (O_647,N_14949,N_14963);
and UO_648 (O_648,N_14961,N_14941);
nand UO_649 (O_649,N_14915,N_14912);
or UO_650 (O_650,N_14993,N_14898);
and UO_651 (O_651,N_14904,N_14933);
xor UO_652 (O_652,N_14954,N_14900);
xor UO_653 (O_653,N_14942,N_14921);
nand UO_654 (O_654,N_14887,N_14919);
nor UO_655 (O_655,N_14940,N_14891);
nor UO_656 (O_656,N_14901,N_14947);
nand UO_657 (O_657,N_14976,N_14896);
or UO_658 (O_658,N_14892,N_14969);
nand UO_659 (O_659,N_14969,N_14890);
and UO_660 (O_660,N_14889,N_14903);
xor UO_661 (O_661,N_14902,N_14929);
or UO_662 (O_662,N_14998,N_14942);
or UO_663 (O_663,N_14916,N_14920);
nand UO_664 (O_664,N_14966,N_14920);
xnor UO_665 (O_665,N_14959,N_14999);
nor UO_666 (O_666,N_14983,N_14900);
or UO_667 (O_667,N_14930,N_14900);
and UO_668 (O_668,N_14983,N_14997);
or UO_669 (O_669,N_14958,N_14916);
and UO_670 (O_670,N_14971,N_14884);
and UO_671 (O_671,N_14963,N_14928);
nand UO_672 (O_672,N_14877,N_14986);
or UO_673 (O_673,N_14894,N_14946);
nor UO_674 (O_674,N_14936,N_14893);
nor UO_675 (O_675,N_14899,N_14900);
xor UO_676 (O_676,N_14877,N_14931);
or UO_677 (O_677,N_14964,N_14963);
and UO_678 (O_678,N_14924,N_14927);
or UO_679 (O_679,N_14929,N_14927);
or UO_680 (O_680,N_14875,N_14980);
xor UO_681 (O_681,N_14985,N_14929);
nor UO_682 (O_682,N_14882,N_14939);
or UO_683 (O_683,N_14941,N_14906);
xnor UO_684 (O_684,N_14949,N_14970);
nor UO_685 (O_685,N_14921,N_14994);
nor UO_686 (O_686,N_14943,N_14919);
nand UO_687 (O_687,N_14990,N_14944);
nor UO_688 (O_688,N_14896,N_14938);
or UO_689 (O_689,N_14887,N_14932);
and UO_690 (O_690,N_14973,N_14963);
nand UO_691 (O_691,N_14963,N_14935);
xnor UO_692 (O_692,N_14899,N_14954);
xor UO_693 (O_693,N_14962,N_14955);
nand UO_694 (O_694,N_14922,N_14912);
and UO_695 (O_695,N_14979,N_14972);
or UO_696 (O_696,N_14891,N_14947);
nor UO_697 (O_697,N_14908,N_14991);
xor UO_698 (O_698,N_14961,N_14908);
xnor UO_699 (O_699,N_14945,N_14934);
xnor UO_700 (O_700,N_14997,N_14936);
or UO_701 (O_701,N_14969,N_14988);
xor UO_702 (O_702,N_14952,N_14962);
nor UO_703 (O_703,N_14946,N_14943);
nor UO_704 (O_704,N_14917,N_14925);
or UO_705 (O_705,N_14876,N_14987);
or UO_706 (O_706,N_14880,N_14883);
and UO_707 (O_707,N_14990,N_14924);
or UO_708 (O_708,N_14931,N_14880);
nand UO_709 (O_709,N_14882,N_14953);
and UO_710 (O_710,N_14892,N_14972);
nor UO_711 (O_711,N_14889,N_14906);
and UO_712 (O_712,N_14909,N_14983);
nand UO_713 (O_713,N_14935,N_14992);
or UO_714 (O_714,N_14922,N_14908);
nor UO_715 (O_715,N_14876,N_14912);
and UO_716 (O_716,N_14997,N_14960);
nor UO_717 (O_717,N_14877,N_14891);
xnor UO_718 (O_718,N_14914,N_14978);
nand UO_719 (O_719,N_14975,N_14947);
or UO_720 (O_720,N_14910,N_14997);
nand UO_721 (O_721,N_14962,N_14892);
or UO_722 (O_722,N_14921,N_14967);
or UO_723 (O_723,N_14892,N_14982);
nand UO_724 (O_724,N_14998,N_14964);
nor UO_725 (O_725,N_14968,N_14931);
nor UO_726 (O_726,N_14875,N_14976);
or UO_727 (O_727,N_14976,N_14999);
and UO_728 (O_728,N_14944,N_14896);
and UO_729 (O_729,N_14962,N_14905);
nor UO_730 (O_730,N_14992,N_14925);
nand UO_731 (O_731,N_14896,N_14929);
and UO_732 (O_732,N_14958,N_14942);
xnor UO_733 (O_733,N_14968,N_14926);
xor UO_734 (O_734,N_14973,N_14954);
xnor UO_735 (O_735,N_14883,N_14997);
and UO_736 (O_736,N_14944,N_14960);
nor UO_737 (O_737,N_14962,N_14968);
nor UO_738 (O_738,N_14878,N_14968);
nand UO_739 (O_739,N_14908,N_14915);
or UO_740 (O_740,N_14896,N_14875);
nor UO_741 (O_741,N_14914,N_14975);
nand UO_742 (O_742,N_14955,N_14881);
nand UO_743 (O_743,N_14930,N_14928);
xnor UO_744 (O_744,N_14879,N_14971);
nand UO_745 (O_745,N_14951,N_14979);
or UO_746 (O_746,N_14930,N_14933);
or UO_747 (O_747,N_14906,N_14902);
nor UO_748 (O_748,N_14905,N_14925);
or UO_749 (O_749,N_14959,N_14876);
and UO_750 (O_750,N_14936,N_14968);
and UO_751 (O_751,N_14882,N_14998);
xnor UO_752 (O_752,N_14902,N_14963);
xor UO_753 (O_753,N_14965,N_14906);
nand UO_754 (O_754,N_14993,N_14925);
and UO_755 (O_755,N_14897,N_14970);
xor UO_756 (O_756,N_14903,N_14975);
nand UO_757 (O_757,N_14903,N_14998);
xnor UO_758 (O_758,N_14972,N_14917);
nand UO_759 (O_759,N_14889,N_14895);
or UO_760 (O_760,N_14944,N_14901);
nor UO_761 (O_761,N_14901,N_14917);
nor UO_762 (O_762,N_14950,N_14988);
nand UO_763 (O_763,N_14979,N_14976);
and UO_764 (O_764,N_14881,N_14941);
nor UO_765 (O_765,N_14938,N_14900);
and UO_766 (O_766,N_14910,N_14891);
and UO_767 (O_767,N_14946,N_14947);
and UO_768 (O_768,N_14950,N_14967);
or UO_769 (O_769,N_14946,N_14877);
or UO_770 (O_770,N_14946,N_14983);
nor UO_771 (O_771,N_14931,N_14884);
xor UO_772 (O_772,N_14968,N_14915);
or UO_773 (O_773,N_14911,N_14909);
and UO_774 (O_774,N_14877,N_14962);
or UO_775 (O_775,N_14944,N_14937);
or UO_776 (O_776,N_14974,N_14896);
nor UO_777 (O_777,N_14897,N_14876);
nand UO_778 (O_778,N_14911,N_14962);
nor UO_779 (O_779,N_14909,N_14960);
or UO_780 (O_780,N_14984,N_14890);
nor UO_781 (O_781,N_14938,N_14976);
or UO_782 (O_782,N_14963,N_14913);
nor UO_783 (O_783,N_14922,N_14925);
nor UO_784 (O_784,N_14911,N_14904);
and UO_785 (O_785,N_14949,N_14994);
nor UO_786 (O_786,N_14954,N_14982);
and UO_787 (O_787,N_14963,N_14922);
and UO_788 (O_788,N_14975,N_14927);
nand UO_789 (O_789,N_14958,N_14938);
and UO_790 (O_790,N_14937,N_14886);
or UO_791 (O_791,N_14962,N_14939);
nand UO_792 (O_792,N_14910,N_14934);
or UO_793 (O_793,N_14946,N_14984);
and UO_794 (O_794,N_14895,N_14976);
nor UO_795 (O_795,N_14881,N_14917);
nand UO_796 (O_796,N_14949,N_14916);
xnor UO_797 (O_797,N_14933,N_14891);
nor UO_798 (O_798,N_14916,N_14966);
and UO_799 (O_799,N_14952,N_14980);
nand UO_800 (O_800,N_14889,N_14910);
nand UO_801 (O_801,N_14972,N_14961);
nand UO_802 (O_802,N_14977,N_14902);
or UO_803 (O_803,N_14885,N_14928);
xor UO_804 (O_804,N_14955,N_14929);
nor UO_805 (O_805,N_14881,N_14912);
nand UO_806 (O_806,N_14924,N_14895);
or UO_807 (O_807,N_14944,N_14904);
or UO_808 (O_808,N_14918,N_14877);
or UO_809 (O_809,N_14975,N_14920);
xnor UO_810 (O_810,N_14990,N_14881);
and UO_811 (O_811,N_14927,N_14993);
xor UO_812 (O_812,N_14955,N_14891);
or UO_813 (O_813,N_14943,N_14995);
xor UO_814 (O_814,N_14996,N_14927);
xnor UO_815 (O_815,N_14924,N_14913);
xor UO_816 (O_816,N_14950,N_14907);
xnor UO_817 (O_817,N_14913,N_14999);
xnor UO_818 (O_818,N_14966,N_14977);
nor UO_819 (O_819,N_14956,N_14896);
nor UO_820 (O_820,N_14958,N_14945);
nor UO_821 (O_821,N_14887,N_14898);
nand UO_822 (O_822,N_14893,N_14890);
and UO_823 (O_823,N_14883,N_14914);
or UO_824 (O_824,N_14881,N_14907);
nor UO_825 (O_825,N_14953,N_14979);
or UO_826 (O_826,N_14980,N_14972);
nor UO_827 (O_827,N_14877,N_14900);
xnor UO_828 (O_828,N_14961,N_14882);
nand UO_829 (O_829,N_14951,N_14997);
nand UO_830 (O_830,N_14924,N_14956);
nand UO_831 (O_831,N_14985,N_14882);
nand UO_832 (O_832,N_14988,N_14986);
nand UO_833 (O_833,N_14989,N_14954);
and UO_834 (O_834,N_14950,N_14957);
xor UO_835 (O_835,N_14902,N_14936);
or UO_836 (O_836,N_14991,N_14998);
nand UO_837 (O_837,N_14877,N_14875);
nand UO_838 (O_838,N_14907,N_14961);
and UO_839 (O_839,N_14918,N_14952);
or UO_840 (O_840,N_14989,N_14939);
nand UO_841 (O_841,N_14892,N_14979);
nor UO_842 (O_842,N_14908,N_14983);
nand UO_843 (O_843,N_14944,N_14947);
and UO_844 (O_844,N_14966,N_14899);
xor UO_845 (O_845,N_14942,N_14969);
nand UO_846 (O_846,N_14901,N_14966);
and UO_847 (O_847,N_14922,N_14889);
nand UO_848 (O_848,N_14929,N_14939);
nand UO_849 (O_849,N_14967,N_14906);
nor UO_850 (O_850,N_14946,N_14954);
nor UO_851 (O_851,N_14896,N_14877);
or UO_852 (O_852,N_14999,N_14939);
or UO_853 (O_853,N_14955,N_14922);
nand UO_854 (O_854,N_14942,N_14993);
nand UO_855 (O_855,N_14947,N_14964);
nor UO_856 (O_856,N_14876,N_14920);
nand UO_857 (O_857,N_14983,N_14907);
or UO_858 (O_858,N_14905,N_14933);
and UO_859 (O_859,N_14999,N_14961);
nand UO_860 (O_860,N_14939,N_14932);
nor UO_861 (O_861,N_14916,N_14994);
and UO_862 (O_862,N_14978,N_14918);
and UO_863 (O_863,N_14916,N_14908);
or UO_864 (O_864,N_14954,N_14961);
xnor UO_865 (O_865,N_14961,N_14965);
and UO_866 (O_866,N_14935,N_14922);
nand UO_867 (O_867,N_14975,N_14901);
or UO_868 (O_868,N_14897,N_14947);
nor UO_869 (O_869,N_14916,N_14885);
nand UO_870 (O_870,N_14893,N_14919);
xnor UO_871 (O_871,N_14918,N_14883);
nand UO_872 (O_872,N_14945,N_14949);
xor UO_873 (O_873,N_14997,N_14909);
xor UO_874 (O_874,N_14953,N_14988);
and UO_875 (O_875,N_14966,N_14968);
and UO_876 (O_876,N_14929,N_14875);
and UO_877 (O_877,N_14876,N_14988);
and UO_878 (O_878,N_14922,N_14926);
and UO_879 (O_879,N_14992,N_14932);
xor UO_880 (O_880,N_14953,N_14922);
or UO_881 (O_881,N_14939,N_14972);
nor UO_882 (O_882,N_14877,N_14903);
nor UO_883 (O_883,N_14992,N_14966);
and UO_884 (O_884,N_14992,N_14931);
nor UO_885 (O_885,N_14937,N_14911);
nand UO_886 (O_886,N_14968,N_14970);
xor UO_887 (O_887,N_14893,N_14894);
or UO_888 (O_888,N_14884,N_14877);
or UO_889 (O_889,N_14957,N_14968);
xnor UO_890 (O_890,N_14878,N_14963);
nand UO_891 (O_891,N_14894,N_14902);
xor UO_892 (O_892,N_14979,N_14886);
nand UO_893 (O_893,N_14988,N_14983);
nor UO_894 (O_894,N_14918,N_14908);
nor UO_895 (O_895,N_14935,N_14961);
nor UO_896 (O_896,N_14991,N_14924);
xor UO_897 (O_897,N_14974,N_14925);
or UO_898 (O_898,N_14979,N_14896);
or UO_899 (O_899,N_14984,N_14922);
nand UO_900 (O_900,N_14943,N_14904);
and UO_901 (O_901,N_14952,N_14999);
nand UO_902 (O_902,N_14995,N_14934);
nand UO_903 (O_903,N_14953,N_14875);
nand UO_904 (O_904,N_14976,N_14919);
and UO_905 (O_905,N_14909,N_14908);
and UO_906 (O_906,N_14931,N_14981);
and UO_907 (O_907,N_14995,N_14987);
nor UO_908 (O_908,N_14975,N_14883);
nand UO_909 (O_909,N_14895,N_14947);
nand UO_910 (O_910,N_14965,N_14998);
and UO_911 (O_911,N_14951,N_14878);
nor UO_912 (O_912,N_14885,N_14935);
and UO_913 (O_913,N_14928,N_14975);
and UO_914 (O_914,N_14907,N_14897);
nand UO_915 (O_915,N_14962,N_14991);
and UO_916 (O_916,N_14993,N_14957);
or UO_917 (O_917,N_14882,N_14949);
or UO_918 (O_918,N_14936,N_14949);
nor UO_919 (O_919,N_14914,N_14917);
xnor UO_920 (O_920,N_14980,N_14896);
or UO_921 (O_921,N_14882,N_14988);
nand UO_922 (O_922,N_14948,N_14991);
and UO_923 (O_923,N_14893,N_14898);
and UO_924 (O_924,N_14879,N_14981);
nor UO_925 (O_925,N_14878,N_14974);
and UO_926 (O_926,N_14970,N_14937);
nor UO_927 (O_927,N_14985,N_14897);
or UO_928 (O_928,N_14899,N_14906);
nor UO_929 (O_929,N_14983,N_14998);
xnor UO_930 (O_930,N_14958,N_14896);
or UO_931 (O_931,N_14955,N_14923);
and UO_932 (O_932,N_14979,N_14910);
xor UO_933 (O_933,N_14888,N_14998);
and UO_934 (O_934,N_14893,N_14953);
and UO_935 (O_935,N_14927,N_14969);
and UO_936 (O_936,N_14909,N_14967);
nand UO_937 (O_937,N_14952,N_14910);
xnor UO_938 (O_938,N_14907,N_14958);
or UO_939 (O_939,N_14908,N_14975);
or UO_940 (O_940,N_14978,N_14887);
nand UO_941 (O_941,N_14902,N_14947);
xnor UO_942 (O_942,N_14991,N_14935);
and UO_943 (O_943,N_14899,N_14919);
or UO_944 (O_944,N_14930,N_14888);
and UO_945 (O_945,N_14988,N_14968);
and UO_946 (O_946,N_14992,N_14886);
and UO_947 (O_947,N_14964,N_14932);
and UO_948 (O_948,N_14888,N_14960);
xor UO_949 (O_949,N_14897,N_14968);
or UO_950 (O_950,N_14953,N_14918);
nor UO_951 (O_951,N_14941,N_14891);
xnor UO_952 (O_952,N_14942,N_14960);
nand UO_953 (O_953,N_14930,N_14984);
nor UO_954 (O_954,N_14959,N_14899);
nor UO_955 (O_955,N_14922,N_14911);
nand UO_956 (O_956,N_14879,N_14905);
and UO_957 (O_957,N_14969,N_14915);
nor UO_958 (O_958,N_14988,N_14952);
or UO_959 (O_959,N_14984,N_14997);
xor UO_960 (O_960,N_14966,N_14928);
nand UO_961 (O_961,N_14978,N_14945);
and UO_962 (O_962,N_14896,N_14972);
nand UO_963 (O_963,N_14910,N_14914);
xor UO_964 (O_964,N_14967,N_14889);
nand UO_965 (O_965,N_14928,N_14979);
and UO_966 (O_966,N_14978,N_14889);
and UO_967 (O_967,N_14885,N_14913);
nand UO_968 (O_968,N_14995,N_14909);
and UO_969 (O_969,N_14947,N_14980);
xor UO_970 (O_970,N_14957,N_14958);
nand UO_971 (O_971,N_14991,N_14981);
or UO_972 (O_972,N_14969,N_14981);
nand UO_973 (O_973,N_14892,N_14996);
or UO_974 (O_974,N_14988,N_14891);
xnor UO_975 (O_975,N_14885,N_14989);
nor UO_976 (O_976,N_14876,N_14996);
nand UO_977 (O_977,N_14882,N_14922);
nor UO_978 (O_978,N_14967,N_14901);
or UO_979 (O_979,N_14983,N_14978);
xor UO_980 (O_980,N_14975,N_14911);
or UO_981 (O_981,N_14905,N_14881);
nand UO_982 (O_982,N_14924,N_14987);
xor UO_983 (O_983,N_14990,N_14986);
nor UO_984 (O_984,N_14992,N_14880);
and UO_985 (O_985,N_14911,N_14992);
xnor UO_986 (O_986,N_14971,N_14965);
or UO_987 (O_987,N_14911,N_14959);
nor UO_988 (O_988,N_14877,N_14960);
nor UO_989 (O_989,N_14994,N_14989);
xnor UO_990 (O_990,N_14949,N_14951);
and UO_991 (O_991,N_14875,N_14885);
xor UO_992 (O_992,N_14943,N_14914);
or UO_993 (O_993,N_14988,N_14989);
nor UO_994 (O_994,N_14936,N_14975);
and UO_995 (O_995,N_14994,N_14902);
nand UO_996 (O_996,N_14896,N_14989);
or UO_997 (O_997,N_14907,N_14875);
nor UO_998 (O_998,N_14999,N_14993);
and UO_999 (O_999,N_14993,N_14918);
xor UO_1000 (O_1000,N_14944,N_14913);
or UO_1001 (O_1001,N_14990,N_14971);
or UO_1002 (O_1002,N_14876,N_14938);
xor UO_1003 (O_1003,N_14919,N_14986);
or UO_1004 (O_1004,N_14979,N_14950);
nor UO_1005 (O_1005,N_14876,N_14961);
nor UO_1006 (O_1006,N_14940,N_14945);
and UO_1007 (O_1007,N_14964,N_14896);
xor UO_1008 (O_1008,N_14915,N_14924);
nand UO_1009 (O_1009,N_14991,N_14918);
nand UO_1010 (O_1010,N_14896,N_14886);
nor UO_1011 (O_1011,N_14921,N_14911);
or UO_1012 (O_1012,N_14995,N_14982);
and UO_1013 (O_1013,N_14888,N_14989);
xnor UO_1014 (O_1014,N_14919,N_14937);
nor UO_1015 (O_1015,N_14912,N_14914);
nand UO_1016 (O_1016,N_14921,N_14939);
nor UO_1017 (O_1017,N_14942,N_14996);
nor UO_1018 (O_1018,N_14906,N_14904);
nor UO_1019 (O_1019,N_14946,N_14975);
nand UO_1020 (O_1020,N_14932,N_14885);
or UO_1021 (O_1021,N_14912,N_14921);
nand UO_1022 (O_1022,N_14960,N_14875);
or UO_1023 (O_1023,N_14955,N_14936);
nor UO_1024 (O_1024,N_14930,N_14938);
xnor UO_1025 (O_1025,N_14955,N_14879);
nor UO_1026 (O_1026,N_14909,N_14942);
or UO_1027 (O_1027,N_14932,N_14943);
nand UO_1028 (O_1028,N_14959,N_14912);
and UO_1029 (O_1029,N_14989,N_14930);
or UO_1030 (O_1030,N_14979,N_14991);
nand UO_1031 (O_1031,N_14969,N_14956);
and UO_1032 (O_1032,N_14970,N_14958);
nand UO_1033 (O_1033,N_14934,N_14944);
xor UO_1034 (O_1034,N_14877,N_14902);
nor UO_1035 (O_1035,N_14879,N_14898);
nand UO_1036 (O_1036,N_14937,N_14951);
nand UO_1037 (O_1037,N_14947,N_14925);
xnor UO_1038 (O_1038,N_14967,N_14976);
or UO_1039 (O_1039,N_14896,N_14982);
and UO_1040 (O_1040,N_14993,N_14969);
xnor UO_1041 (O_1041,N_14928,N_14978);
or UO_1042 (O_1042,N_14908,N_14932);
nand UO_1043 (O_1043,N_14923,N_14887);
and UO_1044 (O_1044,N_14901,N_14897);
and UO_1045 (O_1045,N_14928,N_14968);
and UO_1046 (O_1046,N_14974,N_14969);
xnor UO_1047 (O_1047,N_14911,N_14905);
xor UO_1048 (O_1048,N_14927,N_14895);
or UO_1049 (O_1049,N_14991,N_14922);
nand UO_1050 (O_1050,N_14895,N_14928);
and UO_1051 (O_1051,N_14895,N_14899);
and UO_1052 (O_1052,N_14927,N_14881);
nor UO_1053 (O_1053,N_14963,N_14954);
and UO_1054 (O_1054,N_14945,N_14924);
or UO_1055 (O_1055,N_14957,N_14909);
xor UO_1056 (O_1056,N_14972,N_14927);
and UO_1057 (O_1057,N_14996,N_14910);
and UO_1058 (O_1058,N_14913,N_14938);
and UO_1059 (O_1059,N_14986,N_14896);
and UO_1060 (O_1060,N_14965,N_14928);
nand UO_1061 (O_1061,N_14893,N_14987);
nand UO_1062 (O_1062,N_14972,N_14893);
or UO_1063 (O_1063,N_14925,N_14883);
nand UO_1064 (O_1064,N_14916,N_14905);
nand UO_1065 (O_1065,N_14944,N_14971);
or UO_1066 (O_1066,N_14929,N_14974);
nor UO_1067 (O_1067,N_14876,N_14985);
nor UO_1068 (O_1068,N_14932,N_14940);
xnor UO_1069 (O_1069,N_14994,N_14927);
nand UO_1070 (O_1070,N_14975,N_14876);
xor UO_1071 (O_1071,N_14993,N_14963);
xor UO_1072 (O_1072,N_14922,N_14968);
nand UO_1073 (O_1073,N_14949,N_14979);
nor UO_1074 (O_1074,N_14940,N_14914);
xor UO_1075 (O_1075,N_14933,N_14993);
and UO_1076 (O_1076,N_14933,N_14999);
and UO_1077 (O_1077,N_14897,N_14940);
nor UO_1078 (O_1078,N_14887,N_14990);
nor UO_1079 (O_1079,N_14910,N_14930);
nand UO_1080 (O_1080,N_14894,N_14937);
or UO_1081 (O_1081,N_14961,N_14975);
xnor UO_1082 (O_1082,N_14941,N_14952);
xnor UO_1083 (O_1083,N_14910,N_14911);
and UO_1084 (O_1084,N_14923,N_14967);
nor UO_1085 (O_1085,N_14898,N_14895);
nand UO_1086 (O_1086,N_14934,N_14940);
xor UO_1087 (O_1087,N_14997,N_14950);
nand UO_1088 (O_1088,N_14902,N_14941);
or UO_1089 (O_1089,N_14992,N_14970);
or UO_1090 (O_1090,N_14884,N_14978);
and UO_1091 (O_1091,N_14975,N_14962);
and UO_1092 (O_1092,N_14883,N_14987);
or UO_1093 (O_1093,N_14995,N_14891);
or UO_1094 (O_1094,N_14886,N_14920);
or UO_1095 (O_1095,N_14993,N_14951);
xor UO_1096 (O_1096,N_14917,N_14903);
nand UO_1097 (O_1097,N_14974,N_14928);
or UO_1098 (O_1098,N_14898,N_14907);
or UO_1099 (O_1099,N_14994,N_14953);
and UO_1100 (O_1100,N_14930,N_14954);
nand UO_1101 (O_1101,N_14897,N_14976);
or UO_1102 (O_1102,N_14882,N_14931);
xor UO_1103 (O_1103,N_14915,N_14962);
nor UO_1104 (O_1104,N_14948,N_14894);
nand UO_1105 (O_1105,N_14932,N_14902);
nor UO_1106 (O_1106,N_14884,N_14928);
or UO_1107 (O_1107,N_14902,N_14914);
or UO_1108 (O_1108,N_14994,N_14962);
or UO_1109 (O_1109,N_14883,N_14908);
or UO_1110 (O_1110,N_14987,N_14965);
xor UO_1111 (O_1111,N_14964,N_14989);
and UO_1112 (O_1112,N_14886,N_14963);
nor UO_1113 (O_1113,N_14900,N_14894);
nand UO_1114 (O_1114,N_14927,N_14890);
or UO_1115 (O_1115,N_14967,N_14886);
nand UO_1116 (O_1116,N_14930,N_14962);
nor UO_1117 (O_1117,N_14881,N_14987);
and UO_1118 (O_1118,N_14876,N_14924);
nor UO_1119 (O_1119,N_14962,N_14875);
xor UO_1120 (O_1120,N_14992,N_14994);
and UO_1121 (O_1121,N_14924,N_14939);
nand UO_1122 (O_1122,N_14889,N_14994);
nand UO_1123 (O_1123,N_14986,N_14980);
xnor UO_1124 (O_1124,N_14877,N_14889);
or UO_1125 (O_1125,N_14878,N_14939);
and UO_1126 (O_1126,N_14890,N_14998);
and UO_1127 (O_1127,N_14886,N_14908);
nand UO_1128 (O_1128,N_14893,N_14962);
or UO_1129 (O_1129,N_14948,N_14999);
or UO_1130 (O_1130,N_14920,N_14957);
and UO_1131 (O_1131,N_14898,N_14982);
nor UO_1132 (O_1132,N_14926,N_14974);
xnor UO_1133 (O_1133,N_14882,N_14929);
or UO_1134 (O_1134,N_14916,N_14985);
and UO_1135 (O_1135,N_14918,N_14932);
xnor UO_1136 (O_1136,N_14903,N_14933);
nor UO_1137 (O_1137,N_14907,N_14921);
xnor UO_1138 (O_1138,N_14965,N_14907);
xor UO_1139 (O_1139,N_14986,N_14954);
and UO_1140 (O_1140,N_14905,N_14884);
xor UO_1141 (O_1141,N_14941,N_14875);
or UO_1142 (O_1142,N_14887,N_14877);
nor UO_1143 (O_1143,N_14884,N_14983);
or UO_1144 (O_1144,N_14948,N_14982);
or UO_1145 (O_1145,N_14902,N_14921);
or UO_1146 (O_1146,N_14953,N_14991);
or UO_1147 (O_1147,N_14965,N_14930);
and UO_1148 (O_1148,N_14978,N_14922);
nor UO_1149 (O_1149,N_14945,N_14927);
or UO_1150 (O_1150,N_14880,N_14996);
or UO_1151 (O_1151,N_14952,N_14897);
nand UO_1152 (O_1152,N_14876,N_14946);
nor UO_1153 (O_1153,N_14925,N_14914);
nor UO_1154 (O_1154,N_14935,N_14877);
and UO_1155 (O_1155,N_14911,N_14982);
xnor UO_1156 (O_1156,N_14891,N_14887);
nor UO_1157 (O_1157,N_14977,N_14997);
or UO_1158 (O_1158,N_14923,N_14999);
nand UO_1159 (O_1159,N_14963,N_14982);
and UO_1160 (O_1160,N_14916,N_14909);
nand UO_1161 (O_1161,N_14931,N_14922);
or UO_1162 (O_1162,N_14981,N_14970);
nor UO_1163 (O_1163,N_14890,N_14973);
nor UO_1164 (O_1164,N_14898,N_14919);
and UO_1165 (O_1165,N_14903,N_14902);
or UO_1166 (O_1166,N_14980,N_14991);
nor UO_1167 (O_1167,N_14916,N_14893);
and UO_1168 (O_1168,N_14930,N_14875);
and UO_1169 (O_1169,N_14944,N_14939);
or UO_1170 (O_1170,N_14974,N_14910);
xnor UO_1171 (O_1171,N_14945,N_14984);
and UO_1172 (O_1172,N_14929,N_14967);
or UO_1173 (O_1173,N_14916,N_14978);
and UO_1174 (O_1174,N_14895,N_14956);
xor UO_1175 (O_1175,N_14959,N_14949);
nor UO_1176 (O_1176,N_14932,N_14924);
and UO_1177 (O_1177,N_14953,N_14923);
nand UO_1178 (O_1178,N_14909,N_14937);
or UO_1179 (O_1179,N_14955,N_14907);
nand UO_1180 (O_1180,N_14884,N_14900);
nand UO_1181 (O_1181,N_14993,N_14926);
and UO_1182 (O_1182,N_14942,N_14881);
nand UO_1183 (O_1183,N_14897,N_14890);
or UO_1184 (O_1184,N_14884,N_14934);
or UO_1185 (O_1185,N_14880,N_14933);
nand UO_1186 (O_1186,N_14939,N_14902);
nor UO_1187 (O_1187,N_14938,N_14922);
nand UO_1188 (O_1188,N_14987,N_14915);
and UO_1189 (O_1189,N_14953,N_14920);
or UO_1190 (O_1190,N_14964,N_14960);
nand UO_1191 (O_1191,N_14995,N_14988);
xor UO_1192 (O_1192,N_14945,N_14931);
and UO_1193 (O_1193,N_14975,N_14984);
and UO_1194 (O_1194,N_14919,N_14875);
xor UO_1195 (O_1195,N_14896,N_14930);
or UO_1196 (O_1196,N_14962,N_14960);
and UO_1197 (O_1197,N_14993,N_14937);
or UO_1198 (O_1198,N_14881,N_14926);
nor UO_1199 (O_1199,N_14938,N_14984);
and UO_1200 (O_1200,N_14978,N_14897);
and UO_1201 (O_1201,N_14895,N_14968);
and UO_1202 (O_1202,N_14970,N_14906);
or UO_1203 (O_1203,N_14888,N_14967);
xor UO_1204 (O_1204,N_14912,N_14990);
nand UO_1205 (O_1205,N_14891,N_14897);
and UO_1206 (O_1206,N_14915,N_14993);
nand UO_1207 (O_1207,N_14948,N_14880);
nand UO_1208 (O_1208,N_14931,N_14881);
nand UO_1209 (O_1209,N_14950,N_14989);
and UO_1210 (O_1210,N_14891,N_14900);
nand UO_1211 (O_1211,N_14992,N_14958);
or UO_1212 (O_1212,N_14996,N_14945);
nand UO_1213 (O_1213,N_14885,N_14958);
nor UO_1214 (O_1214,N_14934,N_14899);
nand UO_1215 (O_1215,N_14900,N_14920);
xor UO_1216 (O_1216,N_14943,N_14899);
or UO_1217 (O_1217,N_14880,N_14964);
or UO_1218 (O_1218,N_14943,N_14896);
or UO_1219 (O_1219,N_14940,N_14921);
nor UO_1220 (O_1220,N_14996,N_14970);
nor UO_1221 (O_1221,N_14924,N_14891);
and UO_1222 (O_1222,N_14893,N_14964);
nor UO_1223 (O_1223,N_14992,N_14948);
xor UO_1224 (O_1224,N_14914,N_14941);
and UO_1225 (O_1225,N_14951,N_14954);
or UO_1226 (O_1226,N_14942,N_14930);
nand UO_1227 (O_1227,N_14967,N_14884);
nand UO_1228 (O_1228,N_14975,N_14892);
nor UO_1229 (O_1229,N_14999,N_14934);
xor UO_1230 (O_1230,N_14996,N_14950);
xnor UO_1231 (O_1231,N_14999,N_14911);
nor UO_1232 (O_1232,N_14877,N_14881);
nand UO_1233 (O_1233,N_14988,N_14974);
and UO_1234 (O_1234,N_14913,N_14940);
and UO_1235 (O_1235,N_14917,N_14949);
or UO_1236 (O_1236,N_14961,N_14951);
xor UO_1237 (O_1237,N_14894,N_14955);
xnor UO_1238 (O_1238,N_14968,N_14982);
xor UO_1239 (O_1239,N_14973,N_14879);
nor UO_1240 (O_1240,N_14976,N_14947);
nor UO_1241 (O_1241,N_14964,N_14995);
or UO_1242 (O_1242,N_14918,N_14985);
nor UO_1243 (O_1243,N_14921,N_14964);
nor UO_1244 (O_1244,N_14997,N_14957);
nor UO_1245 (O_1245,N_14902,N_14908);
or UO_1246 (O_1246,N_14932,N_14916);
or UO_1247 (O_1247,N_14996,N_14887);
and UO_1248 (O_1248,N_14907,N_14977);
and UO_1249 (O_1249,N_14997,N_14927);
nand UO_1250 (O_1250,N_14901,N_14906);
nand UO_1251 (O_1251,N_14979,N_14937);
xnor UO_1252 (O_1252,N_14939,N_14879);
xor UO_1253 (O_1253,N_14907,N_14889);
nand UO_1254 (O_1254,N_14941,N_14901);
and UO_1255 (O_1255,N_14894,N_14983);
xnor UO_1256 (O_1256,N_14974,N_14893);
or UO_1257 (O_1257,N_14905,N_14995);
and UO_1258 (O_1258,N_14972,N_14956);
nand UO_1259 (O_1259,N_14903,N_14943);
xor UO_1260 (O_1260,N_14981,N_14904);
or UO_1261 (O_1261,N_14994,N_14891);
and UO_1262 (O_1262,N_14969,N_14991);
and UO_1263 (O_1263,N_14980,N_14992);
and UO_1264 (O_1264,N_14945,N_14899);
and UO_1265 (O_1265,N_14970,N_14969);
nor UO_1266 (O_1266,N_14988,N_14944);
and UO_1267 (O_1267,N_14988,N_14975);
nand UO_1268 (O_1268,N_14920,N_14969);
nor UO_1269 (O_1269,N_14882,N_14965);
or UO_1270 (O_1270,N_14998,N_14935);
and UO_1271 (O_1271,N_14913,N_14935);
nand UO_1272 (O_1272,N_14929,N_14930);
nor UO_1273 (O_1273,N_14924,N_14937);
or UO_1274 (O_1274,N_14975,N_14993);
and UO_1275 (O_1275,N_14955,N_14900);
nor UO_1276 (O_1276,N_14936,N_14912);
and UO_1277 (O_1277,N_14897,N_14964);
nor UO_1278 (O_1278,N_14973,N_14962);
nand UO_1279 (O_1279,N_14949,N_14905);
or UO_1280 (O_1280,N_14892,N_14930);
or UO_1281 (O_1281,N_14931,N_14929);
nor UO_1282 (O_1282,N_14987,N_14997);
xnor UO_1283 (O_1283,N_14923,N_14943);
and UO_1284 (O_1284,N_14917,N_14981);
or UO_1285 (O_1285,N_14908,N_14985);
xor UO_1286 (O_1286,N_14908,N_14945);
or UO_1287 (O_1287,N_14905,N_14932);
or UO_1288 (O_1288,N_14929,N_14883);
or UO_1289 (O_1289,N_14958,N_14893);
nor UO_1290 (O_1290,N_14879,N_14915);
nand UO_1291 (O_1291,N_14967,N_14965);
xnor UO_1292 (O_1292,N_14978,N_14937);
nand UO_1293 (O_1293,N_14941,N_14888);
nor UO_1294 (O_1294,N_14924,N_14934);
nor UO_1295 (O_1295,N_14885,N_14900);
or UO_1296 (O_1296,N_14895,N_14958);
or UO_1297 (O_1297,N_14883,N_14989);
nand UO_1298 (O_1298,N_14938,N_14889);
nand UO_1299 (O_1299,N_14963,N_14991);
xor UO_1300 (O_1300,N_14994,N_14885);
and UO_1301 (O_1301,N_14942,N_14931);
nand UO_1302 (O_1302,N_14902,N_14917);
nand UO_1303 (O_1303,N_14991,N_14882);
xnor UO_1304 (O_1304,N_14975,N_14912);
xnor UO_1305 (O_1305,N_14918,N_14888);
nand UO_1306 (O_1306,N_14947,N_14914);
xor UO_1307 (O_1307,N_14991,N_14946);
nand UO_1308 (O_1308,N_14941,N_14900);
xnor UO_1309 (O_1309,N_14936,N_14996);
and UO_1310 (O_1310,N_14970,N_14956);
or UO_1311 (O_1311,N_14985,N_14962);
xnor UO_1312 (O_1312,N_14931,N_14892);
nand UO_1313 (O_1313,N_14994,N_14906);
or UO_1314 (O_1314,N_14958,N_14948);
or UO_1315 (O_1315,N_14908,N_14998);
xor UO_1316 (O_1316,N_14945,N_14906);
or UO_1317 (O_1317,N_14887,N_14988);
and UO_1318 (O_1318,N_14945,N_14913);
or UO_1319 (O_1319,N_14976,N_14982);
and UO_1320 (O_1320,N_14961,N_14892);
xnor UO_1321 (O_1321,N_14989,N_14940);
and UO_1322 (O_1322,N_14906,N_14958);
or UO_1323 (O_1323,N_14888,N_14939);
or UO_1324 (O_1324,N_14947,N_14893);
and UO_1325 (O_1325,N_14964,N_14967);
nor UO_1326 (O_1326,N_14980,N_14944);
or UO_1327 (O_1327,N_14957,N_14973);
or UO_1328 (O_1328,N_14972,N_14996);
nand UO_1329 (O_1329,N_14978,N_14940);
or UO_1330 (O_1330,N_14959,N_14948);
xor UO_1331 (O_1331,N_14939,N_14903);
nor UO_1332 (O_1332,N_14967,N_14944);
nand UO_1333 (O_1333,N_14958,N_14965);
and UO_1334 (O_1334,N_14888,N_14956);
xor UO_1335 (O_1335,N_14947,N_14915);
xnor UO_1336 (O_1336,N_14961,N_14912);
and UO_1337 (O_1337,N_14965,N_14948);
nand UO_1338 (O_1338,N_14876,N_14954);
and UO_1339 (O_1339,N_14969,N_14921);
xor UO_1340 (O_1340,N_14996,N_14890);
nor UO_1341 (O_1341,N_14898,N_14891);
nand UO_1342 (O_1342,N_14959,N_14976);
or UO_1343 (O_1343,N_14912,N_14927);
nand UO_1344 (O_1344,N_14904,N_14955);
or UO_1345 (O_1345,N_14966,N_14983);
or UO_1346 (O_1346,N_14968,N_14964);
xnor UO_1347 (O_1347,N_14984,N_14911);
or UO_1348 (O_1348,N_14913,N_14987);
and UO_1349 (O_1349,N_14923,N_14894);
nor UO_1350 (O_1350,N_14978,N_14909);
nand UO_1351 (O_1351,N_14944,N_14905);
xor UO_1352 (O_1352,N_14928,N_14915);
nand UO_1353 (O_1353,N_14892,N_14997);
or UO_1354 (O_1354,N_14997,N_14898);
nand UO_1355 (O_1355,N_14944,N_14941);
xnor UO_1356 (O_1356,N_14920,N_14923);
and UO_1357 (O_1357,N_14897,N_14919);
nor UO_1358 (O_1358,N_14994,N_14951);
and UO_1359 (O_1359,N_14889,N_14880);
or UO_1360 (O_1360,N_14877,N_14950);
nor UO_1361 (O_1361,N_14923,N_14884);
nand UO_1362 (O_1362,N_14941,N_14895);
and UO_1363 (O_1363,N_14991,N_14934);
and UO_1364 (O_1364,N_14957,N_14942);
nand UO_1365 (O_1365,N_14971,N_14922);
and UO_1366 (O_1366,N_14933,N_14879);
nand UO_1367 (O_1367,N_14914,N_14895);
nor UO_1368 (O_1368,N_14921,N_14890);
xnor UO_1369 (O_1369,N_14934,N_14983);
or UO_1370 (O_1370,N_14933,N_14964);
xnor UO_1371 (O_1371,N_14902,N_14880);
and UO_1372 (O_1372,N_14943,N_14941);
nand UO_1373 (O_1373,N_14958,N_14923);
nand UO_1374 (O_1374,N_14948,N_14911);
and UO_1375 (O_1375,N_14988,N_14971);
nand UO_1376 (O_1376,N_14982,N_14881);
nand UO_1377 (O_1377,N_14925,N_14932);
xnor UO_1378 (O_1378,N_14961,N_14994);
nand UO_1379 (O_1379,N_14984,N_14995);
or UO_1380 (O_1380,N_14908,N_14987);
xor UO_1381 (O_1381,N_14939,N_14954);
nor UO_1382 (O_1382,N_14881,N_14923);
xnor UO_1383 (O_1383,N_14881,N_14906);
nor UO_1384 (O_1384,N_14894,N_14986);
and UO_1385 (O_1385,N_14977,N_14980);
nor UO_1386 (O_1386,N_14876,N_14914);
nand UO_1387 (O_1387,N_14995,N_14974);
and UO_1388 (O_1388,N_14912,N_14963);
xor UO_1389 (O_1389,N_14990,N_14982);
nor UO_1390 (O_1390,N_14977,N_14912);
nand UO_1391 (O_1391,N_14983,N_14984);
nand UO_1392 (O_1392,N_14988,N_14878);
or UO_1393 (O_1393,N_14912,N_14932);
or UO_1394 (O_1394,N_14926,N_14996);
and UO_1395 (O_1395,N_14952,N_14972);
nor UO_1396 (O_1396,N_14895,N_14969);
or UO_1397 (O_1397,N_14961,N_14934);
nor UO_1398 (O_1398,N_14879,N_14903);
nand UO_1399 (O_1399,N_14938,N_14904);
or UO_1400 (O_1400,N_14939,N_14963);
nand UO_1401 (O_1401,N_14928,N_14882);
xnor UO_1402 (O_1402,N_14938,N_14989);
or UO_1403 (O_1403,N_14875,N_14947);
or UO_1404 (O_1404,N_14946,N_14883);
nand UO_1405 (O_1405,N_14948,N_14892);
or UO_1406 (O_1406,N_14914,N_14919);
nor UO_1407 (O_1407,N_14931,N_14921);
and UO_1408 (O_1408,N_14891,N_14968);
xnor UO_1409 (O_1409,N_14936,N_14976);
nand UO_1410 (O_1410,N_14933,N_14894);
nand UO_1411 (O_1411,N_14995,N_14898);
nor UO_1412 (O_1412,N_14906,N_14927);
nand UO_1413 (O_1413,N_14905,N_14959);
and UO_1414 (O_1414,N_14941,N_14925);
nand UO_1415 (O_1415,N_14901,N_14903);
and UO_1416 (O_1416,N_14980,N_14993);
xnor UO_1417 (O_1417,N_14881,N_14944);
xor UO_1418 (O_1418,N_14893,N_14955);
nand UO_1419 (O_1419,N_14975,N_14933);
and UO_1420 (O_1420,N_14946,N_14979);
or UO_1421 (O_1421,N_14875,N_14958);
nand UO_1422 (O_1422,N_14954,N_14929);
xnor UO_1423 (O_1423,N_14986,N_14921);
nand UO_1424 (O_1424,N_14963,N_14953);
nand UO_1425 (O_1425,N_14969,N_14931);
and UO_1426 (O_1426,N_14919,N_14949);
or UO_1427 (O_1427,N_14976,N_14941);
xnor UO_1428 (O_1428,N_14904,N_14958);
nand UO_1429 (O_1429,N_14893,N_14903);
xnor UO_1430 (O_1430,N_14936,N_14939);
or UO_1431 (O_1431,N_14971,N_14887);
xor UO_1432 (O_1432,N_14891,N_14931);
nand UO_1433 (O_1433,N_14967,N_14953);
or UO_1434 (O_1434,N_14898,N_14901);
xor UO_1435 (O_1435,N_14883,N_14947);
nand UO_1436 (O_1436,N_14912,N_14895);
and UO_1437 (O_1437,N_14910,N_14899);
or UO_1438 (O_1438,N_14930,N_14920);
and UO_1439 (O_1439,N_14937,N_14945);
nor UO_1440 (O_1440,N_14888,N_14982);
and UO_1441 (O_1441,N_14963,N_14879);
nor UO_1442 (O_1442,N_14902,N_14984);
and UO_1443 (O_1443,N_14958,N_14911);
xor UO_1444 (O_1444,N_14894,N_14995);
and UO_1445 (O_1445,N_14952,N_14960);
or UO_1446 (O_1446,N_14932,N_14893);
nor UO_1447 (O_1447,N_14908,N_14876);
and UO_1448 (O_1448,N_14998,N_14931);
nor UO_1449 (O_1449,N_14963,N_14884);
xnor UO_1450 (O_1450,N_14918,N_14930);
and UO_1451 (O_1451,N_14918,N_14924);
nor UO_1452 (O_1452,N_14938,N_14885);
nand UO_1453 (O_1453,N_14917,N_14995);
nor UO_1454 (O_1454,N_14990,N_14908);
or UO_1455 (O_1455,N_14937,N_14902);
or UO_1456 (O_1456,N_14996,N_14883);
and UO_1457 (O_1457,N_14893,N_14930);
and UO_1458 (O_1458,N_14949,N_14939);
or UO_1459 (O_1459,N_14894,N_14901);
xnor UO_1460 (O_1460,N_14931,N_14995);
or UO_1461 (O_1461,N_14891,N_14926);
nand UO_1462 (O_1462,N_14914,N_14986);
and UO_1463 (O_1463,N_14918,N_14974);
xor UO_1464 (O_1464,N_14929,N_14986);
xor UO_1465 (O_1465,N_14948,N_14985);
and UO_1466 (O_1466,N_14928,N_14896);
or UO_1467 (O_1467,N_14918,N_14984);
nand UO_1468 (O_1468,N_14958,N_14935);
and UO_1469 (O_1469,N_14979,N_14913);
or UO_1470 (O_1470,N_14917,N_14884);
or UO_1471 (O_1471,N_14992,N_14950);
nor UO_1472 (O_1472,N_14969,N_14945);
and UO_1473 (O_1473,N_14915,N_14974);
nand UO_1474 (O_1474,N_14875,N_14999);
or UO_1475 (O_1475,N_14903,N_14882);
xor UO_1476 (O_1476,N_14985,N_14947);
or UO_1477 (O_1477,N_14923,N_14931);
nand UO_1478 (O_1478,N_14998,N_14918);
nor UO_1479 (O_1479,N_14899,N_14904);
and UO_1480 (O_1480,N_14898,N_14999);
and UO_1481 (O_1481,N_14888,N_14943);
and UO_1482 (O_1482,N_14949,N_14934);
xor UO_1483 (O_1483,N_14887,N_14973);
nor UO_1484 (O_1484,N_14994,N_14919);
nor UO_1485 (O_1485,N_14905,N_14878);
nand UO_1486 (O_1486,N_14932,N_14946);
nor UO_1487 (O_1487,N_14950,N_14956);
xor UO_1488 (O_1488,N_14988,N_14885);
or UO_1489 (O_1489,N_14904,N_14939);
nor UO_1490 (O_1490,N_14953,N_14878);
and UO_1491 (O_1491,N_14984,N_14910);
nor UO_1492 (O_1492,N_14897,N_14913);
nand UO_1493 (O_1493,N_14881,N_14916);
or UO_1494 (O_1494,N_14955,N_14897);
xor UO_1495 (O_1495,N_14908,N_14897);
or UO_1496 (O_1496,N_14967,N_14919);
and UO_1497 (O_1497,N_14982,N_14973);
nand UO_1498 (O_1498,N_14979,N_14985);
or UO_1499 (O_1499,N_14987,N_14886);
nor UO_1500 (O_1500,N_14970,N_14909);
or UO_1501 (O_1501,N_14931,N_14979);
nor UO_1502 (O_1502,N_14970,N_14960);
or UO_1503 (O_1503,N_14999,N_14935);
or UO_1504 (O_1504,N_14893,N_14943);
or UO_1505 (O_1505,N_14985,N_14917);
and UO_1506 (O_1506,N_14908,N_14981);
nand UO_1507 (O_1507,N_14927,N_14966);
or UO_1508 (O_1508,N_14904,N_14886);
nor UO_1509 (O_1509,N_14913,N_14936);
nand UO_1510 (O_1510,N_14932,N_14917);
nand UO_1511 (O_1511,N_14994,N_14920);
nand UO_1512 (O_1512,N_14968,N_14996);
nor UO_1513 (O_1513,N_14985,N_14905);
nor UO_1514 (O_1514,N_14980,N_14907);
and UO_1515 (O_1515,N_14927,N_14995);
nor UO_1516 (O_1516,N_14988,N_14875);
and UO_1517 (O_1517,N_14985,N_14923);
nand UO_1518 (O_1518,N_14896,N_14894);
and UO_1519 (O_1519,N_14952,N_14997);
nand UO_1520 (O_1520,N_14896,N_14889);
xnor UO_1521 (O_1521,N_14975,N_14905);
xor UO_1522 (O_1522,N_14886,N_14922);
or UO_1523 (O_1523,N_14927,N_14901);
or UO_1524 (O_1524,N_14956,N_14904);
or UO_1525 (O_1525,N_14992,N_14888);
and UO_1526 (O_1526,N_14968,N_14984);
and UO_1527 (O_1527,N_14984,N_14955);
or UO_1528 (O_1528,N_14890,N_14879);
nand UO_1529 (O_1529,N_14921,N_14909);
or UO_1530 (O_1530,N_14943,N_14998);
nand UO_1531 (O_1531,N_14917,N_14889);
and UO_1532 (O_1532,N_14902,N_14973);
and UO_1533 (O_1533,N_14988,N_14982);
nor UO_1534 (O_1534,N_14917,N_14956);
nor UO_1535 (O_1535,N_14953,N_14989);
and UO_1536 (O_1536,N_14938,N_14932);
nor UO_1537 (O_1537,N_14941,N_14938);
and UO_1538 (O_1538,N_14879,N_14951);
or UO_1539 (O_1539,N_14918,N_14904);
nor UO_1540 (O_1540,N_14936,N_14933);
xor UO_1541 (O_1541,N_14962,N_14961);
and UO_1542 (O_1542,N_14990,N_14937);
nand UO_1543 (O_1543,N_14979,N_14977);
nor UO_1544 (O_1544,N_14983,N_14888);
xor UO_1545 (O_1545,N_14907,N_14934);
or UO_1546 (O_1546,N_14952,N_14929);
nand UO_1547 (O_1547,N_14983,N_14921);
nor UO_1548 (O_1548,N_14895,N_14904);
xnor UO_1549 (O_1549,N_14910,N_14894);
nand UO_1550 (O_1550,N_14952,N_14924);
or UO_1551 (O_1551,N_14925,N_14972);
or UO_1552 (O_1552,N_14905,N_14919);
nand UO_1553 (O_1553,N_14897,N_14912);
and UO_1554 (O_1554,N_14972,N_14989);
nand UO_1555 (O_1555,N_14899,N_14875);
xor UO_1556 (O_1556,N_14885,N_14922);
or UO_1557 (O_1557,N_14880,N_14895);
nor UO_1558 (O_1558,N_14909,N_14876);
nand UO_1559 (O_1559,N_14946,N_14931);
nand UO_1560 (O_1560,N_14942,N_14994);
or UO_1561 (O_1561,N_14877,N_14934);
and UO_1562 (O_1562,N_14930,N_14907);
or UO_1563 (O_1563,N_14979,N_14943);
and UO_1564 (O_1564,N_14975,N_14931);
nand UO_1565 (O_1565,N_14939,N_14994);
nor UO_1566 (O_1566,N_14959,N_14955);
and UO_1567 (O_1567,N_14973,N_14915);
or UO_1568 (O_1568,N_14959,N_14882);
and UO_1569 (O_1569,N_14967,N_14936);
or UO_1570 (O_1570,N_14926,N_14995);
or UO_1571 (O_1571,N_14886,N_14972);
nand UO_1572 (O_1572,N_14948,N_14900);
and UO_1573 (O_1573,N_14875,N_14921);
xnor UO_1574 (O_1574,N_14987,N_14897);
nand UO_1575 (O_1575,N_14886,N_14957);
or UO_1576 (O_1576,N_14954,N_14977);
or UO_1577 (O_1577,N_14927,N_14980);
and UO_1578 (O_1578,N_14976,N_14917);
nor UO_1579 (O_1579,N_14981,N_14954);
or UO_1580 (O_1580,N_14936,N_14900);
and UO_1581 (O_1581,N_14881,N_14880);
or UO_1582 (O_1582,N_14905,N_14982);
or UO_1583 (O_1583,N_14963,N_14972);
xnor UO_1584 (O_1584,N_14984,N_14879);
and UO_1585 (O_1585,N_14954,N_14931);
xor UO_1586 (O_1586,N_14916,N_14891);
or UO_1587 (O_1587,N_14965,N_14973);
or UO_1588 (O_1588,N_14916,N_14986);
nor UO_1589 (O_1589,N_14993,N_14939);
nand UO_1590 (O_1590,N_14959,N_14891);
and UO_1591 (O_1591,N_14933,N_14968);
and UO_1592 (O_1592,N_14910,N_14994);
and UO_1593 (O_1593,N_14992,N_14984);
or UO_1594 (O_1594,N_14918,N_14917);
nand UO_1595 (O_1595,N_14927,N_14884);
nand UO_1596 (O_1596,N_14993,N_14921);
and UO_1597 (O_1597,N_14996,N_14938);
xnor UO_1598 (O_1598,N_14915,N_14904);
or UO_1599 (O_1599,N_14966,N_14991);
and UO_1600 (O_1600,N_14980,N_14984);
nand UO_1601 (O_1601,N_14978,N_14968);
or UO_1602 (O_1602,N_14972,N_14973);
nor UO_1603 (O_1603,N_14925,N_14958);
nor UO_1604 (O_1604,N_14899,N_14932);
or UO_1605 (O_1605,N_14902,N_14981);
nor UO_1606 (O_1606,N_14921,N_14968);
nand UO_1607 (O_1607,N_14956,N_14902);
or UO_1608 (O_1608,N_14945,N_14875);
and UO_1609 (O_1609,N_14927,N_14953);
and UO_1610 (O_1610,N_14942,N_14973);
nand UO_1611 (O_1611,N_14937,N_14994);
xnor UO_1612 (O_1612,N_14993,N_14959);
nand UO_1613 (O_1613,N_14926,N_14961);
xnor UO_1614 (O_1614,N_14902,N_14920);
nand UO_1615 (O_1615,N_14972,N_14889);
and UO_1616 (O_1616,N_14913,N_14880);
nand UO_1617 (O_1617,N_14946,N_14880);
nand UO_1618 (O_1618,N_14897,N_14899);
nand UO_1619 (O_1619,N_14987,N_14937);
and UO_1620 (O_1620,N_14980,N_14911);
and UO_1621 (O_1621,N_14940,N_14903);
or UO_1622 (O_1622,N_14982,N_14924);
xor UO_1623 (O_1623,N_14937,N_14930);
nor UO_1624 (O_1624,N_14937,N_14995);
or UO_1625 (O_1625,N_14985,N_14883);
nor UO_1626 (O_1626,N_14952,N_14902);
nor UO_1627 (O_1627,N_14938,N_14966);
nand UO_1628 (O_1628,N_14959,N_14998);
nor UO_1629 (O_1629,N_14996,N_14917);
and UO_1630 (O_1630,N_14947,N_14911);
or UO_1631 (O_1631,N_14915,N_14939);
nand UO_1632 (O_1632,N_14954,N_14996);
nand UO_1633 (O_1633,N_14995,N_14940);
and UO_1634 (O_1634,N_14978,N_14896);
nand UO_1635 (O_1635,N_14983,N_14939);
and UO_1636 (O_1636,N_14949,N_14937);
xnor UO_1637 (O_1637,N_14972,N_14982);
xor UO_1638 (O_1638,N_14966,N_14965);
or UO_1639 (O_1639,N_14892,N_14991);
nand UO_1640 (O_1640,N_14902,N_14895);
nor UO_1641 (O_1641,N_14891,N_14921);
nand UO_1642 (O_1642,N_14906,N_14915);
and UO_1643 (O_1643,N_14894,N_14884);
or UO_1644 (O_1644,N_14917,N_14909);
or UO_1645 (O_1645,N_14995,N_14876);
or UO_1646 (O_1646,N_14976,N_14943);
nand UO_1647 (O_1647,N_14896,N_14892);
nand UO_1648 (O_1648,N_14927,N_14877);
nand UO_1649 (O_1649,N_14932,N_14962);
xnor UO_1650 (O_1650,N_14918,N_14966);
and UO_1651 (O_1651,N_14992,N_14956);
nand UO_1652 (O_1652,N_14989,N_14914);
nor UO_1653 (O_1653,N_14888,N_14993);
nand UO_1654 (O_1654,N_14980,N_14983);
nand UO_1655 (O_1655,N_14937,N_14967);
nand UO_1656 (O_1656,N_14930,N_14905);
xnor UO_1657 (O_1657,N_14926,N_14932);
nand UO_1658 (O_1658,N_14910,N_14991);
or UO_1659 (O_1659,N_14956,N_14984);
and UO_1660 (O_1660,N_14910,N_14966);
and UO_1661 (O_1661,N_14943,N_14883);
and UO_1662 (O_1662,N_14898,N_14928);
nand UO_1663 (O_1663,N_14883,N_14899);
or UO_1664 (O_1664,N_14923,N_14892);
xor UO_1665 (O_1665,N_14980,N_14918);
nor UO_1666 (O_1666,N_14888,N_14903);
nand UO_1667 (O_1667,N_14936,N_14924);
and UO_1668 (O_1668,N_14931,N_14967);
nor UO_1669 (O_1669,N_14959,N_14893);
and UO_1670 (O_1670,N_14985,N_14922);
and UO_1671 (O_1671,N_14986,N_14884);
nand UO_1672 (O_1672,N_14992,N_14927);
and UO_1673 (O_1673,N_14912,N_14950);
nand UO_1674 (O_1674,N_14953,N_14944);
nor UO_1675 (O_1675,N_14942,N_14951);
xnor UO_1676 (O_1676,N_14889,N_14979);
nand UO_1677 (O_1677,N_14882,N_14938);
nor UO_1678 (O_1678,N_14990,N_14911);
nor UO_1679 (O_1679,N_14972,N_14978);
or UO_1680 (O_1680,N_14880,N_14896);
and UO_1681 (O_1681,N_14879,N_14897);
or UO_1682 (O_1682,N_14924,N_14961);
xor UO_1683 (O_1683,N_14886,N_14952);
xnor UO_1684 (O_1684,N_14996,N_14997);
xor UO_1685 (O_1685,N_14939,N_14943);
nand UO_1686 (O_1686,N_14989,N_14893);
or UO_1687 (O_1687,N_14923,N_14925);
nand UO_1688 (O_1688,N_14995,N_14953);
nor UO_1689 (O_1689,N_14906,N_14969);
nand UO_1690 (O_1690,N_14933,N_14981);
and UO_1691 (O_1691,N_14996,N_14975);
nand UO_1692 (O_1692,N_14912,N_14937);
nand UO_1693 (O_1693,N_14999,N_14938);
or UO_1694 (O_1694,N_14893,N_14908);
nor UO_1695 (O_1695,N_14877,N_14965);
nand UO_1696 (O_1696,N_14886,N_14889);
nor UO_1697 (O_1697,N_14892,N_14967);
nand UO_1698 (O_1698,N_14932,N_14975);
xnor UO_1699 (O_1699,N_14999,N_14885);
nand UO_1700 (O_1700,N_14945,N_14994);
or UO_1701 (O_1701,N_14901,N_14996);
xor UO_1702 (O_1702,N_14911,N_14979);
nand UO_1703 (O_1703,N_14984,N_14921);
or UO_1704 (O_1704,N_14934,N_14955);
nor UO_1705 (O_1705,N_14983,N_14876);
or UO_1706 (O_1706,N_14954,N_14959);
and UO_1707 (O_1707,N_14955,N_14889);
nand UO_1708 (O_1708,N_14890,N_14989);
and UO_1709 (O_1709,N_14910,N_14957);
or UO_1710 (O_1710,N_14911,N_14938);
nor UO_1711 (O_1711,N_14950,N_14910);
xnor UO_1712 (O_1712,N_14969,N_14878);
and UO_1713 (O_1713,N_14899,N_14929);
xnor UO_1714 (O_1714,N_14889,N_14997);
nor UO_1715 (O_1715,N_14894,N_14944);
xnor UO_1716 (O_1716,N_14921,N_14971);
or UO_1717 (O_1717,N_14924,N_14960);
xnor UO_1718 (O_1718,N_14900,N_14957);
xor UO_1719 (O_1719,N_14969,N_14951);
nor UO_1720 (O_1720,N_14962,N_14886);
or UO_1721 (O_1721,N_14908,N_14919);
and UO_1722 (O_1722,N_14965,N_14954);
xnor UO_1723 (O_1723,N_14986,N_14882);
xnor UO_1724 (O_1724,N_14937,N_14950);
and UO_1725 (O_1725,N_14991,N_14995);
or UO_1726 (O_1726,N_14918,N_14958);
and UO_1727 (O_1727,N_14921,N_14926);
or UO_1728 (O_1728,N_14989,N_14897);
nor UO_1729 (O_1729,N_14958,N_14983);
nand UO_1730 (O_1730,N_14875,N_14914);
nor UO_1731 (O_1731,N_14944,N_14981);
and UO_1732 (O_1732,N_14935,N_14888);
nand UO_1733 (O_1733,N_14979,N_14935);
nor UO_1734 (O_1734,N_14968,N_14918);
nor UO_1735 (O_1735,N_14911,N_14993);
xnor UO_1736 (O_1736,N_14921,N_14904);
and UO_1737 (O_1737,N_14932,N_14936);
or UO_1738 (O_1738,N_14896,N_14898);
and UO_1739 (O_1739,N_14930,N_14992);
nand UO_1740 (O_1740,N_14988,N_14905);
or UO_1741 (O_1741,N_14917,N_14905);
xnor UO_1742 (O_1742,N_14992,N_14947);
xnor UO_1743 (O_1743,N_14964,N_14961);
or UO_1744 (O_1744,N_14930,N_14974);
or UO_1745 (O_1745,N_14969,N_14984);
xor UO_1746 (O_1746,N_14941,N_14973);
or UO_1747 (O_1747,N_14949,N_14889);
nor UO_1748 (O_1748,N_14875,N_14968);
or UO_1749 (O_1749,N_14958,N_14928);
nand UO_1750 (O_1750,N_14946,N_14941);
nor UO_1751 (O_1751,N_14918,N_14912);
or UO_1752 (O_1752,N_14918,N_14929);
and UO_1753 (O_1753,N_14913,N_14916);
or UO_1754 (O_1754,N_14899,N_14894);
and UO_1755 (O_1755,N_14907,N_14924);
and UO_1756 (O_1756,N_14908,N_14939);
nor UO_1757 (O_1757,N_14933,N_14924);
nand UO_1758 (O_1758,N_14978,N_14941);
xor UO_1759 (O_1759,N_14939,N_14984);
and UO_1760 (O_1760,N_14971,N_14963);
or UO_1761 (O_1761,N_14935,N_14895);
and UO_1762 (O_1762,N_14929,N_14958);
or UO_1763 (O_1763,N_14971,N_14905);
nand UO_1764 (O_1764,N_14964,N_14918);
and UO_1765 (O_1765,N_14967,N_14876);
nor UO_1766 (O_1766,N_14882,N_14967);
nand UO_1767 (O_1767,N_14960,N_14995);
xnor UO_1768 (O_1768,N_14883,N_14915);
xnor UO_1769 (O_1769,N_14920,N_14887);
and UO_1770 (O_1770,N_14955,N_14880);
nand UO_1771 (O_1771,N_14980,N_14879);
or UO_1772 (O_1772,N_14903,N_14986);
xor UO_1773 (O_1773,N_14978,N_14891);
and UO_1774 (O_1774,N_14965,N_14912);
nor UO_1775 (O_1775,N_14984,N_14919);
nand UO_1776 (O_1776,N_14995,N_14946);
xnor UO_1777 (O_1777,N_14992,N_14996);
nand UO_1778 (O_1778,N_14940,N_14948);
xnor UO_1779 (O_1779,N_14997,N_14942);
and UO_1780 (O_1780,N_14899,N_14880);
or UO_1781 (O_1781,N_14927,N_14937);
nor UO_1782 (O_1782,N_14948,N_14970);
or UO_1783 (O_1783,N_14897,N_14956);
nor UO_1784 (O_1784,N_14888,N_14895);
or UO_1785 (O_1785,N_14964,N_14987);
xnor UO_1786 (O_1786,N_14936,N_14875);
and UO_1787 (O_1787,N_14898,N_14929);
and UO_1788 (O_1788,N_14958,N_14980);
and UO_1789 (O_1789,N_14938,N_14937);
or UO_1790 (O_1790,N_14926,N_14890);
xor UO_1791 (O_1791,N_14950,N_14983);
or UO_1792 (O_1792,N_14949,N_14875);
or UO_1793 (O_1793,N_14994,N_14940);
nor UO_1794 (O_1794,N_14976,N_14880);
and UO_1795 (O_1795,N_14997,N_14931);
and UO_1796 (O_1796,N_14930,N_14915);
or UO_1797 (O_1797,N_14902,N_14882);
and UO_1798 (O_1798,N_14992,N_14988);
and UO_1799 (O_1799,N_14900,N_14931);
nor UO_1800 (O_1800,N_14945,N_14998);
nand UO_1801 (O_1801,N_14880,N_14993);
and UO_1802 (O_1802,N_14985,N_14957);
xnor UO_1803 (O_1803,N_14908,N_14926);
xor UO_1804 (O_1804,N_14948,N_14955);
nand UO_1805 (O_1805,N_14927,N_14952);
nand UO_1806 (O_1806,N_14994,N_14947);
nor UO_1807 (O_1807,N_14953,N_14935);
and UO_1808 (O_1808,N_14951,N_14987);
nand UO_1809 (O_1809,N_14975,N_14890);
nor UO_1810 (O_1810,N_14965,N_14935);
or UO_1811 (O_1811,N_14992,N_14949);
xnor UO_1812 (O_1812,N_14929,N_14940);
xor UO_1813 (O_1813,N_14990,N_14987);
and UO_1814 (O_1814,N_14895,N_14984);
xor UO_1815 (O_1815,N_14961,N_14963);
nor UO_1816 (O_1816,N_14886,N_14905);
xnor UO_1817 (O_1817,N_14967,N_14935);
or UO_1818 (O_1818,N_14939,N_14953);
nand UO_1819 (O_1819,N_14932,N_14952);
and UO_1820 (O_1820,N_14993,N_14917);
nand UO_1821 (O_1821,N_14998,N_14996);
xor UO_1822 (O_1822,N_14980,N_14913);
and UO_1823 (O_1823,N_14886,N_14974);
and UO_1824 (O_1824,N_14913,N_14955);
or UO_1825 (O_1825,N_14951,N_14924);
xor UO_1826 (O_1826,N_14891,N_14909);
and UO_1827 (O_1827,N_14992,N_14920);
xnor UO_1828 (O_1828,N_14927,N_14978);
nor UO_1829 (O_1829,N_14889,N_14876);
and UO_1830 (O_1830,N_14981,N_14948);
or UO_1831 (O_1831,N_14951,N_14920);
nor UO_1832 (O_1832,N_14886,N_14901);
xnor UO_1833 (O_1833,N_14931,N_14915);
or UO_1834 (O_1834,N_14892,N_14901);
or UO_1835 (O_1835,N_14944,N_14910);
xor UO_1836 (O_1836,N_14981,N_14889);
xnor UO_1837 (O_1837,N_14952,N_14965);
or UO_1838 (O_1838,N_14968,N_14955);
and UO_1839 (O_1839,N_14904,N_14989);
and UO_1840 (O_1840,N_14903,N_14992);
nor UO_1841 (O_1841,N_14979,N_14978);
xnor UO_1842 (O_1842,N_14900,N_14991);
nand UO_1843 (O_1843,N_14997,N_14962);
and UO_1844 (O_1844,N_14888,N_14996);
or UO_1845 (O_1845,N_14891,N_14925);
and UO_1846 (O_1846,N_14941,N_14999);
and UO_1847 (O_1847,N_14924,N_14900);
nand UO_1848 (O_1848,N_14925,N_14881);
xnor UO_1849 (O_1849,N_14918,N_14962);
or UO_1850 (O_1850,N_14969,N_14966);
xor UO_1851 (O_1851,N_14945,N_14946);
xnor UO_1852 (O_1852,N_14898,N_14948);
xor UO_1853 (O_1853,N_14974,N_14885);
xnor UO_1854 (O_1854,N_14900,N_14993);
or UO_1855 (O_1855,N_14981,N_14999);
xor UO_1856 (O_1856,N_14892,N_14907);
nand UO_1857 (O_1857,N_14915,N_14900);
xnor UO_1858 (O_1858,N_14909,N_14892);
nor UO_1859 (O_1859,N_14931,N_14950);
nor UO_1860 (O_1860,N_14906,N_14949);
xnor UO_1861 (O_1861,N_14960,N_14999);
nand UO_1862 (O_1862,N_14984,N_14966);
and UO_1863 (O_1863,N_14969,N_14985);
xnor UO_1864 (O_1864,N_14985,N_14981);
nor UO_1865 (O_1865,N_14886,N_14971);
xor UO_1866 (O_1866,N_14933,N_14967);
and UO_1867 (O_1867,N_14982,N_14904);
and UO_1868 (O_1868,N_14980,N_14942);
nor UO_1869 (O_1869,N_14884,N_14897);
xnor UO_1870 (O_1870,N_14976,N_14882);
or UO_1871 (O_1871,N_14962,N_14891);
xor UO_1872 (O_1872,N_14990,N_14927);
and UO_1873 (O_1873,N_14927,N_14962);
xor UO_1874 (O_1874,N_14970,N_14952);
xor UO_1875 (O_1875,N_14916,N_14917);
or UO_1876 (O_1876,N_14889,N_14990);
nand UO_1877 (O_1877,N_14909,N_14883);
and UO_1878 (O_1878,N_14934,N_14979);
or UO_1879 (O_1879,N_14986,N_14915);
or UO_1880 (O_1880,N_14987,N_14887);
nand UO_1881 (O_1881,N_14922,N_14921);
nor UO_1882 (O_1882,N_14996,N_14935);
nand UO_1883 (O_1883,N_14890,N_14980);
or UO_1884 (O_1884,N_14912,N_14951);
nand UO_1885 (O_1885,N_14956,N_14933);
or UO_1886 (O_1886,N_14986,N_14895);
nor UO_1887 (O_1887,N_14995,N_14924);
and UO_1888 (O_1888,N_14881,N_14999);
xor UO_1889 (O_1889,N_14902,N_14998);
xor UO_1890 (O_1890,N_14882,N_14946);
or UO_1891 (O_1891,N_14944,N_14961);
and UO_1892 (O_1892,N_14917,N_14948);
and UO_1893 (O_1893,N_14977,N_14913);
xnor UO_1894 (O_1894,N_14934,N_14980);
or UO_1895 (O_1895,N_14944,N_14926);
nor UO_1896 (O_1896,N_14983,N_14993);
nor UO_1897 (O_1897,N_14935,N_14902);
and UO_1898 (O_1898,N_14876,N_14974);
or UO_1899 (O_1899,N_14907,N_14933);
nor UO_1900 (O_1900,N_14949,N_14993);
or UO_1901 (O_1901,N_14875,N_14880);
xor UO_1902 (O_1902,N_14992,N_14978);
or UO_1903 (O_1903,N_14991,N_14890);
nand UO_1904 (O_1904,N_14988,N_14920);
xnor UO_1905 (O_1905,N_14925,N_14901);
xnor UO_1906 (O_1906,N_14891,N_14922);
or UO_1907 (O_1907,N_14878,N_14947);
xor UO_1908 (O_1908,N_14905,N_14938);
nor UO_1909 (O_1909,N_14988,N_14900);
nand UO_1910 (O_1910,N_14912,N_14989);
and UO_1911 (O_1911,N_14990,N_14963);
nor UO_1912 (O_1912,N_14914,N_14983);
nor UO_1913 (O_1913,N_14928,N_14934);
nor UO_1914 (O_1914,N_14997,N_14923);
nand UO_1915 (O_1915,N_14957,N_14999);
nand UO_1916 (O_1916,N_14936,N_14946);
or UO_1917 (O_1917,N_14876,N_14878);
and UO_1918 (O_1918,N_14892,N_14935);
nand UO_1919 (O_1919,N_14914,N_14879);
nand UO_1920 (O_1920,N_14990,N_14947);
xnor UO_1921 (O_1921,N_14962,N_14907);
nand UO_1922 (O_1922,N_14964,N_14940);
nor UO_1923 (O_1923,N_14887,N_14966);
and UO_1924 (O_1924,N_14939,N_14951);
or UO_1925 (O_1925,N_14876,N_14936);
nand UO_1926 (O_1926,N_14984,N_14954);
or UO_1927 (O_1927,N_14920,N_14955);
and UO_1928 (O_1928,N_14935,N_14984);
nor UO_1929 (O_1929,N_14902,N_14971);
and UO_1930 (O_1930,N_14974,N_14982);
or UO_1931 (O_1931,N_14897,N_14889);
and UO_1932 (O_1932,N_14931,N_14885);
or UO_1933 (O_1933,N_14940,N_14896);
xor UO_1934 (O_1934,N_14883,N_14924);
or UO_1935 (O_1935,N_14886,N_14966);
and UO_1936 (O_1936,N_14933,N_14922);
nor UO_1937 (O_1937,N_14903,N_14878);
and UO_1938 (O_1938,N_14989,N_14924);
nor UO_1939 (O_1939,N_14971,N_14906);
xor UO_1940 (O_1940,N_14944,N_14946);
xnor UO_1941 (O_1941,N_14943,N_14917);
nor UO_1942 (O_1942,N_14923,N_14899);
nand UO_1943 (O_1943,N_14946,N_14953);
nand UO_1944 (O_1944,N_14895,N_14921);
or UO_1945 (O_1945,N_14968,N_14985);
xnor UO_1946 (O_1946,N_14912,N_14916);
nor UO_1947 (O_1947,N_14960,N_14890);
and UO_1948 (O_1948,N_14986,N_14924);
and UO_1949 (O_1949,N_14968,N_14902);
and UO_1950 (O_1950,N_14900,N_14912);
nor UO_1951 (O_1951,N_14972,N_14953);
nor UO_1952 (O_1952,N_14898,N_14957);
xor UO_1953 (O_1953,N_14927,N_14947);
and UO_1954 (O_1954,N_14999,N_14920);
or UO_1955 (O_1955,N_14895,N_14929);
and UO_1956 (O_1956,N_14921,N_14913);
nand UO_1957 (O_1957,N_14969,N_14967);
nor UO_1958 (O_1958,N_14964,N_14920);
nand UO_1959 (O_1959,N_14905,N_14960);
nor UO_1960 (O_1960,N_14944,N_14959);
xnor UO_1961 (O_1961,N_14982,N_14971);
or UO_1962 (O_1962,N_14929,N_14988);
nor UO_1963 (O_1963,N_14876,N_14890);
xnor UO_1964 (O_1964,N_14957,N_14992);
or UO_1965 (O_1965,N_14969,N_14930);
nor UO_1966 (O_1966,N_14985,N_14875);
nor UO_1967 (O_1967,N_14927,N_14985);
xor UO_1968 (O_1968,N_14919,N_14951);
xor UO_1969 (O_1969,N_14940,N_14991);
xor UO_1970 (O_1970,N_14875,N_14963);
and UO_1971 (O_1971,N_14894,N_14931);
and UO_1972 (O_1972,N_14922,N_14966);
nand UO_1973 (O_1973,N_14936,N_14929);
or UO_1974 (O_1974,N_14931,N_14983);
nor UO_1975 (O_1975,N_14875,N_14957);
and UO_1976 (O_1976,N_14881,N_14904);
and UO_1977 (O_1977,N_14952,N_14955);
xnor UO_1978 (O_1978,N_14882,N_14972);
xor UO_1979 (O_1979,N_14957,N_14928);
and UO_1980 (O_1980,N_14895,N_14907);
nand UO_1981 (O_1981,N_14917,N_14911);
xnor UO_1982 (O_1982,N_14964,N_14891);
nor UO_1983 (O_1983,N_14950,N_14954);
xnor UO_1984 (O_1984,N_14904,N_14930);
nor UO_1985 (O_1985,N_14909,N_14974);
nand UO_1986 (O_1986,N_14992,N_14906);
xor UO_1987 (O_1987,N_14898,N_14974);
and UO_1988 (O_1988,N_14931,N_14918);
nor UO_1989 (O_1989,N_14923,N_14879);
nand UO_1990 (O_1990,N_14986,N_14939);
and UO_1991 (O_1991,N_14973,N_14885);
nand UO_1992 (O_1992,N_14903,N_14927);
nor UO_1993 (O_1993,N_14993,N_14936);
xor UO_1994 (O_1994,N_14938,N_14987);
or UO_1995 (O_1995,N_14882,N_14970);
nand UO_1996 (O_1996,N_14984,N_14982);
nor UO_1997 (O_1997,N_14961,N_14936);
and UO_1998 (O_1998,N_14990,N_14930);
and UO_1999 (O_1999,N_14988,N_14962);
endmodule