module basic_500_3000_500_3_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_335,In_298);
and U1 (N_1,In_333,In_356);
or U2 (N_2,In_80,In_191);
or U3 (N_3,In_284,In_125);
or U4 (N_4,In_343,In_468);
nor U5 (N_5,In_370,In_39);
and U6 (N_6,In_411,In_102);
and U7 (N_7,In_262,In_320);
or U8 (N_8,In_239,In_96);
nor U9 (N_9,In_364,In_62);
or U10 (N_10,In_342,In_279);
xor U11 (N_11,In_214,In_120);
or U12 (N_12,In_372,In_105);
nor U13 (N_13,In_290,In_18);
nand U14 (N_14,In_168,In_206);
nand U15 (N_15,In_166,In_440);
nand U16 (N_16,In_149,In_382);
nor U17 (N_17,In_272,In_400);
or U18 (N_18,In_365,In_115);
and U19 (N_19,In_188,In_480);
or U20 (N_20,In_455,In_375);
nand U21 (N_21,In_27,In_386);
and U22 (N_22,In_133,In_67);
nand U23 (N_23,In_453,In_371);
nor U24 (N_24,In_70,In_11);
nand U25 (N_25,In_212,In_38);
xor U26 (N_26,In_387,In_492);
xor U27 (N_27,In_286,In_267);
or U28 (N_28,In_173,In_99);
nand U29 (N_29,In_146,In_285);
or U30 (N_30,In_297,In_463);
nor U31 (N_31,In_276,In_199);
nand U32 (N_32,In_68,In_454);
xor U33 (N_33,In_295,In_402);
nor U34 (N_34,In_477,In_202);
nor U35 (N_35,In_247,In_160);
nand U36 (N_36,In_449,In_167);
and U37 (N_37,In_313,In_117);
nor U38 (N_38,In_21,In_497);
nor U39 (N_39,In_24,In_350);
nand U40 (N_40,In_434,In_479);
and U41 (N_41,In_104,In_180);
nand U42 (N_42,In_281,In_315);
and U43 (N_43,In_197,In_347);
or U44 (N_44,In_139,In_194);
nand U45 (N_45,In_491,In_140);
or U46 (N_46,In_116,In_263);
xnor U47 (N_47,In_12,In_15);
or U48 (N_48,In_78,In_69);
nand U49 (N_49,In_181,In_123);
nor U50 (N_50,In_427,In_63);
nand U51 (N_51,In_421,In_476);
xor U52 (N_52,In_448,In_470);
xor U53 (N_53,In_441,In_6);
xnor U54 (N_54,In_465,In_29);
and U55 (N_55,In_221,In_458);
or U56 (N_56,In_251,In_327);
xnor U57 (N_57,In_131,In_107);
or U58 (N_58,In_486,In_368);
nand U59 (N_59,In_236,In_494);
nand U60 (N_60,In_226,In_308);
and U61 (N_61,In_225,In_48);
xnor U62 (N_62,In_134,In_64);
nor U63 (N_63,In_363,In_159);
or U64 (N_64,In_113,In_355);
or U65 (N_65,In_437,In_446);
xnor U66 (N_66,In_360,In_178);
nand U67 (N_67,In_293,In_256);
nand U68 (N_68,In_359,In_329);
and U69 (N_69,In_229,In_302);
nor U70 (N_70,In_249,In_259);
nand U71 (N_71,In_367,In_124);
nor U72 (N_72,In_42,In_9);
nand U73 (N_73,In_144,In_274);
xnor U74 (N_74,In_300,In_143);
nand U75 (N_75,In_129,In_184);
xor U76 (N_76,In_353,In_325);
and U77 (N_77,In_424,In_459);
and U78 (N_78,In_156,In_86);
xor U79 (N_79,In_339,In_151);
nor U80 (N_80,In_106,In_378);
and U81 (N_81,In_444,In_340);
and U82 (N_82,In_472,In_310);
xnor U83 (N_83,In_224,In_161);
xor U84 (N_84,In_100,In_358);
nand U85 (N_85,In_1,In_33);
or U86 (N_86,In_436,In_257);
and U87 (N_87,In_54,In_208);
or U88 (N_88,In_255,In_130);
nor U89 (N_89,In_79,In_403);
or U90 (N_90,In_362,In_270);
or U91 (N_91,In_451,In_152);
and U92 (N_92,In_25,In_485);
xor U93 (N_93,In_176,In_243);
nor U94 (N_94,In_391,In_205);
and U95 (N_95,In_75,In_457);
xnor U96 (N_96,In_396,In_162);
or U97 (N_97,In_269,In_461);
and U98 (N_98,In_182,In_264);
nand U99 (N_99,In_85,In_307);
xor U100 (N_100,In_58,In_228);
and U101 (N_101,In_142,In_338);
xnor U102 (N_102,In_336,In_482);
nand U103 (N_103,In_471,In_488);
and U104 (N_104,In_217,In_489);
or U105 (N_105,In_397,In_433);
and U106 (N_106,In_345,In_413);
nand U107 (N_107,In_341,In_244);
nor U108 (N_108,In_108,In_373);
or U109 (N_109,In_201,In_288);
nand U110 (N_110,In_45,In_137);
or U111 (N_111,In_32,In_61);
xor U112 (N_112,In_443,In_462);
and U113 (N_113,In_369,In_204);
xor U114 (N_114,In_237,In_496);
nand U115 (N_115,In_31,In_16);
or U116 (N_116,In_381,In_393);
nand U117 (N_117,In_495,In_498);
nand U118 (N_118,In_410,In_73);
xor U119 (N_119,In_445,In_154);
nor U120 (N_120,In_493,In_44);
or U121 (N_121,In_261,In_322);
nand U122 (N_122,In_87,In_55);
xnor U123 (N_123,In_401,In_211);
xor U124 (N_124,In_442,In_50);
and U125 (N_125,In_289,In_303);
nor U126 (N_126,In_409,In_392);
nand U127 (N_127,In_394,In_474);
or U128 (N_128,In_98,In_379);
xor U129 (N_129,In_59,In_291);
xor U130 (N_130,In_323,In_418);
or U131 (N_131,In_28,In_245);
xor U132 (N_132,In_95,In_384);
and U133 (N_133,In_428,In_405);
xnor U134 (N_134,In_385,In_109);
or U135 (N_135,In_121,In_450);
or U136 (N_136,In_216,In_135);
or U137 (N_137,In_57,In_438);
and U138 (N_138,In_304,In_20);
and U139 (N_139,In_399,In_432);
nor U140 (N_140,In_114,In_253);
xor U141 (N_141,In_469,In_155);
and U142 (N_142,In_83,In_84);
or U143 (N_143,In_17,In_53);
or U144 (N_144,In_318,In_74);
xor U145 (N_145,In_334,In_157);
xor U146 (N_146,In_346,In_447);
nand U147 (N_147,In_150,In_41);
xor U148 (N_148,In_314,In_223);
or U149 (N_149,In_337,In_52);
or U150 (N_150,In_282,In_275);
or U151 (N_151,In_317,In_219);
nand U152 (N_152,In_273,In_250);
nand U153 (N_153,In_435,In_296);
and U154 (N_154,In_490,In_390);
nor U155 (N_155,In_283,In_254);
and U156 (N_156,In_40,In_158);
nand U157 (N_157,In_8,In_252);
nand U158 (N_158,In_127,In_89);
or U159 (N_159,In_136,In_278);
nand U160 (N_160,In_326,In_90);
and U161 (N_161,In_431,In_311);
and U162 (N_162,In_148,In_404);
nor U163 (N_163,In_215,In_195);
and U164 (N_164,In_280,In_380);
xnor U165 (N_165,In_232,In_88);
xor U166 (N_166,In_110,In_321);
and U167 (N_167,In_316,In_287);
or U168 (N_168,In_171,In_141);
and U169 (N_169,In_51,In_357);
xnor U170 (N_170,In_13,In_344);
and U171 (N_171,In_101,In_60);
xor U172 (N_172,In_126,In_30);
nand U173 (N_173,In_260,In_354);
nand U174 (N_174,In_305,In_376);
or U175 (N_175,In_266,In_153);
xnor U176 (N_176,In_77,In_189);
or U177 (N_177,In_456,In_499);
nand U178 (N_178,In_242,In_420);
or U179 (N_179,In_193,In_395);
or U180 (N_180,In_198,In_72);
and U181 (N_181,In_233,In_332);
and U182 (N_182,In_473,In_309);
or U183 (N_183,In_3,In_430);
or U184 (N_184,In_349,In_377);
and U185 (N_185,In_200,In_423);
nand U186 (N_186,In_147,In_172);
nor U187 (N_187,In_294,In_118);
xor U188 (N_188,In_122,In_5);
and U189 (N_189,In_111,In_170);
nand U190 (N_190,In_460,In_163);
xnor U191 (N_191,In_234,In_426);
or U192 (N_192,In_227,In_132);
nor U193 (N_193,In_419,In_478);
xnor U194 (N_194,In_422,In_417);
nor U195 (N_195,In_467,In_91);
nand U196 (N_196,In_128,In_203);
xor U197 (N_197,In_220,In_22);
nand U198 (N_198,In_165,In_174);
xnor U199 (N_199,In_92,In_240);
and U200 (N_200,In_425,In_383);
nand U201 (N_201,In_277,In_175);
and U202 (N_202,In_408,In_265);
xor U203 (N_203,In_268,In_179);
or U204 (N_204,In_483,In_312);
or U205 (N_205,In_439,In_352);
nand U206 (N_206,In_93,In_112);
nor U207 (N_207,In_164,In_415);
or U208 (N_208,In_10,In_196);
nor U209 (N_209,In_429,In_319);
and U210 (N_210,In_388,In_7);
xnor U211 (N_211,In_481,In_119);
and U212 (N_212,In_487,In_389);
nor U213 (N_213,In_475,In_76);
nor U214 (N_214,In_218,In_0);
nor U215 (N_215,In_97,In_37);
or U216 (N_216,In_26,In_398);
nor U217 (N_217,In_258,In_49);
nand U218 (N_218,In_412,In_464);
nor U219 (N_219,In_330,In_222);
or U220 (N_220,In_2,In_81);
or U221 (N_221,In_94,In_71);
and U222 (N_222,In_169,In_187);
nand U223 (N_223,In_452,In_65);
or U224 (N_224,In_331,In_248);
nor U225 (N_225,In_190,In_66);
nand U226 (N_226,In_348,In_484);
nand U227 (N_227,In_235,In_407);
nor U228 (N_228,In_466,In_238);
nor U229 (N_229,In_246,In_23);
xor U230 (N_230,In_406,In_324);
nor U231 (N_231,In_4,In_292);
nand U232 (N_232,In_416,In_192);
nor U233 (N_233,In_230,In_271);
or U234 (N_234,In_14,In_82);
xor U235 (N_235,In_328,In_306);
or U236 (N_236,In_46,In_301);
xnor U237 (N_237,In_374,In_231);
nand U238 (N_238,In_366,In_299);
or U239 (N_239,In_145,In_177);
or U240 (N_240,In_103,In_361);
or U241 (N_241,In_19,In_185);
nand U242 (N_242,In_47,In_209);
nor U243 (N_243,In_56,In_34);
nor U244 (N_244,In_43,In_414);
and U245 (N_245,In_35,In_207);
nor U246 (N_246,In_138,In_241);
nand U247 (N_247,In_183,In_36);
or U248 (N_248,In_186,In_351);
xor U249 (N_249,In_210,In_213);
nand U250 (N_250,In_11,In_310);
xor U251 (N_251,In_324,In_81);
nand U252 (N_252,In_185,In_199);
nand U253 (N_253,In_10,In_409);
nand U254 (N_254,In_318,In_264);
xnor U255 (N_255,In_198,In_399);
xor U256 (N_256,In_160,In_297);
and U257 (N_257,In_150,In_471);
nand U258 (N_258,In_440,In_12);
and U259 (N_259,In_369,In_77);
xnor U260 (N_260,In_136,In_271);
nand U261 (N_261,In_440,In_113);
nand U262 (N_262,In_258,In_465);
nor U263 (N_263,In_99,In_183);
and U264 (N_264,In_487,In_345);
or U265 (N_265,In_156,In_293);
nor U266 (N_266,In_253,In_475);
nand U267 (N_267,In_496,In_38);
nor U268 (N_268,In_195,In_384);
xor U269 (N_269,In_70,In_41);
nor U270 (N_270,In_350,In_16);
or U271 (N_271,In_51,In_91);
or U272 (N_272,In_294,In_361);
xor U273 (N_273,In_359,In_325);
and U274 (N_274,In_108,In_327);
or U275 (N_275,In_132,In_163);
nand U276 (N_276,In_50,In_78);
or U277 (N_277,In_326,In_273);
or U278 (N_278,In_360,In_291);
nand U279 (N_279,In_251,In_148);
nand U280 (N_280,In_488,In_148);
nand U281 (N_281,In_179,In_413);
xor U282 (N_282,In_107,In_113);
nor U283 (N_283,In_297,In_373);
xnor U284 (N_284,In_82,In_305);
nor U285 (N_285,In_161,In_45);
nor U286 (N_286,In_432,In_341);
xor U287 (N_287,In_227,In_432);
or U288 (N_288,In_223,In_34);
nor U289 (N_289,In_422,In_231);
and U290 (N_290,In_265,In_475);
nand U291 (N_291,In_430,In_378);
nor U292 (N_292,In_317,In_160);
nor U293 (N_293,In_136,In_361);
xor U294 (N_294,In_177,In_373);
xnor U295 (N_295,In_192,In_196);
and U296 (N_296,In_379,In_92);
xnor U297 (N_297,In_174,In_78);
and U298 (N_298,In_337,In_357);
or U299 (N_299,In_183,In_341);
nand U300 (N_300,In_166,In_141);
or U301 (N_301,In_276,In_408);
and U302 (N_302,In_72,In_137);
nand U303 (N_303,In_361,In_259);
xnor U304 (N_304,In_132,In_307);
xnor U305 (N_305,In_433,In_352);
and U306 (N_306,In_413,In_279);
nor U307 (N_307,In_128,In_428);
or U308 (N_308,In_62,In_111);
nor U309 (N_309,In_175,In_74);
and U310 (N_310,In_65,In_457);
or U311 (N_311,In_70,In_216);
and U312 (N_312,In_86,In_407);
xnor U313 (N_313,In_27,In_156);
nand U314 (N_314,In_6,In_336);
xor U315 (N_315,In_286,In_270);
and U316 (N_316,In_170,In_196);
nor U317 (N_317,In_337,In_348);
or U318 (N_318,In_402,In_26);
and U319 (N_319,In_419,In_407);
nand U320 (N_320,In_413,In_273);
nand U321 (N_321,In_111,In_302);
and U322 (N_322,In_229,In_232);
nor U323 (N_323,In_468,In_345);
xnor U324 (N_324,In_109,In_111);
nand U325 (N_325,In_139,In_310);
and U326 (N_326,In_363,In_430);
nor U327 (N_327,In_464,In_295);
xor U328 (N_328,In_229,In_388);
and U329 (N_329,In_452,In_220);
nand U330 (N_330,In_238,In_25);
or U331 (N_331,In_119,In_193);
nor U332 (N_332,In_22,In_167);
nand U333 (N_333,In_351,In_429);
nor U334 (N_334,In_77,In_402);
xor U335 (N_335,In_438,In_171);
and U336 (N_336,In_425,In_459);
nand U337 (N_337,In_499,In_396);
nand U338 (N_338,In_26,In_211);
nand U339 (N_339,In_409,In_264);
or U340 (N_340,In_296,In_8);
nand U341 (N_341,In_282,In_238);
nor U342 (N_342,In_245,In_120);
nor U343 (N_343,In_113,In_124);
nand U344 (N_344,In_204,In_264);
nand U345 (N_345,In_375,In_339);
nor U346 (N_346,In_91,In_84);
xor U347 (N_347,In_373,In_399);
or U348 (N_348,In_104,In_222);
nor U349 (N_349,In_87,In_415);
nand U350 (N_350,In_255,In_258);
nand U351 (N_351,In_310,In_13);
nor U352 (N_352,In_247,In_103);
nand U353 (N_353,In_426,In_469);
nand U354 (N_354,In_293,In_183);
xor U355 (N_355,In_54,In_337);
nand U356 (N_356,In_463,In_261);
nand U357 (N_357,In_247,In_147);
nor U358 (N_358,In_281,In_265);
nand U359 (N_359,In_240,In_147);
nor U360 (N_360,In_373,In_294);
or U361 (N_361,In_172,In_465);
or U362 (N_362,In_236,In_68);
xor U363 (N_363,In_334,In_247);
or U364 (N_364,In_344,In_394);
or U365 (N_365,In_128,In_365);
and U366 (N_366,In_64,In_236);
and U367 (N_367,In_97,In_69);
or U368 (N_368,In_328,In_329);
xor U369 (N_369,In_423,In_72);
and U370 (N_370,In_101,In_273);
nor U371 (N_371,In_291,In_286);
xnor U372 (N_372,In_201,In_379);
nand U373 (N_373,In_377,In_179);
nor U374 (N_374,In_12,In_476);
nand U375 (N_375,In_353,In_367);
nor U376 (N_376,In_406,In_263);
nand U377 (N_377,In_395,In_43);
nand U378 (N_378,In_211,In_430);
nand U379 (N_379,In_39,In_105);
nor U380 (N_380,In_276,In_58);
and U381 (N_381,In_86,In_122);
nor U382 (N_382,In_21,In_153);
or U383 (N_383,In_403,In_195);
nand U384 (N_384,In_334,In_470);
nand U385 (N_385,In_162,In_253);
or U386 (N_386,In_175,In_309);
nor U387 (N_387,In_376,In_7);
xnor U388 (N_388,In_68,In_155);
and U389 (N_389,In_62,In_127);
or U390 (N_390,In_363,In_406);
nand U391 (N_391,In_39,In_374);
xor U392 (N_392,In_62,In_492);
xnor U393 (N_393,In_62,In_164);
and U394 (N_394,In_128,In_90);
or U395 (N_395,In_24,In_144);
or U396 (N_396,In_426,In_61);
nand U397 (N_397,In_230,In_386);
and U398 (N_398,In_277,In_302);
nor U399 (N_399,In_21,In_114);
nand U400 (N_400,In_428,In_369);
or U401 (N_401,In_460,In_173);
or U402 (N_402,In_206,In_401);
nor U403 (N_403,In_240,In_280);
nor U404 (N_404,In_432,In_433);
xor U405 (N_405,In_59,In_362);
and U406 (N_406,In_45,In_104);
nand U407 (N_407,In_105,In_362);
and U408 (N_408,In_21,In_398);
and U409 (N_409,In_156,In_232);
xor U410 (N_410,In_177,In_287);
and U411 (N_411,In_104,In_340);
xnor U412 (N_412,In_325,In_249);
nor U413 (N_413,In_363,In_377);
nand U414 (N_414,In_203,In_468);
and U415 (N_415,In_81,In_326);
or U416 (N_416,In_413,In_288);
xor U417 (N_417,In_122,In_422);
nand U418 (N_418,In_442,In_268);
or U419 (N_419,In_444,In_156);
or U420 (N_420,In_228,In_463);
nand U421 (N_421,In_449,In_23);
nor U422 (N_422,In_488,In_318);
and U423 (N_423,In_338,In_192);
nand U424 (N_424,In_101,In_478);
nand U425 (N_425,In_313,In_141);
or U426 (N_426,In_250,In_56);
nand U427 (N_427,In_79,In_341);
nand U428 (N_428,In_395,In_192);
and U429 (N_429,In_143,In_14);
nand U430 (N_430,In_123,In_26);
nor U431 (N_431,In_71,In_364);
nor U432 (N_432,In_316,In_308);
xnor U433 (N_433,In_90,In_230);
nand U434 (N_434,In_205,In_490);
and U435 (N_435,In_157,In_229);
nand U436 (N_436,In_158,In_455);
xor U437 (N_437,In_141,In_15);
or U438 (N_438,In_293,In_240);
xnor U439 (N_439,In_142,In_143);
and U440 (N_440,In_472,In_118);
nor U441 (N_441,In_349,In_222);
nor U442 (N_442,In_143,In_200);
or U443 (N_443,In_136,In_171);
or U444 (N_444,In_67,In_326);
nor U445 (N_445,In_70,In_496);
and U446 (N_446,In_236,In_184);
nand U447 (N_447,In_369,In_419);
and U448 (N_448,In_245,In_451);
and U449 (N_449,In_322,In_42);
nor U450 (N_450,In_304,In_224);
nand U451 (N_451,In_465,In_355);
and U452 (N_452,In_454,In_498);
nand U453 (N_453,In_440,In_219);
nand U454 (N_454,In_480,In_436);
or U455 (N_455,In_456,In_67);
xor U456 (N_456,In_471,In_194);
nor U457 (N_457,In_275,In_211);
nand U458 (N_458,In_31,In_356);
nand U459 (N_459,In_365,In_82);
xor U460 (N_460,In_207,In_56);
and U461 (N_461,In_289,In_86);
and U462 (N_462,In_327,In_328);
xnor U463 (N_463,In_403,In_432);
or U464 (N_464,In_155,In_332);
and U465 (N_465,In_225,In_162);
nand U466 (N_466,In_383,In_18);
nor U467 (N_467,In_340,In_12);
nor U468 (N_468,In_173,In_158);
or U469 (N_469,In_300,In_448);
or U470 (N_470,In_27,In_90);
and U471 (N_471,In_15,In_262);
nand U472 (N_472,In_165,In_373);
or U473 (N_473,In_468,In_91);
nor U474 (N_474,In_263,In_472);
nor U475 (N_475,In_90,In_337);
nand U476 (N_476,In_209,In_136);
xnor U477 (N_477,In_112,In_12);
nor U478 (N_478,In_241,In_398);
or U479 (N_479,In_332,In_107);
nor U480 (N_480,In_406,In_137);
and U481 (N_481,In_428,In_233);
nor U482 (N_482,In_177,In_397);
xor U483 (N_483,In_183,In_360);
and U484 (N_484,In_459,In_60);
nor U485 (N_485,In_149,In_250);
nand U486 (N_486,In_424,In_148);
or U487 (N_487,In_164,In_281);
nor U488 (N_488,In_396,In_146);
and U489 (N_489,In_285,In_37);
nor U490 (N_490,In_151,In_288);
and U491 (N_491,In_470,In_202);
nand U492 (N_492,In_433,In_116);
nand U493 (N_493,In_263,In_180);
and U494 (N_494,In_414,In_377);
nor U495 (N_495,In_72,In_499);
and U496 (N_496,In_450,In_255);
nand U497 (N_497,In_44,In_146);
and U498 (N_498,In_104,In_267);
or U499 (N_499,In_342,In_129);
xnor U500 (N_500,In_209,In_12);
nand U501 (N_501,In_443,In_340);
or U502 (N_502,In_282,In_412);
nand U503 (N_503,In_352,In_399);
nand U504 (N_504,In_296,In_37);
nand U505 (N_505,In_65,In_146);
nor U506 (N_506,In_35,In_173);
and U507 (N_507,In_306,In_122);
and U508 (N_508,In_234,In_97);
nand U509 (N_509,In_328,In_366);
or U510 (N_510,In_343,In_300);
xnor U511 (N_511,In_479,In_388);
xnor U512 (N_512,In_210,In_270);
and U513 (N_513,In_131,In_395);
and U514 (N_514,In_380,In_401);
nor U515 (N_515,In_359,In_298);
and U516 (N_516,In_53,In_372);
and U517 (N_517,In_303,In_200);
nand U518 (N_518,In_304,In_80);
nor U519 (N_519,In_389,In_420);
or U520 (N_520,In_420,In_97);
xor U521 (N_521,In_487,In_451);
nand U522 (N_522,In_450,In_34);
xnor U523 (N_523,In_83,In_64);
nand U524 (N_524,In_156,In_278);
xor U525 (N_525,In_178,In_210);
nand U526 (N_526,In_138,In_109);
or U527 (N_527,In_213,In_197);
nor U528 (N_528,In_273,In_313);
and U529 (N_529,In_364,In_394);
xor U530 (N_530,In_134,In_26);
xor U531 (N_531,In_325,In_87);
and U532 (N_532,In_364,In_145);
nor U533 (N_533,In_283,In_410);
nor U534 (N_534,In_416,In_385);
nand U535 (N_535,In_60,In_69);
nand U536 (N_536,In_463,In_153);
or U537 (N_537,In_483,In_424);
nand U538 (N_538,In_431,In_283);
nand U539 (N_539,In_198,In_220);
nand U540 (N_540,In_178,In_388);
nand U541 (N_541,In_163,In_453);
xnor U542 (N_542,In_344,In_105);
and U543 (N_543,In_26,In_72);
nor U544 (N_544,In_358,In_172);
nor U545 (N_545,In_411,In_384);
and U546 (N_546,In_19,In_482);
and U547 (N_547,In_195,In_114);
xor U548 (N_548,In_260,In_226);
xnor U549 (N_549,In_409,In_413);
nor U550 (N_550,In_309,In_450);
nand U551 (N_551,In_0,In_11);
and U552 (N_552,In_42,In_252);
nand U553 (N_553,In_182,In_475);
nand U554 (N_554,In_36,In_48);
nand U555 (N_555,In_111,In_358);
and U556 (N_556,In_340,In_269);
xor U557 (N_557,In_64,In_308);
and U558 (N_558,In_371,In_221);
nor U559 (N_559,In_471,In_327);
xnor U560 (N_560,In_143,In_195);
and U561 (N_561,In_380,In_29);
or U562 (N_562,In_16,In_464);
and U563 (N_563,In_160,In_461);
nor U564 (N_564,In_217,In_41);
or U565 (N_565,In_234,In_410);
nor U566 (N_566,In_254,In_133);
xor U567 (N_567,In_146,In_297);
nand U568 (N_568,In_447,In_405);
nor U569 (N_569,In_462,In_403);
nand U570 (N_570,In_243,In_151);
or U571 (N_571,In_305,In_363);
nor U572 (N_572,In_354,In_163);
xnor U573 (N_573,In_217,In_73);
and U574 (N_574,In_256,In_387);
nand U575 (N_575,In_43,In_99);
xor U576 (N_576,In_283,In_273);
nor U577 (N_577,In_252,In_174);
or U578 (N_578,In_198,In_339);
nand U579 (N_579,In_13,In_271);
xnor U580 (N_580,In_413,In_219);
nor U581 (N_581,In_348,In_163);
or U582 (N_582,In_136,In_472);
xor U583 (N_583,In_286,In_442);
nor U584 (N_584,In_155,In_203);
nor U585 (N_585,In_222,In_300);
nor U586 (N_586,In_173,In_315);
nor U587 (N_587,In_464,In_151);
nor U588 (N_588,In_309,In_413);
xor U589 (N_589,In_240,In_23);
and U590 (N_590,In_297,In_382);
nand U591 (N_591,In_495,In_473);
nand U592 (N_592,In_212,In_483);
or U593 (N_593,In_215,In_18);
xor U594 (N_594,In_226,In_486);
or U595 (N_595,In_129,In_51);
or U596 (N_596,In_463,In_421);
and U597 (N_597,In_455,In_190);
and U598 (N_598,In_21,In_265);
nor U599 (N_599,In_423,In_271);
or U600 (N_600,In_338,In_44);
xnor U601 (N_601,In_182,In_13);
xor U602 (N_602,In_260,In_321);
xor U603 (N_603,In_449,In_276);
or U604 (N_604,In_23,In_337);
xor U605 (N_605,In_10,In_163);
nor U606 (N_606,In_61,In_270);
and U607 (N_607,In_439,In_359);
xnor U608 (N_608,In_32,In_142);
nand U609 (N_609,In_284,In_357);
or U610 (N_610,In_490,In_285);
xor U611 (N_611,In_200,In_408);
xor U612 (N_612,In_298,In_313);
and U613 (N_613,In_192,In_75);
and U614 (N_614,In_106,In_495);
nor U615 (N_615,In_145,In_31);
xnor U616 (N_616,In_180,In_220);
nand U617 (N_617,In_480,In_311);
or U618 (N_618,In_368,In_149);
or U619 (N_619,In_216,In_492);
xnor U620 (N_620,In_90,In_356);
or U621 (N_621,In_432,In_353);
nand U622 (N_622,In_307,In_152);
or U623 (N_623,In_165,In_253);
nor U624 (N_624,In_28,In_330);
or U625 (N_625,In_443,In_85);
or U626 (N_626,In_267,In_15);
nand U627 (N_627,In_423,In_341);
xor U628 (N_628,In_148,In_320);
and U629 (N_629,In_233,In_373);
xor U630 (N_630,In_350,In_91);
nor U631 (N_631,In_418,In_335);
and U632 (N_632,In_108,In_266);
nor U633 (N_633,In_150,In_400);
xor U634 (N_634,In_32,In_429);
or U635 (N_635,In_198,In_272);
nor U636 (N_636,In_336,In_407);
nand U637 (N_637,In_198,In_346);
nand U638 (N_638,In_85,In_211);
nor U639 (N_639,In_490,In_325);
xor U640 (N_640,In_334,In_84);
or U641 (N_641,In_179,In_354);
or U642 (N_642,In_337,In_181);
nand U643 (N_643,In_3,In_444);
xnor U644 (N_644,In_263,In_330);
nand U645 (N_645,In_282,In_449);
nand U646 (N_646,In_207,In_90);
or U647 (N_647,In_364,In_321);
nand U648 (N_648,In_72,In_307);
or U649 (N_649,In_80,In_182);
nand U650 (N_650,In_87,In_267);
xor U651 (N_651,In_322,In_204);
and U652 (N_652,In_340,In_409);
and U653 (N_653,In_171,In_123);
xnor U654 (N_654,In_15,In_8);
nor U655 (N_655,In_282,In_130);
or U656 (N_656,In_202,In_290);
nand U657 (N_657,In_477,In_65);
nor U658 (N_658,In_138,In_51);
nand U659 (N_659,In_333,In_414);
and U660 (N_660,In_490,In_249);
or U661 (N_661,In_444,In_24);
or U662 (N_662,In_61,In_443);
xor U663 (N_663,In_488,In_212);
nor U664 (N_664,In_293,In_371);
nand U665 (N_665,In_408,In_363);
xnor U666 (N_666,In_183,In_161);
xnor U667 (N_667,In_165,In_374);
nor U668 (N_668,In_27,In_119);
nor U669 (N_669,In_271,In_462);
or U670 (N_670,In_321,In_381);
nor U671 (N_671,In_383,In_353);
xnor U672 (N_672,In_224,In_464);
or U673 (N_673,In_487,In_393);
xnor U674 (N_674,In_255,In_191);
nand U675 (N_675,In_419,In_463);
xnor U676 (N_676,In_179,In_132);
and U677 (N_677,In_286,In_435);
xor U678 (N_678,In_230,In_289);
or U679 (N_679,In_483,In_325);
nand U680 (N_680,In_192,In_354);
or U681 (N_681,In_386,In_22);
or U682 (N_682,In_426,In_161);
or U683 (N_683,In_431,In_479);
xnor U684 (N_684,In_275,In_249);
nor U685 (N_685,In_420,In_255);
and U686 (N_686,In_154,In_485);
nand U687 (N_687,In_219,In_324);
xnor U688 (N_688,In_7,In_464);
or U689 (N_689,In_231,In_460);
or U690 (N_690,In_24,In_193);
nor U691 (N_691,In_427,In_202);
and U692 (N_692,In_438,In_440);
or U693 (N_693,In_209,In_121);
nand U694 (N_694,In_60,In_461);
and U695 (N_695,In_242,In_75);
nor U696 (N_696,In_70,In_74);
and U697 (N_697,In_106,In_192);
nor U698 (N_698,In_64,In_144);
and U699 (N_699,In_163,In_155);
xor U700 (N_700,In_165,In_351);
and U701 (N_701,In_273,In_302);
xnor U702 (N_702,In_291,In_104);
xor U703 (N_703,In_58,In_167);
nand U704 (N_704,In_66,In_288);
nand U705 (N_705,In_200,In_233);
and U706 (N_706,In_109,In_291);
nor U707 (N_707,In_266,In_230);
and U708 (N_708,In_478,In_384);
and U709 (N_709,In_464,In_175);
nand U710 (N_710,In_338,In_344);
xor U711 (N_711,In_97,In_211);
nor U712 (N_712,In_22,In_322);
nor U713 (N_713,In_395,In_22);
and U714 (N_714,In_379,In_43);
nand U715 (N_715,In_69,In_434);
nor U716 (N_716,In_119,In_174);
nand U717 (N_717,In_400,In_35);
nor U718 (N_718,In_450,In_264);
xnor U719 (N_719,In_232,In_407);
or U720 (N_720,In_194,In_359);
nand U721 (N_721,In_126,In_430);
nor U722 (N_722,In_197,In_282);
xnor U723 (N_723,In_421,In_388);
or U724 (N_724,In_384,In_464);
or U725 (N_725,In_45,In_483);
nand U726 (N_726,In_211,In_182);
nand U727 (N_727,In_246,In_124);
nor U728 (N_728,In_190,In_406);
nand U729 (N_729,In_454,In_117);
and U730 (N_730,In_25,In_75);
xor U731 (N_731,In_334,In_413);
xnor U732 (N_732,In_418,In_242);
nor U733 (N_733,In_121,In_406);
or U734 (N_734,In_30,In_353);
or U735 (N_735,In_406,In_177);
and U736 (N_736,In_416,In_97);
and U737 (N_737,In_414,In_297);
or U738 (N_738,In_412,In_99);
xnor U739 (N_739,In_233,In_102);
and U740 (N_740,In_497,In_409);
and U741 (N_741,In_390,In_320);
nand U742 (N_742,In_160,In_48);
nor U743 (N_743,In_379,In_480);
nand U744 (N_744,In_483,In_458);
nand U745 (N_745,In_486,In_117);
nor U746 (N_746,In_241,In_450);
nand U747 (N_747,In_9,In_129);
and U748 (N_748,In_367,In_462);
or U749 (N_749,In_67,In_404);
or U750 (N_750,In_85,In_13);
and U751 (N_751,In_132,In_15);
nand U752 (N_752,In_242,In_190);
and U753 (N_753,In_458,In_355);
xor U754 (N_754,In_427,In_333);
nand U755 (N_755,In_169,In_238);
nand U756 (N_756,In_64,In_429);
nand U757 (N_757,In_462,In_299);
nand U758 (N_758,In_415,In_66);
and U759 (N_759,In_419,In_345);
and U760 (N_760,In_169,In_417);
and U761 (N_761,In_441,In_94);
xnor U762 (N_762,In_435,In_189);
xor U763 (N_763,In_401,In_442);
nor U764 (N_764,In_202,In_281);
or U765 (N_765,In_187,In_478);
nor U766 (N_766,In_70,In_29);
xnor U767 (N_767,In_243,In_50);
and U768 (N_768,In_299,In_336);
and U769 (N_769,In_175,In_449);
nand U770 (N_770,In_168,In_459);
xor U771 (N_771,In_173,In_265);
and U772 (N_772,In_435,In_323);
nand U773 (N_773,In_100,In_257);
nor U774 (N_774,In_460,In_232);
or U775 (N_775,In_215,In_361);
or U776 (N_776,In_253,In_415);
or U777 (N_777,In_130,In_223);
xnor U778 (N_778,In_399,In_467);
nor U779 (N_779,In_484,In_489);
or U780 (N_780,In_188,In_125);
or U781 (N_781,In_131,In_345);
xnor U782 (N_782,In_325,In_329);
nand U783 (N_783,In_232,In_451);
and U784 (N_784,In_415,In_441);
and U785 (N_785,In_437,In_85);
and U786 (N_786,In_154,In_360);
xor U787 (N_787,In_251,In_20);
nand U788 (N_788,In_408,In_329);
nor U789 (N_789,In_12,In_365);
or U790 (N_790,In_68,In_190);
xnor U791 (N_791,In_484,In_185);
and U792 (N_792,In_44,In_300);
xnor U793 (N_793,In_216,In_315);
or U794 (N_794,In_136,In_459);
xor U795 (N_795,In_316,In_493);
xnor U796 (N_796,In_140,In_434);
xor U797 (N_797,In_341,In_415);
xnor U798 (N_798,In_283,In_55);
nand U799 (N_799,In_428,In_214);
and U800 (N_800,In_8,In_308);
xnor U801 (N_801,In_128,In_143);
nor U802 (N_802,In_353,In_318);
or U803 (N_803,In_9,In_463);
and U804 (N_804,In_224,In_330);
xnor U805 (N_805,In_299,In_189);
or U806 (N_806,In_456,In_312);
or U807 (N_807,In_242,In_494);
and U808 (N_808,In_477,In_81);
nor U809 (N_809,In_426,In_327);
xor U810 (N_810,In_208,In_238);
or U811 (N_811,In_404,In_177);
and U812 (N_812,In_223,In_242);
nor U813 (N_813,In_448,In_489);
xnor U814 (N_814,In_198,In_147);
nand U815 (N_815,In_289,In_71);
and U816 (N_816,In_445,In_56);
nor U817 (N_817,In_399,In_171);
nor U818 (N_818,In_155,In_110);
nand U819 (N_819,In_301,In_399);
and U820 (N_820,In_385,In_319);
nand U821 (N_821,In_103,In_443);
or U822 (N_822,In_321,In_236);
and U823 (N_823,In_348,In_260);
nor U824 (N_824,In_462,In_445);
nor U825 (N_825,In_27,In_495);
xor U826 (N_826,In_325,In_182);
xor U827 (N_827,In_342,In_376);
xor U828 (N_828,In_310,In_413);
and U829 (N_829,In_232,In_189);
nand U830 (N_830,In_216,In_409);
xnor U831 (N_831,In_327,In_81);
and U832 (N_832,In_478,In_150);
and U833 (N_833,In_452,In_419);
and U834 (N_834,In_271,In_115);
and U835 (N_835,In_57,In_99);
xor U836 (N_836,In_473,In_228);
and U837 (N_837,In_33,In_220);
xnor U838 (N_838,In_94,In_474);
and U839 (N_839,In_305,In_57);
xnor U840 (N_840,In_93,In_65);
nor U841 (N_841,In_94,In_228);
and U842 (N_842,In_148,In_95);
nand U843 (N_843,In_352,In_4);
and U844 (N_844,In_178,In_84);
xnor U845 (N_845,In_301,In_471);
and U846 (N_846,In_470,In_153);
nand U847 (N_847,In_251,In_272);
or U848 (N_848,In_287,In_123);
nand U849 (N_849,In_179,In_407);
nand U850 (N_850,In_162,In_391);
xor U851 (N_851,In_9,In_124);
nor U852 (N_852,In_140,In_249);
and U853 (N_853,In_246,In_21);
and U854 (N_854,In_405,In_195);
and U855 (N_855,In_408,In_165);
or U856 (N_856,In_219,In_116);
or U857 (N_857,In_112,In_62);
nor U858 (N_858,In_72,In_278);
nor U859 (N_859,In_351,In_436);
or U860 (N_860,In_383,In_340);
or U861 (N_861,In_28,In_441);
or U862 (N_862,In_111,In_402);
xor U863 (N_863,In_396,In_97);
and U864 (N_864,In_256,In_445);
xor U865 (N_865,In_391,In_80);
nor U866 (N_866,In_104,In_288);
or U867 (N_867,In_59,In_97);
xnor U868 (N_868,In_467,In_221);
or U869 (N_869,In_421,In_446);
xnor U870 (N_870,In_101,In_371);
and U871 (N_871,In_155,In_465);
and U872 (N_872,In_1,In_74);
nand U873 (N_873,In_323,In_249);
nand U874 (N_874,In_392,In_198);
or U875 (N_875,In_476,In_456);
and U876 (N_876,In_281,In_181);
xnor U877 (N_877,In_134,In_201);
xor U878 (N_878,In_6,In_462);
and U879 (N_879,In_476,In_466);
nand U880 (N_880,In_42,In_107);
or U881 (N_881,In_329,In_255);
or U882 (N_882,In_100,In_18);
nand U883 (N_883,In_108,In_1);
or U884 (N_884,In_242,In_439);
nor U885 (N_885,In_231,In_51);
xnor U886 (N_886,In_249,In_169);
nor U887 (N_887,In_299,In_286);
xnor U888 (N_888,In_41,In_130);
nor U889 (N_889,In_241,In_81);
and U890 (N_890,In_9,In_96);
xor U891 (N_891,In_417,In_324);
nor U892 (N_892,In_239,In_398);
xor U893 (N_893,In_91,In_8);
nor U894 (N_894,In_485,In_162);
or U895 (N_895,In_402,In_280);
or U896 (N_896,In_233,In_473);
nand U897 (N_897,In_37,In_3);
nand U898 (N_898,In_46,In_337);
nand U899 (N_899,In_327,In_184);
nor U900 (N_900,In_214,In_212);
nor U901 (N_901,In_58,In_113);
nand U902 (N_902,In_235,In_470);
nand U903 (N_903,In_53,In_370);
or U904 (N_904,In_5,In_368);
xnor U905 (N_905,In_210,In_418);
xor U906 (N_906,In_336,In_210);
or U907 (N_907,In_417,In_185);
and U908 (N_908,In_309,In_335);
nand U909 (N_909,In_149,In_422);
xnor U910 (N_910,In_454,In_343);
nand U911 (N_911,In_88,In_48);
and U912 (N_912,In_468,In_421);
nor U913 (N_913,In_301,In_69);
nor U914 (N_914,In_267,In_316);
nor U915 (N_915,In_492,In_1);
xnor U916 (N_916,In_471,In_207);
nor U917 (N_917,In_272,In_403);
nor U918 (N_918,In_294,In_286);
nand U919 (N_919,In_200,In_228);
and U920 (N_920,In_268,In_160);
and U921 (N_921,In_336,In_394);
nor U922 (N_922,In_316,In_496);
and U923 (N_923,In_113,In_20);
and U924 (N_924,In_477,In_208);
and U925 (N_925,In_171,In_29);
nor U926 (N_926,In_315,In_233);
nor U927 (N_927,In_96,In_189);
nand U928 (N_928,In_245,In_466);
nor U929 (N_929,In_210,In_483);
or U930 (N_930,In_459,In_341);
or U931 (N_931,In_489,In_122);
or U932 (N_932,In_145,In_342);
or U933 (N_933,In_449,In_258);
nor U934 (N_934,In_57,In_214);
or U935 (N_935,In_486,In_43);
nand U936 (N_936,In_489,In_370);
nand U937 (N_937,In_68,In_15);
nand U938 (N_938,In_275,In_160);
nand U939 (N_939,In_335,In_145);
nand U940 (N_940,In_437,In_470);
nor U941 (N_941,In_497,In_453);
nand U942 (N_942,In_271,In_219);
and U943 (N_943,In_292,In_173);
nand U944 (N_944,In_408,In_492);
nand U945 (N_945,In_42,In_149);
nor U946 (N_946,In_250,In_158);
xor U947 (N_947,In_406,In_340);
nand U948 (N_948,In_464,In_309);
nand U949 (N_949,In_346,In_483);
and U950 (N_950,In_255,In_299);
nand U951 (N_951,In_470,In_400);
or U952 (N_952,In_24,In_163);
xor U953 (N_953,In_126,In_319);
nand U954 (N_954,In_298,In_67);
nand U955 (N_955,In_232,In_227);
nand U956 (N_956,In_198,In_101);
or U957 (N_957,In_355,In_163);
or U958 (N_958,In_195,In_76);
or U959 (N_959,In_444,In_392);
xor U960 (N_960,In_48,In_377);
and U961 (N_961,In_44,In_65);
and U962 (N_962,In_454,In_208);
nand U963 (N_963,In_251,In_350);
or U964 (N_964,In_135,In_155);
nand U965 (N_965,In_333,In_116);
nand U966 (N_966,In_290,In_426);
and U967 (N_967,In_347,In_211);
nand U968 (N_968,In_193,In_176);
nor U969 (N_969,In_13,In_489);
and U970 (N_970,In_349,In_490);
or U971 (N_971,In_266,In_156);
or U972 (N_972,In_481,In_76);
nand U973 (N_973,In_386,In_1);
nand U974 (N_974,In_12,In_45);
xor U975 (N_975,In_185,In_328);
nor U976 (N_976,In_198,In_274);
xor U977 (N_977,In_313,In_254);
xor U978 (N_978,In_105,In_461);
xor U979 (N_979,In_52,In_169);
xnor U980 (N_980,In_135,In_74);
and U981 (N_981,In_438,In_311);
nor U982 (N_982,In_181,In_62);
nor U983 (N_983,In_331,In_4);
or U984 (N_984,In_117,In_178);
or U985 (N_985,In_14,In_409);
and U986 (N_986,In_179,In_422);
xor U987 (N_987,In_189,In_254);
xnor U988 (N_988,In_236,In_105);
nand U989 (N_989,In_182,In_44);
nand U990 (N_990,In_172,In_279);
or U991 (N_991,In_448,In_226);
nor U992 (N_992,In_351,In_251);
or U993 (N_993,In_195,In_240);
xor U994 (N_994,In_217,In_54);
or U995 (N_995,In_109,In_413);
xor U996 (N_996,In_313,In_6);
or U997 (N_997,In_340,In_351);
xnor U998 (N_998,In_9,In_481);
xnor U999 (N_999,In_409,In_103);
xnor U1000 (N_1000,N_162,N_610);
xor U1001 (N_1001,N_246,N_625);
xnor U1002 (N_1002,N_488,N_928);
or U1003 (N_1003,N_409,N_662);
and U1004 (N_1004,N_795,N_211);
or U1005 (N_1005,N_580,N_512);
or U1006 (N_1006,N_865,N_345);
or U1007 (N_1007,N_612,N_283);
nand U1008 (N_1008,N_584,N_650);
nand U1009 (N_1009,N_78,N_820);
nor U1010 (N_1010,N_915,N_407);
xor U1011 (N_1011,N_517,N_875);
xor U1012 (N_1012,N_989,N_482);
nor U1013 (N_1013,N_722,N_51);
xor U1014 (N_1014,N_567,N_449);
nor U1015 (N_1015,N_961,N_481);
xnor U1016 (N_1016,N_579,N_30);
nor U1017 (N_1017,N_144,N_430);
nor U1018 (N_1018,N_737,N_770);
or U1019 (N_1019,N_901,N_976);
or U1020 (N_1020,N_575,N_745);
or U1021 (N_1021,N_158,N_997);
nor U1022 (N_1022,N_11,N_728);
and U1023 (N_1023,N_359,N_63);
xnor U1024 (N_1024,N_823,N_185);
nand U1025 (N_1025,N_643,N_186);
and U1026 (N_1026,N_548,N_590);
and U1027 (N_1027,N_883,N_787);
or U1028 (N_1028,N_251,N_959);
nor U1029 (N_1029,N_759,N_425);
and U1030 (N_1030,N_635,N_805);
and U1031 (N_1031,N_206,N_431);
and U1032 (N_1032,N_896,N_131);
and U1033 (N_1033,N_320,N_258);
and U1034 (N_1034,N_726,N_80);
and U1035 (N_1035,N_421,N_515);
and U1036 (N_1036,N_478,N_862);
or U1037 (N_1037,N_853,N_767);
xnor U1038 (N_1038,N_744,N_781);
or U1039 (N_1039,N_221,N_957);
xor U1040 (N_1040,N_255,N_557);
xor U1041 (N_1041,N_659,N_10);
nor U1042 (N_1042,N_911,N_236);
nor U1043 (N_1043,N_129,N_536);
and U1044 (N_1044,N_760,N_943);
or U1045 (N_1045,N_688,N_969);
and U1046 (N_1046,N_285,N_968);
or U1047 (N_1047,N_631,N_748);
and U1048 (N_1048,N_429,N_125);
xor U1049 (N_1049,N_72,N_730);
or U1050 (N_1050,N_32,N_35);
nor U1051 (N_1051,N_237,N_462);
nor U1052 (N_1052,N_617,N_633);
or U1053 (N_1053,N_403,N_360);
or U1054 (N_1054,N_215,N_471);
nand U1055 (N_1055,N_97,N_323);
or U1056 (N_1056,N_279,N_134);
nand U1057 (N_1057,N_920,N_783);
xor U1058 (N_1058,N_167,N_61);
nand U1059 (N_1059,N_514,N_970);
xor U1060 (N_1060,N_9,N_898);
xnor U1061 (N_1061,N_543,N_739);
or U1062 (N_1062,N_933,N_428);
or U1063 (N_1063,N_127,N_678);
or U1064 (N_1064,N_302,N_480);
or U1065 (N_1065,N_982,N_519);
and U1066 (N_1066,N_333,N_20);
and U1067 (N_1067,N_484,N_367);
or U1068 (N_1068,N_287,N_460);
xor U1069 (N_1069,N_347,N_294);
and U1070 (N_1070,N_469,N_310);
nor U1071 (N_1071,N_395,N_582);
and U1072 (N_1072,N_855,N_570);
or U1073 (N_1073,N_538,N_335);
nor U1074 (N_1074,N_467,N_504);
and U1075 (N_1075,N_521,N_904);
nand U1076 (N_1076,N_38,N_379);
xnor U1077 (N_1077,N_498,N_723);
and U1078 (N_1078,N_241,N_50);
nor U1079 (N_1079,N_293,N_919);
nor U1080 (N_1080,N_275,N_792);
nand U1081 (N_1081,N_161,N_712);
nand U1082 (N_1082,N_905,N_160);
nor U1083 (N_1083,N_159,N_942);
nor U1084 (N_1084,N_363,N_43);
xor U1085 (N_1085,N_637,N_269);
xnor U1086 (N_1086,N_668,N_581);
nor U1087 (N_1087,N_205,N_235);
xnor U1088 (N_1088,N_48,N_846);
xnor U1089 (N_1089,N_966,N_117);
nand U1090 (N_1090,N_630,N_417);
or U1091 (N_1091,N_690,N_743);
or U1092 (N_1092,N_472,N_714);
and U1093 (N_1093,N_442,N_277);
or U1094 (N_1094,N_41,N_344);
nor U1095 (N_1095,N_910,N_150);
nand U1096 (N_1096,N_500,N_252);
and U1097 (N_1097,N_595,N_863);
xnor U1098 (N_1098,N_94,N_667);
xnor U1099 (N_1099,N_278,N_921);
and U1100 (N_1100,N_243,N_376);
and U1101 (N_1101,N_647,N_719);
nand U1102 (N_1102,N_636,N_326);
nand U1103 (N_1103,N_420,N_939);
nor U1104 (N_1104,N_308,N_785);
or U1105 (N_1105,N_300,N_353);
and U1106 (N_1106,N_151,N_180);
or U1107 (N_1107,N_374,N_149);
and U1108 (N_1108,N_571,N_291);
and U1109 (N_1109,N_172,N_842);
nor U1110 (N_1110,N_39,N_356);
or U1111 (N_1111,N_53,N_837);
and U1112 (N_1112,N_383,N_870);
xnor U1113 (N_1113,N_57,N_495);
nor U1114 (N_1114,N_272,N_746);
xor U1115 (N_1115,N_541,N_950);
nor U1116 (N_1116,N_917,N_819);
xnor U1117 (N_1117,N_537,N_700);
nand U1118 (N_1118,N_434,N_124);
nand U1119 (N_1119,N_156,N_13);
or U1120 (N_1120,N_96,N_49);
xnor U1121 (N_1121,N_104,N_711);
nand U1122 (N_1122,N_187,N_314);
xor U1123 (N_1123,N_847,N_660);
and U1124 (N_1124,N_200,N_193);
xnor U1125 (N_1125,N_720,N_16);
xnor U1126 (N_1126,N_486,N_796);
nand U1127 (N_1127,N_249,N_408);
xor U1128 (N_1128,N_192,N_598);
and U1129 (N_1129,N_317,N_591);
xnor U1130 (N_1130,N_142,N_299);
and U1131 (N_1131,N_544,N_228);
nor U1132 (N_1132,N_814,N_618);
and U1133 (N_1133,N_130,N_105);
xor U1134 (N_1134,N_756,N_262);
xor U1135 (N_1135,N_47,N_520);
xnor U1136 (N_1136,N_75,N_422);
and U1137 (N_1137,N_59,N_68);
nor U1138 (N_1138,N_600,N_931);
nor U1139 (N_1139,N_912,N_766);
and U1140 (N_1140,N_804,N_574);
nand U1141 (N_1141,N_138,N_392);
nand U1142 (N_1142,N_747,N_717);
nor U1143 (N_1143,N_807,N_736);
nor U1144 (N_1144,N_621,N_455);
nand U1145 (N_1145,N_112,N_485);
xor U1146 (N_1146,N_163,N_316);
or U1147 (N_1147,N_466,N_527);
or U1148 (N_1148,N_679,N_704);
and U1149 (N_1149,N_852,N_616);
nand U1150 (N_1150,N_450,N_17);
nand U1151 (N_1151,N_2,N_531);
nor U1152 (N_1152,N_542,N_860);
xor U1153 (N_1153,N_83,N_639);
and U1154 (N_1154,N_391,N_168);
and U1155 (N_1155,N_250,N_828);
or U1156 (N_1156,N_330,N_708);
nand U1157 (N_1157,N_476,N_705);
nor U1158 (N_1158,N_508,N_216);
or U1159 (N_1159,N_406,N_627);
nand U1160 (N_1160,N_812,N_588);
nor U1161 (N_1161,N_682,N_733);
and U1162 (N_1162,N_93,N_0);
nand U1163 (N_1163,N_967,N_390);
nand U1164 (N_1164,N_977,N_419);
xor U1165 (N_1165,N_114,N_809);
nand U1166 (N_1166,N_701,N_55);
nand U1167 (N_1167,N_735,N_622);
nand U1168 (N_1168,N_882,N_348);
or U1169 (N_1169,N_932,N_769);
xnor U1170 (N_1170,N_295,N_926);
xor U1171 (N_1171,N_751,N_410);
and U1172 (N_1172,N_398,N_597);
nor U1173 (N_1173,N_505,N_341);
and U1174 (N_1174,N_899,N_208);
xnor U1175 (N_1175,N_689,N_790);
nand U1176 (N_1176,N_468,N_128);
xnor U1177 (N_1177,N_85,N_585);
or U1178 (N_1178,N_568,N_534);
nand U1179 (N_1179,N_210,N_493);
or U1180 (N_1180,N_135,N_857);
nor U1181 (N_1181,N_451,N_841);
xor U1182 (N_1182,N_626,N_964);
and U1183 (N_1183,N_835,N_593);
and U1184 (N_1184,N_724,N_902);
or U1185 (N_1185,N_411,N_608);
nand U1186 (N_1186,N_141,N_439);
xor U1187 (N_1187,N_780,N_143);
nand U1188 (N_1188,N_492,N_992);
nand U1189 (N_1189,N_350,N_979);
nand U1190 (N_1190,N_753,N_290);
nor U1191 (N_1191,N_757,N_473);
nor U1192 (N_1192,N_586,N_818);
xnor U1193 (N_1193,N_65,N_895);
nand U1194 (N_1194,N_336,N_634);
nand U1195 (N_1195,N_664,N_803);
and U1196 (N_1196,N_424,N_975);
and U1197 (N_1197,N_132,N_303);
nand U1198 (N_1198,N_884,N_672);
or U1199 (N_1199,N_92,N_569);
nand U1200 (N_1200,N_201,N_264);
or U1201 (N_1201,N_87,N_553);
and U1202 (N_1202,N_872,N_599);
or U1203 (N_1203,N_697,N_242);
nand U1204 (N_1204,N_653,N_503);
xnor U1205 (N_1205,N_772,N_980);
and U1206 (N_1206,N_827,N_988);
or U1207 (N_1207,N_893,N_764);
xnor U1208 (N_1208,N_64,N_227);
xnor U1209 (N_1209,N_873,N_324);
and U1210 (N_1210,N_154,N_373);
nand U1211 (N_1211,N_233,N_958);
or U1212 (N_1212,N_540,N_686);
and U1213 (N_1213,N_266,N_220);
xnor U1214 (N_1214,N_171,N_611);
and U1215 (N_1215,N_256,N_869);
nand U1216 (N_1216,N_620,N_362);
nand U1217 (N_1217,N_123,N_522);
or U1218 (N_1218,N_489,N_497);
nor U1219 (N_1219,N_773,N_765);
xnor U1220 (N_1220,N_995,N_725);
and U1221 (N_1221,N_762,N_196);
nor U1222 (N_1222,N_42,N_673);
xor U1223 (N_1223,N_589,N_111);
or U1224 (N_1224,N_157,N_954);
or U1225 (N_1225,N_868,N_122);
xor U1226 (N_1226,N_176,N_808);
xnor U1227 (N_1227,N_399,N_754);
nor U1228 (N_1228,N_306,N_240);
or U1229 (N_1229,N_602,N_576);
nand U1230 (N_1230,N_385,N_716);
nand U1231 (N_1231,N_229,N_118);
nand U1232 (N_1232,N_22,N_331);
nor U1233 (N_1233,N_60,N_935);
xnor U1234 (N_1234,N_758,N_908);
nor U1235 (N_1235,N_632,N_29);
nand U1236 (N_1236,N_800,N_594);
nand U1237 (N_1237,N_121,N_5);
xnor U1238 (N_1238,N_402,N_661);
or U1239 (N_1239,N_839,N_934);
or U1240 (N_1240,N_509,N_26);
and U1241 (N_1241,N_784,N_596);
xor U1242 (N_1242,N_327,N_671);
xnor U1243 (N_1243,N_365,N_502);
nor U1244 (N_1244,N_831,N_448);
nand U1245 (N_1245,N_197,N_603);
or U1246 (N_1246,N_73,N_925);
xnor U1247 (N_1247,N_674,N_707);
or U1248 (N_1248,N_28,N_95);
nand U1249 (N_1249,N_226,N_445);
and U1250 (N_1250,N_381,N_179);
or U1251 (N_1251,N_761,N_427);
nor U1252 (N_1252,N_774,N_271);
and U1253 (N_1253,N_414,N_194);
xnor U1254 (N_1254,N_566,N_742);
nor U1255 (N_1255,N_551,N_101);
and U1256 (N_1256,N_413,N_940);
and U1257 (N_1257,N_230,N_254);
or U1258 (N_1258,N_401,N_532);
xor U1259 (N_1259,N_972,N_558);
nor U1260 (N_1260,N_535,N_483);
and U1261 (N_1261,N_793,N_153);
nor U1262 (N_1262,N_789,N_510);
xor U1263 (N_1263,N_552,N_821);
or U1264 (N_1264,N_801,N_811);
nor U1265 (N_1265,N_182,N_311);
xnor U1266 (N_1266,N_328,N_525);
xnor U1267 (N_1267,N_457,N_877);
and U1268 (N_1268,N_177,N_443);
and U1269 (N_1269,N_209,N_88);
nand U1270 (N_1270,N_866,N_990);
and U1271 (N_1271,N_775,N_786);
nor U1272 (N_1272,N_296,N_313);
nor U1273 (N_1273,N_885,N_874);
xor U1274 (N_1274,N_684,N_788);
or U1275 (N_1275,N_628,N_945);
xnor U1276 (N_1276,N_338,N_438);
xor U1277 (N_1277,N_948,N_152);
nand U1278 (N_1278,N_40,N_985);
and U1279 (N_1279,N_54,N_559);
or U1280 (N_1280,N_560,N_231);
and U1281 (N_1281,N_530,N_499);
nand U1282 (N_1282,N_477,N_393);
and U1283 (N_1283,N_415,N_223);
or U1284 (N_1284,N_76,N_273);
and U1285 (N_1285,N_378,N_346);
and U1286 (N_1286,N_507,N_691);
xnor U1287 (N_1287,N_369,N_366);
and U1288 (N_1288,N_609,N_46);
nand U1289 (N_1289,N_991,N_315);
or U1290 (N_1290,N_615,N_960);
and U1291 (N_1291,N_944,N_444);
nor U1292 (N_1292,N_386,N_98);
nor U1293 (N_1293,N_687,N_918);
nand U1294 (N_1294,N_71,N_802);
xor U1295 (N_1295,N_859,N_815);
nor U1296 (N_1296,N_810,N_305);
or U1297 (N_1297,N_528,N_994);
nand U1298 (N_1298,N_613,N_261);
xnor U1299 (N_1299,N_511,N_974);
nor U1300 (N_1300,N_973,N_562);
or U1301 (N_1301,N_694,N_851);
and U1302 (N_1302,N_195,N_833);
or U1303 (N_1303,N_490,N_494);
nor U1304 (N_1304,N_377,N_955);
xnor U1305 (N_1305,N_234,N_867);
nor U1306 (N_1306,N_693,N_307);
nor U1307 (N_1307,N_861,N_265);
nand U1308 (N_1308,N_993,N_267);
xnor U1309 (N_1309,N_782,N_849);
nor U1310 (N_1310,N_268,N_665);
xnor U1311 (N_1311,N_394,N_706);
nand U1312 (N_1312,N_550,N_147);
xor U1313 (N_1313,N_24,N_830);
and U1314 (N_1314,N_946,N_914);
xor U1315 (N_1315,N_930,N_212);
and U1316 (N_1316,N_642,N_836);
xor U1317 (N_1317,N_126,N_583);
or U1318 (N_1318,N_139,N_282);
nor U1319 (N_1319,N_843,N_458);
and U1320 (N_1320,N_813,N_52);
or U1321 (N_1321,N_19,N_337);
nor U1322 (N_1322,N_604,N_198);
nand U1323 (N_1323,N_343,N_965);
nor U1324 (N_1324,N_654,N_213);
or U1325 (N_1325,N_4,N_368);
xor U1326 (N_1326,N_881,N_644);
or U1327 (N_1327,N_913,N_82);
nand U1328 (N_1328,N_446,N_380);
and U1329 (N_1329,N_189,N_794);
nor U1330 (N_1330,N_685,N_909);
xor U1331 (N_1331,N_916,N_69);
and U1332 (N_1332,N_734,N_937);
nor U1333 (N_1333,N_718,N_845);
nor U1334 (N_1334,N_938,N_396);
nand U1335 (N_1335,N_70,N_222);
nor U1336 (N_1336,N_33,N_826);
and U1337 (N_1337,N_155,N_680);
xor U1338 (N_1338,N_288,N_81);
xnor U1339 (N_1339,N_702,N_703);
nand U1340 (N_1340,N_854,N_217);
nand U1341 (N_1341,N_470,N_832);
or U1342 (N_1342,N_165,N_318);
nand U1343 (N_1343,N_113,N_166);
or U1344 (N_1344,N_983,N_436);
nor U1345 (N_1345,N_297,N_270);
nor U1346 (N_1346,N_136,N_645);
nand U1347 (N_1347,N_669,N_658);
nor U1348 (N_1348,N_715,N_732);
and U1349 (N_1349,N_418,N_100);
xor U1350 (N_1350,N_892,N_204);
xnor U1351 (N_1351,N_397,N_607);
nor U1352 (N_1352,N_641,N_646);
nand U1353 (N_1353,N_14,N_174);
nor U1354 (N_1354,N_453,N_922);
nor U1355 (N_1355,N_66,N_452);
xnor U1356 (N_1356,N_247,N_244);
xnor U1357 (N_1357,N_798,N_304);
nor U1358 (N_1358,N_533,N_286);
nand U1359 (N_1359,N_103,N_190);
and U1360 (N_1360,N_322,N_349);
nor U1361 (N_1361,N_546,N_137);
or U1362 (N_1362,N_806,N_962);
and U1363 (N_1363,N_239,N_999);
nand U1364 (N_1364,N_140,N_663);
nand U1365 (N_1365,N_695,N_888);
nand U1366 (N_1366,N_108,N_58);
xnor U1367 (N_1367,N_437,N_740);
and U1368 (N_1368,N_191,N_624);
and U1369 (N_1369,N_894,N_25);
or U1370 (N_1370,N_840,N_464);
nand U1371 (N_1371,N_683,N_120);
xnor U1372 (N_1372,N_890,N_84);
or U1373 (N_1373,N_924,N_698);
nand U1374 (N_1374,N_173,N_292);
xor U1375 (N_1375,N_109,N_332);
or U1376 (N_1376,N_146,N_99);
nand U1377 (N_1377,N_440,N_325);
nor U1378 (N_1378,N_184,N_214);
or U1379 (N_1379,N_44,N_253);
nand U1380 (N_1380,N_8,N_459);
nor U1381 (N_1381,N_987,N_880);
and U1382 (N_1382,N_879,N_465);
or U1383 (N_1383,N_677,N_829);
or U1384 (N_1384,N_578,N_479);
and U1385 (N_1385,N_433,N_986);
or U1386 (N_1386,N_648,N_856);
nor U1387 (N_1387,N_768,N_750);
or U1388 (N_1388,N_963,N_947);
and U1389 (N_1389,N_412,N_281);
nand U1390 (N_1390,N_903,N_148);
xnor U1391 (N_1391,N_441,N_956);
or U1392 (N_1392,N_79,N_727);
nand U1393 (N_1393,N_729,N_886);
and U1394 (N_1394,N_501,N_513);
nand U1395 (N_1395,N_91,N_878);
xor U1396 (N_1396,N_848,N_876);
nand U1397 (N_1397,N_749,N_529);
or U1398 (N_1398,N_655,N_423);
nand U1399 (N_1399,N_547,N_565);
or U1400 (N_1400,N_941,N_629);
nand U1401 (N_1401,N_797,N_906);
nand U1402 (N_1402,N_86,N_850);
and U1403 (N_1403,N_432,N_822);
nor U1404 (N_1404,N_203,N_889);
nand U1405 (N_1405,N_670,N_996);
or U1406 (N_1406,N_526,N_907);
xor U1407 (N_1407,N_372,N_755);
and U1408 (N_1408,N_340,N_900);
nor U1409 (N_1409,N_649,N_110);
nand U1410 (N_1410,N_825,N_516);
or U1411 (N_1411,N_188,N_183);
nand U1412 (N_1412,N_454,N_936);
or U1413 (N_1413,N_864,N_280);
nand U1414 (N_1414,N_404,N_107);
and U1415 (N_1415,N_834,N_334);
or U1416 (N_1416,N_248,N_358);
nand U1417 (N_1417,N_518,N_27);
nor U1418 (N_1418,N_496,N_34);
nand U1419 (N_1419,N_657,N_354);
or U1420 (N_1420,N_555,N_232);
xnor U1421 (N_1421,N_321,N_351);
xnor U1422 (N_1422,N_752,N_572);
nor U1423 (N_1423,N_21,N_384);
nor U1424 (N_1424,N_981,N_36);
xor U1425 (N_1425,N_435,N_897);
nand U1426 (N_1426,N_676,N_426);
xnor U1427 (N_1427,N_319,N_289);
and U1428 (N_1428,N_927,N_67);
or U1429 (N_1429,N_984,N_224);
nor U1430 (N_1430,N_219,N_587);
nand U1431 (N_1431,N_89,N_355);
nor U1432 (N_1432,N_31,N_799);
xnor U1433 (N_1433,N_606,N_692);
nor U1434 (N_1434,N_699,N_475);
or U1435 (N_1435,N_312,N_656);
or U1436 (N_1436,N_77,N_563);
xnor U1437 (N_1437,N_45,N_474);
and U1438 (N_1438,N_116,N_738);
and U1439 (N_1439,N_556,N_309);
xnor U1440 (N_1440,N_858,N_952);
nand U1441 (N_1441,N_561,N_605);
nor U1442 (N_1442,N_175,N_257);
nand U1443 (N_1443,N_545,N_169);
nor U1444 (N_1444,N_524,N_953);
and U1445 (N_1445,N_284,N_923);
and U1446 (N_1446,N_577,N_721);
nor U1447 (N_1447,N_342,N_106);
nor U1448 (N_1448,N_298,N_145);
nor U1449 (N_1449,N_640,N_929);
or U1450 (N_1450,N_15,N_259);
and U1451 (N_1451,N_709,N_115);
and U1452 (N_1452,N_405,N_549);
xnor U1453 (N_1453,N_564,N_276);
and U1454 (N_1454,N_6,N_978);
nor U1455 (N_1455,N_90,N_388);
nor U1456 (N_1456,N_400,N_731);
and U1457 (N_1457,N_681,N_181);
or U1458 (N_1458,N_971,N_871);
nand U1459 (N_1459,N_218,N_202);
and U1460 (N_1460,N_652,N_416);
and U1461 (N_1461,N_771,N_891);
or U1462 (N_1462,N_506,N_37);
nand U1463 (N_1463,N_824,N_675);
nor U1464 (N_1464,N_352,N_463);
nor U1465 (N_1465,N_18,N_178);
xnor U1466 (N_1466,N_949,N_447);
and U1467 (N_1467,N_998,N_778);
and U1468 (N_1468,N_62,N_329);
xor U1469 (N_1469,N_12,N_741);
xor U1470 (N_1470,N_887,N_523);
and U1471 (N_1471,N_357,N_614);
nor U1472 (N_1472,N_164,N_238);
xnor U1473 (N_1473,N_554,N_619);
nor U1474 (N_1474,N_696,N_776);
xnor U1475 (N_1475,N_816,N_274);
xor U1476 (N_1476,N_199,N_651);
and U1477 (N_1477,N_119,N_387);
nor U1478 (N_1478,N_456,N_491);
nand U1479 (N_1479,N_539,N_361);
nand U1480 (N_1480,N_638,N_370);
xnor U1481 (N_1481,N_844,N_710);
nand U1482 (N_1482,N_102,N_623);
nor U1483 (N_1483,N_339,N_375);
xor U1484 (N_1484,N_23,N_487);
nor U1485 (N_1485,N_389,N_207);
and U1486 (N_1486,N_666,N_777);
xnor U1487 (N_1487,N_371,N_74);
or U1488 (N_1488,N_1,N_170);
xnor U1489 (N_1489,N_7,N_601);
or U1490 (N_1490,N_763,N_245);
xor U1491 (N_1491,N_382,N_713);
xnor U1492 (N_1492,N_951,N_133);
xnor U1493 (N_1493,N_838,N_364);
xor U1494 (N_1494,N_779,N_225);
and U1495 (N_1495,N_573,N_3);
nand U1496 (N_1496,N_260,N_592);
nand U1497 (N_1497,N_791,N_301);
nor U1498 (N_1498,N_56,N_263);
and U1499 (N_1499,N_461,N_817);
or U1500 (N_1500,N_71,N_645);
xor U1501 (N_1501,N_681,N_287);
nand U1502 (N_1502,N_59,N_144);
nand U1503 (N_1503,N_570,N_560);
nor U1504 (N_1504,N_882,N_747);
and U1505 (N_1505,N_575,N_225);
and U1506 (N_1506,N_718,N_690);
and U1507 (N_1507,N_759,N_705);
nor U1508 (N_1508,N_869,N_437);
nand U1509 (N_1509,N_451,N_916);
nor U1510 (N_1510,N_581,N_630);
or U1511 (N_1511,N_381,N_264);
nand U1512 (N_1512,N_611,N_139);
or U1513 (N_1513,N_705,N_933);
nor U1514 (N_1514,N_0,N_217);
nand U1515 (N_1515,N_151,N_647);
and U1516 (N_1516,N_472,N_544);
and U1517 (N_1517,N_541,N_376);
or U1518 (N_1518,N_36,N_456);
or U1519 (N_1519,N_403,N_781);
xor U1520 (N_1520,N_726,N_803);
nor U1521 (N_1521,N_480,N_200);
nor U1522 (N_1522,N_952,N_496);
or U1523 (N_1523,N_445,N_224);
nor U1524 (N_1524,N_329,N_375);
xnor U1525 (N_1525,N_182,N_427);
nand U1526 (N_1526,N_54,N_212);
and U1527 (N_1527,N_135,N_497);
xnor U1528 (N_1528,N_823,N_676);
or U1529 (N_1529,N_139,N_846);
nand U1530 (N_1530,N_928,N_497);
xor U1531 (N_1531,N_322,N_829);
or U1532 (N_1532,N_447,N_129);
nand U1533 (N_1533,N_301,N_651);
nor U1534 (N_1534,N_839,N_200);
xnor U1535 (N_1535,N_877,N_490);
nand U1536 (N_1536,N_236,N_553);
nor U1537 (N_1537,N_583,N_576);
or U1538 (N_1538,N_637,N_360);
and U1539 (N_1539,N_509,N_418);
xnor U1540 (N_1540,N_335,N_628);
or U1541 (N_1541,N_272,N_598);
nand U1542 (N_1542,N_714,N_494);
and U1543 (N_1543,N_600,N_520);
and U1544 (N_1544,N_714,N_925);
and U1545 (N_1545,N_720,N_879);
and U1546 (N_1546,N_731,N_482);
and U1547 (N_1547,N_350,N_778);
and U1548 (N_1548,N_272,N_930);
or U1549 (N_1549,N_105,N_3);
nand U1550 (N_1550,N_16,N_773);
xor U1551 (N_1551,N_737,N_971);
or U1552 (N_1552,N_735,N_194);
xnor U1553 (N_1553,N_893,N_233);
xnor U1554 (N_1554,N_163,N_973);
and U1555 (N_1555,N_520,N_991);
nor U1556 (N_1556,N_213,N_922);
xor U1557 (N_1557,N_552,N_387);
or U1558 (N_1558,N_518,N_943);
nand U1559 (N_1559,N_848,N_315);
xnor U1560 (N_1560,N_10,N_674);
xor U1561 (N_1561,N_44,N_942);
xnor U1562 (N_1562,N_656,N_775);
and U1563 (N_1563,N_14,N_212);
nor U1564 (N_1564,N_669,N_510);
xnor U1565 (N_1565,N_859,N_614);
xor U1566 (N_1566,N_634,N_183);
or U1567 (N_1567,N_867,N_487);
nand U1568 (N_1568,N_384,N_821);
or U1569 (N_1569,N_657,N_203);
nand U1570 (N_1570,N_29,N_124);
xor U1571 (N_1571,N_372,N_915);
nand U1572 (N_1572,N_757,N_514);
nand U1573 (N_1573,N_375,N_337);
nand U1574 (N_1574,N_353,N_813);
and U1575 (N_1575,N_260,N_367);
nor U1576 (N_1576,N_715,N_988);
xnor U1577 (N_1577,N_508,N_518);
nor U1578 (N_1578,N_457,N_437);
nand U1579 (N_1579,N_720,N_220);
or U1580 (N_1580,N_234,N_215);
xnor U1581 (N_1581,N_509,N_530);
and U1582 (N_1582,N_710,N_489);
and U1583 (N_1583,N_308,N_285);
nand U1584 (N_1584,N_836,N_189);
or U1585 (N_1585,N_925,N_591);
and U1586 (N_1586,N_168,N_952);
xnor U1587 (N_1587,N_88,N_950);
nand U1588 (N_1588,N_326,N_658);
nand U1589 (N_1589,N_159,N_856);
and U1590 (N_1590,N_68,N_407);
nor U1591 (N_1591,N_988,N_682);
nand U1592 (N_1592,N_751,N_288);
xnor U1593 (N_1593,N_407,N_300);
xnor U1594 (N_1594,N_744,N_348);
nand U1595 (N_1595,N_609,N_242);
or U1596 (N_1596,N_817,N_408);
xnor U1597 (N_1597,N_13,N_867);
nand U1598 (N_1598,N_777,N_352);
and U1599 (N_1599,N_4,N_407);
nand U1600 (N_1600,N_188,N_277);
xnor U1601 (N_1601,N_289,N_629);
and U1602 (N_1602,N_171,N_183);
and U1603 (N_1603,N_236,N_455);
or U1604 (N_1604,N_402,N_869);
and U1605 (N_1605,N_936,N_277);
xor U1606 (N_1606,N_124,N_869);
nand U1607 (N_1607,N_639,N_323);
or U1608 (N_1608,N_621,N_642);
or U1609 (N_1609,N_176,N_833);
nor U1610 (N_1610,N_564,N_502);
xor U1611 (N_1611,N_979,N_472);
and U1612 (N_1612,N_89,N_447);
xor U1613 (N_1613,N_76,N_73);
nor U1614 (N_1614,N_916,N_727);
nor U1615 (N_1615,N_975,N_394);
nand U1616 (N_1616,N_838,N_872);
or U1617 (N_1617,N_503,N_912);
and U1618 (N_1618,N_498,N_415);
nand U1619 (N_1619,N_653,N_393);
xnor U1620 (N_1620,N_486,N_825);
or U1621 (N_1621,N_581,N_86);
and U1622 (N_1622,N_314,N_527);
xor U1623 (N_1623,N_254,N_167);
xnor U1624 (N_1624,N_955,N_76);
and U1625 (N_1625,N_301,N_727);
nor U1626 (N_1626,N_980,N_414);
xnor U1627 (N_1627,N_212,N_135);
nor U1628 (N_1628,N_115,N_155);
nor U1629 (N_1629,N_548,N_309);
or U1630 (N_1630,N_275,N_648);
or U1631 (N_1631,N_452,N_793);
nand U1632 (N_1632,N_924,N_951);
and U1633 (N_1633,N_592,N_606);
xnor U1634 (N_1634,N_964,N_310);
nor U1635 (N_1635,N_227,N_515);
or U1636 (N_1636,N_269,N_253);
nor U1637 (N_1637,N_757,N_658);
and U1638 (N_1638,N_548,N_318);
or U1639 (N_1639,N_32,N_817);
nor U1640 (N_1640,N_145,N_574);
nor U1641 (N_1641,N_756,N_146);
nor U1642 (N_1642,N_921,N_295);
and U1643 (N_1643,N_566,N_338);
nand U1644 (N_1644,N_283,N_957);
and U1645 (N_1645,N_913,N_416);
and U1646 (N_1646,N_616,N_403);
nor U1647 (N_1647,N_298,N_283);
and U1648 (N_1648,N_838,N_507);
xnor U1649 (N_1649,N_910,N_645);
nand U1650 (N_1650,N_959,N_640);
nor U1651 (N_1651,N_234,N_754);
nand U1652 (N_1652,N_565,N_671);
nor U1653 (N_1653,N_140,N_709);
xnor U1654 (N_1654,N_85,N_275);
nand U1655 (N_1655,N_437,N_11);
xnor U1656 (N_1656,N_645,N_852);
nor U1657 (N_1657,N_142,N_975);
or U1658 (N_1658,N_942,N_522);
and U1659 (N_1659,N_962,N_110);
xor U1660 (N_1660,N_227,N_971);
and U1661 (N_1661,N_638,N_991);
nand U1662 (N_1662,N_309,N_1);
nor U1663 (N_1663,N_170,N_208);
xnor U1664 (N_1664,N_519,N_732);
or U1665 (N_1665,N_936,N_170);
or U1666 (N_1666,N_423,N_277);
xnor U1667 (N_1667,N_296,N_516);
or U1668 (N_1668,N_144,N_328);
nor U1669 (N_1669,N_10,N_885);
nor U1670 (N_1670,N_707,N_358);
and U1671 (N_1671,N_35,N_515);
and U1672 (N_1672,N_696,N_146);
xor U1673 (N_1673,N_487,N_243);
or U1674 (N_1674,N_81,N_829);
and U1675 (N_1675,N_647,N_805);
and U1676 (N_1676,N_53,N_257);
or U1677 (N_1677,N_94,N_968);
and U1678 (N_1678,N_949,N_213);
nand U1679 (N_1679,N_674,N_729);
xor U1680 (N_1680,N_909,N_248);
nand U1681 (N_1681,N_11,N_325);
and U1682 (N_1682,N_782,N_4);
or U1683 (N_1683,N_663,N_986);
nor U1684 (N_1684,N_336,N_402);
or U1685 (N_1685,N_525,N_152);
nand U1686 (N_1686,N_437,N_617);
nand U1687 (N_1687,N_95,N_925);
nor U1688 (N_1688,N_559,N_455);
xnor U1689 (N_1689,N_725,N_235);
or U1690 (N_1690,N_783,N_651);
xor U1691 (N_1691,N_52,N_956);
xor U1692 (N_1692,N_256,N_328);
and U1693 (N_1693,N_996,N_667);
nand U1694 (N_1694,N_618,N_831);
xor U1695 (N_1695,N_475,N_463);
nand U1696 (N_1696,N_287,N_229);
and U1697 (N_1697,N_548,N_897);
nor U1698 (N_1698,N_575,N_46);
or U1699 (N_1699,N_767,N_404);
xnor U1700 (N_1700,N_797,N_885);
nor U1701 (N_1701,N_819,N_147);
and U1702 (N_1702,N_583,N_605);
xnor U1703 (N_1703,N_998,N_712);
and U1704 (N_1704,N_470,N_516);
and U1705 (N_1705,N_768,N_376);
xnor U1706 (N_1706,N_841,N_847);
xor U1707 (N_1707,N_90,N_631);
and U1708 (N_1708,N_602,N_779);
nor U1709 (N_1709,N_401,N_992);
nand U1710 (N_1710,N_274,N_497);
nand U1711 (N_1711,N_361,N_646);
and U1712 (N_1712,N_616,N_83);
nor U1713 (N_1713,N_890,N_936);
or U1714 (N_1714,N_367,N_146);
or U1715 (N_1715,N_241,N_936);
nor U1716 (N_1716,N_594,N_821);
and U1717 (N_1717,N_792,N_198);
or U1718 (N_1718,N_142,N_611);
nor U1719 (N_1719,N_350,N_902);
or U1720 (N_1720,N_183,N_101);
nor U1721 (N_1721,N_746,N_811);
nand U1722 (N_1722,N_262,N_957);
xnor U1723 (N_1723,N_349,N_472);
and U1724 (N_1724,N_835,N_789);
and U1725 (N_1725,N_963,N_206);
or U1726 (N_1726,N_29,N_56);
xor U1727 (N_1727,N_333,N_876);
nand U1728 (N_1728,N_41,N_392);
or U1729 (N_1729,N_424,N_833);
xor U1730 (N_1730,N_660,N_55);
or U1731 (N_1731,N_445,N_338);
nor U1732 (N_1732,N_980,N_149);
nand U1733 (N_1733,N_366,N_25);
nand U1734 (N_1734,N_339,N_215);
xor U1735 (N_1735,N_324,N_183);
or U1736 (N_1736,N_589,N_536);
and U1737 (N_1737,N_534,N_581);
or U1738 (N_1738,N_127,N_445);
nor U1739 (N_1739,N_497,N_791);
and U1740 (N_1740,N_501,N_416);
nor U1741 (N_1741,N_801,N_7);
or U1742 (N_1742,N_677,N_161);
nor U1743 (N_1743,N_715,N_701);
or U1744 (N_1744,N_619,N_652);
nand U1745 (N_1745,N_930,N_102);
or U1746 (N_1746,N_583,N_20);
and U1747 (N_1747,N_318,N_380);
and U1748 (N_1748,N_769,N_834);
nand U1749 (N_1749,N_98,N_661);
xor U1750 (N_1750,N_860,N_939);
nand U1751 (N_1751,N_100,N_118);
nand U1752 (N_1752,N_975,N_598);
or U1753 (N_1753,N_64,N_575);
and U1754 (N_1754,N_631,N_904);
xnor U1755 (N_1755,N_923,N_448);
xnor U1756 (N_1756,N_521,N_469);
nand U1757 (N_1757,N_43,N_305);
xor U1758 (N_1758,N_802,N_840);
nor U1759 (N_1759,N_183,N_640);
or U1760 (N_1760,N_488,N_632);
or U1761 (N_1761,N_231,N_110);
nor U1762 (N_1762,N_282,N_229);
xor U1763 (N_1763,N_955,N_791);
xor U1764 (N_1764,N_316,N_13);
nor U1765 (N_1765,N_7,N_782);
nand U1766 (N_1766,N_999,N_537);
and U1767 (N_1767,N_69,N_632);
nand U1768 (N_1768,N_478,N_732);
and U1769 (N_1769,N_13,N_162);
xor U1770 (N_1770,N_155,N_725);
and U1771 (N_1771,N_619,N_351);
nor U1772 (N_1772,N_794,N_113);
or U1773 (N_1773,N_14,N_589);
xnor U1774 (N_1774,N_141,N_178);
or U1775 (N_1775,N_191,N_322);
or U1776 (N_1776,N_986,N_156);
and U1777 (N_1777,N_697,N_415);
nand U1778 (N_1778,N_538,N_407);
and U1779 (N_1779,N_185,N_46);
or U1780 (N_1780,N_39,N_717);
and U1781 (N_1781,N_531,N_276);
nor U1782 (N_1782,N_991,N_487);
or U1783 (N_1783,N_628,N_438);
xnor U1784 (N_1784,N_82,N_517);
nor U1785 (N_1785,N_230,N_928);
or U1786 (N_1786,N_194,N_82);
and U1787 (N_1787,N_342,N_41);
or U1788 (N_1788,N_657,N_408);
xnor U1789 (N_1789,N_490,N_708);
or U1790 (N_1790,N_927,N_8);
or U1791 (N_1791,N_426,N_990);
nand U1792 (N_1792,N_80,N_894);
and U1793 (N_1793,N_24,N_479);
or U1794 (N_1794,N_755,N_859);
nor U1795 (N_1795,N_725,N_194);
nand U1796 (N_1796,N_831,N_573);
and U1797 (N_1797,N_869,N_144);
nand U1798 (N_1798,N_416,N_78);
nand U1799 (N_1799,N_795,N_864);
xor U1800 (N_1800,N_515,N_843);
or U1801 (N_1801,N_759,N_398);
nand U1802 (N_1802,N_835,N_51);
or U1803 (N_1803,N_761,N_249);
xor U1804 (N_1804,N_530,N_955);
nor U1805 (N_1805,N_614,N_323);
nor U1806 (N_1806,N_712,N_398);
nor U1807 (N_1807,N_795,N_903);
or U1808 (N_1808,N_134,N_678);
and U1809 (N_1809,N_434,N_118);
nand U1810 (N_1810,N_857,N_568);
and U1811 (N_1811,N_95,N_951);
nand U1812 (N_1812,N_949,N_831);
and U1813 (N_1813,N_111,N_142);
nor U1814 (N_1814,N_935,N_167);
nand U1815 (N_1815,N_711,N_557);
nand U1816 (N_1816,N_824,N_290);
or U1817 (N_1817,N_16,N_346);
or U1818 (N_1818,N_428,N_588);
xnor U1819 (N_1819,N_751,N_869);
nand U1820 (N_1820,N_842,N_530);
and U1821 (N_1821,N_847,N_350);
xnor U1822 (N_1822,N_508,N_872);
or U1823 (N_1823,N_800,N_967);
nand U1824 (N_1824,N_301,N_858);
or U1825 (N_1825,N_168,N_69);
and U1826 (N_1826,N_557,N_230);
nand U1827 (N_1827,N_739,N_35);
or U1828 (N_1828,N_486,N_601);
xnor U1829 (N_1829,N_274,N_146);
nor U1830 (N_1830,N_146,N_433);
nand U1831 (N_1831,N_409,N_71);
xor U1832 (N_1832,N_730,N_507);
xor U1833 (N_1833,N_60,N_66);
xnor U1834 (N_1834,N_874,N_69);
and U1835 (N_1835,N_52,N_951);
xnor U1836 (N_1836,N_890,N_786);
nand U1837 (N_1837,N_932,N_633);
nor U1838 (N_1838,N_514,N_650);
and U1839 (N_1839,N_763,N_344);
xor U1840 (N_1840,N_967,N_293);
nor U1841 (N_1841,N_931,N_644);
and U1842 (N_1842,N_560,N_168);
and U1843 (N_1843,N_141,N_898);
nand U1844 (N_1844,N_333,N_386);
or U1845 (N_1845,N_694,N_828);
xnor U1846 (N_1846,N_593,N_182);
xor U1847 (N_1847,N_512,N_689);
or U1848 (N_1848,N_365,N_497);
xor U1849 (N_1849,N_519,N_26);
nor U1850 (N_1850,N_583,N_972);
nor U1851 (N_1851,N_115,N_695);
or U1852 (N_1852,N_553,N_790);
or U1853 (N_1853,N_90,N_971);
or U1854 (N_1854,N_381,N_492);
xnor U1855 (N_1855,N_281,N_818);
and U1856 (N_1856,N_686,N_572);
nand U1857 (N_1857,N_683,N_710);
nor U1858 (N_1858,N_543,N_667);
nor U1859 (N_1859,N_589,N_845);
xnor U1860 (N_1860,N_785,N_420);
nand U1861 (N_1861,N_942,N_31);
nand U1862 (N_1862,N_691,N_835);
or U1863 (N_1863,N_495,N_332);
xnor U1864 (N_1864,N_312,N_928);
xnor U1865 (N_1865,N_198,N_721);
nor U1866 (N_1866,N_864,N_504);
or U1867 (N_1867,N_64,N_848);
nand U1868 (N_1868,N_333,N_786);
nor U1869 (N_1869,N_297,N_535);
xor U1870 (N_1870,N_57,N_519);
nor U1871 (N_1871,N_760,N_516);
and U1872 (N_1872,N_123,N_882);
nor U1873 (N_1873,N_772,N_928);
nand U1874 (N_1874,N_658,N_130);
and U1875 (N_1875,N_76,N_994);
nor U1876 (N_1876,N_647,N_43);
nor U1877 (N_1877,N_361,N_454);
or U1878 (N_1878,N_653,N_988);
xnor U1879 (N_1879,N_487,N_264);
or U1880 (N_1880,N_603,N_959);
nand U1881 (N_1881,N_665,N_694);
xnor U1882 (N_1882,N_940,N_663);
or U1883 (N_1883,N_424,N_425);
nor U1884 (N_1884,N_408,N_763);
nor U1885 (N_1885,N_679,N_751);
and U1886 (N_1886,N_584,N_419);
nand U1887 (N_1887,N_891,N_586);
or U1888 (N_1888,N_671,N_536);
or U1889 (N_1889,N_657,N_64);
xnor U1890 (N_1890,N_741,N_279);
and U1891 (N_1891,N_616,N_838);
or U1892 (N_1892,N_654,N_703);
nor U1893 (N_1893,N_938,N_785);
nand U1894 (N_1894,N_129,N_603);
and U1895 (N_1895,N_315,N_470);
nor U1896 (N_1896,N_989,N_474);
nand U1897 (N_1897,N_484,N_677);
or U1898 (N_1898,N_824,N_807);
and U1899 (N_1899,N_147,N_207);
nor U1900 (N_1900,N_60,N_578);
xor U1901 (N_1901,N_47,N_355);
and U1902 (N_1902,N_524,N_799);
or U1903 (N_1903,N_652,N_377);
nor U1904 (N_1904,N_370,N_70);
and U1905 (N_1905,N_262,N_484);
xor U1906 (N_1906,N_26,N_684);
and U1907 (N_1907,N_156,N_917);
nor U1908 (N_1908,N_101,N_325);
nand U1909 (N_1909,N_607,N_819);
nand U1910 (N_1910,N_195,N_311);
or U1911 (N_1911,N_677,N_926);
and U1912 (N_1912,N_764,N_713);
nand U1913 (N_1913,N_16,N_355);
and U1914 (N_1914,N_942,N_624);
xor U1915 (N_1915,N_95,N_177);
nor U1916 (N_1916,N_760,N_806);
and U1917 (N_1917,N_101,N_345);
nor U1918 (N_1918,N_3,N_135);
xor U1919 (N_1919,N_855,N_501);
nor U1920 (N_1920,N_502,N_976);
and U1921 (N_1921,N_178,N_990);
and U1922 (N_1922,N_180,N_915);
xnor U1923 (N_1923,N_540,N_305);
or U1924 (N_1924,N_194,N_161);
or U1925 (N_1925,N_6,N_697);
or U1926 (N_1926,N_270,N_975);
or U1927 (N_1927,N_134,N_68);
xnor U1928 (N_1928,N_459,N_471);
or U1929 (N_1929,N_921,N_386);
or U1930 (N_1930,N_905,N_754);
or U1931 (N_1931,N_709,N_517);
nand U1932 (N_1932,N_33,N_24);
xnor U1933 (N_1933,N_411,N_38);
nand U1934 (N_1934,N_445,N_681);
and U1935 (N_1935,N_622,N_188);
or U1936 (N_1936,N_374,N_453);
nand U1937 (N_1937,N_638,N_578);
or U1938 (N_1938,N_866,N_986);
xor U1939 (N_1939,N_425,N_60);
nor U1940 (N_1940,N_518,N_480);
xor U1941 (N_1941,N_8,N_618);
nor U1942 (N_1942,N_560,N_850);
nand U1943 (N_1943,N_377,N_666);
and U1944 (N_1944,N_691,N_615);
and U1945 (N_1945,N_476,N_971);
nand U1946 (N_1946,N_501,N_11);
xor U1947 (N_1947,N_469,N_783);
xnor U1948 (N_1948,N_192,N_315);
xor U1949 (N_1949,N_997,N_926);
nand U1950 (N_1950,N_802,N_84);
or U1951 (N_1951,N_468,N_143);
nand U1952 (N_1952,N_385,N_908);
nor U1953 (N_1953,N_862,N_15);
and U1954 (N_1954,N_18,N_529);
xor U1955 (N_1955,N_85,N_33);
nor U1956 (N_1956,N_362,N_159);
or U1957 (N_1957,N_364,N_191);
nand U1958 (N_1958,N_695,N_20);
nor U1959 (N_1959,N_58,N_555);
nor U1960 (N_1960,N_620,N_876);
nor U1961 (N_1961,N_73,N_439);
and U1962 (N_1962,N_486,N_593);
nor U1963 (N_1963,N_974,N_333);
or U1964 (N_1964,N_892,N_244);
nand U1965 (N_1965,N_378,N_544);
nand U1966 (N_1966,N_802,N_738);
or U1967 (N_1967,N_826,N_740);
or U1968 (N_1968,N_361,N_205);
and U1969 (N_1969,N_708,N_105);
nand U1970 (N_1970,N_343,N_454);
or U1971 (N_1971,N_924,N_842);
xor U1972 (N_1972,N_340,N_758);
and U1973 (N_1973,N_192,N_439);
nand U1974 (N_1974,N_346,N_874);
xnor U1975 (N_1975,N_826,N_61);
nor U1976 (N_1976,N_729,N_188);
nor U1977 (N_1977,N_921,N_78);
nor U1978 (N_1978,N_848,N_814);
xor U1979 (N_1979,N_189,N_471);
or U1980 (N_1980,N_776,N_811);
xor U1981 (N_1981,N_912,N_575);
nand U1982 (N_1982,N_29,N_28);
or U1983 (N_1983,N_482,N_839);
and U1984 (N_1984,N_978,N_333);
nor U1985 (N_1985,N_680,N_118);
xor U1986 (N_1986,N_782,N_804);
or U1987 (N_1987,N_961,N_926);
nand U1988 (N_1988,N_580,N_702);
xor U1989 (N_1989,N_479,N_988);
nand U1990 (N_1990,N_946,N_195);
and U1991 (N_1991,N_200,N_345);
or U1992 (N_1992,N_861,N_890);
nand U1993 (N_1993,N_556,N_929);
nor U1994 (N_1994,N_596,N_82);
or U1995 (N_1995,N_503,N_489);
nor U1996 (N_1996,N_500,N_294);
nand U1997 (N_1997,N_784,N_669);
nor U1998 (N_1998,N_524,N_654);
nor U1999 (N_1999,N_706,N_995);
or U2000 (N_2000,N_1586,N_1314);
nor U2001 (N_2001,N_1000,N_1342);
xor U2002 (N_2002,N_1644,N_1281);
nor U2003 (N_2003,N_1002,N_1946);
nor U2004 (N_2004,N_1578,N_1435);
nand U2005 (N_2005,N_1358,N_1369);
nand U2006 (N_2006,N_1088,N_1080);
nor U2007 (N_2007,N_1001,N_1013);
nor U2008 (N_2008,N_1187,N_1818);
xor U2009 (N_2009,N_1915,N_1200);
nor U2010 (N_2010,N_1326,N_1964);
nand U2011 (N_2011,N_1635,N_1424);
xor U2012 (N_2012,N_1830,N_1693);
nor U2013 (N_2013,N_1023,N_1202);
nor U2014 (N_2014,N_1348,N_1502);
or U2015 (N_2015,N_1816,N_1735);
and U2016 (N_2016,N_1323,N_1584);
and U2017 (N_2017,N_1163,N_1570);
nand U2018 (N_2018,N_1804,N_1381);
nor U2019 (N_2019,N_1135,N_1351);
nand U2020 (N_2020,N_1188,N_1926);
and U2021 (N_2021,N_1535,N_1919);
nor U2022 (N_2022,N_1506,N_1815);
xor U2023 (N_2023,N_1364,N_1254);
or U2024 (N_2024,N_1030,N_1726);
xnor U2025 (N_2025,N_1451,N_1597);
and U2026 (N_2026,N_1972,N_1923);
and U2027 (N_2027,N_1180,N_1302);
or U2028 (N_2028,N_1654,N_1207);
and U2029 (N_2029,N_1363,N_1712);
xor U2030 (N_2030,N_1691,N_1466);
and U2031 (N_2031,N_1990,N_1474);
nor U2032 (N_2032,N_1718,N_1368);
nor U2033 (N_2033,N_1575,N_1507);
nor U2034 (N_2034,N_1067,N_1995);
or U2035 (N_2035,N_1497,N_1076);
nor U2036 (N_2036,N_1897,N_1929);
nor U2037 (N_2037,N_1702,N_1218);
or U2038 (N_2038,N_1128,N_1925);
nand U2039 (N_2039,N_1111,N_1914);
or U2040 (N_2040,N_1836,N_1296);
xnor U2041 (N_2041,N_1922,N_1489);
xnor U2042 (N_2042,N_1463,N_1063);
or U2043 (N_2043,N_1394,N_1231);
nor U2044 (N_2044,N_1663,N_1630);
and U2045 (N_2045,N_1861,N_1731);
or U2046 (N_2046,N_1796,N_1376);
and U2047 (N_2047,N_1215,N_1638);
xnor U2048 (N_2048,N_1835,N_1641);
or U2049 (N_2049,N_1588,N_1567);
xnor U2050 (N_2050,N_1931,N_1283);
nor U2051 (N_2051,N_1012,N_1725);
xor U2052 (N_2052,N_1869,N_1800);
and U2053 (N_2053,N_1624,N_1059);
xor U2054 (N_2054,N_1060,N_1711);
nor U2055 (N_2055,N_1403,N_1426);
nor U2056 (N_2056,N_1872,N_1477);
and U2057 (N_2057,N_1798,N_1340);
or U2058 (N_2058,N_1015,N_1881);
xor U2059 (N_2059,N_1388,N_1083);
nor U2060 (N_2060,N_1515,N_1958);
or U2061 (N_2061,N_1344,N_1677);
nand U2062 (N_2062,N_1406,N_1255);
nand U2063 (N_2063,N_1096,N_1636);
or U2064 (N_2064,N_1960,N_1849);
nor U2065 (N_2065,N_1189,N_1170);
or U2066 (N_2066,N_1593,N_1320);
xor U2067 (N_2067,N_1680,N_1687);
nor U2068 (N_2068,N_1449,N_1688);
xor U2069 (N_2069,N_1117,N_1829);
nand U2070 (N_2070,N_1970,N_1138);
nand U2071 (N_2071,N_1632,N_1555);
nor U2072 (N_2072,N_1452,N_1405);
or U2073 (N_2073,N_1446,N_1309);
xor U2074 (N_2074,N_1284,N_1674);
nand U2075 (N_2075,N_1757,N_1025);
and U2076 (N_2076,N_1885,N_1679);
nor U2077 (N_2077,N_1606,N_1203);
nand U2078 (N_2078,N_1873,N_1014);
or U2079 (N_2079,N_1476,N_1143);
nor U2080 (N_2080,N_1879,N_1429);
nand U2081 (N_2081,N_1759,N_1459);
and U2082 (N_2082,N_1007,N_1890);
or U2083 (N_2083,N_1949,N_1623);
or U2084 (N_2084,N_1387,N_1736);
or U2085 (N_2085,N_1916,N_1303);
xnor U2086 (N_2086,N_1658,N_1269);
nor U2087 (N_2087,N_1542,N_1602);
and U2088 (N_2088,N_1587,N_1045);
or U2089 (N_2089,N_1647,N_1753);
nand U2090 (N_2090,N_1662,N_1942);
nand U2091 (N_2091,N_1653,N_1582);
and U2092 (N_2092,N_1973,N_1825);
nor U2093 (N_2093,N_1004,N_1617);
and U2094 (N_2094,N_1565,N_1445);
and U2095 (N_2095,N_1159,N_1383);
nor U2096 (N_2096,N_1948,N_1047);
nor U2097 (N_2097,N_1543,N_1036);
nand U2098 (N_2098,N_1402,N_1856);
xor U2099 (N_2099,N_1895,N_1197);
nand U2100 (N_2100,N_1902,N_1907);
xor U2101 (N_2101,N_1029,N_1675);
xor U2102 (N_2102,N_1289,N_1775);
or U2103 (N_2103,N_1758,N_1051);
nor U2104 (N_2104,N_1604,N_1136);
nor U2105 (N_2105,N_1304,N_1749);
xor U2106 (N_2106,N_1470,N_1589);
nor U2107 (N_2107,N_1713,N_1934);
nor U2108 (N_2108,N_1266,N_1954);
or U2109 (N_2109,N_1247,N_1058);
and U2110 (N_2110,N_1892,N_1338);
xnor U2111 (N_2111,N_1720,N_1761);
and U2112 (N_2112,N_1724,N_1290);
nor U2113 (N_2113,N_1386,N_1528);
and U2114 (N_2114,N_1397,N_1114);
or U2115 (N_2115,N_1886,N_1107);
nand U2116 (N_2116,N_1353,N_1104);
nand U2117 (N_2117,N_1992,N_1772);
xor U2118 (N_2118,N_1211,N_1053);
and U2119 (N_2119,N_1837,N_1622);
xor U2120 (N_2120,N_1074,N_1035);
and U2121 (N_2121,N_1300,N_1158);
nand U2122 (N_2122,N_1119,N_1618);
nand U2123 (N_2123,N_1652,N_1840);
nand U2124 (N_2124,N_1657,N_1823);
nand U2125 (N_2125,N_1982,N_1750);
or U2126 (N_2126,N_1410,N_1645);
and U2127 (N_2127,N_1295,N_1969);
nand U2128 (N_2128,N_1493,N_1486);
xor U2129 (N_2129,N_1473,N_1245);
nor U2130 (N_2130,N_1171,N_1105);
nand U2131 (N_2131,N_1611,N_1468);
or U2132 (N_2132,N_1744,N_1172);
nand U2133 (N_2133,N_1722,N_1407);
and U2134 (N_2134,N_1462,N_1723);
or U2135 (N_2135,N_1077,N_1637);
and U2136 (N_2136,N_1971,N_1062);
nand U2137 (N_2137,N_1692,N_1249);
and U2138 (N_2138,N_1102,N_1305);
and U2139 (N_2139,N_1144,N_1975);
or U2140 (N_2140,N_1150,N_1701);
nand U2141 (N_2141,N_1549,N_1317);
or U2142 (N_2142,N_1616,N_1913);
or U2143 (N_2143,N_1766,N_1748);
xnor U2144 (N_2144,N_1838,N_1983);
or U2145 (N_2145,N_1998,N_1437);
xor U2146 (N_2146,N_1086,N_1808);
nand U2147 (N_2147,N_1057,N_1742);
nand U2148 (N_2148,N_1075,N_1959);
or U2149 (N_2149,N_1771,N_1504);
nor U2150 (N_2150,N_1009,N_1087);
nand U2151 (N_2151,N_1793,N_1626);
xnor U2152 (N_2152,N_1167,N_1268);
or U2153 (N_2153,N_1858,N_1994);
or U2154 (N_2154,N_1777,N_1208);
nand U2155 (N_2155,N_1494,N_1439);
nand U2156 (N_2156,N_1380,N_1500);
nand U2157 (N_2157,N_1115,N_1548);
xor U2158 (N_2158,N_1416,N_1017);
or U2159 (N_2159,N_1503,N_1794);
nor U2160 (N_2160,N_1336,N_1235);
and U2161 (N_2161,N_1554,N_1178);
xor U2162 (N_2162,N_1953,N_1374);
xor U2163 (N_2163,N_1517,N_1061);
or U2164 (N_2164,N_1393,N_1870);
nand U2165 (N_2165,N_1252,N_1279);
xor U2166 (N_2166,N_1366,N_1571);
or U2167 (N_2167,N_1887,N_1988);
nand U2168 (N_2168,N_1531,N_1556);
nor U2169 (N_2169,N_1471,N_1475);
or U2170 (N_2170,N_1774,N_1073);
nand U2171 (N_2171,N_1665,N_1454);
nor U2172 (N_2172,N_1193,N_1220);
nand U2173 (N_2173,N_1780,N_1656);
and U2174 (N_2174,N_1776,N_1423);
and U2175 (N_2175,N_1469,N_1993);
and U2176 (N_2176,N_1359,N_1868);
nand U2177 (N_2177,N_1650,N_1118);
nor U2178 (N_2178,N_1299,N_1529);
nand U2179 (N_2179,N_1544,N_1933);
nor U2180 (N_2180,N_1223,N_1884);
nand U2181 (N_2181,N_1401,N_1129);
xnor U2182 (N_2182,N_1275,N_1642);
and U2183 (N_2183,N_1545,N_1109);
and U2184 (N_2184,N_1044,N_1160);
and U2185 (N_2185,N_1259,N_1910);
or U2186 (N_2186,N_1843,N_1018);
and U2187 (N_2187,N_1425,N_1217);
or U2188 (N_2188,N_1669,N_1694);
xor U2189 (N_2189,N_1824,N_1541);
nand U2190 (N_2190,N_1716,N_1989);
nand U2191 (N_2191,N_1501,N_1173);
nor U2192 (N_2192,N_1224,N_1276);
or U2193 (N_2193,N_1746,N_1037);
nor U2194 (N_2194,N_1627,N_1600);
nand U2195 (N_2195,N_1137,N_1799);
or U2196 (N_2196,N_1607,N_1605);
nand U2197 (N_2197,N_1226,N_1041);
nor U2198 (N_2198,N_1003,N_1871);
or U2199 (N_2199,N_1513,N_1999);
nor U2200 (N_2200,N_1801,N_1773);
and U2201 (N_2201,N_1455,N_1537);
and U2202 (N_2202,N_1920,N_1412);
xnor U2203 (N_2203,N_1893,N_1464);
or U2204 (N_2204,N_1390,N_1113);
and U2205 (N_2205,N_1098,N_1272);
xor U2206 (N_2206,N_1956,N_1043);
and U2207 (N_2207,N_1034,N_1768);
nand U2208 (N_2208,N_1832,N_1708);
or U2209 (N_2209,N_1730,N_1700);
nand U2210 (N_2210,N_1262,N_1192);
nand U2211 (N_2211,N_1005,N_1236);
nor U2212 (N_2212,N_1066,N_1696);
nor U2213 (N_2213,N_1293,N_1943);
xnor U2214 (N_2214,N_1332,N_1966);
or U2215 (N_2215,N_1559,N_1698);
nand U2216 (N_2216,N_1227,N_1198);
and U2217 (N_2217,N_1442,N_1976);
or U2218 (N_2218,N_1286,N_1924);
nor U2219 (N_2219,N_1078,N_1085);
nand U2220 (N_2220,N_1328,N_1093);
nand U2221 (N_2221,N_1710,N_1448);
nor U2222 (N_2222,N_1027,N_1467);
and U2223 (N_2223,N_1530,N_1209);
or U2224 (N_2224,N_1154,N_1450);
xor U2225 (N_2225,N_1590,N_1151);
or U2226 (N_2226,N_1951,N_1557);
xor U2227 (N_2227,N_1755,N_1081);
and U2228 (N_2228,N_1182,N_1979);
nor U2229 (N_2229,N_1146,N_1148);
nand U2230 (N_2230,N_1094,N_1905);
and U2231 (N_2231,N_1620,N_1056);
and U2232 (N_2232,N_1024,N_1697);
nand U2233 (N_2233,N_1360,N_1125);
and U2234 (N_2234,N_1633,N_1514);
nor U2235 (N_2235,N_1882,N_1789);
nand U2236 (N_2236,N_1329,N_1149);
or U2237 (N_2237,N_1572,N_1228);
nand U2238 (N_2238,N_1496,N_1261);
or U2239 (N_2239,N_1860,N_1715);
xor U2240 (N_2240,N_1516,N_1655);
nand U2241 (N_2241,N_1996,N_1327);
nand U2242 (N_2242,N_1909,N_1977);
nor U2243 (N_2243,N_1727,N_1846);
nand U2244 (N_2244,N_1048,N_1912);
nand U2245 (N_2245,N_1532,N_1256);
or U2246 (N_2246,N_1760,N_1404);
or U2247 (N_2247,N_1398,N_1222);
nor U2248 (N_2248,N_1985,N_1097);
or U2249 (N_2249,N_1330,N_1482);
nor U2250 (N_2250,N_1661,N_1273);
or U2251 (N_2251,N_1225,N_1229);
and U2252 (N_2252,N_1240,N_1945);
and U2253 (N_2253,N_1569,N_1221);
or U2254 (N_2254,N_1857,N_1016);
nand U2255 (N_2255,N_1518,N_1684);
nand U2256 (N_2256,N_1123,N_1553);
or U2257 (N_2257,N_1490,N_1560);
nand U2258 (N_2258,N_1291,N_1010);
xnor U2259 (N_2259,N_1441,N_1277);
or U2260 (N_2260,N_1084,N_1333);
nand U2261 (N_2261,N_1349,N_1312);
xor U2262 (N_2262,N_1596,N_1997);
xnor U2263 (N_2263,N_1288,N_1643);
or U2264 (N_2264,N_1049,N_1629);
and U2265 (N_2265,N_1512,N_1831);
xor U2266 (N_2266,N_1903,N_1161);
or U2267 (N_2267,N_1282,N_1628);
nor U2268 (N_2268,N_1558,N_1659);
and U2269 (N_2269,N_1899,N_1765);
or U2270 (N_2270,N_1522,N_1216);
or U2271 (N_2271,N_1510,N_1298);
and U2272 (N_2272,N_1134,N_1311);
or U2273 (N_2273,N_1592,N_1438);
nor U2274 (N_2274,N_1784,N_1008);
or U2275 (N_2275,N_1099,N_1365);
xnor U2276 (N_2276,N_1705,N_1511);
and U2277 (N_2277,N_1343,N_1483);
nor U2278 (N_2278,N_1239,N_1599);
xnor U2279 (N_2279,N_1373,N_1585);
nor U2280 (N_2280,N_1420,N_1274);
nand U2281 (N_2281,N_1963,N_1610);
nand U2282 (N_2282,N_1552,N_1769);
nand U2283 (N_2283,N_1709,N_1706);
nand U2284 (N_2284,N_1385,N_1069);
or U2285 (N_2285,N_1867,N_1950);
nor U2286 (N_2286,N_1120,N_1246);
or U2287 (N_2287,N_1938,N_1921);
xor U2288 (N_2288,N_1020,N_1457);
nor U2289 (N_2289,N_1743,N_1244);
nor U2290 (N_2290,N_1265,N_1499);
nor U2291 (N_2291,N_1176,N_1301);
xor U2292 (N_2292,N_1807,N_1667);
or U2293 (N_2293,N_1666,N_1901);
nor U2294 (N_2294,N_1480,N_1573);
nand U2295 (N_2295,N_1196,N_1539);
nor U2296 (N_2296,N_1889,N_1621);
or U2297 (N_2297,N_1714,N_1270);
or U2298 (N_2298,N_1375,N_1140);
and U2299 (N_2299,N_1121,N_1595);
and U2300 (N_2300,N_1377,N_1054);
and U2301 (N_2301,N_1206,N_1853);
or U2302 (N_2302,N_1157,N_1052);
and U2303 (N_2303,N_1795,N_1318);
xnor U2304 (N_2304,N_1527,N_1928);
or U2305 (N_2305,N_1465,N_1619);
and U2306 (N_2306,N_1155,N_1930);
and U2307 (N_2307,N_1417,N_1703);
or U2308 (N_2308,N_1389,N_1767);
and U2309 (N_2309,N_1201,N_1574);
or U2310 (N_2310,N_1370,N_1937);
nor U2311 (N_2311,N_1660,N_1447);
nand U2312 (N_2312,N_1428,N_1790);
xnor U2313 (N_2313,N_1781,N_1354);
nand U2314 (N_2314,N_1022,N_1686);
and U2315 (N_2315,N_1162,N_1952);
and U2316 (N_2316,N_1126,N_1851);
nand U2317 (N_2317,N_1232,N_1936);
and U2318 (N_2318,N_1478,N_1166);
nand U2319 (N_2319,N_1908,N_1649);
or U2320 (N_2320,N_1230,N_1826);
xnor U2321 (N_2321,N_1112,N_1770);
nor U2322 (N_2322,N_1717,N_1028);
or U2323 (N_2323,N_1440,N_1734);
nor U2324 (N_2324,N_1400,N_1689);
nand U2325 (N_2325,N_1891,N_1116);
and U2326 (N_2326,N_1601,N_1763);
nor U2327 (N_2327,N_1285,N_1874);
nand U2328 (N_2328,N_1350,N_1175);
or U2329 (N_2329,N_1615,N_1190);
and U2330 (N_2330,N_1878,N_1681);
xnor U2331 (N_2331,N_1064,N_1839);
nor U2332 (N_2332,N_1568,N_1392);
and U2333 (N_2333,N_1673,N_1443);
nor U2334 (N_2334,N_1820,N_1550);
xnor U2335 (N_2335,N_1719,N_1880);
nand U2336 (N_2336,N_1803,N_1894);
nand U2337 (N_2337,N_1184,N_1263);
nand U2338 (N_2338,N_1614,N_1234);
xor U2339 (N_2339,N_1070,N_1536);
and U2340 (N_2340,N_1357,N_1613);
or U2341 (N_2341,N_1019,N_1651);
or U2342 (N_2342,N_1210,N_1177);
nand U2343 (N_2343,N_1458,N_1699);
xor U2344 (N_2344,N_1127,N_1728);
or U2345 (N_2345,N_1491,N_1855);
or U2346 (N_2346,N_1991,N_1243);
nand U2347 (N_2347,N_1631,N_1183);
or U2348 (N_2348,N_1594,N_1546);
nor U2349 (N_2349,N_1564,N_1310);
nand U2350 (N_2350,N_1174,N_1095);
or U2351 (N_2351,N_1817,N_1740);
nor U2352 (N_2352,N_1384,N_1737);
or U2353 (N_2353,N_1006,N_1100);
nand U2354 (N_2354,N_1785,N_1355);
xnor U2355 (N_2355,N_1509,N_1391);
xor U2356 (N_2356,N_1521,N_1371);
nand U2357 (N_2357,N_1453,N_1292);
and U2358 (N_2358,N_1822,N_1212);
and U2359 (N_2359,N_1181,N_1538);
nor U2360 (N_2360,N_1257,N_1779);
xor U2361 (N_2361,N_1347,N_1186);
nor U2362 (N_2362,N_1813,N_1850);
or U2363 (N_2363,N_1888,N_1050);
and U2364 (N_2364,N_1356,N_1248);
nand U2365 (N_2365,N_1382,N_1540);
or U2366 (N_2366,N_1409,N_1091);
or U2367 (N_2367,N_1747,N_1864);
and U2368 (N_2368,N_1828,N_1788);
or U2369 (N_2369,N_1414,N_1124);
nand U2370 (N_2370,N_1579,N_1898);
or U2371 (N_2371,N_1133,N_1152);
or U2372 (N_2372,N_1046,N_1561);
or U2373 (N_2373,N_1092,N_1704);
nor U2374 (N_2374,N_1110,N_1955);
xnor U2375 (N_2375,N_1754,N_1169);
xor U2376 (N_2376,N_1238,N_1947);
or U2377 (N_2377,N_1233,N_1812);
or U2378 (N_2378,N_1806,N_1101);
nand U2379 (N_2379,N_1130,N_1676);
nor U2380 (N_2380,N_1859,N_1191);
xnor U2381 (N_2381,N_1313,N_1819);
or U2382 (N_2382,N_1419,N_1325);
nor U2383 (N_2383,N_1346,N_1646);
xnor U2384 (N_2384,N_1562,N_1738);
nand U2385 (N_2385,N_1865,N_1141);
nor U2386 (N_2386,N_1707,N_1981);
or U2387 (N_2387,N_1508,N_1762);
or U2388 (N_2388,N_1576,N_1786);
or U2389 (N_2389,N_1852,N_1845);
nor U2390 (N_2390,N_1103,N_1145);
nor U2391 (N_2391,N_1042,N_1844);
nand U2392 (N_2392,N_1219,N_1783);
nand U2393 (N_2393,N_1978,N_1566);
nor U2394 (N_2394,N_1460,N_1917);
nor U2395 (N_2395,N_1598,N_1577);
nor U2396 (N_2396,N_1732,N_1782);
and U2397 (N_2397,N_1413,N_1962);
and U2398 (N_2398,N_1682,N_1827);
or U2399 (N_2399,N_1911,N_1258);
and U2400 (N_2400,N_1751,N_1854);
nor U2401 (N_2401,N_1608,N_1065);
nor U2402 (N_2402,N_1011,N_1433);
nand U2403 (N_2403,N_1833,N_1213);
nand U2404 (N_2404,N_1487,N_1372);
xnor U2405 (N_2405,N_1927,N_1287);
nor U2406 (N_2406,N_1436,N_1523);
nor U2407 (N_2407,N_1307,N_1683);
or U2408 (N_2408,N_1791,N_1408);
or U2409 (N_2409,N_1179,N_1308);
nand U2410 (N_2410,N_1316,N_1935);
or U2411 (N_2411,N_1671,N_1253);
or U2412 (N_2412,N_1805,N_1315);
nor U2413 (N_2413,N_1421,N_1205);
xnor U2414 (N_2414,N_1362,N_1980);
xor U2415 (N_2415,N_1153,N_1339);
and U2416 (N_2416,N_1814,N_1108);
or U2417 (N_2417,N_1668,N_1896);
and U2418 (N_2418,N_1481,N_1237);
and U2419 (N_2419,N_1739,N_1877);
nor U2420 (N_2420,N_1974,N_1147);
and U2421 (N_2421,N_1271,N_1640);
and U2422 (N_2422,N_1670,N_1484);
or U2423 (N_2423,N_1488,N_1106);
nand U2424 (N_2424,N_1378,N_1089);
or U2425 (N_2425,N_1957,N_1031);
and U2426 (N_2426,N_1625,N_1581);
or U2427 (N_2427,N_1764,N_1241);
nand U2428 (N_2428,N_1583,N_1431);
nor U2429 (N_2429,N_1547,N_1194);
nand U2430 (N_2430,N_1379,N_1906);
xor U2431 (N_2431,N_1809,N_1242);
or U2432 (N_2432,N_1866,N_1164);
or U2433 (N_2433,N_1741,N_1396);
and U2434 (N_2434,N_1361,N_1399);
nor U2435 (N_2435,N_1634,N_1729);
and U2436 (N_2436,N_1664,N_1341);
nor U2437 (N_2437,N_1883,N_1944);
nand U2438 (N_2438,N_1519,N_1648);
or U2439 (N_2439,N_1260,N_1422);
and U2440 (N_2440,N_1294,N_1032);
nor U2441 (N_2441,N_1337,N_1987);
nor U2442 (N_2442,N_1778,N_1082);
nand U2443 (N_2443,N_1940,N_1068);
or U2444 (N_2444,N_1609,N_1297);
or U2445 (N_2445,N_1461,N_1132);
nor U2446 (N_2446,N_1168,N_1802);
or U2447 (N_2447,N_1456,N_1427);
and U2448 (N_2448,N_1352,N_1904);
and U2449 (N_2449,N_1472,N_1033);
and U2450 (N_2450,N_1411,N_1038);
nand U2451 (N_2451,N_1863,N_1444);
and U2452 (N_2452,N_1185,N_1842);
xnor U2453 (N_2453,N_1334,N_1485);
and U2454 (N_2454,N_1165,N_1479);
xor U2455 (N_2455,N_1331,N_1672);
nor U2456 (N_2456,N_1685,N_1841);
nor U2457 (N_2457,N_1967,N_1072);
and U2458 (N_2458,N_1591,N_1278);
and U2459 (N_2459,N_1695,N_1321);
xnor U2460 (N_2460,N_1524,N_1199);
xnor U2461 (N_2461,N_1345,N_1322);
xor U2462 (N_2462,N_1900,N_1214);
or U2463 (N_2463,N_1026,N_1195);
and U2464 (N_2464,N_1811,N_1721);
or U2465 (N_2465,N_1418,N_1678);
nor U2466 (N_2466,N_1319,N_1984);
xor U2467 (N_2467,N_1251,N_1862);
and U2468 (N_2468,N_1055,N_1834);
and U2469 (N_2469,N_1495,N_1432);
or U2470 (N_2470,N_1079,N_1821);
nor U2471 (N_2471,N_1324,N_1876);
xnor U2472 (N_2472,N_1918,N_1071);
nor U2473 (N_2473,N_1264,N_1520);
nor U2474 (N_2474,N_1250,N_1787);
nor U2475 (N_2475,N_1810,N_1395);
xnor U2476 (N_2476,N_1280,N_1122);
or U2477 (N_2477,N_1142,N_1756);
and U2478 (N_2478,N_1965,N_1752);
or U2479 (N_2479,N_1939,N_1430);
or U2480 (N_2480,N_1986,N_1090);
nor U2481 (N_2481,N_1434,N_1792);
nor U2482 (N_2482,N_1335,N_1961);
or U2483 (N_2483,N_1505,N_1267);
nand U2484 (N_2484,N_1690,N_1131);
xnor U2485 (N_2485,N_1551,N_1797);
nand U2486 (N_2486,N_1875,N_1040);
nor U2487 (N_2487,N_1533,N_1968);
xor U2488 (N_2488,N_1745,N_1367);
nand U2489 (N_2489,N_1021,N_1492);
xor U2490 (N_2490,N_1039,N_1733);
xor U2491 (N_2491,N_1156,N_1534);
or U2492 (N_2492,N_1306,N_1848);
or U2493 (N_2493,N_1932,N_1139);
nand U2494 (N_2494,N_1941,N_1525);
nor U2495 (N_2495,N_1204,N_1526);
nand U2496 (N_2496,N_1498,N_1563);
nor U2497 (N_2497,N_1639,N_1580);
or U2498 (N_2498,N_1612,N_1603);
or U2499 (N_2499,N_1847,N_1415);
nand U2500 (N_2500,N_1527,N_1382);
and U2501 (N_2501,N_1480,N_1599);
nand U2502 (N_2502,N_1321,N_1072);
and U2503 (N_2503,N_1884,N_1449);
xor U2504 (N_2504,N_1857,N_1646);
and U2505 (N_2505,N_1855,N_1377);
and U2506 (N_2506,N_1194,N_1441);
and U2507 (N_2507,N_1226,N_1085);
or U2508 (N_2508,N_1461,N_1680);
xnor U2509 (N_2509,N_1019,N_1702);
nor U2510 (N_2510,N_1418,N_1785);
or U2511 (N_2511,N_1122,N_1582);
and U2512 (N_2512,N_1529,N_1667);
or U2513 (N_2513,N_1985,N_1629);
nor U2514 (N_2514,N_1779,N_1672);
nor U2515 (N_2515,N_1194,N_1505);
or U2516 (N_2516,N_1950,N_1057);
and U2517 (N_2517,N_1227,N_1489);
nor U2518 (N_2518,N_1340,N_1274);
xor U2519 (N_2519,N_1503,N_1242);
and U2520 (N_2520,N_1950,N_1271);
or U2521 (N_2521,N_1338,N_1054);
nand U2522 (N_2522,N_1463,N_1076);
nor U2523 (N_2523,N_1936,N_1019);
nor U2524 (N_2524,N_1720,N_1471);
nor U2525 (N_2525,N_1646,N_1540);
xor U2526 (N_2526,N_1346,N_1058);
and U2527 (N_2527,N_1847,N_1836);
nand U2528 (N_2528,N_1103,N_1813);
xnor U2529 (N_2529,N_1148,N_1304);
or U2530 (N_2530,N_1207,N_1563);
and U2531 (N_2531,N_1632,N_1369);
nor U2532 (N_2532,N_1512,N_1875);
nor U2533 (N_2533,N_1288,N_1298);
nand U2534 (N_2534,N_1872,N_1836);
or U2535 (N_2535,N_1458,N_1682);
and U2536 (N_2536,N_1549,N_1817);
and U2537 (N_2537,N_1030,N_1221);
and U2538 (N_2538,N_1812,N_1360);
nand U2539 (N_2539,N_1987,N_1110);
nand U2540 (N_2540,N_1741,N_1093);
and U2541 (N_2541,N_1737,N_1838);
and U2542 (N_2542,N_1904,N_1946);
xor U2543 (N_2543,N_1506,N_1914);
or U2544 (N_2544,N_1498,N_1751);
and U2545 (N_2545,N_1652,N_1748);
xor U2546 (N_2546,N_1263,N_1388);
and U2547 (N_2547,N_1341,N_1655);
nand U2548 (N_2548,N_1305,N_1468);
nor U2549 (N_2549,N_1988,N_1338);
xor U2550 (N_2550,N_1937,N_1150);
and U2551 (N_2551,N_1159,N_1262);
nand U2552 (N_2552,N_1670,N_1809);
nand U2553 (N_2553,N_1877,N_1184);
and U2554 (N_2554,N_1759,N_1498);
or U2555 (N_2555,N_1083,N_1549);
or U2556 (N_2556,N_1977,N_1777);
nand U2557 (N_2557,N_1319,N_1554);
xnor U2558 (N_2558,N_1260,N_1229);
nand U2559 (N_2559,N_1031,N_1338);
and U2560 (N_2560,N_1357,N_1130);
or U2561 (N_2561,N_1698,N_1959);
or U2562 (N_2562,N_1521,N_1610);
nand U2563 (N_2563,N_1134,N_1907);
xnor U2564 (N_2564,N_1428,N_1548);
nand U2565 (N_2565,N_1705,N_1399);
nand U2566 (N_2566,N_1370,N_1588);
xor U2567 (N_2567,N_1775,N_1102);
nand U2568 (N_2568,N_1079,N_1034);
and U2569 (N_2569,N_1974,N_1275);
xnor U2570 (N_2570,N_1480,N_1741);
and U2571 (N_2571,N_1261,N_1308);
or U2572 (N_2572,N_1616,N_1160);
xnor U2573 (N_2573,N_1499,N_1326);
nor U2574 (N_2574,N_1348,N_1870);
or U2575 (N_2575,N_1810,N_1208);
xnor U2576 (N_2576,N_1498,N_1399);
xor U2577 (N_2577,N_1939,N_1145);
or U2578 (N_2578,N_1636,N_1128);
xor U2579 (N_2579,N_1067,N_1749);
nor U2580 (N_2580,N_1337,N_1022);
and U2581 (N_2581,N_1041,N_1673);
and U2582 (N_2582,N_1633,N_1890);
xor U2583 (N_2583,N_1873,N_1987);
nor U2584 (N_2584,N_1353,N_1291);
xor U2585 (N_2585,N_1787,N_1368);
xor U2586 (N_2586,N_1921,N_1467);
xnor U2587 (N_2587,N_1128,N_1521);
nor U2588 (N_2588,N_1728,N_1672);
xnor U2589 (N_2589,N_1048,N_1728);
and U2590 (N_2590,N_1805,N_1602);
xor U2591 (N_2591,N_1365,N_1327);
nor U2592 (N_2592,N_1464,N_1940);
xnor U2593 (N_2593,N_1042,N_1153);
or U2594 (N_2594,N_1201,N_1811);
nand U2595 (N_2595,N_1987,N_1004);
xnor U2596 (N_2596,N_1622,N_1755);
nand U2597 (N_2597,N_1283,N_1336);
nor U2598 (N_2598,N_1007,N_1215);
nand U2599 (N_2599,N_1139,N_1037);
nor U2600 (N_2600,N_1619,N_1530);
nor U2601 (N_2601,N_1347,N_1029);
nor U2602 (N_2602,N_1316,N_1178);
or U2603 (N_2603,N_1603,N_1617);
nor U2604 (N_2604,N_1360,N_1527);
xor U2605 (N_2605,N_1228,N_1972);
or U2606 (N_2606,N_1651,N_1702);
nand U2607 (N_2607,N_1563,N_1616);
or U2608 (N_2608,N_1506,N_1820);
nand U2609 (N_2609,N_1749,N_1547);
nand U2610 (N_2610,N_1475,N_1504);
and U2611 (N_2611,N_1390,N_1118);
nand U2612 (N_2612,N_1968,N_1183);
xnor U2613 (N_2613,N_1617,N_1781);
or U2614 (N_2614,N_1960,N_1989);
and U2615 (N_2615,N_1455,N_1442);
and U2616 (N_2616,N_1018,N_1670);
nor U2617 (N_2617,N_1591,N_1360);
nand U2618 (N_2618,N_1210,N_1720);
or U2619 (N_2619,N_1388,N_1929);
and U2620 (N_2620,N_1640,N_1830);
and U2621 (N_2621,N_1019,N_1134);
nor U2622 (N_2622,N_1540,N_1847);
and U2623 (N_2623,N_1523,N_1085);
xnor U2624 (N_2624,N_1447,N_1351);
or U2625 (N_2625,N_1315,N_1811);
or U2626 (N_2626,N_1200,N_1638);
nor U2627 (N_2627,N_1369,N_1149);
xnor U2628 (N_2628,N_1115,N_1695);
or U2629 (N_2629,N_1297,N_1909);
or U2630 (N_2630,N_1172,N_1722);
xor U2631 (N_2631,N_1659,N_1922);
xnor U2632 (N_2632,N_1694,N_1516);
or U2633 (N_2633,N_1364,N_1749);
nor U2634 (N_2634,N_1326,N_1311);
nand U2635 (N_2635,N_1427,N_1320);
or U2636 (N_2636,N_1252,N_1377);
nand U2637 (N_2637,N_1658,N_1641);
nand U2638 (N_2638,N_1975,N_1669);
nor U2639 (N_2639,N_1844,N_1474);
xor U2640 (N_2640,N_1932,N_1252);
nor U2641 (N_2641,N_1205,N_1087);
or U2642 (N_2642,N_1846,N_1280);
or U2643 (N_2643,N_1181,N_1652);
nand U2644 (N_2644,N_1346,N_1191);
xor U2645 (N_2645,N_1030,N_1971);
and U2646 (N_2646,N_1783,N_1525);
and U2647 (N_2647,N_1219,N_1916);
or U2648 (N_2648,N_1513,N_1605);
nand U2649 (N_2649,N_1392,N_1448);
or U2650 (N_2650,N_1536,N_1565);
nor U2651 (N_2651,N_1874,N_1827);
nor U2652 (N_2652,N_1118,N_1369);
nand U2653 (N_2653,N_1158,N_1177);
xnor U2654 (N_2654,N_1189,N_1989);
nand U2655 (N_2655,N_1897,N_1520);
and U2656 (N_2656,N_1531,N_1079);
nor U2657 (N_2657,N_1037,N_1482);
nor U2658 (N_2658,N_1954,N_1064);
nor U2659 (N_2659,N_1044,N_1066);
nand U2660 (N_2660,N_1525,N_1511);
nand U2661 (N_2661,N_1236,N_1647);
nand U2662 (N_2662,N_1178,N_1818);
nor U2663 (N_2663,N_1077,N_1507);
or U2664 (N_2664,N_1274,N_1384);
xor U2665 (N_2665,N_1755,N_1627);
or U2666 (N_2666,N_1280,N_1220);
nor U2667 (N_2667,N_1111,N_1476);
nand U2668 (N_2668,N_1442,N_1658);
xnor U2669 (N_2669,N_1829,N_1907);
and U2670 (N_2670,N_1395,N_1309);
nor U2671 (N_2671,N_1474,N_1307);
nand U2672 (N_2672,N_1080,N_1010);
nor U2673 (N_2673,N_1815,N_1229);
and U2674 (N_2674,N_1218,N_1534);
nor U2675 (N_2675,N_1593,N_1717);
or U2676 (N_2676,N_1919,N_1585);
nand U2677 (N_2677,N_1546,N_1254);
and U2678 (N_2678,N_1933,N_1367);
nor U2679 (N_2679,N_1846,N_1343);
xnor U2680 (N_2680,N_1359,N_1213);
xnor U2681 (N_2681,N_1733,N_1429);
nand U2682 (N_2682,N_1153,N_1166);
nor U2683 (N_2683,N_1288,N_1046);
or U2684 (N_2684,N_1993,N_1666);
xor U2685 (N_2685,N_1276,N_1447);
nand U2686 (N_2686,N_1053,N_1606);
or U2687 (N_2687,N_1181,N_1777);
nand U2688 (N_2688,N_1762,N_1836);
nand U2689 (N_2689,N_1710,N_1935);
or U2690 (N_2690,N_1908,N_1171);
nor U2691 (N_2691,N_1024,N_1363);
nand U2692 (N_2692,N_1347,N_1419);
and U2693 (N_2693,N_1579,N_1243);
or U2694 (N_2694,N_1644,N_1784);
xnor U2695 (N_2695,N_1534,N_1079);
xnor U2696 (N_2696,N_1084,N_1527);
and U2697 (N_2697,N_1491,N_1000);
xnor U2698 (N_2698,N_1784,N_1456);
and U2699 (N_2699,N_1777,N_1241);
or U2700 (N_2700,N_1674,N_1626);
or U2701 (N_2701,N_1082,N_1392);
and U2702 (N_2702,N_1798,N_1879);
or U2703 (N_2703,N_1020,N_1248);
and U2704 (N_2704,N_1137,N_1630);
nor U2705 (N_2705,N_1061,N_1635);
xor U2706 (N_2706,N_1906,N_1787);
xor U2707 (N_2707,N_1657,N_1925);
and U2708 (N_2708,N_1683,N_1349);
nor U2709 (N_2709,N_1833,N_1104);
nor U2710 (N_2710,N_1486,N_1506);
and U2711 (N_2711,N_1920,N_1197);
xor U2712 (N_2712,N_1138,N_1258);
nor U2713 (N_2713,N_1172,N_1573);
nor U2714 (N_2714,N_1045,N_1249);
xnor U2715 (N_2715,N_1406,N_1507);
or U2716 (N_2716,N_1812,N_1939);
nor U2717 (N_2717,N_1303,N_1907);
or U2718 (N_2718,N_1347,N_1190);
nand U2719 (N_2719,N_1124,N_1936);
nor U2720 (N_2720,N_1169,N_1678);
nand U2721 (N_2721,N_1742,N_1574);
and U2722 (N_2722,N_1096,N_1498);
nor U2723 (N_2723,N_1449,N_1074);
nand U2724 (N_2724,N_1541,N_1075);
nand U2725 (N_2725,N_1125,N_1696);
xor U2726 (N_2726,N_1856,N_1567);
nand U2727 (N_2727,N_1168,N_1907);
or U2728 (N_2728,N_1792,N_1136);
xnor U2729 (N_2729,N_1088,N_1682);
nor U2730 (N_2730,N_1442,N_1250);
and U2731 (N_2731,N_1749,N_1543);
xor U2732 (N_2732,N_1096,N_1190);
nor U2733 (N_2733,N_1033,N_1286);
nand U2734 (N_2734,N_1112,N_1238);
nor U2735 (N_2735,N_1413,N_1645);
nand U2736 (N_2736,N_1769,N_1598);
and U2737 (N_2737,N_1565,N_1204);
and U2738 (N_2738,N_1652,N_1097);
nand U2739 (N_2739,N_1556,N_1540);
or U2740 (N_2740,N_1663,N_1225);
nor U2741 (N_2741,N_1558,N_1535);
xor U2742 (N_2742,N_1902,N_1178);
nor U2743 (N_2743,N_1847,N_1406);
nand U2744 (N_2744,N_1505,N_1588);
nor U2745 (N_2745,N_1904,N_1363);
or U2746 (N_2746,N_1935,N_1983);
xnor U2747 (N_2747,N_1466,N_1786);
nor U2748 (N_2748,N_1069,N_1516);
and U2749 (N_2749,N_1683,N_1547);
or U2750 (N_2750,N_1711,N_1432);
or U2751 (N_2751,N_1871,N_1357);
nor U2752 (N_2752,N_1959,N_1099);
or U2753 (N_2753,N_1257,N_1834);
nor U2754 (N_2754,N_1637,N_1945);
xnor U2755 (N_2755,N_1608,N_1353);
nor U2756 (N_2756,N_1227,N_1484);
nor U2757 (N_2757,N_1424,N_1055);
xnor U2758 (N_2758,N_1347,N_1899);
or U2759 (N_2759,N_1591,N_1903);
or U2760 (N_2760,N_1053,N_1681);
and U2761 (N_2761,N_1290,N_1805);
and U2762 (N_2762,N_1874,N_1489);
nand U2763 (N_2763,N_1705,N_1397);
xor U2764 (N_2764,N_1767,N_1038);
or U2765 (N_2765,N_1100,N_1047);
or U2766 (N_2766,N_1970,N_1377);
or U2767 (N_2767,N_1911,N_1596);
xnor U2768 (N_2768,N_1028,N_1616);
xnor U2769 (N_2769,N_1543,N_1201);
xnor U2770 (N_2770,N_1339,N_1218);
and U2771 (N_2771,N_1389,N_1963);
xor U2772 (N_2772,N_1568,N_1709);
or U2773 (N_2773,N_1491,N_1592);
nand U2774 (N_2774,N_1329,N_1998);
and U2775 (N_2775,N_1566,N_1581);
nand U2776 (N_2776,N_1508,N_1321);
nor U2777 (N_2777,N_1844,N_1373);
or U2778 (N_2778,N_1684,N_1570);
or U2779 (N_2779,N_1039,N_1969);
xor U2780 (N_2780,N_1033,N_1020);
xor U2781 (N_2781,N_1710,N_1042);
or U2782 (N_2782,N_1675,N_1883);
nand U2783 (N_2783,N_1067,N_1864);
nor U2784 (N_2784,N_1510,N_1091);
and U2785 (N_2785,N_1330,N_1858);
or U2786 (N_2786,N_1850,N_1589);
xnor U2787 (N_2787,N_1100,N_1126);
nand U2788 (N_2788,N_1987,N_1432);
nor U2789 (N_2789,N_1139,N_1323);
and U2790 (N_2790,N_1823,N_1973);
nand U2791 (N_2791,N_1599,N_1477);
and U2792 (N_2792,N_1912,N_1254);
and U2793 (N_2793,N_1155,N_1591);
nor U2794 (N_2794,N_1023,N_1924);
nor U2795 (N_2795,N_1333,N_1775);
nand U2796 (N_2796,N_1662,N_1488);
nand U2797 (N_2797,N_1102,N_1860);
or U2798 (N_2798,N_1147,N_1886);
or U2799 (N_2799,N_1952,N_1815);
xnor U2800 (N_2800,N_1525,N_1368);
xor U2801 (N_2801,N_1284,N_1372);
nand U2802 (N_2802,N_1397,N_1625);
or U2803 (N_2803,N_1879,N_1679);
xor U2804 (N_2804,N_1491,N_1103);
nor U2805 (N_2805,N_1601,N_1345);
and U2806 (N_2806,N_1354,N_1139);
and U2807 (N_2807,N_1755,N_1271);
nor U2808 (N_2808,N_1171,N_1148);
nand U2809 (N_2809,N_1247,N_1835);
and U2810 (N_2810,N_1756,N_1874);
or U2811 (N_2811,N_1880,N_1547);
and U2812 (N_2812,N_1772,N_1848);
nor U2813 (N_2813,N_1638,N_1737);
or U2814 (N_2814,N_1129,N_1752);
nand U2815 (N_2815,N_1245,N_1571);
and U2816 (N_2816,N_1505,N_1865);
or U2817 (N_2817,N_1063,N_1621);
or U2818 (N_2818,N_1612,N_1494);
xnor U2819 (N_2819,N_1739,N_1430);
nand U2820 (N_2820,N_1539,N_1474);
nand U2821 (N_2821,N_1125,N_1018);
or U2822 (N_2822,N_1850,N_1545);
nor U2823 (N_2823,N_1816,N_1940);
or U2824 (N_2824,N_1116,N_1249);
nand U2825 (N_2825,N_1669,N_1643);
xor U2826 (N_2826,N_1642,N_1254);
and U2827 (N_2827,N_1952,N_1989);
xor U2828 (N_2828,N_1745,N_1074);
or U2829 (N_2829,N_1090,N_1312);
or U2830 (N_2830,N_1998,N_1537);
xnor U2831 (N_2831,N_1137,N_1649);
nor U2832 (N_2832,N_1381,N_1810);
and U2833 (N_2833,N_1063,N_1406);
nand U2834 (N_2834,N_1666,N_1842);
or U2835 (N_2835,N_1343,N_1679);
xnor U2836 (N_2836,N_1390,N_1095);
nand U2837 (N_2837,N_1881,N_1408);
nor U2838 (N_2838,N_1780,N_1418);
nor U2839 (N_2839,N_1249,N_1659);
or U2840 (N_2840,N_1741,N_1432);
and U2841 (N_2841,N_1560,N_1425);
nor U2842 (N_2842,N_1716,N_1254);
nor U2843 (N_2843,N_1601,N_1093);
nor U2844 (N_2844,N_1614,N_1981);
or U2845 (N_2845,N_1519,N_1824);
and U2846 (N_2846,N_1385,N_1700);
xnor U2847 (N_2847,N_1901,N_1904);
nand U2848 (N_2848,N_1831,N_1565);
nand U2849 (N_2849,N_1587,N_1116);
and U2850 (N_2850,N_1558,N_1287);
or U2851 (N_2851,N_1884,N_1978);
and U2852 (N_2852,N_1748,N_1854);
nor U2853 (N_2853,N_1124,N_1437);
xor U2854 (N_2854,N_1255,N_1628);
xor U2855 (N_2855,N_1922,N_1203);
xnor U2856 (N_2856,N_1860,N_1844);
or U2857 (N_2857,N_1694,N_1478);
nand U2858 (N_2858,N_1800,N_1318);
nand U2859 (N_2859,N_1132,N_1919);
xor U2860 (N_2860,N_1038,N_1347);
or U2861 (N_2861,N_1674,N_1499);
xnor U2862 (N_2862,N_1861,N_1042);
nor U2863 (N_2863,N_1725,N_1722);
xor U2864 (N_2864,N_1483,N_1045);
nand U2865 (N_2865,N_1977,N_1939);
nor U2866 (N_2866,N_1338,N_1070);
xnor U2867 (N_2867,N_1604,N_1292);
nor U2868 (N_2868,N_1580,N_1030);
nand U2869 (N_2869,N_1524,N_1247);
xnor U2870 (N_2870,N_1713,N_1832);
nor U2871 (N_2871,N_1638,N_1004);
or U2872 (N_2872,N_1901,N_1706);
or U2873 (N_2873,N_1626,N_1338);
and U2874 (N_2874,N_1551,N_1352);
xnor U2875 (N_2875,N_1108,N_1572);
and U2876 (N_2876,N_1625,N_1815);
xor U2877 (N_2877,N_1862,N_1099);
and U2878 (N_2878,N_1160,N_1707);
xnor U2879 (N_2879,N_1323,N_1066);
or U2880 (N_2880,N_1927,N_1086);
xor U2881 (N_2881,N_1083,N_1809);
and U2882 (N_2882,N_1922,N_1830);
xor U2883 (N_2883,N_1185,N_1464);
xor U2884 (N_2884,N_1897,N_1866);
and U2885 (N_2885,N_1986,N_1216);
nand U2886 (N_2886,N_1952,N_1122);
or U2887 (N_2887,N_1953,N_1619);
nand U2888 (N_2888,N_1065,N_1232);
or U2889 (N_2889,N_1310,N_1925);
nor U2890 (N_2890,N_1522,N_1872);
and U2891 (N_2891,N_1866,N_1489);
nand U2892 (N_2892,N_1463,N_1386);
xor U2893 (N_2893,N_1553,N_1188);
xnor U2894 (N_2894,N_1198,N_1898);
or U2895 (N_2895,N_1876,N_1917);
nand U2896 (N_2896,N_1247,N_1556);
or U2897 (N_2897,N_1950,N_1711);
nand U2898 (N_2898,N_1142,N_1464);
and U2899 (N_2899,N_1377,N_1096);
and U2900 (N_2900,N_1410,N_1613);
nand U2901 (N_2901,N_1170,N_1701);
or U2902 (N_2902,N_1132,N_1821);
nand U2903 (N_2903,N_1480,N_1477);
and U2904 (N_2904,N_1781,N_1135);
or U2905 (N_2905,N_1068,N_1686);
and U2906 (N_2906,N_1774,N_1453);
xor U2907 (N_2907,N_1184,N_1246);
nor U2908 (N_2908,N_1538,N_1235);
nand U2909 (N_2909,N_1363,N_1788);
or U2910 (N_2910,N_1391,N_1571);
and U2911 (N_2911,N_1463,N_1801);
xnor U2912 (N_2912,N_1085,N_1375);
nor U2913 (N_2913,N_1519,N_1386);
or U2914 (N_2914,N_1158,N_1755);
nor U2915 (N_2915,N_1601,N_1481);
nand U2916 (N_2916,N_1171,N_1776);
and U2917 (N_2917,N_1580,N_1721);
nand U2918 (N_2918,N_1901,N_1469);
and U2919 (N_2919,N_1940,N_1349);
nor U2920 (N_2920,N_1745,N_1223);
nor U2921 (N_2921,N_1408,N_1699);
nand U2922 (N_2922,N_1954,N_1392);
and U2923 (N_2923,N_1708,N_1075);
and U2924 (N_2924,N_1876,N_1638);
or U2925 (N_2925,N_1521,N_1734);
xnor U2926 (N_2926,N_1481,N_1757);
xnor U2927 (N_2927,N_1082,N_1302);
xor U2928 (N_2928,N_1479,N_1767);
nor U2929 (N_2929,N_1907,N_1761);
nand U2930 (N_2930,N_1799,N_1432);
nand U2931 (N_2931,N_1822,N_1306);
nand U2932 (N_2932,N_1534,N_1727);
nor U2933 (N_2933,N_1350,N_1232);
xnor U2934 (N_2934,N_1040,N_1026);
nor U2935 (N_2935,N_1395,N_1471);
xor U2936 (N_2936,N_1975,N_1019);
or U2937 (N_2937,N_1436,N_1300);
nor U2938 (N_2938,N_1254,N_1115);
or U2939 (N_2939,N_1798,N_1529);
nor U2940 (N_2940,N_1152,N_1170);
or U2941 (N_2941,N_1381,N_1565);
or U2942 (N_2942,N_1239,N_1862);
nand U2943 (N_2943,N_1422,N_1686);
nand U2944 (N_2944,N_1819,N_1531);
nor U2945 (N_2945,N_1548,N_1389);
and U2946 (N_2946,N_1766,N_1266);
or U2947 (N_2947,N_1387,N_1401);
and U2948 (N_2948,N_1978,N_1419);
and U2949 (N_2949,N_1937,N_1215);
nand U2950 (N_2950,N_1576,N_1283);
and U2951 (N_2951,N_1136,N_1672);
nand U2952 (N_2952,N_1702,N_1623);
and U2953 (N_2953,N_1985,N_1671);
xnor U2954 (N_2954,N_1092,N_1579);
xnor U2955 (N_2955,N_1434,N_1341);
xor U2956 (N_2956,N_1355,N_1341);
xnor U2957 (N_2957,N_1221,N_1757);
xnor U2958 (N_2958,N_1878,N_1065);
nor U2959 (N_2959,N_1622,N_1500);
nand U2960 (N_2960,N_1047,N_1085);
nand U2961 (N_2961,N_1775,N_1010);
nor U2962 (N_2962,N_1446,N_1475);
or U2963 (N_2963,N_1555,N_1001);
xnor U2964 (N_2964,N_1865,N_1190);
and U2965 (N_2965,N_1449,N_1098);
nor U2966 (N_2966,N_1987,N_1660);
and U2967 (N_2967,N_1051,N_1190);
nand U2968 (N_2968,N_1721,N_1695);
nand U2969 (N_2969,N_1984,N_1690);
nor U2970 (N_2970,N_1109,N_1847);
and U2971 (N_2971,N_1770,N_1513);
nor U2972 (N_2972,N_1350,N_1910);
and U2973 (N_2973,N_1087,N_1121);
nand U2974 (N_2974,N_1654,N_1158);
nand U2975 (N_2975,N_1579,N_1250);
nor U2976 (N_2976,N_1723,N_1918);
xor U2977 (N_2977,N_1667,N_1677);
or U2978 (N_2978,N_1198,N_1009);
nor U2979 (N_2979,N_1852,N_1600);
nand U2980 (N_2980,N_1103,N_1169);
nor U2981 (N_2981,N_1090,N_1733);
nand U2982 (N_2982,N_1034,N_1877);
nor U2983 (N_2983,N_1679,N_1990);
nor U2984 (N_2984,N_1950,N_1622);
and U2985 (N_2985,N_1072,N_1170);
nand U2986 (N_2986,N_1252,N_1103);
xor U2987 (N_2987,N_1444,N_1490);
or U2988 (N_2988,N_1565,N_1265);
or U2989 (N_2989,N_1166,N_1841);
or U2990 (N_2990,N_1627,N_1793);
or U2991 (N_2991,N_1734,N_1461);
xor U2992 (N_2992,N_1532,N_1723);
and U2993 (N_2993,N_1808,N_1486);
xnor U2994 (N_2994,N_1195,N_1334);
or U2995 (N_2995,N_1352,N_1389);
nand U2996 (N_2996,N_1389,N_1152);
and U2997 (N_2997,N_1158,N_1508);
and U2998 (N_2998,N_1684,N_1077);
and U2999 (N_2999,N_1022,N_1648);
and UO_0 (O_0,N_2544,N_2848);
nand UO_1 (O_1,N_2057,N_2134);
and UO_2 (O_2,N_2071,N_2437);
xnor UO_3 (O_3,N_2809,N_2035);
or UO_4 (O_4,N_2102,N_2395);
nand UO_5 (O_5,N_2937,N_2367);
or UO_6 (O_6,N_2581,N_2323);
and UO_7 (O_7,N_2750,N_2006);
or UO_8 (O_8,N_2267,N_2992);
and UO_9 (O_9,N_2791,N_2608);
nand UO_10 (O_10,N_2115,N_2675);
nand UO_11 (O_11,N_2386,N_2228);
or UO_12 (O_12,N_2986,N_2441);
nand UO_13 (O_13,N_2348,N_2227);
nor UO_14 (O_14,N_2664,N_2201);
nand UO_15 (O_15,N_2210,N_2368);
xor UO_16 (O_16,N_2512,N_2040);
and UO_17 (O_17,N_2967,N_2553);
nor UO_18 (O_18,N_2221,N_2128);
and UO_19 (O_19,N_2351,N_2379);
nor UO_20 (O_20,N_2516,N_2604);
nor UO_21 (O_21,N_2744,N_2823);
and UO_22 (O_22,N_2660,N_2854);
nor UO_23 (O_23,N_2162,N_2981);
xor UO_24 (O_24,N_2794,N_2335);
nand UO_25 (O_25,N_2959,N_2229);
or UO_26 (O_26,N_2277,N_2732);
or UO_27 (O_27,N_2977,N_2887);
nor UO_28 (O_28,N_2763,N_2725);
or UO_29 (O_29,N_2352,N_2853);
and UO_30 (O_30,N_2189,N_2574);
and UO_31 (O_31,N_2956,N_2826);
or UO_32 (O_32,N_2097,N_2421);
xor UO_33 (O_33,N_2394,N_2968);
nor UO_34 (O_34,N_2143,N_2105);
nand UO_35 (O_35,N_2655,N_2139);
nor UO_36 (O_36,N_2947,N_2401);
or UO_37 (O_37,N_2314,N_2775);
xor UO_38 (O_38,N_2007,N_2662);
and UO_39 (O_39,N_2031,N_2244);
xor UO_40 (O_40,N_2813,N_2797);
nor UO_41 (O_41,N_2837,N_2739);
xor UO_42 (O_42,N_2148,N_2643);
nor UO_43 (O_43,N_2987,N_2249);
nand UO_44 (O_44,N_2436,N_2418);
or UO_45 (O_45,N_2788,N_2188);
nand UO_46 (O_46,N_2685,N_2708);
and UO_47 (O_47,N_2173,N_2883);
or UO_48 (O_48,N_2215,N_2142);
nor UO_49 (O_49,N_2601,N_2485);
or UO_50 (O_50,N_2353,N_2336);
nand UO_51 (O_51,N_2058,N_2312);
and UO_52 (O_52,N_2338,N_2690);
xor UO_53 (O_53,N_2478,N_2202);
nand UO_54 (O_54,N_2735,N_2002);
and UO_55 (O_55,N_2181,N_2811);
xnor UO_56 (O_56,N_2941,N_2784);
or UO_57 (O_57,N_2442,N_2546);
or UO_58 (O_58,N_2077,N_2266);
nor UO_59 (O_59,N_2378,N_2587);
xor UO_60 (O_60,N_2480,N_2617);
nor UO_61 (O_61,N_2157,N_2796);
nand UO_62 (O_62,N_2107,N_2344);
or UO_63 (O_63,N_2501,N_2955);
nor UO_64 (O_64,N_2554,N_2108);
and UO_65 (O_65,N_2166,N_2673);
xor UO_66 (O_66,N_2745,N_2785);
nand UO_67 (O_67,N_2817,N_2046);
nor UO_68 (O_68,N_2424,N_2576);
nor UO_69 (O_69,N_2892,N_2905);
nor UO_70 (O_70,N_2078,N_2165);
or UO_71 (O_71,N_2877,N_2779);
xnor UO_72 (O_72,N_2023,N_2524);
and UO_73 (O_73,N_2680,N_2857);
nand UO_74 (O_74,N_2464,N_2993);
nand UO_75 (O_75,N_2384,N_2320);
and UO_76 (O_76,N_2275,N_2702);
xnor UO_77 (O_77,N_2237,N_2907);
nor UO_78 (O_78,N_2559,N_2774);
nor UO_79 (O_79,N_2253,N_2717);
or UO_80 (O_80,N_2677,N_2371);
nor UO_81 (O_81,N_2961,N_2783);
or UO_82 (O_82,N_2593,N_2549);
xnor UO_83 (O_83,N_2646,N_2505);
xor UO_84 (O_84,N_2451,N_2592);
nand UO_85 (O_85,N_2679,N_2220);
nor UO_86 (O_86,N_2532,N_2484);
nor UO_87 (O_87,N_2402,N_2607);
xor UO_88 (O_88,N_2814,N_2771);
nor UO_89 (O_89,N_2276,N_2152);
or UO_90 (O_90,N_2836,N_2610);
nor UO_91 (O_91,N_2649,N_2509);
nand UO_92 (O_92,N_2911,N_2120);
and UO_93 (O_93,N_2503,N_2880);
or UO_94 (O_94,N_2940,N_2493);
nor UO_95 (O_95,N_2316,N_2780);
nor UO_96 (O_96,N_2870,N_2197);
or UO_97 (O_97,N_2294,N_2518);
nor UO_98 (O_98,N_2236,N_2787);
nor UO_99 (O_99,N_2951,N_2869);
nand UO_100 (O_100,N_2766,N_2026);
and UO_101 (O_101,N_2241,N_2557);
xnor UO_102 (O_102,N_2531,N_2710);
and UO_103 (O_103,N_2223,N_2100);
xor UO_104 (O_104,N_2627,N_2900);
nand UO_105 (O_105,N_2109,N_2008);
or UO_106 (O_106,N_2271,N_2547);
and UO_107 (O_107,N_2714,N_2716);
or UO_108 (O_108,N_2431,N_2615);
and UO_109 (O_109,N_2370,N_2663);
or UO_110 (O_110,N_2471,N_2591);
nor UO_111 (O_111,N_2460,N_2399);
xnor UO_112 (O_112,N_2678,N_2828);
nand UO_113 (O_113,N_2552,N_2555);
nor UO_114 (O_114,N_2050,N_2467);
nand UO_115 (O_115,N_2003,N_2313);
nand UO_116 (O_116,N_2667,N_2160);
nand UO_117 (O_117,N_2124,N_2778);
and UO_118 (O_118,N_2706,N_2974);
or UO_119 (O_119,N_2123,N_2170);
nand UO_120 (O_120,N_2133,N_2332);
and UO_121 (O_121,N_2688,N_2825);
nor UO_122 (O_122,N_2930,N_2203);
or UO_123 (O_123,N_2920,N_2965);
xnor UO_124 (O_124,N_2843,N_2789);
or UO_125 (O_125,N_2259,N_2866);
nor UO_126 (O_126,N_2440,N_2328);
nand UO_127 (O_127,N_2758,N_2749);
or UO_128 (O_128,N_2186,N_2948);
and UO_129 (O_129,N_2021,N_2225);
xnor UO_130 (O_130,N_2438,N_2302);
or UO_131 (O_131,N_2863,N_2536);
or UO_132 (O_132,N_2453,N_2723);
or UO_133 (O_133,N_2738,N_2962);
or UO_134 (O_134,N_2747,N_2208);
nor UO_135 (O_135,N_2632,N_2537);
nand UO_136 (O_136,N_2855,N_2268);
nor UO_137 (O_137,N_2497,N_2594);
nand UO_138 (O_138,N_2469,N_2769);
xnor UO_139 (O_139,N_2448,N_2740);
or UO_140 (O_140,N_2751,N_2994);
nor UO_141 (O_141,N_2560,N_2326);
xnor UO_142 (O_142,N_2209,N_2430);
or UO_143 (O_143,N_2178,N_2248);
xnor UO_144 (O_144,N_2207,N_2693);
nand UO_145 (O_145,N_2444,N_2898);
xnor UO_146 (O_146,N_2985,N_2899);
nand UO_147 (O_147,N_2099,N_2342);
xnor UO_148 (O_148,N_2599,N_2017);
nand UO_149 (O_149,N_2807,N_2315);
xnor UO_150 (O_150,N_2199,N_2283);
or UO_151 (O_151,N_2080,N_2952);
nor UO_152 (O_152,N_2988,N_2458);
nand UO_153 (O_153,N_2568,N_2116);
nand UO_154 (O_154,N_2192,N_2647);
nor UO_155 (O_155,N_2297,N_2614);
nand UO_156 (O_156,N_2412,N_2310);
nor UO_157 (O_157,N_2092,N_2770);
xor UO_158 (O_158,N_2629,N_2694);
nand UO_159 (O_159,N_2403,N_2474);
xnor UO_160 (O_160,N_2616,N_2243);
nand UO_161 (O_161,N_2571,N_2895);
and UO_162 (O_162,N_2971,N_2341);
and UO_163 (O_163,N_2047,N_2976);
and UO_164 (O_164,N_2489,N_2175);
xnor UO_165 (O_165,N_2041,N_2978);
nand UO_166 (O_166,N_2079,N_2411);
nand UO_167 (O_167,N_2765,N_2185);
or UO_168 (O_168,N_2292,N_2748);
and UO_169 (O_169,N_2212,N_2681);
and UO_170 (O_170,N_2908,N_2069);
xnor UO_171 (O_171,N_2343,N_2713);
nor UO_172 (O_172,N_2393,N_2004);
nor UO_173 (O_173,N_2942,N_2037);
nor UO_174 (O_174,N_2578,N_2640);
nor UO_175 (O_175,N_2645,N_2269);
xor UO_176 (O_176,N_2762,N_2890);
xor UO_177 (O_177,N_2609,N_2729);
and UO_178 (O_178,N_2226,N_2300);
or UO_179 (O_179,N_2802,N_2874);
and UO_180 (O_180,N_2272,N_2760);
nor UO_181 (O_181,N_2492,N_2076);
nor UO_182 (O_182,N_2915,N_2598);
nand UO_183 (O_183,N_2198,N_2672);
or UO_184 (O_184,N_2818,N_2999);
or UO_185 (O_185,N_2290,N_2149);
nand UO_186 (O_186,N_2051,N_2700);
and UO_187 (O_187,N_2415,N_2439);
or UO_188 (O_188,N_2864,N_2795);
xnor UO_189 (O_189,N_2131,N_2445);
nor UO_190 (O_190,N_2299,N_2801);
or UO_191 (O_191,N_2695,N_2712);
or UO_192 (O_192,N_2768,N_2345);
or UO_193 (O_193,N_2245,N_2205);
xor UO_194 (O_194,N_2580,N_2465);
nor UO_195 (O_195,N_2168,N_2840);
nand UO_196 (O_196,N_2298,N_2112);
nand UO_197 (O_197,N_2325,N_2856);
and UO_198 (O_198,N_2910,N_2586);
nand UO_199 (O_199,N_2846,N_2566);
xor UO_200 (O_200,N_2011,N_2456);
xnor UO_201 (O_201,N_2838,N_2065);
xor UO_202 (O_202,N_2666,N_2096);
nand UO_203 (O_203,N_2287,N_2125);
xor UO_204 (O_204,N_2637,N_2240);
xor UO_205 (O_205,N_2638,N_2180);
nor UO_206 (O_206,N_2603,N_2126);
nor UO_207 (O_207,N_2129,N_2264);
nand UO_208 (O_208,N_2691,N_2319);
nor UO_209 (O_209,N_2921,N_2340);
and UO_210 (O_210,N_2511,N_2155);
and UO_211 (O_211,N_2879,N_2318);
nor UO_212 (O_212,N_2564,N_2958);
nand UO_213 (O_213,N_2251,N_2565);
and UO_214 (O_214,N_2064,N_2377);
nor UO_215 (O_215,N_2039,N_2365);
and UO_216 (O_216,N_2528,N_2285);
and UO_217 (O_217,N_2334,N_2466);
xor UO_218 (O_218,N_2792,N_2432);
xor UO_219 (O_219,N_2522,N_2746);
nor UO_220 (O_220,N_2254,N_2491);
or UO_221 (O_221,N_2665,N_2904);
or UO_222 (O_222,N_2376,N_2075);
nand UO_223 (O_223,N_2233,N_2945);
nor UO_224 (O_224,N_2117,N_2514);
nand UO_225 (O_225,N_2301,N_2246);
nand UO_226 (O_226,N_2824,N_2731);
xor UO_227 (O_227,N_2206,N_2709);
nand UO_228 (O_228,N_2705,N_2671);
nand UO_229 (O_229,N_2262,N_2946);
nor UO_230 (O_230,N_2816,N_2426);
or UO_231 (O_231,N_2293,N_2850);
or UO_232 (O_232,N_2606,N_2844);
nand UO_233 (O_233,N_2670,N_2585);
xnor UO_234 (O_234,N_2960,N_2966);
xnor UO_235 (O_235,N_2085,N_2933);
xnor UO_236 (O_236,N_2786,N_2841);
xor UO_237 (O_237,N_2589,N_2525);
or UO_238 (O_238,N_2094,N_2304);
xor UO_239 (O_239,N_2296,N_2582);
xor UO_240 (O_240,N_2383,N_2648);
nand UO_241 (O_241,N_2538,N_2569);
nor UO_242 (O_242,N_2095,N_2835);
or UO_243 (O_243,N_2799,N_2027);
xnor UO_244 (O_244,N_2742,N_2623);
and UO_245 (O_245,N_2406,N_2288);
and UO_246 (O_246,N_2903,N_2234);
nand UO_247 (O_247,N_2036,N_2833);
or UO_248 (O_248,N_2500,N_2000);
or UO_249 (O_249,N_2043,N_2303);
nand UO_250 (O_250,N_2274,N_2450);
and UO_251 (O_251,N_2972,N_2380);
xnor UO_252 (O_252,N_2683,N_2156);
or UO_253 (O_253,N_2238,N_2169);
nand UO_254 (O_254,N_2263,N_2888);
and UO_255 (O_255,N_2333,N_2182);
nand UO_256 (O_256,N_2996,N_2074);
or UO_257 (O_257,N_2545,N_2053);
and UO_258 (O_258,N_2917,N_2490);
or UO_259 (O_259,N_2889,N_2849);
nand UO_260 (O_260,N_2330,N_2286);
xnor UO_261 (O_261,N_2446,N_2405);
or UO_262 (O_262,N_2943,N_2692);
xnor UO_263 (O_263,N_2550,N_2410);
nor UO_264 (O_264,N_2281,N_2776);
nor UO_265 (O_265,N_2349,N_2523);
xnor UO_266 (O_266,N_2652,N_2113);
xnor UO_267 (O_267,N_2392,N_2009);
and UO_268 (O_268,N_2687,N_2455);
xnor UO_269 (O_269,N_2231,N_2867);
nor UO_270 (O_270,N_2258,N_2827);
xnor UO_271 (O_271,N_2515,N_2054);
nand UO_272 (O_272,N_2669,N_2756);
or UO_273 (O_273,N_2193,N_2567);
and UO_274 (O_274,N_2147,N_2216);
xnor UO_275 (O_275,N_2183,N_2218);
nand UO_276 (O_276,N_2468,N_2337);
nand UO_277 (O_277,N_2991,N_2804);
and UO_278 (O_278,N_2620,N_2195);
nor UO_279 (O_279,N_2289,N_2030);
or UO_280 (O_280,N_2761,N_2927);
xor UO_281 (O_281,N_2934,N_2306);
nand UO_282 (O_282,N_2499,N_2419);
nor UO_283 (O_283,N_2261,N_2540);
nand UO_284 (O_284,N_2815,N_2519);
xor UO_285 (O_285,N_2158,N_2689);
xor UO_286 (O_286,N_2101,N_2472);
nor UO_287 (O_287,N_2820,N_2382);
nor UO_288 (O_288,N_2390,N_2014);
xnor UO_289 (O_289,N_2005,N_2726);
nor UO_290 (O_290,N_2388,N_2016);
xnor UO_291 (O_291,N_2878,N_2896);
and UO_292 (O_292,N_2916,N_2164);
nand UO_293 (O_293,N_2084,N_2482);
nand UO_294 (O_294,N_2707,N_2324);
xor UO_295 (O_295,N_2372,N_2798);
or UO_296 (O_296,N_2089,N_2953);
xnor UO_297 (O_297,N_2481,N_2682);
xnor UO_298 (O_298,N_2473,N_2730);
xor UO_299 (O_299,N_2479,N_2529);
or UO_300 (O_300,N_2963,N_2872);
nand UO_301 (O_301,N_2964,N_2805);
nor UO_302 (O_302,N_2839,N_2360);
and UO_303 (O_303,N_2906,N_2772);
nor UO_304 (O_304,N_2881,N_2653);
xor UO_305 (O_305,N_2684,N_2154);
nor UO_306 (O_306,N_2048,N_2612);
nor UO_307 (O_307,N_2224,N_2416);
or UO_308 (O_308,N_2020,N_2361);
and UO_309 (O_309,N_2808,N_2171);
nor UO_310 (O_310,N_2433,N_2222);
and UO_311 (O_311,N_2032,N_2597);
and UO_312 (O_312,N_2362,N_2018);
nor UO_313 (O_313,N_2639,N_2435);
xnor UO_314 (O_314,N_2347,N_2111);
xor UO_315 (O_315,N_2728,N_2423);
nand UO_316 (O_316,N_2704,N_2502);
nand UO_317 (O_317,N_2374,N_2029);
and UO_318 (O_318,N_2061,N_2625);
or UO_319 (O_319,N_2308,N_2819);
nand UO_320 (O_320,N_2936,N_2132);
nand UO_321 (O_321,N_2630,N_2136);
nor UO_322 (O_322,N_2425,N_2659);
xor UO_323 (O_323,N_2494,N_2350);
and UO_324 (O_324,N_2862,N_2369);
or UO_325 (O_325,N_2914,N_2408);
and UO_326 (O_326,N_2548,N_2429);
and UO_327 (O_327,N_2534,N_2176);
nand UO_328 (O_328,N_2506,N_2357);
xor UO_329 (O_329,N_2950,N_2722);
xor UO_330 (O_330,N_2641,N_2159);
or UO_331 (O_331,N_2397,N_2068);
xor UO_332 (O_332,N_2483,N_2187);
xnor UO_333 (O_333,N_2174,N_2982);
xor UO_334 (O_334,N_2909,N_2457);
and UO_335 (O_335,N_2385,N_2056);
nand UO_336 (O_336,N_2618,N_2926);
or UO_337 (O_337,N_2624,N_2894);
or UO_338 (O_338,N_2504,N_2720);
and UO_339 (O_339,N_2860,N_2517);
or UO_340 (O_340,N_2590,N_2389);
xor UO_341 (O_341,N_2082,N_2321);
and UO_342 (O_342,N_2521,N_2773);
or UO_343 (O_343,N_2701,N_2635);
nand UO_344 (O_344,N_2781,N_2034);
nor UO_345 (O_345,N_2755,N_2575);
nor UO_346 (O_346,N_2535,N_2543);
xor UO_347 (O_347,N_2363,N_2759);
nor UO_348 (O_348,N_2656,N_2790);
nand UO_349 (O_349,N_2417,N_2600);
nand UO_350 (O_350,N_2280,N_2777);
xor UO_351 (O_351,N_2676,N_2724);
nor UO_352 (O_352,N_2256,N_2434);
nor UO_353 (O_353,N_2052,N_2355);
xor UO_354 (O_354,N_2970,N_2821);
xor UO_355 (O_355,N_2734,N_2114);
nor UO_356 (O_356,N_2719,N_2727);
or UO_357 (O_357,N_2613,N_2686);
or UO_358 (O_358,N_2153,N_2845);
or UO_359 (O_359,N_2997,N_2452);
and UO_360 (O_360,N_2214,N_2087);
nor UO_361 (O_361,N_2563,N_2010);
nor UO_362 (O_362,N_2404,N_2470);
or UO_363 (O_363,N_2194,N_2110);
and UO_364 (O_364,N_2885,N_2400);
nand UO_365 (O_365,N_2721,N_2918);
nand UO_366 (O_366,N_2366,N_2462);
and UO_367 (O_367,N_2414,N_2875);
nand UO_368 (O_368,N_2239,N_2167);
or UO_369 (O_369,N_2127,N_2868);
nand UO_370 (O_370,N_2086,N_2980);
nor UO_371 (O_371,N_2033,N_2830);
and UO_372 (O_372,N_2584,N_2104);
nor UO_373 (O_373,N_2847,N_2923);
nand UO_374 (O_374,N_2718,N_2703);
nor UO_375 (O_375,N_2711,N_2939);
and UO_376 (O_376,N_2358,N_2375);
and UO_377 (O_377,N_2024,N_2486);
nand UO_378 (O_378,N_2449,N_2806);
and UO_379 (O_379,N_2741,N_2307);
and UO_380 (O_380,N_2044,N_2886);
nand UO_381 (O_381,N_2475,N_2583);
and UO_382 (O_382,N_2882,N_2901);
xor UO_383 (O_383,N_2346,N_2969);
and UO_384 (O_384,N_2413,N_2252);
or UO_385 (O_385,N_2364,N_2995);
or UO_386 (O_386,N_2073,N_2902);
and UO_387 (O_387,N_2539,N_2998);
xnor UO_388 (O_388,N_2217,N_2083);
xnor UO_389 (O_389,N_2602,N_2919);
or UO_390 (O_390,N_2001,N_2737);
or UO_391 (O_391,N_2572,N_2088);
xnor UO_392 (O_392,N_2232,N_2957);
xnor UO_393 (O_393,N_2527,N_2752);
nor UO_394 (O_394,N_2831,N_2144);
nand UO_395 (O_395,N_2924,N_2513);
nand UO_396 (O_396,N_2767,N_2260);
or UO_397 (O_397,N_2764,N_2605);
xor UO_398 (O_398,N_2295,N_2339);
nor UO_399 (O_399,N_2477,N_2990);
or UO_400 (O_400,N_2628,N_2636);
xnor UO_401 (O_401,N_2851,N_2698);
and UO_402 (O_402,N_2699,N_2526);
nor UO_403 (O_403,N_2311,N_2573);
xnor UO_404 (O_404,N_2931,N_2496);
or UO_405 (O_405,N_2447,N_2151);
or UO_406 (O_406,N_2913,N_2242);
xor UO_407 (O_407,N_2279,N_2858);
nand UO_408 (O_408,N_2803,N_2063);
xor UO_409 (O_409,N_2331,N_2622);
and UO_410 (O_410,N_2422,N_2327);
nand UO_411 (O_411,N_2278,N_2211);
xnor UO_412 (O_412,N_2782,N_2562);
xor UO_413 (O_413,N_2658,N_2674);
nand UO_414 (O_414,N_2697,N_2081);
or UO_415 (O_415,N_2498,N_2019);
and UO_416 (O_416,N_2654,N_2595);
nand UO_417 (O_417,N_2255,N_2510);
xor UO_418 (O_418,N_2055,N_2025);
or UO_419 (O_419,N_2396,N_2661);
nand UO_420 (O_420,N_2938,N_2873);
xnor UO_421 (O_421,N_2631,N_2066);
and UO_422 (O_422,N_2743,N_2038);
xor UO_423 (O_423,N_2891,N_2213);
and UO_424 (O_424,N_2247,N_2530);
nand UO_425 (O_425,N_2949,N_2059);
or UO_426 (O_426,N_2884,N_2928);
xor UO_427 (O_427,N_2257,N_2570);
xor UO_428 (O_428,N_2579,N_2508);
nand UO_429 (O_429,N_2122,N_2265);
and UO_430 (O_430,N_2443,N_2812);
or UO_431 (O_431,N_2067,N_2753);
xor UO_432 (O_432,N_2893,N_2551);
and UO_433 (O_433,N_2196,N_2138);
or UO_434 (O_434,N_2596,N_2190);
nor UO_435 (O_435,N_2495,N_2822);
or UO_436 (O_436,N_2091,N_2533);
or UO_437 (O_437,N_2644,N_2463);
xnor UO_438 (O_438,N_2106,N_2219);
or UO_439 (O_439,N_2420,N_2975);
nand UO_440 (O_440,N_2250,N_2634);
or UO_441 (O_441,N_2626,N_2398);
nor UO_442 (O_442,N_2045,N_2409);
and UO_443 (O_443,N_2150,N_2179);
xnor UO_444 (O_444,N_2935,N_2177);
nor UO_445 (O_445,N_2042,N_2049);
nor UO_446 (O_446,N_2135,N_2373);
nor UO_447 (O_447,N_2932,N_2954);
nand UO_448 (O_448,N_2556,N_2354);
nand UO_449 (O_449,N_2984,N_2487);
nor UO_450 (O_450,N_2090,N_2381);
and UO_451 (O_451,N_2633,N_2387);
nor UO_452 (O_452,N_2842,N_2093);
nor UO_453 (O_453,N_2103,N_2507);
or UO_454 (O_454,N_2929,N_2284);
xor UO_455 (O_455,N_2163,N_2922);
xnor UO_456 (O_456,N_2161,N_2611);
and UO_457 (O_457,N_2118,N_2461);
and UO_458 (O_458,N_2172,N_2651);
nand UO_459 (O_459,N_2621,N_2619);
and UO_460 (O_460,N_2829,N_2897);
nand UO_461 (O_461,N_2852,N_2642);
and UO_462 (O_462,N_2588,N_2072);
nor UO_463 (O_463,N_2012,N_2561);
nor UO_464 (O_464,N_2859,N_2200);
xor UO_465 (O_465,N_2488,N_2356);
nor UO_466 (O_466,N_2121,N_2119);
nor UO_467 (O_467,N_2800,N_2070);
or UO_468 (O_468,N_2015,N_2098);
and UO_469 (O_469,N_2542,N_2832);
xnor UO_470 (O_470,N_2979,N_2305);
or UO_471 (O_471,N_2391,N_2925);
nor UO_472 (O_472,N_2476,N_2329);
and UO_473 (O_473,N_2696,N_2204);
nor UO_474 (O_474,N_2973,N_2754);
nand UO_475 (O_475,N_2282,N_2141);
nor UO_476 (O_476,N_2145,N_2427);
nor UO_477 (O_477,N_2577,N_2668);
nor UO_478 (O_478,N_2022,N_2317);
or UO_479 (O_479,N_2865,N_2520);
nand UO_480 (O_480,N_2558,N_2013);
xnor UO_481 (O_481,N_2060,N_2541);
and UO_482 (O_482,N_2459,N_2650);
nand UO_483 (O_483,N_2322,N_2757);
nor UO_484 (O_484,N_2454,N_2137);
nand UO_485 (O_485,N_2235,N_2184);
nand UO_486 (O_486,N_2230,N_2291);
or UO_487 (O_487,N_2944,N_2989);
or UO_488 (O_488,N_2140,N_2130);
nor UO_489 (O_489,N_2270,N_2810);
nand UO_490 (O_490,N_2146,N_2428);
nor UO_491 (O_491,N_2273,N_2657);
nor UO_492 (O_492,N_2834,N_2407);
nand UO_493 (O_493,N_2736,N_2191);
nor UO_494 (O_494,N_2876,N_2983);
and UO_495 (O_495,N_2912,N_2793);
nand UO_496 (O_496,N_2359,N_2062);
nor UO_497 (O_497,N_2715,N_2028);
and UO_498 (O_498,N_2309,N_2861);
xnor UO_499 (O_499,N_2733,N_2871);
endmodule