module basic_750_5000_1000_2_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2503,N_2505,N_2506,N_2507,N_2509,N_2510,N_2512,N_2513,N_2514,N_2515,N_2516,N_2518,N_2519,N_2520,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2529,N_2530,N_2531,N_2533,N_2534,N_2535,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2545,N_2546,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2555,N_2556,N_2557,N_2559,N_2560,N_2561,N_2563,N_2564,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2578,N_2579,N_2580,N_2582,N_2583,N_2584,N_2587,N_2589,N_2592,N_2593,N_2595,N_2596,N_2598,N_2599,N_2600,N_2601,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2616,N_2617,N_2618,N_2619,N_2621,N_2622,N_2623,N_2625,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2644,N_2645,N_2646,N_2647,N_2648,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2659,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2668,N_2669,N_2670,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2681,N_2682,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2692,N_2693,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2705,N_2706,N_2707,N_2708,N_2709,N_2711,N_2712,N_2713,N_2714,N_2716,N_2717,N_2718,N_2720,N_2721,N_2722,N_2724,N_2725,N_2726,N_2727,N_2730,N_2731,N_2732,N_2733,N_2734,N_2736,N_2737,N_2738,N_2739,N_2740,N_2742,N_2743,N_2744,N_2746,N_2747,N_2748,N_2750,N_2752,N_2753,N_2754,N_2756,N_2757,N_2758,N_2759,N_2760,N_2762,N_2763,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2775,N_2776,N_2777,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2813,N_2814,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2824,N_2826,N_2828,N_2829,N_2830,N_2831,N_2832,N_2834,N_2835,N_2836,N_2838,N_2839,N_2840,N_2845,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2854,N_2855,N_2857,N_2858,N_2859,N_2860,N_2863,N_2864,N_2865,N_2867,N_2869,N_2870,N_2871,N_2872,N_2874,N_2875,N_2876,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2885,N_2886,N_2887,N_2888,N_2889,N_2891,N_2893,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2913,N_2914,N_2915,N_2916,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2941,N_2942,N_2945,N_2947,N_2948,N_2949,N_2950,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2962,N_2963,N_2964,N_2965,N_2966,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2979,N_2980,N_2981,N_2982,N_2985,N_2986,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3027,N_3029,N_3030,N_3032,N_3033,N_3034,N_3036,N_3037,N_3039,N_3041,N_3042,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3060,N_3061,N_3062,N_3063,N_3065,N_3066,N_3068,N_3069,N_3070,N_3071,N_3072,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3124,N_3128,N_3129,N_3131,N_3132,N_3135,N_3136,N_3137,N_3138,N_3139,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3151,N_3153,N_3154,N_3156,N_3157,N_3158,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3208,N_3209,N_3211,N_3212,N_3213,N_3214,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3247,N_3248,N_3250,N_3251,N_3252,N_3253,N_3255,N_3256,N_3257,N_3258,N_3260,N_3261,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3273,N_3274,N_3276,N_3277,N_3278,N_3280,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3338,N_3340,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3354,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3395,N_3396,N_3397,N_3398,N_3399,N_3401,N_3402,N_3403,N_3405,N_3406,N_3408,N_3409,N_3411,N_3413,N_3414,N_3415,N_3416,N_3417,N_3419,N_3420,N_3421,N_3423,N_3424,N_3425,N_3426,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3435,N_3436,N_3437,N_3439,N_3440,N_3441,N_3442,N_3443,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3463,N_3464,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3479,N_3480,N_3482,N_3483,N_3484,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3496,N_3498,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3523,N_3524,N_3525,N_3526,N_3528,N_3529,N_3530,N_3531,N_3532,N_3534,N_3535,N_3537,N_3538,N_3539,N_3540,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3559,N_3561,N_3563,N_3564,N_3565,N_3568,N_3569,N_3571,N_3573,N_3574,N_3575,N_3577,N_3578,N_3579,N_3580,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3589,N_3590,N_3591,N_3592,N_3593,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3609,N_3610,N_3611,N_3613,N_3614,N_3616,N_3618,N_3619,N_3620,N_3621,N_3622,N_3624,N_3625,N_3626,N_3628,N_3629,N_3630,N_3632,N_3634,N_3635,N_3638,N_3639,N_3641,N_3642,N_3643,N_3644,N_3645,N_3647,N_3648,N_3649,N_3650,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3661,N_3662,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3680,N_3681,N_3683,N_3684,N_3685,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3695,N_3696,N_3697,N_3698,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3728,N_3729,N_3731,N_3732,N_3734,N_3735,N_3736,N_3737,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3768,N_3769,N_3770,N_3772,N_3773,N_3774,N_3775,N_3776,N_3778,N_3780,N_3781,N_3783,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3814,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3834,N_3836,N_3837,N_3838,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3851,N_3852,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3862,N_3865,N_3866,N_3867,N_3868,N_3869,N_3872,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3903,N_3904,N_3906,N_3907,N_3908,N_3909,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3918,N_3920,N_3921,N_3923,N_3924,N_3928,N_3930,N_3932,N_3934,N_3936,N_3937,N_3938,N_3939,N_3941,N_3943,N_3944,N_3945,N_3946,N_3947,N_3949,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3967,N_3968,N_3969,N_3970,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3986,N_3987,N_3989,N_3990,N_3992,N_3993,N_3994,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4005,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4015,N_4016,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4025,N_4028,N_4029,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4039,N_4040,N_4042,N_4044,N_4045,N_4046,N_4047,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4057,N_4058,N_4059,N_4061,N_4062,N_4065,N_4066,N_4068,N_4069,N_4070,N_4071,N_4072,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4083,N_4084,N_4085,N_4087,N_4088,N_4089,N_4090,N_4091,N_4093,N_4094,N_4095,N_4096,N_4097,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4109,N_4110,N_4111,N_4113,N_4115,N_4117,N_4118,N_4119,N_4120,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4131,N_4132,N_4133,N_4136,N_4137,N_4138,N_4139,N_4140,N_4142,N_4143,N_4144,N_4145,N_4147,N_4148,N_4150,N_4151,N_4152,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4161,N_4162,N_4163,N_4164,N_4166,N_4167,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4194,N_4197,N_4198,N_4200,N_4201,N_4203,N_4204,N_4205,N_4206,N_4207,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4225,N_4226,N_4227,N_4229,N_4230,N_4231,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4240,N_4241,N_4242,N_4243,N_4245,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4263,N_4264,N_4267,N_4268,N_4269,N_4270,N_4274,N_4275,N_4276,N_4277,N_4279,N_4280,N_4281,N_4283,N_4284,N_4285,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4295,N_4298,N_4299,N_4302,N_4303,N_4304,N_4307,N_4308,N_4310,N_4311,N_4312,N_4313,N_4314,N_4316,N_4317,N_4318,N_4319,N_4320,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4332,N_4333,N_4334,N_4335,N_4336,N_4338,N_4340,N_4341,N_4342,N_4345,N_4346,N_4348,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4370,N_4371,N_4372,N_4373,N_4377,N_4378,N_4379,N_4380,N_4381,N_4383,N_4385,N_4386,N_4388,N_4389,N_4390,N_4391,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4402,N_4404,N_4405,N_4406,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4478,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4505,N_4506,N_4507,N_4508,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4517,N_4518,N_4519,N_4522,N_4523,N_4524,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4541,N_4542,N_4543,N_4545,N_4546,N_4548,N_4550,N_4551,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4614,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4634,N_4635,N_4636,N_4639,N_4640,N_4641,N_4642,N_4644,N_4646,N_4647,N_4649,N_4650,N_4651,N_4652,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4675,N_4677,N_4678,N_4679,N_4680,N_4684,N_4686,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4695,N_4696,N_4697,N_4698,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4739,N_4740,N_4745,N_4747,N_4749,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4762,N_4766,N_4767,N_4768,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4786,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4808,N_4809,N_4811,N_4812,N_4813,N_4814,N_4815,N_4818,N_4819,N_4820,N_4821,N_4822,N_4824,N_4825,N_4826,N_4827,N_4828,N_4832,N_4833,N_4834,N_4835,N_4836,N_4840,N_4841,N_4842,N_4845,N_4847,N_4848,N_4849,N_4851,N_4852,N_4853,N_4854,N_4855,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4870,N_4871,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4884,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4899,N_4900,N_4901,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4917,N_4919,N_4921,N_4922,N_4923,N_4924,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4937,N_4938,N_4939,N_4942,N_4943,N_4944,N_4945,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4979,N_4983,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4998,N_4999;
nand U0 (N_0,In_250,In_649);
nor U1 (N_1,In_681,In_563);
nand U2 (N_2,In_59,In_748);
nand U3 (N_3,In_429,In_679);
nor U4 (N_4,In_643,In_50);
nor U5 (N_5,In_283,In_249);
and U6 (N_6,In_530,In_339);
nand U7 (N_7,In_452,In_722);
nor U8 (N_8,In_96,In_98);
xnor U9 (N_9,In_324,In_585);
nand U10 (N_10,In_160,In_354);
nand U11 (N_11,In_86,In_221);
and U12 (N_12,In_64,In_177);
and U13 (N_13,In_277,In_32);
nor U14 (N_14,In_149,In_708);
nor U15 (N_15,In_77,In_731);
or U16 (N_16,In_484,In_472);
xnor U17 (N_17,In_22,In_12);
or U18 (N_18,In_686,In_516);
nor U19 (N_19,In_533,In_45);
xor U20 (N_20,In_402,In_519);
or U21 (N_21,In_747,In_348);
nand U22 (N_22,In_364,In_636);
or U23 (N_23,In_743,In_670);
nor U24 (N_24,In_235,In_280);
and U25 (N_25,In_721,In_38);
and U26 (N_26,In_40,In_596);
and U27 (N_27,In_198,In_203);
nand U28 (N_28,In_180,In_661);
xnor U29 (N_29,In_410,In_209);
nand U30 (N_30,In_674,In_434);
and U31 (N_31,In_702,In_78);
or U32 (N_32,In_729,In_610);
or U33 (N_33,In_181,In_246);
and U34 (N_34,In_468,In_659);
xor U35 (N_35,In_311,In_33);
nor U36 (N_36,In_145,In_122);
xnor U37 (N_37,In_44,In_407);
nand U38 (N_38,In_243,In_475);
nand U39 (N_39,In_505,In_453);
nand U40 (N_40,In_346,In_626);
xor U41 (N_41,In_361,In_606);
nand U42 (N_42,In_598,In_321);
nand U43 (N_43,In_683,In_213);
xnor U44 (N_44,In_25,In_546);
xor U45 (N_45,In_138,In_171);
xnor U46 (N_46,In_706,In_673);
and U47 (N_47,In_230,In_603);
nor U48 (N_48,In_545,In_318);
and U49 (N_49,In_539,In_624);
nor U50 (N_50,In_133,In_582);
nand U51 (N_51,In_46,In_501);
and U52 (N_52,In_100,In_615);
nand U53 (N_53,In_455,In_314);
nand U54 (N_54,In_34,In_581);
nand U55 (N_55,In_335,In_61);
xnor U56 (N_56,In_552,In_657);
or U57 (N_57,In_337,In_68);
xor U58 (N_58,In_294,In_675);
or U59 (N_59,In_279,In_597);
xnor U60 (N_60,In_144,In_668);
or U61 (N_61,In_471,In_24);
nand U62 (N_62,In_518,In_489);
or U63 (N_63,In_586,In_602);
and U64 (N_64,In_51,In_423);
and U65 (N_65,In_616,In_166);
nand U66 (N_66,In_744,In_469);
or U67 (N_67,In_334,In_634);
xor U68 (N_68,In_111,In_730);
and U69 (N_69,In_89,In_413);
nor U70 (N_70,In_608,In_349);
and U71 (N_71,In_91,In_291);
or U72 (N_72,In_698,In_225);
xor U73 (N_73,In_232,In_80);
nand U74 (N_74,In_266,In_384);
nand U75 (N_75,In_537,In_151);
and U76 (N_76,In_503,In_693);
and U77 (N_77,In_49,In_633);
nor U78 (N_78,In_264,In_58);
nand U79 (N_79,In_67,In_543);
xnor U80 (N_80,In_477,In_255);
nand U81 (N_81,In_415,In_742);
nor U82 (N_82,In_15,In_688);
xnor U83 (N_83,In_142,In_482);
and U84 (N_84,In_82,In_214);
nand U85 (N_85,In_701,In_116);
nand U86 (N_86,In_196,In_385);
and U87 (N_87,In_726,In_92);
nor U88 (N_88,In_493,In_135);
xnor U89 (N_89,In_589,In_382);
xnor U90 (N_90,In_548,In_593);
or U91 (N_91,In_449,In_247);
nor U92 (N_92,In_445,In_363);
xnor U93 (N_93,In_320,In_682);
and U94 (N_94,In_3,In_262);
xnor U95 (N_95,In_558,In_669);
xnor U96 (N_96,In_459,In_28);
xnor U97 (N_97,In_454,In_511);
and U98 (N_98,In_513,In_226);
xnor U99 (N_99,In_672,In_336);
xnor U100 (N_100,In_719,In_35);
xor U101 (N_101,In_442,In_430);
and U102 (N_102,In_26,In_724);
and U103 (N_103,In_458,In_6);
or U104 (N_104,In_551,In_689);
nor U105 (N_105,In_605,In_451);
xnor U106 (N_106,In_141,In_562);
nand U107 (N_107,In_467,In_717);
nor U108 (N_108,In_161,In_23);
and U109 (N_109,In_660,In_486);
and U110 (N_110,In_319,In_491);
or U111 (N_111,In_43,In_400);
xor U112 (N_112,In_515,In_658);
xnor U113 (N_113,In_268,In_441);
xnor U114 (N_114,In_139,In_535);
nand U115 (N_115,In_715,In_611);
nand U116 (N_116,In_465,In_179);
or U117 (N_117,In_323,In_749);
nor U118 (N_118,In_432,In_295);
xnor U119 (N_119,In_200,In_736);
nor U120 (N_120,In_549,In_547);
or U121 (N_121,In_147,In_114);
and U122 (N_122,In_222,In_576);
or U123 (N_123,In_521,In_629);
and U124 (N_124,In_732,In_508);
nand U125 (N_125,In_165,In_63);
or U126 (N_126,In_307,In_368);
and U127 (N_127,In_630,In_322);
nand U128 (N_128,In_375,In_527);
nand U129 (N_129,In_446,In_102);
and U130 (N_130,In_480,In_297);
or U131 (N_131,In_374,In_263);
xor U132 (N_132,In_261,In_298);
nand U133 (N_133,In_716,In_478);
or U134 (N_134,In_189,In_350);
xnor U135 (N_135,In_639,In_456);
or U136 (N_136,In_276,In_65);
nand U137 (N_137,In_14,In_542);
or U138 (N_138,In_627,In_176);
and U139 (N_139,In_56,In_424);
xor U140 (N_140,In_403,In_207);
xor U141 (N_141,In_245,In_281);
nor U142 (N_142,In_740,In_461);
and U143 (N_143,In_571,In_391);
or U144 (N_144,In_621,In_671);
xnor U145 (N_145,In_257,In_388);
or U146 (N_146,In_488,In_162);
nand U147 (N_147,In_330,In_574);
nor U148 (N_148,In_405,In_306);
or U149 (N_149,In_328,In_310);
or U150 (N_150,In_417,In_378);
or U151 (N_151,In_308,In_696);
and U152 (N_152,In_316,In_664);
or U153 (N_153,In_199,In_218);
xor U154 (N_154,In_395,In_398);
and U155 (N_155,In_228,In_396);
or U156 (N_156,In_631,In_329);
xnor U157 (N_157,In_191,In_399);
nor U158 (N_158,In_258,In_437);
nor U159 (N_159,In_460,In_473);
nor U160 (N_160,In_103,In_483);
nor U161 (N_161,In_514,In_8);
nor U162 (N_162,In_19,In_20);
nand U163 (N_163,In_57,In_691);
or U164 (N_164,In_565,In_344);
or U165 (N_165,In_738,In_409);
nand U166 (N_166,In_231,In_99);
and U167 (N_167,In_520,In_587);
nor U168 (N_168,In_408,In_739);
nand U169 (N_169,In_112,In_617);
and U170 (N_170,In_566,In_287);
nor U171 (N_171,In_13,In_416);
or U172 (N_172,In_41,In_108);
and U173 (N_173,In_684,In_609);
nand U174 (N_174,In_87,In_700);
nand U175 (N_175,In_187,In_599);
xnor U176 (N_176,In_544,In_590);
and U177 (N_177,In_367,In_340);
nand U178 (N_178,In_619,In_169);
nor U179 (N_179,In_663,In_522);
and U180 (N_180,In_278,In_97);
or U181 (N_181,In_685,In_284);
xnor U182 (N_182,In_433,In_564);
and U183 (N_183,In_677,In_241);
xnor U184 (N_184,In_79,In_105);
nand U185 (N_185,In_302,In_130);
and U186 (N_186,In_267,In_140);
and U187 (N_187,In_389,In_195);
xor U188 (N_188,In_123,In_369);
nor U189 (N_189,In_632,In_440);
xnor U190 (N_190,In_260,In_353);
nand U191 (N_191,In_327,In_252);
and U192 (N_192,In_583,In_131);
and U193 (N_193,In_652,In_259);
nand U194 (N_194,In_366,In_418);
or U195 (N_195,In_604,In_338);
and U196 (N_196,In_536,In_746);
or U197 (N_197,In_269,In_342);
or U198 (N_198,In_466,In_600);
and U199 (N_199,In_81,In_175);
and U200 (N_200,In_153,In_271);
or U201 (N_201,In_110,In_325);
or U202 (N_202,In_370,In_601);
or U203 (N_203,In_372,In_224);
and U204 (N_204,In_2,In_220);
nand U205 (N_205,In_376,In_579);
or U206 (N_206,In_301,In_642);
nand U207 (N_207,In_83,In_412);
nand U208 (N_208,In_72,In_404);
nor U209 (N_209,In_431,In_55);
and U210 (N_210,In_186,In_251);
nor U211 (N_211,In_435,In_554);
nor U212 (N_212,In_5,In_705);
xor U213 (N_213,In_494,In_359);
nand U214 (N_214,In_623,In_448);
or U215 (N_215,In_377,In_242);
nand U216 (N_216,In_90,In_383);
nor U217 (N_217,In_580,In_578);
nor U218 (N_218,In_290,In_293);
and U219 (N_219,In_463,In_299);
or U220 (N_220,In_572,In_436);
and U221 (N_221,In_524,In_9);
xor U222 (N_222,In_690,In_421);
nor U223 (N_223,In_365,In_113);
and U224 (N_224,In_733,In_227);
nor U225 (N_225,In_504,In_355);
nand U226 (N_226,In_206,In_317);
or U227 (N_227,In_561,In_714);
and U228 (N_228,In_728,In_397);
nand U229 (N_229,In_592,In_347);
or U230 (N_230,In_18,In_699);
or U231 (N_231,In_735,In_39);
nand U232 (N_232,In_119,In_305);
xnor U233 (N_233,In_115,In_644);
or U234 (N_234,In_233,In_725);
nor U235 (N_235,In_124,In_737);
nand U236 (N_236,In_69,In_635);
xor U237 (N_237,In_553,In_595);
and U238 (N_238,In_183,In_204);
nor U239 (N_239,In_95,In_170);
nand U240 (N_240,In_93,In_156);
nand U241 (N_241,In_439,In_387);
and U242 (N_242,In_358,In_4);
and U243 (N_243,In_628,In_155);
and U244 (N_244,In_202,In_695);
nor U245 (N_245,In_31,In_568);
nor U246 (N_246,In_326,In_485);
nor U247 (N_247,In_680,In_531);
xor U248 (N_248,In_289,In_625);
nor U249 (N_249,In_237,In_622);
and U250 (N_250,In_136,In_534);
or U251 (N_251,In_205,In_29);
or U252 (N_252,In_117,In_517);
nand U253 (N_253,In_379,In_178);
nand U254 (N_254,In_154,In_502);
xnor U255 (N_255,In_345,In_666);
nor U256 (N_256,In_723,In_727);
or U257 (N_257,In_0,In_219);
nor U258 (N_258,In_148,In_647);
nand U259 (N_259,In_497,In_125);
nand U260 (N_260,In_60,In_47);
xnor U261 (N_261,In_272,In_185);
xor U262 (N_262,In_357,In_17);
and U263 (N_263,In_425,In_498);
nor U264 (N_264,In_406,In_7);
or U265 (N_265,In_174,In_66);
nor U266 (N_266,In_697,In_720);
nand U267 (N_267,In_238,In_16);
and U268 (N_268,In_381,In_270);
or U269 (N_269,In_236,In_392);
or U270 (N_270,In_573,In_30);
or U271 (N_271,In_464,In_168);
nor U272 (N_272,In_193,In_152);
xor U273 (N_273,In_470,In_481);
and U274 (N_274,In_710,In_303);
nand U275 (N_275,In_490,In_665);
or U276 (N_276,In_27,In_532);
nand U277 (N_277,In_704,In_687);
nand U278 (N_278,In_127,In_134);
nor U279 (N_279,In_76,In_10);
or U280 (N_280,In_640,In_215);
or U281 (N_281,In_645,In_496);
and U282 (N_282,In_394,In_248);
nor U283 (N_283,In_707,In_618);
nand U284 (N_284,In_343,In_438);
or U285 (N_285,In_75,In_285);
nor U286 (N_286,In_555,In_653);
and U287 (N_287,In_510,In_159);
nand U288 (N_288,In_507,In_157);
xor U289 (N_289,In_300,In_709);
nand U290 (N_290,In_201,In_254);
xnor U291 (N_291,In_584,In_120);
nand U292 (N_292,In_309,In_210);
xor U293 (N_293,In_462,In_256);
or U294 (N_294,In_362,In_208);
nor U295 (N_295,In_393,In_651);
and U296 (N_296,In_286,In_655);
nor U297 (N_297,In_85,In_73);
and U298 (N_298,In_426,In_620);
and U299 (N_299,In_487,In_70);
nor U300 (N_300,In_692,In_234);
nor U301 (N_301,In_331,In_275);
or U302 (N_302,In_229,In_648);
and U303 (N_303,In_182,In_457);
and U304 (N_304,In_380,In_495);
nand U305 (N_305,In_559,In_313);
or U306 (N_306,In_273,In_474);
or U307 (N_307,In_713,In_101);
xnor U308 (N_308,In_121,In_21);
xor U309 (N_309,In_447,In_575);
and U310 (N_310,In_567,In_570);
or U311 (N_311,In_741,In_332);
nand U312 (N_312,In_500,In_656);
nand U313 (N_313,In_499,In_126);
xnor U314 (N_314,In_54,In_37);
xor U315 (N_315,In_253,In_74);
xnor U316 (N_316,In_167,In_163);
or U317 (N_317,In_509,In_386);
and U318 (N_318,In_239,In_712);
xnor U319 (N_319,In_591,In_107);
and U320 (N_320,In_282,In_212);
and U321 (N_321,In_312,In_641);
xor U322 (N_322,In_476,In_612);
xnor U323 (N_323,In_146,In_443);
xnor U324 (N_324,In_694,In_42);
or U325 (N_325,In_654,In_390);
nor U326 (N_326,In_373,In_192);
nand U327 (N_327,In_676,In_703);
or U328 (N_328,In_211,In_428);
nand U329 (N_329,In_52,In_745);
xor U330 (N_330,In_184,In_734);
or U331 (N_331,In_718,In_678);
xnor U332 (N_332,In_506,In_128);
or U333 (N_333,In_352,In_173);
or U334 (N_334,In_371,In_197);
or U335 (N_335,In_104,In_129);
xnor U336 (N_336,In_288,In_164);
xnor U337 (N_337,In_109,In_444);
nand U338 (N_338,In_240,In_557);
nor U339 (N_339,In_646,In_190);
nand U340 (N_340,In_84,In_143);
or U341 (N_341,In_150,In_172);
nor U342 (N_342,In_296,In_223);
or U343 (N_343,In_62,In_333);
nor U344 (N_344,In_427,In_132);
xor U345 (N_345,In_422,In_550);
or U346 (N_346,In_53,In_137);
or U347 (N_347,In_613,In_217);
nand U348 (N_348,In_304,In_492);
or U349 (N_349,In_401,In_526);
xnor U350 (N_350,In_411,In_414);
and U351 (N_351,In_711,In_538);
xnor U352 (N_352,In_351,In_594);
or U353 (N_353,In_419,In_560);
xor U354 (N_354,In_529,In_274);
or U355 (N_355,In_360,In_94);
nand U356 (N_356,In_1,In_88);
or U357 (N_357,In_71,In_244);
nor U358 (N_358,In_194,In_479);
nand U359 (N_359,In_588,In_607);
xor U360 (N_360,In_569,In_637);
and U361 (N_361,In_158,In_667);
nor U362 (N_362,In_356,In_265);
xor U363 (N_363,In_577,In_292);
and U364 (N_364,In_540,In_525);
nor U365 (N_365,In_11,In_662);
nor U366 (N_366,In_614,In_118);
xor U367 (N_367,In_556,In_528);
nand U368 (N_368,In_48,In_106);
xor U369 (N_369,In_315,In_188);
or U370 (N_370,In_512,In_638);
or U371 (N_371,In_216,In_523);
and U372 (N_372,In_450,In_341);
xor U373 (N_373,In_36,In_650);
or U374 (N_374,In_541,In_420);
xor U375 (N_375,In_99,In_629);
nand U376 (N_376,In_444,In_300);
or U377 (N_377,In_701,In_363);
nand U378 (N_378,In_578,In_297);
xor U379 (N_379,In_321,In_660);
nand U380 (N_380,In_177,In_262);
or U381 (N_381,In_288,In_446);
or U382 (N_382,In_51,In_176);
xor U383 (N_383,In_11,In_37);
nand U384 (N_384,In_100,In_470);
or U385 (N_385,In_491,In_174);
and U386 (N_386,In_668,In_346);
nand U387 (N_387,In_388,In_482);
nor U388 (N_388,In_615,In_614);
nand U389 (N_389,In_486,In_289);
nand U390 (N_390,In_422,In_354);
nand U391 (N_391,In_229,In_465);
xnor U392 (N_392,In_558,In_710);
nor U393 (N_393,In_375,In_659);
or U394 (N_394,In_723,In_332);
or U395 (N_395,In_479,In_136);
xnor U396 (N_396,In_29,In_584);
and U397 (N_397,In_248,In_208);
nor U398 (N_398,In_594,In_749);
and U399 (N_399,In_128,In_720);
or U400 (N_400,In_575,In_88);
nor U401 (N_401,In_29,In_428);
and U402 (N_402,In_527,In_400);
or U403 (N_403,In_92,In_592);
and U404 (N_404,In_569,In_400);
and U405 (N_405,In_722,In_305);
or U406 (N_406,In_550,In_600);
or U407 (N_407,In_527,In_133);
nor U408 (N_408,In_588,In_246);
and U409 (N_409,In_736,In_90);
or U410 (N_410,In_607,In_38);
nor U411 (N_411,In_11,In_548);
nand U412 (N_412,In_562,In_310);
xnor U413 (N_413,In_159,In_631);
xnor U414 (N_414,In_157,In_195);
xor U415 (N_415,In_33,In_510);
or U416 (N_416,In_614,In_216);
xnor U417 (N_417,In_623,In_323);
and U418 (N_418,In_323,In_39);
xnor U419 (N_419,In_627,In_240);
or U420 (N_420,In_359,In_580);
nand U421 (N_421,In_76,In_678);
nand U422 (N_422,In_38,In_741);
or U423 (N_423,In_391,In_710);
nand U424 (N_424,In_414,In_630);
and U425 (N_425,In_660,In_372);
nand U426 (N_426,In_438,In_745);
xnor U427 (N_427,In_261,In_296);
and U428 (N_428,In_529,In_227);
xnor U429 (N_429,In_547,In_668);
nor U430 (N_430,In_264,In_673);
nand U431 (N_431,In_105,In_219);
or U432 (N_432,In_569,In_712);
nor U433 (N_433,In_108,In_525);
nor U434 (N_434,In_414,In_66);
or U435 (N_435,In_615,In_536);
nand U436 (N_436,In_255,In_294);
nor U437 (N_437,In_368,In_156);
nand U438 (N_438,In_284,In_515);
and U439 (N_439,In_111,In_138);
or U440 (N_440,In_674,In_369);
or U441 (N_441,In_70,In_68);
or U442 (N_442,In_97,In_648);
or U443 (N_443,In_600,In_357);
or U444 (N_444,In_266,In_221);
xor U445 (N_445,In_355,In_264);
nor U446 (N_446,In_630,In_551);
and U447 (N_447,In_102,In_625);
xor U448 (N_448,In_82,In_342);
nand U449 (N_449,In_175,In_598);
and U450 (N_450,In_52,In_561);
nor U451 (N_451,In_575,In_354);
nor U452 (N_452,In_622,In_500);
nand U453 (N_453,In_486,In_176);
or U454 (N_454,In_275,In_120);
nand U455 (N_455,In_578,In_231);
nor U456 (N_456,In_16,In_103);
nand U457 (N_457,In_243,In_738);
xor U458 (N_458,In_91,In_322);
and U459 (N_459,In_532,In_224);
nand U460 (N_460,In_354,In_172);
xnor U461 (N_461,In_454,In_393);
nor U462 (N_462,In_143,In_292);
and U463 (N_463,In_43,In_666);
xnor U464 (N_464,In_195,In_357);
nand U465 (N_465,In_749,In_581);
nor U466 (N_466,In_214,In_306);
nor U467 (N_467,In_716,In_229);
nor U468 (N_468,In_294,In_400);
nand U469 (N_469,In_405,In_542);
nand U470 (N_470,In_109,In_520);
and U471 (N_471,In_724,In_544);
and U472 (N_472,In_342,In_47);
nand U473 (N_473,In_696,In_613);
nor U474 (N_474,In_518,In_423);
nand U475 (N_475,In_180,In_592);
xor U476 (N_476,In_13,In_443);
xnor U477 (N_477,In_351,In_638);
nand U478 (N_478,In_14,In_117);
or U479 (N_479,In_283,In_122);
and U480 (N_480,In_266,In_297);
xor U481 (N_481,In_12,In_722);
and U482 (N_482,In_722,In_233);
or U483 (N_483,In_35,In_536);
xnor U484 (N_484,In_510,In_81);
or U485 (N_485,In_222,In_645);
nor U486 (N_486,In_334,In_369);
and U487 (N_487,In_741,In_374);
and U488 (N_488,In_700,In_622);
xor U489 (N_489,In_481,In_305);
and U490 (N_490,In_418,In_175);
xor U491 (N_491,In_139,In_263);
xor U492 (N_492,In_694,In_459);
nand U493 (N_493,In_616,In_190);
nand U494 (N_494,In_633,In_147);
nor U495 (N_495,In_660,In_8);
or U496 (N_496,In_584,In_83);
nand U497 (N_497,In_735,In_586);
xor U498 (N_498,In_465,In_718);
and U499 (N_499,In_479,In_130);
nor U500 (N_500,In_363,In_432);
nand U501 (N_501,In_29,In_481);
and U502 (N_502,In_419,In_615);
and U503 (N_503,In_11,In_624);
or U504 (N_504,In_435,In_321);
nor U505 (N_505,In_709,In_91);
or U506 (N_506,In_321,In_466);
nor U507 (N_507,In_85,In_595);
xor U508 (N_508,In_275,In_486);
and U509 (N_509,In_416,In_706);
nor U510 (N_510,In_283,In_623);
nor U511 (N_511,In_396,In_666);
and U512 (N_512,In_421,In_96);
or U513 (N_513,In_460,In_447);
or U514 (N_514,In_522,In_21);
xnor U515 (N_515,In_321,In_451);
or U516 (N_516,In_478,In_167);
nor U517 (N_517,In_76,In_290);
nand U518 (N_518,In_32,In_301);
and U519 (N_519,In_206,In_522);
and U520 (N_520,In_4,In_70);
nor U521 (N_521,In_193,In_271);
and U522 (N_522,In_367,In_496);
and U523 (N_523,In_248,In_679);
or U524 (N_524,In_365,In_517);
and U525 (N_525,In_105,In_359);
nor U526 (N_526,In_322,In_189);
nand U527 (N_527,In_656,In_501);
nand U528 (N_528,In_433,In_509);
nor U529 (N_529,In_85,In_699);
xnor U530 (N_530,In_335,In_143);
and U531 (N_531,In_549,In_154);
nor U532 (N_532,In_368,In_698);
xnor U533 (N_533,In_678,In_629);
and U534 (N_534,In_700,In_135);
nor U535 (N_535,In_170,In_105);
or U536 (N_536,In_536,In_403);
xor U537 (N_537,In_284,In_250);
or U538 (N_538,In_343,In_362);
nand U539 (N_539,In_511,In_574);
and U540 (N_540,In_707,In_551);
or U541 (N_541,In_133,In_346);
xnor U542 (N_542,In_392,In_263);
nand U543 (N_543,In_145,In_238);
nand U544 (N_544,In_429,In_661);
nand U545 (N_545,In_312,In_566);
nand U546 (N_546,In_120,In_668);
nor U547 (N_547,In_64,In_226);
nor U548 (N_548,In_44,In_561);
or U549 (N_549,In_468,In_217);
nor U550 (N_550,In_61,In_316);
and U551 (N_551,In_407,In_53);
and U552 (N_552,In_698,In_474);
nor U553 (N_553,In_721,In_428);
or U554 (N_554,In_400,In_385);
and U555 (N_555,In_365,In_635);
xnor U556 (N_556,In_340,In_702);
nand U557 (N_557,In_34,In_484);
xor U558 (N_558,In_325,In_614);
nor U559 (N_559,In_460,In_145);
and U560 (N_560,In_195,In_719);
nand U561 (N_561,In_481,In_635);
xor U562 (N_562,In_499,In_568);
and U563 (N_563,In_313,In_6);
xnor U564 (N_564,In_164,In_284);
nand U565 (N_565,In_325,In_520);
xnor U566 (N_566,In_647,In_89);
nand U567 (N_567,In_693,In_144);
xnor U568 (N_568,In_103,In_445);
nand U569 (N_569,In_209,In_172);
nand U570 (N_570,In_728,In_511);
and U571 (N_571,In_533,In_690);
and U572 (N_572,In_233,In_339);
and U573 (N_573,In_30,In_67);
or U574 (N_574,In_425,In_482);
or U575 (N_575,In_194,In_174);
or U576 (N_576,In_124,In_528);
or U577 (N_577,In_475,In_421);
nand U578 (N_578,In_258,In_377);
or U579 (N_579,In_545,In_28);
and U580 (N_580,In_635,In_448);
or U581 (N_581,In_678,In_201);
xor U582 (N_582,In_258,In_70);
and U583 (N_583,In_253,In_110);
or U584 (N_584,In_115,In_153);
and U585 (N_585,In_73,In_29);
and U586 (N_586,In_320,In_399);
xor U587 (N_587,In_37,In_144);
nor U588 (N_588,In_72,In_655);
and U589 (N_589,In_650,In_737);
nand U590 (N_590,In_522,In_428);
and U591 (N_591,In_326,In_275);
nand U592 (N_592,In_261,In_143);
nor U593 (N_593,In_707,In_415);
xnor U594 (N_594,In_292,In_615);
nor U595 (N_595,In_533,In_302);
and U596 (N_596,In_560,In_295);
nor U597 (N_597,In_103,In_399);
or U598 (N_598,In_498,In_370);
and U599 (N_599,In_650,In_735);
nand U600 (N_600,In_55,In_97);
and U601 (N_601,In_92,In_637);
or U602 (N_602,In_595,In_333);
nor U603 (N_603,In_621,In_320);
and U604 (N_604,In_47,In_585);
nor U605 (N_605,In_411,In_300);
xnor U606 (N_606,In_231,In_548);
or U607 (N_607,In_469,In_341);
xor U608 (N_608,In_161,In_125);
or U609 (N_609,In_678,In_504);
and U610 (N_610,In_699,In_618);
nor U611 (N_611,In_569,In_85);
or U612 (N_612,In_126,In_260);
nand U613 (N_613,In_93,In_330);
or U614 (N_614,In_462,In_631);
xnor U615 (N_615,In_342,In_549);
nand U616 (N_616,In_447,In_310);
and U617 (N_617,In_390,In_154);
nand U618 (N_618,In_60,In_694);
xor U619 (N_619,In_745,In_737);
or U620 (N_620,In_30,In_556);
nor U621 (N_621,In_75,In_29);
or U622 (N_622,In_97,In_58);
xnor U623 (N_623,In_630,In_666);
or U624 (N_624,In_311,In_712);
and U625 (N_625,In_331,In_593);
and U626 (N_626,In_328,In_443);
xnor U627 (N_627,In_60,In_713);
and U628 (N_628,In_355,In_319);
and U629 (N_629,In_722,In_176);
and U630 (N_630,In_293,In_40);
xor U631 (N_631,In_228,In_725);
or U632 (N_632,In_673,In_424);
and U633 (N_633,In_379,In_573);
xnor U634 (N_634,In_533,In_650);
nand U635 (N_635,In_477,In_109);
nor U636 (N_636,In_352,In_498);
and U637 (N_637,In_589,In_604);
or U638 (N_638,In_189,In_125);
nand U639 (N_639,In_250,In_244);
or U640 (N_640,In_219,In_13);
or U641 (N_641,In_175,In_203);
or U642 (N_642,In_563,In_426);
or U643 (N_643,In_383,In_276);
or U644 (N_644,In_288,In_115);
and U645 (N_645,In_447,In_364);
nand U646 (N_646,In_660,In_545);
nand U647 (N_647,In_140,In_656);
nor U648 (N_648,In_742,In_543);
nor U649 (N_649,In_378,In_107);
and U650 (N_650,In_363,In_395);
nand U651 (N_651,In_513,In_205);
nor U652 (N_652,In_254,In_612);
or U653 (N_653,In_35,In_116);
nor U654 (N_654,In_394,In_330);
or U655 (N_655,In_636,In_64);
nor U656 (N_656,In_253,In_167);
xnor U657 (N_657,In_463,In_311);
nand U658 (N_658,In_291,In_63);
and U659 (N_659,In_9,In_261);
nand U660 (N_660,In_241,In_645);
nand U661 (N_661,In_39,In_370);
nor U662 (N_662,In_639,In_97);
nor U663 (N_663,In_186,In_545);
and U664 (N_664,In_502,In_549);
or U665 (N_665,In_548,In_290);
xor U666 (N_666,In_226,In_48);
or U667 (N_667,In_599,In_591);
nand U668 (N_668,In_253,In_749);
and U669 (N_669,In_492,In_498);
and U670 (N_670,In_575,In_353);
or U671 (N_671,In_339,In_545);
xor U672 (N_672,In_571,In_572);
or U673 (N_673,In_130,In_105);
and U674 (N_674,In_284,In_724);
or U675 (N_675,In_50,In_359);
nor U676 (N_676,In_340,In_616);
and U677 (N_677,In_86,In_669);
and U678 (N_678,In_441,In_156);
or U679 (N_679,In_546,In_131);
nor U680 (N_680,In_450,In_157);
xor U681 (N_681,In_518,In_84);
xnor U682 (N_682,In_267,In_414);
nand U683 (N_683,In_175,In_622);
xnor U684 (N_684,In_532,In_450);
nand U685 (N_685,In_558,In_251);
xnor U686 (N_686,In_418,In_388);
xnor U687 (N_687,In_109,In_647);
or U688 (N_688,In_588,In_687);
nand U689 (N_689,In_655,In_508);
xor U690 (N_690,In_632,In_656);
xnor U691 (N_691,In_0,In_412);
nand U692 (N_692,In_171,In_262);
and U693 (N_693,In_459,In_256);
nor U694 (N_694,In_213,In_618);
nand U695 (N_695,In_424,In_333);
nor U696 (N_696,In_467,In_43);
xor U697 (N_697,In_233,In_683);
or U698 (N_698,In_9,In_735);
and U699 (N_699,In_260,In_244);
or U700 (N_700,In_714,In_223);
and U701 (N_701,In_412,In_596);
and U702 (N_702,In_473,In_396);
nor U703 (N_703,In_221,In_146);
nand U704 (N_704,In_477,In_103);
and U705 (N_705,In_86,In_225);
xnor U706 (N_706,In_304,In_306);
and U707 (N_707,In_260,In_720);
and U708 (N_708,In_228,In_339);
xor U709 (N_709,In_260,In_295);
xnor U710 (N_710,In_19,In_9);
nand U711 (N_711,In_188,In_683);
nor U712 (N_712,In_454,In_476);
nand U713 (N_713,In_3,In_225);
or U714 (N_714,In_284,In_720);
or U715 (N_715,In_293,In_93);
xor U716 (N_716,In_635,In_226);
nor U717 (N_717,In_448,In_400);
nand U718 (N_718,In_132,In_584);
nor U719 (N_719,In_25,In_674);
nand U720 (N_720,In_531,In_45);
or U721 (N_721,In_705,In_645);
nand U722 (N_722,In_506,In_347);
and U723 (N_723,In_368,In_243);
and U724 (N_724,In_525,In_599);
nand U725 (N_725,In_145,In_22);
and U726 (N_726,In_561,In_8);
and U727 (N_727,In_300,In_340);
nor U728 (N_728,In_453,In_604);
nand U729 (N_729,In_51,In_207);
xor U730 (N_730,In_469,In_269);
or U731 (N_731,In_537,In_433);
nand U732 (N_732,In_658,In_79);
nand U733 (N_733,In_222,In_44);
and U734 (N_734,In_434,In_307);
xor U735 (N_735,In_727,In_142);
nand U736 (N_736,In_733,In_592);
xnor U737 (N_737,In_735,In_690);
and U738 (N_738,In_213,In_307);
nand U739 (N_739,In_132,In_332);
nor U740 (N_740,In_1,In_561);
nand U741 (N_741,In_652,In_626);
nand U742 (N_742,In_429,In_344);
and U743 (N_743,In_644,In_431);
xor U744 (N_744,In_259,In_622);
nor U745 (N_745,In_547,In_105);
and U746 (N_746,In_278,In_684);
and U747 (N_747,In_430,In_249);
xnor U748 (N_748,In_562,In_418);
nor U749 (N_749,In_460,In_571);
or U750 (N_750,In_583,In_343);
or U751 (N_751,In_695,In_237);
xor U752 (N_752,In_424,In_87);
nand U753 (N_753,In_6,In_418);
or U754 (N_754,In_710,In_108);
and U755 (N_755,In_738,In_688);
xnor U756 (N_756,In_16,In_701);
xnor U757 (N_757,In_619,In_98);
nor U758 (N_758,In_741,In_224);
xnor U759 (N_759,In_41,In_450);
and U760 (N_760,In_577,In_456);
or U761 (N_761,In_397,In_636);
nand U762 (N_762,In_204,In_623);
xnor U763 (N_763,In_146,In_389);
nand U764 (N_764,In_111,In_291);
nand U765 (N_765,In_353,In_246);
and U766 (N_766,In_472,In_313);
nand U767 (N_767,In_14,In_238);
or U768 (N_768,In_463,In_64);
or U769 (N_769,In_592,In_729);
nand U770 (N_770,In_204,In_100);
or U771 (N_771,In_502,In_57);
nor U772 (N_772,In_685,In_581);
nor U773 (N_773,In_553,In_395);
xnor U774 (N_774,In_472,In_243);
or U775 (N_775,In_143,In_589);
nor U776 (N_776,In_356,In_309);
xnor U777 (N_777,In_321,In_470);
xor U778 (N_778,In_581,In_491);
and U779 (N_779,In_195,In_33);
nand U780 (N_780,In_719,In_186);
nand U781 (N_781,In_285,In_106);
and U782 (N_782,In_93,In_252);
nor U783 (N_783,In_140,In_322);
nor U784 (N_784,In_283,In_727);
or U785 (N_785,In_453,In_496);
or U786 (N_786,In_352,In_544);
nand U787 (N_787,In_650,In_200);
xnor U788 (N_788,In_446,In_738);
nor U789 (N_789,In_338,In_414);
or U790 (N_790,In_433,In_511);
xor U791 (N_791,In_36,In_451);
nor U792 (N_792,In_137,In_85);
xnor U793 (N_793,In_399,In_187);
and U794 (N_794,In_159,In_635);
nand U795 (N_795,In_363,In_617);
nor U796 (N_796,In_472,In_290);
nor U797 (N_797,In_637,In_680);
nand U798 (N_798,In_77,In_119);
and U799 (N_799,In_447,In_506);
nor U800 (N_800,In_715,In_200);
nor U801 (N_801,In_72,In_523);
and U802 (N_802,In_705,In_84);
and U803 (N_803,In_45,In_97);
nand U804 (N_804,In_702,In_507);
nand U805 (N_805,In_169,In_23);
and U806 (N_806,In_540,In_573);
nor U807 (N_807,In_640,In_146);
nor U808 (N_808,In_494,In_706);
xor U809 (N_809,In_635,In_456);
xor U810 (N_810,In_519,In_592);
nand U811 (N_811,In_269,In_373);
xor U812 (N_812,In_690,In_634);
or U813 (N_813,In_180,In_131);
xor U814 (N_814,In_164,In_179);
nand U815 (N_815,In_592,In_678);
xor U816 (N_816,In_228,In_397);
and U817 (N_817,In_297,In_170);
or U818 (N_818,In_168,In_183);
nor U819 (N_819,In_392,In_64);
nand U820 (N_820,In_233,In_632);
xor U821 (N_821,In_117,In_647);
or U822 (N_822,In_213,In_590);
or U823 (N_823,In_21,In_513);
and U824 (N_824,In_283,In_93);
and U825 (N_825,In_102,In_342);
nor U826 (N_826,In_94,In_83);
nand U827 (N_827,In_568,In_519);
or U828 (N_828,In_601,In_620);
or U829 (N_829,In_139,In_294);
xor U830 (N_830,In_160,In_731);
xor U831 (N_831,In_743,In_208);
nor U832 (N_832,In_272,In_651);
or U833 (N_833,In_200,In_488);
xor U834 (N_834,In_58,In_52);
or U835 (N_835,In_425,In_616);
or U836 (N_836,In_243,In_113);
xnor U837 (N_837,In_334,In_141);
and U838 (N_838,In_208,In_259);
or U839 (N_839,In_487,In_455);
nor U840 (N_840,In_474,In_615);
nand U841 (N_841,In_16,In_474);
and U842 (N_842,In_370,In_49);
and U843 (N_843,In_530,In_568);
nor U844 (N_844,In_196,In_663);
xnor U845 (N_845,In_272,In_209);
nand U846 (N_846,In_486,In_320);
xnor U847 (N_847,In_201,In_135);
and U848 (N_848,In_271,In_145);
nand U849 (N_849,In_230,In_682);
xor U850 (N_850,In_702,In_165);
and U851 (N_851,In_201,In_241);
nor U852 (N_852,In_664,In_304);
xor U853 (N_853,In_152,In_16);
and U854 (N_854,In_283,In_291);
xnor U855 (N_855,In_576,In_185);
and U856 (N_856,In_662,In_547);
nand U857 (N_857,In_21,In_482);
or U858 (N_858,In_340,In_681);
and U859 (N_859,In_306,In_35);
nand U860 (N_860,In_298,In_28);
or U861 (N_861,In_199,In_358);
or U862 (N_862,In_177,In_541);
or U863 (N_863,In_33,In_70);
or U864 (N_864,In_260,In_583);
nor U865 (N_865,In_155,In_565);
nand U866 (N_866,In_157,In_182);
nand U867 (N_867,In_280,In_715);
xor U868 (N_868,In_224,In_222);
nor U869 (N_869,In_260,In_494);
xnor U870 (N_870,In_269,In_132);
and U871 (N_871,In_388,In_139);
and U872 (N_872,In_353,In_689);
nand U873 (N_873,In_620,In_307);
nor U874 (N_874,In_608,In_632);
or U875 (N_875,In_654,In_413);
and U876 (N_876,In_86,In_695);
or U877 (N_877,In_192,In_561);
nand U878 (N_878,In_295,In_372);
and U879 (N_879,In_737,In_239);
nand U880 (N_880,In_564,In_68);
nand U881 (N_881,In_709,In_503);
or U882 (N_882,In_424,In_677);
or U883 (N_883,In_143,In_259);
nand U884 (N_884,In_704,In_613);
xor U885 (N_885,In_199,In_555);
and U886 (N_886,In_461,In_274);
xor U887 (N_887,In_698,In_460);
or U888 (N_888,In_347,In_373);
nor U889 (N_889,In_212,In_429);
nor U890 (N_890,In_114,In_266);
nor U891 (N_891,In_662,In_256);
and U892 (N_892,In_361,In_237);
or U893 (N_893,In_24,In_546);
and U894 (N_894,In_672,In_263);
xor U895 (N_895,In_292,In_201);
or U896 (N_896,In_617,In_45);
xor U897 (N_897,In_89,In_333);
or U898 (N_898,In_650,In_546);
nor U899 (N_899,In_288,In_433);
and U900 (N_900,In_367,In_433);
nand U901 (N_901,In_290,In_171);
nand U902 (N_902,In_392,In_192);
nor U903 (N_903,In_97,In_567);
or U904 (N_904,In_339,In_43);
or U905 (N_905,In_174,In_724);
or U906 (N_906,In_129,In_132);
and U907 (N_907,In_573,In_694);
nand U908 (N_908,In_668,In_73);
nand U909 (N_909,In_425,In_640);
nor U910 (N_910,In_606,In_247);
and U911 (N_911,In_417,In_165);
nor U912 (N_912,In_37,In_192);
and U913 (N_913,In_98,In_78);
nor U914 (N_914,In_377,In_665);
nand U915 (N_915,In_544,In_723);
and U916 (N_916,In_725,In_695);
or U917 (N_917,In_199,In_225);
xor U918 (N_918,In_277,In_330);
nand U919 (N_919,In_383,In_635);
xor U920 (N_920,In_525,In_60);
or U921 (N_921,In_264,In_698);
and U922 (N_922,In_197,In_163);
and U923 (N_923,In_441,In_504);
and U924 (N_924,In_535,In_110);
or U925 (N_925,In_430,In_737);
nor U926 (N_926,In_246,In_554);
xnor U927 (N_927,In_137,In_362);
and U928 (N_928,In_292,In_294);
or U929 (N_929,In_205,In_74);
or U930 (N_930,In_47,In_285);
or U931 (N_931,In_641,In_672);
or U932 (N_932,In_640,In_128);
or U933 (N_933,In_610,In_338);
nor U934 (N_934,In_650,In_183);
nand U935 (N_935,In_474,In_265);
and U936 (N_936,In_620,In_105);
nor U937 (N_937,In_507,In_619);
nor U938 (N_938,In_231,In_588);
and U939 (N_939,In_628,In_432);
or U940 (N_940,In_549,In_505);
or U941 (N_941,In_224,In_463);
xnor U942 (N_942,In_209,In_481);
or U943 (N_943,In_299,In_469);
nor U944 (N_944,In_534,In_346);
and U945 (N_945,In_447,In_290);
and U946 (N_946,In_123,In_199);
xnor U947 (N_947,In_621,In_515);
and U948 (N_948,In_85,In_106);
nor U949 (N_949,In_152,In_499);
xnor U950 (N_950,In_290,In_605);
or U951 (N_951,In_9,In_393);
and U952 (N_952,In_98,In_572);
nor U953 (N_953,In_248,In_133);
or U954 (N_954,In_637,In_643);
xnor U955 (N_955,In_679,In_337);
nand U956 (N_956,In_377,In_549);
nor U957 (N_957,In_16,In_297);
nor U958 (N_958,In_512,In_585);
nor U959 (N_959,In_91,In_580);
or U960 (N_960,In_457,In_64);
nor U961 (N_961,In_662,In_105);
nand U962 (N_962,In_721,In_142);
or U963 (N_963,In_29,In_576);
nor U964 (N_964,In_555,In_729);
nand U965 (N_965,In_120,In_431);
or U966 (N_966,In_236,In_333);
nor U967 (N_967,In_661,In_484);
or U968 (N_968,In_47,In_63);
nor U969 (N_969,In_181,In_570);
or U970 (N_970,In_624,In_108);
nor U971 (N_971,In_104,In_502);
nor U972 (N_972,In_112,In_562);
and U973 (N_973,In_259,In_198);
or U974 (N_974,In_735,In_687);
or U975 (N_975,In_575,In_264);
nor U976 (N_976,In_265,In_482);
nor U977 (N_977,In_298,In_250);
nand U978 (N_978,In_479,In_638);
or U979 (N_979,In_562,In_677);
and U980 (N_980,In_2,In_394);
nor U981 (N_981,In_504,In_228);
and U982 (N_982,In_585,In_274);
nor U983 (N_983,In_44,In_311);
xor U984 (N_984,In_276,In_163);
xnor U985 (N_985,In_290,In_220);
and U986 (N_986,In_356,In_287);
nor U987 (N_987,In_305,In_279);
and U988 (N_988,In_42,In_59);
or U989 (N_989,In_415,In_203);
nand U990 (N_990,In_434,In_579);
and U991 (N_991,In_18,In_193);
or U992 (N_992,In_180,In_101);
nand U993 (N_993,In_38,In_106);
and U994 (N_994,In_675,In_603);
nand U995 (N_995,In_199,In_296);
or U996 (N_996,In_658,In_652);
nand U997 (N_997,In_292,In_50);
xor U998 (N_998,In_526,In_747);
nand U999 (N_999,In_326,In_565);
and U1000 (N_1000,In_626,In_672);
nor U1001 (N_1001,In_176,In_526);
xnor U1002 (N_1002,In_562,In_56);
xor U1003 (N_1003,In_123,In_251);
xor U1004 (N_1004,In_669,In_552);
nand U1005 (N_1005,In_476,In_555);
xnor U1006 (N_1006,In_260,In_411);
xor U1007 (N_1007,In_457,In_346);
and U1008 (N_1008,In_43,In_33);
nand U1009 (N_1009,In_748,In_4);
nor U1010 (N_1010,In_379,In_698);
xor U1011 (N_1011,In_35,In_663);
xor U1012 (N_1012,In_403,In_514);
or U1013 (N_1013,In_735,In_246);
and U1014 (N_1014,In_292,In_69);
and U1015 (N_1015,In_289,In_207);
xor U1016 (N_1016,In_72,In_327);
nand U1017 (N_1017,In_54,In_583);
and U1018 (N_1018,In_584,In_399);
nand U1019 (N_1019,In_241,In_445);
and U1020 (N_1020,In_416,In_699);
nor U1021 (N_1021,In_429,In_485);
and U1022 (N_1022,In_260,In_678);
or U1023 (N_1023,In_244,In_695);
or U1024 (N_1024,In_255,In_167);
nor U1025 (N_1025,In_520,In_162);
xnor U1026 (N_1026,In_480,In_688);
nor U1027 (N_1027,In_275,In_609);
nand U1028 (N_1028,In_88,In_26);
nor U1029 (N_1029,In_309,In_693);
nor U1030 (N_1030,In_341,In_746);
xnor U1031 (N_1031,In_14,In_662);
or U1032 (N_1032,In_2,In_742);
nor U1033 (N_1033,In_210,In_429);
nand U1034 (N_1034,In_384,In_233);
nand U1035 (N_1035,In_548,In_102);
nand U1036 (N_1036,In_466,In_480);
xnor U1037 (N_1037,In_435,In_735);
xnor U1038 (N_1038,In_32,In_499);
or U1039 (N_1039,In_308,In_489);
xnor U1040 (N_1040,In_608,In_327);
nor U1041 (N_1041,In_415,In_456);
or U1042 (N_1042,In_599,In_369);
or U1043 (N_1043,In_371,In_581);
xor U1044 (N_1044,In_321,In_744);
or U1045 (N_1045,In_77,In_745);
or U1046 (N_1046,In_253,In_41);
and U1047 (N_1047,In_392,In_399);
nor U1048 (N_1048,In_357,In_150);
nor U1049 (N_1049,In_378,In_445);
and U1050 (N_1050,In_70,In_314);
xnor U1051 (N_1051,In_677,In_492);
or U1052 (N_1052,In_711,In_18);
nand U1053 (N_1053,In_713,In_352);
or U1054 (N_1054,In_88,In_558);
and U1055 (N_1055,In_307,In_32);
nand U1056 (N_1056,In_467,In_166);
or U1057 (N_1057,In_476,In_489);
nor U1058 (N_1058,In_368,In_345);
xnor U1059 (N_1059,In_145,In_481);
nand U1060 (N_1060,In_65,In_241);
nand U1061 (N_1061,In_395,In_35);
nor U1062 (N_1062,In_639,In_12);
nand U1063 (N_1063,In_568,In_539);
or U1064 (N_1064,In_521,In_235);
nand U1065 (N_1065,In_124,In_299);
and U1066 (N_1066,In_548,In_339);
xnor U1067 (N_1067,In_119,In_105);
xnor U1068 (N_1068,In_102,In_10);
nor U1069 (N_1069,In_498,In_622);
nor U1070 (N_1070,In_74,In_705);
nor U1071 (N_1071,In_665,In_680);
and U1072 (N_1072,In_338,In_714);
nand U1073 (N_1073,In_96,In_181);
nor U1074 (N_1074,In_563,In_742);
xnor U1075 (N_1075,In_704,In_304);
or U1076 (N_1076,In_625,In_454);
nand U1077 (N_1077,In_469,In_470);
nand U1078 (N_1078,In_604,In_137);
or U1079 (N_1079,In_90,In_367);
xnor U1080 (N_1080,In_592,In_745);
or U1081 (N_1081,In_513,In_18);
or U1082 (N_1082,In_339,In_559);
xnor U1083 (N_1083,In_727,In_160);
xnor U1084 (N_1084,In_99,In_243);
nand U1085 (N_1085,In_367,In_696);
or U1086 (N_1086,In_666,In_511);
and U1087 (N_1087,In_409,In_733);
nand U1088 (N_1088,In_80,In_425);
nor U1089 (N_1089,In_54,In_299);
nor U1090 (N_1090,In_671,In_659);
nor U1091 (N_1091,In_551,In_570);
nand U1092 (N_1092,In_694,In_333);
nor U1093 (N_1093,In_518,In_67);
nor U1094 (N_1094,In_699,In_242);
xnor U1095 (N_1095,In_406,In_523);
or U1096 (N_1096,In_190,In_218);
nand U1097 (N_1097,In_294,In_0);
and U1098 (N_1098,In_157,In_236);
and U1099 (N_1099,In_624,In_66);
nand U1100 (N_1100,In_191,In_692);
or U1101 (N_1101,In_561,In_400);
nor U1102 (N_1102,In_134,In_546);
nand U1103 (N_1103,In_504,In_674);
nor U1104 (N_1104,In_223,In_319);
xor U1105 (N_1105,In_119,In_469);
nand U1106 (N_1106,In_410,In_717);
or U1107 (N_1107,In_550,In_296);
or U1108 (N_1108,In_738,In_11);
nand U1109 (N_1109,In_302,In_739);
xnor U1110 (N_1110,In_53,In_342);
or U1111 (N_1111,In_260,In_537);
xnor U1112 (N_1112,In_194,In_530);
nand U1113 (N_1113,In_70,In_360);
or U1114 (N_1114,In_548,In_699);
nor U1115 (N_1115,In_54,In_649);
nor U1116 (N_1116,In_726,In_554);
and U1117 (N_1117,In_233,In_26);
or U1118 (N_1118,In_595,In_68);
nor U1119 (N_1119,In_643,In_152);
nor U1120 (N_1120,In_21,In_142);
nand U1121 (N_1121,In_677,In_253);
or U1122 (N_1122,In_278,In_162);
nor U1123 (N_1123,In_659,In_59);
nor U1124 (N_1124,In_287,In_662);
and U1125 (N_1125,In_628,In_490);
and U1126 (N_1126,In_147,In_267);
and U1127 (N_1127,In_547,In_65);
nand U1128 (N_1128,In_670,In_317);
nand U1129 (N_1129,In_143,In_640);
or U1130 (N_1130,In_457,In_248);
or U1131 (N_1131,In_74,In_12);
or U1132 (N_1132,In_170,In_551);
xnor U1133 (N_1133,In_452,In_450);
or U1134 (N_1134,In_359,In_219);
nand U1135 (N_1135,In_83,In_299);
xor U1136 (N_1136,In_620,In_114);
and U1137 (N_1137,In_380,In_189);
xnor U1138 (N_1138,In_349,In_655);
xnor U1139 (N_1139,In_120,In_554);
and U1140 (N_1140,In_383,In_524);
xnor U1141 (N_1141,In_677,In_205);
nand U1142 (N_1142,In_86,In_207);
nand U1143 (N_1143,In_40,In_187);
nand U1144 (N_1144,In_324,In_321);
nor U1145 (N_1145,In_360,In_394);
nor U1146 (N_1146,In_188,In_529);
or U1147 (N_1147,In_568,In_450);
nor U1148 (N_1148,In_413,In_37);
xor U1149 (N_1149,In_54,In_611);
nand U1150 (N_1150,In_666,In_300);
xor U1151 (N_1151,In_134,In_278);
nand U1152 (N_1152,In_547,In_716);
nand U1153 (N_1153,In_338,In_507);
and U1154 (N_1154,In_731,In_621);
nor U1155 (N_1155,In_539,In_255);
and U1156 (N_1156,In_432,In_463);
xor U1157 (N_1157,In_111,In_200);
xnor U1158 (N_1158,In_352,In_505);
and U1159 (N_1159,In_360,In_455);
xor U1160 (N_1160,In_192,In_93);
nor U1161 (N_1161,In_337,In_397);
nor U1162 (N_1162,In_411,In_279);
nor U1163 (N_1163,In_480,In_90);
nand U1164 (N_1164,In_553,In_381);
xnor U1165 (N_1165,In_503,In_531);
xnor U1166 (N_1166,In_381,In_15);
or U1167 (N_1167,In_705,In_13);
nand U1168 (N_1168,In_402,In_697);
nand U1169 (N_1169,In_250,In_469);
or U1170 (N_1170,In_264,In_201);
or U1171 (N_1171,In_434,In_140);
nand U1172 (N_1172,In_27,In_204);
and U1173 (N_1173,In_703,In_509);
nor U1174 (N_1174,In_60,In_444);
nor U1175 (N_1175,In_383,In_495);
xor U1176 (N_1176,In_602,In_402);
xor U1177 (N_1177,In_535,In_347);
nor U1178 (N_1178,In_1,In_343);
nor U1179 (N_1179,In_343,In_672);
xor U1180 (N_1180,In_307,In_82);
nand U1181 (N_1181,In_60,In_215);
or U1182 (N_1182,In_310,In_265);
xnor U1183 (N_1183,In_644,In_560);
xor U1184 (N_1184,In_737,In_327);
xnor U1185 (N_1185,In_160,In_269);
xnor U1186 (N_1186,In_186,In_284);
or U1187 (N_1187,In_130,In_238);
or U1188 (N_1188,In_484,In_226);
nand U1189 (N_1189,In_419,In_552);
nand U1190 (N_1190,In_380,In_557);
and U1191 (N_1191,In_240,In_626);
or U1192 (N_1192,In_412,In_400);
nand U1193 (N_1193,In_581,In_266);
or U1194 (N_1194,In_252,In_157);
or U1195 (N_1195,In_419,In_171);
and U1196 (N_1196,In_329,In_336);
and U1197 (N_1197,In_266,In_162);
xnor U1198 (N_1198,In_713,In_268);
nand U1199 (N_1199,In_710,In_132);
xor U1200 (N_1200,In_544,In_446);
nor U1201 (N_1201,In_189,In_372);
nand U1202 (N_1202,In_498,In_58);
xor U1203 (N_1203,In_734,In_428);
and U1204 (N_1204,In_58,In_62);
or U1205 (N_1205,In_582,In_538);
nand U1206 (N_1206,In_634,In_466);
or U1207 (N_1207,In_532,In_111);
nor U1208 (N_1208,In_560,In_20);
nor U1209 (N_1209,In_83,In_195);
xnor U1210 (N_1210,In_736,In_487);
and U1211 (N_1211,In_387,In_14);
xnor U1212 (N_1212,In_717,In_261);
and U1213 (N_1213,In_466,In_311);
or U1214 (N_1214,In_394,In_69);
nand U1215 (N_1215,In_507,In_725);
or U1216 (N_1216,In_355,In_638);
nand U1217 (N_1217,In_536,In_715);
xor U1218 (N_1218,In_414,In_572);
and U1219 (N_1219,In_279,In_208);
nor U1220 (N_1220,In_210,In_38);
nand U1221 (N_1221,In_369,In_729);
and U1222 (N_1222,In_520,In_99);
xnor U1223 (N_1223,In_203,In_12);
xor U1224 (N_1224,In_556,In_707);
nor U1225 (N_1225,In_405,In_558);
nand U1226 (N_1226,In_303,In_321);
or U1227 (N_1227,In_188,In_338);
and U1228 (N_1228,In_293,In_713);
or U1229 (N_1229,In_496,In_154);
or U1230 (N_1230,In_559,In_734);
nor U1231 (N_1231,In_79,In_201);
nand U1232 (N_1232,In_145,In_253);
nor U1233 (N_1233,In_532,In_660);
and U1234 (N_1234,In_466,In_727);
nor U1235 (N_1235,In_548,In_302);
or U1236 (N_1236,In_240,In_382);
or U1237 (N_1237,In_746,In_251);
or U1238 (N_1238,In_656,In_607);
xnor U1239 (N_1239,In_608,In_168);
or U1240 (N_1240,In_616,In_746);
or U1241 (N_1241,In_585,In_1);
nor U1242 (N_1242,In_663,In_115);
and U1243 (N_1243,In_104,In_618);
nor U1244 (N_1244,In_100,In_618);
nor U1245 (N_1245,In_89,In_121);
nor U1246 (N_1246,In_648,In_607);
and U1247 (N_1247,In_142,In_732);
and U1248 (N_1248,In_504,In_722);
nand U1249 (N_1249,In_534,In_562);
nand U1250 (N_1250,In_67,In_9);
nor U1251 (N_1251,In_357,In_710);
or U1252 (N_1252,In_75,In_81);
nor U1253 (N_1253,In_287,In_584);
and U1254 (N_1254,In_652,In_34);
xnor U1255 (N_1255,In_364,In_459);
nand U1256 (N_1256,In_280,In_625);
or U1257 (N_1257,In_538,In_539);
or U1258 (N_1258,In_5,In_286);
nor U1259 (N_1259,In_386,In_337);
or U1260 (N_1260,In_254,In_293);
nor U1261 (N_1261,In_586,In_80);
nor U1262 (N_1262,In_239,In_749);
nor U1263 (N_1263,In_377,In_161);
nor U1264 (N_1264,In_550,In_140);
or U1265 (N_1265,In_172,In_63);
and U1266 (N_1266,In_471,In_720);
or U1267 (N_1267,In_476,In_35);
nor U1268 (N_1268,In_458,In_201);
and U1269 (N_1269,In_260,In_415);
and U1270 (N_1270,In_500,In_494);
or U1271 (N_1271,In_393,In_35);
and U1272 (N_1272,In_724,In_681);
xnor U1273 (N_1273,In_48,In_497);
xor U1274 (N_1274,In_210,In_630);
nand U1275 (N_1275,In_199,In_534);
xnor U1276 (N_1276,In_533,In_175);
or U1277 (N_1277,In_713,In_427);
nand U1278 (N_1278,In_116,In_748);
xnor U1279 (N_1279,In_36,In_386);
nor U1280 (N_1280,In_722,In_296);
nand U1281 (N_1281,In_97,In_318);
or U1282 (N_1282,In_382,In_300);
xor U1283 (N_1283,In_63,In_162);
and U1284 (N_1284,In_742,In_560);
and U1285 (N_1285,In_435,In_208);
and U1286 (N_1286,In_449,In_377);
and U1287 (N_1287,In_616,In_310);
or U1288 (N_1288,In_583,In_12);
nor U1289 (N_1289,In_369,In_264);
nor U1290 (N_1290,In_223,In_603);
xor U1291 (N_1291,In_599,In_551);
or U1292 (N_1292,In_427,In_691);
nand U1293 (N_1293,In_470,In_305);
or U1294 (N_1294,In_6,In_612);
nand U1295 (N_1295,In_702,In_654);
and U1296 (N_1296,In_489,In_299);
or U1297 (N_1297,In_450,In_600);
xnor U1298 (N_1298,In_377,In_640);
nand U1299 (N_1299,In_500,In_150);
xnor U1300 (N_1300,In_149,In_733);
nand U1301 (N_1301,In_587,In_335);
or U1302 (N_1302,In_392,In_321);
and U1303 (N_1303,In_28,In_370);
nor U1304 (N_1304,In_157,In_241);
and U1305 (N_1305,In_302,In_161);
nand U1306 (N_1306,In_226,In_307);
nand U1307 (N_1307,In_338,In_110);
nand U1308 (N_1308,In_128,In_431);
or U1309 (N_1309,In_173,In_545);
and U1310 (N_1310,In_75,In_203);
nand U1311 (N_1311,In_303,In_386);
nor U1312 (N_1312,In_688,In_95);
nand U1313 (N_1313,In_398,In_233);
xnor U1314 (N_1314,In_10,In_615);
and U1315 (N_1315,In_575,In_178);
nor U1316 (N_1316,In_7,In_12);
nand U1317 (N_1317,In_637,In_241);
nand U1318 (N_1318,In_37,In_308);
xnor U1319 (N_1319,In_344,In_300);
nand U1320 (N_1320,In_275,In_363);
nand U1321 (N_1321,In_735,In_310);
xor U1322 (N_1322,In_669,In_345);
or U1323 (N_1323,In_401,In_128);
nand U1324 (N_1324,In_263,In_730);
nand U1325 (N_1325,In_321,In_385);
nand U1326 (N_1326,In_618,In_206);
nor U1327 (N_1327,In_402,In_640);
or U1328 (N_1328,In_205,In_554);
nand U1329 (N_1329,In_584,In_613);
and U1330 (N_1330,In_515,In_546);
xnor U1331 (N_1331,In_320,In_90);
nand U1332 (N_1332,In_471,In_82);
or U1333 (N_1333,In_644,In_196);
or U1334 (N_1334,In_493,In_4);
or U1335 (N_1335,In_346,In_564);
or U1336 (N_1336,In_12,In_320);
and U1337 (N_1337,In_512,In_628);
xor U1338 (N_1338,In_633,In_638);
and U1339 (N_1339,In_502,In_64);
and U1340 (N_1340,In_716,In_677);
xnor U1341 (N_1341,In_370,In_449);
or U1342 (N_1342,In_236,In_381);
nor U1343 (N_1343,In_503,In_559);
nor U1344 (N_1344,In_386,In_489);
xnor U1345 (N_1345,In_720,In_164);
and U1346 (N_1346,In_449,In_434);
and U1347 (N_1347,In_220,In_79);
or U1348 (N_1348,In_735,In_222);
nor U1349 (N_1349,In_451,In_364);
nand U1350 (N_1350,In_355,In_158);
and U1351 (N_1351,In_627,In_283);
and U1352 (N_1352,In_198,In_505);
xnor U1353 (N_1353,In_517,In_383);
or U1354 (N_1354,In_323,In_97);
and U1355 (N_1355,In_535,In_198);
nor U1356 (N_1356,In_474,In_14);
nor U1357 (N_1357,In_224,In_604);
and U1358 (N_1358,In_282,In_351);
xnor U1359 (N_1359,In_542,In_196);
xnor U1360 (N_1360,In_170,In_747);
and U1361 (N_1361,In_560,In_719);
nor U1362 (N_1362,In_44,In_346);
nor U1363 (N_1363,In_36,In_202);
nor U1364 (N_1364,In_387,In_214);
nor U1365 (N_1365,In_665,In_654);
xor U1366 (N_1366,In_590,In_596);
xor U1367 (N_1367,In_408,In_465);
nand U1368 (N_1368,In_24,In_101);
or U1369 (N_1369,In_399,In_665);
xor U1370 (N_1370,In_278,In_676);
and U1371 (N_1371,In_13,In_252);
and U1372 (N_1372,In_268,In_336);
nor U1373 (N_1373,In_405,In_61);
xnor U1374 (N_1374,In_75,In_196);
nand U1375 (N_1375,In_717,In_182);
xnor U1376 (N_1376,In_552,In_673);
nor U1377 (N_1377,In_106,In_172);
nand U1378 (N_1378,In_250,In_229);
or U1379 (N_1379,In_480,In_193);
and U1380 (N_1380,In_119,In_116);
nand U1381 (N_1381,In_426,In_542);
nand U1382 (N_1382,In_209,In_539);
or U1383 (N_1383,In_535,In_404);
nor U1384 (N_1384,In_607,In_674);
nand U1385 (N_1385,In_727,In_552);
and U1386 (N_1386,In_303,In_283);
or U1387 (N_1387,In_742,In_53);
nand U1388 (N_1388,In_723,In_679);
nand U1389 (N_1389,In_250,In_452);
nand U1390 (N_1390,In_58,In_216);
nand U1391 (N_1391,In_119,In_9);
or U1392 (N_1392,In_584,In_27);
nor U1393 (N_1393,In_96,In_606);
nand U1394 (N_1394,In_365,In_115);
xor U1395 (N_1395,In_264,In_393);
nand U1396 (N_1396,In_546,In_390);
xnor U1397 (N_1397,In_137,In_204);
nor U1398 (N_1398,In_190,In_261);
xnor U1399 (N_1399,In_72,In_586);
nand U1400 (N_1400,In_655,In_618);
nand U1401 (N_1401,In_43,In_326);
or U1402 (N_1402,In_614,In_655);
nand U1403 (N_1403,In_604,In_627);
nand U1404 (N_1404,In_585,In_621);
nand U1405 (N_1405,In_327,In_1);
xnor U1406 (N_1406,In_530,In_500);
nor U1407 (N_1407,In_93,In_204);
and U1408 (N_1408,In_348,In_12);
nor U1409 (N_1409,In_677,In_58);
xor U1410 (N_1410,In_22,In_7);
nand U1411 (N_1411,In_102,In_160);
xnor U1412 (N_1412,In_176,In_668);
nand U1413 (N_1413,In_631,In_373);
and U1414 (N_1414,In_658,In_359);
xor U1415 (N_1415,In_627,In_99);
nor U1416 (N_1416,In_639,In_104);
xnor U1417 (N_1417,In_115,In_577);
or U1418 (N_1418,In_516,In_645);
or U1419 (N_1419,In_158,In_234);
or U1420 (N_1420,In_3,In_267);
and U1421 (N_1421,In_308,In_61);
nor U1422 (N_1422,In_325,In_214);
nand U1423 (N_1423,In_113,In_484);
xor U1424 (N_1424,In_245,In_236);
xnor U1425 (N_1425,In_7,In_623);
xnor U1426 (N_1426,In_248,In_429);
nor U1427 (N_1427,In_623,In_685);
nand U1428 (N_1428,In_57,In_52);
and U1429 (N_1429,In_221,In_321);
nor U1430 (N_1430,In_148,In_55);
or U1431 (N_1431,In_420,In_432);
or U1432 (N_1432,In_504,In_329);
xnor U1433 (N_1433,In_572,In_587);
and U1434 (N_1434,In_700,In_62);
or U1435 (N_1435,In_562,In_95);
nand U1436 (N_1436,In_477,In_73);
and U1437 (N_1437,In_74,In_85);
nand U1438 (N_1438,In_553,In_662);
and U1439 (N_1439,In_415,In_322);
nand U1440 (N_1440,In_703,In_383);
or U1441 (N_1441,In_477,In_346);
nand U1442 (N_1442,In_227,In_289);
xnor U1443 (N_1443,In_646,In_606);
xor U1444 (N_1444,In_733,In_230);
nand U1445 (N_1445,In_658,In_289);
nand U1446 (N_1446,In_581,In_19);
nand U1447 (N_1447,In_36,In_99);
and U1448 (N_1448,In_363,In_143);
nand U1449 (N_1449,In_304,In_250);
and U1450 (N_1450,In_278,In_394);
nor U1451 (N_1451,In_469,In_315);
nand U1452 (N_1452,In_6,In_242);
and U1453 (N_1453,In_335,In_440);
nand U1454 (N_1454,In_355,In_443);
nand U1455 (N_1455,In_170,In_223);
xor U1456 (N_1456,In_139,In_394);
and U1457 (N_1457,In_666,In_689);
nor U1458 (N_1458,In_174,In_182);
or U1459 (N_1459,In_235,In_335);
xor U1460 (N_1460,In_598,In_160);
and U1461 (N_1461,In_84,In_393);
nor U1462 (N_1462,In_505,In_708);
nor U1463 (N_1463,In_61,In_273);
and U1464 (N_1464,In_243,In_463);
nand U1465 (N_1465,In_547,In_317);
xnor U1466 (N_1466,In_453,In_686);
nor U1467 (N_1467,In_98,In_310);
nor U1468 (N_1468,In_315,In_337);
or U1469 (N_1469,In_39,In_538);
nand U1470 (N_1470,In_264,In_290);
nor U1471 (N_1471,In_155,In_219);
nand U1472 (N_1472,In_154,In_681);
nand U1473 (N_1473,In_607,In_191);
nor U1474 (N_1474,In_476,In_209);
nand U1475 (N_1475,In_341,In_228);
nand U1476 (N_1476,In_58,In_552);
nand U1477 (N_1477,In_523,In_733);
nand U1478 (N_1478,In_509,In_8);
nor U1479 (N_1479,In_418,In_229);
nor U1480 (N_1480,In_91,In_66);
and U1481 (N_1481,In_269,In_310);
or U1482 (N_1482,In_258,In_250);
and U1483 (N_1483,In_62,In_449);
xor U1484 (N_1484,In_432,In_112);
xnor U1485 (N_1485,In_621,In_255);
xor U1486 (N_1486,In_506,In_559);
nand U1487 (N_1487,In_403,In_308);
nor U1488 (N_1488,In_23,In_553);
nand U1489 (N_1489,In_393,In_578);
nand U1490 (N_1490,In_736,In_214);
nand U1491 (N_1491,In_648,In_472);
xor U1492 (N_1492,In_245,In_442);
and U1493 (N_1493,In_384,In_310);
and U1494 (N_1494,In_612,In_202);
nor U1495 (N_1495,In_624,In_207);
or U1496 (N_1496,In_550,In_358);
nor U1497 (N_1497,In_176,In_675);
xor U1498 (N_1498,In_642,In_285);
or U1499 (N_1499,In_648,In_238);
nand U1500 (N_1500,In_73,In_742);
nor U1501 (N_1501,In_550,In_433);
nor U1502 (N_1502,In_632,In_518);
xor U1503 (N_1503,In_49,In_678);
or U1504 (N_1504,In_226,In_598);
xor U1505 (N_1505,In_324,In_546);
nor U1506 (N_1506,In_300,In_30);
nand U1507 (N_1507,In_549,In_132);
or U1508 (N_1508,In_654,In_244);
and U1509 (N_1509,In_505,In_454);
nand U1510 (N_1510,In_8,In_302);
nand U1511 (N_1511,In_700,In_400);
or U1512 (N_1512,In_642,In_367);
nand U1513 (N_1513,In_169,In_727);
or U1514 (N_1514,In_687,In_618);
nand U1515 (N_1515,In_92,In_70);
nand U1516 (N_1516,In_267,In_138);
or U1517 (N_1517,In_22,In_214);
or U1518 (N_1518,In_339,In_182);
xor U1519 (N_1519,In_181,In_718);
or U1520 (N_1520,In_213,In_412);
or U1521 (N_1521,In_574,In_142);
nor U1522 (N_1522,In_110,In_672);
or U1523 (N_1523,In_262,In_387);
and U1524 (N_1524,In_302,In_337);
xnor U1525 (N_1525,In_631,In_70);
nand U1526 (N_1526,In_142,In_417);
or U1527 (N_1527,In_591,In_76);
xnor U1528 (N_1528,In_709,In_58);
and U1529 (N_1529,In_606,In_654);
or U1530 (N_1530,In_689,In_149);
and U1531 (N_1531,In_621,In_99);
and U1532 (N_1532,In_698,In_432);
nand U1533 (N_1533,In_23,In_309);
nand U1534 (N_1534,In_367,In_484);
or U1535 (N_1535,In_382,In_193);
or U1536 (N_1536,In_439,In_623);
or U1537 (N_1537,In_300,In_621);
or U1538 (N_1538,In_24,In_381);
and U1539 (N_1539,In_627,In_525);
and U1540 (N_1540,In_551,In_567);
or U1541 (N_1541,In_439,In_223);
nand U1542 (N_1542,In_520,In_40);
nand U1543 (N_1543,In_474,In_518);
or U1544 (N_1544,In_188,In_437);
or U1545 (N_1545,In_302,In_282);
nor U1546 (N_1546,In_209,In_455);
or U1547 (N_1547,In_358,In_406);
and U1548 (N_1548,In_605,In_642);
or U1549 (N_1549,In_573,In_1);
nand U1550 (N_1550,In_530,In_465);
nor U1551 (N_1551,In_618,In_207);
and U1552 (N_1552,In_156,In_534);
and U1553 (N_1553,In_211,In_359);
nor U1554 (N_1554,In_632,In_306);
nand U1555 (N_1555,In_198,In_19);
xor U1556 (N_1556,In_238,In_426);
xor U1557 (N_1557,In_626,In_107);
nand U1558 (N_1558,In_573,In_156);
nand U1559 (N_1559,In_576,In_377);
xor U1560 (N_1560,In_71,In_470);
nor U1561 (N_1561,In_400,In_677);
xnor U1562 (N_1562,In_508,In_610);
or U1563 (N_1563,In_545,In_512);
nor U1564 (N_1564,In_579,In_351);
nor U1565 (N_1565,In_449,In_663);
nand U1566 (N_1566,In_265,In_545);
nor U1567 (N_1567,In_364,In_531);
nor U1568 (N_1568,In_555,In_303);
nor U1569 (N_1569,In_740,In_699);
nand U1570 (N_1570,In_317,In_542);
or U1571 (N_1571,In_645,In_224);
nand U1572 (N_1572,In_105,In_729);
xnor U1573 (N_1573,In_271,In_110);
and U1574 (N_1574,In_176,In_11);
and U1575 (N_1575,In_603,In_164);
and U1576 (N_1576,In_82,In_255);
nor U1577 (N_1577,In_401,In_560);
and U1578 (N_1578,In_299,In_321);
or U1579 (N_1579,In_464,In_297);
nor U1580 (N_1580,In_508,In_405);
or U1581 (N_1581,In_80,In_319);
and U1582 (N_1582,In_250,In_321);
nand U1583 (N_1583,In_104,In_37);
and U1584 (N_1584,In_739,In_106);
nor U1585 (N_1585,In_599,In_223);
nand U1586 (N_1586,In_4,In_95);
xnor U1587 (N_1587,In_662,In_670);
and U1588 (N_1588,In_631,In_147);
xnor U1589 (N_1589,In_363,In_719);
or U1590 (N_1590,In_48,In_687);
xnor U1591 (N_1591,In_658,In_100);
nor U1592 (N_1592,In_605,In_487);
and U1593 (N_1593,In_321,In_158);
nand U1594 (N_1594,In_493,In_568);
xnor U1595 (N_1595,In_254,In_257);
nor U1596 (N_1596,In_608,In_132);
and U1597 (N_1597,In_637,In_659);
or U1598 (N_1598,In_54,In_76);
xor U1599 (N_1599,In_524,In_735);
nor U1600 (N_1600,In_413,In_182);
nor U1601 (N_1601,In_544,In_409);
or U1602 (N_1602,In_566,In_98);
and U1603 (N_1603,In_454,In_544);
or U1604 (N_1604,In_1,In_34);
and U1605 (N_1605,In_589,In_726);
or U1606 (N_1606,In_675,In_674);
nand U1607 (N_1607,In_657,In_662);
or U1608 (N_1608,In_207,In_128);
and U1609 (N_1609,In_63,In_496);
or U1610 (N_1610,In_496,In_34);
xnor U1611 (N_1611,In_578,In_517);
nor U1612 (N_1612,In_70,In_120);
and U1613 (N_1613,In_60,In_626);
or U1614 (N_1614,In_96,In_435);
nand U1615 (N_1615,In_595,In_312);
nand U1616 (N_1616,In_667,In_571);
nand U1617 (N_1617,In_4,In_51);
nand U1618 (N_1618,In_265,In_480);
nand U1619 (N_1619,In_501,In_56);
xnor U1620 (N_1620,In_666,In_87);
and U1621 (N_1621,In_246,In_58);
or U1622 (N_1622,In_473,In_744);
and U1623 (N_1623,In_349,In_365);
nor U1624 (N_1624,In_49,In_219);
or U1625 (N_1625,In_47,In_299);
nor U1626 (N_1626,In_685,In_557);
and U1627 (N_1627,In_338,In_534);
xnor U1628 (N_1628,In_83,In_4);
nand U1629 (N_1629,In_414,In_389);
xnor U1630 (N_1630,In_250,In_177);
nand U1631 (N_1631,In_563,In_70);
nor U1632 (N_1632,In_603,In_406);
and U1633 (N_1633,In_398,In_160);
nand U1634 (N_1634,In_372,In_736);
and U1635 (N_1635,In_521,In_632);
and U1636 (N_1636,In_503,In_232);
nand U1637 (N_1637,In_736,In_568);
xnor U1638 (N_1638,In_678,In_3);
nor U1639 (N_1639,In_356,In_368);
and U1640 (N_1640,In_591,In_242);
nand U1641 (N_1641,In_452,In_104);
nor U1642 (N_1642,In_652,In_539);
nand U1643 (N_1643,In_495,In_141);
nand U1644 (N_1644,In_273,In_642);
xnor U1645 (N_1645,In_593,In_559);
nand U1646 (N_1646,In_421,In_579);
and U1647 (N_1647,In_582,In_364);
nand U1648 (N_1648,In_370,In_432);
or U1649 (N_1649,In_606,In_742);
nand U1650 (N_1650,In_376,In_234);
nand U1651 (N_1651,In_151,In_731);
xnor U1652 (N_1652,In_376,In_395);
nor U1653 (N_1653,In_716,In_225);
and U1654 (N_1654,In_215,In_67);
nor U1655 (N_1655,In_417,In_457);
nand U1656 (N_1656,In_587,In_607);
and U1657 (N_1657,In_665,In_421);
or U1658 (N_1658,In_279,In_670);
and U1659 (N_1659,In_151,In_143);
nand U1660 (N_1660,In_593,In_116);
xor U1661 (N_1661,In_175,In_6);
or U1662 (N_1662,In_703,In_713);
nor U1663 (N_1663,In_378,In_294);
nand U1664 (N_1664,In_303,In_413);
nand U1665 (N_1665,In_405,In_514);
xor U1666 (N_1666,In_11,In_319);
and U1667 (N_1667,In_549,In_645);
nor U1668 (N_1668,In_78,In_219);
xnor U1669 (N_1669,In_319,In_239);
nand U1670 (N_1670,In_462,In_32);
nor U1671 (N_1671,In_626,In_419);
xnor U1672 (N_1672,In_636,In_520);
nand U1673 (N_1673,In_448,In_39);
nand U1674 (N_1674,In_603,In_597);
xnor U1675 (N_1675,In_93,In_605);
and U1676 (N_1676,In_672,In_465);
and U1677 (N_1677,In_685,In_454);
nand U1678 (N_1678,In_360,In_71);
nor U1679 (N_1679,In_723,In_371);
or U1680 (N_1680,In_276,In_11);
and U1681 (N_1681,In_147,In_54);
nor U1682 (N_1682,In_492,In_320);
nor U1683 (N_1683,In_719,In_84);
nor U1684 (N_1684,In_344,In_631);
xor U1685 (N_1685,In_146,In_525);
xor U1686 (N_1686,In_672,In_317);
xor U1687 (N_1687,In_699,In_370);
or U1688 (N_1688,In_394,In_546);
nand U1689 (N_1689,In_54,In_198);
nand U1690 (N_1690,In_131,In_402);
and U1691 (N_1691,In_392,In_709);
nand U1692 (N_1692,In_29,In_300);
or U1693 (N_1693,In_738,In_393);
or U1694 (N_1694,In_203,In_163);
xor U1695 (N_1695,In_270,In_449);
nand U1696 (N_1696,In_537,In_133);
nand U1697 (N_1697,In_402,In_520);
nor U1698 (N_1698,In_562,In_130);
and U1699 (N_1699,In_136,In_129);
or U1700 (N_1700,In_741,In_261);
and U1701 (N_1701,In_161,In_604);
and U1702 (N_1702,In_174,In_13);
nor U1703 (N_1703,In_32,In_340);
or U1704 (N_1704,In_325,In_608);
nor U1705 (N_1705,In_417,In_124);
nand U1706 (N_1706,In_36,In_308);
nand U1707 (N_1707,In_162,In_286);
or U1708 (N_1708,In_284,In_383);
nor U1709 (N_1709,In_66,In_101);
nand U1710 (N_1710,In_325,In_65);
or U1711 (N_1711,In_282,In_452);
nand U1712 (N_1712,In_732,In_719);
nor U1713 (N_1713,In_686,In_288);
or U1714 (N_1714,In_495,In_84);
nand U1715 (N_1715,In_433,In_436);
and U1716 (N_1716,In_404,In_380);
or U1717 (N_1717,In_699,In_590);
and U1718 (N_1718,In_323,In_355);
or U1719 (N_1719,In_8,In_20);
nand U1720 (N_1720,In_154,In_13);
xor U1721 (N_1721,In_429,In_42);
nand U1722 (N_1722,In_206,In_22);
nor U1723 (N_1723,In_180,In_541);
nor U1724 (N_1724,In_232,In_79);
nand U1725 (N_1725,In_471,In_534);
and U1726 (N_1726,In_495,In_505);
and U1727 (N_1727,In_58,In_10);
and U1728 (N_1728,In_246,In_727);
and U1729 (N_1729,In_366,In_702);
nor U1730 (N_1730,In_203,In_712);
nand U1731 (N_1731,In_4,In_664);
nand U1732 (N_1732,In_178,In_580);
or U1733 (N_1733,In_163,In_562);
nand U1734 (N_1734,In_382,In_710);
nand U1735 (N_1735,In_187,In_318);
nor U1736 (N_1736,In_297,In_358);
and U1737 (N_1737,In_355,In_541);
nand U1738 (N_1738,In_247,In_52);
and U1739 (N_1739,In_386,In_134);
nand U1740 (N_1740,In_591,In_378);
xnor U1741 (N_1741,In_326,In_282);
and U1742 (N_1742,In_721,In_211);
nor U1743 (N_1743,In_450,In_336);
and U1744 (N_1744,In_588,In_71);
xnor U1745 (N_1745,In_643,In_653);
nor U1746 (N_1746,In_153,In_709);
nand U1747 (N_1747,In_589,In_317);
nand U1748 (N_1748,In_435,In_676);
or U1749 (N_1749,In_276,In_697);
nand U1750 (N_1750,In_510,In_310);
and U1751 (N_1751,In_589,In_701);
nand U1752 (N_1752,In_287,In_747);
nand U1753 (N_1753,In_69,In_150);
nand U1754 (N_1754,In_334,In_297);
xor U1755 (N_1755,In_571,In_330);
nor U1756 (N_1756,In_167,In_501);
and U1757 (N_1757,In_214,In_365);
xor U1758 (N_1758,In_116,In_517);
or U1759 (N_1759,In_307,In_129);
or U1760 (N_1760,In_545,In_344);
or U1761 (N_1761,In_439,In_611);
and U1762 (N_1762,In_621,In_557);
xnor U1763 (N_1763,In_35,In_210);
nand U1764 (N_1764,In_658,In_284);
and U1765 (N_1765,In_345,In_553);
nor U1766 (N_1766,In_503,In_322);
and U1767 (N_1767,In_360,In_32);
nor U1768 (N_1768,In_222,In_500);
nand U1769 (N_1769,In_368,In_640);
xnor U1770 (N_1770,In_341,In_639);
nor U1771 (N_1771,In_97,In_217);
and U1772 (N_1772,In_693,In_146);
nor U1773 (N_1773,In_454,In_365);
nand U1774 (N_1774,In_499,In_322);
nor U1775 (N_1775,In_256,In_469);
nor U1776 (N_1776,In_562,In_693);
nand U1777 (N_1777,In_99,In_528);
and U1778 (N_1778,In_643,In_516);
and U1779 (N_1779,In_118,In_479);
xor U1780 (N_1780,In_192,In_395);
and U1781 (N_1781,In_158,In_451);
nand U1782 (N_1782,In_659,In_324);
or U1783 (N_1783,In_617,In_433);
nor U1784 (N_1784,In_224,In_494);
and U1785 (N_1785,In_372,In_465);
and U1786 (N_1786,In_361,In_444);
nand U1787 (N_1787,In_31,In_480);
xnor U1788 (N_1788,In_13,In_162);
and U1789 (N_1789,In_17,In_175);
or U1790 (N_1790,In_634,In_710);
xnor U1791 (N_1791,In_576,In_231);
nor U1792 (N_1792,In_641,In_600);
xor U1793 (N_1793,In_603,In_1);
xnor U1794 (N_1794,In_712,In_522);
and U1795 (N_1795,In_702,In_349);
and U1796 (N_1796,In_256,In_298);
nor U1797 (N_1797,In_353,In_75);
nor U1798 (N_1798,In_149,In_184);
and U1799 (N_1799,In_242,In_669);
xor U1800 (N_1800,In_672,In_702);
xor U1801 (N_1801,In_733,In_706);
xnor U1802 (N_1802,In_56,In_81);
and U1803 (N_1803,In_713,In_388);
and U1804 (N_1804,In_41,In_136);
nand U1805 (N_1805,In_328,In_424);
nand U1806 (N_1806,In_572,In_132);
or U1807 (N_1807,In_124,In_215);
and U1808 (N_1808,In_323,In_516);
xnor U1809 (N_1809,In_416,In_498);
and U1810 (N_1810,In_557,In_541);
or U1811 (N_1811,In_631,In_689);
and U1812 (N_1812,In_245,In_684);
and U1813 (N_1813,In_69,In_250);
nor U1814 (N_1814,In_425,In_120);
nand U1815 (N_1815,In_225,In_340);
or U1816 (N_1816,In_190,In_282);
xnor U1817 (N_1817,In_0,In_586);
nand U1818 (N_1818,In_359,In_45);
or U1819 (N_1819,In_76,In_58);
nor U1820 (N_1820,In_349,In_111);
or U1821 (N_1821,In_104,In_33);
or U1822 (N_1822,In_485,In_142);
or U1823 (N_1823,In_736,In_472);
nor U1824 (N_1824,In_386,In_348);
or U1825 (N_1825,In_182,In_386);
nand U1826 (N_1826,In_256,In_231);
xor U1827 (N_1827,In_68,In_351);
nand U1828 (N_1828,In_502,In_102);
nand U1829 (N_1829,In_191,In_479);
xor U1830 (N_1830,In_3,In_224);
or U1831 (N_1831,In_343,In_199);
nor U1832 (N_1832,In_628,In_216);
and U1833 (N_1833,In_66,In_591);
nor U1834 (N_1834,In_76,In_350);
nor U1835 (N_1835,In_243,In_522);
nor U1836 (N_1836,In_191,In_563);
nand U1837 (N_1837,In_653,In_122);
or U1838 (N_1838,In_105,In_289);
or U1839 (N_1839,In_454,In_478);
and U1840 (N_1840,In_404,In_56);
xor U1841 (N_1841,In_355,In_207);
xnor U1842 (N_1842,In_389,In_472);
nand U1843 (N_1843,In_419,In_291);
nor U1844 (N_1844,In_410,In_617);
or U1845 (N_1845,In_179,In_416);
nand U1846 (N_1846,In_741,In_64);
nor U1847 (N_1847,In_553,In_371);
nand U1848 (N_1848,In_660,In_236);
nor U1849 (N_1849,In_718,In_376);
or U1850 (N_1850,In_300,In_133);
nand U1851 (N_1851,In_201,In_43);
and U1852 (N_1852,In_673,In_455);
nand U1853 (N_1853,In_453,In_564);
nand U1854 (N_1854,In_526,In_499);
nand U1855 (N_1855,In_215,In_643);
and U1856 (N_1856,In_100,In_395);
or U1857 (N_1857,In_53,In_538);
and U1858 (N_1858,In_162,In_1);
and U1859 (N_1859,In_23,In_451);
and U1860 (N_1860,In_50,In_554);
nor U1861 (N_1861,In_257,In_165);
nand U1862 (N_1862,In_51,In_159);
or U1863 (N_1863,In_2,In_586);
and U1864 (N_1864,In_720,In_174);
and U1865 (N_1865,In_430,In_721);
or U1866 (N_1866,In_145,In_16);
nand U1867 (N_1867,In_94,In_533);
xor U1868 (N_1868,In_573,In_727);
nor U1869 (N_1869,In_105,In_281);
nand U1870 (N_1870,In_412,In_1);
nand U1871 (N_1871,In_427,In_87);
nor U1872 (N_1872,In_698,In_596);
nand U1873 (N_1873,In_351,In_664);
nor U1874 (N_1874,In_499,In_91);
xor U1875 (N_1875,In_13,In_666);
nor U1876 (N_1876,In_287,In_276);
xnor U1877 (N_1877,In_530,In_273);
xnor U1878 (N_1878,In_110,In_405);
nand U1879 (N_1879,In_591,In_351);
xnor U1880 (N_1880,In_344,In_239);
and U1881 (N_1881,In_475,In_412);
xnor U1882 (N_1882,In_233,In_314);
nand U1883 (N_1883,In_303,In_398);
nand U1884 (N_1884,In_42,In_249);
xor U1885 (N_1885,In_281,In_456);
nand U1886 (N_1886,In_173,In_625);
or U1887 (N_1887,In_450,In_228);
xnor U1888 (N_1888,In_303,In_94);
or U1889 (N_1889,In_125,In_186);
xor U1890 (N_1890,In_188,In_522);
and U1891 (N_1891,In_271,In_148);
or U1892 (N_1892,In_410,In_279);
xor U1893 (N_1893,In_445,In_653);
xnor U1894 (N_1894,In_624,In_619);
nor U1895 (N_1895,In_96,In_521);
and U1896 (N_1896,In_36,In_601);
xor U1897 (N_1897,In_515,In_529);
and U1898 (N_1898,In_244,In_167);
nor U1899 (N_1899,In_632,In_547);
nor U1900 (N_1900,In_504,In_324);
and U1901 (N_1901,In_690,In_481);
or U1902 (N_1902,In_77,In_361);
nand U1903 (N_1903,In_32,In_27);
xnor U1904 (N_1904,In_311,In_11);
nand U1905 (N_1905,In_267,In_219);
xor U1906 (N_1906,In_672,In_628);
nor U1907 (N_1907,In_749,In_640);
nor U1908 (N_1908,In_298,In_559);
and U1909 (N_1909,In_386,In_699);
nand U1910 (N_1910,In_737,In_565);
xor U1911 (N_1911,In_62,In_490);
or U1912 (N_1912,In_290,In_232);
nor U1913 (N_1913,In_745,In_444);
or U1914 (N_1914,In_623,In_524);
xnor U1915 (N_1915,In_468,In_582);
and U1916 (N_1916,In_337,In_533);
or U1917 (N_1917,In_80,In_37);
nor U1918 (N_1918,In_353,In_32);
nand U1919 (N_1919,In_132,In_428);
nor U1920 (N_1920,In_657,In_284);
nor U1921 (N_1921,In_544,In_175);
xor U1922 (N_1922,In_711,In_66);
and U1923 (N_1923,In_426,In_135);
nor U1924 (N_1924,In_567,In_444);
xnor U1925 (N_1925,In_543,In_576);
nor U1926 (N_1926,In_467,In_479);
nor U1927 (N_1927,In_311,In_275);
and U1928 (N_1928,In_252,In_403);
xor U1929 (N_1929,In_617,In_610);
or U1930 (N_1930,In_380,In_394);
nand U1931 (N_1931,In_634,In_107);
nor U1932 (N_1932,In_209,In_102);
and U1933 (N_1933,In_5,In_312);
nand U1934 (N_1934,In_151,In_52);
or U1935 (N_1935,In_47,In_522);
and U1936 (N_1936,In_537,In_662);
xor U1937 (N_1937,In_470,In_543);
nor U1938 (N_1938,In_591,In_502);
and U1939 (N_1939,In_692,In_129);
xor U1940 (N_1940,In_467,In_393);
or U1941 (N_1941,In_97,In_313);
and U1942 (N_1942,In_248,In_732);
nor U1943 (N_1943,In_324,In_560);
nand U1944 (N_1944,In_193,In_117);
or U1945 (N_1945,In_571,In_684);
xor U1946 (N_1946,In_428,In_535);
nor U1947 (N_1947,In_222,In_509);
or U1948 (N_1948,In_617,In_119);
nor U1949 (N_1949,In_459,In_442);
xnor U1950 (N_1950,In_286,In_218);
xor U1951 (N_1951,In_473,In_195);
or U1952 (N_1952,In_100,In_447);
or U1953 (N_1953,In_696,In_260);
or U1954 (N_1954,In_744,In_629);
xor U1955 (N_1955,In_268,In_136);
nor U1956 (N_1956,In_688,In_518);
nand U1957 (N_1957,In_98,In_170);
and U1958 (N_1958,In_578,In_504);
nand U1959 (N_1959,In_157,In_654);
xnor U1960 (N_1960,In_162,In_615);
or U1961 (N_1961,In_555,In_166);
nand U1962 (N_1962,In_439,In_687);
xnor U1963 (N_1963,In_193,In_166);
xor U1964 (N_1964,In_133,In_603);
xnor U1965 (N_1965,In_604,In_489);
or U1966 (N_1966,In_235,In_122);
and U1967 (N_1967,In_41,In_619);
nor U1968 (N_1968,In_648,In_464);
or U1969 (N_1969,In_279,In_331);
xnor U1970 (N_1970,In_516,In_354);
or U1971 (N_1971,In_55,In_58);
nand U1972 (N_1972,In_172,In_139);
and U1973 (N_1973,In_631,In_552);
nand U1974 (N_1974,In_475,In_572);
xor U1975 (N_1975,In_98,In_525);
nor U1976 (N_1976,In_455,In_64);
nor U1977 (N_1977,In_582,In_463);
xor U1978 (N_1978,In_61,In_42);
nor U1979 (N_1979,In_463,In_321);
and U1980 (N_1980,In_312,In_250);
nand U1981 (N_1981,In_383,In_489);
nor U1982 (N_1982,In_466,In_91);
or U1983 (N_1983,In_499,In_645);
xnor U1984 (N_1984,In_27,In_242);
or U1985 (N_1985,In_638,In_730);
nor U1986 (N_1986,In_22,In_739);
xor U1987 (N_1987,In_713,In_575);
and U1988 (N_1988,In_665,In_25);
nand U1989 (N_1989,In_260,In_402);
and U1990 (N_1990,In_208,In_462);
xnor U1991 (N_1991,In_514,In_526);
xor U1992 (N_1992,In_590,In_166);
or U1993 (N_1993,In_387,In_516);
nand U1994 (N_1994,In_502,In_1);
or U1995 (N_1995,In_385,In_408);
xnor U1996 (N_1996,In_314,In_720);
and U1997 (N_1997,In_133,In_109);
nand U1998 (N_1998,In_175,In_237);
nand U1999 (N_1999,In_428,In_404);
nor U2000 (N_2000,In_659,In_371);
and U2001 (N_2001,In_280,In_458);
xor U2002 (N_2002,In_445,In_384);
nor U2003 (N_2003,In_205,In_440);
or U2004 (N_2004,In_425,In_145);
and U2005 (N_2005,In_482,In_597);
xnor U2006 (N_2006,In_304,In_176);
xor U2007 (N_2007,In_18,In_149);
xnor U2008 (N_2008,In_258,In_103);
nor U2009 (N_2009,In_336,In_413);
or U2010 (N_2010,In_683,In_743);
or U2011 (N_2011,In_382,In_133);
nand U2012 (N_2012,In_520,In_597);
nand U2013 (N_2013,In_338,In_60);
and U2014 (N_2014,In_1,In_713);
xnor U2015 (N_2015,In_299,In_481);
and U2016 (N_2016,In_81,In_550);
xor U2017 (N_2017,In_692,In_79);
and U2018 (N_2018,In_516,In_119);
and U2019 (N_2019,In_120,In_49);
nor U2020 (N_2020,In_136,In_485);
nand U2021 (N_2021,In_409,In_211);
nand U2022 (N_2022,In_94,In_596);
xor U2023 (N_2023,In_516,In_183);
nor U2024 (N_2024,In_747,In_688);
nor U2025 (N_2025,In_522,In_449);
and U2026 (N_2026,In_212,In_11);
or U2027 (N_2027,In_702,In_740);
nor U2028 (N_2028,In_347,In_454);
and U2029 (N_2029,In_427,In_613);
and U2030 (N_2030,In_15,In_529);
and U2031 (N_2031,In_516,In_139);
or U2032 (N_2032,In_702,In_394);
xor U2033 (N_2033,In_429,In_297);
nor U2034 (N_2034,In_635,In_731);
nor U2035 (N_2035,In_246,In_300);
nand U2036 (N_2036,In_416,In_214);
xnor U2037 (N_2037,In_428,In_261);
nand U2038 (N_2038,In_423,In_446);
xor U2039 (N_2039,In_687,In_477);
and U2040 (N_2040,In_89,In_543);
nand U2041 (N_2041,In_325,In_684);
xor U2042 (N_2042,In_189,In_108);
or U2043 (N_2043,In_263,In_681);
and U2044 (N_2044,In_436,In_162);
xor U2045 (N_2045,In_249,In_207);
and U2046 (N_2046,In_316,In_32);
nand U2047 (N_2047,In_76,In_534);
nor U2048 (N_2048,In_79,In_465);
xor U2049 (N_2049,In_217,In_354);
nand U2050 (N_2050,In_736,In_434);
xor U2051 (N_2051,In_566,In_111);
or U2052 (N_2052,In_237,In_681);
xor U2053 (N_2053,In_132,In_249);
nor U2054 (N_2054,In_494,In_367);
and U2055 (N_2055,In_504,In_63);
nand U2056 (N_2056,In_290,In_366);
nand U2057 (N_2057,In_346,In_508);
and U2058 (N_2058,In_259,In_413);
or U2059 (N_2059,In_623,In_460);
or U2060 (N_2060,In_437,In_151);
nand U2061 (N_2061,In_65,In_124);
or U2062 (N_2062,In_486,In_208);
and U2063 (N_2063,In_148,In_299);
and U2064 (N_2064,In_463,In_67);
or U2065 (N_2065,In_434,In_629);
nor U2066 (N_2066,In_34,In_626);
nand U2067 (N_2067,In_419,In_607);
nor U2068 (N_2068,In_87,In_655);
and U2069 (N_2069,In_507,In_85);
or U2070 (N_2070,In_521,In_626);
nand U2071 (N_2071,In_331,In_470);
and U2072 (N_2072,In_728,In_525);
nor U2073 (N_2073,In_705,In_308);
nand U2074 (N_2074,In_144,In_143);
xnor U2075 (N_2075,In_594,In_547);
or U2076 (N_2076,In_447,In_483);
and U2077 (N_2077,In_611,In_449);
xnor U2078 (N_2078,In_117,In_355);
nand U2079 (N_2079,In_662,In_646);
nand U2080 (N_2080,In_403,In_353);
xor U2081 (N_2081,In_80,In_97);
nor U2082 (N_2082,In_421,In_666);
nand U2083 (N_2083,In_472,In_72);
nor U2084 (N_2084,In_727,In_198);
nor U2085 (N_2085,In_90,In_424);
nand U2086 (N_2086,In_436,In_92);
or U2087 (N_2087,In_532,In_307);
nor U2088 (N_2088,In_666,In_729);
nand U2089 (N_2089,In_542,In_214);
nand U2090 (N_2090,In_14,In_196);
nand U2091 (N_2091,In_435,In_665);
xor U2092 (N_2092,In_742,In_292);
nand U2093 (N_2093,In_107,In_621);
and U2094 (N_2094,In_408,In_644);
or U2095 (N_2095,In_45,In_478);
nor U2096 (N_2096,In_450,In_329);
nor U2097 (N_2097,In_202,In_365);
nor U2098 (N_2098,In_107,In_196);
or U2099 (N_2099,In_150,In_168);
nand U2100 (N_2100,In_180,In_516);
xnor U2101 (N_2101,In_615,In_261);
or U2102 (N_2102,In_489,In_20);
and U2103 (N_2103,In_680,In_258);
nor U2104 (N_2104,In_183,In_81);
or U2105 (N_2105,In_293,In_255);
nand U2106 (N_2106,In_22,In_417);
nand U2107 (N_2107,In_197,In_279);
nand U2108 (N_2108,In_332,In_80);
nand U2109 (N_2109,In_331,In_712);
or U2110 (N_2110,In_337,In_17);
or U2111 (N_2111,In_127,In_256);
or U2112 (N_2112,In_671,In_574);
nor U2113 (N_2113,In_89,In_399);
nand U2114 (N_2114,In_456,In_116);
nand U2115 (N_2115,In_320,In_735);
nand U2116 (N_2116,In_575,In_3);
and U2117 (N_2117,In_146,In_406);
nor U2118 (N_2118,In_211,In_352);
and U2119 (N_2119,In_18,In_454);
and U2120 (N_2120,In_725,In_254);
nor U2121 (N_2121,In_306,In_185);
nor U2122 (N_2122,In_626,In_648);
nor U2123 (N_2123,In_657,In_122);
nor U2124 (N_2124,In_103,In_586);
xnor U2125 (N_2125,In_456,In_416);
and U2126 (N_2126,In_326,In_105);
and U2127 (N_2127,In_375,In_463);
nor U2128 (N_2128,In_54,In_613);
or U2129 (N_2129,In_335,In_433);
nand U2130 (N_2130,In_140,In_658);
xor U2131 (N_2131,In_680,In_372);
nor U2132 (N_2132,In_736,In_299);
nand U2133 (N_2133,In_345,In_567);
nand U2134 (N_2134,In_406,In_142);
and U2135 (N_2135,In_377,In_671);
nor U2136 (N_2136,In_207,In_165);
nand U2137 (N_2137,In_356,In_454);
or U2138 (N_2138,In_576,In_331);
nor U2139 (N_2139,In_22,In_337);
nor U2140 (N_2140,In_269,In_82);
xor U2141 (N_2141,In_444,In_119);
xor U2142 (N_2142,In_548,In_142);
and U2143 (N_2143,In_617,In_471);
nand U2144 (N_2144,In_440,In_736);
nand U2145 (N_2145,In_611,In_448);
nand U2146 (N_2146,In_66,In_520);
xor U2147 (N_2147,In_685,In_715);
nand U2148 (N_2148,In_388,In_524);
or U2149 (N_2149,In_450,In_680);
or U2150 (N_2150,In_263,In_675);
nand U2151 (N_2151,In_172,In_79);
nor U2152 (N_2152,In_323,In_336);
or U2153 (N_2153,In_704,In_17);
xnor U2154 (N_2154,In_516,In_76);
nand U2155 (N_2155,In_397,In_606);
or U2156 (N_2156,In_200,In_254);
and U2157 (N_2157,In_460,In_521);
or U2158 (N_2158,In_721,In_316);
xor U2159 (N_2159,In_548,In_12);
nor U2160 (N_2160,In_456,In_144);
and U2161 (N_2161,In_108,In_66);
nor U2162 (N_2162,In_118,In_268);
xnor U2163 (N_2163,In_240,In_439);
and U2164 (N_2164,In_103,In_368);
nand U2165 (N_2165,In_485,In_682);
xor U2166 (N_2166,In_377,In_644);
xnor U2167 (N_2167,In_488,In_7);
nand U2168 (N_2168,In_617,In_120);
or U2169 (N_2169,In_706,In_325);
nor U2170 (N_2170,In_54,In_333);
nand U2171 (N_2171,In_273,In_657);
and U2172 (N_2172,In_243,In_344);
xnor U2173 (N_2173,In_669,In_39);
xnor U2174 (N_2174,In_556,In_446);
nand U2175 (N_2175,In_38,In_515);
nand U2176 (N_2176,In_161,In_701);
or U2177 (N_2177,In_338,In_68);
nand U2178 (N_2178,In_491,In_599);
xnor U2179 (N_2179,In_75,In_518);
or U2180 (N_2180,In_203,In_312);
nand U2181 (N_2181,In_118,In_636);
xnor U2182 (N_2182,In_482,In_109);
xor U2183 (N_2183,In_9,In_584);
nor U2184 (N_2184,In_677,In_542);
or U2185 (N_2185,In_391,In_638);
and U2186 (N_2186,In_521,In_746);
xor U2187 (N_2187,In_556,In_697);
xnor U2188 (N_2188,In_142,In_14);
nand U2189 (N_2189,In_477,In_589);
nand U2190 (N_2190,In_6,In_577);
nor U2191 (N_2191,In_692,In_21);
and U2192 (N_2192,In_324,In_292);
and U2193 (N_2193,In_463,In_279);
xnor U2194 (N_2194,In_156,In_660);
xnor U2195 (N_2195,In_651,In_681);
or U2196 (N_2196,In_398,In_657);
xnor U2197 (N_2197,In_153,In_529);
or U2198 (N_2198,In_217,In_629);
xnor U2199 (N_2199,In_476,In_146);
nor U2200 (N_2200,In_61,In_69);
and U2201 (N_2201,In_531,In_552);
and U2202 (N_2202,In_648,In_293);
nor U2203 (N_2203,In_85,In_722);
nor U2204 (N_2204,In_215,In_437);
nand U2205 (N_2205,In_347,In_715);
or U2206 (N_2206,In_270,In_87);
or U2207 (N_2207,In_482,In_728);
nand U2208 (N_2208,In_79,In_58);
nor U2209 (N_2209,In_197,In_126);
nor U2210 (N_2210,In_323,In_524);
and U2211 (N_2211,In_638,In_49);
nand U2212 (N_2212,In_652,In_490);
nor U2213 (N_2213,In_613,In_397);
nor U2214 (N_2214,In_501,In_102);
xnor U2215 (N_2215,In_521,In_455);
nor U2216 (N_2216,In_687,In_567);
and U2217 (N_2217,In_387,In_740);
and U2218 (N_2218,In_465,In_107);
nand U2219 (N_2219,In_334,In_56);
and U2220 (N_2220,In_400,In_649);
nor U2221 (N_2221,In_21,In_421);
nor U2222 (N_2222,In_268,In_602);
nor U2223 (N_2223,In_533,In_432);
or U2224 (N_2224,In_361,In_666);
nor U2225 (N_2225,In_425,In_684);
xor U2226 (N_2226,In_440,In_69);
and U2227 (N_2227,In_168,In_630);
nand U2228 (N_2228,In_277,In_479);
nor U2229 (N_2229,In_591,In_300);
or U2230 (N_2230,In_666,In_390);
or U2231 (N_2231,In_716,In_719);
or U2232 (N_2232,In_394,In_146);
xnor U2233 (N_2233,In_509,In_470);
xor U2234 (N_2234,In_672,In_261);
xor U2235 (N_2235,In_214,In_718);
or U2236 (N_2236,In_313,In_259);
xnor U2237 (N_2237,In_125,In_44);
nor U2238 (N_2238,In_306,In_456);
nand U2239 (N_2239,In_650,In_88);
nor U2240 (N_2240,In_111,In_631);
nor U2241 (N_2241,In_437,In_748);
and U2242 (N_2242,In_709,In_537);
or U2243 (N_2243,In_479,In_608);
nand U2244 (N_2244,In_724,In_309);
xnor U2245 (N_2245,In_362,In_68);
and U2246 (N_2246,In_556,In_28);
nor U2247 (N_2247,In_527,In_188);
xor U2248 (N_2248,In_554,In_229);
or U2249 (N_2249,In_218,In_247);
or U2250 (N_2250,In_455,In_620);
or U2251 (N_2251,In_170,In_532);
nor U2252 (N_2252,In_211,In_434);
and U2253 (N_2253,In_245,In_173);
xor U2254 (N_2254,In_137,In_645);
nand U2255 (N_2255,In_546,In_190);
nand U2256 (N_2256,In_599,In_706);
xnor U2257 (N_2257,In_328,In_511);
or U2258 (N_2258,In_372,In_8);
or U2259 (N_2259,In_31,In_217);
or U2260 (N_2260,In_352,In_331);
and U2261 (N_2261,In_10,In_440);
or U2262 (N_2262,In_489,In_347);
nand U2263 (N_2263,In_693,In_706);
and U2264 (N_2264,In_241,In_733);
nand U2265 (N_2265,In_336,In_376);
xnor U2266 (N_2266,In_11,In_201);
and U2267 (N_2267,In_16,In_370);
or U2268 (N_2268,In_723,In_253);
xor U2269 (N_2269,In_330,In_669);
nand U2270 (N_2270,In_619,In_589);
or U2271 (N_2271,In_429,In_649);
and U2272 (N_2272,In_554,In_585);
or U2273 (N_2273,In_657,In_700);
or U2274 (N_2274,In_733,In_97);
nor U2275 (N_2275,In_46,In_683);
nand U2276 (N_2276,In_740,In_652);
and U2277 (N_2277,In_712,In_206);
and U2278 (N_2278,In_76,In_8);
nor U2279 (N_2279,In_483,In_745);
xnor U2280 (N_2280,In_2,In_725);
nand U2281 (N_2281,In_359,In_527);
and U2282 (N_2282,In_562,In_594);
or U2283 (N_2283,In_674,In_538);
xnor U2284 (N_2284,In_287,In_555);
xnor U2285 (N_2285,In_610,In_262);
and U2286 (N_2286,In_422,In_706);
xnor U2287 (N_2287,In_200,In_179);
xnor U2288 (N_2288,In_479,In_47);
or U2289 (N_2289,In_158,In_427);
nand U2290 (N_2290,In_307,In_325);
nand U2291 (N_2291,In_687,In_438);
and U2292 (N_2292,In_444,In_743);
and U2293 (N_2293,In_595,In_435);
and U2294 (N_2294,In_558,In_324);
or U2295 (N_2295,In_746,In_268);
or U2296 (N_2296,In_285,In_644);
nor U2297 (N_2297,In_468,In_26);
and U2298 (N_2298,In_21,In_174);
xor U2299 (N_2299,In_437,In_99);
nand U2300 (N_2300,In_351,In_648);
nor U2301 (N_2301,In_607,In_128);
nand U2302 (N_2302,In_493,In_572);
or U2303 (N_2303,In_554,In_483);
or U2304 (N_2304,In_530,In_710);
nor U2305 (N_2305,In_34,In_197);
and U2306 (N_2306,In_45,In_401);
nand U2307 (N_2307,In_240,In_480);
nand U2308 (N_2308,In_23,In_80);
xnor U2309 (N_2309,In_568,In_588);
or U2310 (N_2310,In_621,In_60);
nor U2311 (N_2311,In_331,In_412);
or U2312 (N_2312,In_148,In_116);
xor U2313 (N_2313,In_366,In_697);
nand U2314 (N_2314,In_360,In_438);
xor U2315 (N_2315,In_228,In_175);
nand U2316 (N_2316,In_414,In_233);
and U2317 (N_2317,In_580,In_535);
nand U2318 (N_2318,In_530,In_691);
or U2319 (N_2319,In_648,In_230);
or U2320 (N_2320,In_132,In_462);
and U2321 (N_2321,In_696,In_213);
and U2322 (N_2322,In_579,In_666);
xnor U2323 (N_2323,In_479,In_200);
or U2324 (N_2324,In_496,In_579);
nor U2325 (N_2325,In_122,In_210);
and U2326 (N_2326,In_577,In_670);
xor U2327 (N_2327,In_340,In_559);
xnor U2328 (N_2328,In_421,In_457);
and U2329 (N_2329,In_285,In_534);
xnor U2330 (N_2330,In_33,In_562);
and U2331 (N_2331,In_474,In_278);
or U2332 (N_2332,In_534,In_366);
nor U2333 (N_2333,In_40,In_664);
xor U2334 (N_2334,In_601,In_646);
or U2335 (N_2335,In_359,In_726);
nor U2336 (N_2336,In_553,In_62);
nand U2337 (N_2337,In_371,In_406);
nand U2338 (N_2338,In_470,In_44);
and U2339 (N_2339,In_310,In_456);
nor U2340 (N_2340,In_321,In_545);
nor U2341 (N_2341,In_337,In_691);
xor U2342 (N_2342,In_146,In_679);
xnor U2343 (N_2343,In_156,In_391);
nor U2344 (N_2344,In_569,In_688);
or U2345 (N_2345,In_455,In_180);
xnor U2346 (N_2346,In_416,In_601);
nand U2347 (N_2347,In_256,In_522);
nand U2348 (N_2348,In_543,In_328);
nand U2349 (N_2349,In_437,In_345);
nor U2350 (N_2350,In_80,In_162);
xor U2351 (N_2351,In_112,In_550);
nor U2352 (N_2352,In_427,In_572);
nand U2353 (N_2353,In_307,In_663);
xor U2354 (N_2354,In_218,In_403);
nor U2355 (N_2355,In_616,In_491);
nor U2356 (N_2356,In_107,In_692);
and U2357 (N_2357,In_84,In_630);
and U2358 (N_2358,In_0,In_668);
nor U2359 (N_2359,In_689,In_725);
nor U2360 (N_2360,In_161,In_191);
and U2361 (N_2361,In_21,In_407);
xnor U2362 (N_2362,In_367,In_627);
nor U2363 (N_2363,In_193,In_326);
and U2364 (N_2364,In_332,In_448);
or U2365 (N_2365,In_464,In_274);
xor U2366 (N_2366,In_473,In_397);
xor U2367 (N_2367,In_279,In_592);
nor U2368 (N_2368,In_495,In_145);
or U2369 (N_2369,In_393,In_310);
and U2370 (N_2370,In_328,In_274);
and U2371 (N_2371,In_163,In_313);
nand U2372 (N_2372,In_253,In_329);
or U2373 (N_2373,In_139,In_304);
or U2374 (N_2374,In_151,In_69);
nand U2375 (N_2375,In_107,In_666);
xnor U2376 (N_2376,In_666,In_97);
or U2377 (N_2377,In_41,In_643);
xnor U2378 (N_2378,In_22,In_336);
nor U2379 (N_2379,In_652,In_297);
xnor U2380 (N_2380,In_587,In_179);
or U2381 (N_2381,In_526,In_736);
xor U2382 (N_2382,In_265,In_572);
nand U2383 (N_2383,In_515,In_112);
and U2384 (N_2384,In_361,In_513);
and U2385 (N_2385,In_551,In_132);
nor U2386 (N_2386,In_549,In_210);
nand U2387 (N_2387,In_198,In_389);
nor U2388 (N_2388,In_314,In_516);
and U2389 (N_2389,In_24,In_9);
nand U2390 (N_2390,In_740,In_475);
and U2391 (N_2391,In_401,In_320);
nand U2392 (N_2392,In_699,In_569);
xnor U2393 (N_2393,In_662,In_331);
and U2394 (N_2394,In_590,In_713);
xnor U2395 (N_2395,In_581,In_113);
and U2396 (N_2396,In_551,In_673);
nor U2397 (N_2397,In_683,In_517);
and U2398 (N_2398,In_733,In_157);
nor U2399 (N_2399,In_16,In_571);
and U2400 (N_2400,In_731,In_616);
and U2401 (N_2401,In_189,In_271);
and U2402 (N_2402,In_124,In_281);
xnor U2403 (N_2403,In_25,In_190);
and U2404 (N_2404,In_353,In_592);
nor U2405 (N_2405,In_520,In_582);
and U2406 (N_2406,In_45,In_152);
and U2407 (N_2407,In_2,In_335);
nor U2408 (N_2408,In_105,In_506);
xnor U2409 (N_2409,In_731,In_602);
nor U2410 (N_2410,In_725,In_102);
xnor U2411 (N_2411,In_288,In_589);
nor U2412 (N_2412,In_202,In_589);
nand U2413 (N_2413,In_729,In_45);
nand U2414 (N_2414,In_36,In_466);
nor U2415 (N_2415,In_240,In_306);
nand U2416 (N_2416,In_489,In_680);
nand U2417 (N_2417,In_82,In_654);
or U2418 (N_2418,In_73,In_378);
nand U2419 (N_2419,In_447,In_613);
nand U2420 (N_2420,In_575,In_226);
nand U2421 (N_2421,In_35,In_616);
or U2422 (N_2422,In_415,In_695);
xor U2423 (N_2423,In_545,In_437);
or U2424 (N_2424,In_57,In_179);
xnor U2425 (N_2425,In_269,In_329);
xor U2426 (N_2426,In_509,In_432);
xor U2427 (N_2427,In_289,In_746);
nand U2428 (N_2428,In_500,In_357);
nor U2429 (N_2429,In_180,In_715);
nor U2430 (N_2430,In_310,In_698);
xor U2431 (N_2431,In_479,In_601);
and U2432 (N_2432,In_607,In_578);
xnor U2433 (N_2433,In_559,In_662);
or U2434 (N_2434,In_654,In_255);
xnor U2435 (N_2435,In_243,In_574);
xor U2436 (N_2436,In_594,In_76);
or U2437 (N_2437,In_211,In_213);
nand U2438 (N_2438,In_600,In_451);
xnor U2439 (N_2439,In_273,In_643);
or U2440 (N_2440,In_482,In_548);
nand U2441 (N_2441,In_577,In_12);
nor U2442 (N_2442,In_338,In_229);
nand U2443 (N_2443,In_99,In_381);
nand U2444 (N_2444,In_648,In_131);
nor U2445 (N_2445,In_307,In_40);
nor U2446 (N_2446,In_238,In_175);
nor U2447 (N_2447,In_388,In_294);
nand U2448 (N_2448,In_389,In_311);
nand U2449 (N_2449,In_324,In_697);
or U2450 (N_2450,In_398,In_87);
or U2451 (N_2451,In_349,In_357);
or U2452 (N_2452,In_497,In_436);
or U2453 (N_2453,In_696,In_560);
nor U2454 (N_2454,In_483,In_286);
nor U2455 (N_2455,In_297,In_674);
or U2456 (N_2456,In_588,In_195);
nor U2457 (N_2457,In_543,In_670);
nand U2458 (N_2458,In_286,In_174);
xnor U2459 (N_2459,In_181,In_586);
and U2460 (N_2460,In_656,In_602);
xnor U2461 (N_2461,In_123,In_747);
xor U2462 (N_2462,In_384,In_710);
or U2463 (N_2463,In_210,In_51);
nand U2464 (N_2464,In_371,In_435);
or U2465 (N_2465,In_717,In_553);
nor U2466 (N_2466,In_474,In_30);
nand U2467 (N_2467,In_227,In_301);
or U2468 (N_2468,In_572,In_328);
nand U2469 (N_2469,In_377,In_592);
or U2470 (N_2470,In_444,In_283);
nor U2471 (N_2471,In_48,In_716);
xor U2472 (N_2472,In_435,In_249);
xnor U2473 (N_2473,In_352,In_30);
nor U2474 (N_2474,In_400,In_56);
and U2475 (N_2475,In_45,In_264);
or U2476 (N_2476,In_11,In_532);
xnor U2477 (N_2477,In_261,In_328);
xor U2478 (N_2478,In_680,In_383);
nand U2479 (N_2479,In_622,In_212);
or U2480 (N_2480,In_534,In_289);
or U2481 (N_2481,In_340,In_121);
xor U2482 (N_2482,In_716,In_172);
or U2483 (N_2483,In_188,In_582);
or U2484 (N_2484,In_352,In_348);
nand U2485 (N_2485,In_164,In_447);
xor U2486 (N_2486,In_557,In_476);
nor U2487 (N_2487,In_62,In_287);
nand U2488 (N_2488,In_591,In_701);
xor U2489 (N_2489,In_444,In_677);
xor U2490 (N_2490,In_734,In_185);
nor U2491 (N_2491,In_471,In_75);
nand U2492 (N_2492,In_704,In_130);
and U2493 (N_2493,In_243,In_598);
xor U2494 (N_2494,In_663,In_264);
nor U2495 (N_2495,In_328,In_45);
or U2496 (N_2496,In_719,In_541);
nor U2497 (N_2497,In_176,In_674);
nand U2498 (N_2498,In_530,In_380);
nand U2499 (N_2499,In_11,In_527);
nor U2500 (N_2500,N_633,N_711);
xor U2501 (N_2501,N_1121,N_2469);
nor U2502 (N_2502,N_240,N_2326);
nand U2503 (N_2503,N_323,N_792);
or U2504 (N_2504,N_125,N_423);
xnor U2505 (N_2505,N_2487,N_758);
nand U2506 (N_2506,N_1655,N_1408);
nor U2507 (N_2507,N_311,N_640);
nand U2508 (N_2508,N_582,N_2018);
xor U2509 (N_2509,N_190,N_1403);
nor U2510 (N_2510,N_2481,N_1821);
or U2511 (N_2511,N_570,N_1664);
nor U2512 (N_2512,N_2112,N_845);
or U2513 (N_2513,N_676,N_150);
nand U2514 (N_2514,N_1266,N_1443);
or U2515 (N_2515,N_838,N_732);
nand U2516 (N_2516,N_1240,N_1162);
xnor U2517 (N_2517,N_1004,N_210);
or U2518 (N_2518,N_77,N_1741);
and U2519 (N_2519,N_1380,N_927);
and U2520 (N_2520,N_218,N_348);
nand U2521 (N_2521,N_186,N_565);
and U2522 (N_2522,N_894,N_2460);
and U2523 (N_2523,N_1848,N_951);
xor U2524 (N_2524,N_1491,N_1826);
or U2525 (N_2525,N_607,N_1393);
xnor U2526 (N_2526,N_244,N_2003);
xnor U2527 (N_2527,N_1983,N_1563);
and U2528 (N_2528,N_841,N_2103);
nor U2529 (N_2529,N_1610,N_1493);
nor U2530 (N_2530,N_1918,N_117);
nand U2531 (N_2531,N_2447,N_2206);
xor U2532 (N_2532,N_2221,N_1994);
or U2533 (N_2533,N_2417,N_2352);
and U2534 (N_2534,N_655,N_1614);
xnor U2535 (N_2535,N_1310,N_664);
xor U2536 (N_2536,N_1750,N_2028);
xnor U2537 (N_2537,N_1947,N_1376);
and U2538 (N_2538,N_2023,N_1564);
and U2539 (N_2539,N_442,N_933);
or U2540 (N_2540,N_2466,N_1416);
or U2541 (N_2541,N_1718,N_1772);
or U2542 (N_2542,N_1690,N_384);
or U2543 (N_2543,N_2266,N_153);
or U2544 (N_2544,N_2302,N_174);
and U2545 (N_2545,N_1765,N_725);
xnor U2546 (N_2546,N_1253,N_2483);
and U2547 (N_2547,N_1836,N_2231);
or U2548 (N_2548,N_748,N_128);
nand U2549 (N_2549,N_2415,N_36);
nand U2550 (N_2550,N_372,N_1753);
or U2551 (N_2551,N_280,N_2060);
and U2552 (N_2552,N_394,N_945);
xor U2553 (N_2553,N_797,N_1406);
and U2554 (N_2554,N_245,N_1835);
and U2555 (N_2555,N_737,N_1845);
and U2556 (N_2556,N_2181,N_521);
xor U2557 (N_2557,N_928,N_177);
xor U2558 (N_2558,N_2226,N_512);
or U2559 (N_2559,N_1808,N_2342);
nor U2560 (N_2560,N_1472,N_445);
xnor U2561 (N_2561,N_1144,N_2201);
nor U2562 (N_2562,N_1878,N_662);
and U2563 (N_2563,N_1246,N_2457);
or U2564 (N_2564,N_182,N_1775);
or U2565 (N_2565,N_1239,N_2285);
or U2566 (N_2566,N_2488,N_1979);
nand U2567 (N_2567,N_784,N_843);
xnor U2568 (N_2568,N_2380,N_1801);
or U2569 (N_2569,N_538,N_2337);
or U2570 (N_2570,N_1041,N_1797);
xor U2571 (N_2571,N_1796,N_1489);
or U2572 (N_2572,N_2240,N_1023);
xnor U2573 (N_2573,N_226,N_249);
and U2574 (N_2574,N_2154,N_579);
nand U2575 (N_2575,N_149,N_2057);
or U2576 (N_2576,N_1386,N_411);
nor U2577 (N_2577,N_317,N_1701);
and U2578 (N_2578,N_357,N_2345);
nand U2579 (N_2579,N_2267,N_105);
nor U2580 (N_2580,N_808,N_28);
nor U2581 (N_2581,N_1577,N_1779);
nor U2582 (N_2582,N_287,N_2473);
nand U2583 (N_2583,N_1875,N_1851);
nand U2584 (N_2584,N_2413,N_1151);
and U2585 (N_2585,N_828,N_1462);
and U2586 (N_2586,N_984,N_1274);
xor U2587 (N_2587,N_704,N_624);
nand U2588 (N_2588,N_1748,N_1702);
xor U2589 (N_2589,N_1734,N_2127);
nand U2590 (N_2590,N_2051,N_1042);
xor U2591 (N_2591,N_740,N_1378);
xnor U2592 (N_2592,N_692,N_2265);
and U2593 (N_2593,N_449,N_1937);
nand U2594 (N_2594,N_453,N_284);
or U2595 (N_2595,N_2247,N_1817);
nand U2596 (N_2596,N_1375,N_681);
nor U2597 (N_2597,N_2261,N_212);
or U2598 (N_2598,N_1328,N_422);
and U2599 (N_2599,N_232,N_461);
nand U2600 (N_2600,N_2243,N_2048);
xnor U2601 (N_2601,N_1372,N_523);
nand U2602 (N_2602,N_2166,N_950);
nand U2603 (N_2603,N_2152,N_362);
and U2604 (N_2604,N_480,N_1663);
nor U2605 (N_2605,N_2377,N_638);
or U2606 (N_2606,N_2116,N_45);
xnor U2607 (N_2607,N_352,N_65);
or U2608 (N_2608,N_1357,N_266);
nor U2609 (N_2609,N_1215,N_1165);
nand U2610 (N_2610,N_1288,N_1658);
nor U2611 (N_2611,N_1133,N_1615);
nand U2612 (N_2612,N_1441,N_2188);
xnor U2613 (N_2613,N_1619,N_1620);
xnor U2614 (N_2614,N_1944,N_2349);
nor U2615 (N_2615,N_1930,N_248);
nand U2616 (N_2616,N_2066,N_650);
xnor U2617 (N_2617,N_1167,N_243);
and U2618 (N_2618,N_2210,N_2289);
nand U2619 (N_2619,N_1339,N_2427);
and U2620 (N_2620,N_1333,N_2096);
nand U2621 (N_2621,N_1127,N_691);
and U2622 (N_2622,N_626,N_499);
nand U2623 (N_2623,N_2175,N_654);
or U2624 (N_2624,N_1849,N_1833);
xor U2625 (N_2625,N_2128,N_1629);
nor U2626 (N_2626,N_2204,N_2219);
or U2627 (N_2627,N_645,N_421);
nand U2628 (N_2628,N_627,N_1208);
nor U2629 (N_2629,N_973,N_2043);
nor U2630 (N_2630,N_2198,N_1884);
and U2631 (N_2631,N_569,N_1649);
or U2632 (N_2632,N_388,N_0);
nand U2633 (N_2633,N_548,N_574);
nand U2634 (N_2634,N_269,N_2435);
nor U2635 (N_2635,N_2495,N_2085);
nand U2636 (N_2636,N_1461,N_800);
or U2637 (N_2637,N_1759,N_819);
and U2638 (N_2638,N_468,N_839);
xor U2639 (N_2639,N_1977,N_1975);
xor U2640 (N_2640,N_2179,N_1843);
nor U2641 (N_2641,N_630,N_1885);
and U2642 (N_2642,N_982,N_276);
nor U2643 (N_2643,N_549,N_519);
and U2644 (N_2644,N_223,N_333);
or U2645 (N_2645,N_884,N_1217);
nor U2646 (N_2646,N_134,N_1928);
and U2647 (N_2647,N_554,N_1680);
xor U2648 (N_2648,N_48,N_763);
and U2649 (N_2649,N_641,N_178);
and U2650 (N_2650,N_1300,N_2340);
nand U2651 (N_2651,N_169,N_1573);
xnor U2652 (N_2652,N_329,N_625);
and U2653 (N_2653,N_1017,N_1504);
xor U2654 (N_2654,N_1325,N_2133);
nand U2655 (N_2655,N_1738,N_2160);
or U2656 (N_2656,N_1621,N_899);
xor U2657 (N_2657,N_367,N_1400);
nand U2658 (N_2658,N_1883,N_215);
and U2659 (N_2659,N_2104,N_1374);
nand U2660 (N_2660,N_493,N_1128);
and U2661 (N_2661,N_1805,N_382);
and U2662 (N_2662,N_1496,N_404);
nand U2663 (N_2663,N_1929,N_917);
nand U2664 (N_2664,N_733,N_900);
nor U2665 (N_2665,N_990,N_619);
xor U2666 (N_2666,N_559,N_837);
or U2667 (N_2667,N_972,N_2109);
xnor U2668 (N_2668,N_4,N_1652);
and U2669 (N_2669,N_298,N_2017);
or U2670 (N_2670,N_1898,N_1784);
nor U2671 (N_2671,N_804,N_940);
or U2672 (N_2672,N_1897,N_386);
and U2673 (N_2673,N_1965,N_531);
xor U2674 (N_2674,N_2132,N_434);
nand U2675 (N_2675,N_1488,N_2189);
or U2676 (N_2676,N_1294,N_443);
nand U2677 (N_2677,N_2012,N_1896);
nor U2678 (N_2678,N_2455,N_1497);
nand U2679 (N_2679,N_987,N_255);
or U2680 (N_2680,N_2250,N_1740);
or U2681 (N_2681,N_330,N_482);
nor U2682 (N_2682,N_948,N_370);
or U2683 (N_2683,N_2329,N_1719);
xor U2684 (N_2684,N_2442,N_1671);
nor U2685 (N_2685,N_1450,N_1886);
and U2686 (N_2686,N_273,N_926);
and U2687 (N_2687,N_2262,N_809);
nor U2688 (N_2688,N_1440,N_2213);
nor U2689 (N_2689,N_206,N_1705);
or U2690 (N_2690,N_492,N_2004);
or U2691 (N_2691,N_889,N_2405);
nor U2692 (N_2692,N_1419,N_1478);
nor U2693 (N_2693,N_924,N_2429);
nor U2694 (N_2694,N_874,N_2007);
nand U2695 (N_2695,N_848,N_179);
and U2696 (N_2696,N_1551,N_1584);
and U2697 (N_2697,N_1685,N_974);
xnor U2698 (N_2698,N_1770,N_1180);
or U2699 (N_2699,N_2363,N_925);
or U2700 (N_2700,N_764,N_1911);
and U2701 (N_2701,N_2033,N_156);
xnor U2702 (N_2702,N_420,N_160);
nor U2703 (N_2703,N_1946,N_2387);
nor U2704 (N_2704,N_2318,N_198);
xor U2705 (N_2705,N_1430,N_199);
nor U2706 (N_2706,N_2046,N_1184);
nand U2707 (N_2707,N_1413,N_728);
nor U2708 (N_2708,N_2047,N_430);
and U2709 (N_2709,N_806,N_968);
or U2710 (N_2710,N_817,N_594);
or U2711 (N_2711,N_2426,N_1547);
and U2712 (N_2712,N_1308,N_1320);
xor U2713 (N_2713,N_1579,N_507);
nand U2714 (N_2714,N_2119,N_853);
nand U2715 (N_2715,N_349,N_458);
xor U2716 (N_2716,N_137,N_814);
nor U2717 (N_2717,N_490,N_257);
xnor U2718 (N_2718,N_2184,N_1495);
or U2719 (N_2719,N_1628,N_1316);
nor U2720 (N_2720,N_844,N_2145);
nor U2721 (N_2721,N_1192,N_1910);
or U2722 (N_2722,N_1912,N_1653);
nand U2723 (N_2723,N_660,N_1005);
nor U2724 (N_2724,N_1301,N_932);
nand U2725 (N_2725,N_2464,N_2183);
xnor U2726 (N_2726,N_2434,N_395);
nand U2727 (N_2727,N_673,N_2064);
xnor U2728 (N_2728,N_575,N_1455);
nor U2729 (N_2729,N_2063,N_1439);
or U2730 (N_2730,N_1263,N_376);
nand U2731 (N_2731,N_999,N_1029);
nor U2732 (N_2732,N_1353,N_605);
or U2733 (N_2733,N_913,N_1802);
xnor U2734 (N_2734,N_1974,N_428);
nand U2735 (N_2735,N_74,N_1035);
nand U2736 (N_2736,N_2115,N_1095);
xor U2737 (N_2737,N_82,N_2432);
or U2738 (N_2738,N_41,N_816);
xnor U2739 (N_2739,N_1703,N_1155);
xor U2740 (N_2740,N_2331,N_2146);
or U2741 (N_2741,N_2490,N_1732);
nand U2742 (N_2742,N_2208,N_425);
nor U2743 (N_2743,N_239,N_2238);
and U2744 (N_2744,N_2268,N_1346);
xor U2745 (N_2745,N_1199,N_868);
or U2746 (N_2746,N_2372,N_2304);
nand U2747 (N_2747,N_1526,N_1252);
nor U2748 (N_2748,N_2241,N_2344);
nor U2749 (N_2749,N_2348,N_229);
xor U2750 (N_2750,N_1140,N_1433);
and U2751 (N_2751,N_2290,N_447);
and U2752 (N_2752,N_791,N_1079);
and U2753 (N_2753,N_46,N_659);
nand U2754 (N_2754,N_1825,N_1656);
and U2755 (N_2755,N_2011,N_1053);
or U2756 (N_2756,N_50,N_354);
and U2757 (N_2757,N_258,N_1509);
xnor U2758 (N_2758,N_1395,N_405);
nor U2759 (N_2759,N_886,N_1880);
xnor U2760 (N_2760,N_1901,N_1587);
nand U2761 (N_2761,N_1015,N_862);
nand U2762 (N_2762,N_1694,N_43);
nand U2763 (N_2763,N_155,N_1137);
and U2764 (N_2764,N_2259,N_2379);
or U2765 (N_2765,N_885,N_1554);
nand U2766 (N_2766,N_2335,N_1210);
or U2767 (N_2767,N_1838,N_2359);
xnor U2768 (N_2768,N_2327,N_595);
nand U2769 (N_2769,N_55,N_1988);
or U2770 (N_2770,N_304,N_1613);
nand U2771 (N_2771,N_1066,N_1241);
and U2772 (N_2772,N_789,N_2232);
xnor U2773 (N_2773,N_1588,N_1641);
and U2774 (N_2774,N_1292,N_426);
nand U2775 (N_2775,N_1049,N_687);
nor U2776 (N_2776,N_1006,N_122);
nor U2777 (N_2777,N_2392,N_775);
nand U2778 (N_2778,N_2030,N_1752);
xnor U2779 (N_2779,N_558,N_1098);
or U2780 (N_2780,N_380,N_1695);
nor U2781 (N_2781,N_419,N_1742);
xor U2782 (N_2782,N_165,N_1224);
xnor U2783 (N_2783,N_1726,N_2217);
xor U2784 (N_2784,N_1962,N_2301);
and U2785 (N_2785,N_1206,N_1484);
or U2786 (N_2786,N_898,N_2026);
or U2787 (N_2787,N_344,N_242);
and U2788 (N_2788,N_441,N_1090);
and U2789 (N_2789,N_281,N_1307);
nand U2790 (N_2790,N_947,N_724);
and U2791 (N_2791,N_1948,N_1037);
or U2792 (N_2792,N_760,N_1211);
or U2793 (N_2793,N_985,N_1524);
or U2794 (N_2794,N_1687,N_1578);
nor U2795 (N_2795,N_157,N_1264);
nand U2796 (N_2796,N_38,N_1708);
nand U2797 (N_2797,N_1172,N_715);
xnor U2798 (N_2798,N_233,N_1560);
nor U2799 (N_2799,N_2177,N_1063);
xor U2800 (N_2800,N_1338,N_869);
or U2801 (N_2801,N_902,N_1113);
or U2802 (N_2802,N_1089,N_417);
or U2803 (N_2803,N_802,N_1340);
and U2804 (N_2804,N_342,N_1535);
nor U2805 (N_2805,N_589,N_1174);
or U2806 (N_2806,N_1754,N_1943);
xnor U2807 (N_2807,N_1200,N_592);
and U2808 (N_2808,N_1223,N_616);
nor U2809 (N_2809,N_2260,N_1709);
nand U2810 (N_2810,N_759,N_1635);
nor U2811 (N_2811,N_699,N_975);
nor U2812 (N_2812,N_992,N_37);
nand U2813 (N_2813,N_464,N_364);
nand U2814 (N_2814,N_345,N_1469);
xor U2815 (N_2815,N_259,N_1778);
xnor U2816 (N_2816,N_2126,N_1036);
or U2817 (N_2817,N_1024,N_251);
and U2818 (N_2818,N_998,N_1985);
nand U2819 (N_2819,N_1018,N_978);
nor U2820 (N_2820,N_912,N_1561);
and U2821 (N_2821,N_922,N_1360);
or U2822 (N_2822,N_92,N_2253);
xnor U2823 (N_2823,N_666,N_2167);
nor U2824 (N_2824,N_2074,N_256);
or U2825 (N_2825,N_1394,N_1522);
nor U2826 (N_2826,N_794,N_278);
and U2827 (N_2827,N_2422,N_2131);
nand U2828 (N_2828,N_1717,N_1899);
nor U2829 (N_2829,N_2092,N_1370);
nand U2830 (N_2830,N_846,N_1905);
and U2831 (N_2831,N_1030,N_562);
xnor U2832 (N_2832,N_221,N_2270);
or U2833 (N_2833,N_477,N_2022);
nand U2834 (N_2834,N_2255,N_587);
and U2835 (N_2835,N_2373,N_1214);
and U2836 (N_2836,N_66,N_1410);
nor U2837 (N_2837,N_2008,N_2078);
nand U2838 (N_2838,N_1083,N_2279);
and U2839 (N_2839,N_790,N_1069);
or U2840 (N_2840,N_1028,N_2484);
or U2841 (N_2841,N_306,N_339);
and U2842 (N_2842,N_1550,N_374);
or U2843 (N_2843,N_981,N_1618);
nand U2844 (N_2844,N_722,N_1026);
nor U2845 (N_2845,N_1016,N_811);
xnor U2846 (N_2846,N_2212,N_220);
and U2847 (N_2847,N_1764,N_1362);
or U2848 (N_2848,N_450,N_935);
and U2849 (N_2849,N_350,N_2376);
or U2850 (N_2850,N_942,N_2199);
xnor U2851 (N_2851,N_15,N_2273);
nand U2852 (N_2852,N_2052,N_1600);
nand U2853 (N_2853,N_1402,N_1681);
nand U2854 (N_2854,N_2358,N_1146);
or U2855 (N_2855,N_2263,N_668);
nor U2856 (N_2856,N_2401,N_2316);
and U2857 (N_2857,N_1860,N_861);
xor U2858 (N_2858,N_1534,N_2136);
xnor U2859 (N_2859,N_1429,N_54);
or U2860 (N_2860,N_1409,N_2264);
nand U2861 (N_2861,N_1303,N_1768);
xnor U2862 (N_2862,N_1583,N_2200);
nand U2863 (N_2863,N_1330,N_8);
and U2864 (N_2864,N_2411,N_1870);
or U2865 (N_2865,N_1516,N_1092);
nor U2866 (N_2866,N_1527,N_389);
nand U2867 (N_2867,N_327,N_1225);
nor U2868 (N_2868,N_1617,N_1706);
nand U2869 (N_2869,N_678,N_322);
or U2870 (N_2870,N_414,N_1660);
xnor U2871 (N_2871,N_1056,N_163);
xor U2872 (N_2872,N_871,N_2151);
nand U2873 (N_2873,N_980,N_2010);
xnor U2874 (N_2874,N_2142,N_2418);
nor U2875 (N_2875,N_1737,N_880);
or U2876 (N_2876,N_191,N_713);
nor U2877 (N_2877,N_2140,N_1071);
xor U2878 (N_2878,N_2024,N_2305);
xor U2879 (N_2879,N_695,N_2034);
nand U2880 (N_2880,N_1725,N_936);
xor U2881 (N_2881,N_2338,N_739);
and U2882 (N_2882,N_2328,N_1668);
xnor U2883 (N_2883,N_1099,N_1955);
nand U2884 (N_2884,N_1088,N_631);
and U2885 (N_2885,N_2367,N_1272);
nand U2886 (N_2886,N_1081,N_2158);
and U2887 (N_2887,N_69,N_738);
nand U2888 (N_2888,N_1281,N_1444);
or U2889 (N_2889,N_812,N_1842);
nand U2890 (N_2890,N_1730,N_1259);
or U2891 (N_2891,N_192,N_491);
and U2892 (N_2892,N_1463,N_14);
nor U2893 (N_2893,N_1574,N_200);
and U2894 (N_2894,N_1103,N_803);
nor U2895 (N_2895,N_2002,N_1058);
nand U2896 (N_2896,N_1729,N_2430);
nor U2897 (N_2897,N_1290,N_590);
or U2898 (N_2898,N_1492,N_1745);
xor U2899 (N_2899,N_1161,N_1);
nor U2900 (N_2900,N_1625,N_2317);
nand U2901 (N_2901,N_1498,N_1158);
nor U2902 (N_2902,N_1645,N_368);
or U2903 (N_2903,N_2229,N_2220);
xor U2904 (N_2904,N_866,N_1767);
and U2905 (N_2905,N_1822,N_700);
xnor U2906 (N_2906,N_2170,N_85);
nor U2907 (N_2907,N_1384,N_1149);
or U2908 (N_2908,N_1153,N_1830);
and U2909 (N_2909,N_1371,N_2439);
and U2910 (N_2910,N_2105,N_44);
nor U2911 (N_2911,N_543,N_1892);
or U2912 (N_2912,N_1157,N_2205);
or U2913 (N_2913,N_1917,N_247);
and U2914 (N_2914,N_164,N_1366);
and U2915 (N_2915,N_753,N_1939);
nand U2916 (N_2916,N_949,N_787);
or U2917 (N_2917,N_2006,N_2251);
and U2918 (N_2918,N_697,N_1420);
xnor U2919 (N_2919,N_2195,N_1335);
or U2920 (N_2920,N_2100,N_400);
nand U2921 (N_2921,N_1627,N_252);
nor U2922 (N_2922,N_1799,N_1879);
nand U2923 (N_2923,N_222,N_1678);
and U2924 (N_2924,N_1392,N_2203);
nand U2925 (N_2925,N_217,N_139);
or U2926 (N_2926,N_2339,N_2137);
nor U2927 (N_2927,N_2361,N_1093);
or U2928 (N_2928,N_636,N_675);
or U2929 (N_2929,N_2368,N_916);
nor U2930 (N_2930,N_1971,N_295);
nor U2931 (N_2931,N_1474,N_1397);
xor U2932 (N_2932,N_494,N_1841);
or U2933 (N_2933,N_1677,N_1204);
nand U2934 (N_2934,N_1611,N_1827);
nand U2935 (N_2935,N_1623,N_550);
and U2936 (N_2936,N_373,N_1033);
xor U2937 (N_2937,N_546,N_197);
and U2938 (N_2938,N_1811,N_2246);
and U2939 (N_2939,N_1934,N_1595);
xor U2940 (N_2940,N_873,N_1479);
nor U2941 (N_2941,N_1218,N_1072);
and U2942 (N_2942,N_392,N_771);
nand U2943 (N_2943,N_326,N_2468);
nand U2944 (N_2944,N_770,N_1604);
or U2945 (N_2945,N_285,N_1205);
nand U2946 (N_2946,N_1909,N_2300);
xnor U2947 (N_2947,N_1135,N_1227);
and U2948 (N_2948,N_1603,N_847);
nand U2949 (N_2949,N_1115,N_1508);
nor U2950 (N_2950,N_1993,N_189);
nand U2951 (N_2951,N_752,N_568);
nand U2952 (N_2952,N_2061,N_561);
nand U2953 (N_2953,N_1048,N_1987);
or U2954 (N_2954,N_24,N_1980);
xnor U2955 (N_2955,N_315,N_556);
and U2956 (N_2956,N_904,N_622);
nor U2957 (N_2957,N_1967,N_51);
nor U2958 (N_2958,N_1720,N_1916);
or U2959 (N_2959,N_765,N_166);
and U2960 (N_2960,N_923,N_1989);
and U2961 (N_2961,N_1565,N_402);
and U2962 (N_2962,N_1318,N_403);
and U2963 (N_2963,N_721,N_2465);
or U2964 (N_2964,N_1931,N_2117);
nand U2965 (N_2965,N_463,N_535);
nand U2966 (N_2966,N_2176,N_522);
or U2967 (N_2967,N_2347,N_93);
or U2968 (N_2968,N_1589,N_540);
and U2969 (N_2969,N_524,N_2248);
xor U2970 (N_2970,N_1874,N_1515);
xor U2971 (N_2971,N_2134,N_1052);
and U2972 (N_2972,N_286,N_11);
and U2973 (N_2973,N_822,N_986);
and U2974 (N_2974,N_9,N_1662);
or U2975 (N_2975,N_1887,N_623);
and U2976 (N_2976,N_1760,N_1519);
and U2977 (N_2977,N_2448,N_716);
nor U2978 (N_2978,N_892,N_1543);
xor U2979 (N_2979,N_16,N_1122);
xnor U2980 (N_2980,N_1986,N_1597);
and U2981 (N_2981,N_1721,N_1299);
or U2982 (N_2982,N_1859,N_2235);
xor U2983 (N_2983,N_1289,N_995);
nand U2984 (N_2984,N_2478,N_1130);
and U2985 (N_2985,N_2399,N_465);
nor U2986 (N_2986,N_509,N_1666);
or U2987 (N_2987,N_2333,N_112);
and U2988 (N_2988,N_1644,N_401);
xnor U2989 (N_2989,N_1234,N_56);
xor U2990 (N_2990,N_1156,N_130);
xor U2991 (N_2991,N_685,N_1132);
or U2992 (N_2992,N_920,N_1902);
and U2993 (N_2993,N_1869,N_1996);
xnor U2994 (N_2994,N_1755,N_1580);
and U2995 (N_2995,N_1216,N_1815);
nand U2996 (N_2996,N_635,N_573);
nor U2997 (N_2997,N_705,N_1511);
and U2998 (N_2998,N_1942,N_1735);
xor U2999 (N_2999,N_2313,N_291);
xor U3000 (N_3000,N_1990,N_639);
nor U3001 (N_3001,N_337,N_121);
nor U3002 (N_3002,N_1451,N_833);
and U3003 (N_3003,N_72,N_855);
nor U3004 (N_3004,N_1207,N_1776);
xnor U3005 (N_3005,N_444,N_416);
nor U3006 (N_3006,N_2297,N_823);
and U3007 (N_3007,N_1691,N_1314);
or U3008 (N_3008,N_1984,N_432);
xnor U3009 (N_3009,N_1958,N_1723);
nor U3010 (N_3010,N_1812,N_1659);
and U3011 (N_3011,N_282,N_647);
or U3012 (N_3012,N_882,N_1143);
nand U3013 (N_3013,N_1904,N_1185);
nand U3014 (N_3014,N_2293,N_718);
nor U3015 (N_3015,N_801,N_152);
nand U3016 (N_3016,N_727,N_1229);
nand U3017 (N_3017,N_1067,N_469);
or U3018 (N_3018,N_1693,N_1531);
or U3019 (N_3019,N_1387,N_864);
xor U3020 (N_3020,N_307,N_1782);
or U3021 (N_3021,N_661,N_653);
nor U3022 (N_3022,N_1622,N_1437);
or U3023 (N_3023,N_2089,N_17);
and U3024 (N_3024,N_473,N_346);
xor U3025 (N_3025,N_310,N_1514);
and U3026 (N_3026,N_476,N_827);
and U3027 (N_3027,N_1676,N_2314);
and U3028 (N_3028,N_994,N_1854);
and U3029 (N_3029,N_1852,N_1117);
xnor U3030 (N_3030,N_1548,N_964);
nand U3031 (N_3031,N_1293,N_27);
and U3032 (N_3032,N_1486,N_1178);
nor U3033 (N_3033,N_462,N_504);
nor U3034 (N_3034,N_1385,N_1139);
or U3035 (N_3035,N_2001,N_1698);
nor U3036 (N_3036,N_1555,N_1114);
and U3037 (N_3037,N_921,N_1201);
or U3038 (N_3038,N_541,N_993);
nand U3039 (N_3039,N_1212,N_1997);
xor U3040 (N_3040,N_195,N_2381);
and U3041 (N_3041,N_1170,N_2163);
nand U3042 (N_3042,N_496,N_1000);
nor U3043 (N_3043,N_263,N_415);
nand U3044 (N_3044,N_1173,N_1452);
xor U3045 (N_3045,N_2234,N_1256);
nand U3046 (N_3046,N_674,N_1327);
nand U3047 (N_3047,N_788,N_598);
nor U3048 (N_3048,N_2068,N_1710);
xnor U3049 (N_3049,N_183,N_1101);
nor U3050 (N_3050,N_293,N_966);
nor U3051 (N_3051,N_958,N_98);
and U3052 (N_3052,N_308,N_2303);
nand U3053 (N_3053,N_1481,N_1448);
nand U3054 (N_3054,N_2135,N_1168);
and U3055 (N_3055,N_1949,N_505);
and U3056 (N_3056,N_2106,N_96);
or U3057 (N_3057,N_749,N_2364);
nand U3058 (N_3058,N_1244,N_133);
xnor U3059 (N_3059,N_1570,N_1242);
nand U3060 (N_3060,N_2114,N_1945);
nor U3061 (N_3061,N_113,N_954);
xnor U3062 (N_3062,N_2065,N_1819);
xor U3063 (N_3063,N_1311,N_634);
nand U3064 (N_3064,N_1598,N_957);
or U3065 (N_3065,N_90,N_1104);
nor U3066 (N_3066,N_1341,N_1136);
or U3067 (N_3067,N_2282,N_318);
nor U3068 (N_3068,N_1190,N_1936);
and U3069 (N_3069,N_1536,N_498);
nor U3070 (N_3070,N_2071,N_1650);
or U3071 (N_3071,N_2271,N_1034);
or U3072 (N_3072,N_1935,N_850);
xnor U3073 (N_3073,N_2403,N_471);
nor U3074 (N_3074,N_95,N_1634);
nand U3075 (N_3075,N_1567,N_109);
xor U3076 (N_3076,N_1351,N_1425);
nand U3077 (N_3077,N_611,N_955);
nand U3078 (N_3078,N_881,N_2485);
nand U3079 (N_3079,N_825,N_2032);
xor U3080 (N_3080,N_2443,N_2389);
nand U3081 (N_3081,N_956,N_148);
or U3082 (N_3082,N_1633,N_1976);
or U3083 (N_3083,N_79,N_332);
nand U3084 (N_3084,N_2407,N_246);
nand U3085 (N_3085,N_983,N_1867);
and U3086 (N_3086,N_2121,N_102);
nor U3087 (N_3087,N_1715,N_919);
nand U3088 (N_3088,N_2312,N_2053);
nand U3089 (N_3089,N_511,N_2295);
and U3090 (N_3090,N_2366,N_1179);
nor U3091 (N_3091,N_1120,N_782);
xor U3092 (N_3092,N_601,N_409);
nand U3093 (N_3093,N_865,N_1692);
nand U3094 (N_3094,N_918,N_1468);
or U3095 (N_3095,N_2031,N_2130);
and U3096 (N_3096,N_2141,N_2182);
nand U3097 (N_3097,N_2491,N_2049);
nor U3098 (N_3098,N_1142,N_116);
xor U3099 (N_3099,N_383,N_1926);
nand U3100 (N_3100,N_366,N_1057);
nor U3101 (N_3101,N_2084,N_717);
xnor U3102 (N_3102,N_620,N_1840);
nand U3103 (N_3103,N_303,N_162);
xor U3104 (N_3104,N_1853,N_2088);
and U3105 (N_3105,N_2,N_1119);
and U3106 (N_3106,N_399,N_1435);
and U3107 (N_3107,N_667,N_474);
xnor U3108 (N_3108,N_632,N_1722);
nor U3109 (N_3109,N_1528,N_1038);
xor U3110 (N_3110,N_2230,N_1348);
or U3111 (N_3111,N_2185,N_515);
xor U3112 (N_3112,N_2284,N_2120);
xor U3113 (N_3113,N_1343,N_32);
nor U3114 (N_3114,N_140,N_343);
and U3115 (N_3115,N_867,N_1920);
nand U3116 (N_3116,N_446,N_2394);
nor U3117 (N_3117,N_1465,N_2336);
nand U3118 (N_3118,N_1591,N_860);
nor U3119 (N_3119,N_196,N_1800);
nand U3120 (N_3120,N_64,N_78);
nor U3121 (N_3121,N_67,N_1221);
and U3122 (N_3122,N_2471,N_580);
nand U3123 (N_3123,N_173,N_234);
nor U3124 (N_3124,N_1383,N_726);
nand U3125 (N_3125,N_617,N_2237);
xnor U3126 (N_3126,N_1739,N_1517);
nor U3127 (N_3127,N_1810,N_1027);
and U3128 (N_3128,N_365,N_1927);
or U3129 (N_3129,N_1183,N_1642);
xor U3130 (N_3130,N_1367,N_652);
or U3131 (N_3131,N_1585,N_2308);
and U3132 (N_3132,N_1107,N_1863);
xor U3133 (N_3133,N_840,N_241);
and U3134 (N_3134,N_2058,N_745);
or U3135 (N_3135,N_2187,N_1969);
or U3136 (N_3136,N_780,N_84);
xnor U3137 (N_3137,N_483,N_151);
xor U3138 (N_3138,N_120,N_300);
nor U3139 (N_3139,N_1485,N_381);
nand U3140 (N_3140,N_289,N_682);
and U3141 (N_3141,N_1972,N_1831);
or U3142 (N_3142,N_497,N_513);
nor U3143 (N_3143,N_1025,N_967);
xnor U3144 (N_3144,N_2402,N_1513);
xor U3145 (N_3145,N_1262,N_930);
xor U3146 (N_3146,N_2451,N_2014);
nor U3147 (N_3147,N_42,N_1674);
and U3148 (N_3148,N_988,N_187);
nand U3149 (N_3149,N_361,N_747);
nand U3150 (N_3150,N_2144,N_533);
nor U3151 (N_3151,N_2441,N_1590);
nand U3152 (N_3152,N_698,N_1607);
nor U3153 (N_3153,N_1537,N_2497);
nor U3154 (N_3154,N_1258,N_439);
and U3155 (N_3155,N_2498,N_21);
nor U3156 (N_3156,N_829,N_769);
nand U3157 (N_3157,N_1686,N_907);
xnor U3158 (N_3158,N_1487,N_1804);
nor U3159 (N_3159,N_2384,N_1950);
or U3160 (N_3160,N_1999,N_1606);
nor U3161 (N_3161,N_1321,N_325);
or U3162 (N_3162,N_888,N_1552);
nand U3163 (N_3163,N_2272,N_107);
nand U3164 (N_3164,N_1868,N_2445);
nand U3165 (N_3165,N_1781,N_2009);
nor U3166 (N_3166,N_1540,N_2281);
xor U3167 (N_3167,N_703,N_213);
xnor U3168 (N_3168,N_2207,N_887);
xor U3169 (N_3169,N_1544,N_714);
xor U3170 (N_3170,N_2147,N_1925);
nand U3171 (N_3171,N_1601,N_1315);
nand U3172 (N_3172,N_938,N_1291);
xnor U3173 (N_3173,N_1238,N_1297);
nor U3174 (N_3174,N_1814,N_2087);
or U3175 (N_3175,N_2156,N_2258);
nor U3176 (N_3176,N_262,N_2174);
nand U3177 (N_3177,N_2159,N_1533);
nor U3178 (N_3178,N_1070,N_1889);
xor U3179 (N_3179,N_876,N_2072);
or U3180 (N_3180,N_2287,N_2000);
nand U3181 (N_3181,N_1193,N_1744);
and U3182 (N_3182,N_1992,N_500);
nor U3183 (N_3183,N_895,N_1872);
nor U3184 (N_3184,N_1834,N_1235);
and U3185 (N_3185,N_1275,N_1746);
nor U3186 (N_3186,N_2013,N_1047);
nand U3187 (N_3187,N_205,N_34);
xor U3188 (N_3188,N_438,N_2076);
nand U3189 (N_3189,N_2178,N_106);
nand U3190 (N_3190,N_901,N_1636);
nor U3191 (N_3191,N_2041,N_750);
xor U3192 (N_3192,N_2165,N_1546);
nor U3193 (N_3193,N_776,N_1317);
and U3194 (N_3194,N_1941,N_1940);
nor U3195 (N_3195,N_2406,N_88);
xnor U3196 (N_3196,N_1302,N_1254);
xor U3197 (N_3197,N_1453,N_2249);
xnor U3198 (N_3198,N_1019,N_1922);
nand U3199 (N_3199,N_1756,N_2216);
nand U3200 (N_3200,N_970,N_1243);
and U3201 (N_3201,N_1045,N_2292);
and U3202 (N_3202,N_1464,N_1131);
nand U3203 (N_3203,N_1921,N_658);
xnor U3204 (N_3204,N_1747,N_1230);
nand U3205 (N_3205,N_1186,N_470);
and U3206 (N_3206,N_224,N_2351);
xor U3207 (N_3207,N_1358,N_1890);
and U3208 (N_3208,N_2493,N_2035);
and U3209 (N_3209,N_2256,N_2444);
nor U3210 (N_3210,N_1696,N_1365);
nand U3211 (N_3211,N_670,N_1347);
xor U3212 (N_3212,N_584,N_1247);
and U3213 (N_3213,N_1202,N_254);
nand U3214 (N_3214,N_2191,N_1806);
xor U3215 (N_3215,N_2080,N_1952);
xor U3216 (N_3216,N_1352,N_953);
or U3217 (N_3217,N_684,N_1159);
and U3218 (N_3218,N_2390,N_1777);
and U3219 (N_3219,N_1228,N_1111);
or U3220 (N_3220,N_2045,N_1457);
or U3221 (N_3221,N_99,N_2197);
nor U3222 (N_3222,N_1043,N_277);
or U3223 (N_3223,N_1900,N_883);
xnor U3224 (N_3224,N_2227,N_1388);
nor U3225 (N_3225,N_2244,N_911);
or U3226 (N_3226,N_597,N_997);
or U3227 (N_3227,N_407,N_831);
xor U3228 (N_3228,N_479,N_1631);
nor U3229 (N_3229,N_1039,N_1616);
xnor U3230 (N_3230,N_1427,N_2269);
xnor U3231 (N_3231,N_2218,N_710);
or U3232 (N_3232,N_893,N_1438);
xnor U3233 (N_3233,N_663,N_1684);
xor U3234 (N_3234,N_756,N_387);
xnor U3235 (N_3235,N_1332,N_1505);
nor U3236 (N_3236,N_830,N_746);
nor U3237 (N_3237,N_33,N_526);
xnor U3238 (N_3238,N_2019,N_610);
or U3239 (N_3239,N_111,N_679);
nand U3240 (N_3240,N_1296,N_1700);
nor U3241 (N_3241,N_1138,N_2157);
or U3242 (N_3242,N_1557,N_1689);
nand U3243 (N_3243,N_1682,N_94);
nor U3244 (N_3244,N_672,N_1471);
or U3245 (N_3245,N_1907,N_1426);
nor U3246 (N_3246,N_1350,N_1411);
nor U3247 (N_3247,N_1507,N_1542);
xor U3248 (N_3248,N_536,N_734);
nor U3249 (N_3249,N_2332,N_680);
nor U3250 (N_3250,N_2320,N_2067);
or U3251 (N_3251,N_578,N_2462);
and U3252 (N_3252,N_1003,N_910);
nor U3253 (N_3253,N_1198,N_2143);
or U3254 (N_3254,N_472,N_2382);
xor U3255 (N_3255,N_1231,N_1837);
xor U3256 (N_3256,N_1105,N_2306);
nor U3257 (N_3257,N_2474,N_144);
nor U3258 (N_3258,N_1084,N_460);
or U3259 (N_3259,N_2450,N_2391);
nand U3260 (N_3260,N_1189,N_851);
nor U3261 (N_3261,N_390,N_320);
or U3262 (N_3262,N_618,N_115);
or U3263 (N_3263,N_271,N_786);
xor U3264 (N_3264,N_762,N_1232);
nand U3265 (N_3265,N_1865,N_1319);
or U3266 (N_3266,N_502,N_1364);
nand U3267 (N_3267,N_1978,N_1787);
xor U3268 (N_3268,N_2412,N_1309);
xnor U3269 (N_3269,N_2298,N_1285);
nor U3270 (N_3270,N_1337,N_1991);
nor U3271 (N_3271,N_835,N_2428);
or U3272 (N_3272,N_1283,N_934);
xnor U3273 (N_3273,N_1373,N_1171);
nor U3274 (N_3274,N_1082,N_2343);
nand U3275 (N_3275,N_359,N_2162);
nor U3276 (N_3276,N_628,N_260);
or U3277 (N_3277,N_2192,N_71);
nor U3278 (N_3278,N_612,N_1475);
or U3279 (N_3279,N_1828,N_2118);
xor U3280 (N_3280,N_2409,N_1074);
and U3281 (N_3281,N_525,N_2330);
nand U3282 (N_3282,N_694,N_475);
or U3283 (N_3283,N_944,N_599);
xnor U3284 (N_3284,N_1771,N_1728);
or U3285 (N_3285,N_1749,N_1790);
and U3286 (N_3286,N_1342,N_1857);
or U3287 (N_3287,N_1418,N_2209);
xnor U3288 (N_3288,N_1431,N_2456);
nand U3289 (N_3289,N_1273,N_834);
or U3290 (N_3290,N_274,N_2423);
nor U3291 (N_3291,N_1602,N_2476);
and U3292 (N_3292,N_40,N_1704);
nor U3293 (N_3293,N_996,N_103);
nand U3294 (N_3294,N_1998,N_971);
or U3295 (N_3295,N_340,N_755);
and U3296 (N_3296,N_2388,N_859);
or U3297 (N_3297,N_730,N_2449);
or U3298 (N_3298,N_1882,N_1665);
nand U3299 (N_3299,N_962,N_1445);
nand U3300 (N_3300,N_591,N_532);
nor U3301 (N_3301,N_1336,N_1888);
and U3302 (N_3302,N_1525,N_1669);
nor U3303 (N_3303,N_1421,N_1582);
nor U3304 (N_3304,N_1009,N_646);
nor U3305 (N_3305,N_76,N_1279);
xor U3306 (N_3306,N_2094,N_1331);
nor U3307 (N_3307,N_793,N_1539);
and U3308 (N_3308,N_1575,N_1237);
xor U3309 (N_3309,N_1076,N_2055);
nand U3310 (N_3310,N_2395,N_671);
xor U3311 (N_3311,N_528,N_184);
nand U3312 (N_3312,N_637,N_1345);
nand U3313 (N_3313,N_572,N_2044);
and U3314 (N_3314,N_97,N_1713);
nor U3315 (N_3315,N_1792,N_914);
or U3316 (N_3316,N_1177,N_706);
nand U3317 (N_3317,N_1368,N_83);
and U3318 (N_3318,N_355,N_931);
and U3319 (N_3319,N_1398,N_2436);
nor U3320 (N_3320,N_237,N_1609);
xnor U3321 (N_3321,N_1097,N_1334);
xnor U3322 (N_3322,N_2223,N_451);
xor U3323 (N_3323,N_1401,N_2150);
nor U3324 (N_3324,N_288,N_2452);
and U3325 (N_3325,N_1716,N_2311);
nor U3326 (N_3326,N_1282,N_585);
xor U3327 (N_3327,N_1761,N_1995);
xor U3328 (N_3328,N_2425,N_1203);
xnor U3329 (N_3329,N_818,N_378);
nor U3330 (N_3330,N_1001,N_905);
and U3331 (N_3331,N_1306,N_1871);
or U3332 (N_3332,N_1672,N_2122);
nand U3333 (N_3333,N_1123,N_204);
xnor U3334 (N_3334,N_669,N_506);
nand U3335 (N_3335,N_1261,N_1793);
xnor U3336 (N_3336,N_2275,N_2321);
xor U3337 (N_3337,N_1040,N_2102);
nand U3338 (N_3338,N_1529,N_1683);
nand U3339 (N_3339,N_1415,N_302);
or U3340 (N_3340,N_2277,N_353);
and U3341 (N_3341,N_649,N_1512);
or U3342 (N_3342,N_1894,N_707);
nand U3343 (N_3343,N_778,N_2233);
and U3344 (N_3344,N_1954,N_517);
xor U3345 (N_3345,N_2486,N_1163);
and U3346 (N_3346,N_977,N_613);
nor U3347 (N_3347,N_170,N_1091);
nor U3348 (N_3348,N_1824,N_1236);
xnor U3349 (N_3349,N_2027,N_826);
nor U3350 (N_3350,N_2437,N_1654);
xnor U3351 (N_3351,N_2398,N_360);
and U3352 (N_3352,N_1846,N_454);
xor U3353 (N_3353,N_2360,N_172);
or U3354 (N_3354,N_397,N_1530);
or U3355 (N_3355,N_527,N_6);
nor U3356 (N_3356,N_118,N_1646);
and U3357 (N_3357,N_614,N_261);
nor U3358 (N_3358,N_135,N_1769);
and U3359 (N_3359,N_1592,N_1798);
xor U3360 (N_3360,N_2020,N_1124);
nand U3361 (N_3361,N_267,N_30);
and U3362 (N_3362,N_1521,N_608);
nand U3363 (N_3363,N_301,N_2355);
and U3364 (N_3364,N_70,N_406);
or U3365 (N_3365,N_331,N_25);
xor U3366 (N_3366,N_101,N_216);
nand U3367 (N_3367,N_227,N_1809);
xor U3368 (N_3368,N_2242,N_1112);
nand U3369 (N_3369,N_379,N_1807);
nor U3370 (N_3370,N_1458,N_396);
xor U3371 (N_3371,N_1304,N_2062);
nor U3372 (N_3372,N_1456,N_1449);
or U3373 (N_3373,N_2374,N_796);
nor U3374 (N_3374,N_294,N_1785);
nand U3375 (N_3375,N_1640,N_159);
or U3376 (N_3376,N_1571,N_2280);
nor U3377 (N_3377,N_188,N_1324);
and U3378 (N_3378,N_943,N_341);
or U3379 (N_3379,N_773,N_2393);
or U3380 (N_3380,N_1538,N_433);
and U3381 (N_3381,N_2470,N_1913);
nand U3382 (N_3382,N_1923,N_751);
xnor U3383 (N_3383,N_1788,N_1599);
xnor U3384 (N_3384,N_2499,N_2161);
nand U3385 (N_3385,N_1847,N_1423);
nor U3386 (N_3386,N_2149,N_1220);
nor U3387 (N_3387,N_2274,N_781);
nand U3388 (N_3388,N_604,N_566);
or U3389 (N_3389,N_2101,N_723);
nor U3390 (N_3390,N_1326,N_854);
xnor U3391 (N_3391,N_236,N_126);
nand U3392 (N_3392,N_503,N_486);
and U3393 (N_3393,N_1050,N_1109);
xor U3394 (N_3394,N_2059,N_2356);
or U3395 (N_3395,N_299,N_124);
nor U3396 (N_3396,N_1568,N_815);
or U3397 (N_3397,N_2309,N_2077);
nor U3398 (N_3398,N_731,N_143);
or U3399 (N_3399,N_1046,N_202);
and U3400 (N_3400,N_1844,N_1277);
nand U3401 (N_3401,N_1377,N_1818);
or U3402 (N_3402,N_1194,N_1724);
and U3403 (N_3403,N_2310,N_297);
or U3404 (N_3404,N_208,N_2056);
nor U3405 (N_3405,N_1391,N_1476);
and U3406 (N_3406,N_596,N_648);
nor U3407 (N_3407,N_1855,N_1699);
nand U3408 (N_3408,N_1280,N_1532);
nand U3409 (N_3409,N_129,N_238);
xor U3410 (N_3410,N_1490,N_313);
and U3411 (N_3411,N_1399,N_171);
nand U3412 (N_3412,N_2440,N_2424);
nand U3413 (N_3413,N_1803,N_1096);
or U3414 (N_3414,N_1981,N_2397);
nor U3415 (N_3415,N_363,N_1518);
xor U3416 (N_3416,N_1094,N_693);
or U3417 (N_3417,N_1670,N_1305);
xor U3418 (N_3418,N_466,N_2354);
xnor U3419 (N_3419,N_897,N_1866);
nand U3420 (N_3420,N_896,N_358);
nand U3421 (N_3421,N_1973,N_1477);
or U3422 (N_3422,N_2257,N_2083);
nor U3423 (N_3423,N_2016,N_767);
and U3424 (N_3424,N_1011,N_1502);
nand U3425 (N_3425,N_1250,N_1751);
or U3426 (N_3426,N_2431,N_720);
xor U3427 (N_3427,N_795,N_1510);
xnor U3428 (N_3428,N_1651,N_1219);
and U3429 (N_3429,N_2186,N_1593);
and U3430 (N_3430,N_1780,N_228);
and U3431 (N_3431,N_1446,N_534);
and U3432 (N_3432,N_1118,N_1382);
and U3433 (N_3433,N_2239,N_547);
xor U3434 (N_3434,N_1813,N_742);
or U3435 (N_3435,N_448,N_459);
and U3436 (N_3436,N_209,N_2042);
nand U3437 (N_3437,N_1245,N_1483);
or U3438 (N_3438,N_1964,N_193);
and U3439 (N_3439,N_856,N_1428);
and U3440 (N_3440,N_741,N_2021);
xor U3441 (N_3441,N_1520,N_1085);
or U3442 (N_3442,N_455,N_516);
nor U3443 (N_3443,N_1862,N_1356);
and U3444 (N_3444,N_564,N_1626);
and U3445 (N_3445,N_1482,N_1010);
and U3446 (N_3446,N_201,N_696);
xor U3447 (N_3447,N_1960,N_690);
nand U3448 (N_3448,N_219,N_1956);
or U3449 (N_3449,N_10,N_2369);
and U3450 (N_3450,N_1014,N_1032);
and U3451 (N_3451,N_2370,N_2324);
or U3452 (N_3452,N_1675,N_712);
or U3453 (N_3453,N_2172,N_452);
xnor U3454 (N_3454,N_136,N_35);
and U3455 (N_3455,N_1963,N_73);
and U3456 (N_3456,N_1915,N_1624);
nor U3457 (N_3457,N_2433,N_849);
nand U3458 (N_3458,N_960,N_832);
nand U3459 (N_3459,N_709,N_272);
or U3460 (N_3460,N_1313,N_1829);
xor U3461 (N_3461,N_61,N_18);
xor U3462 (N_3462,N_552,N_1166);
nand U3463 (N_3463,N_487,N_729);
nand U3464 (N_3464,N_963,N_427);
or U3465 (N_3465,N_1612,N_1816);
and U3466 (N_3466,N_1466,N_2416);
nor U3467 (N_3467,N_283,N_230);
or U3468 (N_3468,N_2438,N_408);
and U3469 (N_3469,N_1417,N_385);
xor U3470 (N_3470,N_2086,N_132);
nor U3471 (N_3471,N_1379,N_2168);
nor U3472 (N_3472,N_185,N_544);
and U3473 (N_3473,N_1044,N_2005);
nand U3474 (N_3474,N_754,N_26);
xnor U3475 (N_3475,N_976,N_1116);
or U3476 (N_3476,N_2245,N_131);
xnor U3477 (N_3477,N_321,N_813);
or U3478 (N_3478,N_2288,N_1774);
nand U3479 (N_3479,N_2383,N_2453);
nor U3480 (N_3480,N_2283,N_1638);
xnor U3481 (N_3481,N_1460,N_772);
nand U3482 (N_3482,N_1763,N_314);
nand U3483 (N_3483,N_2419,N_1637);
and U3484 (N_3484,N_60,N_154);
and U3485 (N_3485,N_49,N_583);
nand U3486 (N_3486,N_1322,N_2458);
nand U3487 (N_3487,N_1390,N_1251);
or U3488 (N_3488,N_1007,N_1459);
nand U3489 (N_3489,N_2073,N_100);
and U3490 (N_3490,N_1354,N_563);
or U3491 (N_3491,N_1657,N_1523);
or U3492 (N_3492,N_1148,N_1639);
nor U3493 (N_3493,N_2252,N_890);
xnor U3494 (N_3494,N_657,N_1298);
or U3495 (N_3495,N_296,N_316);
nand U3496 (N_3496,N_81,N_1447);
nand U3497 (N_3497,N_1647,N_104);
nand U3498 (N_3498,N_312,N_1953);
nand U3499 (N_3499,N_1160,N_2362);
xor U3500 (N_3500,N_551,N_766);
xnor U3501 (N_3501,N_1503,N_588);
xor U3502 (N_3502,N_161,N_961);
nor U3503 (N_3503,N_5,N_292);
nor U3504 (N_3504,N_1020,N_1667);
xnor U3505 (N_3505,N_2299,N_2463);
or U3506 (N_3506,N_456,N_1404);
or U3507 (N_3507,N_2236,N_265);
or U3508 (N_3508,N_2171,N_520);
or U3509 (N_3509,N_484,N_761);
and U3510 (N_3510,N_375,N_19);
or U3511 (N_3511,N_2420,N_2286);
xor U3512 (N_3512,N_478,N_824);
xnor U3513 (N_3513,N_2054,N_702);
nor U3514 (N_3514,N_1494,N_1506);
nor U3515 (N_3515,N_1970,N_665);
nand U3516 (N_3516,N_1500,N_991);
or U3517 (N_3517,N_1002,N_2025);
or U3518 (N_3518,N_2482,N_2494);
and U3519 (N_3519,N_1697,N_412);
nor U3520 (N_3520,N_1569,N_1197);
nand U3521 (N_3521,N_488,N_576);
nand U3522 (N_3522,N_2069,N_2029);
xor U3523 (N_3523,N_1608,N_2404);
nor U3524 (N_3524,N_1012,N_2472);
xor U3525 (N_3525,N_1268,N_878);
or U3526 (N_3526,N_2093,N_147);
nor U3527 (N_3527,N_602,N_264);
nand U3528 (N_3528,N_615,N_2479);
or U3529 (N_3529,N_110,N_1078);
or U3530 (N_3530,N_47,N_1850);
and U3531 (N_3531,N_398,N_39);
or U3532 (N_3532,N_1312,N_80);
or U3533 (N_3533,N_2353,N_119);
nand U3534 (N_3534,N_677,N_1549);
and U3535 (N_3535,N_593,N_1369);
and U3536 (N_3536,N_1576,N_2291);
nor U3537 (N_3537,N_437,N_2386);
nor U3538 (N_3538,N_1766,N_467);
xnor U3539 (N_3539,N_127,N_1422);
xor U3540 (N_3540,N_1267,N_1643);
or U3541 (N_3541,N_2040,N_1856);
nor U3542 (N_3542,N_1087,N_557);
and U3543 (N_3543,N_1714,N_2113);
or U3544 (N_3544,N_2139,N_12);
and U3545 (N_3545,N_1959,N_903);
nand U3546 (N_3546,N_145,N_424);
xnor U3547 (N_3547,N_2467,N_1594);
and U3548 (N_3548,N_1154,N_858);
nand U3549 (N_3549,N_909,N_501);
nand U3550 (N_3550,N_872,N_2346);
nor U3551 (N_3551,N_621,N_952);
xor U3552 (N_3552,N_270,N_2496);
and U3553 (N_3553,N_1982,N_807);
and U3554 (N_3554,N_2222,N_2400);
nand U3555 (N_3555,N_175,N_2153);
and U3556 (N_3556,N_440,N_1396);
or U3557 (N_3557,N_377,N_1467);
nor U3558 (N_3558,N_1541,N_2070);
nand U3559 (N_3559,N_1924,N_180);
or U3560 (N_3560,N_768,N_719);
xor U3561 (N_3561,N_744,N_1176);
and U3562 (N_3562,N_1733,N_2164);
and U3563 (N_3563,N_1432,N_1255);
or U3564 (N_3564,N_1270,N_959);
xnor U3565 (N_3565,N_581,N_1249);
or U3566 (N_3566,N_2079,N_309);
xor U3567 (N_3567,N_1213,N_1932);
nand U3568 (N_3568,N_1061,N_2211);
and U3569 (N_3569,N_1414,N_1661);
and U3570 (N_3570,N_606,N_810);
nand U3571 (N_3571,N_168,N_1820);
nand U3572 (N_3572,N_1858,N_820);
nor U3573 (N_3573,N_836,N_1791);
or U3574 (N_3574,N_1175,N_1269);
nor U3575 (N_3575,N_2341,N_1966);
or U3576 (N_3576,N_2148,N_1073);
or U3577 (N_3577,N_2446,N_1068);
or U3578 (N_3578,N_52,N_821);
and U3579 (N_3579,N_877,N_937);
xnor U3580 (N_3580,N_1581,N_2111);
or U3581 (N_3581,N_324,N_2224);
and U3582 (N_3582,N_1265,N_686);
nand U3583 (N_3583,N_89,N_1271);
xnor U3584 (N_3584,N_785,N_1596);
and U3585 (N_3585,N_2107,N_2123);
nand U3586 (N_3586,N_2015,N_194);
xnor U3587 (N_3587,N_1182,N_644);
and U3588 (N_3588,N_1773,N_537);
xor U3589 (N_3589,N_908,N_1126);
xnor U3590 (N_3590,N_542,N_1054);
and U3591 (N_3591,N_351,N_1679);
nand U3592 (N_3592,N_2202,N_1233);
or U3593 (N_3593,N_2036,N_915);
nor U3594 (N_3594,N_1389,N_481);
nor U3595 (N_3595,N_736,N_2180);
nand U3596 (N_3596,N_777,N_2480);
xnor U3597 (N_3597,N_530,N_1630);
nand U3598 (N_3598,N_1473,N_1553);
or U3599 (N_3599,N_2276,N_603);
nand U3600 (N_3600,N_1075,N_1147);
xnor U3601 (N_3601,N_1260,N_1454);
xor U3602 (N_3602,N_2138,N_2489);
nand U3603 (N_3603,N_1839,N_508);
xnor U3604 (N_3604,N_906,N_1295);
nand U3605 (N_3605,N_1480,N_857);
and U3606 (N_3606,N_1903,N_290);
nor U3607 (N_3607,N_1442,N_2278);
or U3608 (N_3608,N_2414,N_435);
or U3609 (N_3609,N_1344,N_1794);
xnor U3610 (N_3610,N_2365,N_1381);
nor U3611 (N_3611,N_2190,N_1743);
nand U3612 (N_3612,N_1558,N_2169);
and U3613 (N_3613,N_2129,N_2214);
nand U3614 (N_3614,N_31,N_1169);
nand U3615 (N_3615,N_1876,N_567);
xnor U3616 (N_3616,N_1731,N_2410);
or U3617 (N_3617,N_1187,N_138);
or U3618 (N_3618,N_1957,N_1873);
xnor U3619 (N_3619,N_1736,N_231);
nand U3620 (N_3620,N_891,N_2421);
nor U3621 (N_3621,N_207,N_1586);
or U3622 (N_3622,N_1864,N_1908);
or U3623 (N_3623,N_1572,N_1795);
or U3624 (N_3624,N_1919,N_2098);
or U3625 (N_3625,N_600,N_391);
nor U3626 (N_3626,N_68,N_1191);
and U3627 (N_3627,N_1021,N_1059);
xnor U3628 (N_3628,N_336,N_356);
nand U3629 (N_3629,N_22,N_1758);
and U3630 (N_3630,N_1110,N_1424);
xor U3631 (N_3631,N_1893,N_743);
and U3632 (N_3632,N_1501,N_1951);
nor U3633 (N_3633,N_2095,N_842);
or U3634 (N_3634,N_560,N_2228);
xor U3635 (N_3635,N_2357,N_2196);
and U3636 (N_3636,N_2039,N_1757);
nor U3637 (N_3637,N_1906,N_1181);
xnor U3638 (N_3638,N_2296,N_689);
or U3639 (N_3639,N_53,N_1361);
and U3640 (N_3640,N_1141,N_1355);
and U3641 (N_3641,N_929,N_20);
nand U3642 (N_3642,N_2075,N_969);
nand U3643 (N_3643,N_2215,N_1881);
xor U3644 (N_3644,N_1861,N_1832);
and U3645 (N_3645,N_708,N_495);
or U3646 (N_3646,N_779,N_989);
nor U3647 (N_3647,N_2461,N_1823);
nand U3648 (N_3648,N_2385,N_2254);
and U3649 (N_3649,N_852,N_176);
nor U3650 (N_3650,N_13,N_2108);
and U3651 (N_3651,N_1013,N_2371);
nor U3652 (N_3652,N_870,N_181);
and U3653 (N_3653,N_609,N_418);
nand U3654 (N_3654,N_879,N_1164);
nor U3655 (N_3655,N_863,N_319);
and U3656 (N_3656,N_683,N_1407);
and U3657 (N_3657,N_1961,N_1707);
nor U3658 (N_3658,N_146,N_1008);
and U3659 (N_3659,N_489,N_1145);
nor U3660 (N_3660,N_1257,N_1064);
xnor U3661 (N_3661,N_2097,N_2173);
nand U3662 (N_3662,N_2408,N_141);
xnor U3663 (N_3663,N_1673,N_1031);
and U3664 (N_3664,N_757,N_1278);
nand U3665 (N_3665,N_58,N_553);
nand U3666 (N_3666,N_369,N_2315);
or U3667 (N_3667,N_1129,N_586);
nand U3668 (N_3668,N_1329,N_235);
nor U3669 (N_3669,N_108,N_23);
and U3670 (N_3670,N_1727,N_275);
nand U3671 (N_3671,N_2091,N_571);
xnor U3672 (N_3672,N_75,N_1648);
and U3673 (N_3673,N_643,N_334);
or U3674 (N_3674,N_2375,N_2378);
nor U3675 (N_3675,N_2350,N_1363);
and U3676 (N_3676,N_735,N_86);
xor U3677 (N_3677,N_1022,N_518);
or U3678 (N_3678,N_142,N_1559);
xor U3679 (N_3679,N_1712,N_3);
or U3680 (N_3680,N_965,N_413);
nor U3681 (N_3681,N_253,N_268);
and U3682 (N_3682,N_875,N_1566);
nand U3683 (N_3683,N_1222,N_1323);
and U3684 (N_3684,N_1783,N_2323);
and U3685 (N_3685,N_1789,N_1108);
nor U3686 (N_3686,N_1150,N_1077);
xnor U3687 (N_3687,N_1349,N_158);
nand U3688 (N_3688,N_2325,N_123);
nand U3689 (N_3689,N_1914,N_1152);
nor U3690 (N_3690,N_2125,N_2193);
or U3691 (N_3691,N_1632,N_2322);
nor U3692 (N_3692,N_2081,N_941);
nor U3693 (N_3693,N_1762,N_1499);
xor U3694 (N_3694,N_29,N_1051);
nand U3695 (N_3695,N_2038,N_2307);
nor U3696 (N_3696,N_1188,N_87);
nand U3697 (N_3697,N_431,N_1287);
xnor U3698 (N_3698,N_2082,N_1102);
nor U3699 (N_3699,N_167,N_2155);
nor U3700 (N_3700,N_979,N_2124);
and U3701 (N_3701,N_62,N_2492);
nand U3702 (N_3702,N_1086,N_279);
nor U3703 (N_3703,N_1436,N_2090);
or U3704 (N_3704,N_2477,N_783);
nand U3705 (N_3705,N_1786,N_2294);
nor U3706 (N_3706,N_1286,N_1412);
nor U3707 (N_3707,N_1196,N_328);
xor U3708 (N_3708,N_688,N_1877);
nor U3709 (N_3709,N_7,N_1405);
nor U3710 (N_3710,N_1711,N_1891);
nor U3711 (N_3711,N_799,N_1195);
nand U3712 (N_3712,N_214,N_2459);
xor U3713 (N_3713,N_1968,N_57);
and U3714 (N_3714,N_393,N_1545);
xor U3715 (N_3715,N_1556,N_545);
nand U3716 (N_3716,N_1060,N_629);
xor U3717 (N_3717,N_63,N_1938);
and U3718 (N_3718,N_1688,N_114);
xor U3719 (N_3719,N_2475,N_798);
and U3720 (N_3720,N_347,N_939);
xnor U3721 (N_3721,N_211,N_371);
and U3722 (N_3722,N_91,N_555);
xor U3723 (N_3723,N_2225,N_1359);
xnor U3724 (N_3724,N_2396,N_1080);
xnor U3725 (N_3725,N_1933,N_1895);
nor U3726 (N_3726,N_1434,N_1125);
or U3727 (N_3727,N_1605,N_2454);
xnor U3728 (N_3728,N_59,N_1055);
and U3729 (N_3729,N_305,N_1134);
xnor U3730 (N_3730,N_1248,N_805);
xor U3731 (N_3731,N_1226,N_946);
or U3732 (N_3732,N_1209,N_429);
xnor U3733 (N_3733,N_1065,N_539);
xor U3734 (N_3734,N_701,N_577);
or U3735 (N_3735,N_1106,N_2110);
nor U3736 (N_3736,N_436,N_656);
nand U3737 (N_3737,N_485,N_1276);
and U3738 (N_3738,N_510,N_2099);
xor U3739 (N_3739,N_529,N_642);
xnor U3740 (N_3740,N_2319,N_1062);
nand U3741 (N_3741,N_2037,N_335);
nor U3742 (N_3742,N_1100,N_250);
or U3743 (N_3743,N_338,N_1470);
and U3744 (N_3744,N_514,N_203);
xnor U3745 (N_3745,N_1284,N_410);
xnor U3746 (N_3746,N_225,N_2194);
nor U3747 (N_3747,N_1562,N_2050);
nor U3748 (N_3748,N_774,N_457);
nand U3749 (N_3749,N_651,N_2334);
nor U3750 (N_3750,N_619,N_2489);
nor U3751 (N_3751,N_47,N_1234);
nand U3752 (N_3752,N_447,N_1193);
nor U3753 (N_3753,N_369,N_719);
nor U3754 (N_3754,N_1965,N_2388);
xnor U3755 (N_3755,N_1450,N_358);
xor U3756 (N_3756,N_402,N_1435);
nand U3757 (N_3757,N_1461,N_1951);
or U3758 (N_3758,N_385,N_2399);
or U3759 (N_3759,N_2015,N_863);
and U3760 (N_3760,N_2185,N_1176);
xnor U3761 (N_3761,N_661,N_1418);
and U3762 (N_3762,N_618,N_1736);
nor U3763 (N_3763,N_2181,N_682);
xnor U3764 (N_3764,N_2497,N_2324);
xor U3765 (N_3765,N_1822,N_1636);
and U3766 (N_3766,N_1962,N_2282);
nor U3767 (N_3767,N_1210,N_1498);
or U3768 (N_3768,N_1584,N_1749);
or U3769 (N_3769,N_1882,N_1278);
nor U3770 (N_3770,N_1935,N_106);
xor U3771 (N_3771,N_2310,N_1391);
nor U3772 (N_3772,N_1929,N_1991);
xor U3773 (N_3773,N_1790,N_600);
and U3774 (N_3774,N_31,N_1998);
or U3775 (N_3775,N_2469,N_2126);
xnor U3776 (N_3776,N_2286,N_642);
or U3777 (N_3777,N_1096,N_2316);
xor U3778 (N_3778,N_1722,N_189);
and U3779 (N_3779,N_1713,N_1468);
and U3780 (N_3780,N_179,N_312);
or U3781 (N_3781,N_2427,N_815);
or U3782 (N_3782,N_1115,N_1602);
nor U3783 (N_3783,N_1094,N_1581);
or U3784 (N_3784,N_793,N_1445);
or U3785 (N_3785,N_1053,N_1402);
and U3786 (N_3786,N_1186,N_973);
or U3787 (N_3787,N_1958,N_877);
or U3788 (N_3788,N_2109,N_1225);
and U3789 (N_3789,N_682,N_1855);
nor U3790 (N_3790,N_1050,N_1507);
xnor U3791 (N_3791,N_1394,N_1225);
nand U3792 (N_3792,N_454,N_1758);
or U3793 (N_3793,N_778,N_2349);
xnor U3794 (N_3794,N_891,N_1310);
nor U3795 (N_3795,N_499,N_1433);
xnor U3796 (N_3796,N_405,N_2131);
or U3797 (N_3797,N_1966,N_1725);
and U3798 (N_3798,N_2231,N_1319);
or U3799 (N_3799,N_2387,N_2433);
nor U3800 (N_3800,N_915,N_333);
and U3801 (N_3801,N_1344,N_171);
xor U3802 (N_3802,N_1152,N_427);
or U3803 (N_3803,N_2172,N_1229);
and U3804 (N_3804,N_958,N_123);
nand U3805 (N_3805,N_1255,N_1500);
nand U3806 (N_3806,N_154,N_1979);
and U3807 (N_3807,N_876,N_1805);
or U3808 (N_3808,N_2273,N_564);
nand U3809 (N_3809,N_1852,N_740);
nor U3810 (N_3810,N_2478,N_2302);
and U3811 (N_3811,N_1992,N_421);
or U3812 (N_3812,N_1867,N_1544);
and U3813 (N_3813,N_371,N_241);
nor U3814 (N_3814,N_943,N_266);
or U3815 (N_3815,N_1466,N_2002);
xor U3816 (N_3816,N_1787,N_2265);
nand U3817 (N_3817,N_749,N_2489);
or U3818 (N_3818,N_1584,N_2289);
and U3819 (N_3819,N_801,N_1960);
nand U3820 (N_3820,N_855,N_1165);
nand U3821 (N_3821,N_1369,N_179);
nor U3822 (N_3822,N_2053,N_1474);
nand U3823 (N_3823,N_1300,N_200);
nand U3824 (N_3824,N_1895,N_2155);
xnor U3825 (N_3825,N_905,N_2351);
or U3826 (N_3826,N_1592,N_1468);
nand U3827 (N_3827,N_1421,N_1745);
and U3828 (N_3828,N_2306,N_385);
nor U3829 (N_3829,N_573,N_853);
nand U3830 (N_3830,N_716,N_203);
nand U3831 (N_3831,N_1002,N_1502);
nor U3832 (N_3832,N_1737,N_896);
nand U3833 (N_3833,N_1161,N_784);
xnor U3834 (N_3834,N_1469,N_1382);
or U3835 (N_3835,N_786,N_1404);
or U3836 (N_3836,N_2166,N_1449);
xnor U3837 (N_3837,N_1011,N_941);
and U3838 (N_3838,N_2225,N_808);
nor U3839 (N_3839,N_749,N_2212);
xor U3840 (N_3840,N_854,N_1621);
xor U3841 (N_3841,N_2012,N_2202);
and U3842 (N_3842,N_544,N_2383);
or U3843 (N_3843,N_168,N_1042);
or U3844 (N_3844,N_1907,N_1465);
or U3845 (N_3845,N_1451,N_525);
or U3846 (N_3846,N_348,N_803);
or U3847 (N_3847,N_1980,N_1157);
xor U3848 (N_3848,N_1430,N_913);
nor U3849 (N_3849,N_1780,N_322);
nor U3850 (N_3850,N_2476,N_2393);
xnor U3851 (N_3851,N_1330,N_851);
nor U3852 (N_3852,N_1767,N_439);
nor U3853 (N_3853,N_1734,N_252);
and U3854 (N_3854,N_2237,N_555);
and U3855 (N_3855,N_498,N_2029);
nand U3856 (N_3856,N_65,N_2284);
nor U3857 (N_3857,N_1271,N_467);
nand U3858 (N_3858,N_287,N_635);
nand U3859 (N_3859,N_1400,N_1830);
or U3860 (N_3860,N_889,N_1523);
xor U3861 (N_3861,N_1691,N_1991);
xor U3862 (N_3862,N_749,N_2211);
nand U3863 (N_3863,N_6,N_1270);
nor U3864 (N_3864,N_2054,N_485);
or U3865 (N_3865,N_1146,N_1047);
nand U3866 (N_3866,N_1398,N_884);
xnor U3867 (N_3867,N_1848,N_208);
and U3868 (N_3868,N_389,N_1422);
nor U3869 (N_3869,N_2321,N_703);
xor U3870 (N_3870,N_1271,N_830);
nand U3871 (N_3871,N_2433,N_2235);
and U3872 (N_3872,N_966,N_385);
or U3873 (N_3873,N_1824,N_148);
xnor U3874 (N_3874,N_2178,N_2392);
nand U3875 (N_3875,N_1497,N_7);
and U3876 (N_3876,N_1600,N_1028);
nor U3877 (N_3877,N_2026,N_1234);
and U3878 (N_3878,N_851,N_193);
and U3879 (N_3879,N_1902,N_1552);
nor U3880 (N_3880,N_2272,N_2180);
and U3881 (N_3881,N_2065,N_957);
or U3882 (N_3882,N_1320,N_1556);
nor U3883 (N_3883,N_629,N_823);
xnor U3884 (N_3884,N_2398,N_475);
nor U3885 (N_3885,N_1763,N_299);
or U3886 (N_3886,N_909,N_327);
and U3887 (N_3887,N_1258,N_1684);
or U3888 (N_3888,N_2346,N_703);
and U3889 (N_3889,N_642,N_1864);
nor U3890 (N_3890,N_2287,N_22);
nor U3891 (N_3891,N_1610,N_822);
and U3892 (N_3892,N_545,N_478);
nand U3893 (N_3893,N_2401,N_2479);
nand U3894 (N_3894,N_2469,N_1877);
or U3895 (N_3895,N_746,N_1836);
nor U3896 (N_3896,N_378,N_1043);
nand U3897 (N_3897,N_362,N_222);
and U3898 (N_3898,N_2060,N_83);
nor U3899 (N_3899,N_1278,N_408);
and U3900 (N_3900,N_1834,N_1367);
xor U3901 (N_3901,N_10,N_1261);
and U3902 (N_3902,N_377,N_645);
or U3903 (N_3903,N_251,N_1012);
nand U3904 (N_3904,N_103,N_2262);
and U3905 (N_3905,N_17,N_2276);
or U3906 (N_3906,N_228,N_1976);
nor U3907 (N_3907,N_910,N_756);
xnor U3908 (N_3908,N_333,N_546);
nor U3909 (N_3909,N_2335,N_1687);
and U3910 (N_3910,N_1133,N_1173);
xor U3911 (N_3911,N_833,N_925);
nand U3912 (N_3912,N_660,N_175);
and U3913 (N_3913,N_109,N_2043);
nor U3914 (N_3914,N_1498,N_1569);
nor U3915 (N_3915,N_1193,N_1796);
nand U3916 (N_3916,N_977,N_19);
nor U3917 (N_3917,N_55,N_898);
and U3918 (N_3918,N_1472,N_1388);
and U3919 (N_3919,N_1802,N_755);
or U3920 (N_3920,N_2144,N_1261);
xor U3921 (N_3921,N_1081,N_957);
xnor U3922 (N_3922,N_1314,N_2434);
nor U3923 (N_3923,N_2257,N_2013);
and U3924 (N_3924,N_1294,N_885);
and U3925 (N_3925,N_1918,N_353);
nand U3926 (N_3926,N_647,N_469);
nand U3927 (N_3927,N_1110,N_2385);
nor U3928 (N_3928,N_1336,N_1515);
or U3929 (N_3929,N_1961,N_8);
nand U3930 (N_3930,N_95,N_2388);
and U3931 (N_3931,N_251,N_1847);
nand U3932 (N_3932,N_803,N_911);
and U3933 (N_3933,N_929,N_580);
nor U3934 (N_3934,N_734,N_1868);
xor U3935 (N_3935,N_951,N_600);
and U3936 (N_3936,N_665,N_860);
nor U3937 (N_3937,N_535,N_2081);
nand U3938 (N_3938,N_392,N_1766);
and U3939 (N_3939,N_1076,N_50);
nor U3940 (N_3940,N_1422,N_1994);
nand U3941 (N_3941,N_1199,N_2211);
nand U3942 (N_3942,N_147,N_970);
xnor U3943 (N_3943,N_1151,N_781);
nand U3944 (N_3944,N_433,N_1371);
xor U3945 (N_3945,N_2481,N_1361);
or U3946 (N_3946,N_895,N_1263);
xor U3947 (N_3947,N_2142,N_987);
nor U3948 (N_3948,N_570,N_1483);
nand U3949 (N_3949,N_2490,N_2288);
or U3950 (N_3950,N_1033,N_64);
xnor U3951 (N_3951,N_1106,N_634);
nor U3952 (N_3952,N_2280,N_431);
nand U3953 (N_3953,N_600,N_584);
nor U3954 (N_3954,N_1578,N_144);
or U3955 (N_3955,N_784,N_26);
nand U3956 (N_3956,N_472,N_455);
and U3957 (N_3957,N_360,N_1287);
xor U3958 (N_3958,N_1401,N_623);
or U3959 (N_3959,N_2380,N_433);
or U3960 (N_3960,N_1661,N_305);
nor U3961 (N_3961,N_1000,N_573);
and U3962 (N_3962,N_2328,N_829);
or U3963 (N_3963,N_1260,N_757);
and U3964 (N_3964,N_60,N_1327);
nor U3965 (N_3965,N_700,N_810);
or U3966 (N_3966,N_448,N_2332);
or U3967 (N_3967,N_2239,N_739);
nand U3968 (N_3968,N_1105,N_1442);
or U3969 (N_3969,N_1252,N_480);
nand U3970 (N_3970,N_1070,N_1820);
nand U3971 (N_3971,N_368,N_900);
nor U3972 (N_3972,N_1287,N_518);
or U3973 (N_3973,N_943,N_1892);
or U3974 (N_3974,N_621,N_1140);
xnor U3975 (N_3975,N_2085,N_874);
nand U3976 (N_3976,N_147,N_1734);
xor U3977 (N_3977,N_2140,N_134);
xnor U3978 (N_3978,N_1623,N_1466);
and U3979 (N_3979,N_1991,N_451);
nor U3980 (N_3980,N_2045,N_471);
nand U3981 (N_3981,N_1973,N_351);
or U3982 (N_3982,N_1397,N_1268);
or U3983 (N_3983,N_294,N_1327);
and U3984 (N_3984,N_642,N_2334);
or U3985 (N_3985,N_108,N_676);
nor U3986 (N_3986,N_1253,N_1705);
nor U3987 (N_3987,N_434,N_163);
xor U3988 (N_3988,N_1404,N_2349);
xor U3989 (N_3989,N_1289,N_1673);
nor U3990 (N_3990,N_1514,N_621);
xnor U3991 (N_3991,N_2081,N_1427);
xnor U3992 (N_3992,N_1544,N_998);
and U3993 (N_3993,N_1019,N_1481);
nand U3994 (N_3994,N_2092,N_166);
or U3995 (N_3995,N_1668,N_1838);
nor U3996 (N_3996,N_677,N_954);
and U3997 (N_3997,N_1037,N_200);
xor U3998 (N_3998,N_1537,N_442);
or U3999 (N_3999,N_2150,N_316);
and U4000 (N_4000,N_473,N_571);
nand U4001 (N_4001,N_483,N_2138);
or U4002 (N_4002,N_1815,N_1317);
and U4003 (N_4003,N_684,N_1587);
nor U4004 (N_4004,N_741,N_38);
or U4005 (N_4005,N_517,N_2181);
and U4006 (N_4006,N_2201,N_784);
xnor U4007 (N_4007,N_509,N_1138);
or U4008 (N_4008,N_1368,N_953);
xor U4009 (N_4009,N_2248,N_2455);
nand U4010 (N_4010,N_2212,N_2289);
nand U4011 (N_4011,N_631,N_1697);
or U4012 (N_4012,N_343,N_2170);
and U4013 (N_4013,N_1713,N_1031);
xor U4014 (N_4014,N_1089,N_1364);
xnor U4015 (N_4015,N_1502,N_2318);
nor U4016 (N_4016,N_344,N_961);
xnor U4017 (N_4017,N_2184,N_511);
and U4018 (N_4018,N_1921,N_1676);
or U4019 (N_4019,N_1848,N_304);
nor U4020 (N_4020,N_1948,N_2131);
xnor U4021 (N_4021,N_991,N_2043);
xor U4022 (N_4022,N_118,N_393);
xnor U4023 (N_4023,N_2026,N_1553);
nor U4024 (N_4024,N_2493,N_2104);
and U4025 (N_4025,N_1488,N_2387);
and U4026 (N_4026,N_1343,N_1632);
nor U4027 (N_4027,N_730,N_2482);
xor U4028 (N_4028,N_939,N_1129);
nand U4029 (N_4029,N_814,N_404);
xor U4030 (N_4030,N_35,N_1380);
xor U4031 (N_4031,N_1301,N_1274);
nor U4032 (N_4032,N_1399,N_342);
nor U4033 (N_4033,N_1214,N_876);
and U4034 (N_4034,N_1854,N_861);
and U4035 (N_4035,N_1519,N_1523);
nor U4036 (N_4036,N_2250,N_387);
xnor U4037 (N_4037,N_215,N_2334);
nand U4038 (N_4038,N_2253,N_1054);
xnor U4039 (N_4039,N_1775,N_1318);
nand U4040 (N_4040,N_1015,N_658);
nor U4041 (N_4041,N_2224,N_1976);
nand U4042 (N_4042,N_1048,N_37);
or U4043 (N_4043,N_640,N_1611);
xnor U4044 (N_4044,N_1663,N_1937);
and U4045 (N_4045,N_111,N_120);
or U4046 (N_4046,N_2247,N_869);
and U4047 (N_4047,N_978,N_1851);
or U4048 (N_4048,N_1920,N_780);
or U4049 (N_4049,N_812,N_630);
or U4050 (N_4050,N_48,N_923);
xor U4051 (N_4051,N_994,N_741);
and U4052 (N_4052,N_921,N_1187);
nor U4053 (N_4053,N_1522,N_387);
nand U4054 (N_4054,N_1840,N_1172);
or U4055 (N_4055,N_1354,N_1033);
nand U4056 (N_4056,N_2037,N_663);
nand U4057 (N_4057,N_1995,N_1403);
or U4058 (N_4058,N_807,N_1251);
nor U4059 (N_4059,N_253,N_486);
xnor U4060 (N_4060,N_1072,N_1246);
nor U4061 (N_4061,N_21,N_100);
nand U4062 (N_4062,N_565,N_1697);
and U4063 (N_4063,N_269,N_2110);
xor U4064 (N_4064,N_2224,N_1467);
and U4065 (N_4065,N_1592,N_563);
nand U4066 (N_4066,N_1741,N_1924);
nor U4067 (N_4067,N_2005,N_2235);
or U4068 (N_4068,N_1649,N_1551);
and U4069 (N_4069,N_190,N_542);
xor U4070 (N_4070,N_730,N_2343);
or U4071 (N_4071,N_63,N_479);
or U4072 (N_4072,N_2224,N_1453);
or U4073 (N_4073,N_1965,N_1020);
nand U4074 (N_4074,N_1809,N_1852);
and U4075 (N_4075,N_316,N_2397);
or U4076 (N_4076,N_272,N_2461);
nand U4077 (N_4077,N_1776,N_1947);
or U4078 (N_4078,N_1581,N_1920);
nand U4079 (N_4079,N_555,N_1742);
nand U4080 (N_4080,N_558,N_2467);
or U4081 (N_4081,N_1640,N_85);
nor U4082 (N_4082,N_1281,N_537);
or U4083 (N_4083,N_304,N_1479);
nand U4084 (N_4084,N_671,N_619);
nand U4085 (N_4085,N_1868,N_1644);
nand U4086 (N_4086,N_1380,N_147);
nand U4087 (N_4087,N_1114,N_1393);
nand U4088 (N_4088,N_380,N_2145);
nor U4089 (N_4089,N_1898,N_1668);
nor U4090 (N_4090,N_770,N_1889);
or U4091 (N_4091,N_2193,N_1366);
or U4092 (N_4092,N_557,N_1959);
nand U4093 (N_4093,N_1199,N_1591);
and U4094 (N_4094,N_2305,N_2093);
xor U4095 (N_4095,N_1050,N_2037);
nor U4096 (N_4096,N_2007,N_460);
nor U4097 (N_4097,N_1977,N_1389);
nand U4098 (N_4098,N_2471,N_115);
and U4099 (N_4099,N_2127,N_549);
nor U4100 (N_4100,N_1688,N_2204);
nor U4101 (N_4101,N_193,N_808);
nand U4102 (N_4102,N_2058,N_1363);
nand U4103 (N_4103,N_1203,N_990);
nor U4104 (N_4104,N_1304,N_1678);
xnor U4105 (N_4105,N_1764,N_1165);
and U4106 (N_4106,N_203,N_86);
and U4107 (N_4107,N_1533,N_1185);
or U4108 (N_4108,N_1021,N_1993);
nand U4109 (N_4109,N_462,N_1358);
and U4110 (N_4110,N_904,N_415);
nand U4111 (N_4111,N_883,N_167);
and U4112 (N_4112,N_438,N_1804);
and U4113 (N_4113,N_2353,N_521);
and U4114 (N_4114,N_1123,N_158);
nand U4115 (N_4115,N_1368,N_121);
and U4116 (N_4116,N_242,N_2079);
nand U4117 (N_4117,N_945,N_326);
or U4118 (N_4118,N_568,N_2224);
and U4119 (N_4119,N_771,N_462);
nor U4120 (N_4120,N_619,N_1913);
nand U4121 (N_4121,N_1155,N_1998);
nand U4122 (N_4122,N_2021,N_816);
or U4123 (N_4123,N_1050,N_2459);
and U4124 (N_4124,N_2328,N_293);
or U4125 (N_4125,N_1213,N_1357);
xor U4126 (N_4126,N_1160,N_440);
xnor U4127 (N_4127,N_629,N_1899);
nand U4128 (N_4128,N_2136,N_627);
or U4129 (N_4129,N_1737,N_1054);
and U4130 (N_4130,N_2268,N_188);
nor U4131 (N_4131,N_644,N_810);
nand U4132 (N_4132,N_2317,N_494);
and U4133 (N_4133,N_2166,N_111);
nor U4134 (N_4134,N_1653,N_451);
or U4135 (N_4135,N_1841,N_567);
nor U4136 (N_4136,N_617,N_549);
nand U4137 (N_4137,N_975,N_2207);
and U4138 (N_4138,N_557,N_145);
xor U4139 (N_4139,N_122,N_1065);
or U4140 (N_4140,N_260,N_2155);
nand U4141 (N_4141,N_222,N_976);
xor U4142 (N_4142,N_1578,N_580);
and U4143 (N_4143,N_1950,N_319);
and U4144 (N_4144,N_936,N_1347);
xnor U4145 (N_4145,N_635,N_1508);
nor U4146 (N_4146,N_159,N_2494);
xor U4147 (N_4147,N_902,N_2245);
nor U4148 (N_4148,N_1588,N_550);
nand U4149 (N_4149,N_1683,N_1811);
xnor U4150 (N_4150,N_2217,N_303);
xnor U4151 (N_4151,N_1123,N_1725);
xnor U4152 (N_4152,N_2074,N_795);
or U4153 (N_4153,N_1633,N_308);
or U4154 (N_4154,N_964,N_1940);
nor U4155 (N_4155,N_1841,N_362);
xnor U4156 (N_4156,N_535,N_2090);
or U4157 (N_4157,N_581,N_2015);
xnor U4158 (N_4158,N_583,N_392);
xnor U4159 (N_4159,N_1210,N_972);
and U4160 (N_4160,N_1963,N_1145);
nor U4161 (N_4161,N_349,N_1749);
xnor U4162 (N_4162,N_1415,N_1075);
xnor U4163 (N_4163,N_251,N_1700);
and U4164 (N_4164,N_2217,N_697);
and U4165 (N_4165,N_563,N_1758);
nor U4166 (N_4166,N_571,N_2100);
nor U4167 (N_4167,N_1881,N_1305);
nor U4168 (N_4168,N_322,N_902);
xnor U4169 (N_4169,N_289,N_564);
nand U4170 (N_4170,N_352,N_511);
nand U4171 (N_4171,N_260,N_1663);
nand U4172 (N_4172,N_543,N_1078);
or U4173 (N_4173,N_2424,N_2403);
nand U4174 (N_4174,N_246,N_1359);
and U4175 (N_4175,N_1238,N_1127);
nand U4176 (N_4176,N_2390,N_1437);
xnor U4177 (N_4177,N_202,N_1979);
nand U4178 (N_4178,N_1967,N_549);
or U4179 (N_4179,N_2136,N_1759);
or U4180 (N_4180,N_449,N_1511);
or U4181 (N_4181,N_2244,N_1889);
and U4182 (N_4182,N_2173,N_2181);
nand U4183 (N_4183,N_320,N_1523);
or U4184 (N_4184,N_1539,N_2139);
and U4185 (N_4185,N_1139,N_205);
and U4186 (N_4186,N_906,N_1524);
xor U4187 (N_4187,N_1916,N_406);
nor U4188 (N_4188,N_534,N_184);
nor U4189 (N_4189,N_794,N_1583);
and U4190 (N_4190,N_1393,N_2411);
nand U4191 (N_4191,N_530,N_477);
xnor U4192 (N_4192,N_1128,N_2044);
and U4193 (N_4193,N_2353,N_892);
nor U4194 (N_4194,N_612,N_1443);
nor U4195 (N_4195,N_2439,N_905);
nand U4196 (N_4196,N_1086,N_723);
nor U4197 (N_4197,N_1550,N_1745);
and U4198 (N_4198,N_291,N_526);
nand U4199 (N_4199,N_2350,N_178);
nand U4200 (N_4200,N_2020,N_590);
nor U4201 (N_4201,N_1149,N_2483);
nor U4202 (N_4202,N_659,N_1644);
or U4203 (N_4203,N_1199,N_1372);
nand U4204 (N_4204,N_1826,N_1355);
nor U4205 (N_4205,N_1874,N_827);
nand U4206 (N_4206,N_1442,N_843);
or U4207 (N_4207,N_1333,N_2177);
xor U4208 (N_4208,N_1113,N_2192);
or U4209 (N_4209,N_519,N_2166);
nor U4210 (N_4210,N_928,N_830);
nand U4211 (N_4211,N_2374,N_454);
or U4212 (N_4212,N_1600,N_31);
and U4213 (N_4213,N_927,N_2156);
or U4214 (N_4214,N_262,N_535);
nand U4215 (N_4215,N_1999,N_847);
or U4216 (N_4216,N_1426,N_935);
nor U4217 (N_4217,N_870,N_2412);
or U4218 (N_4218,N_2061,N_1706);
or U4219 (N_4219,N_482,N_873);
nor U4220 (N_4220,N_209,N_587);
xnor U4221 (N_4221,N_417,N_2494);
xor U4222 (N_4222,N_771,N_1312);
nor U4223 (N_4223,N_718,N_2201);
and U4224 (N_4224,N_2389,N_62);
and U4225 (N_4225,N_12,N_2207);
or U4226 (N_4226,N_407,N_2207);
and U4227 (N_4227,N_2057,N_1561);
and U4228 (N_4228,N_804,N_718);
and U4229 (N_4229,N_468,N_1663);
nand U4230 (N_4230,N_662,N_1142);
nand U4231 (N_4231,N_1767,N_282);
nor U4232 (N_4232,N_676,N_2089);
xnor U4233 (N_4233,N_796,N_1407);
or U4234 (N_4234,N_927,N_1496);
nand U4235 (N_4235,N_1608,N_2180);
xor U4236 (N_4236,N_2170,N_1294);
nor U4237 (N_4237,N_1209,N_549);
or U4238 (N_4238,N_573,N_1431);
xor U4239 (N_4239,N_2003,N_2444);
xnor U4240 (N_4240,N_2080,N_1434);
nand U4241 (N_4241,N_128,N_425);
xor U4242 (N_4242,N_1804,N_1816);
nand U4243 (N_4243,N_2405,N_1113);
or U4244 (N_4244,N_777,N_819);
nor U4245 (N_4245,N_615,N_856);
xnor U4246 (N_4246,N_1319,N_29);
and U4247 (N_4247,N_959,N_117);
and U4248 (N_4248,N_1650,N_737);
xor U4249 (N_4249,N_413,N_2098);
xnor U4250 (N_4250,N_1602,N_112);
nor U4251 (N_4251,N_887,N_791);
xor U4252 (N_4252,N_2097,N_2277);
or U4253 (N_4253,N_389,N_288);
and U4254 (N_4254,N_349,N_217);
xor U4255 (N_4255,N_1748,N_1202);
nor U4256 (N_4256,N_1829,N_2250);
nand U4257 (N_4257,N_898,N_712);
nor U4258 (N_4258,N_261,N_1152);
and U4259 (N_4259,N_2061,N_2164);
or U4260 (N_4260,N_107,N_1986);
nor U4261 (N_4261,N_1606,N_1022);
nand U4262 (N_4262,N_2150,N_67);
and U4263 (N_4263,N_734,N_1626);
nand U4264 (N_4264,N_246,N_628);
nand U4265 (N_4265,N_1133,N_886);
and U4266 (N_4266,N_1024,N_1967);
and U4267 (N_4267,N_1394,N_22);
and U4268 (N_4268,N_758,N_168);
xor U4269 (N_4269,N_198,N_1613);
nor U4270 (N_4270,N_950,N_1003);
nand U4271 (N_4271,N_323,N_329);
and U4272 (N_4272,N_844,N_147);
or U4273 (N_4273,N_1750,N_2073);
and U4274 (N_4274,N_1185,N_585);
nand U4275 (N_4275,N_773,N_2187);
nor U4276 (N_4276,N_2261,N_43);
and U4277 (N_4277,N_2104,N_1955);
nor U4278 (N_4278,N_306,N_1565);
and U4279 (N_4279,N_1190,N_164);
nor U4280 (N_4280,N_793,N_2291);
nand U4281 (N_4281,N_281,N_844);
and U4282 (N_4282,N_2474,N_1936);
xnor U4283 (N_4283,N_126,N_851);
xnor U4284 (N_4284,N_1123,N_833);
or U4285 (N_4285,N_668,N_1549);
or U4286 (N_4286,N_689,N_1875);
nor U4287 (N_4287,N_894,N_778);
or U4288 (N_4288,N_36,N_2349);
nor U4289 (N_4289,N_151,N_2439);
and U4290 (N_4290,N_2233,N_1811);
or U4291 (N_4291,N_1295,N_2373);
or U4292 (N_4292,N_417,N_584);
or U4293 (N_4293,N_1293,N_1082);
nand U4294 (N_4294,N_1571,N_1681);
and U4295 (N_4295,N_1517,N_2345);
xnor U4296 (N_4296,N_1607,N_407);
nor U4297 (N_4297,N_240,N_1975);
nor U4298 (N_4298,N_2358,N_1470);
nand U4299 (N_4299,N_785,N_1915);
nor U4300 (N_4300,N_1167,N_1381);
xor U4301 (N_4301,N_724,N_1181);
xor U4302 (N_4302,N_1337,N_394);
nand U4303 (N_4303,N_24,N_2128);
and U4304 (N_4304,N_2277,N_980);
or U4305 (N_4305,N_2260,N_318);
xnor U4306 (N_4306,N_792,N_1552);
xor U4307 (N_4307,N_808,N_1936);
nor U4308 (N_4308,N_2310,N_1691);
xor U4309 (N_4309,N_1357,N_1215);
and U4310 (N_4310,N_2108,N_265);
or U4311 (N_4311,N_1441,N_2369);
nor U4312 (N_4312,N_2110,N_1600);
xor U4313 (N_4313,N_1961,N_96);
or U4314 (N_4314,N_1863,N_587);
nand U4315 (N_4315,N_1116,N_1267);
nand U4316 (N_4316,N_1882,N_741);
nand U4317 (N_4317,N_2335,N_397);
or U4318 (N_4318,N_218,N_2357);
or U4319 (N_4319,N_132,N_974);
or U4320 (N_4320,N_308,N_2472);
nand U4321 (N_4321,N_2145,N_2430);
xnor U4322 (N_4322,N_2486,N_427);
or U4323 (N_4323,N_1855,N_1083);
nand U4324 (N_4324,N_1546,N_484);
and U4325 (N_4325,N_1435,N_880);
nand U4326 (N_4326,N_199,N_1997);
xor U4327 (N_4327,N_2001,N_449);
nor U4328 (N_4328,N_884,N_248);
xnor U4329 (N_4329,N_2154,N_271);
nand U4330 (N_4330,N_1723,N_1265);
and U4331 (N_4331,N_1882,N_1724);
or U4332 (N_4332,N_114,N_739);
and U4333 (N_4333,N_1775,N_1652);
and U4334 (N_4334,N_1523,N_2098);
nor U4335 (N_4335,N_2388,N_1286);
or U4336 (N_4336,N_1456,N_2431);
or U4337 (N_4337,N_1875,N_1048);
xnor U4338 (N_4338,N_87,N_1692);
or U4339 (N_4339,N_197,N_1099);
xnor U4340 (N_4340,N_936,N_1340);
or U4341 (N_4341,N_1004,N_310);
nor U4342 (N_4342,N_50,N_595);
nor U4343 (N_4343,N_626,N_1318);
and U4344 (N_4344,N_765,N_1777);
xor U4345 (N_4345,N_1515,N_2138);
and U4346 (N_4346,N_183,N_1406);
nor U4347 (N_4347,N_902,N_1562);
nor U4348 (N_4348,N_2064,N_1283);
nor U4349 (N_4349,N_844,N_50);
nand U4350 (N_4350,N_99,N_1649);
or U4351 (N_4351,N_45,N_1055);
nand U4352 (N_4352,N_850,N_2122);
nor U4353 (N_4353,N_1773,N_1420);
or U4354 (N_4354,N_741,N_2420);
and U4355 (N_4355,N_1034,N_1075);
nor U4356 (N_4356,N_2178,N_1947);
xor U4357 (N_4357,N_1641,N_389);
nor U4358 (N_4358,N_2344,N_1601);
nor U4359 (N_4359,N_414,N_1308);
and U4360 (N_4360,N_278,N_2065);
or U4361 (N_4361,N_28,N_1165);
or U4362 (N_4362,N_1460,N_1621);
nand U4363 (N_4363,N_1125,N_1667);
or U4364 (N_4364,N_1899,N_1193);
nor U4365 (N_4365,N_428,N_2375);
nand U4366 (N_4366,N_2099,N_1551);
nor U4367 (N_4367,N_2134,N_63);
and U4368 (N_4368,N_388,N_594);
or U4369 (N_4369,N_1372,N_1904);
xnor U4370 (N_4370,N_1310,N_2170);
nand U4371 (N_4371,N_403,N_95);
or U4372 (N_4372,N_434,N_2110);
and U4373 (N_4373,N_269,N_1006);
or U4374 (N_4374,N_1537,N_2175);
and U4375 (N_4375,N_1990,N_2156);
or U4376 (N_4376,N_1473,N_1486);
and U4377 (N_4377,N_462,N_1863);
xnor U4378 (N_4378,N_696,N_1189);
or U4379 (N_4379,N_170,N_1289);
nand U4380 (N_4380,N_154,N_1616);
nor U4381 (N_4381,N_2258,N_333);
and U4382 (N_4382,N_2455,N_2385);
and U4383 (N_4383,N_704,N_1621);
xor U4384 (N_4384,N_812,N_2432);
or U4385 (N_4385,N_2096,N_1566);
nor U4386 (N_4386,N_2119,N_272);
nand U4387 (N_4387,N_1178,N_1929);
nor U4388 (N_4388,N_1459,N_1778);
nand U4389 (N_4389,N_1251,N_1825);
and U4390 (N_4390,N_328,N_1508);
xnor U4391 (N_4391,N_1376,N_1495);
nand U4392 (N_4392,N_998,N_2476);
nand U4393 (N_4393,N_2293,N_367);
xor U4394 (N_4394,N_524,N_1147);
nor U4395 (N_4395,N_1688,N_2063);
nand U4396 (N_4396,N_1556,N_911);
xor U4397 (N_4397,N_405,N_1099);
nor U4398 (N_4398,N_1417,N_1560);
and U4399 (N_4399,N_755,N_426);
nand U4400 (N_4400,N_289,N_1033);
nand U4401 (N_4401,N_31,N_1981);
and U4402 (N_4402,N_845,N_1118);
nor U4403 (N_4403,N_307,N_1300);
nand U4404 (N_4404,N_642,N_913);
nor U4405 (N_4405,N_1268,N_541);
and U4406 (N_4406,N_1529,N_321);
and U4407 (N_4407,N_581,N_999);
or U4408 (N_4408,N_875,N_1299);
nor U4409 (N_4409,N_512,N_480);
or U4410 (N_4410,N_1460,N_959);
nor U4411 (N_4411,N_1647,N_142);
or U4412 (N_4412,N_748,N_2306);
and U4413 (N_4413,N_2481,N_781);
nand U4414 (N_4414,N_830,N_1599);
nand U4415 (N_4415,N_1284,N_1957);
nor U4416 (N_4416,N_1734,N_1404);
nor U4417 (N_4417,N_988,N_2244);
nor U4418 (N_4418,N_1152,N_1563);
nor U4419 (N_4419,N_2120,N_217);
nor U4420 (N_4420,N_1413,N_2448);
and U4421 (N_4421,N_2125,N_2461);
nand U4422 (N_4422,N_57,N_1543);
and U4423 (N_4423,N_2447,N_765);
xor U4424 (N_4424,N_2460,N_1021);
or U4425 (N_4425,N_913,N_2238);
nand U4426 (N_4426,N_708,N_623);
nor U4427 (N_4427,N_1487,N_797);
or U4428 (N_4428,N_610,N_1272);
nand U4429 (N_4429,N_2428,N_2227);
nor U4430 (N_4430,N_998,N_1059);
nor U4431 (N_4431,N_139,N_2051);
or U4432 (N_4432,N_1800,N_1399);
or U4433 (N_4433,N_1265,N_1789);
nand U4434 (N_4434,N_594,N_1165);
nand U4435 (N_4435,N_392,N_2381);
or U4436 (N_4436,N_2422,N_148);
nor U4437 (N_4437,N_133,N_2120);
and U4438 (N_4438,N_772,N_857);
xor U4439 (N_4439,N_2392,N_2153);
and U4440 (N_4440,N_1770,N_2089);
nand U4441 (N_4441,N_512,N_338);
nor U4442 (N_4442,N_402,N_168);
xor U4443 (N_4443,N_1447,N_439);
or U4444 (N_4444,N_684,N_2170);
nand U4445 (N_4445,N_2332,N_2171);
or U4446 (N_4446,N_1950,N_1237);
or U4447 (N_4447,N_1878,N_249);
xnor U4448 (N_4448,N_96,N_1153);
or U4449 (N_4449,N_2065,N_1503);
and U4450 (N_4450,N_2095,N_1108);
nor U4451 (N_4451,N_1075,N_1799);
xor U4452 (N_4452,N_2204,N_1245);
or U4453 (N_4453,N_1149,N_1754);
and U4454 (N_4454,N_1420,N_1687);
nor U4455 (N_4455,N_1499,N_864);
nor U4456 (N_4456,N_1184,N_1444);
nor U4457 (N_4457,N_1538,N_2358);
and U4458 (N_4458,N_2274,N_132);
nor U4459 (N_4459,N_1163,N_864);
nand U4460 (N_4460,N_2086,N_1086);
or U4461 (N_4461,N_1346,N_476);
nor U4462 (N_4462,N_2076,N_2494);
nand U4463 (N_4463,N_1672,N_2015);
xor U4464 (N_4464,N_2144,N_1307);
nand U4465 (N_4465,N_2334,N_1236);
nor U4466 (N_4466,N_2265,N_79);
and U4467 (N_4467,N_875,N_1454);
nand U4468 (N_4468,N_1570,N_965);
and U4469 (N_4469,N_729,N_2265);
nand U4470 (N_4470,N_1847,N_722);
and U4471 (N_4471,N_1323,N_1152);
or U4472 (N_4472,N_917,N_281);
nand U4473 (N_4473,N_1468,N_31);
nor U4474 (N_4474,N_1064,N_133);
nand U4475 (N_4475,N_608,N_998);
or U4476 (N_4476,N_1385,N_1098);
nor U4477 (N_4477,N_1579,N_1991);
xnor U4478 (N_4478,N_945,N_1963);
xnor U4479 (N_4479,N_2068,N_1439);
nand U4480 (N_4480,N_2386,N_1341);
or U4481 (N_4481,N_2079,N_62);
nor U4482 (N_4482,N_292,N_239);
nand U4483 (N_4483,N_1206,N_1878);
nand U4484 (N_4484,N_1061,N_997);
nor U4485 (N_4485,N_2330,N_1220);
nor U4486 (N_4486,N_1450,N_2086);
xor U4487 (N_4487,N_1726,N_1643);
xor U4488 (N_4488,N_321,N_694);
nand U4489 (N_4489,N_1131,N_457);
nand U4490 (N_4490,N_217,N_1875);
nand U4491 (N_4491,N_1769,N_2326);
nor U4492 (N_4492,N_2106,N_1663);
nand U4493 (N_4493,N_2191,N_2091);
nand U4494 (N_4494,N_1571,N_906);
xor U4495 (N_4495,N_1354,N_1870);
or U4496 (N_4496,N_1231,N_1744);
nand U4497 (N_4497,N_1940,N_2076);
nand U4498 (N_4498,N_1047,N_1606);
nor U4499 (N_4499,N_2268,N_138);
nand U4500 (N_4500,N_1766,N_504);
xor U4501 (N_4501,N_1779,N_2037);
nor U4502 (N_4502,N_181,N_784);
or U4503 (N_4503,N_887,N_2100);
nor U4504 (N_4504,N_401,N_768);
or U4505 (N_4505,N_745,N_749);
xor U4506 (N_4506,N_968,N_626);
and U4507 (N_4507,N_1326,N_621);
or U4508 (N_4508,N_2493,N_1987);
and U4509 (N_4509,N_1891,N_166);
nor U4510 (N_4510,N_472,N_700);
nor U4511 (N_4511,N_978,N_725);
or U4512 (N_4512,N_541,N_1587);
or U4513 (N_4513,N_570,N_1211);
or U4514 (N_4514,N_832,N_1427);
or U4515 (N_4515,N_2398,N_1153);
nand U4516 (N_4516,N_2216,N_1732);
and U4517 (N_4517,N_1273,N_618);
nand U4518 (N_4518,N_2383,N_1972);
and U4519 (N_4519,N_2462,N_2184);
nor U4520 (N_4520,N_2028,N_481);
nand U4521 (N_4521,N_928,N_2113);
nand U4522 (N_4522,N_904,N_2364);
or U4523 (N_4523,N_1843,N_203);
nor U4524 (N_4524,N_61,N_457);
nor U4525 (N_4525,N_535,N_1698);
or U4526 (N_4526,N_1973,N_1139);
and U4527 (N_4527,N_1093,N_2306);
nor U4528 (N_4528,N_2104,N_695);
nand U4529 (N_4529,N_805,N_574);
xor U4530 (N_4530,N_900,N_251);
or U4531 (N_4531,N_1019,N_1715);
nor U4532 (N_4532,N_1844,N_367);
and U4533 (N_4533,N_1561,N_231);
and U4534 (N_4534,N_80,N_1301);
and U4535 (N_4535,N_384,N_2037);
nor U4536 (N_4536,N_2356,N_1173);
xor U4537 (N_4537,N_1482,N_1305);
and U4538 (N_4538,N_332,N_906);
nand U4539 (N_4539,N_2149,N_1410);
xnor U4540 (N_4540,N_824,N_43);
or U4541 (N_4541,N_2377,N_2357);
and U4542 (N_4542,N_888,N_1175);
nand U4543 (N_4543,N_2446,N_2496);
nand U4544 (N_4544,N_746,N_1301);
or U4545 (N_4545,N_1916,N_138);
nand U4546 (N_4546,N_1186,N_1450);
nand U4547 (N_4547,N_320,N_768);
nor U4548 (N_4548,N_1666,N_2125);
xnor U4549 (N_4549,N_2145,N_1343);
nand U4550 (N_4550,N_749,N_1996);
and U4551 (N_4551,N_3,N_1205);
or U4552 (N_4552,N_1961,N_733);
nand U4553 (N_4553,N_262,N_2290);
xnor U4554 (N_4554,N_56,N_1729);
nor U4555 (N_4555,N_2338,N_1975);
nand U4556 (N_4556,N_118,N_271);
xor U4557 (N_4557,N_1851,N_477);
xnor U4558 (N_4558,N_1433,N_1389);
xor U4559 (N_4559,N_571,N_2089);
or U4560 (N_4560,N_942,N_1748);
xor U4561 (N_4561,N_509,N_377);
xnor U4562 (N_4562,N_914,N_29);
or U4563 (N_4563,N_208,N_629);
nand U4564 (N_4564,N_930,N_2123);
nand U4565 (N_4565,N_799,N_431);
nand U4566 (N_4566,N_196,N_1756);
or U4567 (N_4567,N_780,N_1843);
or U4568 (N_4568,N_538,N_1903);
nand U4569 (N_4569,N_1231,N_1092);
xnor U4570 (N_4570,N_138,N_1102);
or U4571 (N_4571,N_1009,N_1810);
and U4572 (N_4572,N_1472,N_2348);
and U4573 (N_4573,N_199,N_889);
or U4574 (N_4574,N_1018,N_2090);
xor U4575 (N_4575,N_85,N_938);
nor U4576 (N_4576,N_2235,N_1092);
nand U4577 (N_4577,N_626,N_611);
nand U4578 (N_4578,N_2108,N_1930);
nand U4579 (N_4579,N_2492,N_1978);
or U4580 (N_4580,N_639,N_1702);
xnor U4581 (N_4581,N_497,N_1071);
and U4582 (N_4582,N_724,N_1575);
xnor U4583 (N_4583,N_313,N_1645);
nor U4584 (N_4584,N_1762,N_2200);
nand U4585 (N_4585,N_448,N_1749);
nor U4586 (N_4586,N_1786,N_1564);
and U4587 (N_4587,N_909,N_663);
nand U4588 (N_4588,N_2325,N_882);
xnor U4589 (N_4589,N_2064,N_907);
and U4590 (N_4590,N_1342,N_1647);
or U4591 (N_4591,N_1981,N_205);
or U4592 (N_4592,N_22,N_1699);
nor U4593 (N_4593,N_345,N_1619);
and U4594 (N_4594,N_605,N_1893);
xnor U4595 (N_4595,N_1818,N_1189);
nor U4596 (N_4596,N_1133,N_1830);
nand U4597 (N_4597,N_2246,N_96);
nor U4598 (N_4598,N_2269,N_1265);
or U4599 (N_4599,N_998,N_1194);
nor U4600 (N_4600,N_112,N_1456);
nand U4601 (N_4601,N_1348,N_286);
nor U4602 (N_4602,N_724,N_890);
and U4603 (N_4603,N_1459,N_1306);
nand U4604 (N_4604,N_2114,N_2235);
or U4605 (N_4605,N_677,N_840);
xnor U4606 (N_4606,N_144,N_548);
nor U4607 (N_4607,N_2382,N_1780);
and U4608 (N_4608,N_1448,N_109);
or U4609 (N_4609,N_2325,N_2020);
nor U4610 (N_4610,N_783,N_524);
and U4611 (N_4611,N_98,N_439);
and U4612 (N_4612,N_655,N_1379);
and U4613 (N_4613,N_1860,N_1703);
xor U4614 (N_4614,N_405,N_1117);
or U4615 (N_4615,N_2381,N_1739);
and U4616 (N_4616,N_1086,N_1475);
or U4617 (N_4617,N_47,N_591);
or U4618 (N_4618,N_297,N_50);
nand U4619 (N_4619,N_579,N_1934);
nand U4620 (N_4620,N_2409,N_195);
nor U4621 (N_4621,N_79,N_1464);
or U4622 (N_4622,N_1143,N_1476);
xnor U4623 (N_4623,N_2436,N_213);
or U4624 (N_4624,N_1181,N_458);
xnor U4625 (N_4625,N_1466,N_1891);
nor U4626 (N_4626,N_2454,N_379);
or U4627 (N_4627,N_1872,N_616);
xnor U4628 (N_4628,N_159,N_941);
or U4629 (N_4629,N_958,N_107);
xnor U4630 (N_4630,N_1552,N_1926);
xnor U4631 (N_4631,N_285,N_2369);
or U4632 (N_4632,N_1701,N_1884);
or U4633 (N_4633,N_2133,N_1411);
and U4634 (N_4634,N_2171,N_1314);
and U4635 (N_4635,N_1851,N_1033);
xnor U4636 (N_4636,N_1610,N_476);
and U4637 (N_4637,N_244,N_1354);
or U4638 (N_4638,N_883,N_2262);
xnor U4639 (N_4639,N_1553,N_613);
and U4640 (N_4640,N_1985,N_521);
and U4641 (N_4641,N_1349,N_1519);
xnor U4642 (N_4642,N_1411,N_1506);
nor U4643 (N_4643,N_368,N_741);
or U4644 (N_4644,N_79,N_128);
and U4645 (N_4645,N_1181,N_216);
and U4646 (N_4646,N_2032,N_863);
nand U4647 (N_4647,N_1575,N_2078);
and U4648 (N_4648,N_1236,N_530);
nand U4649 (N_4649,N_2447,N_2449);
and U4650 (N_4650,N_1465,N_1890);
or U4651 (N_4651,N_319,N_938);
xnor U4652 (N_4652,N_2442,N_940);
and U4653 (N_4653,N_1523,N_33);
xnor U4654 (N_4654,N_168,N_965);
xor U4655 (N_4655,N_927,N_1046);
nand U4656 (N_4656,N_1374,N_2315);
or U4657 (N_4657,N_1138,N_2060);
and U4658 (N_4658,N_39,N_929);
xor U4659 (N_4659,N_1810,N_2111);
or U4660 (N_4660,N_1549,N_416);
nor U4661 (N_4661,N_1023,N_499);
nand U4662 (N_4662,N_1545,N_1753);
xor U4663 (N_4663,N_481,N_11);
xor U4664 (N_4664,N_1045,N_2302);
nor U4665 (N_4665,N_545,N_974);
nand U4666 (N_4666,N_1711,N_2049);
and U4667 (N_4667,N_1012,N_2473);
and U4668 (N_4668,N_500,N_2310);
or U4669 (N_4669,N_2227,N_1272);
or U4670 (N_4670,N_719,N_1046);
nor U4671 (N_4671,N_2121,N_1055);
and U4672 (N_4672,N_2466,N_1011);
or U4673 (N_4673,N_325,N_1390);
xor U4674 (N_4674,N_1299,N_1757);
and U4675 (N_4675,N_85,N_315);
nand U4676 (N_4676,N_166,N_1519);
and U4677 (N_4677,N_1101,N_2290);
nor U4678 (N_4678,N_798,N_400);
xor U4679 (N_4679,N_2432,N_706);
or U4680 (N_4680,N_2273,N_1135);
or U4681 (N_4681,N_2430,N_1484);
nand U4682 (N_4682,N_1683,N_1100);
or U4683 (N_4683,N_2400,N_1781);
and U4684 (N_4684,N_834,N_1827);
xor U4685 (N_4685,N_625,N_2486);
nor U4686 (N_4686,N_776,N_1491);
xnor U4687 (N_4687,N_504,N_970);
or U4688 (N_4688,N_1218,N_1626);
or U4689 (N_4689,N_1383,N_432);
xor U4690 (N_4690,N_2277,N_1210);
or U4691 (N_4691,N_612,N_582);
and U4692 (N_4692,N_810,N_1699);
and U4693 (N_4693,N_1554,N_884);
xor U4694 (N_4694,N_2206,N_583);
nand U4695 (N_4695,N_1521,N_1595);
and U4696 (N_4696,N_1386,N_887);
nor U4697 (N_4697,N_526,N_1336);
nor U4698 (N_4698,N_369,N_1839);
or U4699 (N_4699,N_1439,N_1273);
xor U4700 (N_4700,N_1466,N_1107);
xnor U4701 (N_4701,N_1110,N_698);
nand U4702 (N_4702,N_2019,N_344);
or U4703 (N_4703,N_480,N_2279);
nor U4704 (N_4704,N_2089,N_679);
xnor U4705 (N_4705,N_869,N_2019);
nor U4706 (N_4706,N_622,N_840);
and U4707 (N_4707,N_756,N_392);
and U4708 (N_4708,N_1452,N_1735);
nand U4709 (N_4709,N_1826,N_654);
or U4710 (N_4710,N_42,N_1633);
xnor U4711 (N_4711,N_70,N_2196);
xor U4712 (N_4712,N_2187,N_1812);
nand U4713 (N_4713,N_2430,N_1279);
nor U4714 (N_4714,N_44,N_2385);
nand U4715 (N_4715,N_2,N_367);
nor U4716 (N_4716,N_2396,N_1597);
or U4717 (N_4717,N_1466,N_1160);
or U4718 (N_4718,N_218,N_1457);
nor U4719 (N_4719,N_818,N_628);
and U4720 (N_4720,N_721,N_2321);
xnor U4721 (N_4721,N_2014,N_617);
or U4722 (N_4722,N_2164,N_2445);
nand U4723 (N_4723,N_2105,N_871);
nand U4724 (N_4724,N_2097,N_693);
and U4725 (N_4725,N_1357,N_1094);
nand U4726 (N_4726,N_340,N_1706);
or U4727 (N_4727,N_339,N_678);
nor U4728 (N_4728,N_1865,N_2429);
xnor U4729 (N_4729,N_1697,N_1969);
nor U4730 (N_4730,N_582,N_1513);
nand U4731 (N_4731,N_1298,N_1950);
xor U4732 (N_4732,N_1715,N_2337);
and U4733 (N_4733,N_2012,N_1746);
xnor U4734 (N_4734,N_2352,N_139);
and U4735 (N_4735,N_1085,N_2396);
or U4736 (N_4736,N_685,N_1874);
nand U4737 (N_4737,N_2285,N_33);
nand U4738 (N_4738,N_1020,N_1355);
nor U4739 (N_4739,N_602,N_701);
nor U4740 (N_4740,N_19,N_2333);
xnor U4741 (N_4741,N_1426,N_71);
nor U4742 (N_4742,N_2289,N_1182);
and U4743 (N_4743,N_2407,N_272);
xor U4744 (N_4744,N_469,N_950);
nor U4745 (N_4745,N_2342,N_695);
xnor U4746 (N_4746,N_1333,N_698);
or U4747 (N_4747,N_1412,N_728);
nand U4748 (N_4748,N_1991,N_1727);
and U4749 (N_4749,N_541,N_90);
xnor U4750 (N_4750,N_1803,N_1868);
and U4751 (N_4751,N_676,N_2461);
and U4752 (N_4752,N_1053,N_1847);
nand U4753 (N_4753,N_1047,N_1241);
or U4754 (N_4754,N_113,N_1837);
xor U4755 (N_4755,N_1706,N_1746);
or U4756 (N_4756,N_328,N_1513);
or U4757 (N_4757,N_1345,N_2401);
nand U4758 (N_4758,N_2289,N_2168);
xnor U4759 (N_4759,N_1122,N_351);
and U4760 (N_4760,N_770,N_2436);
nand U4761 (N_4761,N_1581,N_1185);
and U4762 (N_4762,N_2288,N_1913);
nand U4763 (N_4763,N_2136,N_1269);
nand U4764 (N_4764,N_658,N_1420);
xnor U4765 (N_4765,N_262,N_1369);
nor U4766 (N_4766,N_2337,N_972);
or U4767 (N_4767,N_2093,N_2096);
nand U4768 (N_4768,N_1519,N_1892);
or U4769 (N_4769,N_2308,N_1816);
and U4770 (N_4770,N_1668,N_422);
nor U4771 (N_4771,N_1232,N_1299);
and U4772 (N_4772,N_293,N_1022);
or U4773 (N_4773,N_1656,N_2342);
or U4774 (N_4774,N_515,N_268);
nor U4775 (N_4775,N_968,N_58);
nor U4776 (N_4776,N_2362,N_1892);
nor U4777 (N_4777,N_2487,N_1725);
and U4778 (N_4778,N_989,N_2368);
xor U4779 (N_4779,N_1753,N_1471);
and U4780 (N_4780,N_1506,N_579);
xnor U4781 (N_4781,N_1621,N_413);
or U4782 (N_4782,N_591,N_2218);
nor U4783 (N_4783,N_498,N_2192);
and U4784 (N_4784,N_1931,N_1474);
xor U4785 (N_4785,N_1474,N_887);
nor U4786 (N_4786,N_824,N_298);
nand U4787 (N_4787,N_2045,N_2191);
nand U4788 (N_4788,N_38,N_628);
nor U4789 (N_4789,N_2445,N_2135);
nor U4790 (N_4790,N_1056,N_1425);
nor U4791 (N_4791,N_47,N_1142);
or U4792 (N_4792,N_1037,N_647);
or U4793 (N_4793,N_1551,N_1476);
or U4794 (N_4794,N_959,N_485);
and U4795 (N_4795,N_1941,N_1455);
and U4796 (N_4796,N_2397,N_271);
and U4797 (N_4797,N_875,N_858);
and U4798 (N_4798,N_204,N_2220);
xnor U4799 (N_4799,N_913,N_1141);
nand U4800 (N_4800,N_1724,N_534);
nor U4801 (N_4801,N_1550,N_2113);
and U4802 (N_4802,N_1481,N_507);
nor U4803 (N_4803,N_1601,N_2293);
nand U4804 (N_4804,N_1896,N_744);
nand U4805 (N_4805,N_774,N_431);
nor U4806 (N_4806,N_2173,N_1543);
nor U4807 (N_4807,N_2271,N_1836);
nor U4808 (N_4808,N_1821,N_1524);
nor U4809 (N_4809,N_1106,N_1991);
or U4810 (N_4810,N_958,N_2391);
and U4811 (N_4811,N_2408,N_68);
and U4812 (N_4812,N_201,N_303);
or U4813 (N_4813,N_576,N_1628);
xor U4814 (N_4814,N_911,N_1937);
nor U4815 (N_4815,N_637,N_744);
nor U4816 (N_4816,N_2115,N_303);
nand U4817 (N_4817,N_1227,N_1622);
nand U4818 (N_4818,N_1572,N_911);
nand U4819 (N_4819,N_1249,N_176);
nor U4820 (N_4820,N_357,N_1599);
and U4821 (N_4821,N_252,N_1163);
nor U4822 (N_4822,N_238,N_1371);
or U4823 (N_4823,N_136,N_2006);
xor U4824 (N_4824,N_1124,N_2029);
nor U4825 (N_4825,N_530,N_1193);
or U4826 (N_4826,N_1806,N_2006);
xor U4827 (N_4827,N_783,N_561);
and U4828 (N_4828,N_203,N_787);
nand U4829 (N_4829,N_2341,N_1953);
nand U4830 (N_4830,N_435,N_2163);
and U4831 (N_4831,N_1934,N_1869);
and U4832 (N_4832,N_2024,N_604);
nor U4833 (N_4833,N_1273,N_146);
and U4834 (N_4834,N_719,N_2082);
nor U4835 (N_4835,N_1224,N_852);
nor U4836 (N_4836,N_113,N_1380);
xnor U4837 (N_4837,N_28,N_1090);
and U4838 (N_4838,N_564,N_2460);
xnor U4839 (N_4839,N_591,N_1266);
or U4840 (N_4840,N_1857,N_319);
nor U4841 (N_4841,N_1095,N_134);
and U4842 (N_4842,N_903,N_2093);
nor U4843 (N_4843,N_149,N_1270);
and U4844 (N_4844,N_78,N_33);
nor U4845 (N_4845,N_1541,N_372);
xor U4846 (N_4846,N_2111,N_1914);
or U4847 (N_4847,N_325,N_962);
nand U4848 (N_4848,N_466,N_1163);
nand U4849 (N_4849,N_94,N_1714);
and U4850 (N_4850,N_640,N_237);
xnor U4851 (N_4851,N_876,N_85);
nor U4852 (N_4852,N_2451,N_1258);
xor U4853 (N_4853,N_256,N_186);
or U4854 (N_4854,N_2291,N_871);
xor U4855 (N_4855,N_1329,N_561);
nor U4856 (N_4856,N_2453,N_1301);
xor U4857 (N_4857,N_339,N_1830);
xnor U4858 (N_4858,N_1503,N_1071);
and U4859 (N_4859,N_1933,N_1338);
or U4860 (N_4860,N_592,N_1240);
or U4861 (N_4861,N_2362,N_2267);
nand U4862 (N_4862,N_108,N_2185);
xor U4863 (N_4863,N_2083,N_2359);
xnor U4864 (N_4864,N_1537,N_1870);
and U4865 (N_4865,N_678,N_1378);
nor U4866 (N_4866,N_1249,N_490);
nor U4867 (N_4867,N_1295,N_1387);
xor U4868 (N_4868,N_1632,N_363);
nand U4869 (N_4869,N_2105,N_2422);
nand U4870 (N_4870,N_1931,N_2336);
or U4871 (N_4871,N_2173,N_682);
nor U4872 (N_4872,N_358,N_1316);
or U4873 (N_4873,N_365,N_867);
xor U4874 (N_4874,N_160,N_1465);
xor U4875 (N_4875,N_1599,N_464);
or U4876 (N_4876,N_1791,N_2343);
xor U4877 (N_4877,N_1599,N_942);
nor U4878 (N_4878,N_1901,N_2231);
nor U4879 (N_4879,N_121,N_1136);
nand U4880 (N_4880,N_2325,N_2075);
and U4881 (N_4881,N_2094,N_1368);
nand U4882 (N_4882,N_919,N_2011);
xnor U4883 (N_4883,N_1626,N_2224);
xnor U4884 (N_4884,N_190,N_722);
nor U4885 (N_4885,N_305,N_1932);
xnor U4886 (N_4886,N_1552,N_686);
nor U4887 (N_4887,N_1713,N_1019);
or U4888 (N_4888,N_1376,N_80);
xor U4889 (N_4889,N_1217,N_1646);
xnor U4890 (N_4890,N_1054,N_2428);
nor U4891 (N_4891,N_1222,N_2153);
xor U4892 (N_4892,N_1663,N_2123);
or U4893 (N_4893,N_189,N_1023);
nand U4894 (N_4894,N_883,N_939);
nand U4895 (N_4895,N_1091,N_2194);
xnor U4896 (N_4896,N_1891,N_396);
or U4897 (N_4897,N_2059,N_1034);
nor U4898 (N_4898,N_1325,N_1383);
and U4899 (N_4899,N_1079,N_1763);
or U4900 (N_4900,N_707,N_329);
and U4901 (N_4901,N_1000,N_85);
nand U4902 (N_4902,N_1058,N_1896);
or U4903 (N_4903,N_1108,N_367);
nand U4904 (N_4904,N_1090,N_1049);
nand U4905 (N_4905,N_385,N_1054);
xnor U4906 (N_4906,N_266,N_1348);
nand U4907 (N_4907,N_1608,N_591);
nor U4908 (N_4908,N_512,N_2441);
xor U4909 (N_4909,N_251,N_1733);
nor U4910 (N_4910,N_101,N_1981);
and U4911 (N_4911,N_442,N_1411);
or U4912 (N_4912,N_102,N_2109);
or U4913 (N_4913,N_937,N_5);
nand U4914 (N_4914,N_1608,N_178);
xor U4915 (N_4915,N_1605,N_2422);
nand U4916 (N_4916,N_1341,N_1487);
and U4917 (N_4917,N_2014,N_2112);
xnor U4918 (N_4918,N_1181,N_528);
and U4919 (N_4919,N_682,N_2038);
xnor U4920 (N_4920,N_1690,N_2427);
nor U4921 (N_4921,N_1026,N_1341);
xnor U4922 (N_4922,N_2445,N_529);
and U4923 (N_4923,N_1738,N_2475);
nor U4924 (N_4924,N_1760,N_1131);
xor U4925 (N_4925,N_977,N_639);
and U4926 (N_4926,N_1884,N_925);
nor U4927 (N_4927,N_1161,N_1305);
and U4928 (N_4928,N_1577,N_1723);
nand U4929 (N_4929,N_563,N_1486);
and U4930 (N_4930,N_879,N_1896);
nand U4931 (N_4931,N_619,N_2353);
xnor U4932 (N_4932,N_605,N_1553);
nand U4933 (N_4933,N_2241,N_839);
nand U4934 (N_4934,N_1313,N_2306);
nor U4935 (N_4935,N_326,N_1361);
xor U4936 (N_4936,N_933,N_146);
nand U4937 (N_4937,N_451,N_1172);
and U4938 (N_4938,N_1908,N_2487);
xnor U4939 (N_4939,N_1157,N_1171);
nand U4940 (N_4940,N_178,N_2171);
nor U4941 (N_4941,N_2460,N_1889);
xnor U4942 (N_4942,N_230,N_1366);
and U4943 (N_4943,N_1771,N_860);
nor U4944 (N_4944,N_2291,N_1215);
and U4945 (N_4945,N_1163,N_469);
and U4946 (N_4946,N_1988,N_728);
nor U4947 (N_4947,N_1336,N_161);
and U4948 (N_4948,N_1219,N_396);
or U4949 (N_4949,N_1211,N_2478);
and U4950 (N_4950,N_1813,N_932);
xor U4951 (N_4951,N_1243,N_411);
nand U4952 (N_4952,N_2004,N_616);
or U4953 (N_4953,N_93,N_300);
nor U4954 (N_4954,N_1594,N_2206);
nand U4955 (N_4955,N_53,N_1795);
nand U4956 (N_4956,N_2016,N_801);
or U4957 (N_4957,N_151,N_1282);
nand U4958 (N_4958,N_1816,N_706);
nor U4959 (N_4959,N_877,N_2279);
and U4960 (N_4960,N_1319,N_412);
or U4961 (N_4961,N_1307,N_54);
nand U4962 (N_4962,N_435,N_263);
and U4963 (N_4963,N_1011,N_1918);
or U4964 (N_4964,N_73,N_2055);
or U4965 (N_4965,N_1485,N_1136);
xor U4966 (N_4966,N_1229,N_1233);
or U4967 (N_4967,N_648,N_2451);
nand U4968 (N_4968,N_1540,N_385);
and U4969 (N_4969,N_395,N_1261);
nor U4970 (N_4970,N_1327,N_1927);
nand U4971 (N_4971,N_1170,N_953);
or U4972 (N_4972,N_1271,N_1801);
nand U4973 (N_4973,N_595,N_680);
nor U4974 (N_4974,N_696,N_1318);
nand U4975 (N_4975,N_820,N_191);
and U4976 (N_4976,N_1462,N_399);
or U4977 (N_4977,N_524,N_367);
or U4978 (N_4978,N_1173,N_2344);
or U4979 (N_4979,N_183,N_733);
xor U4980 (N_4980,N_411,N_2395);
and U4981 (N_4981,N_2264,N_442);
and U4982 (N_4982,N_1482,N_1761);
or U4983 (N_4983,N_1140,N_1264);
and U4984 (N_4984,N_727,N_857);
nor U4985 (N_4985,N_2384,N_1830);
nor U4986 (N_4986,N_2155,N_694);
nor U4987 (N_4987,N_1086,N_1837);
nor U4988 (N_4988,N_1211,N_2441);
or U4989 (N_4989,N_313,N_831);
and U4990 (N_4990,N_767,N_639);
nor U4991 (N_4991,N_762,N_197);
xnor U4992 (N_4992,N_1891,N_2192);
nand U4993 (N_4993,N_1049,N_865);
and U4994 (N_4994,N_1166,N_60);
nor U4995 (N_4995,N_1767,N_1682);
nor U4996 (N_4996,N_276,N_874);
and U4997 (N_4997,N_1223,N_2404);
nor U4998 (N_4998,N_777,N_708);
and U4999 (N_4999,N_1596,N_51);
and UO_0 (O_0,N_2661,N_3083);
xnor UO_1 (O_1,N_3039,N_3289);
xor UO_2 (O_2,N_4314,N_4119);
and UO_3 (O_3,N_3292,N_2519);
or UO_4 (O_4,N_2790,N_3963);
xor UO_5 (O_5,N_2810,N_3882);
xnor UO_6 (O_6,N_4598,N_3058);
and UO_7 (O_7,N_3457,N_3587);
nand UO_8 (O_8,N_4888,N_3006);
nand UO_9 (O_9,N_4565,N_4529);
and UO_10 (O_10,N_4176,N_3411);
or UO_11 (O_11,N_3051,N_3869);
or UO_12 (O_12,N_3661,N_2589);
xor UO_13 (O_13,N_3788,N_2656);
and UO_14 (O_14,N_2552,N_4449);
and UO_15 (O_15,N_3605,N_4541);
nand UO_16 (O_16,N_3619,N_4879);
nor UO_17 (O_17,N_4128,N_3603);
xor UO_18 (O_18,N_4977,N_3696);
nand UO_19 (O_19,N_2796,N_4494);
and UO_20 (O_20,N_3609,N_4150);
nand UO_21 (O_21,N_3227,N_4189);
and UO_22 (O_22,N_4732,N_4342);
and UO_23 (O_23,N_3301,N_2637);
and UO_24 (O_24,N_3482,N_2639);
and UO_25 (O_25,N_2996,N_4040);
xor UO_26 (O_26,N_2819,N_4588);
nor UO_27 (O_27,N_2666,N_4701);
and UO_28 (O_28,N_3367,N_3774);
nand UO_29 (O_29,N_2851,N_3848);
and UO_30 (O_30,N_4353,N_4792);
xor UO_31 (O_31,N_4352,N_3017);
xnor UO_32 (O_32,N_4435,N_3224);
nor UO_33 (O_33,N_2582,N_4833);
nor UO_34 (O_34,N_3918,N_3642);
or UO_35 (O_35,N_4716,N_3620);
xor UO_36 (O_36,N_3537,N_4819);
nand UO_37 (O_37,N_4566,N_4416);
and UO_38 (O_38,N_4550,N_2599);
and UO_39 (O_39,N_4910,N_2553);
xor UO_40 (O_40,N_4791,N_3937);
nand UO_41 (O_41,N_2988,N_4680);
and UO_42 (O_42,N_2610,N_3855);
xor UO_43 (O_43,N_3798,N_2713);
nor UO_44 (O_44,N_3081,N_4075);
nor UO_45 (O_45,N_3732,N_4450);
nor UO_46 (O_46,N_3193,N_3818);
nand UO_47 (O_47,N_3138,N_3186);
or UO_48 (O_48,N_4385,N_4953);
or UO_49 (O_49,N_2895,N_4948);
nor UO_50 (O_50,N_2869,N_3582);
xor UO_51 (O_51,N_4573,N_4610);
nor UO_52 (O_52,N_3852,N_3683);
xor UO_53 (O_53,N_4206,N_3729);
xor UO_54 (O_54,N_3512,N_3097);
or UO_55 (O_55,N_3335,N_4803);
and UO_56 (O_56,N_4720,N_2538);
xor UO_57 (O_57,N_4915,N_4993);
and UO_58 (O_58,N_4779,N_3448);
xnor UO_59 (O_59,N_2712,N_2648);
or UO_60 (O_60,N_3697,N_3895);
or UO_61 (O_61,N_4906,N_3205);
and UO_62 (O_62,N_4197,N_3096);
nor UO_63 (O_63,N_4646,N_2991);
xor UO_64 (O_64,N_4865,N_4989);
or UO_65 (O_65,N_3569,N_4754);
or UO_66 (O_66,N_3409,N_2572);
and UO_67 (O_67,N_3595,N_3243);
nor UO_68 (O_68,N_2687,N_3349);
nand UO_69 (O_69,N_3113,N_4714);
and UO_70 (O_70,N_4204,N_3924);
nor UO_71 (O_71,N_3256,N_3531);
xor UO_72 (O_72,N_3746,N_4907);
and UO_73 (O_73,N_3773,N_4256);
or UO_74 (O_74,N_4625,N_3681);
or UO_75 (O_75,N_3492,N_3034);
nor UO_76 (O_76,N_2510,N_4432);
nand UO_77 (O_77,N_3979,N_4210);
nand UO_78 (O_78,N_3255,N_3808);
and UO_79 (O_79,N_4127,N_4632);
nand UO_80 (O_80,N_4088,N_4447);
and UO_81 (O_81,N_3449,N_4794);
nand UO_82 (O_82,N_2885,N_3618);
nand UO_83 (O_83,N_3351,N_4032);
and UO_84 (O_84,N_3616,N_4753);
or UO_85 (O_85,N_4310,N_2919);
nor UO_86 (O_86,N_2783,N_4083);
nor UO_87 (O_87,N_4345,N_3001);
or UO_88 (O_88,N_3980,N_4011);
or UO_89 (O_89,N_4703,N_4323);
and UO_90 (O_90,N_3333,N_4905);
or UO_91 (O_91,N_3783,N_4316);
nor UO_92 (O_92,N_3897,N_4568);
and UO_93 (O_93,N_3740,N_2824);
nor UO_94 (O_94,N_4094,N_4618);
or UO_95 (O_95,N_3419,N_4721);
nor UO_96 (O_96,N_4890,N_3800);
and UO_97 (O_97,N_3178,N_2670);
and UO_98 (O_98,N_3881,N_3290);
xor UO_99 (O_99,N_3020,N_3552);
or UO_100 (O_100,N_3472,N_4657);
nor UO_101 (O_101,N_4485,N_4583);
or UO_102 (O_102,N_3817,N_2828);
and UO_103 (O_103,N_3674,N_3548);
xnor UO_104 (O_104,N_3856,N_3116);
and UO_105 (O_105,N_3180,N_2512);
or UO_106 (O_106,N_4518,N_3379);
nor UO_107 (O_107,N_3602,N_3089);
nor UO_108 (O_108,N_4304,N_4651);
or UO_109 (O_109,N_3233,N_4226);
xnor UO_110 (O_110,N_3105,N_3414);
or UO_111 (O_111,N_2836,N_3689);
or UO_112 (O_112,N_4700,N_4834);
and UO_113 (O_113,N_2794,N_4355);
and UO_114 (O_114,N_3575,N_3960);
and UO_115 (O_115,N_4969,N_2965);
xor UO_116 (O_116,N_3765,N_4245);
and UO_117 (O_117,N_3607,N_3590);
nand UO_118 (O_118,N_4913,N_3847);
nand UO_119 (O_119,N_3680,N_3720);
nor UO_120 (O_120,N_3439,N_4242);
or UO_121 (O_121,N_4381,N_4842);
nand UO_122 (O_122,N_3072,N_2916);
xor UO_123 (O_123,N_3188,N_4644);
and UO_124 (O_124,N_3842,N_3827);
nor UO_125 (O_125,N_4366,N_3543);
nand UO_126 (O_126,N_4340,N_3593);
nand UO_127 (O_127,N_2963,N_3143);
and UO_128 (O_128,N_4250,N_2501);
nor UO_129 (O_129,N_4489,N_3261);
and UO_130 (O_130,N_2746,N_4985);
or UO_131 (O_131,N_4537,N_3098);
nor UO_132 (O_132,N_2893,N_3310);
xnor UO_133 (O_133,N_3989,N_4747);
xor UO_134 (O_134,N_2909,N_3554);
and UO_135 (O_135,N_3446,N_3913);
or UO_136 (O_136,N_4483,N_3347);
nand UO_137 (O_137,N_3626,N_3781);
or UO_138 (O_138,N_4251,N_3291);
nand UO_139 (O_139,N_4538,N_3378);
nor UO_140 (O_140,N_4470,N_3421);
and UO_141 (O_141,N_4260,N_4418);
or UO_142 (O_142,N_4811,N_4881);
xor UO_143 (O_143,N_4973,N_4696);
nand UO_144 (O_144,N_3085,N_3725);
and UO_145 (O_145,N_3033,N_3723);
or UO_146 (O_146,N_4459,N_3179);
xnor UO_147 (O_147,N_3157,N_4442);
nand UO_148 (O_148,N_3153,N_4364);
nor UO_149 (O_149,N_3420,N_4394);
and UO_150 (O_150,N_3237,N_2773);
nand UO_151 (O_151,N_4990,N_3228);
or UO_152 (O_152,N_4445,N_3996);
xnor UO_153 (O_153,N_3785,N_2578);
or UO_154 (O_154,N_4288,N_3252);
nand UO_155 (O_155,N_2768,N_4182);
nand UO_156 (O_156,N_4723,N_3840);
nand UO_157 (O_157,N_3401,N_4515);
nor UO_158 (O_158,N_2915,N_3684);
or UO_159 (O_159,N_3019,N_4686);
xor UO_160 (O_160,N_3844,N_3789);
or UO_161 (O_161,N_3936,N_4956);
xor UO_162 (O_162,N_4760,N_2818);
xor UO_163 (O_163,N_3114,N_2556);
xnor UO_164 (O_164,N_3111,N_4436);
or UO_165 (O_165,N_3386,N_2874);
or UO_166 (O_166,N_3911,N_4236);
or UO_167 (O_167,N_2816,N_3796);
and UO_168 (O_168,N_3084,N_4148);
or UO_169 (O_169,N_3467,N_4994);
or UO_170 (O_170,N_3502,N_4142);
nor UO_171 (O_171,N_3209,N_3191);
nor UO_172 (O_172,N_4446,N_4372);
nand UO_173 (O_173,N_4855,N_4712);
and UO_174 (O_174,N_2653,N_4368);
or UO_175 (O_175,N_4126,N_4438);
nor UO_176 (O_176,N_2975,N_4584);
nor UO_177 (O_177,N_3435,N_4647);
nand UO_178 (O_178,N_3629,N_3653);
nand UO_179 (O_179,N_4365,N_2811);
xnor UO_180 (O_180,N_4579,N_2934);
or UO_181 (O_181,N_2698,N_3809);
or UO_182 (O_182,N_4996,N_3970);
nor UO_183 (O_183,N_3036,N_2955);
xnor UO_184 (O_184,N_4654,N_3932);
nor UO_185 (O_185,N_3520,N_3164);
nor UO_186 (O_186,N_4373,N_4074);
nand UO_187 (O_187,N_3968,N_3523);
nand UO_188 (O_188,N_4486,N_4054);
nor UO_189 (O_189,N_3717,N_4718);
xor UO_190 (O_190,N_2516,N_4234);
xor UO_191 (O_191,N_2569,N_3577);
or UO_192 (O_192,N_2647,N_3923);
and UO_193 (O_193,N_3350,N_2964);
nor UO_194 (O_194,N_2518,N_4804);
or UO_195 (O_195,N_4955,N_4444);
and UO_196 (O_196,N_3794,N_4706);
and UO_197 (O_197,N_2941,N_3461);
or UO_198 (O_198,N_2593,N_2685);
or UO_199 (O_199,N_4992,N_2673);
xor UO_200 (O_200,N_3220,N_4841);
nor UO_201 (O_201,N_2507,N_3167);
xnor UO_202 (O_202,N_3538,N_2520);
xor UO_203 (O_203,N_4897,N_2936);
nand UO_204 (O_204,N_3455,N_3204);
nor UO_205 (O_205,N_4926,N_4553);
nand UO_206 (O_206,N_3490,N_3876);
or UO_207 (O_207,N_4522,N_3055);
xnor UO_208 (O_208,N_3477,N_3257);
nor UO_209 (O_209,N_3145,N_2938);
xor UO_210 (O_210,N_3219,N_4783);
xor UO_211 (O_211,N_4419,N_4397);
nor UO_212 (O_212,N_4409,N_3806);
nor UO_213 (O_213,N_3837,N_4284);
nand UO_214 (O_214,N_2765,N_3247);
xor UO_215 (O_215,N_4200,N_4766);
or UO_216 (O_216,N_4899,N_4389);
nand UO_217 (O_217,N_3149,N_4689);
nor UO_218 (O_218,N_4534,N_2855);
and UO_219 (O_219,N_3768,N_2706);
and UO_220 (O_220,N_4983,N_4478);
nor UO_221 (O_221,N_2645,N_4324);
nor UO_222 (O_222,N_3556,N_3299);
nand UO_223 (O_223,N_2731,N_4884);
nor UO_224 (O_224,N_3162,N_3345);
or UO_225 (O_225,N_3385,N_4471);
or UO_226 (O_226,N_3088,N_3574);
nand UO_227 (O_227,N_3321,N_2676);
nand UO_228 (O_228,N_3719,N_4205);
nand UO_229 (O_229,N_4317,N_3670);
nand UO_230 (O_230,N_4767,N_4861);
or UO_231 (O_231,N_3479,N_2530);
xnor UO_232 (O_232,N_3390,N_2795);
nand UO_233 (O_233,N_3589,N_3174);
or UO_234 (O_234,N_3008,N_2503);
and UO_235 (O_235,N_4814,N_2738);
xor UO_236 (O_236,N_4768,N_4071);
nand UO_237 (O_237,N_3518,N_4569);
nand UO_238 (O_238,N_4554,N_3731);
xnor UO_239 (O_239,N_2625,N_2545);
or UO_240 (O_240,N_4179,N_4586);
xor UO_241 (O_241,N_4457,N_3921);
xor UO_242 (O_242,N_2928,N_3721);
or UO_243 (O_243,N_3061,N_4258);
and UO_244 (O_244,N_4034,N_3487);
and UO_245 (O_245,N_3845,N_2617);
and UO_246 (O_246,N_2524,N_3854);
nor UO_247 (O_247,N_4152,N_2800);
xor UO_248 (O_248,N_2740,N_2897);
xnor UO_249 (O_249,N_4958,N_2985);
xor UO_250 (O_250,N_2867,N_3319);
xor UO_251 (O_251,N_4998,N_4530);
xnor UO_252 (O_252,N_2678,N_4203);
nor UO_253 (O_253,N_3614,N_3494);
or UO_254 (O_254,N_3392,N_3142);
nand UO_255 (O_255,N_4254,N_2973);
and UO_256 (O_256,N_2506,N_3711);
nand UO_257 (O_257,N_3967,N_3596);
nand UO_258 (O_258,N_3712,N_4016);
nor UO_259 (O_259,N_3076,N_2611);
xnor UO_260 (O_260,N_3430,N_3744);
xor UO_261 (O_261,N_3649,N_4740);
xor UO_262 (O_262,N_4417,N_4558);
nand UO_263 (O_263,N_4231,N_2640);
nand UO_264 (O_264,N_3002,N_3718);
nand UO_265 (O_265,N_3892,N_4667);
xor UO_266 (O_266,N_2609,N_3830);
nor UO_267 (O_267,N_4731,N_2945);
nand UO_268 (O_268,N_4156,N_3325);
and UO_269 (O_269,N_3442,N_3190);
nand UO_270 (O_270,N_3194,N_4882);
and UO_271 (O_271,N_3894,N_4279);
or UO_272 (O_272,N_3389,N_4729);
nand UO_273 (O_273,N_4878,N_4543);
nor UO_274 (O_274,N_2918,N_4055);
and UO_275 (O_275,N_4934,N_3278);
or UO_276 (O_276,N_3786,N_3928);
nor UO_277 (O_277,N_3709,N_3973);
nand UO_278 (O_278,N_3176,N_3778);
or UO_279 (O_279,N_3956,N_3121);
and UO_280 (O_280,N_3643,N_3752);
nor UO_281 (O_281,N_4139,N_3284);
nor UO_282 (O_282,N_2724,N_2889);
xor UO_283 (O_283,N_3547,N_4954);
or UO_284 (O_284,N_3049,N_3825);
and UO_285 (O_285,N_3384,N_3545);
nor UO_286 (O_286,N_2805,N_4557);
or UO_287 (O_287,N_4357,N_4393);
and UO_288 (O_288,N_3580,N_3797);
nor UO_289 (O_289,N_3944,N_3736);
nor UO_290 (O_290,N_2758,N_3906);
nor UO_291 (O_291,N_3086,N_2891);
and UO_292 (O_292,N_4162,N_4551);
or UO_293 (O_293,N_3647,N_4079);
and UO_294 (O_294,N_4967,N_4621);
and UO_295 (O_295,N_2623,N_2717);
nor UO_296 (O_296,N_3476,N_4581);
nand UO_297 (O_297,N_3992,N_4012);
nand UO_298 (O_298,N_2958,N_2632);
or UO_299 (O_299,N_3755,N_4868);
and UO_300 (O_300,N_3371,N_2709);
xnor UO_301 (O_301,N_4964,N_2798);
or UO_302 (O_302,N_3012,N_3011);
nor UO_303 (O_303,N_3092,N_3005);
nand UO_304 (O_304,N_4512,N_4287);
and UO_305 (O_305,N_3610,N_4351);
nand UO_306 (O_306,N_4259,N_4225);
nand UO_307 (O_307,N_3429,N_4931);
xnor UO_308 (O_308,N_2887,N_3196);
xnor UO_309 (O_309,N_3016,N_4630);
nor UO_310 (O_310,N_3090,N_4105);
xor UO_311 (O_311,N_4849,N_4628);
nand UO_312 (O_312,N_3187,N_2974);
and UO_313 (O_313,N_3943,N_4736);
nand UO_314 (O_314,N_4523,N_3287);
or UO_315 (O_315,N_3685,N_3757);
xnor UO_316 (O_316,N_3735,N_2949);
or UO_317 (O_317,N_3846,N_4386);
and UO_318 (O_318,N_3669,N_2969);
or UO_319 (O_319,N_4500,N_3716);
nor UO_320 (O_320,N_3804,N_3158);
and UO_321 (O_321,N_4429,N_3331);
xnor UO_322 (O_322,N_2601,N_2779);
nor UO_323 (O_323,N_4501,N_2555);
nand UO_324 (O_324,N_2743,N_3565);
nand UO_325 (O_325,N_4671,N_3509);
nand UO_326 (O_326,N_3912,N_4475);
and UO_327 (O_327,N_2968,N_3062);
and UO_328 (O_328,N_4257,N_4609);
xor UO_329 (O_329,N_3206,N_2775);
or UO_330 (O_330,N_4413,N_3930);
nand UO_331 (O_331,N_2948,N_3166);
and UO_332 (O_332,N_2557,N_2977);
nor UO_333 (O_333,N_2606,N_3099);
xor UO_334 (O_334,N_4227,N_3819);
and UO_335 (O_335,N_2979,N_3077);
xor UO_336 (O_336,N_4218,N_3505);
xnor UO_337 (O_337,N_4867,N_2574);
xnor UO_338 (O_338,N_3137,N_4456);
or UO_339 (O_339,N_4778,N_4115);
nand UO_340 (O_340,N_3398,N_4122);
and UO_341 (O_341,N_2858,N_3622);
and UO_342 (O_342,N_3486,N_4570);
and UO_343 (O_343,N_3656,N_4895);
and UO_344 (O_344,N_2947,N_4893);
nand UO_345 (O_345,N_4864,N_4836);
or UO_346 (O_346,N_3368,N_3146);
xnor UO_347 (O_347,N_3851,N_3185);
nand UO_348 (O_348,N_2525,N_3294);
nand UO_349 (O_349,N_3489,N_4577);
xor UO_350 (O_350,N_3578,N_3666);
xor UO_351 (O_351,N_4267,N_4951);
or UO_352 (O_352,N_4422,N_3958);
and UO_353 (O_353,N_3591,N_4110);
or UO_354 (O_354,N_3300,N_4292);
and UO_355 (O_355,N_3306,N_3613);
nor UO_356 (O_356,N_2950,N_3454);
nand UO_357 (O_357,N_3483,N_4739);
xnor UO_358 (O_358,N_3480,N_4495);
nand UO_359 (O_359,N_3415,N_2707);
and UO_360 (O_360,N_3296,N_2513);
or UO_361 (O_361,N_2981,N_4045);
or UO_362 (O_362,N_3583,N_4465);
xnor UO_363 (O_363,N_4904,N_3202);
xor UO_364 (O_364,N_3491,N_3795);
xor UO_365 (O_365,N_3790,N_4578);
and UO_366 (O_366,N_2913,N_4923);
or UO_367 (O_367,N_3880,N_3198);
or UO_368 (O_368,N_4170,N_3066);
xor UO_369 (O_369,N_3983,N_4639);
nor UO_370 (O_370,N_3938,N_3812);
or UO_371 (O_371,N_3144,N_3664);
and UO_372 (O_372,N_3050,N_4361);
or UO_373 (O_373,N_3151,N_2613);
or UO_374 (O_374,N_4678,N_4187);
nand UO_375 (O_375,N_4066,N_3994);
nor UO_376 (O_376,N_4561,N_2850);
nand UO_377 (O_377,N_3816,N_2808);
or UO_378 (O_378,N_3443,N_2550);
nor UO_379 (O_379,N_4587,N_4263);
and UO_380 (O_380,N_4589,N_2932);
xnor UO_381 (O_381,N_2781,N_2523);
nand UO_382 (O_382,N_2998,N_2847);
nand UO_383 (O_383,N_3208,N_2568);
or UO_384 (O_384,N_4826,N_4880);
and UO_385 (O_385,N_2994,N_4157);
nor UO_386 (O_386,N_3743,N_3900);
xor UO_387 (O_387,N_2618,N_4608);
or UO_388 (O_388,N_4391,N_4217);
nor UO_389 (O_389,N_4668,N_3737);
xnor UO_390 (O_390,N_4688,N_3658);
and UO_391 (O_391,N_4268,N_3118);
nand UO_392 (O_392,N_4129,N_3365);
xnor UO_393 (O_393,N_2752,N_2659);
nor UO_394 (O_394,N_3754,N_2870);
nor UO_395 (O_395,N_3764,N_4002);
nand UO_396 (O_396,N_4641,N_4574);
or UO_397 (O_397,N_4190,N_4924);
nor UO_398 (O_398,N_3883,N_3772);
nor UO_399 (O_399,N_3399,N_2922);
nor UO_400 (O_400,N_2638,N_4594);
or UO_401 (O_401,N_4591,N_4592);
or UO_402 (O_402,N_4330,N_3517);
and UO_403 (O_403,N_3148,N_2835);
and UO_404 (O_404,N_2672,N_2879);
xor UO_405 (O_405,N_3372,N_4533);
and UO_406 (O_406,N_4235,N_4697);
or UO_407 (O_407,N_2652,N_2682);
nand UO_408 (O_408,N_3369,N_4564);
and UO_409 (O_409,N_3776,N_4582);
xor UO_410 (O_410,N_3117,N_2799);
nor UO_411 (O_411,N_3436,N_3941);
and UO_412 (O_412,N_4874,N_2900);
or UO_413 (O_413,N_3561,N_2972);
or UO_414 (O_414,N_3695,N_4172);
nor UO_415 (O_415,N_3288,N_3802);
nor UO_416 (O_416,N_2786,N_4358);
and UO_417 (O_417,N_2697,N_2925);
and UO_418 (O_418,N_3057,N_3317);
xor UO_419 (O_419,N_4575,N_4102);
xor UO_420 (O_420,N_4517,N_2767);
nand UO_421 (O_421,N_3380,N_4061);
and UO_422 (O_422,N_3009,N_4627);
and UO_423 (O_423,N_3307,N_3318);
and UO_424 (O_424,N_4036,N_3363);
xor UO_425 (O_425,N_4338,N_2787);
nand UO_426 (O_426,N_4859,N_3075);
xnor UO_427 (O_427,N_3805,N_3728);
nor UO_428 (O_428,N_4252,N_4726);
or UO_429 (O_429,N_2865,N_4866);
and UO_430 (O_430,N_2636,N_4007);
and UO_431 (O_431,N_4093,N_4971);
or UO_432 (O_432,N_2514,N_3074);
and UO_433 (O_433,N_4237,N_3242);
nor UO_434 (O_434,N_3976,N_3354);
and UO_435 (O_435,N_4972,N_3692);
and UO_436 (O_436,N_2526,N_4759);
nor UO_437 (O_437,N_3070,N_2631);
or UO_438 (O_438,N_2654,N_4427);
nor UO_439 (O_439,N_2860,N_3893);
nor UO_440 (O_440,N_2999,N_4828);
nor UO_441 (O_441,N_3947,N_2849);
xnor UO_442 (O_442,N_3431,N_4406);
nor UO_443 (O_443,N_3239,N_3165);
and UO_444 (O_444,N_3110,N_3232);
nand UO_445 (O_445,N_3460,N_4889);
and UO_446 (O_446,N_4600,N_3832);
or UO_447 (O_447,N_2701,N_2954);
nor UO_448 (O_448,N_3340,N_2992);
or UO_449 (O_449,N_4398,N_2957);
and UO_450 (O_450,N_4733,N_3763);
nand UO_451 (O_451,N_4692,N_4167);
and UO_452 (O_452,N_4151,N_4109);
nor UO_453 (O_453,N_2543,N_3885);
nand UO_454 (O_454,N_2621,N_2962);
or UO_455 (O_455,N_3469,N_3260);
and UO_456 (O_456,N_3549,N_2732);
or UO_457 (O_457,N_4937,N_4261);
or UO_458 (O_458,N_4943,N_4536);
and UO_459 (O_459,N_3200,N_3192);
and UO_460 (O_460,N_4270,N_2995);
nand UO_461 (O_461,N_3238,N_4396);
and UO_462 (O_462,N_3129,N_4827);
xnor UO_463 (O_463,N_4433,N_2720);
and UO_464 (O_464,N_3964,N_2664);
or UO_465 (O_465,N_3571,N_2739);
nor UO_466 (O_466,N_4140,N_4425);
nor UO_467 (O_467,N_2583,N_2726);
nor UO_468 (O_468,N_4762,N_2980);
and UO_469 (O_469,N_3128,N_3463);
xnor UO_470 (O_470,N_2921,N_4482);
or UO_471 (O_471,N_4607,N_3510);
nor UO_472 (O_472,N_3559,N_3986);
xnor UO_473 (O_473,N_4511,N_3507);
and UO_474 (O_474,N_3673,N_4559);
or UO_475 (O_475,N_2956,N_2785);
xnor UO_476 (O_476,N_4820,N_3687);
and UO_477 (O_477,N_4307,N_4801);
nor UO_478 (O_478,N_2878,N_3360);
and UO_479 (O_479,N_3741,N_4793);
xnor UO_480 (O_480,N_4929,N_3172);
or UO_481 (O_481,N_4325,N_4289);
or UO_482 (O_482,N_3199,N_3550);
nand UO_483 (O_483,N_3645,N_3624);
or UO_484 (O_484,N_3078,N_2690);
nand UO_485 (O_485,N_2716,N_4576);
and UO_486 (O_486,N_3346,N_2990);
xor UO_487 (O_487,N_4230,N_3657);
xor UO_488 (O_488,N_2953,N_4655);
nand UO_489 (O_489,N_4719,N_4118);
nor UO_490 (O_490,N_3177,N_3857);
and UO_491 (O_491,N_3955,N_3903);
or UO_492 (O_492,N_3171,N_3230);
nor UO_493 (O_493,N_3516,N_2699);
xnor UO_494 (O_494,N_3271,N_2662);
nor UO_495 (O_495,N_4914,N_4091);
or UO_496 (O_496,N_3201,N_3498);
or UO_497 (O_497,N_3328,N_3387);
nand UO_498 (O_498,N_4077,N_4665);
nor UO_499 (O_499,N_2852,N_3586);
nor UO_500 (O_500,N_3829,N_4332);
nor UO_501 (O_501,N_4752,N_4854);
nor UO_502 (O_502,N_4184,N_2563);
nor UO_503 (O_503,N_4303,N_3959);
nand UO_504 (O_504,N_4620,N_3285);
nand UO_505 (O_505,N_2854,N_3513);
or UO_506 (O_506,N_3023,N_3014);
or UO_507 (O_507,N_3573,N_4451);
and UO_508 (O_508,N_3849,N_3330);
nor UO_509 (O_509,N_4089,N_2559);
xnor UO_510 (O_510,N_3048,N_4524);
or UO_511 (O_511,N_2838,N_4602);
xnor UO_512 (O_512,N_3592,N_2571);
and UO_513 (O_513,N_2663,N_4212);
nand UO_514 (O_514,N_4050,N_4840);
xnor UO_515 (O_515,N_2848,N_3183);
and UO_516 (O_516,N_4690,N_3108);
and UO_517 (O_517,N_2937,N_4318);
xor UO_518 (O_518,N_3470,N_3969);
or UO_519 (O_519,N_2959,N_3742);
and UO_520 (O_520,N_3107,N_4022);
nand UO_521 (O_521,N_4707,N_3276);
or UO_522 (O_522,N_2580,N_4010);
nand UO_523 (O_523,N_4362,N_4320);
or UO_524 (O_524,N_2817,N_2677);
and UO_525 (O_525,N_4896,N_3364);
xnor UO_526 (O_526,N_3791,N_2750);
xor UO_527 (O_527,N_4460,N_3320);
and UO_528 (O_528,N_3888,N_4945);
nor UO_529 (O_529,N_2939,N_4756);
and UO_530 (O_530,N_4069,N_4892);
nand UO_531 (O_531,N_4711,N_4240);
and UO_532 (O_532,N_3007,N_3053);
nor UO_533 (O_533,N_2527,N_2834);
or UO_534 (O_534,N_3221,N_2757);
and UO_535 (O_535,N_3308,N_2595);
or UO_536 (O_536,N_4528,N_2721);
and UO_537 (O_537,N_2634,N_4546);
xor UO_538 (O_538,N_3635,N_4812);
nor UO_539 (O_539,N_2821,N_3710);
or UO_540 (O_540,N_2789,N_3867);
or UO_541 (O_541,N_3056,N_4277);
xnor UO_542 (O_542,N_3311,N_2607);
nor UO_543 (O_543,N_4132,N_4214);
nor UO_544 (O_544,N_4497,N_4961);
and UO_545 (O_545,N_4137,N_3223);
nor UO_546 (O_546,N_4000,N_4311);
xnor UO_547 (O_547,N_3997,N_2679);
and UO_548 (O_548,N_2807,N_2539);
nor UO_549 (O_549,N_3822,N_2628);
nand UO_550 (O_550,N_4782,N_3405);
nand UO_551 (O_551,N_4285,N_4835);
and UO_552 (O_552,N_4815,N_2931);
nor UO_553 (O_553,N_3756,N_2771);
xor UO_554 (O_554,N_4341,N_4120);
xor UO_555 (O_555,N_3691,N_4932);
xnor UO_556 (O_556,N_4173,N_3456);
and UO_557 (O_557,N_4476,N_4213);
nand UO_558 (O_558,N_3704,N_2788);
or UO_559 (O_559,N_3803,N_3464);
nand UO_560 (O_560,N_4377,N_2903);
xnor UO_561 (O_561,N_2696,N_2753);
nand UO_562 (O_562,N_4514,N_3500);
xor UO_563 (O_563,N_3722,N_4410);
and UO_564 (O_564,N_4033,N_3901);
nor UO_565 (O_565,N_4999,N_2881);
nand UO_566 (O_566,N_3748,N_3584);
xor UO_567 (O_567,N_3700,N_4356);
nand UO_568 (O_568,N_3274,N_4072);
nand UO_569 (O_569,N_2734,N_4013);
xor UO_570 (O_570,N_4917,N_3211);
nand UO_571 (O_571,N_3356,N_2910);
nor UO_572 (O_572,N_2646,N_2935);
xor UO_573 (O_573,N_2509,N_4400);
and UO_574 (O_574,N_2777,N_4950);
nor UO_575 (O_575,N_4661,N_3156);
xnor UO_576 (O_576,N_3326,N_3904);
nor UO_577 (O_577,N_4774,N_4635);
nand UO_578 (O_578,N_4664,N_3222);
nand UO_579 (O_579,N_4965,N_3799);
and UO_580 (O_580,N_4503,N_4253);
nand UO_581 (O_581,N_2533,N_2886);
nand UO_582 (O_582,N_3949,N_4019);
nand UO_583 (O_583,N_3091,N_3004);
and UO_584 (O_584,N_2551,N_2896);
and UO_585 (O_585,N_4367,N_2564);
and UO_586 (O_586,N_4308,N_3546);
nor UO_587 (O_587,N_3381,N_4291);
nor UO_588 (O_588,N_4051,N_3359);
or UO_589 (O_589,N_3361,N_4669);
xnor UO_590 (O_590,N_4281,N_4496);
and UO_591 (O_591,N_4085,N_4161);
or UO_592 (O_592,N_4046,N_4111);
nand UO_593 (O_593,N_3212,N_4595);
nand UO_594 (O_594,N_4818,N_4220);
xnor UO_595 (O_595,N_4155,N_3676);
xor UO_596 (O_596,N_3659,N_3747);
or UO_597 (O_597,N_3226,N_3762);
nor UO_598 (O_598,N_3951,N_3690);
xnor UO_599 (O_599,N_3024,N_3101);
or UO_600 (O_600,N_3283,N_4070);
nor UO_601 (O_601,N_4666,N_3323);
or UO_602 (O_602,N_4100,N_4329);
nand UO_603 (O_603,N_4611,N_4663);
and UO_604 (O_604,N_2641,N_4775);
or UO_605 (O_605,N_3154,N_4599);
nor UO_606 (O_606,N_3539,N_3298);
or UO_607 (O_607,N_4949,N_4624);
nor UO_608 (O_608,N_3898,N_3132);
or UO_609 (O_609,N_4322,N_4704);
nand UO_610 (O_610,N_2882,N_4057);
nor UO_611 (O_611,N_4959,N_2813);
xnor UO_612 (O_612,N_4542,N_4921);
or UO_613 (O_613,N_3216,N_3042);
xnor UO_614 (O_614,N_2714,N_4851);
and UO_615 (O_615,N_3450,N_4087);
nor UO_616 (O_616,N_3896,N_4614);
xnor UO_617 (O_617,N_4283,N_4420);
and UO_618 (O_618,N_4772,N_3770);
and UO_619 (O_619,N_3879,N_2548);
and UO_620 (O_620,N_3961,N_4472);
or UO_621 (O_621,N_3229,N_2871);
nand UO_622 (O_622,N_3655,N_4059);
and UO_623 (O_623,N_4947,N_4545);
or UO_624 (O_624,N_2686,N_2642);
nand UO_625 (O_625,N_2633,N_3775);
and UO_626 (O_626,N_4987,N_3425);
nor UO_627 (O_627,N_4789,N_2888);
or UO_628 (O_628,N_2902,N_4604);
nand UO_629 (O_629,N_3396,N_3267);
nor UO_630 (O_630,N_3920,N_3312);
nand UO_631 (O_631,N_4491,N_4481);
and UO_632 (O_632,N_3236,N_3828);
and UO_633 (O_633,N_4428,N_4728);
or UO_634 (O_634,N_4821,N_3280);
nor UO_635 (O_635,N_4749,N_4028);
nand UO_636 (O_636,N_4873,N_4957);
nor UO_637 (O_637,N_3484,N_3751);
and UO_638 (O_638,N_3241,N_3698);
and UO_639 (O_639,N_2923,N_2797);
nand UO_640 (O_640,N_4832,N_3270);
and UO_641 (O_641,N_3750,N_3391);
nand UO_642 (O_642,N_3068,N_2820);
or UO_643 (O_643,N_4488,N_4679);
and UO_644 (O_644,N_4634,N_4813);
xnor UO_645 (O_645,N_3811,N_3052);
nand UO_646 (O_646,N_2675,N_3831);
and UO_647 (O_647,N_4619,N_2872);
and UO_648 (O_648,N_4183,N_3305);
nor UO_649 (O_649,N_3393,N_4670);
nor UO_650 (O_650,N_3993,N_4388);
and UO_651 (O_651,N_4572,N_4968);
or UO_652 (O_652,N_3273,N_3063);
or UO_653 (O_653,N_4622,N_3625);
and UO_654 (O_654,N_3136,N_3250);
or UO_655 (O_655,N_4001,N_2742);
or UO_656 (O_656,N_4437,N_4424);
xnor UO_657 (O_657,N_4970,N_2608);
or UO_658 (O_658,N_2584,N_4326);
nand UO_659 (O_659,N_4163,N_4453);
nor UO_660 (O_660,N_2930,N_4927);
xnor UO_661 (O_661,N_4264,N_3217);
nand UO_662 (O_662,N_3975,N_3563);
and UO_663 (O_663,N_4976,N_4562);
or UO_664 (O_664,N_3604,N_3473);
or UO_665 (O_665,N_4241,N_3688);
or UO_666 (O_666,N_4131,N_2718);
or UO_667 (O_667,N_4900,N_3868);
nand UO_668 (O_668,N_4201,N_2831);
and UO_669 (O_669,N_4675,N_3244);
nand UO_670 (O_670,N_3135,N_4822);
and UO_671 (O_671,N_3675,N_3041);
or UO_672 (O_672,N_4346,N_4215);
and UO_673 (O_673,N_3102,N_4383);
nand UO_674 (O_674,N_4008,N_3823);
and UO_675 (O_675,N_3872,N_3060);
nand UO_676 (O_676,N_4677,N_2535);
nand UO_677 (O_677,N_4629,N_4194);
or UO_678 (O_678,N_4660,N_3962);
or UO_679 (O_679,N_4023,N_4166);
xor UO_680 (O_680,N_3702,N_3514);
xor UO_681 (O_681,N_3214,N_3598);
nor UO_682 (O_682,N_4363,N_3329);
xor UO_683 (O_683,N_2924,N_2665);
nand UO_684 (O_684,N_3293,N_4443);
or UO_685 (O_685,N_3861,N_4068);
nor UO_686 (O_686,N_2832,N_4191);
or UO_687 (O_687,N_4029,N_3891);
or UO_688 (O_688,N_3352,N_4164);
or UO_689 (O_689,N_2573,N_3521);
or UO_690 (O_690,N_4858,N_3030);
nor UO_691 (O_691,N_3501,N_4009);
or UO_692 (O_692,N_4887,N_3769);
xor UO_693 (O_693,N_4223,N_4052);
nor UO_694 (O_694,N_4415,N_4255);
xor UO_695 (O_695,N_4507,N_3761);
xor UO_696 (O_696,N_2976,N_3071);
nor UO_697 (O_697,N_4612,N_3376);
xnor UO_698 (O_698,N_2766,N_3141);
nor UO_699 (O_699,N_4563,N_3734);
xnor UO_700 (O_700,N_4493,N_2692);
nand UO_701 (O_701,N_4464,N_4335);
nand UO_702 (O_702,N_3677,N_3416);
nand UO_703 (O_703,N_3662,N_4035);
or UO_704 (O_704,N_3047,N_4454);
and UO_705 (O_705,N_3021,N_4379);
and UO_706 (O_706,N_2700,N_3639);
or UO_707 (O_707,N_3403,N_3003);
or UO_708 (O_708,N_4238,N_2971);
and UO_709 (O_709,N_4986,N_2688);
xor UO_710 (O_710,N_3124,N_2596);
or UO_711 (O_711,N_4065,N_4044);
xnor UO_712 (O_712,N_2864,N_3406);
nor UO_713 (O_713,N_3915,N_3173);
xnor UO_714 (O_714,N_4101,N_4018);
nand UO_715 (O_715,N_2829,N_3466);
or UO_716 (O_716,N_2579,N_4147);
nor UO_717 (O_717,N_3564,N_2592);
or UO_718 (O_718,N_2776,N_4159);
xnor UO_719 (O_719,N_3475,N_4154);
or UO_720 (O_720,N_4784,N_3235);
nand UO_721 (O_721,N_2674,N_4169);
and UO_722 (O_722,N_3758,N_4402);
and UO_723 (O_723,N_4601,N_4799);
nor UO_724 (O_724,N_3109,N_2904);
and UO_725 (O_725,N_3324,N_4871);
nor UO_726 (O_726,N_2911,N_3082);
and UO_727 (O_727,N_4468,N_3665);
and UO_728 (O_728,N_3585,N_3899);
and UO_729 (O_729,N_4672,N_3945);
or UO_730 (O_730,N_3946,N_3459);
or UO_731 (O_731,N_4359,N_2542);
nand UO_732 (O_732,N_2784,N_2515);
and UO_733 (O_733,N_3939,N_4708);
nand UO_734 (O_734,N_3568,N_2612);
nand UO_735 (O_735,N_4441,N_2927);
nand UO_736 (O_736,N_2711,N_4585);
and UO_737 (O_737,N_2791,N_2500);
and UO_738 (O_738,N_3370,N_3161);
xnor UO_739 (O_739,N_4757,N_2782);
xor UO_740 (O_740,N_3977,N_3838);
and UO_741 (O_741,N_4698,N_4788);
xnor UO_742 (O_742,N_4966,N_4911);
xor UO_743 (O_743,N_4636,N_2733);
nand UO_744 (O_744,N_4930,N_4180);
xnor UO_745 (O_745,N_3515,N_4458);
or UO_746 (O_746,N_3015,N_4502);
and UO_747 (O_747,N_3046,N_3984);
and UO_748 (O_748,N_4039,N_4722);
xnor UO_749 (O_749,N_4003,N_4290);
nand UO_750 (O_750,N_4336,N_4695);
and UO_751 (O_751,N_3606,N_3724);
and UO_752 (O_752,N_3175,N_3029);
or UO_753 (O_753,N_4378,N_4090);
nor UO_754 (O_754,N_4080,N_4421);
nor UO_755 (O_755,N_3972,N_3423);
and UO_756 (O_756,N_3982,N_3316);
nor UO_757 (O_757,N_4198,N_3428);
or UO_758 (O_758,N_2806,N_3553);
nor UO_759 (O_759,N_3843,N_4952);
nand UO_760 (O_760,N_4499,N_4021);
xnor UO_761 (O_761,N_4440,N_3395);
xnor UO_762 (O_762,N_4894,N_4875);
xor UO_763 (O_763,N_4181,N_3544);
nand UO_764 (O_764,N_4505,N_2993);
and UO_765 (O_765,N_3889,N_4248);
xor UO_766 (O_766,N_4058,N_3506);
xnor UO_767 (O_767,N_3377,N_2997);
nor UO_768 (O_768,N_3859,N_3634);
xor UO_769 (O_769,N_3203,N_3862);
nand UO_770 (O_770,N_4498,N_3820);
or UO_771 (O_771,N_4078,N_3714);
and UO_772 (O_772,N_3441,N_4596);
or UO_773 (O_773,N_4207,N_3471);
xor UO_774 (O_774,N_2770,N_2744);
nor UO_775 (O_775,N_3630,N_2540);
xor UO_776 (O_776,N_2914,N_3706);
nand UO_777 (O_777,N_3253,N_2730);
nand UO_778 (O_778,N_3120,N_3726);
nor UO_779 (O_779,N_4755,N_3181);
nor UO_780 (O_780,N_3934,N_4684);
nor UO_781 (O_781,N_2616,N_3131);
xor UO_782 (O_782,N_2737,N_3999);
nand UO_783 (O_783,N_3652,N_4928);
and UO_784 (O_784,N_3334,N_4870);
or UO_785 (O_785,N_4298,N_2566);
and UO_786 (O_786,N_4158,N_3474);
nand UO_787 (O_787,N_4580,N_4047);
xnor UO_788 (O_788,N_4650,N_3468);
nor UO_789 (O_789,N_4623,N_3648);
nand UO_790 (O_790,N_4177,N_4605);
nor UO_791 (O_791,N_4848,N_4144);
xor UO_792 (O_792,N_4942,N_2883);
nand UO_793 (O_793,N_3453,N_3488);
nand UO_794 (O_794,N_4275,N_3810);
nand UO_795 (O_795,N_3908,N_3650);
nand UO_796 (O_796,N_4901,N_3245);
xor UO_797 (O_797,N_3974,N_4532);
or UO_798 (O_798,N_2905,N_2780);
and UO_799 (O_799,N_2560,N_4233);
and UO_800 (O_800,N_4412,N_3821);
nor UO_801 (O_801,N_3705,N_3358);
nand UO_802 (O_802,N_2587,N_3954);
nand UO_803 (O_803,N_2970,N_4192);
xnor UO_804 (O_804,N_2920,N_2830);
and UO_805 (O_805,N_2759,N_4042);
nand UO_806 (O_806,N_3493,N_4922);
or UO_807 (O_807,N_2570,N_3437);
nor UO_808 (O_808,N_4786,N_3877);
xor UO_809 (O_809,N_4174,N_4295);
or UO_810 (O_810,N_3106,N_4171);
and UO_811 (O_811,N_4390,N_2622);
nor UO_812 (O_812,N_4737,N_4467);
xnor UO_813 (O_813,N_3160,N_4455);
and UO_814 (O_814,N_4658,N_2626);
and UO_815 (O_815,N_3433,N_2650);
and UO_816 (O_816,N_4758,N_4806);
and UO_817 (O_817,N_4860,N_4448);
xnor UO_818 (O_818,N_2763,N_4903);
or UO_819 (O_819,N_2747,N_3248);
or UO_820 (O_820,N_3807,N_2531);
and UO_821 (O_821,N_3981,N_4399);
nand UO_822 (O_822,N_2705,N_4853);
or UO_823 (O_823,N_4380,N_3037);
nand UO_824 (O_824,N_4274,N_4790);
nand UO_825 (O_825,N_2899,N_4995);
xor UO_826 (O_826,N_4908,N_4243);
and UO_827 (O_827,N_4062,N_4617);
xor UO_828 (O_828,N_3841,N_4991);
xor UO_829 (O_829,N_3315,N_2541);
or UO_830 (O_830,N_3440,N_4219);
xnor UO_831 (O_831,N_4312,N_3348);
or UO_832 (O_832,N_4730,N_3555);
or UO_833 (O_833,N_2801,N_4037);
and UO_834 (O_834,N_4474,N_4229);
nor UO_835 (O_835,N_4123,N_3528);
and UO_836 (O_836,N_2986,N_3987);
and UO_837 (O_837,N_4548,N_2857);
nand UO_838 (O_838,N_3953,N_2748);
nor UO_839 (O_839,N_4117,N_2989);
nand UO_840 (O_840,N_3112,N_4247);
or UO_841 (O_841,N_4809,N_3452);
nor UO_842 (O_842,N_4988,N_4125);
and UO_843 (O_843,N_4348,N_4824);
nand UO_844 (O_844,N_2942,N_2567);
or UO_845 (O_845,N_4103,N_3225);
or UO_846 (O_846,N_3122,N_2529);
xor UO_847 (O_847,N_4702,N_2839);
or UO_848 (O_848,N_2756,N_4466);
xnor UO_849 (O_849,N_4136,N_2982);
and UO_850 (O_850,N_3266,N_3169);
and UO_851 (O_851,N_4593,N_3874);
xor UO_852 (O_852,N_3104,N_4862);
xnor UO_853 (O_853,N_3998,N_3535);
or UO_854 (O_854,N_4852,N_3632);
or UO_855 (O_855,N_4411,N_3027);
nor UO_856 (O_856,N_4606,N_3766);
nor UO_857 (O_857,N_4735,N_4642);
nand UO_858 (O_858,N_3309,N_4912);
nand UO_859 (O_859,N_4020,N_4802);
nand UO_860 (O_860,N_3263,N_3297);
nand UO_861 (O_861,N_2926,N_4211);
nand UO_862 (O_862,N_3115,N_4863);
xnor UO_863 (O_863,N_2693,N_4780);
nand UO_864 (O_864,N_2933,N_4302);
xor UO_865 (O_865,N_3638,N_2549);
or UO_866 (O_866,N_3519,N_3524);
or UO_867 (O_867,N_3644,N_4556);
and UO_868 (O_868,N_3139,N_4939);
or UO_869 (O_869,N_4713,N_2859);
xnor UO_870 (O_870,N_3054,N_3397);
nor UO_871 (O_871,N_4143,N_2505);
nand UO_872 (O_872,N_3277,N_3357);
nor UO_873 (O_873,N_4084,N_3990);
and UO_874 (O_874,N_4800,N_4178);
nor UO_875 (O_875,N_4492,N_4186);
nand UO_876 (O_876,N_4590,N_4745);
or UO_877 (O_877,N_4404,N_2695);
nand UO_878 (O_878,N_4513,N_3065);
nor UO_879 (O_879,N_4662,N_2681);
and UO_880 (O_880,N_3079,N_2598);
xnor UO_881 (O_881,N_3417,N_3814);
nand UO_882 (O_882,N_3628,N_2876);
or UO_883 (O_883,N_2803,N_2534);
xnor UO_884 (O_884,N_3251,N_4960);
nor UO_885 (O_885,N_4891,N_4519);
nand UO_886 (O_886,N_4280,N_3713);
nor UO_887 (O_887,N_3022,N_4909);
nor UO_888 (O_888,N_2814,N_3753);
xnor UO_889 (O_889,N_3532,N_4276);
nand UO_890 (O_890,N_3836,N_4877);
xnor UO_891 (O_891,N_3760,N_3957);
nor UO_892 (O_892,N_4313,N_3579);
xor UO_893 (O_893,N_4249,N_2668);
or UO_894 (O_894,N_2689,N_4487);
and UO_895 (O_895,N_3265,N_3667);
xnor UO_896 (O_896,N_4145,N_3668);
or UO_897 (O_897,N_3916,N_4555);
nand UO_898 (O_898,N_3269,N_3100);
nand UO_899 (O_899,N_4371,N_3093);
or UO_900 (O_900,N_3195,N_3551);
or UO_901 (O_901,N_3503,N_4776);
nand UO_902 (O_902,N_4053,N_2863);
xor UO_903 (O_903,N_4825,N_4025);
nor UO_904 (O_904,N_3432,N_4076);
and UO_905 (O_905,N_3402,N_4005);
and UO_906 (O_906,N_2727,N_3032);
or UO_907 (O_907,N_3426,N_4334);
xnor UO_908 (O_908,N_4659,N_4299);
nand UO_909 (O_909,N_2906,N_4805);
or UO_910 (O_910,N_2966,N_4944);
xor UO_911 (O_911,N_4876,N_4333);
nand UO_912 (O_912,N_3388,N_4095);
nand UO_913 (O_913,N_4188,N_4104);
xor UO_914 (O_914,N_3366,N_2722);
xnor UO_915 (O_915,N_4857,N_3525);
and UO_916 (O_916,N_4461,N_4269);
or UO_917 (O_917,N_2754,N_3597);
nor UO_918 (O_918,N_3600,N_2792);
nor UO_919 (O_919,N_4656,N_4221);
and UO_920 (O_920,N_2736,N_3373);
nand UO_921 (O_921,N_3914,N_3701);
nand UO_922 (O_922,N_4360,N_2762);
nand UO_923 (O_923,N_4771,N_4531);
or UO_924 (O_924,N_3069,N_2708);
nor UO_925 (O_925,N_2772,N_2802);
nand UO_926 (O_926,N_3304,N_2875);
and UO_927 (O_927,N_3787,N_2826);
nor UO_928 (O_928,N_4405,N_4408);
nor UO_929 (O_929,N_4770,N_4847);
or UO_930 (O_930,N_3413,N_4473);
nand UO_931 (O_931,N_2644,N_3824);
or UO_932 (O_932,N_4808,N_3865);
nand UO_933 (O_933,N_3240,N_4709);
xnor UO_934 (O_934,N_2655,N_4506);
or UO_935 (O_935,N_4734,N_3878);
or UO_936 (O_936,N_2725,N_3866);
and UO_937 (O_937,N_3611,N_4724);
and UO_938 (O_938,N_4354,N_4845);
and UO_939 (O_939,N_4777,N_2845);
or UO_940 (O_940,N_4781,N_3526);
and UO_941 (O_941,N_2600,N_3601);
nand UO_942 (O_942,N_4773,N_4640);
or UO_943 (O_943,N_3013,N_4185);
or UO_944 (O_944,N_4124,N_3749);
and UO_945 (O_945,N_3094,N_4113);
nand UO_946 (O_946,N_3511,N_4426);
nand UO_947 (O_947,N_4938,N_3534);
nand UO_948 (O_948,N_2629,N_2627);
nand UO_949 (O_949,N_3362,N_3234);
nor UO_950 (O_950,N_4431,N_2760);
nor UO_951 (O_951,N_2907,N_3327);
nor UO_952 (O_952,N_2929,N_4463);
nor UO_953 (O_953,N_4133,N_3458);
nand UO_954 (O_954,N_3884,N_4434);
nor UO_955 (O_955,N_3103,N_3424);
or UO_956 (O_956,N_4510,N_2669);
xnor UO_957 (O_957,N_4715,N_3952);
and UO_958 (O_958,N_2898,N_4107);
nor UO_959 (O_959,N_3264,N_4725);
xnor UO_960 (O_960,N_4535,N_4979);
nand UO_961 (O_961,N_4567,N_3445);
or UO_962 (O_962,N_4975,N_2908);
and UO_963 (O_963,N_3739,N_4795);
xor UO_964 (O_964,N_3213,N_4319);
xnor UO_965 (O_965,N_2880,N_4328);
or UO_966 (O_966,N_3119,N_2840);
or UO_967 (O_967,N_3672,N_4096);
nor UO_968 (O_968,N_3504,N_3168);
nand UO_969 (O_969,N_4649,N_4370);
and UO_970 (O_970,N_3621,N_2546);
or UO_971 (O_971,N_3018,N_3529);
nand UO_972 (O_972,N_3182,N_3890);
or UO_973 (O_973,N_3654,N_4395);
nor UO_974 (O_974,N_2522,N_2809);
or UO_975 (O_975,N_4652,N_3887);
nand UO_976 (O_976,N_2619,N_3909);
nand UO_977 (O_977,N_3258,N_3703);
or UO_978 (O_978,N_3496,N_4222);
or UO_979 (O_979,N_3302,N_4414);
or UO_980 (O_980,N_2769,N_3000);
nand UO_981 (O_981,N_3780,N_4974);
or UO_982 (O_982,N_3010,N_2657);
nand UO_983 (O_983,N_4138,N_4015);
and UO_984 (O_984,N_3858,N_3834);
xnor UO_985 (O_985,N_3540,N_2635);
and UO_986 (O_986,N_3408,N_4508);
nor UO_987 (O_987,N_3338,N_3332);
xor UO_988 (O_988,N_4919,N_4097);
and UO_989 (O_989,N_3218,N_3875);
or UO_990 (O_990,N_4106,N_4705);
xor UO_991 (O_991,N_4430,N_3147);
xnor UO_992 (O_992,N_3268,N_3599);
nor UO_993 (O_993,N_4484,N_3530);
and UO_994 (O_994,N_3163,N_4480);
nand UO_995 (O_995,N_3447,N_4691);
or UO_996 (O_996,N_2561,N_4327);
nand UO_997 (O_997,N_3189,N_4693);
nor UO_998 (O_998,N_3907,N_4933);
nand UO_999 (O_999,N_3641,N_4631);
endmodule