module basic_1000_10000_1500_4_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_972,In_93);
nand U1 (N_1,In_567,In_401);
or U2 (N_2,In_445,In_45);
or U3 (N_3,In_11,In_510);
or U4 (N_4,In_193,In_880);
and U5 (N_5,In_147,In_209);
or U6 (N_6,In_678,In_149);
nor U7 (N_7,In_592,In_270);
or U8 (N_8,In_719,In_117);
nand U9 (N_9,In_708,In_480);
nand U10 (N_10,In_145,In_832);
and U11 (N_11,In_562,In_724);
nand U12 (N_12,In_604,In_98);
and U13 (N_13,In_860,In_84);
and U14 (N_14,In_721,In_677);
nand U15 (N_15,In_561,In_17);
nand U16 (N_16,In_371,In_375);
nor U17 (N_17,In_213,In_126);
nand U18 (N_18,In_57,In_827);
and U19 (N_19,In_778,In_261);
nand U20 (N_20,In_840,In_785);
nor U21 (N_21,In_535,In_389);
xnor U22 (N_22,In_484,In_771);
nor U23 (N_23,In_78,In_517);
or U24 (N_24,In_596,In_743);
or U25 (N_25,In_881,In_920);
nand U26 (N_26,In_140,In_173);
nand U27 (N_27,In_685,In_988);
nand U28 (N_28,In_781,In_965);
xor U29 (N_29,In_593,In_528);
or U30 (N_30,In_710,In_157);
xor U31 (N_31,In_674,In_862);
or U32 (N_32,In_887,In_791);
nand U33 (N_33,In_668,In_956);
and U34 (N_34,In_660,In_536);
or U35 (N_35,In_357,In_856);
nor U36 (N_36,In_489,In_493);
nand U37 (N_37,In_706,In_231);
and U38 (N_38,In_21,In_423);
nor U39 (N_39,In_699,In_795);
and U40 (N_40,In_946,In_806);
nand U41 (N_41,In_284,In_986);
nand U42 (N_42,In_717,In_430);
or U43 (N_43,In_749,In_443);
nand U44 (N_44,In_485,In_487);
and U45 (N_45,In_967,In_542);
nor U46 (N_46,In_970,In_235);
or U47 (N_47,In_899,In_886);
nand U48 (N_48,In_683,In_110);
and U49 (N_49,In_521,In_684);
nand U50 (N_50,In_306,In_702);
and U51 (N_51,In_120,In_250);
or U52 (N_52,In_625,In_419);
and U53 (N_53,In_618,In_958);
or U54 (N_54,In_633,In_497);
or U55 (N_55,In_560,In_893);
nor U56 (N_56,In_242,In_365);
nor U57 (N_57,In_488,In_913);
xor U58 (N_58,In_697,In_56);
nor U59 (N_59,In_367,In_704);
nand U60 (N_60,In_763,In_124);
nand U61 (N_61,In_324,In_449);
nand U62 (N_62,In_727,In_68);
or U63 (N_63,In_650,In_753);
nor U64 (N_64,In_969,In_470);
nor U65 (N_65,In_171,In_386);
nor U66 (N_66,In_415,In_39);
and U67 (N_67,In_450,In_595);
or U68 (N_68,In_890,In_410);
nor U69 (N_69,In_529,In_728);
or U70 (N_70,In_808,In_918);
nor U71 (N_71,In_40,In_854);
nor U72 (N_72,In_418,In_566);
and U73 (N_73,In_349,In_648);
or U74 (N_74,In_962,In_770);
and U75 (N_75,In_963,In_444);
or U76 (N_76,In_971,In_611);
nand U77 (N_77,In_281,In_514);
nor U78 (N_78,In_258,In_649);
nor U79 (N_79,In_819,In_516);
or U80 (N_80,In_764,In_119);
or U81 (N_81,In_826,In_413);
nor U82 (N_82,In_309,In_909);
and U83 (N_83,In_420,In_506);
nor U84 (N_84,In_564,In_709);
nand U85 (N_85,In_374,In_999);
nor U86 (N_86,In_786,In_533);
nand U87 (N_87,In_552,In_316);
nor U88 (N_88,In_251,In_559);
nand U89 (N_89,In_897,In_196);
and U90 (N_90,In_644,In_169);
and U91 (N_91,In_3,In_614);
and U92 (N_92,In_989,In_384);
and U93 (N_93,In_974,In_621);
and U94 (N_94,In_712,In_464);
nor U95 (N_95,In_977,In_333);
nor U96 (N_96,In_524,In_424);
nand U97 (N_97,In_328,In_898);
and U98 (N_98,In_613,In_733);
and U99 (N_99,In_782,In_872);
or U100 (N_100,In_41,In_393);
and U101 (N_101,In_900,In_783);
and U102 (N_102,In_975,In_342);
nor U103 (N_103,In_479,In_458);
nor U104 (N_104,In_50,In_576);
and U105 (N_105,In_923,In_421);
nand U106 (N_106,In_574,In_148);
and U107 (N_107,In_657,In_902);
nor U108 (N_108,In_651,In_851);
nor U109 (N_109,In_264,In_549);
nand U110 (N_110,In_65,In_315);
nand U111 (N_111,In_940,In_937);
and U112 (N_112,In_426,In_679);
or U113 (N_113,In_591,In_109);
and U114 (N_114,In_737,In_14);
and U115 (N_115,In_234,In_305);
nor U116 (N_116,In_186,In_159);
and U117 (N_117,In_780,In_994);
nor U118 (N_118,In_601,In_336);
nor U119 (N_119,In_575,In_698);
and U120 (N_120,In_757,In_500);
nand U121 (N_121,In_184,In_957);
nor U122 (N_122,In_652,In_345);
nand U123 (N_123,In_790,In_441);
and U124 (N_124,In_232,In_195);
nor U125 (N_125,In_643,In_817);
and U126 (N_126,In_486,In_891);
and U127 (N_127,In_914,In_537);
and U128 (N_128,In_285,In_278);
nor U129 (N_129,In_134,In_955);
nand U130 (N_130,In_414,In_571);
nor U131 (N_131,In_658,In_942);
or U132 (N_132,In_792,In_245);
nand U133 (N_133,In_555,In_32);
or U134 (N_134,In_387,In_432);
or U135 (N_135,In_198,In_52);
or U136 (N_136,In_118,In_948);
nand U137 (N_137,In_870,In_587);
nand U138 (N_138,In_187,In_846);
nand U139 (N_139,In_314,In_113);
nor U140 (N_140,In_277,In_578);
or U141 (N_141,In_689,In_168);
or U142 (N_142,In_824,In_20);
or U143 (N_143,In_211,In_463);
and U144 (N_144,In_615,In_908);
nand U145 (N_145,In_569,In_164);
nand U146 (N_146,In_271,In_579);
or U147 (N_147,In_54,In_176);
or U148 (N_148,In_170,In_327);
nand U149 (N_149,In_842,In_318);
nand U150 (N_150,In_453,In_473);
nor U151 (N_151,In_992,In_155);
nand U152 (N_152,In_895,In_411);
or U153 (N_153,In_539,In_835);
and U154 (N_154,In_51,In_707);
xor U155 (N_155,In_705,In_362);
or U156 (N_156,In_12,In_356);
or U157 (N_157,In_280,In_758);
or U158 (N_158,In_203,In_355);
and U159 (N_159,In_116,In_744);
nor U160 (N_160,In_274,In_761);
or U161 (N_161,In_548,In_610);
or U162 (N_162,In_976,In_404);
nor U163 (N_163,In_359,In_812);
or U164 (N_164,In_166,In_300);
and U165 (N_165,In_192,In_312);
or U166 (N_166,In_28,In_713);
nand U167 (N_167,In_291,In_563);
and U168 (N_168,In_889,In_991);
nor U169 (N_169,In_457,In_260);
or U170 (N_170,In_793,In_208);
or U171 (N_171,In_392,In_645);
nor U172 (N_172,In_153,In_1);
nand U173 (N_173,In_104,In_904);
or U174 (N_174,In_585,In_545);
nand U175 (N_175,In_804,In_233);
or U176 (N_176,In_541,In_400);
or U177 (N_177,In_573,In_163);
and U178 (N_178,In_869,In_123);
nand U179 (N_179,In_694,In_317);
nor U180 (N_180,In_935,In_960);
or U181 (N_181,In_238,In_647);
nor U182 (N_182,In_875,In_476);
nor U183 (N_183,In_547,In_538);
or U184 (N_184,In_219,In_125);
nor U185 (N_185,In_378,In_205);
and U186 (N_186,In_282,In_222);
or U187 (N_187,In_368,In_672);
xor U188 (N_188,In_48,In_332);
or U189 (N_189,In_322,In_254);
or U190 (N_190,In_436,In_105);
nand U191 (N_191,In_570,In_112);
and U192 (N_192,In_622,In_688);
nand U193 (N_193,In_326,In_814);
or U194 (N_194,In_29,In_848);
or U195 (N_195,In_304,In_402);
nor U196 (N_196,In_941,In_550);
or U197 (N_197,In_325,In_794);
nor U198 (N_198,In_691,In_616);
and U199 (N_199,In_87,In_397);
nor U200 (N_200,In_467,In_439);
nand U201 (N_201,In_24,In_228);
or U202 (N_202,In_132,In_143);
xnor U203 (N_203,In_216,In_797);
and U204 (N_204,In_917,In_929);
nor U205 (N_205,In_624,In_70);
or U206 (N_206,In_437,In_276);
and U207 (N_207,In_405,In_490);
or U208 (N_208,In_810,In_438);
nor U209 (N_209,In_36,In_221);
and U210 (N_210,In_868,In_805);
nor U211 (N_211,In_466,In_468);
or U212 (N_212,In_686,In_71);
and U213 (N_213,In_83,In_630);
nor U214 (N_214,In_499,In_952);
nand U215 (N_215,In_403,In_543);
nand U216 (N_216,In_892,In_588);
nand U217 (N_217,In_179,In_752);
nand U218 (N_218,In_653,In_383);
or U219 (N_219,In_244,In_218);
nor U220 (N_220,In_864,In_828);
nor U221 (N_221,In_905,In_509);
and U222 (N_222,In_475,In_376);
and U223 (N_223,In_504,In_428);
and U224 (N_224,In_871,In_152);
nand U225 (N_225,In_131,In_811);
or U226 (N_226,In_544,In_107);
nand U227 (N_227,In_477,In_337);
or U228 (N_228,In_617,In_982);
or U229 (N_229,In_813,In_850);
nor U230 (N_230,In_716,In_682);
and U231 (N_231,In_638,In_412);
nand U232 (N_232,In_268,In_74);
and U233 (N_233,In_460,In_101);
nand U234 (N_234,In_431,In_272);
or U235 (N_235,In_416,In_609);
and U236 (N_236,In_474,In_978);
nor U237 (N_237,In_103,In_736);
nand U238 (N_238,In_711,In_925);
nand U239 (N_239,In_354,In_767);
nand U240 (N_240,In_448,In_878);
nor U241 (N_241,In_551,In_600);
and U242 (N_242,In_247,In_725);
nor U243 (N_243,In_788,In_964);
nand U244 (N_244,In_180,In_997);
nand U245 (N_245,In_5,In_635);
or U246 (N_246,In_729,In_921);
nor U247 (N_247,In_253,In_884);
nand U248 (N_248,In_847,In_519);
or U249 (N_249,In_55,In_61);
xnor U250 (N_250,In_370,In_311);
or U251 (N_251,In_99,In_565);
xor U252 (N_252,In_755,In_321);
or U253 (N_253,In_96,In_142);
nand U254 (N_254,In_815,In_220);
and U255 (N_255,In_16,In_901);
nand U256 (N_256,In_248,In_745);
nand U257 (N_257,In_910,In_19);
nor U258 (N_258,In_602,In_252);
or U259 (N_259,In_746,In_26);
or U260 (N_260,In_382,In_523);
nor U261 (N_261,In_796,In_911);
and U262 (N_262,In_731,In_313);
and U263 (N_263,In_703,In_750);
or U264 (N_264,In_201,In_307);
nand U265 (N_265,In_557,In_27);
xor U266 (N_266,In_772,In_606);
or U267 (N_267,In_654,In_603);
nor U268 (N_268,In_135,In_379);
and U269 (N_269,In_995,In_896);
and U270 (N_270,In_993,In_25);
nor U271 (N_271,In_966,In_462);
or U272 (N_272,In_210,In_63);
nor U273 (N_273,In_531,In_390);
nand U274 (N_274,In_214,In_572);
or U275 (N_275,In_844,In_215);
and U276 (N_276,In_631,In_348);
or U277 (N_277,In_256,In_76);
and U278 (N_278,In_417,In_372);
and U279 (N_279,In_894,In_396);
or U280 (N_280,In_931,In_299);
or U281 (N_281,In_161,In_241);
or U282 (N_282,In_598,In_665);
nor U283 (N_283,In_329,In_30);
xor U284 (N_284,In_478,In_292);
nor U285 (N_285,In_381,In_515);
nand U286 (N_286,In_37,In_398);
nand U287 (N_287,In_406,In_936);
and U288 (N_288,In_69,In_81);
or U289 (N_289,In_998,In_715);
and U290 (N_290,In_18,In_175);
or U291 (N_291,In_903,In_472);
nand U292 (N_292,In_507,In_310);
xor U293 (N_293,In_446,In_89);
and U294 (N_294,In_720,In_129);
nor U295 (N_295,In_151,In_769);
nor U296 (N_296,In_366,In_915);
and U297 (N_297,In_407,In_23);
nand U298 (N_298,In_246,In_206);
nor U299 (N_299,In_380,In_981);
and U300 (N_300,In_663,In_503);
or U301 (N_301,In_287,In_738);
nor U302 (N_302,In_589,In_723);
nor U303 (N_303,In_47,In_225);
nor U304 (N_304,In_754,In_255);
and U305 (N_305,In_496,In_127);
and U306 (N_306,In_556,In_742);
and U307 (N_307,In_62,In_58);
nand U308 (N_308,In_352,In_605);
or U309 (N_309,In_774,In_773);
and U310 (N_310,In_838,In_106);
nor U311 (N_311,In_240,In_558);
nor U312 (N_312,In_154,In_434);
or U313 (N_313,In_491,In_756);
and U314 (N_314,In_79,In_294);
and U315 (N_315,In_269,In_341);
nor U316 (N_316,In_320,In_150);
or U317 (N_317,In_907,In_361);
or U318 (N_318,In_293,In_926);
and U319 (N_319,In_217,In_298);
nor U320 (N_320,In_798,In_289);
nand U321 (N_321,In_760,In_823);
nor U322 (N_322,In_695,In_237);
and U323 (N_323,In_122,In_985);
and U324 (N_324,In_227,In_130);
nand U325 (N_325,In_31,In_987);
nand U326 (N_326,In_72,In_599);
nand U327 (N_327,In_659,In_620);
nor U328 (N_328,In_641,In_953);
or U329 (N_329,In_944,In_182);
nand U330 (N_330,In_102,In_7);
or U331 (N_331,In_15,In_800);
and U332 (N_332,In_38,In_197);
nand U333 (N_333,In_865,In_673);
and U334 (N_334,In_747,In_360);
and U335 (N_335,In_459,In_94);
xor U336 (N_336,In_88,In_91);
or U337 (N_337,In_288,In_732);
nand U338 (N_338,In_836,In_303);
nor U339 (N_339,In_597,In_748);
nand U340 (N_340,In_849,In_534);
nand U341 (N_341,In_308,In_973);
nand U342 (N_342,In_816,In_980);
xor U343 (N_343,In_863,In_223);
nand U344 (N_344,In_801,In_492);
and U345 (N_345,In_111,In_671);
nand U346 (N_346,In_498,In_857);
nor U347 (N_347,In_799,In_687);
or U348 (N_348,In_158,In_640);
or U349 (N_349,In_740,In_73);
and U350 (N_350,In_821,In_162);
or U351 (N_351,In_373,In_273);
and U352 (N_352,In_353,In_789);
and U353 (N_353,In_133,In_207);
nand U354 (N_354,In_584,In_820);
or U355 (N_355,In_67,In_347);
nand U356 (N_356,In_2,In_984);
nor U357 (N_357,In_581,In_114);
and U358 (N_358,In_199,In_178);
xnor U359 (N_359,In_204,In_66);
xnor U360 (N_360,In_42,In_85);
xnor U361 (N_361,In_136,In_714);
xor U362 (N_362,In_751,In_961);
or U363 (N_363,In_185,In_825);
or U364 (N_364,In_239,In_950);
nand U365 (N_365,In_391,In_331);
nand U366 (N_366,In_979,In_661);
nor U367 (N_367,In_249,In_730);
and U368 (N_368,In_520,In_577);
and U369 (N_369,In_676,In_667);
and U370 (N_370,In_666,In_4);
nand U371 (N_371,In_831,In_646);
or U372 (N_372,In_43,In_634);
nor U373 (N_373,In_885,In_837);
nor U374 (N_374,In_481,In_809);
nor U375 (N_375,In_664,In_363);
nand U376 (N_376,In_283,In_90);
nand U377 (N_377,In_302,In_339);
nand U378 (N_378,In_934,In_422);
or U379 (N_379,In_874,In_526);
xor U380 (N_380,In_82,In_429);
or U381 (N_381,In_59,In_843);
and U382 (N_382,In_922,In_512);
nand U383 (N_383,In_696,In_912);
or U384 (N_384,In_335,In_718);
nand U385 (N_385,In_121,In_642);
nor U386 (N_386,In_295,In_834);
or U387 (N_387,In_160,In_983);
nand U388 (N_388,In_167,In_177);
or U389 (N_389,In_330,In_408);
nand U390 (N_390,In_334,In_959);
and U391 (N_391,In_968,In_680);
and U392 (N_392,In_97,In_230);
nor U393 (N_393,In_628,In_852);
or U394 (N_394,In_833,In_859);
nor U395 (N_395,In_933,In_637);
nor U396 (N_396,In_845,In_582);
nor U397 (N_397,In_626,In_80);
nor U398 (N_398,In_165,In_511);
nor U399 (N_399,In_469,In_266);
and U400 (N_400,In_141,In_346);
nand U401 (N_401,In_358,In_802);
xnor U402 (N_402,In_279,In_409);
and U403 (N_403,In_8,In_435);
or U404 (N_404,In_456,In_619);
nor U405 (N_405,In_873,In_92);
or U406 (N_406,In_505,In_632);
and U407 (N_407,In_275,In_265);
nand U408 (N_408,In_0,In_191);
or U409 (N_409,In_49,In_501);
or U410 (N_410,In_882,In_267);
and U411 (N_411,In_340,In_629);
xnor U412 (N_412,In_768,In_440);
and U413 (N_413,In_947,In_452);
nand U414 (N_414,In_156,In_675);
and U415 (N_415,In_427,In_943);
or U416 (N_416,In_766,In_447);
and U417 (N_417,In_951,In_369);
and U418 (N_418,In_385,In_181);
nand U419 (N_419,In_494,In_502);
or U420 (N_420,In_338,In_229);
or U421 (N_421,In_35,In_46);
nand U422 (N_422,In_351,In_739);
or U423 (N_423,In_701,In_442);
and U424 (N_424,In_779,In_879);
and U425 (N_425,In_286,In_829);
nand U426 (N_426,In_513,In_77);
xor U427 (N_427,In_323,In_741);
nand U428 (N_428,In_855,In_395);
xor U429 (N_429,In_692,In_734);
and U430 (N_430,In_95,In_100);
nand U431 (N_431,In_669,In_930);
nand U432 (N_432,In_44,In_906);
nand U433 (N_433,In_656,In_568);
and U434 (N_434,In_916,In_13);
nor U435 (N_435,In_700,In_224);
nand U436 (N_436,In_482,In_296);
nor U437 (N_437,In_670,In_853);
nor U438 (N_438,In_841,In_939);
nand U439 (N_439,In_867,In_608);
nor U440 (N_440,In_454,In_919);
or U441 (N_441,In_583,In_425);
nor U442 (N_442,In_580,In_33);
nor U443 (N_443,In_188,In_590);
and U444 (N_444,In_259,In_818);
and U445 (N_445,In_144,In_839);
or U446 (N_446,In_928,In_722);
nor U447 (N_447,In_607,In_433);
nor U448 (N_448,In_861,In_257);
nor U449 (N_449,In_344,In_927);
nor U450 (N_450,In_765,In_471);
and U451 (N_451,In_525,In_190);
nand U452 (N_452,In_877,In_301);
nor U453 (N_453,In_639,In_775);
or U454 (N_454,In_532,In_949);
nand U455 (N_455,In_586,In_866);
or U456 (N_456,In_681,In_726);
nor U457 (N_457,In_461,In_522);
nor U458 (N_458,In_212,In_954);
nor U459 (N_459,In_350,In_693);
nand U460 (N_460,In_262,In_495);
nand U461 (N_461,In_60,In_655);
or U462 (N_462,In_394,In_777);
nor U463 (N_463,In_858,In_75);
or U464 (N_464,In_183,In_388);
nand U465 (N_465,In_759,In_883);
nor U466 (N_466,In_172,In_189);
or U467 (N_467,In_876,In_465);
nand U468 (N_468,In_996,In_451);
or U469 (N_469,In_623,In_594);
nor U470 (N_470,In_9,In_128);
or U471 (N_471,In_787,In_822);
xor U472 (N_472,In_53,In_6);
nor U473 (N_473,In_86,In_762);
nand U474 (N_474,In_200,In_662);
nor U475 (N_475,In_34,In_319);
nand U476 (N_476,In_945,In_553);
or U477 (N_477,In_139,In_364);
nor U478 (N_478,In_137,In_612);
nor U479 (N_479,In_22,In_636);
or U480 (N_480,In_932,In_830);
or U481 (N_481,In_455,In_735);
nor U482 (N_482,In_174,In_297);
and U483 (N_483,In_243,In_546);
and U484 (N_484,In_377,In_924);
and U485 (N_485,In_108,In_236);
nor U486 (N_486,In_690,In_290);
or U487 (N_487,In_64,In_938);
or U488 (N_488,In_888,In_115);
xor U489 (N_489,In_226,In_138);
or U490 (N_490,In_554,In_527);
and U491 (N_491,In_803,In_483);
or U492 (N_492,In_146,In_627);
nor U493 (N_493,In_530,In_508);
or U494 (N_494,In_784,In_263);
nor U495 (N_495,In_202,In_399);
and U496 (N_496,In_990,In_540);
and U497 (N_497,In_807,In_10);
or U498 (N_498,In_194,In_518);
nand U499 (N_499,In_343,In_776);
or U500 (N_500,In_303,In_306);
and U501 (N_501,In_682,In_310);
or U502 (N_502,In_321,In_4);
nand U503 (N_503,In_587,In_344);
and U504 (N_504,In_546,In_833);
or U505 (N_505,In_508,In_917);
and U506 (N_506,In_740,In_844);
nor U507 (N_507,In_785,In_842);
and U508 (N_508,In_531,In_2);
nand U509 (N_509,In_620,In_678);
or U510 (N_510,In_655,In_532);
nand U511 (N_511,In_385,In_520);
xnor U512 (N_512,In_525,In_969);
and U513 (N_513,In_465,In_26);
and U514 (N_514,In_420,In_359);
and U515 (N_515,In_422,In_663);
or U516 (N_516,In_549,In_554);
nor U517 (N_517,In_558,In_178);
nor U518 (N_518,In_468,In_705);
nand U519 (N_519,In_971,In_559);
and U520 (N_520,In_98,In_979);
and U521 (N_521,In_850,In_505);
or U522 (N_522,In_338,In_43);
nand U523 (N_523,In_611,In_709);
nand U524 (N_524,In_426,In_665);
and U525 (N_525,In_889,In_585);
and U526 (N_526,In_353,In_888);
nor U527 (N_527,In_832,In_228);
or U528 (N_528,In_570,In_509);
and U529 (N_529,In_9,In_930);
nand U530 (N_530,In_33,In_173);
and U531 (N_531,In_664,In_956);
and U532 (N_532,In_941,In_750);
or U533 (N_533,In_853,In_927);
or U534 (N_534,In_476,In_492);
and U535 (N_535,In_151,In_344);
nor U536 (N_536,In_731,In_942);
nor U537 (N_537,In_13,In_547);
nor U538 (N_538,In_574,In_559);
nor U539 (N_539,In_409,In_515);
nand U540 (N_540,In_819,In_287);
or U541 (N_541,In_663,In_19);
or U542 (N_542,In_511,In_625);
nand U543 (N_543,In_778,In_194);
nand U544 (N_544,In_437,In_700);
or U545 (N_545,In_724,In_633);
nor U546 (N_546,In_592,In_107);
or U547 (N_547,In_194,In_266);
nand U548 (N_548,In_557,In_766);
and U549 (N_549,In_602,In_150);
nor U550 (N_550,In_371,In_836);
and U551 (N_551,In_109,In_206);
or U552 (N_552,In_820,In_732);
or U553 (N_553,In_519,In_555);
and U554 (N_554,In_485,In_403);
or U555 (N_555,In_500,In_669);
nor U556 (N_556,In_833,In_221);
or U557 (N_557,In_784,In_475);
or U558 (N_558,In_413,In_383);
nor U559 (N_559,In_839,In_31);
or U560 (N_560,In_738,In_167);
or U561 (N_561,In_576,In_851);
xor U562 (N_562,In_688,In_16);
or U563 (N_563,In_158,In_232);
xnor U564 (N_564,In_603,In_21);
or U565 (N_565,In_427,In_579);
xor U566 (N_566,In_422,In_627);
or U567 (N_567,In_94,In_349);
nand U568 (N_568,In_599,In_627);
and U569 (N_569,In_924,In_804);
or U570 (N_570,In_163,In_361);
nor U571 (N_571,In_243,In_96);
nor U572 (N_572,In_255,In_196);
and U573 (N_573,In_761,In_604);
nor U574 (N_574,In_572,In_138);
nor U575 (N_575,In_683,In_522);
nand U576 (N_576,In_917,In_711);
nor U577 (N_577,In_154,In_848);
nand U578 (N_578,In_209,In_41);
or U579 (N_579,In_324,In_669);
nand U580 (N_580,In_859,In_820);
and U581 (N_581,In_749,In_132);
or U582 (N_582,In_284,In_447);
or U583 (N_583,In_74,In_237);
or U584 (N_584,In_626,In_821);
nor U585 (N_585,In_499,In_847);
nand U586 (N_586,In_804,In_252);
and U587 (N_587,In_735,In_391);
nor U588 (N_588,In_671,In_292);
nor U589 (N_589,In_955,In_791);
nor U590 (N_590,In_788,In_936);
and U591 (N_591,In_363,In_390);
and U592 (N_592,In_345,In_815);
or U593 (N_593,In_213,In_348);
or U594 (N_594,In_382,In_647);
nor U595 (N_595,In_677,In_702);
nor U596 (N_596,In_835,In_70);
and U597 (N_597,In_840,In_674);
or U598 (N_598,In_642,In_208);
nand U599 (N_599,In_944,In_40);
nor U600 (N_600,In_750,In_788);
nand U601 (N_601,In_986,In_348);
and U602 (N_602,In_258,In_624);
nor U603 (N_603,In_682,In_554);
and U604 (N_604,In_939,In_109);
nand U605 (N_605,In_114,In_512);
nor U606 (N_606,In_674,In_324);
or U607 (N_607,In_503,In_746);
or U608 (N_608,In_678,In_390);
nand U609 (N_609,In_637,In_854);
or U610 (N_610,In_338,In_90);
nand U611 (N_611,In_914,In_936);
and U612 (N_612,In_330,In_393);
or U613 (N_613,In_178,In_914);
or U614 (N_614,In_338,In_547);
nor U615 (N_615,In_329,In_996);
or U616 (N_616,In_60,In_515);
and U617 (N_617,In_215,In_689);
or U618 (N_618,In_640,In_282);
and U619 (N_619,In_402,In_136);
and U620 (N_620,In_236,In_995);
or U621 (N_621,In_850,In_259);
nor U622 (N_622,In_724,In_13);
or U623 (N_623,In_79,In_326);
or U624 (N_624,In_732,In_836);
nand U625 (N_625,In_488,In_557);
nand U626 (N_626,In_837,In_60);
nand U627 (N_627,In_377,In_538);
or U628 (N_628,In_127,In_951);
nand U629 (N_629,In_648,In_278);
nand U630 (N_630,In_971,In_585);
nor U631 (N_631,In_443,In_864);
nor U632 (N_632,In_559,In_614);
nand U633 (N_633,In_714,In_754);
or U634 (N_634,In_669,In_817);
nand U635 (N_635,In_799,In_910);
or U636 (N_636,In_21,In_515);
and U637 (N_637,In_232,In_373);
nor U638 (N_638,In_965,In_340);
or U639 (N_639,In_445,In_657);
and U640 (N_640,In_290,In_553);
and U641 (N_641,In_571,In_137);
nor U642 (N_642,In_749,In_807);
nand U643 (N_643,In_131,In_979);
nor U644 (N_644,In_117,In_19);
nor U645 (N_645,In_561,In_980);
nand U646 (N_646,In_781,In_300);
and U647 (N_647,In_176,In_25);
and U648 (N_648,In_199,In_373);
nand U649 (N_649,In_399,In_746);
and U650 (N_650,In_760,In_221);
nand U651 (N_651,In_373,In_141);
nand U652 (N_652,In_597,In_71);
nand U653 (N_653,In_396,In_810);
nand U654 (N_654,In_632,In_341);
nand U655 (N_655,In_725,In_228);
nor U656 (N_656,In_15,In_331);
or U657 (N_657,In_614,In_634);
nor U658 (N_658,In_238,In_676);
nand U659 (N_659,In_651,In_116);
nand U660 (N_660,In_701,In_539);
nand U661 (N_661,In_485,In_636);
xnor U662 (N_662,In_808,In_220);
nor U663 (N_663,In_796,In_533);
nand U664 (N_664,In_200,In_960);
or U665 (N_665,In_56,In_367);
nor U666 (N_666,In_244,In_142);
or U667 (N_667,In_243,In_128);
nor U668 (N_668,In_442,In_828);
and U669 (N_669,In_377,In_244);
nand U670 (N_670,In_981,In_153);
nand U671 (N_671,In_262,In_100);
nand U672 (N_672,In_143,In_270);
nor U673 (N_673,In_816,In_204);
nor U674 (N_674,In_22,In_12);
nor U675 (N_675,In_630,In_96);
or U676 (N_676,In_970,In_640);
and U677 (N_677,In_815,In_38);
and U678 (N_678,In_180,In_798);
nor U679 (N_679,In_235,In_43);
nor U680 (N_680,In_923,In_864);
and U681 (N_681,In_540,In_963);
and U682 (N_682,In_218,In_394);
nand U683 (N_683,In_453,In_63);
nor U684 (N_684,In_409,In_641);
nand U685 (N_685,In_120,In_910);
or U686 (N_686,In_118,In_613);
nor U687 (N_687,In_827,In_714);
or U688 (N_688,In_58,In_302);
nand U689 (N_689,In_789,In_565);
nand U690 (N_690,In_513,In_942);
or U691 (N_691,In_910,In_273);
nor U692 (N_692,In_176,In_622);
and U693 (N_693,In_653,In_148);
and U694 (N_694,In_605,In_129);
nand U695 (N_695,In_48,In_899);
nor U696 (N_696,In_211,In_77);
or U697 (N_697,In_283,In_846);
nor U698 (N_698,In_996,In_161);
nor U699 (N_699,In_317,In_324);
or U700 (N_700,In_278,In_923);
or U701 (N_701,In_855,In_902);
nand U702 (N_702,In_508,In_834);
nand U703 (N_703,In_662,In_265);
xnor U704 (N_704,In_433,In_288);
nand U705 (N_705,In_461,In_620);
nand U706 (N_706,In_515,In_605);
nand U707 (N_707,In_831,In_292);
or U708 (N_708,In_80,In_44);
or U709 (N_709,In_574,In_684);
nor U710 (N_710,In_931,In_93);
nand U711 (N_711,In_337,In_7);
and U712 (N_712,In_416,In_299);
and U713 (N_713,In_550,In_661);
and U714 (N_714,In_829,In_468);
and U715 (N_715,In_817,In_903);
and U716 (N_716,In_189,In_380);
and U717 (N_717,In_238,In_511);
nor U718 (N_718,In_995,In_214);
nand U719 (N_719,In_650,In_756);
nor U720 (N_720,In_673,In_339);
nor U721 (N_721,In_662,In_552);
nand U722 (N_722,In_258,In_517);
xnor U723 (N_723,In_95,In_628);
or U724 (N_724,In_406,In_241);
nand U725 (N_725,In_373,In_731);
xor U726 (N_726,In_967,In_720);
nor U727 (N_727,In_137,In_315);
nand U728 (N_728,In_883,In_443);
nand U729 (N_729,In_850,In_957);
nor U730 (N_730,In_835,In_148);
nor U731 (N_731,In_621,In_853);
nor U732 (N_732,In_953,In_946);
nor U733 (N_733,In_224,In_970);
nor U734 (N_734,In_301,In_705);
nor U735 (N_735,In_347,In_297);
or U736 (N_736,In_517,In_884);
nand U737 (N_737,In_761,In_303);
nand U738 (N_738,In_319,In_817);
or U739 (N_739,In_320,In_382);
and U740 (N_740,In_757,In_847);
nand U741 (N_741,In_218,In_776);
nand U742 (N_742,In_519,In_447);
nand U743 (N_743,In_135,In_182);
or U744 (N_744,In_204,In_451);
nor U745 (N_745,In_34,In_640);
xnor U746 (N_746,In_711,In_132);
nor U747 (N_747,In_768,In_783);
and U748 (N_748,In_945,In_977);
and U749 (N_749,In_97,In_40);
nand U750 (N_750,In_932,In_238);
nand U751 (N_751,In_165,In_320);
nor U752 (N_752,In_328,In_643);
or U753 (N_753,In_478,In_757);
nand U754 (N_754,In_886,In_752);
and U755 (N_755,In_739,In_113);
and U756 (N_756,In_355,In_358);
xnor U757 (N_757,In_842,In_739);
nand U758 (N_758,In_329,In_656);
nor U759 (N_759,In_207,In_825);
and U760 (N_760,In_203,In_354);
nand U761 (N_761,In_126,In_184);
and U762 (N_762,In_804,In_45);
or U763 (N_763,In_79,In_533);
nor U764 (N_764,In_865,In_112);
and U765 (N_765,In_112,In_232);
nand U766 (N_766,In_127,In_871);
nand U767 (N_767,In_661,In_101);
and U768 (N_768,In_992,In_693);
and U769 (N_769,In_362,In_75);
or U770 (N_770,In_241,In_609);
xnor U771 (N_771,In_754,In_955);
or U772 (N_772,In_377,In_965);
nor U773 (N_773,In_702,In_601);
or U774 (N_774,In_16,In_595);
nor U775 (N_775,In_406,In_437);
nor U776 (N_776,In_349,In_614);
nand U777 (N_777,In_761,In_327);
or U778 (N_778,In_124,In_146);
and U779 (N_779,In_972,In_684);
or U780 (N_780,In_432,In_408);
and U781 (N_781,In_85,In_169);
and U782 (N_782,In_774,In_309);
and U783 (N_783,In_931,In_978);
and U784 (N_784,In_858,In_512);
or U785 (N_785,In_534,In_349);
nor U786 (N_786,In_119,In_901);
nand U787 (N_787,In_829,In_525);
nor U788 (N_788,In_845,In_416);
nor U789 (N_789,In_609,In_227);
nand U790 (N_790,In_734,In_693);
or U791 (N_791,In_318,In_110);
nor U792 (N_792,In_631,In_124);
and U793 (N_793,In_765,In_77);
nand U794 (N_794,In_594,In_555);
nor U795 (N_795,In_626,In_696);
and U796 (N_796,In_729,In_273);
nand U797 (N_797,In_342,In_247);
and U798 (N_798,In_17,In_867);
nor U799 (N_799,In_475,In_626);
or U800 (N_800,In_973,In_923);
nor U801 (N_801,In_539,In_834);
nor U802 (N_802,In_3,In_575);
or U803 (N_803,In_886,In_285);
and U804 (N_804,In_54,In_964);
nand U805 (N_805,In_269,In_32);
or U806 (N_806,In_857,In_429);
or U807 (N_807,In_100,In_146);
or U808 (N_808,In_251,In_495);
or U809 (N_809,In_883,In_815);
nand U810 (N_810,In_327,In_910);
nand U811 (N_811,In_213,In_848);
nor U812 (N_812,In_545,In_582);
and U813 (N_813,In_57,In_957);
and U814 (N_814,In_85,In_179);
or U815 (N_815,In_289,In_990);
and U816 (N_816,In_578,In_395);
nand U817 (N_817,In_650,In_589);
or U818 (N_818,In_191,In_491);
and U819 (N_819,In_455,In_505);
or U820 (N_820,In_40,In_666);
and U821 (N_821,In_20,In_985);
nand U822 (N_822,In_1,In_660);
or U823 (N_823,In_768,In_227);
nand U824 (N_824,In_77,In_934);
and U825 (N_825,In_409,In_76);
and U826 (N_826,In_722,In_10);
and U827 (N_827,In_602,In_393);
and U828 (N_828,In_873,In_598);
and U829 (N_829,In_298,In_348);
and U830 (N_830,In_733,In_124);
nand U831 (N_831,In_950,In_406);
nand U832 (N_832,In_229,In_908);
or U833 (N_833,In_732,In_821);
nor U834 (N_834,In_640,In_693);
nor U835 (N_835,In_954,In_999);
nand U836 (N_836,In_785,In_295);
and U837 (N_837,In_630,In_238);
nor U838 (N_838,In_840,In_456);
nand U839 (N_839,In_855,In_664);
nand U840 (N_840,In_152,In_863);
nor U841 (N_841,In_638,In_904);
nor U842 (N_842,In_587,In_528);
or U843 (N_843,In_418,In_128);
nand U844 (N_844,In_113,In_238);
or U845 (N_845,In_518,In_43);
nand U846 (N_846,In_102,In_786);
or U847 (N_847,In_938,In_189);
or U848 (N_848,In_858,In_259);
or U849 (N_849,In_957,In_672);
nor U850 (N_850,In_5,In_700);
nor U851 (N_851,In_844,In_999);
nand U852 (N_852,In_240,In_416);
nand U853 (N_853,In_308,In_796);
nand U854 (N_854,In_699,In_349);
nor U855 (N_855,In_100,In_433);
or U856 (N_856,In_104,In_389);
nand U857 (N_857,In_199,In_862);
nand U858 (N_858,In_822,In_868);
or U859 (N_859,In_826,In_225);
nor U860 (N_860,In_915,In_37);
nor U861 (N_861,In_24,In_13);
nor U862 (N_862,In_696,In_316);
xor U863 (N_863,In_640,In_779);
and U864 (N_864,In_478,In_701);
nor U865 (N_865,In_627,In_910);
xor U866 (N_866,In_429,In_909);
and U867 (N_867,In_603,In_818);
and U868 (N_868,In_839,In_900);
and U869 (N_869,In_478,In_158);
and U870 (N_870,In_744,In_816);
and U871 (N_871,In_418,In_659);
nor U872 (N_872,In_620,In_384);
or U873 (N_873,In_198,In_904);
or U874 (N_874,In_41,In_537);
nor U875 (N_875,In_851,In_910);
or U876 (N_876,In_145,In_708);
nand U877 (N_877,In_975,In_39);
and U878 (N_878,In_357,In_396);
or U879 (N_879,In_789,In_156);
and U880 (N_880,In_563,In_706);
and U881 (N_881,In_331,In_950);
nand U882 (N_882,In_670,In_522);
nand U883 (N_883,In_135,In_547);
or U884 (N_884,In_546,In_113);
nor U885 (N_885,In_632,In_968);
nand U886 (N_886,In_264,In_584);
or U887 (N_887,In_525,In_251);
or U888 (N_888,In_760,In_572);
nand U889 (N_889,In_109,In_291);
nor U890 (N_890,In_917,In_306);
and U891 (N_891,In_968,In_778);
nor U892 (N_892,In_831,In_182);
nor U893 (N_893,In_382,In_898);
and U894 (N_894,In_825,In_215);
nor U895 (N_895,In_174,In_973);
and U896 (N_896,In_206,In_370);
nand U897 (N_897,In_919,In_374);
nand U898 (N_898,In_865,In_885);
or U899 (N_899,In_224,In_76);
or U900 (N_900,In_232,In_968);
and U901 (N_901,In_444,In_418);
nand U902 (N_902,In_595,In_423);
nor U903 (N_903,In_760,In_934);
and U904 (N_904,In_304,In_969);
nand U905 (N_905,In_303,In_543);
and U906 (N_906,In_463,In_449);
or U907 (N_907,In_770,In_643);
and U908 (N_908,In_478,In_129);
or U909 (N_909,In_58,In_915);
nand U910 (N_910,In_488,In_516);
or U911 (N_911,In_344,In_449);
nor U912 (N_912,In_830,In_971);
nand U913 (N_913,In_677,In_276);
or U914 (N_914,In_994,In_633);
nand U915 (N_915,In_324,In_161);
and U916 (N_916,In_310,In_938);
nand U917 (N_917,In_194,In_294);
and U918 (N_918,In_471,In_775);
nand U919 (N_919,In_38,In_144);
nor U920 (N_920,In_53,In_988);
nor U921 (N_921,In_862,In_436);
or U922 (N_922,In_761,In_314);
nand U923 (N_923,In_187,In_517);
nand U924 (N_924,In_54,In_373);
and U925 (N_925,In_899,In_941);
nor U926 (N_926,In_244,In_108);
and U927 (N_927,In_55,In_947);
or U928 (N_928,In_120,In_688);
and U929 (N_929,In_505,In_325);
nor U930 (N_930,In_215,In_657);
nor U931 (N_931,In_254,In_967);
or U932 (N_932,In_396,In_489);
nand U933 (N_933,In_219,In_43);
nand U934 (N_934,In_434,In_766);
and U935 (N_935,In_323,In_868);
or U936 (N_936,In_168,In_593);
and U937 (N_937,In_328,In_105);
nor U938 (N_938,In_352,In_34);
nor U939 (N_939,In_305,In_383);
nor U940 (N_940,In_228,In_4);
and U941 (N_941,In_103,In_861);
nor U942 (N_942,In_595,In_280);
nand U943 (N_943,In_271,In_1);
nand U944 (N_944,In_583,In_266);
and U945 (N_945,In_428,In_62);
and U946 (N_946,In_704,In_564);
and U947 (N_947,In_109,In_133);
and U948 (N_948,In_11,In_276);
or U949 (N_949,In_520,In_961);
nor U950 (N_950,In_93,In_342);
nor U951 (N_951,In_140,In_698);
nor U952 (N_952,In_270,In_867);
nand U953 (N_953,In_702,In_224);
nor U954 (N_954,In_65,In_147);
or U955 (N_955,In_807,In_409);
xnor U956 (N_956,In_967,In_849);
nor U957 (N_957,In_106,In_898);
nand U958 (N_958,In_111,In_934);
or U959 (N_959,In_446,In_643);
xor U960 (N_960,In_41,In_124);
or U961 (N_961,In_315,In_349);
nor U962 (N_962,In_154,In_632);
and U963 (N_963,In_585,In_324);
and U964 (N_964,In_574,In_264);
nor U965 (N_965,In_814,In_277);
or U966 (N_966,In_172,In_361);
and U967 (N_967,In_219,In_257);
or U968 (N_968,In_64,In_445);
and U969 (N_969,In_810,In_204);
nand U970 (N_970,In_926,In_476);
and U971 (N_971,In_455,In_269);
and U972 (N_972,In_553,In_530);
or U973 (N_973,In_546,In_952);
or U974 (N_974,In_413,In_104);
or U975 (N_975,In_671,In_467);
and U976 (N_976,In_888,In_569);
nand U977 (N_977,In_115,In_338);
nor U978 (N_978,In_747,In_764);
or U979 (N_979,In_845,In_231);
nand U980 (N_980,In_482,In_768);
nand U981 (N_981,In_388,In_810);
nand U982 (N_982,In_573,In_590);
or U983 (N_983,In_901,In_925);
nand U984 (N_984,In_250,In_72);
nand U985 (N_985,In_944,In_721);
and U986 (N_986,In_121,In_510);
nand U987 (N_987,In_571,In_994);
nor U988 (N_988,In_297,In_636);
nor U989 (N_989,In_75,In_211);
nor U990 (N_990,In_540,In_542);
nand U991 (N_991,In_211,In_500);
nand U992 (N_992,In_388,In_609);
nor U993 (N_993,In_918,In_632);
nor U994 (N_994,In_135,In_27);
xnor U995 (N_995,In_438,In_784);
nor U996 (N_996,In_721,In_146);
and U997 (N_997,In_361,In_335);
nor U998 (N_998,In_87,In_284);
nor U999 (N_999,In_525,In_203);
nor U1000 (N_1000,In_939,In_44);
nand U1001 (N_1001,In_62,In_769);
nor U1002 (N_1002,In_136,In_306);
nand U1003 (N_1003,In_785,In_487);
and U1004 (N_1004,In_586,In_287);
xor U1005 (N_1005,In_344,In_467);
nand U1006 (N_1006,In_698,In_284);
nor U1007 (N_1007,In_617,In_944);
nand U1008 (N_1008,In_162,In_205);
nor U1009 (N_1009,In_542,In_254);
nor U1010 (N_1010,In_928,In_102);
nand U1011 (N_1011,In_645,In_837);
or U1012 (N_1012,In_224,In_498);
nor U1013 (N_1013,In_752,In_127);
and U1014 (N_1014,In_595,In_713);
or U1015 (N_1015,In_26,In_979);
nand U1016 (N_1016,In_693,In_752);
nor U1017 (N_1017,In_723,In_712);
nand U1018 (N_1018,In_916,In_327);
nand U1019 (N_1019,In_982,In_336);
nand U1020 (N_1020,In_755,In_323);
nor U1021 (N_1021,In_61,In_372);
nor U1022 (N_1022,In_505,In_460);
or U1023 (N_1023,In_147,In_110);
nand U1024 (N_1024,In_883,In_473);
or U1025 (N_1025,In_437,In_351);
and U1026 (N_1026,In_556,In_81);
nand U1027 (N_1027,In_988,In_3);
or U1028 (N_1028,In_513,In_645);
and U1029 (N_1029,In_154,In_857);
and U1030 (N_1030,In_530,In_514);
and U1031 (N_1031,In_826,In_877);
nor U1032 (N_1032,In_837,In_855);
or U1033 (N_1033,In_677,In_975);
or U1034 (N_1034,In_734,In_875);
and U1035 (N_1035,In_394,In_58);
and U1036 (N_1036,In_102,In_675);
nand U1037 (N_1037,In_938,In_859);
nor U1038 (N_1038,In_228,In_912);
nor U1039 (N_1039,In_224,In_20);
and U1040 (N_1040,In_32,In_820);
or U1041 (N_1041,In_118,In_947);
and U1042 (N_1042,In_622,In_848);
nand U1043 (N_1043,In_465,In_169);
or U1044 (N_1044,In_484,In_987);
nor U1045 (N_1045,In_580,In_150);
nand U1046 (N_1046,In_944,In_129);
or U1047 (N_1047,In_649,In_861);
nand U1048 (N_1048,In_807,In_523);
and U1049 (N_1049,In_842,In_403);
or U1050 (N_1050,In_313,In_716);
nor U1051 (N_1051,In_351,In_404);
nand U1052 (N_1052,In_388,In_727);
or U1053 (N_1053,In_507,In_609);
xor U1054 (N_1054,In_243,In_933);
nand U1055 (N_1055,In_205,In_606);
and U1056 (N_1056,In_13,In_159);
nor U1057 (N_1057,In_470,In_417);
nand U1058 (N_1058,In_890,In_545);
nand U1059 (N_1059,In_604,In_43);
or U1060 (N_1060,In_188,In_289);
nand U1061 (N_1061,In_718,In_647);
and U1062 (N_1062,In_685,In_451);
nand U1063 (N_1063,In_474,In_75);
nor U1064 (N_1064,In_926,In_893);
xnor U1065 (N_1065,In_443,In_868);
and U1066 (N_1066,In_453,In_556);
or U1067 (N_1067,In_166,In_625);
nand U1068 (N_1068,In_107,In_275);
xnor U1069 (N_1069,In_156,In_878);
and U1070 (N_1070,In_172,In_653);
nand U1071 (N_1071,In_479,In_228);
and U1072 (N_1072,In_357,In_395);
nor U1073 (N_1073,In_346,In_836);
or U1074 (N_1074,In_468,In_605);
or U1075 (N_1075,In_566,In_776);
nor U1076 (N_1076,In_733,In_909);
or U1077 (N_1077,In_998,In_190);
nand U1078 (N_1078,In_734,In_757);
nand U1079 (N_1079,In_980,In_941);
nand U1080 (N_1080,In_410,In_203);
or U1081 (N_1081,In_994,In_287);
or U1082 (N_1082,In_794,In_769);
and U1083 (N_1083,In_339,In_91);
and U1084 (N_1084,In_8,In_707);
nor U1085 (N_1085,In_599,In_27);
or U1086 (N_1086,In_239,In_246);
and U1087 (N_1087,In_260,In_880);
nor U1088 (N_1088,In_89,In_384);
nor U1089 (N_1089,In_953,In_987);
and U1090 (N_1090,In_502,In_927);
nor U1091 (N_1091,In_845,In_810);
nand U1092 (N_1092,In_71,In_389);
and U1093 (N_1093,In_580,In_273);
or U1094 (N_1094,In_292,In_918);
nor U1095 (N_1095,In_90,In_51);
nand U1096 (N_1096,In_390,In_771);
or U1097 (N_1097,In_623,In_467);
and U1098 (N_1098,In_505,In_491);
nand U1099 (N_1099,In_970,In_930);
and U1100 (N_1100,In_215,In_554);
nand U1101 (N_1101,In_708,In_63);
or U1102 (N_1102,In_443,In_19);
xnor U1103 (N_1103,In_283,In_145);
nand U1104 (N_1104,In_904,In_297);
or U1105 (N_1105,In_438,In_981);
and U1106 (N_1106,In_978,In_394);
nor U1107 (N_1107,In_594,In_334);
nor U1108 (N_1108,In_767,In_50);
nand U1109 (N_1109,In_691,In_518);
nand U1110 (N_1110,In_416,In_690);
and U1111 (N_1111,In_714,In_290);
and U1112 (N_1112,In_592,In_973);
or U1113 (N_1113,In_625,In_263);
or U1114 (N_1114,In_558,In_593);
nor U1115 (N_1115,In_251,In_545);
xnor U1116 (N_1116,In_766,In_908);
or U1117 (N_1117,In_937,In_769);
nand U1118 (N_1118,In_398,In_127);
or U1119 (N_1119,In_469,In_18);
or U1120 (N_1120,In_732,In_117);
or U1121 (N_1121,In_715,In_801);
nand U1122 (N_1122,In_687,In_121);
or U1123 (N_1123,In_392,In_475);
nor U1124 (N_1124,In_24,In_725);
or U1125 (N_1125,In_764,In_982);
nand U1126 (N_1126,In_562,In_773);
nand U1127 (N_1127,In_495,In_345);
and U1128 (N_1128,In_605,In_197);
or U1129 (N_1129,In_655,In_160);
or U1130 (N_1130,In_793,In_610);
nor U1131 (N_1131,In_440,In_814);
nor U1132 (N_1132,In_689,In_374);
or U1133 (N_1133,In_719,In_730);
and U1134 (N_1134,In_109,In_977);
nand U1135 (N_1135,In_167,In_777);
and U1136 (N_1136,In_417,In_494);
and U1137 (N_1137,In_212,In_686);
and U1138 (N_1138,In_789,In_410);
or U1139 (N_1139,In_601,In_455);
nor U1140 (N_1140,In_483,In_701);
nand U1141 (N_1141,In_561,In_697);
or U1142 (N_1142,In_361,In_142);
nor U1143 (N_1143,In_472,In_67);
or U1144 (N_1144,In_506,In_372);
or U1145 (N_1145,In_509,In_962);
xnor U1146 (N_1146,In_943,In_105);
nor U1147 (N_1147,In_305,In_46);
or U1148 (N_1148,In_295,In_960);
or U1149 (N_1149,In_696,In_522);
xnor U1150 (N_1150,In_171,In_474);
nand U1151 (N_1151,In_560,In_367);
or U1152 (N_1152,In_288,In_523);
and U1153 (N_1153,In_877,In_835);
and U1154 (N_1154,In_737,In_307);
or U1155 (N_1155,In_243,In_451);
or U1156 (N_1156,In_725,In_803);
nor U1157 (N_1157,In_791,In_698);
nor U1158 (N_1158,In_14,In_35);
and U1159 (N_1159,In_845,In_412);
and U1160 (N_1160,In_58,In_713);
and U1161 (N_1161,In_818,In_454);
or U1162 (N_1162,In_237,In_284);
nor U1163 (N_1163,In_66,In_249);
xnor U1164 (N_1164,In_377,In_156);
and U1165 (N_1165,In_277,In_994);
or U1166 (N_1166,In_829,In_974);
nand U1167 (N_1167,In_178,In_374);
nand U1168 (N_1168,In_377,In_633);
nor U1169 (N_1169,In_911,In_339);
nand U1170 (N_1170,In_163,In_918);
and U1171 (N_1171,In_279,In_737);
and U1172 (N_1172,In_947,In_61);
or U1173 (N_1173,In_681,In_863);
or U1174 (N_1174,In_509,In_953);
nand U1175 (N_1175,In_762,In_40);
nand U1176 (N_1176,In_537,In_146);
nor U1177 (N_1177,In_531,In_829);
nor U1178 (N_1178,In_864,In_72);
or U1179 (N_1179,In_764,In_879);
nand U1180 (N_1180,In_42,In_663);
nor U1181 (N_1181,In_145,In_984);
or U1182 (N_1182,In_191,In_980);
nand U1183 (N_1183,In_88,In_330);
nor U1184 (N_1184,In_879,In_21);
xnor U1185 (N_1185,In_853,In_244);
nor U1186 (N_1186,In_134,In_809);
or U1187 (N_1187,In_243,In_529);
nand U1188 (N_1188,In_724,In_630);
or U1189 (N_1189,In_688,In_94);
nor U1190 (N_1190,In_885,In_227);
nor U1191 (N_1191,In_874,In_863);
nand U1192 (N_1192,In_930,In_188);
or U1193 (N_1193,In_317,In_575);
nand U1194 (N_1194,In_495,In_713);
or U1195 (N_1195,In_660,In_626);
nor U1196 (N_1196,In_267,In_752);
and U1197 (N_1197,In_263,In_240);
or U1198 (N_1198,In_180,In_623);
or U1199 (N_1199,In_740,In_275);
and U1200 (N_1200,In_695,In_266);
or U1201 (N_1201,In_721,In_683);
and U1202 (N_1202,In_999,In_119);
nand U1203 (N_1203,In_962,In_252);
nand U1204 (N_1204,In_765,In_31);
or U1205 (N_1205,In_910,In_353);
nor U1206 (N_1206,In_324,In_177);
nor U1207 (N_1207,In_418,In_667);
and U1208 (N_1208,In_36,In_920);
or U1209 (N_1209,In_133,In_429);
nand U1210 (N_1210,In_288,In_449);
or U1211 (N_1211,In_409,In_737);
nor U1212 (N_1212,In_637,In_739);
or U1213 (N_1213,In_115,In_187);
or U1214 (N_1214,In_736,In_436);
and U1215 (N_1215,In_993,In_861);
and U1216 (N_1216,In_984,In_139);
nor U1217 (N_1217,In_676,In_428);
and U1218 (N_1218,In_760,In_279);
or U1219 (N_1219,In_821,In_723);
or U1220 (N_1220,In_508,In_405);
nor U1221 (N_1221,In_427,In_628);
or U1222 (N_1222,In_299,In_543);
nand U1223 (N_1223,In_569,In_1);
and U1224 (N_1224,In_109,In_55);
or U1225 (N_1225,In_62,In_79);
and U1226 (N_1226,In_26,In_859);
nand U1227 (N_1227,In_528,In_106);
nor U1228 (N_1228,In_531,In_295);
and U1229 (N_1229,In_292,In_458);
and U1230 (N_1230,In_608,In_262);
and U1231 (N_1231,In_470,In_548);
or U1232 (N_1232,In_939,In_571);
nor U1233 (N_1233,In_93,In_869);
and U1234 (N_1234,In_873,In_536);
or U1235 (N_1235,In_28,In_715);
and U1236 (N_1236,In_65,In_407);
nand U1237 (N_1237,In_972,In_562);
nand U1238 (N_1238,In_505,In_723);
nand U1239 (N_1239,In_252,In_303);
or U1240 (N_1240,In_47,In_718);
nor U1241 (N_1241,In_935,In_220);
nor U1242 (N_1242,In_264,In_375);
or U1243 (N_1243,In_976,In_687);
or U1244 (N_1244,In_919,In_309);
and U1245 (N_1245,In_1,In_41);
and U1246 (N_1246,In_795,In_875);
nand U1247 (N_1247,In_459,In_839);
nand U1248 (N_1248,In_848,In_863);
nor U1249 (N_1249,In_887,In_977);
or U1250 (N_1250,In_946,In_24);
nor U1251 (N_1251,In_858,In_661);
or U1252 (N_1252,In_404,In_632);
and U1253 (N_1253,In_111,In_163);
and U1254 (N_1254,In_459,In_110);
nand U1255 (N_1255,In_212,In_576);
nor U1256 (N_1256,In_262,In_997);
and U1257 (N_1257,In_938,In_967);
and U1258 (N_1258,In_194,In_596);
or U1259 (N_1259,In_327,In_328);
and U1260 (N_1260,In_909,In_124);
nand U1261 (N_1261,In_720,In_928);
and U1262 (N_1262,In_563,In_889);
and U1263 (N_1263,In_389,In_594);
nor U1264 (N_1264,In_880,In_711);
nand U1265 (N_1265,In_453,In_677);
nand U1266 (N_1266,In_411,In_170);
nand U1267 (N_1267,In_387,In_935);
nand U1268 (N_1268,In_422,In_66);
nand U1269 (N_1269,In_684,In_418);
or U1270 (N_1270,In_369,In_616);
and U1271 (N_1271,In_804,In_809);
or U1272 (N_1272,In_632,In_695);
or U1273 (N_1273,In_105,In_636);
or U1274 (N_1274,In_719,In_763);
or U1275 (N_1275,In_713,In_476);
nand U1276 (N_1276,In_676,In_177);
and U1277 (N_1277,In_231,In_387);
or U1278 (N_1278,In_711,In_698);
or U1279 (N_1279,In_759,In_635);
or U1280 (N_1280,In_496,In_729);
nand U1281 (N_1281,In_946,In_100);
or U1282 (N_1282,In_476,In_519);
or U1283 (N_1283,In_629,In_411);
and U1284 (N_1284,In_398,In_87);
or U1285 (N_1285,In_617,In_415);
xor U1286 (N_1286,In_181,In_113);
nor U1287 (N_1287,In_472,In_647);
or U1288 (N_1288,In_125,In_123);
and U1289 (N_1289,In_981,In_331);
and U1290 (N_1290,In_687,In_619);
or U1291 (N_1291,In_349,In_130);
nor U1292 (N_1292,In_418,In_482);
or U1293 (N_1293,In_316,In_502);
and U1294 (N_1294,In_851,In_399);
nor U1295 (N_1295,In_553,In_435);
and U1296 (N_1296,In_591,In_870);
and U1297 (N_1297,In_830,In_408);
or U1298 (N_1298,In_745,In_851);
nor U1299 (N_1299,In_14,In_611);
nor U1300 (N_1300,In_706,In_906);
or U1301 (N_1301,In_649,In_642);
and U1302 (N_1302,In_958,In_494);
or U1303 (N_1303,In_527,In_788);
nor U1304 (N_1304,In_381,In_622);
or U1305 (N_1305,In_340,In_806);
nand U1306 (N_1306,In_76,In_185);
and U1307 (N_1307,In_117,In_144);
nand U1308 (N_1308,In_534,In_320);
nor U1309 (N_1309,In_67,In_732);
nor U1310 (N_1310,In_529,In_419);
or U1311 (N_1311,In_848,In_548);
nor U1312 (N_1312,In_420,In_278);
nor U1313 (N_1313,In_98,In_95);
and U1314 (N_1314,In_291,In_603);
or U1315 (N_1315,In_879,In_487);
and U1316 (N_1316,In_325,In_713);
nand U1317 (N_1317,In_844,In_465);
and U1318 (N_1318,In_148,In_661);
nand U1319 (N_1319,In_31,In_609);
and U1320 (N_1320,In_662,In_505);
or U1321 (N_1321,In_222,In_82);
nand U1322 (N_1322,In_210,In_597);
and U1323 (N_1323,In_521,In_884);
nor U1324 (N_1324,In_62,In_738);
xor U1325 (N_1325,In_945,In_496);
or U1326 (N_1326,In_906,In_628);
nor U1327 (N_1327,In_401,In_909);
or U1328 (N_1328,In_761,In_610);
and U1329 (N_1329,In_632,In_821);
nor U1330 (N_1330,In_132,In_500);
and U1331 (N_1331,In_59,In_713);
or U1332 (N_1332,In_66,In_858);
or U1333 (N_1333,In_866,In_543);
xor U1334 (N_1334,In_2,In_648);
nor U1335 (N_1335,In_627,In_240);
nand U1336 (N_1336,In_404,In_877);
nor U1337 (N_1337,In_356,In_654);
or U1338 (N_1338,In_551,In_103);
nor U1339 (N_1339,In_389,In_435);
or U1340 (N_1340,In_709,In_872);
nor U1341 (N_1341,In_641,In_190);
nand U1342 (N_1342,In_742,In_95);
xor U1343 (N_1343,In_619,In_665);
or U1344 (N_1344,In_304,In_343);
nor U1345 (N_1345,In_181,In_976);
nor U1346 (N_1346,In_99,In_468);
and U1347 (N_1347,In_690,In_967);
xor U1348 (N_1348,In_922,In_774);
nor U1349 (N_1349,In_778,In_822);
nand U1350 (N_1350,In_571,In_729);
or U1351 (N_1351,In_540,In_560);
xor U1352 (N_1352,In_923,In_440);
nand U1353 (N_1353,In_573,In_35);
and U1354 (N_1354,In_316,In_109);
nor U1355 (N_1355,In_220,In_804);
and U1356 (N_1356,In_754,In_484);
and U1357 (N_1357,In_415,In_643);
nor U1358 (N_1358,In_411,In_952);
nor U1359 (N_1359,In_261,In_460);
or U1360 (N_1360,In_104,In_257);
nor U1361 (N_1361,In_231,In_491);
and U1362 (N_1362,In_445,In_893);
nand U1363 (N_1363,In_781,In_706);
nand U1364 (N_1364,In_779,In_560);
nand U1365 (N_1365,In_847,In_221);
or U1366 (N_1366,In_933,In_717);
nor U1367 (N_1367,In_156,In_265);
or U1368 (N_1368,In_92,In_655);
nand U1369 (N_1369,In_198,In_234);
nand U1370 (N_1370,In_174,In_120);
or U1371 (N_1371,In_521,In_165);
nor U1372 (N_1372,In_559,In_59);
nor U1373 (N_1373,In_39,In_77);
nor U1374 (N_1374,In_555,In_64);
nand U1375 (N_1375,In_871,In_420);
and U1376 (N_1376,In_512,In_992);
nand U1377 (N_1377,In_297,In_7);
nor U1378 (N_1378,In_791,In_215);
nand U1379 (N_1379,In_90,In_234);
or U1380 (N_1380,In_60,In_879);
and U1381 (N_1381,In_421,In_143);
and U1382 (N_1382,In_58,In_620);
nor U1383 (N_1383,In_133,In_477);
or U1384 (N_1384,In_34,In_206);
and U1385 (N_1385,In_830,In_93);
nor U1386 (N_1386,In_987,In_627);
and U1387 (N_1387,In_370,In_171);
xnor U1388 (N_1388,In_347,In_369);
or U1389 (N_1389,In_593,In_938);
nand U1390 (N_1390,In_894,In_115);
or U1391 (N_1391,In_261,In_997);
nand U1392 (N_1392,In_289,In_601);
nor U1393 (N_1393,In_268,In_724);
and U1394 (N_1394,In_231,In_503);
nand U1395 (N_1395,In_893,In_514);
and U1396 (N_1396,In_181,In_957);
and U1397 (N_1397,In_174,In_542);
and U1398 (N_1398,In_420,In_661);
nor U1399 (N_1399,In_756,In_431);
nand U1400 (N_1400,In_981,In_940);
nor U1401 (N_1401,In_748,In_873);
or U1402 (N_1402,In_940,In_197);
nor U1403 (N_1403,In_854,In_929);
and U1404 (N_1404,In_745,In_514);
and U1405 (N_1405,In_505,In_186);
nor U1406 (N_1406,In_511,In_372);
nand U1407 (N_1407,In_281,In_977);
or U1408 (N_1408,In_905,In_144);
and U1409 (N_1409,In_343,In_949);
xor U1410 (N_1410,In_551,In_80);
and U1411 (N_1411,In_432,In_912);
nor U1412 (N_1412,In_411,In_485);
nand U1413 (N_1413,In_918,In_386);
and U1414 (N_1414,In_164,In_633);
and U1415 (N_1415,In_310,In_108);
xnor U1416 (N_1416,In_368,In_755);
or U1417 (N_1417,In_28,In_12);
nor U1418 (N_1418,In_972,In_163);
and U1419 (N_1419,In_364,In_242);
nor U1420 (N_1420,In_534,In_770);
or U1421 (N_1421,In_586,In_212);
nand U1422 (N_1422,In_626,In_543);
or U1423 (N_1423,In_924,In_105);
nand U1424 (N_1424,In_113,In_906);
or U1425 (N_1425,In_614,In_581);
or U1426 (N_1426,In_638,In_674);
nor U1427 (N_1427,In_651,In_947);
and U1428 (N_1428,In_52,In_534);
or U1429 (N_1429,In_420,In_579);
nand U1430 (N_1430,In_550,In_244);
and U1431 (N_1431,In_608,In_323);
nor U1432 (N_1432,In_507,In_135);
and U1433 (N_1433,In_468,In_578);
nor U1434 (N_1434,In_939,In_390);
nand U1435 (N_1435,In_125,In_715);
nand U1436 (N_1436,In_154,In_92);
or U1437 (N_1437,In_745,In_131);
nand U1438 (N_1438,In_523,In_305);
and U1439 (N_1439,In_546,In_941);
or U1440 (N_1440,In_906,In_406);
nand U1441 (N_1441,In_389,In_611);
nor U1442 (N_1442,In_557,In_554);
or U1443 (N_1443,In_779,In_745);
nand U1444 (N_1444,In_426,In_459);
and U1445 (N_1445,In_459,In_610);
or U1446 (N_1446,In_432,In_501);
or U1447 (N_1447,In_809,In_650);
nand U1448 (N_1448,In_713,In_395);
or U1449 (N_1449,In_407,In_832);
nor U1450 (N_1450,In_923,In_213);
and U1451 (N_1451,In_146,In_354);
nor U1452 (N_1452,In_794,In_425);
or U1453 (N_1453,In_912,In_723);
or U1454 (N_1454,In_412,In_171);
nand U1455 (N_1455,In_340,In_194);
or U1456 (N_1456,In_692,In_414);
xnor U1457 (N_1457,In_72,In_796);
or U1458 (N_1458,In_415,In_934);
or U1459 (N_1459,In_391,In_838);
or U1460 (N_1460,In_546,In_307);
nor U1461 (N_1461,In_797,In_330);
or U1462 (N_1462,In_7,In_796);
nor U1463 (N_1463,In_115,In_443);
nor U1464 (N_1464,In_524,In_140);
nor U1465 (N_1465,In_907,In_888);
nand U1466 (N_1466,In_97,In_550);
or U1467 (N_1467,In_487,In_707);
nor U1468 (N_1468,In_939,In_503);
nor U1469 (N_1469,In_159,In_607);
and U1470 (N_1470,In_268,In_759);
or U1471 (N_1471,In_36,In_650);
nor U1472 (N_1472,In_977,In_479);
or U1473 (N_1473,In_302,In_415);
and U1474 (N_1474,In_235,In_666);
nand U1475 (N_1475,In_551,In_647);
nor U1476 (N_1476,In_398,In_467);
and U1477 (N_1477,In_17,In_111);
or U1478 (N_1478,In_211,In_831);
nand U1479 (N_1479,In_95,In_402);
or U1480 (N_1480,In_552,In_559);
or U1481 (N_1481,In_124,In_542);
xnor U1482 (N_1482,In_969,In_266);
nor U1483 (N_1483,In_464,In_546);
nand U1484 (N_1484,In_464,In_701);
nand U1485 (N_1485,In_177,In_13);
nand U1486 (N_1486,In_745,In_658);
or U1487 (N_1487,In_923,In_750);
or U1488 (N_1488,In_352,In_177);
and U1489 (N_1489,In_258,In_932);
nor U1490 (N_1490,In_354,In_897);
or U1491 (N_1491,In_918,In_180);
nor U1492 (N_1492,In_827,In_72);
nand U1493 (N_1493,In_2,In_575);
nor U1494 (N_1494,In_739,In_632);
nand U1495 (N_1495,In_930,In_711);
and U1496 (N_1496,In_206,In_490);
or U1497 (N_1497,In_177,In_138);
nor U1498 (N_1498,In_442,In_295);
nor U1499 (N_1499,In_723,In_706);
or U1500 (N_1500,In_35,In_800);
and U1501 (N_1501,In_92,In_466);
nand U1502 (N_1502,In_649,In_187);
and U1503 (N_1503,In_223,In_528);
and U1504 (N_1504,In_994,In_511);
nand U1505 (N_1505,In_75,In_444);
or U1506 (N_1506,In_658,In_814);
nand U1507 (N_1507,In_583,In_752);
and U1508 (N_1508,In_387,In_287);
nand U1509 (N_1509,In_453,In_492);
nand U1510 (N_1510,In_679,In_646);
nor U1511 (N_1511,In_754,In_64);
or U1512 (N_1512,In_987,In_522);
nand U1513 (N_1513,In_699,In_808);
and U1514 (N_1514,In_679,In_34);
nor U1515 (N_1515,In_746,In_292);
nand U1516 (N_1516,In_774,In_543);
and U1517 (N_1517,In_252,In_733);
nand U1518 (N_1518,In_45,In_473);
nor U1519 (N_1519,In_545,In_281);
or U1520 (N_1520,In_27,In_641);
or U1521 (N_1521,In_672,In_667);
nand U1522 (N_1522,In_325,In_685);
nand U1523 (N_1523,In_818,In_591);
and U1524 (N_1524,In_699,In_149);
nor U1525 (N_1525,In_178,In_369);
or U1526 (N_1526,In_587,In_25);
or U1527 (N_1527,In_712,In_657);
nor U1528 (N_1528,In_821,In_845);
or U1529 (N_1529,In_838,In_99);
nor U1530 (N_1530,In_38,In_255);
nand U1531 (N_1531,In_689,In_708);
nor U1532 (N_1532,In_39,In_204);
nor U1533 (N_1533,In_558,In_426);
nor U1534 (N_1534,In_50,In_14);
and U1535 (N_1535,In_220,In_601);
nand U1536 (N_1536,In_877,In_399);
or U1537 (N_1537,In_352,In_588);
or U1538 (N_1538,In_493,In_607);
and U1539 (N_1539,In_196,In_833);
nor U1540 (N_1540,In_845,In_907);
nand U1541 (N_1541,In_438,In_177);
or U1542 (N_1542,In_445,In_717);
or U1543 (N_1543,In_363,In_36);
or U1544 (N_1544,In_238,In_757);
or U1545 (N_1545,In_466,In_1);
or U1546 (N_1546,In_896,In_274);
and U1547 (N_1547,In_106,In_998);
or U1548 (N_1548,In_687,In_290);
or U1549 (N_1549,In_238,In_94);
nand U1550 (N_1550,In_451,In_413);
nand U1551 (N_1551,In_667,In_616);
nor U1552 (N_1552,In_72,In_416);
or U1553 (N_1553,In_43,In_71);
nand U1554 (N_1554,In_911,In_292);
and U1555 (N_1555,In_528,In_181);
or U1556 (N_1556,In_621,In_457);
and U1557 (N_1557,In_594,In_978);
or U1558 (N_1558,In_306,In_716);
or U1559 (N_1559,In_618,In_455);
nor U1560 (N_1560,In_662,In_508);
and U1561 (N_1561,In_211,In_508);
nor U1562 (N_1562,In_533,In_337);
nand U1563 (N_1563,In_281,In_230);
or U1564 (N_1564,In_401,In_926);
xor U1565 (N_1565,In_468,In_775);
xor U1566 (N_1566,In_65,In_344);
or U1567 (N_1567,In_560,In_848);
nor U1568 (N_1568,In_609,In_175);
and U1569 (N_1569,In_103,In_701);
or U1570 (N_1570,In_475,In_522);
nor U1571 (N_1571,In_461,In_719);
and U1572 (N_1572,In_423,In_461);
nand U1573 (N_1573,In_774,In_416);
or U1574 (N_1574,In_473,In_242);
and U1575 (N_1575,In_167,In_514);
and U1576 (N_1576,In_108,In_54);
nor U1577 (N_1577,In_8,In_860);
nand U1578 (N_1578,In_854,In_363);
and U1579 (N_1579,In_776,In_570);
or U1580 (N_1580,In_741,In_730);
nand U1581 (N_1581,In_872,In_980);
or U1582 (N_1582,In_133,In_625);
and U1583 (N_1583,In_836,In_154);
and U1584 (N_1584,In_224,In_68);
nand U1585 (N_1585,In_70,In_731);
nand U1586 (N_1586,In_530,In_869);
nor U1587 (N_1587,In_382,In_347);
or U1588 (N_1588,In_979,In_983);
or U1589 (N_1589,In_834,In_736);
nand U1590 (N_1590,In_466,In_525);
nand U1591 (N_1591,In_719,In_756);
nor U1592 (N_1592,In_897,In_66);
nor U1593 (N_1593,In_709,In_492);
or U1594 (N_1594,In_74,In_310);
nand U1595 (N_1595,In_509,In_98);
nand U1596 (N_1596,In_683,In_725);
nor U1597 (N_1597,In_332,In_472);
nand U1598 (N_1598,In_204,In_127);
nor U1599 (N_1599,In_931,In_221);
or U1600 (N_1600,In_218,In_493);
xor U1601 (N_1601,In_393,In_603);
nor U1602 (N_1602,In_375,In_15);
nor U1603 (N_1603,In_707,In_95);
or U1604 (N_1604,In_664,In_307);
nor U1605 (N_1605,In_280,In_246);
nor U1606 (N_1606,In_650,In_568);
or U1607 (N_1607,In_419,In_79);
or U1608 (N_1608,In_577,In_266);
nand U1609 (N_1609,In_292,In_319);
nand U1610 (N_1610,In_134,In_987);
or U1611 (N_1611,In_724,In_969);
nand U1612 (N_1612,In_604,In_559);
nand U1613 (N_1613,In_591,In_54);
and U1614 (N_1614,In_625,In_638);
nor U1615 (N_1615,In_658,In_836);
nand U1616 (N_1616,In_534,In_637);
or U1617 (N_1617,In_213,In_829);
or U1618 (N_1618,In_541,In_977);
and U1619 (N_1619,In_20,In_817);
xor U1620 (N_1620,In_146,In_55);
or U1621 (N_1621,In_870,In_107);
nor U1622 (N_1622,In_357,In_349);
nand U1623 (N_1623,In_874,In_494);
nand U1624 (N_1624,In_262,In_790);
nand U1625 (N_1625,In_525,In_121);
nor U1626 (N_1626,In_570,In_259);
or U1627 (N_1627,In_517,In_716);
or U1628 (N_1628,In_373,In_183);
or U1629 (N_1629,In_343,In_788);
nand U1630 (N_1630,In_514,In_610);
xor U1631 (N_1631,In_59,In_612);
nand U1632 (N_1632,In_577,In_944);
and U1633 (N_1633,In_587,In_461);
and U1634 (N_1634,In_731,In_209);
nor U1635 (N_1635,In_102,In_459);
and U1636 (N_1636,In_155,In_181);
and U1637 (N_1637,In_465,In_364);
or U1638 (N_1638,In_110,In_875);
and U1639 (N_1639,In_488,In_832);
nor U1640 (N_1640,In_867,In_708);
nand U1641 (N_1641,In_266,In_455);
or U1642 (N_1642,In_265,In_849);
nand U1643 (N_1643,In_506,In_847);
and U1644 (N_1644,In_318,In_409);
nand U1645 (N_1645,In_149,In_588);
or U1646 (N_1646,In_530,In_177);
nor U1647 (N_1647,In_425,In_499);
nand U1648 (N_1648,In_635,In_349);
and U1649 (N_1649,In_863,In_6);
and U1650 (N_1650,In_981,In_136);
nor U1651 (N_1651,In_420,In_810);
or U1652 (N_1652,In_978,In_769);
and U1653 (N_1653,In_35,In_167);
or U1654 (N_1654,In_58,In_962);
or U1655 (N_1655,In_804,In_543);
and U1656 (N_1656,In_55,In_210);
and U1657 (N_1657,In_821,In_107);
nand U1658 (N_1658,In_916,In_3);
and U1659 (N_1659,In_521,In_979);
nor U1660 (N_1660,In_587,In_66);
nand U1661 (N_1661,In_967,In_616);
and U1662 (N_1662,In_358,In_824);
or U1663 (N_1663,In_69,In_662);
nor U1664 (N_1664,In_643,In_195);
and U1665 (N_1665,In_650,In_87);
or U1666 (N_1666,In_852,In_47);
or U1667 (N_1667,In_380,In_827);
nor U1668 (N_1668,In_626,In_565);
nand U1669 (N_1669,In_775,In_332);
nor U1670 (N_1670,In_927,In_234);
nand U1671 (N_1671,In_415,In_243);
nand U1672 (N_1672,In_580,In_747);
nand U1673 (N_1673,In_534,In_530);
nor U1674 (N_1674,In_676,In_90);
or U1675 (N_1675,In_197,In_512);
or U1676 (N_1676,In_157,In_692);
nand U1677 (N_1677,In_295,In_392);
nor U1678 (N_1678,In_97,In_292);
nor U1679 (N_1679,In_531,In_243);
nand U1680 (N_1680,In_612,In_448);
nand U1681 (N_1681,In_827,In_183);
nor U1682 (N_1682,In_43,In_400);
nand U1683 (N_1683,In_695,In_893);
nand U1684 (N_1684,In_0,In_905);
and U1685 (N_1685,In_622,In_165);
nand U1686 (N_1686,In_442,In_765);
or U1687 (N_1687,In_623,In_869);
nand U1688 (N_1688,In_426,In_387);
nand U1689 (N_1689,In_251,In_25);
or U1690 (N_1690,In_451,In_686);
nor U1691 (N_1691,In_863,In_815);
nand U1692 (N_1692,In_702,In_146);
xor U1693 (N_1693,In_185,In_974);
and U1694 (N_1694,In_767,In_572);
or U1695 (N_1695,In_958,In_766);
nand U1696 (N_1696,In_880,In_151);
xor U1697 (N_1697,In_986,In_366);
or U1698 (N_1698,In_752,In_869);
and U1699 (N_1699,In_755,In_729);
or U1700 (N_1700,In_291,In_932);
nand U1701 (N_1701,In_821,In_648);
nand U1702 (N_1702,In_420,In_116);
and U1703 (N_1703,In_902,In_921);
and U1704 (N_1704,In_18,In_425);
nand U1705 (N_1705,In_368,In_345);
or U1706 (N_1706,In_859,In_766);
nor U1707 (N_1707,In_364,In_309);
and U1708 (N_1708,In_309,In_359);
nand U1709 (N_1709,In_410,In_871);
nor U1710 (N_1710,In_863,In_903);
nand U1711 (N_1711,In_919,In_854);
and U1712 (N_1712,In_983,In_17);
and U1713 (N_1713,In_345,In_643);
and U1714 (N_1714,In_534,In_940);
nand U1715 (N_1715,In_244,In_767);
nor U1716 (N_1716,In_757,In_185);
or U1717 (N_1717,In_429,In_106);
nand U1718 (N_1718,In_419,In_734);
and U1719 (N_1719,In_141,In_547);
or U1720 (N_1720,In_717,In_33);
nor U1721 (N_1721,In_172,In_639);
nand U1722 (N_1722,In_226,In_129);
and U1723 (N_1723,In_926,In_856);
or U1724 (N_1724,In_732,In_7);
xor U1725 (N_1725,In_715,In_176);
nor U1726 (N_1726,In_66,In_870);
nand U1727 (N_1727,In_922,In_838);
and U1728 (N_1728,In_103,In_338);
nand U1729 (N_1729,In_198,In_202);
and U1730 (N_1730,In_601,In_6);
nand U1731 (N_1731,In_279,In_852);
xnor U1732 (N_1732,In_836,In_238);
or U1733 (N_1733,In_457,In_220);
nor U1734 (N_1734,In_488,In_507);
and U1735 (N_1735,In_567,In_437);
nand U1736 (N_1736,In_566,In_558);
nor U1737 (N_1737,In_58,In_465);
and U1738 (N_1738,In_882,In_384);
nor U1739 (N_1739,In_822,In_295);
or U1740 (N_1740,In_177,In_632);
and U1741 (N_1741,In_283,In_139);
nor U1742 (N_1742,In_80,In_895);
or U1743 (N_1743,In_684,In_81);
nor U1744 (N_1744,In_539,In_81);
or U1745 (N_1745,In_649,In_147);
and U1746 (N_1746,In_296,In_981);
or U1747 (N_1747,In_979,In_152);
and U1748 (N_1748,In_423,In_670);
and U1749 (N_1749,In_848,In_2);
nor U1750 (N_1750,In_282,In_108);
xnor U1751 (N_1751,In_358,In_647);
nand U1752 (N_1752,In_725,In_862);
nand U1753 (N_1753,In_619,In_823);
or U1754 (N_1754,In_604,In_745);
and U1755 (N_1755,In_125,In_85);
nor U1756 (N_1756,In_807,In_304);
xnor U1757 (N_1757,In_87,In_704);
and U1758 (N_1758,In_37,In_730);
nor U1759 (N_1759,In_715,In_217);
nand U1760 (N_1760,In_354,In_621);
nand U1761 (N_1761,In_722,In_418);
nor U1762 (N_1762,In_295,In_849);
and U1763 (N_1763,In_170,In_561);
nor U1764 (N_1764,In_508,In_177);
and U1765 (N_1765,In_280,In_965);
nor U1766 (N_1766,In_763,In_564);
nor U1767 (N_1767,In_704,In_487);
and U1768 (N_1768,In_820,In_916);
or U1769 (N_1769,In_42,In_474);
nand U1770 (N_1770,In_775,In_415);
nor U1771 (N_1771,In_611,In_733);
nor U1772 (N_1772,In_922,In_143);
nor U1773 (N_1773,In_466,In_682);
and U1774 (N_1774,In_180,In_748);
and U1775 (N_1775,In_329,In_378);
nor U1776 (N_1776,In_496,In_134);
nand U1777 (N_1777,In_615,In_579);
nand U1778 (N_1778,In_302,In_341);
nand U1779 (N_1779,In_535,In_218);
and U1780 (N_1780,In_834,In_698);
nand U1781 (N_1781,In_634,In_683);
or U1782 (N_1782,In_798,In_56);
nand U1783 (N_1783,In_74,In_460);
and U1784 (N_1784,In_267,In_400);
nor U1785 (N_1785,In_79,In_34);
nand U1786 (N_1786,In_336,In_372);
nand U1787 (N_1787,In_797,In_863);
and U1788 (N_1788,In_929,In_85);
nor U1789 (N_1789,In_690,In_824);
xnor U1790 (N_1790,In_995,In_251);
nand U1791 (N_1791,In_499,In_30);
nand U1792 (N_1792,In_410,In_264);
nand U1793 (N_1793,In_623,In_754);
nand U1794 (N_1794,In_72,In_569);
nand U1795 (N_1795,In_437,In_442);
and U1796 (N_1796,In_357,In_443);
xnor U1797 (N_1797,In_252,In_459);
nand U1798 (N_1798,In_656,In_315);
nor U1799 (N_1799,In_54,In_15);
nand U1800 (N_1800,In_974,In_476);
or U1801 (N_1801,In_323,In_42);
and U1802 (N_1802,In_834,In_43);
nor U1803 (N_1803,In_751,In_444);
or U1804 (N_1804,In_982,In_936);
or U1805 (N_1805,In_516,In_968);
and U1806 (N_1806,In_931,In_784);
nor U1807 (N_1807,In_567,In_800);
nand U1808 (N_1808,In_323,In_328);
or U1809 (N_1809,In_118,In_356);
nor U1810 (N_1810,In_30,In_88);
and U1811 (N_1811,In_588,In_783);
or U1812 (N_1812,In_111,In_295);
or U1813 (N_1813,In_268,In_273);
or U1814 (N_1814,In_521,In_469);
and U1815 (N_1815,In_647,In_65);
nand U1816 (N_1816,In_928,In_414);
and U1817 (N_1817,In_126,In_950);
nand U1818 (N_1818,In_676,In_589);
and U1819 (N_1819,In_528,In_905);
and U1820 (N_1820,In_627,In_507);
nand U1821 (N_1821,In_373,In_396);
nand U1822 (N_1822,In_44,In_255);
nor U1823 (N_1823,In_439,In_11);
nand U1824 (N_1824,In_207,In_237);
or U1825 (N_1825,In_765,In_662);
or U1826 (N_1826,In_640,In_374);
nand U1827 (N_1827,In_678,In_444);
or U1828 (N_1828,In_382,In_56);
nor U1829 (N_1829,In_897,In_560);
nand U1830 (N_1830,In_384,In_985);
nor U1831 (N_1831,In_204,In_417);
nor U1832 (N_1832,In_362,In_198);
nor U1833 (N_1833,In_662,In_506);
nand U1834 (N_1834,In_261,In_420);
nand U1835 (N_1835,In_223,In_288);
and U1836 (N_1836,In_49,In_773);
and U1837 (N_1837,In_84,In_276);
nand U1838 (N_1838,In_380,In_239);
and U1839 (N_1839,In_991,In_701);
nor U1840 (N_1840,In_792,In_124);
or U1841 (N_1841,In_255,In_67);
or U1842 (N_1842,In_615,In_631);
and U1843 (N_1843,In_118,In_0);
and U1844 (N_1844,In_727,In_531);
or U1845 (N_1845,In_725,In_672);
nand U1846 (N_1846,In_357,In_175);
or U1847 (N_1847,In_678,In_880);
nand U1848 (N_1848,In_211,In_203);
and U1849 (N_1849,In_1,In_798);
nor U1850 (N_1850,In_509,In_326);
and U1851 (N_1851,In_74,In_433);
and U1852 (N_1852,In_670,In_280);
xor U1853 (N_1853,In_113,In_705);
nand U1854 (N_1854,In_285,In_275);
nand U1855 (N_1855,In_266,In_789);
nand U1856 (N_1856,In_661,In_98);
nor U1857 (N_1857,In_981,In_351);
or U1858 (N_1858,In_330,In_381);
nor U1859 (N_1859,In_895,In_759);
xnor U1860 (N_1860,In_69,In_373);
and U1861 (N_1861,In_544,In_89);
nand U1862 (N_1862,In_13,In_755);
nand U1863 (N_1863,In_226,In_836);
or U1864 (N_1864,In_27,In_600);
or U1865 (N_1865,In_755,In_70);
nor U1866 (N_1866,In_938,In_383);
nor U1867 (N_1867,In_425,In_854);
and U1868 (N_1868,In_496,In_561);
or U1869 (N_1869,In_924,In_444);
nor U1870 (N_1870,In_689,In_930);
nand U1871 (N_1871,In_626,In_915);
nor U1872 (N_1872,In_238,In_214);
and U1873 (N_1873,In_432,In_762);
nor U1874 (N_1874,In_680,In_109);
or U1875 (N_1875,In_182,In_625);
nand U1876 (N_1876,In_354,In_532);
xnor U1877 (N_1877,In_603,In_986);
nor U1878 (N_1878,In_607,In_76);
nand U1879 (N_1879,In_157,In_644);
nand U1880 (N_1880,In_455,In_57);
nor U1881 (N_1881,In_594,In_833);
or U1882 (N_1882,In_233,In_625);
nor U1883 (N_1883,In_608,In_133);
nor U1884 (N_1884,In_557,In_416);
nor U1885 (N_1885,In_246,In_129);
nor U1886 (N_1886,In_818,In_157);
nand U1887 (N_1887,In_841,In_301);
or U1888 (N_1888,In_681,In_420);
nor U1889 (N_1889,In_597,In_962);
and U1890 (N_1890,In_984,In_278);
nand U1891 (N_1891,In_459,In_607);
nor U1892 (N_1892,In_581,In_739);
nand U1893 (N_1893,In_270,In_550);
and U1894 (N_1894,In_186,In_813);
nand U1895 (N_1895,In_538,In_861);
nor U1896 (N_1896,In_408,In_382);
nand U1897 (N_1897,In_620,In_175);
nand U1898 (N_1898,In_619,In_521);
nor U1899 (N_1899,In_616,In_864);
or U1900 (N_1900,In_513,In_559);
nor U1901 (N_1901,In_635,In_237);
or U1902 (N_1902,In_797,In_326);
nor U1903 (N_1903,In_94,In_903);
nand U1904 (N_1904,In_447,In_393);
and U1905 (N_1905,In_987,In_195);
and U1906 (N_1906,In_57,In_595);
and U1907 (N_1907,In_686,In_983);
or U1908 (N_1908,In_42,In_48);
nor U1909 (N_1909,In_916,In_284);
nand U1910 (N_1910,In_316,In_939);
and U1911 (N_1911,In_807,In_722);
or U1912 (N_1912,In_369,In_389);
nor U1913 (N_1913,In_985,In_299);
or U1914 (N_1914,In_8,In_636);
nor U1915 (N_1915,In_351,In_183);
nand U1916 (N_1916,In_994,In_825);
or U1917 (N_1917,In_687,In_464);
or U1918 (N_1918,In_365,In_565);
or U1919 (N_1919,In_709,In_530);
nor U1920 (N_1920,In_5,In_660);
or U1921 (N_1921,In_990,In_510);
or U1922 (N_1922,In_935,In_754);
or U1923 (N_1923,In_687,In_591);
nand U1924 (N_1924,In_920,In_901);
or U1925 (N_1925,In_725,In_971);
or U1926 (N_1926,In_897,In_724);
or U1927 (N_1927,In_127,In_120);
nand U1928 (N_1928,In_632,In_444);
nand U1929 (N_1929,In_371,In_440);
or U1930 (N_1930,In_672,In_59);
nor U1931 (N_1931,In_735,In_264);
nor U1932 (N_1932,In_195,In_162);
nand U1933 (N_1933,In_120,In_700);
nor U1934 (N_1934,In_250,In_712);
nand U1935 (N_1935,In_769,In_875);
xnor U1936 (N_1936,In_890,In_966);
nand U1937 (N_1937,In_411,In_578);
nand U1938 (N_1938,In_952,In_816);
or U1939 (N_1939,In_325,In_243);
and U1940 (N_1940,In_50,In_818);
nand U1941 (N_1941,In_47,In_574);
xnor U1942 (N_1942,In_499,In_627);
nand U1943 (N_1943,In_601,In_39);
nor U1944 (N_1944,In_274,In_789);
nor U1945 (N_1945,In_469,In_13);
nand U1946 (N_1946,In_721,In_549);
nor U1947 (N_1947,In_597,In_202);
and U1948 (N_1948,In_392,In_86);
and U1949 (N_1949,In_585,In_997);
nor U1950 (N_1950,In_860,In_762);
nor U1951 (N_1951,In_645,In_603);
nand U1952 (N_1952,In_412,In_457);
or U1953 (N_1953,In_986,In_592);
nand U1954 (N_1954,In_294,In_16);
nor U1955 (N_1955,In_365,In_768);
or U1956 (N_1956,In_815,In_730);
or U1957 (N_1957,In_204,In_497);
or U1958 (N_1958,In_21,In_465);
and U1959 (N_1959,In_67,In_259);
and U1960 (N_1960,In_466,In_452);
nor U1961 (N_1961,In_177,In_32);
or U1962 (N_1962,In_427,In_613);
nor U1963 (N_1963,In_636,In_935);
or U1964 (N_1964,In_374,In_122);
and U1965 (N_1965,In_481,In_328);
or U1966 (N_1966,In_973,In_843);
nor U1967 (N_1967,In_978,In_839);
nand U1968 (N_1968,In_523,In_194);
nand U1969 (N_1969,In_102,In_719);
nor U1970 (N_1970,In_398,In_478);
nor U1971 (N_1971,In_182,In_930);
and U1972 (N_1972,In_83,In_133);
nand U1973 (N_1973,In_786,In_941);
or U1974 (N_1974,In_115,In_614);
nor U1975 (N_1975,In_859,In_582);
or U1976 (N_1976,In_282,In_872);
nand U1977 (N_1977,In_932,In_264);
nor U1978 (N_1978,In_0,In_89);
and U1979 (N_1979,In_459,In_393);
and U1980 (N_1980,In_247,In_760);
nor U1981 (N_1981,In_788,In_666);
or U1982 (N_1982,In_741,In_148);
or U1983 (N_1983,In_137,In_387);
nand U1984 (N_1984,In_906,In_776);
nor U1985 (N_1985,In_191,In_740);
nand U1986 (N_1986,In_994,In_711);
nand U1987 (N_1987,In_113,In_30);
or U1988 (N_1988,In_630,In_772);
and U1989 (N_1989,In_215,In_445);
xor U1990 (N_1990,In_148,In_57);
nand U1991 (N_1991,In_872,In_802);
nor U1992 (N_1992,In_673,In_727);
nor U1993 (N_1993,In_427,In_740);
and U1994 (N_1994,In_445,In_304);
and U1995 (N_1995,In_695,In_982);
nand U1996 (N_1996,In_654,In_843);
and U1997 (N_1997,In_683,In_22);
nor U1998 (N_1998,In_612,In_249);
and U1999 (N_1999,In_970,In_931);
nand U2000 (N_2000,In_520,In_424);
nor U2001 (N_2001,In_163,In_893);
nand U2002 (N_2002,In_678,In_689);
nand U2003 (N_2003,In_668,In_903);
nor U2004 (N_2004,In_724,In_597);
nand U2005 (N_2005,In_45,In_563);
nor U2006 (N_2006,In_809,In_318);
or U2007 (N_2007,In_99,In_635);
nor U2008 (N_2008,In_225,In_17);
and U2009 (N_2009,In_927,In_715);
nand U2010 (N_2010,In_995,In_740);
or U2011 (N_2011,In_59,In_580);
xnor U2012 (N_2012,In_539,In_819);
and U2013 (N_2013,In_469,In_216);
nor U2014 (N_2014,In_693,In_114);
nand U2015 (N_2015,In_590,In_825);
and U2016 (N_2016,In_657,In_919);
or U2017 (N_2017,In_336,In_889);
nand U2018 (N_2018,In_229,In_961);
or U2019 (N_2019,In_191,In_277);
nor U2020 (N_2020,In_292,In_962);
nand U2021 (N_2021,In_803,In_141);
and U2022 (N_2022,In_931,In_540);
xnor U2023 (N_2023,In_758,In_76);
xor U2024 (N_2024,In_350,In_863);
nand U2025 (N_2025,In_811,In_353);
nor U2026 (N_2026,In_612,In_892);
nand U2027 (N_2027,In_937,In_779);
nand U2028 (N_2028,In_608,In_949);
nor U2029 (N_2029,In_93,In_238);
and U2030 (N_2030,In_460,In_134);
nand U2031 (N_2031,In_834,In_474);
nor U2032 (N_2032,In_191,In_473);
or U2033 (N_2033,In_483,In_528);
or U2034 (N_2034,In_484,In_629);
xor U2035 (N_2035,In_459,In_873);
or U2036 (N_2036,In_495,In_26);
or U2037 (N_2037,In_111,In_507);
xnor U2038 (N_2038,In_709,In_412);
nand U2039 (N_2039,In_356,In_936);
or U2040 (N_2040,In_401,In_0);
and U2041 (N_2041,In_585,In_284);
and U2042 (N_2042,In_248,In_353);
and U2043 (N_2043,In_633,In_878);
or U2044 (N_2044,In_396,In_541);
and U2045 (N_2045,In_890,In_839);
and U2046 (N_2046,In_614,In_313);
or U2047 (N_2047,In_988,In_485);
or U2048 (N_2048,In_926,In_928);
xnor U2049 (N_2049,In_456,In_254);
nand U2050 (N_2050,In_233,In_907);
or U2051 (N_2051,In_650,In_80);
or U2052 (N_2052,In_18,In_416);
nor U2053 (N_2053,In_272,In_157);
and U2054 (N_2054,In_584,In_238);
or U2055 (N_2055,In_532,In_879);
or U2056 (N_2056,In_533,In_101);
or U2057 (N_2057,In_686,In_599);
nor U2058 (N_2058,In_152,In_685);
and U2059 (N_2059,In_969,In_382);
and U2060 (N_2060,In_446,In_971);
nand U2061 (N_2061,In_53,In_48);
or U2062 (N_2062,In_161,In_126);
nor U2063 (N_2063,In_722,In_986);
nand U2064 (N_2064,In_770,In_934);
and U2065 (N_2065,In_383,In_32);
nand U2066 (N_2066,In_470,In_762);
nor U2067 (N_2067,In_303,In_500);
or U2068 (N_2068,In_342,In_271);
nand U2069 (N_2069,In_617,In_785);
and U2070 (N_2070,In_457,In_774);
or U2071 (N_2071,In_442,In_130);
nor U2072 (N_2072,In_377,In_483);
and U2073 (N_2073,In_628,In_543);
nand U2074 (N_2074,In_982,In_586);
nand U2075 (N_2075,In_372,In_263);
or U2076 (N_2076,In_121,In_993);
and U2077 (N_2077,In_847,In_197);
nand U2078 (N_2078,In_958,In_61);
nand U2079 (N_2079,In_539,In_483);
or U2080 (N_2080,In_204,In_314);
or U2081 (N_2081,In_406,In_569);
nand U2082 (N_2082,In_347,In_494);
and U2083 (N_2083,In_846,In_527);
nand U2084 (N_2084,In_832,In_121);
and U2085 (N_2085,In_73,In_214);
nor U2086 (N_2086,In_906,In_713);
nor U2087 (N_2087,In_484,In_281);
nor U2088 (N_2088,In_747,In_516);
and U2089 (N_2089,In_237,In_598);
nor U2090 (N_2090,In_545,In_339);
nor U2091 (N_2091,In_631,In_481);
nor U2092 (N_2092,In_616,In_971);
and U2093 (N_2093,In_987,In_744);
and U2094 (N_2094,In_46,In_716);
nand U2095 (N_2095,In_680,In_961);
nand U2096 (N_2096,In_93,In_578);
nor U2097 (N_2097,In_995,In_715);
or U2098 (N_2098,In_670,In_340);
nand U2099 (N_2099,In_314,In_655);
nor U2100 (N_2100,In_242,In_337);
nand U2101 (N_2101,In_93,In_237);
or U2102 (N_2102,In_696,In_105);
and U2103 (N_2103,In_511,In_388);
and U2104 (N_2104,In_419,In_373);
nor U2105 (N_2105,In_380,In_401);
and U2106 (N_2106,In_795,In_587);
nand U2107 (N_2107,In_828,In_642);
xnor U2108 (N_2108,In_885,In_440);
nand U2109 (N_2109,In_853,In_831);
and U2110 (N_2110,In_339,In_937);
xor U2111 (N_2111,In_162,In_100);
nand U2112 (N_2112,In_406,In_462);
nor U2113 (N_2113,In_348,In_255);
or U2114 (N_2114,In_578,In_487);
nor U2115 (N_2115,In_181,In_512);
nand U2116 (N_2116,In_849,In_710);
nand U2117 (N_2117,In_333,In_433);
xnor U2118 (N_2118,In_342,In_862);
or U2119 (N_2119,In_748,In_355);
or U2120 (N_2120,In_96,In_146);
nor U2121 (N_2121,In_998,In_253);
nand U2122 (N_2122,In_995,In_812);
nor U2123 (N_2123,In_175,In_826);
nand U2124 (N_2124,In_28,In_880);
nand U2125 (N_2125,In_400,In_955);
nand U2126 (N_2126,In_25,In_943);
or U2127 (N_2127,In_995,In_612);
nor U2128 (N_2128,In_121,In_684);
nand U2129 (N_2129,In_431,In_492);
and U2130 (N_2130,In_413,In_210);
or U2131 (N_2131,In_488,In_181);
and U2132 (N_2132,In_306,In_159);
xor U2133 (N_2133,In_366,In_242);
or U2134 (N_2134,In_164,In_133);
and U2135 (N_2135,In_575,In_455);
nand U2136 (N_2136,In_489,In_240);
and U2137 (N_2137,In_518,In_240);
and U2138 (N_2138,In_960,In_35);
or U2139 (N_2139,In_604,In_820);
nor U2140 (N_2140,In_579,In_905);
or U2141 (N_2141,In_735,In_674);
nand U2142 (N_2142,In_634,In_279);
nand U2143 (N_2143,In_612,In_725);
nand U2144 (N_2144,In_63,In_358);
nand U2145 (N_2145,In_80,In_586);
or U2146 (N_2146,In_846,In_131);
and U2147 (N_2147,In_569,In_877);
nand U2148 (N_2148,In_63,In_800);
xor U2149 (N_2149,In_359,In_74);
or U2150 (N_2150,In_303,In_536);
or U2151 (N_2151,In_980,In_471);
nand U2152 (N_2152,In_7,In_956);
nor U2153 (N_2153,In_81,In_555);
nand U2154 (N_2154,In_720,In_964);
nand U2155 (N_2155,In_556,In_94);
nand U2156 (N_2156,In_124,In_351);
and U2157 (N_2157,In_950,In_396);
and U2158 (N_2158,In_666,In_568);
nor U2159 (N_2159,In_887,In_540);
and U2160 (N_2160,In_179,In_356);
or U2161 (N_2161,In_346,In_362);
xnor U2162 (N_2162,In_179,In_236);
or U2163 (N_2163,In_411,In_265);
xor U2164 (N_2164,In_62,In_1);
or U2165 (N_2165,In_39,In_470);
and U2166 (N_2166,In_791,In_12);
nand U2167 (N_2167,In_737,In_431);
and U2168 (N_2168,In_664,In_375);
and U2169 (N_2169,In_647,In_642);
nor U2170 (N_2170,In_114,In_335);
or U2171 (N_2171,In_703,In_141);
nor U2172 (N_2172,In_332,In_361);
nand U2173 (N_2173,In_22,In_682);
nor U2174 (N_2174,In_516,In_361);
xor U2175 (N_2175,In_630,In_319);
nor U2176 (N_2176,In_396,In_765);
nor U2177 (N_2177,In_688,In_54);
nor U2178 (N_2178,In_194,In_617);
nor U2179 (N_2179,In_326,In_655);
and U2180 (N_2180,In_661,In_359);
nor U2181 (N_2181,In_206,In_408);
nand U2182 (N_2182,In_96,In_856);
nor U2183 (N_2183,In_151,In_94);
nand U2184 (N_2184,In_922,In_974);
nor U2185 (N_2185,In_657,In_203);
or U2186 (N_2186,In_513,In_341);
nand U2187 (N_2187,In_313,In_297);
nor U2188 (N_2188,In_896,In_211);
nand U2189 (N_2189,In_373,In_799);
or U2190 (N_2190,In_270,In_360);
nor U2191 (N_2191,In_351,In_969);
or U2192 (N_2192,In_982,In_279);
or U2193 (N_2193,In_146,In_412);
nor U2194 (N_2194,In_773,In_384);
or U2195 (N_2195,In_422,In_950);
nor U2196 (N_2196,In_642,In_922);
and U2197 (N_2197,In_64,In_338);
or U2198 (N_2198,In_204,In_877);
or U2199 (N_2199,In_899,In_353);
and U2200 (N_2200,In_273,In_470);
nor U2201 (N_2201,In_102,In_733);
nor U2202 (N_2202,In_67,In_376);
nor U2203 (N_2203,In_331,In_48);
and U2204 (N_2204,In_678,In_340);
nor U2205 (N_2205,In_230,In_872);
nand U2206 (N_2206,In_368,In_262);
nand U2207 (N_2207,In_167,In_352);
and U2208 (N_2208,In_863,In_235);
nand U2209 (N_2209,In_170,In_363);
and U2210 (N_2210,In_703,In_675);
or U2211 (N_2211,In_568,In_939);
nor U2212 (N_2212,In_947,In_244);
and U2213 (N_2213,In_447,In_445);
and U2214 (N_2214,In_499,In_571);
nor U2215 (N_2215,In_239,In_650);
nand U2216 (N_2216,In_213,In_426);
and U2217 (N_2217,In_924,In_492);
nand U2218 (N_2218,In_600,In_895);
nor U2219 (N_2219,In_160,In_581);
and U2220 (N_2220,In_620,In_780);
and U2221 (N_2221,In_451,In_229);
or U2222 (N_2222,In_585,In_488);
nand U2223 (N_2223,In_765,In_6);
and U2224 (N_2224,In_930,In_172);
or U2225 (N_2225,In_276,In_423);
nand U2226 (N_2226,In_330,In_491);
or U2227 (N_2227,In_678,In_828);
or U2228 (N_2228,In_680,In_657);
nand U2229 (N_2229,In_618,In_107);
xor U2230 (N_2230,In_826,In_611);
nand U2231 (N_2231,In_861,In_655);
xor U2232 (N_2232,In_91,In_519);
or U2233 (N_2233,In_151,In_331);
or U2234 (N_2234,In_678,In_334);
nor U2235 (N_2235,In_516,In_524);
nor U2236 (N_2236,In_688,In_370);
nor U2237 (N_2237,In_943,In_23);
nand U2238 (N_2238,In_827,In_600);
nand U2239 (N_2239,In_998,In_649);
nor U2240 (N_2240,In_555,In_773);
xnor U2241 (N_2241,In_47,In_526);
nand U2242 (N_2242,In_923,In_575);
nand U2243 (N_2243,In_113,In_921);
and U2244 (N_2244,In_588,In_958);
nor U2245 (N_2245,In_449,In_712);
and U2246 (N_2246,In_952,In_414);
and U2247 (N_2247,In_268,In_359);
or U2248 (N_2248,In_558,In_199);
and U2249 (N_2249,In_587,In_814);
nor U2250 (N_2250,In_138,In_171);
or U2251 (N_2251,In_987,In_961);
or U2252 (N_2252,In_230,In_314);
nand U2253 (N_2253,In_882,In_380);
nand U2254 (N_2254,In_522,In_573);
nand U2255 (N_2255,In_159,In_12);
nor U2256 (N_2256,In_599,In_461);
nand U2257 (N_2257,In_169,In_417);
and U2258 (N_2258,In_325,In_58);
and U2259 (N_2259,In_232,In_346);
or U2260 (N_2260,In_988,In_624);
nor U2261 (N_2261,In_514,In_202);
nand U2262 (N_2262,In_7,In_843);
xor U2263 (N_2263,In_141,In_121);
xnor U2264 (N_2264,In_506,In_540);
and U2265 (N_2265,In_112,In_979);
nor U2266 (N_2266,In_537,In_965);
nor U2267 (N_2267,In_434,In_750);
or U2268 (N_2268,In_917,In_957);
nor U2269 (N_2269,In_297,In_21);
nor U2270 (N_2270,In_999,In_897);
and U2271 (N_2271,In_293,In_146);
nand U2272 (N_2272,In_976,In_324);
or U2273 (N_2273,In_930,In_651);
or U2274 (N_2274,In_819,In_186);
nand U2275 (N_2275,In_42,In_386);
xor U2276 (N_2276,In_251,In_782);
and U2277 (N_2277,In_133,In_236);
nand U2278 (N_2278,In_103,In_29);
nor U2279 (N_2279,In_904,In_192);
nor U2280 (N_2280,In_266,In_925);
or U2281 (N_2281,In_280,In_465);
or U2282 (N_2282,In_803,In_899);
or U2283 (N_2283,In_903,In_743);
nor U2284 (N_2284,In_894,In_40);
and U2285 (N_2285,In_786,In_283);
nand U2286 (N_2286,In_223,In_543);
or U2287 (N_2287,In_860,In_839);
nor U2288 (N_2288,In_530,In_996);
or U2289 (N_2289,In_322,In_310);
and U2290 (N_2290,In_445,In_312);
nand U2291 (N_2291,In_94,In_802);
and U2292 (N_2292,In_290,In_819);
nand U2293 (N_2293,In_71,In_747);
nor U2294 (N_2294,In_859,In_312);
and U2295 (N_2295,In_10,In_785);
or U2296 (N_2296,In_821,In_233);
or U2297 (N_2297,In_468,In_712);
nor U2298 (N_2298,In_913,In_117);
nor U2299 (N_2299,In_833,In_437);
or U2300 (N_2300,In_561,In_611);
or U2301 (N_2301,In_517,In_343);
or U2302 (N_2302,In_150,In_913);
or U2303 (N_2303,In_830,In_2);
nor U2304 (N_2304,In_471,In_391);
and U2305 (N_2305,In_373,In_367);
or U2306 (N_2306,In_581,In_35);
or U2307 (N_2307,In_484,In_526);
and U2308 (N_2308,In_408,In_900);
xnor U2309 (N_2309,In_952,In_712);
xnor U2310 (N_2310,In_189,In_13);
and U2311 (N_2311,In_538,In_940);
and U2312 (N_2312,In_670,In_306);
nand U2313 (N_2313,In_761,In_726);
or U2314 (N_2314,In_113,In_340);
or U2315 (N_2315,In_483,In_209);
nand U2316 (N_2316,In_827,In_640);
nand U2317 (N_2317,In_359,In_715);
nand U2318 (N_2318,In_235,In_552);
or U2319 (N_2319,In_128,In_510);
or U2320 (N_2320,In_435,In_100);
and U2321 (N_2321,In_531,In_953);
and U2322 (N_2322,In_336,In_175);
or U2323 (N_2323,In_641,In_942);
or U2324 (N_2324,In_636,In_889);
nand U2325 (N_2325,In_544,In_951);
or U2326 (N_2326,In_428,In_928);
or U2327 (N_2327,In_477,In_809);
nand U2328 (N_2328,In_415,In_266);
and U2329 (N_2329,In_674,In_765);
nor U2330 (N_2330,In_61,In_857);
nor U2331 (N_2331,In_389,In_112);
or U2332 (N_2332,In_595,In_147);
or U2333 (N_2333,In_694,In_540);
nor U2334 (N_2334,In_585,In_131);
nand U2335 (N_2335,In_638,In_472);
nor U2336 (N_2336,In_436,In_326);
and U2337 (N_2337,In_464,In_422);
and U2338 (N_2338,In_630,In_632);
nor U2339 (N_2339,In_524,In_681);
nand U2340 (N_2340,In_218,In_576);
nor U2341 (N_2341,In_525,In_53);
nand U2342 (N_2342,In_886,In_847);
and U2343 (N_2343,In_771,In_288);
nand U2344 (N_2344,In_356,In_792);
or U2345 (N_2345,In_868,In_490);
and U2346 (N_2346,In_753,In_793);
nor U2347 (N_2347,In_498,In_59);
nand U2348 (N_2348,In_289,In_789);
nor U2349 (N_2349,In_172,In_893);
nor U2350 (N_2350,In_971,In_151);
nand U2351 (N_2351,In_518,In_8);
and U2352 (N_2352,In_327,In_275);
and U2353 (N_2353,In_307,In_998);
and U2354 (N_2354,In_539,In_43);
nand U2355 (N_2355,In_174,In_489);
nand U2356 (N_2356,In_206,In_810);
nand U2357 (N_2357,In_605,In_839);
nand U2358 (N_2358,In_281,In_127);
or U2359 (N_2359,In_692,In_844);
or U2360 (N_2360,In_88,In_350);
nor U2361 (N_2361,In_605,In_131);
nor U2362 (N_2362,In_321,In_77);
and U2363 (N_2363,In_355,In_890);
xor U2364 (N_2364,In_203,In_10);
nand U2365 (N_2365,In_842,In_408);
and U2366 (N_2366,In_522,In_565);
and U2367 (N_2367,In_7,In_920);
nor U2368 (N_2368,In_418,In_702);
and U2369 (N_2369,In_145,In_294);
and U2370 (N_2370,In_416,In_869);
nor U2371 (N_2371,In_132,In_307);
and U2372 (N_2372,In_972,In_457);
nand U2373 (N_2373,In_456,In_887);
or U2374 (N_2374,In_369,In_151);
nor U2375 (N_2375,In_295,In_936);
nand U2376 (N_2376,In_951,In_600);
and U2377 (N_2377,In_988,In_909);
nor U2378 (N_2378,In_393,In_965);
nand U2379 (N_2379,In_507,In_193);
nand U2380 (N_2380,In_916,In_210);
nor U2381 (N_2381,In_314,In_547);
or U2382 (N_2382,In_88,In_931);
and U2383 (N_2383,In_674,In_841);
nor U2384 (N_2384,In_10,In_316);
nand U2385 (N_2385,In_871,In_611);
nor U2386 (N_2386,In_462,In_621);
and U2387 (N_2387,In_653,In_496);
nand U2388 (N_2388,In_729,In_935);
xnor U2389 (N_2389,In_90,In_248);
and U2390 (N_2390,In_746,In_693);
nand U2391 (N_2391,In_565,In_341);
and U2392 (N_2392,In_367,In_161);
and U2393 (N_2393,In_983,In_334);
nor U2394 (N_2394,In_559,In_393);
and U2395 (N_2395,In_297,In_633);
nor U2396 (N_2396,In_715,In_691);
or U2397 (N_2397,In_126,In_374);
nand U2398 (N_2398,In_874,In_985);
or U2399 (N_2399,In_198,In_921);
nand U2400 (N_2400,In_654,In_925);
nand U2401 (N_2401,In_981,In_830);
xnor U2402 (N_2402,In_826,In_30);
nor U2403 (N_2403,In_671,In_694);
nor U2404 (N_2404,In_859,In_675);
nand U2405 (N_2405,In_151,In_74);
and U2406 (N_2406,In_972,In_309);
and U2407 (N_2407,In_517,In_190);
nand U2408 (N_2408,In_620,In_658);
and U2409 (N_2409,In_271,In_469);
or U2410 (N_2410,In_772,In_566);
nand U2411 (N_2411,In_88,In_742);
nor U2412 (N_2412,In_620,In_177);
or U2413 (N_2413,In_521,In_439);
or U2414 (N_2414,In_89,In_72);
and U2415 (N_2415,In_592,In_707);
nand U2416 (N_2416,In_352,In_771);
or U2417 (N_2417,In_520,In_470);
and U2418 (N_2418,In_524,In_250);
xor U2419 (N_2419,In_936,In_53);
or U2420 (N_2420,In_71,In_193);
nand U2421 (N_2421,In_109,In_803);
and U2422 (N_2422,In_586,In_339);
nor U2423 (N_2423,In_953,In_680);
or U2424 (N_2424,In_600,In_681);
or U2425 (N_2425,In_380,In_980);
or U2426 (N_2426,In_131,In_44);
xor U2427 (N_2427,In_421,In_110);
nor U2428 (N_2428,In_524,In_329);
nor U2429 (N_2429,In_518,In_683);
and U2430 (N_2430,In_138,In_731);
or U2431 (N_2431,In_81,In_465);
and U2432 (N_2432,In_315,In_505);
nor U2433 (N_2433,In_498,In_812);
or U2434 (N_2434,In_324,In_566);
nor U2435 (N_2435,In_663,In_365);
nor U2436 (N_2436,In_429,In_806);
nand U2437 (N_2437,In_247,In_245);
nand U2438 (N_2438,In_616,In_334);
or U2439 (N_2439,In_560,In_662);
nor U2440 (N_2440,In_89,In_26);
nor U2441 (N_2441,In_905,In_349);
nand U2442 (N_2442,In_480,In_16);
xnor U2443 (N_2443,In_812,In_155);
nand U2444 (N_2444,In_121,In_532);
or U2445 (N_2445,In_327,In_535);
and U2446 (N_2446,In_423,In_753);
nand U2447 (N_2447,In_484,In_855);
or U2448 (N_2448,In_874,In_236);
or U2449 (N_2449,In_172,In_316);
nand U2450 (N_2450,In_950,In_556);
nand U2451 (N_2451,In_510,In_517);
nand U2452 (N_2452,In_530,In_278);
or U2453 (N_2453,In_688,In_891);
nand U2454 (N_2454,In_304,In_669);
nor U2455 (N_2455,In_864,In_23);
or U2456 (N_2456,In_823,In_881);
or U2457 (N_2457,In_504,In_147);
or U2458 (N_2458,In_319,In_222);
nand U2459 (N_2459,In_872,In_436);
nor U2460 (N_2460,In_570,In_114);
nand U2461 (N_2461,In_436,In_284);
or U2462 (N_2462,In_238,In_174);
and U2463 (N_2463,In_868,In_493);
and U2464 (N_2464,In_995,In_268);
nor U2465 (N_2465,In_355,In_523);
nor U2466 (N_2466,In_39,In_292);
or U2467 (N_2467,In_528,In_393);
or U2468 (N_2468,In_452,In_651);
nor U2469 (N_2469,In_29,In_919);
and U2470 (N_2470,In_63,In_982);
nand U2471 (N_2471,In_854,In_645);
and U2472 (N_2472,In_294,In_595);
nand U2473 (N_2473,In_352,In_975);
and U2474 (N_2474,In_581,In_552);
or U2475 (N_2475,In_273,In_664);
or U2476 (N_2476,In_695,In_890);
or U2477 (N_2477,In_921,In_39);
xnor U2478 (N_2478,In_914,In_84);
nand U2479 (N_2479,In_166,In_381);
nand U2480 (N_2480,In_559,In_962);
or U2481 (N_2481,In_892,In_388);
or U2482 (N_2482,In_360,In_319);
and U2483 (N_2483,In_686,In_58);
or U2484 (N_2484,In_911,In_163);
and U2485 (N_2485,In_438,In_779);
nor U2486 (N_2486,In_945,In_602);
nor U2487 (N_2487,In_74,In_364);
nand U2488 (N_2488,In_256,In_149);
and U2489 (N_2489,In_949,In_898);
nand U2490 (N_2490,In_178,In_175);
nand U2491 (N_2491,In_331,In_420);
or U2492 (N_2492,In_941,In_810);
and U2493 (N_2493,In_411,In_556);
xnor U2494 (N_2494,In_71,In_890);
nand U2495 (N_2495,In_674,In_422);
and U2496 (N_2496,In_911,In_979);
and U2497 (N_2497,In_668,In_842);
nand U2498 (N_2498,In_16,In_213);
and U2499 (N_2499,In_53,In_548);
nand U2500 (N_2500,N_1399,N_1749);
and U2501 (N_2501,N_644,N_27);
or U2502 (N_2502,N_1750,N_2042);
or U2503 (N_2503,N_1932,N_336);
nor U2504 (N_2504,N_1313,N_927);
and U2505 (N_2505,N_1733,N_678);
or U2506 (N_2506,N_379,N_1753);
nand U2507 (N_2507,N_495,N_2493);
and U2508 (N_2508,N_1772,N_797);
nand U2509 (N_2509,N_1017,N_1494);
nor U2510 (N_2510,N_1964,N_610);
nand U2511 (N_2511,N_974,N_1216);
and U2512 (N_2512,N_2110,N_1090);
nor U2513 (N_2513,N_1995,N_2212);
and U2514 (N_2514,N_1320,N_2028);
nor U2515 (N_2515,N_1481,N_1261);
nand U2516 (N_2516,N_554,N_1621);
xnor U2517 (N_2517,N_2352,N_1583);
nor U2518 (N_2518,N_41,N_980);
or U2519 (N_2519,N_194,N_31);
and U2520 (N_2520,N_711,N_1896);
nor U2521 (N_2521,N_988,N_1400);
or U2522 (N_2522,N_71,N_629);
and U2523 (N_2523,N_206,N_1291);
nand U2524 (N_2524,N_6,N_1435);
nor U2525 (N_2525,N_1385,N_2410);
nor U2526 (N_2526,N_640,N_1821);
nor U2527 (N_2527,N_2209,N_1093);
and U2528 (N_2528,N_1800,N_1546);
nand U2529 (N_2529,N_2418,N_1049);
nand U2530 (N_2530,N_1149,N_2302);
or U2531 (N_2531,N_1115,N_933);
nor U2532 (N_2532,N_1707,N_484);
nand U2533 (N_2533,N_734,N_885);
or U2534 (N_2534,N_96,N_2463);
nand U2535 (N_2535,N_2051,N_287);
or U2536 (N_2536,N_305,N_1949);
nor U2537 (N_2537,N_2424,N_462);
nand U2538 (N_2538,N_246,N_1104);
and U2539 (N_2539,N_1831,N_685);
and U2540 (N_2540,N_1010,N_1730);
nor U2541 (N_2541,N_2007,N_2133);
and U2542 (N_2542,N_929,N_1680);
nand U2543 (N_2543,N_45,N_1563);
and U2544 (N_2544,N_370,N_1798);
or U2545 (N_2545,N_1445,N_1705);
nor U2546 (N_2546,N_16,N_924);
or U2547 (N_2547,N_73,N_2091);
nand U2548 (N_2548,N_1453,N_1604);
or U2549 (N_2549,N_2019,N_344);
xor U2550 (N_2550,N_1542,N_91);
nand U2551 (N_2551,N_2322,N_777);
nand U2552 (N_2552,N_532,N_870);
nand U2553 (N_2553,N_319,N_2126);
or U2554 (N_2554,N_1638,N_1071);
nand U2555 (N_2555,N_2130,N_730);
xor U2556 (N_2556,N_848,N_941);
and U2557 (N_2557,N_205,N_1260);
nand U2558 (N_2558,N_2282,N_742);
or U2559 (N_2559,N_1308,N_641);
and U2560 (N_2560,N_1030,N_1124);
nor U2561 (N_2561,N_1819,N_1833);
and U2562 (N_2562,N_2297,N_1020);
nor U2563 (N_2563,N_787,N_167);
and U2564 (N_2564,N_1930,N_850);
or U2565 (N_2565,N_1897,N_512);
xor U2566 (N_2566,N_224,N_1443);
nand U2567 (N_2567,N_2176,N_146);
nor U2568 (N_2568,N_211,N_2279);
or U2569 (N_2569,N_266,N_2129);
nor U2570 (N_2570,N_52,N_2086);
nor U2571 (N_2571,N_338,N_2256);
nor U2572 (N_2572,N_243,N_350);
nand U2573 (N_2573,N_1160,N_1170);
or U2574 (N_2574,N_2355,N_2470);
or U2575 (N_2575,N_355,N_2219);
nor U2576 (N_2576,N_1161,N_949);
and U2577 (N_2577,N_446,N_1468);
nor U2578 (N_2578,N_2085,N_1687);
nand U2579 (N_2579,N_653,N_1873);
or U2580 (N_2580,N_21,N_1770);
nor U2581 (N_2581,N_1200,N_2047);
or U2582 (N_2582,N_1685,N_1540);
and U2583 (N_2583,N_5,N_2494);
or U2584 (N_2584,N_799,N_1719);
nand U2585 (N_2585,N_986,N_544);
and U2586 (N_2586,N_886,N_1289);
or U2587 (N_2587,N_1278,N_1573);
nor U2588 (N_2588,N_1398,N_625);
nor U2589 (N_2589,N_755,N_584);
and U2590 (N_2590,N_839,N_2266);
nor U2591 (N_2591,N_2365,N_1073);
nand U2592 (N_2592,N_1033,N_2068);
nand U2593 (N_2593,N_1001,N_694);
nand U2594 (N_2594,N_1585,N_390);
nand U2595 (N_2595,N_2095,N_2181);
nand U2596 (N_2596,N_1817,N_461);
and U2597 (N_2597,N_1850,N_2313);
or U2598 (N_2598,N_1698,N_2314);
or U2599 (N_2599,N_1013,N_971);
or U2600 (N_2600,N_1900,N_523);
nor U2601 (N_2601,N_505,N_1862);
nand U2602 (N_2602,N_814,N_1467);
nand U2603 (N_2603,N_1598,N_2066);
nand U2604 (N_2604,N_857,N_160);
and U2605 (N_2605,N_1763,N_811);
or U2606 (N_2606,N_1401,N_1882);
or U2607 (N_2607,N_1275,N_1927);
nor U2608 (N_2608,N_1496,N_910);
nor U2609 (N_2609,N_624,N_1866);
nor U2610 (N_2610,N_1381,N_2063);
or U2611 (N_2611,N_2407,N_547);
and U2612 (N_2612,N_1759,N_2213);
nand U2613 (N_2613,N_1863,N_1709);
nand U2614 (N_2614,N_1852,N_903);
nand U2615 (N_2615,N_828,N_1653);
nand U2616 (N_2616,N_558,N_1986);
nor U2617 (N_2617,N_227,N_1777);
nand U2618 (N_2618,N_413,N_2391);
xnor U2619 (N_2619,N_1661,N_743);
nand U2620 (N_2620,N_1396,N_2469);
or U2621 (N_2621,N_1213,N_2408);
and U2622 (N_2622,N_3,N_1879);
and U2623 (N_2623,N_470,N_645);
and U2624 (N_2624,N_1951,N_765);
nand U2625 (N_2625,N_1574,N_1148);
nand U2626 (N_2626,N_1439,N_1710);
nor U2627 (N_2627,N_485,N_578);
xor U2628 (N_2628,N_511,N_2482);
nor U2629 (N_2629,N_76,N_487);
or U2630 (N_2630,N_185,N_1713);
nor U2631 (N_2631,N_2439,N_654);
or U2632 (N_2632,N_1189,N_1885);
or U2633 (N_2633,N_2191,N_2197);
nor U2634 (N_2634,N_771,N_915);
and U2635 (N_2635,N_1605,N_2056);
nand U2636 (N_2636,N_934,N_1910);
and U2637 (N_2637,N_976,N_1279);
nand U2638 (N_2638,N_2349,N_1110);
nor U2639 (N_2639,N_2048,N_1519);
or U2640 (N_2640,N_2427,N_782);
nor U2641 (N_2641,N_136,N_2433);
nor U2642 (N_2642,N_169,N_100);
or U2643 (N_2643,N_1446,N_1393);
or U2644 (N_2644,N_595,N_1190);
or U2645 (N_2645,N_1024,N_662);
and U2646 (N_2646,N_399,N_911);
or U2647 (N_2647,N_1309,N_1361);
nor U2648 (N_2648,N_1069,N_853);
xnor U2649 (N_2649,N_1530,N_868);
nand U2650 (N_2650,N_141,N_535);
nand U2651 (N_2651,N_623,N_2320);
and U2652 (N_2652,N_739,N_435);
and U2653 (N_2653,N_877,N_2000);
nor U2654 (N_2654,N_2026,N_2165);
nor U2655 (N_2655,N_1383,N_1217);
and U2656 (N_2656,N_1622,N_230);
or U2657 (N_2657,N_1688,N_530);
and U2658 (N_2658,N_1324,N_1990);
nor U2659 (N_2659,N_1694,N_1700);
nand U2660 (N_2660,N_1732,N_2190);
and U2661 (N_2661,N_1240,N_2477);
and U2662 (N_2662,N_1989,N_1007);
nand U2663 (N_2663,N_424,N_175);
nand U2664 (N_2664,N_2226,N_1886);
or U2665 (N_2665,N_1871,N_1146);
nand U2666 (N_2666,N_1357,N_2127);
or U2667 (N_2667,N_529,N_833);
nor U2668 (N_2668,N_2441,N_1738);
nand U2669 (N_2669,N_1414,N_199);
nand U2670 (N_2670,N_1697,N_153);
nand U2671 (N_2671,N_113,N_501);
nand U2672 (N_2672,N_674,N_2224);
or U2673 (N_2673,N_513,N_2174);
xnor U2674 (N_2674,N_1619,N_2199);
or U2675 (N_2675,N_2031,N_1230);
or U2676 (N_2676,N_1838,N_1181);
and U2677 (N_2677,N_1865,N_1918);
nor U2678 (N_2678,N_975,N_611);
or U2679 (N_2679,N_187,N_481);
or U2680 (N_2680,N_1447,N_809);
or U2681 (N_2681,N_551,N_2332);
nand U2682 (N_2682,N_1462,N_1239);
nand U2683 (N_2683,N_2220,N_94);
nand U2684 (N_2684,N_506,N_1814);
nand U2685 (N_2685,N_83,N_2317);
nand U2686 (N_2686,N_1174,N_1977);
nand U2687 (N_2687,N_478,N_323);
nand U2688 (N_2688,N_1282,N_1677);
nand U2689 (N_2689,N_790,N_362);
nor U2690 (N_2690,N_1911,N_38);
and U2691 (N_2691,N_1529,N_1437);
nand U2692 (N_2692,N_722,N_1089);
nor U2693 (N_2693,N_202,N_1665);
nand U2694 (N_2694,N_880,N_2497);
nand U2695 (N_2695,N_2468,N_1009);
nor U2696 (N_2696,N_143,N_774);
nor U2697 (N_2697,N_940,N_1664);
nor U2698 (N_2698,N_1133,N_670);
nor U2699 (N_2699,N_208,N_364);
or U2700 (N_2700,N_841,N_1371);
and U2701 (N_2701,N_1011,N_2318);
nor U2702 (N_2702,N_1080,N_631);
or U2703 (N_2703,N_2040,N_1087);
and U2704 (N_2704,N_1431,N_673);
nand U2705 (N_2705,N_1974,N_166);
nor U2706 (N_2706,N_846,N_84);
and U2707 (N_2707,N_895,N_1899);
and U2708 (N_2708,N_1497,N_2443);
xnor U2709 (N_2709,N_322,N_50);
nor U2710 (N_2710,N_1163,N_1512);
nand U2711 (N_2711,N_109,N_842);
nor U2712 (N_2712,N_1648,N_486);
and U2713 (N_2713,N_1894,N_1614);
nand U2714 (N_2714,N_1222,N_1718);
or U2715 (N_2715,N_2276,N_1557);
nor U2716 (N_2716,N_1799,N_2389);
nor U2717 (N_2717,N_1413,N_1156);
or U2718 (N_2718,N_80,N_803);
and U2719 (N_2719,N_1252,N_1144);
nand U2720 (N_2720,N_302,N_689);
or U2721 (N_2721,N_984,N_79);
nand U2722 (N_2722,N_213,N_2461);
nand U2723 (N_2723,N_66,N_560);
and U2724 (N_2724,N_2360,N_1064);
or U2725 (N_2725,N_2221,N_447);
nand U2726 (N_2726,N_994,N_28);
nand U2727 (N_2727,N_1739,N_1241);
and U2728 (N_2728,N_1600,N_460);
nor U2729 (N_2729,N_1844,N_2094);
or U2730 (N_2730,N_1187,N_2310);
nor U2731 (N_2731,N_1036,N_1996);
nor U2732 (N_2732,N_1450,N_1491);
xor U2733 (N_2733,N_1097,N_327);
and U2734 (N_2734,N_1048,N_1988);
nor U2735 (N_2735,N_1803,N_417);
nor U2736 (N_2736,N_2359,N_1926);
and U2737 (N_2737,N_1441,N_1545);
and U2738 (N_2738,N_1589,N_807);
nor U2739 (N_2739,N_1026,N_217);
and U2740 (N_2740,N_1418,N_236);
nor U2741 (N_2741,N_437,N_90);
nand U2742 (N_2742,N_1292,N_878);
nor U2743 (N_2743,N_25,N_65);
or U2744 (N_2744,N_2,N_1535);
and U2745 (N_2745,N_2392,N_1508);
nand U2746 (N_2746,N_691,N_1165);
and U2747 (N_2747,N_749,N_1562);
or U2748 (N_2748,N_2305,N_2012);
nor U2749 (N_2749,N_310,N_2278);
nor U2750 (N_2750,N_1262,N_144);
nor U2751 (N_2751,N_2351,N_705);
or U2752 (N_2752,N_545,N_1483);
and U2753 (N_2753,N_1768,N_1084);
nor U2754 (N_2754,N_7,N_2434);
nor U2755 (N_2755,N_104,N_521);
and U2756 (N_2756,N_2444,N_1220);
and U2757 (N_2757,N_188,N_2152);
or U2758 (N_2758,N_690,N_2018);
nand U2759 (N_2759,N_2373,N_132);
nand U2760 (N_2760,N_262,N_650);
nand U2761 (N_2761,N_527,N_1267);
nor U2762 (N_2762,N_1776,N_464);
and U2763 (N_2763,N_1587,N_411);
nor U2764 (N_2764,N_1055,N_2016);
nand U2765 (N_2765,N_1105,N_655);
nand U2766 (N_2766,N_1311,N_2009);
nor U2767 (N_2767,N_140,N_1281);
nor U2768 (N_2768,N_2123,N_456);
or U2769 (N_2769,N_2485,N_1586);
and U2770 (N_2770,N_1797,N_1625);
nor U2771 (N_2771,N_125,N_982);
nand U2772 (N_2772,N_232,N_2015);
or U2773 (N_2773,N_23,N_427);
and U2774 (N_2774,N_843,N_46);
nor U2775 (N_2775,N_1635,N_769);
nor U2776 (N_2776,N_1360,N_1569);
and U2777 (N_2777,N_873,N_55);
and U2778 (N_2778,N_1000,N_215);
or U2779 (N_2779,N_2036,N_1319);
or U2780 (N_2780,N_747,N_1054);
or U2781 (N_2781,N_2264,N_395);
nand U2782 (N_2782,N_2372,N_1100);
or U2783 (N_2783,N_946,N_1303);
and U2784 (N_2784,N_1404,N_865);
nor U2785 (N_2785,N_533,N_756);
and U2786 (N_2786,N_1344,N_2073);
xnor U2787 (N_2787,N_767,N_1537);
or U2788 (N_2788,N_441,N_1188);
xnor U2789 (N_2789,N_1917,N_1715);
nand U2790 (N_2790,N_1226,N_274);
or U2791 (N_2791,N_1488,N_930);
or U2792 (N_2792,N_1538,N_420);
or U2793 (N_2793,N_1597,N_366);
or U2794 (N_2794,N_2092,N_706);
or U2795 (N_2795,N_1966,N_1847);
and U2796 (N_2796,N_235,N_2106);
nand U2797 (N_2797,N_2013,N_884);
nor U2798 (N_2798,N_2452,N_1933);
nor U2799 (N_2799,N_2377,N_1744);
nand U2800 (N_2800,N_352,N_1352);
and U2801 (N_2801,N_1370,N_837);
nand U2802 (N_2802,N_913,N_1382);
nand U2803 (N_2803,N_1518,N_1666);
and U2804 (N_2804,N_1720,N_1826);
and U2805 (N_2805,N_1526,N_2453);
nor U2806 (N_2806,N_1632,N_2416);
nand U2807 (N_2807,N_2148,N_2251);
and U2808 (N_2808,N_1539,N_661);
nand U2809 (N_2809,N_1658,N_93);
and U2810 (N_2810,N_1489,N_860);
and U2811 (N_2811,N_737,N_316);
nor U2812 (N_2812,N_1214,N_497);
nor U2813 (N_2813,N_1015,N_1994);
or U2814 (N_2814,N_159,N_1890);
and U2815 (N_2815,N_1845,N_2055);
nand U2816 (N_2816,N_1972,N_1039);
nor U2817 (N_2817,N_2324,N_300);
nor U2818 (N_2818,N_1452,N_1854);
or U2819 (N_2819,N_701,N_114);
nor U2820 (N_2820,N_2159,N_2206);
or U2821 (N_2821,N_2033,N_207);
or U2822 (N_2822,N_1126,N_158);
xor U2823 (N_2823,N_134,N_105);
nand U2824 (N_2824,N_1829,N_736);
or U2825 (N_2825,N_1561,N_1329);
nand U2826 (N_2826,N_1460,N_1153);
and U2827 (N_2827,N_520,N_42);
and U2828 (N_2828,N_2411,N_1955);
and U2829 (N_2829,N_1760,N_1642);
and U2830 (N_2830,N_564,N_1078);
nand U2831 (N_2831,N_2300,N_938);
or U2832 (N_2832,N_110,N_469);
nand U2833 (N_2833,N_1456,N_703);
xnor U2834 (N_2834,N_1367,N_2406);
nor U2835 (N_2835,N_119,N_1005);
nor U2836 (N_2836,N_1629,N_1839);
or U2837 (N_2837,N_1334,N_2237);
nand U2838 (N_2838,N_2062,N_1679);
nand U2839 (N_2839,N_1458,N_311);
nand U2840 (N_2840,N_1463,N_1043);
and U2841 (N_2841,N_254,N_58);
and U2842 (N_2842,N_2017,N_612);
nand U2843 (N_2843,N_1433,N_1248);
or U2844 (N_2844,N_493,N_408);
xnor U2845 (N_2845,N_999,N_2379);
nand U2846 (N_2846,N_1081,N_1454);
and U2847 (N_2847,N_567,N_1108);
nand U2848 (N_2848,N_2089,N_2231);
or U2849 (N_2849,N_1276,N_952);
and U2850 (N_2850,N_222,N_1128);
or U2851 (N_2851,N_1063,N_1962);
nor U2852 (N_2852,N_2303,N_1236);
and U2853 (N_2853,N_1690,N_2491);
or U2854 (N_2854,N_707,N_2235);
nor U2855 (N_2855,N_2381,N_1476);
or U2856 (N_2856,N_1135,N_149);
and U2857 (N_2857,N_757,N_1581);
nor U2858 (N_2858,N_574,N_2362);
nor U2859 (N_2859,N_1502,N_808);
nand U2860 (N_2860,N_443,N_1256);
nor U2861 (N_2861,N_2478,N_2021);
and U2862 (N_2862,N_70,N_1416);
and U2863 (N_2863,N_2495,N_2339);
and U2864 (N_2864,N_223,N_360);
nor U2865 (N_2865,N_2401,N_1354);
nor U2866 (N_2866,N_154,N_590);
or U2867 (N_2867,N_192,N_648);
and U2868 (N_2868,N_2053,N_1869);
or U2869 (N_2869,N_1199,N_966);
and U2870 (N_2870,N_2080,N_412);
or U2871 (N_2871,N_238,N_463);
nand U2872 (N_2872,N_2312,N_375);
nand U2873 (N_2873,N_117,N_1116);
and U2874 (N_2874,N_1771,N_2204);
and U2875 (N_2875,N_1480,N_1014);
or U2876 (N_2876,N_1523,N_2208);
and U2877 (N_2877,N_2116,N_1608);
nor U2878 (N_2878,N_1390,N_1981);
nor U2879 (N_2879,N_1593,N_1335);
and U2880 (N_2880,N_1255,N_591);
and U2881 (N_2881,N_2459,N_9);
and U2882 (N_2882,N_1701,N_1902);
nand U2883 (N_2883,N_1492,N_917);
or U2884 (N_2884,N_387,N_1570);
nor U2885 (N_2885,N_2134,N_2088);
nor U2886 (N_2886,N_1599,N_700);
or U2887 (N_2887,N_203,N_1610);
nand U2888 (N_2888,N_2253,N_1347);
nor U2889 (N_2889,N_116,N_1221);
or U2890 (N_2890,N_1975,N_537);
and U2891 (N_2891,N_2409,N_918);
nor U2892 (N_2892,N_549,N_312);
nor U2893 (N_2893,N_32,N_2079);
nand U2894 (N_2894,N_1058,N_1656);
and U2895 (N_2895,N_19,N_921);
nand U2896 (N_2896,N_1544,N_2399);
or U2897 (N_2897,N_1633,N_1389);
nand U2898 (N_2898,N_2366,N_2143);
and U2899 (N_2899,N_1628,N_909);
or U2900 (N_2900,N_431,N_389);
nor U2901 (N_2901,N_252,N_219);
nand U2902 (N_2902,N_1645,N_728);
or U2903 (N_2903,N_1403,N_906);
nand U2904 (N_2904,N_2334,N_509);
nor U2905 (N_2905,N_22,N_1615);
xor U2906 (N_2906,N_400,N_1044);
and U2907 (N_2907,N_465,N_1554);
or U2908 (N_2908,N_2113,N_371);
or U2909 (N_2909,N_821,N_414);
or U2910 (N_2910,N_894,N_597);
nor U2911 (N_2911,N_635,N_1037);
and U2912 (N_2912,N_1059,N_482);
nor U2913 (N_2913,N_2456,N_1388);
nand U2914 (N_2914,N_2203,N_1423);
or U2915 (N_2915,N_2097,N_823);
or U2916 (N_2916,N_2071,N_2075);
and U2917 (N_2917,N_1692,N_75);
nor U2918 (N_2918,N_2150,N_594);
or U2919 (N_2919,N_1032,N_500);
nand U2920 (N_2920,N_1660,N_563);
nand U2921 (N_2921,N_1336,N_1259);
or U2922 (N_2922,N_2098,N_801);
nor U2923 (N_2923,N_1141,N_819);
or U2924 (N_2924,N_1411,N_951);
or U2925 (N_2925,N_643,N_359);
nor U2926 (N_2926,N_785,N_1725);
nand U2927 (N_2927,N_834,N_2388);
nand U2928 (N_2928,N_849,N_896);
nor U2929 (N_2929,N_1397,N_2122);
nand U2930 (N_2930,N_1689,N_1825);
nor U2931 (N_2931,N_1913,N_1325);
or U2932 (N_2932,N_1340,N_292);
nand U2933 (N_2933,N_376,N_2262);
nand U2934 (N_2934,N_1811,N_2440);
nor U2935 (N_2935,N_1410,N_1892);
nand U2936 (N_2936,N_2357,N_321);
nor U2937 (N_2937,N_1970,N_2210);
nand U2938 (N_2938,N_1379,N_2107);
or U2939 (N_2939,N_381,N_864);
or U2940 (N_2940,N_1751,N_1021);
or U2941 (N_2941,N_2222,N_1655);
nand U2942 (N_2942,N_2412,N_245);
and U2943 (N_2943,N_298,N_1843);
and U2944 (N_2944,N_11,N_1130);
and U2945 (N_2945,N_1764,N_1801);
or U2946 (N_2946,N_1806,N_1674);
nand U2947 (N_2947,N_768,N_1793);
nor U2948 (N_2948,N_18,N_72);
and U2949 (N_2949,N_1301,N_2064);
nand U2950 (N_2950,N_133,N_1006);
and U2951 (N_2951,N_2426,N_1673);
and U2952 (N_2952,N_577,N_1057);
or U2953 (N_2953,N_268,N_1306);
and U2954 (N_2954,N_1953,N_1369);
or U2955 (N_2955,N_244,N_363);
nand U2956 (N_2956,N_1830,N_1286);
nand U2957 (N_2957,N_1355,N_748);
nand U2958 (N_2958,N_313,N_139);
nor U2959 (N_2959,N_491,N_2138);
nand U2960 (N_2960,N_1515,N_618);
nand U2961 (N_2961,N_614,N_2230);
and U2962 (N_2962,N_812,N_829);
nand U2963 (N_2963,N_2387,N_2232);
nor U2964 (N_2964,N_525,N_1046);
or U2965 (N_2965,N_1901,N_677);
or U2966 (N_2966,N_1118,N_2299);
nor U2967 (N_2967,N_2192,N_1145);
nor U2968 (N_2968,N_800,N_723);
nand U2969 (N_2969,N_101,N_1867);
nand U2970 (N_2970,N_282,N_1266);
and U2971 (N_2971,N_1532,N_1099);
nor U2972 (N_2972,N_1138,N_2378);
nor U2973 (N_2973,N_422,N_1499);
nor U2974 (N_2974,N_155,N_216);
nand U2975 (N_2975,N_49,N_69);
xor U2976 (N_2976,N_288,N_426);
nor U2977 (N_2977,N_87,N_1113);
or U2978 (N_2978,N_514,N_1004);
nand U2979 (N_2979,N_546,N_679);
or U2980 (N_2980,N_220,N_1878);
nor U2981 (N_2981,N_442,N_2242);
nor U2982 (N_2982,N_2454,N_2155);
nor U2983 (N_2983,N_0,N_1726);
nand U2984 (N_2984,N_522,N_1455);
or U2985 (N_2985,N_1834,N_1272);
nand U2986 (N_2986,N_398,N_1012);
nor U2987 (N_2987,N_1315,N_369);
nand U2988 (N_2988,N_471,N_666);
nand U2989 (N_2989,N_480,N_2402);
and U2990 (N_2990,N_1824,N_2038);
xnor U2991 (N_2991,N_1094,N_1372);
nor U2992 (N_2992,N_2142,N_1157);
or U2993 (N_2993,N_664,N_1716);
nand U2994 (N_2994,N_1755,N_954);
or U2995 (N_2995,N_195,N_892);
or U2996 (N_2996,N_457,N_1415);
nand U2997 (N_2997,N_1940,N_1948);
nand U2998 (N_2998,N_1907,N_2309);
nor U2999 (N_2999,N_2457,N_1180);
nand U3000 (N_3000,N_762,N_620);
nand U3001 (N_3001,N_2321,N_490);
nor U3002 (N_3002,N_357,N_657);
nor U3003 (N_3003,N_2397,N_1358);
and U3004 (N_3004,N_1858,N_1779);
nand U3005 (N_3005,N_531,N_632);
nor U3006 (N_3006,N_1592,N_1510);
and U3007 (N_3007,N_602,N_2466);
and U3008 (N_3008,N_483,N_600);
or U3009 (N_3009,N_1412,N_1968);
and U3010 (N_3010,N_524,N_1350);
nor U3011 (N_3011,N_2249,N_1466);
xor U3012 (N_3012,N_900,N_1072);
or U3013 (N_3013,N_99,N_1470);
and U3014 (N_3014,N_67,N_557);
and U3015 (N_3015,N_1859,N_2488);
nor U3016 (N_3016,N_1297,N_779);
or U3017 (N_3017,N_1774,N_1031);
nor U3018 (N_3018,N_1959,N_1637);
or U3019 (N_3019,N_1908,N_1916);
nand U3020 (N_3020,N_396,N_1438);
xor U3021 (N_3021,N_1928,N_552);
nor U3022 (N_3022,N_1789,N_1003);
nand U3023 (N_3023,N_1368,N_418);
or U3024 (N_3024,N_499,N_1339);
nor U3025 (N_3025,N_1131,N_776);
nand U3026 (N_3026,N_2423,N_296);
nor U3027 (N_3027,N_1812,N_476);
nand U3028 (N_3028,N_2054,N_912);
or U3029 (N_3029,N_1991,N_1691);
or U3030 (N_3030,N_1206,N_1103);
nor U3031 (N_3031,N_2014,N_1983);
and U3032 (N_3032,N_1065,N_646);
nor U3033 (N_3033,N_699,N_2474);
and U3034 (N_3034,N_1695,N_613);
nor U3035 (N_3035,N_1792,N_1419);
nor U3036 (N_3036,N_440,N_97);
or U3037 (N_3037,N_1449,N_2483);
or U3038 (N_3038,N_172,N_280);
nand U3039 (N_3039,N_795,N_2479);
nand U3040 (N_3040,N_135,N_1243);
xor U3041 (N_3041,N_1506,N_393);
nand U3042 (N_3042,N_2294,N_147);
nand U3043 (N_3043,N_286,N_863);
nand U3044 (N_3044,N_1627,N_968);
nand U3045 (N_3045,N_960,N_353);
nor U3046 (N_3046,N_1736,N_1556);
or U3047 (N_3047,N_1495,N_1142);
and U3048 (N_3048,N_1594,N_932);
or U3049 (N_3049,N_1326,N_1931);
and U3050 (N_3050,N_378,N_331);
nand U3051 (N_3051,N_290,N_1937);
and U3052 (N_3052,N_44,N_1219);
or U3053 (N_3053,N_758,N_2257);
or U3054 (N_3054,N_534,N_2254);
or U3055 (N_3055,N_2380,N_955);
nor U3056 (N_3056,N_1212,N_1626);
nand U3057 (N_3057,N_1050,N_1250);
xnor U3058 (N_3058,N_107,N_796);
and U3059 (N_3059,N_1384,N_1804);
xor U3060 (N_3060,N_1992,N_2374);
nand U3061 (N_3061,N_2103,N_1503);
nor U3062 (N_3062,N_1254,N_1253);
nor U3063 (N_3063,N_1516,N_251);
and U3064 (N_3064,N_2298,N_1053);
nand U3065 (N_3065,N_1999,N_794);
or U3066 (N_3066,N_579,N_439);
nand U3067 (N_3067,N_1559,N_278);
or U3068 (N_3068,N_1851,N_2120);
nor U3069 (N_3069,N_168,N_477);
and U3070 (N_3070,N_1247,N_2268);
and U3071 (N_3071,N_1978,N_2347);
nand U3072 (N_3072,N_1883,N_1667);
nand U3073 (N_3073,N_1471,N_303);
and U3074 (N_3074,N_277,N_920);
nor U3075 (N_3075,N_1501,N_1505);
nand U3076 (N_3076,N_751,N_1934);
nor U3077 (N_3077,N_182,N_1207);
or U3078 (N_3078,N_1234,N_1035);
and U3079 (N_3079,N_606,N_508);
and U3080 (N_3080,N_979,N_998);
nand U3081 (N_3081,N_2115,N_1522);
nand U3082 (N_3082,N_433,N_1235);
or U3083 (N_3083,N_1524,N_373);
nand U3084 (N_3084,N_14,N_1376);
nor U3085 (N_3085,N_1708,N_226);
or U3086 (N_3086,N_131,N_2328);
nor U3087 (N_3087,N_1835,N_1969);
or U3088 (N_3088,N_1121,N_764);
or U3089 (N_3089,N_1018,N_2198);
and U3090 (N_3090,N_1722,N_1029);
and U3091 (N_3091,N_1500,N_1294);
or U3092 (N_3092,N_2290,N_1828);
nor U3093 (N_3093,N_142,N_124);
and U3094 (N_3094,N_289,N_2149);
nand U3095 (N_3095,N_638,N_2428);
or U3096 (N_3096,N_556,N_271);
or U3097 (N_3097,N_1083,N_550);
or U3098 (N_3098,N_1998,N_36);
nand U3099 (N_3099,N_184,N_2398);
nor U3100 (N_3100,N_957,N_2214);
xnor U3101 (N_3101,N_2074,N_1699);
and U3102 (N_3102,N_210,N_1425);
nand U3103 (N_3103,N_2272,N_1263);
and U3104 (N_3104,N_1609,N_1051);
nand U3105 (N_3105,N_2480,N_1096);
or U3106 (N_3106,N_82,N_2431);
and U3107 (N_3107,N_1167,N_1238);
or U3108 (N_3108,N_1644,N_1034);
nor U3109 (N_3109,N_103,N_568);
nand U3110 (N_3110,N_332,N_983);
nand U3111 (N_3111,N_1860,N_249);
and U3112 (N_3112,N_1675,N_1417);
nand U3113 (N_3113,N_1066,N_1150);
and U3114 (N_3114,N_2187,N_186);
nor U3115 (N_3115,N_2481,N_330);
nand U3116 (N_3116,N_2259,N_781);
nor U3117 (N_3117,N_745,N_741);
nor U3118 (N_3118,N_201,N_257);
or U3119 (N_3119,N_987,N_1120);
nor U3120 (N_3120,N_1668,N_2102);
and U3121 (N_3121,N_937,N_1293);
or U3122 (N_3122,N_2316,N_281);
and U3123 (N_3123,N_1125,N_598);
nand U3124 (N_3124,N_259,N_221);
nand U3125 (N_3125,N_163,N_1474);
or U3126 (N_3126,N_1560,N_148);
nand U3127 (N_3127,N_1265,N_171);
nand U3128 (N_3128,N_2170,N_1997);
xor U3129 (N_3129,N_1693,N_47);
and U3130 (N_3130,N_1177,N_2002);
nand U3131 (N_3131,N_1342,N_887);
nor U3132 (N_3132,N_1509,N_1650);
or U3133 (N_3133,N_956,N_315);
nand U3134 (N_3134,N_904,N_1676);
nand U3135 (N_3135,N_40,N_448);
nor U3136 (N_3136,N_77,N_622);
nand U3137 (N_3137,N_573,N_1815);
nor U3138 (N_3138,N_179,N_1671);
or U3139 (N_3139,N_792,N_1098);
and U3140 (N_3140,N_1378,N_2177);
and U3141 (N_3141,N_1210,N_733);
nand U3142 (N_3142,N_1363,N_1225);
and U3143 (N_3143,N_2306,N_1086);
or U3144 (N_3144,N_1731,N_1429);
xnor U3145 (N_3145,N_1848,N_687);
and U3146 (N_3146,N_1327,N_798);
or U3147 (N_3147,N_256,N_1657);
nor U3148 (N_3148,N_2233,N_2277);
and U3149 (N_3149,N_430,N_695);
nand U3150 (N_3150,N_1909,N_2383);
and U3151 (N_3151,N_583,N_1233);
or U3152 (N_3152,N_1377,N_908);
nand U3153 (N_3153,N_627,N_59);
and U3154 (N_3154,N_2100,N_601);
and U3155 (N_3155,N_1201,N_329);
or U3156 (N_3156,N_617,N_519);
nor U3157 (N_3157,N_729,N_2022);
nand U3158 (N_3158,N_258,N_856);
nand U3159 (N_3159,N_1528,N_716);
or U3160 (N_3160,N_962,N_1427);
and U3161 (N_3161,N_291,N_1107);
and U3162 (N_3162,N_218,N_1088);
nor U3163 (N_3163,N_1822,N_2325);
and U3164 (N_3164,N_964,N_1040);
and U3165 (N_3165,N_1906,N_862);
xnor U3166 (N_3166,N_1434,N_1469);
and U3167 (N_3167,N_1045,N_1067);
nand U3168 (N_3168,N_1737,N_2039);
and U3169 (N_3169,N_1846,N_1957);
and U3170 (N_3170,N_118,N_416);
nand U3171 (N_3171,N_2263,N_309);
and U3172 (N_3172,N_2420,N_507);
or U3173 (N_3173,N_680,N_2215);
or U3174 (N_3174,N_1123,N_1980);
and U3175 (N_3175,N_510,N_1778);
nand U3176 (N_3176,N_1359,N_1408);
or U3177 (N_3177,N_891,N_269);
and U3178 (N_3178,N_1601,N_1579);
and U3179 (N_3179,N_225,N_1345);
or U3180 (N_3180,N_2189,N_630);
xnor U3181 (N_3181,N_2041,N_2194);
and U3182 (N_3182,N_1919,N_683);
nor U3183 (N_3183,N_1038,N_1205);
or U3184 (N_3184,N_2217,N_2331);
nor U3185 (N_3185,N_1102,N_2471);
or U3186 (N_3186,N_1794,N_713);
or U3187 (N_3187,N_367,N_1493);
and U3188 (N_3188,N_1521,N_543);
nor U3189 (N_3189,N_1285,N_724);
nor U3190 (N_3190,N_1802,N_1960);
nor U3191 (N_3191,N_675,N_2061);
or U3192 (N_3192,N_1490,N_2067);
nand U3193 (N_3193,N_2465,N_2108);
nor U3194 (N_3194,N_2137,N_1392);
or U3195 (N_3195,N_1178,N_804);
nand U3196 (N_3196,N_735,N_2358);
and U3197 (N_3197,N_1832,N_1316);
or U3198 (N_3198,N_37,N_449);
xnor U3199 (N_3199,N_283,N_2057);
nor U3200 (N_3200,N_1507,N_173);
nand U3201 (N_3201,N_1984,N_717);
or U3202 (N_3202,N_2006,N_2323);
or U3203 (N_3203,N_1743,N_548);
nor U3204 (N_3204,N_1042,N_333);
nand U3205 (N_3205,N_2340,N_2104);
nor U3206 (N_3206,N_816,N_1158);
or U3207 (N_3207,N_466,N_335);
nor U3208 (N_3208,N_324,N_474);
or U3209 (N_3209,N_1111,N_341);
nor U3210 (N_3210,N_1312,N_2371);
nand U3211 (N_3211,N_2315,N_438);
and U3212 (N_3212,N_2195,N_397);
nor U3213 (N_3213,N_2034,N_772);
xor U3214 (N_3214,N_926,N_888);
or U3215 (N_3215,N_2437,N_372);
nor U3216 (N_3216,N_1119,N_35);
xnor U3217 (N_3217,N_2346,N_2163);
nand U3218 (N_3218,N_1192,N_24);
or U3219 (N_3219,N_1218,N_2460);
nor U3220 (N_3220,N_2442,N_2455);
nor U3221 (N_3221,N_2072,N_492);
nand U3222 (N_3222,N_1270,N_1639);
and U3223 (N_3223,N_62,N_2211);
nor U3224 (N_3224,N_68,N_2157);
nand U3225 (N_3225,N_61,N_1555);
or U3226 (N_3226,N_671,N_1577);
and U3227 (N_3227,N_1436,N_818);
and U3228 (N_3228,N_265,N_2244);
and U3229 (N_3229,N_57,N_2271);
or U3230 (N_3230,N_1607,N_51);
nand U3231 (N_3231,N_2390,N_1204);
nand U3232 (N_3232,N_1172,N_1582);
or U3233 (N_3233,N_1386,N_279);
nand U3234 (N_3234,N_308,N_1300);
nand U3235 (N_3235,N_1602,N_174);
nand U3236 (N_3236,N_2008,N_1473);
nand U3237 (N_3237,N_1696,N_2490);
nor U3238 (N_3238,N_1328,N_1606);
or U3239 (N_3239,N_897,N_392);
nor U3240 (N_3240,N_354,N_191);
or U3241 (N_3241,N_1823,N_615);
nand U3242 (N_3242,N_1808,N_2369);
nand U3243 (N_3243,N_1391,N_1155);
nor U3244 (N_3244,N_33,N_2333);
nor U3245 (N_3245,N_450,N_2201);
and U3246 (N_3246,N_56,N_1724);
nand U3247 (N_3247,N_2498,N_2430);
or U3248 (N_3248,N_936,N_2188);
or U3249 (N_3249,N_343,N_2273);
nand U3250 (N_3250,N_98,N_1935);
nor U3251 (N_3251,N_2337,N_1773);
xnor U3252 (N_3252,N_882,N_1888);
or U3253 (N_3253,N_651,N_1681);
and U3254 (N_3254,N_2178,N_1889);
and U3255 (N_3255,N_170,N_815);
xor U3256 (N_3256,N_784,N_1482);
nor U3257 (N_3257,N_1877,N_1603);
or U3258 (N_3258,N_374,N_2241);
nor U3259 (N_3259,N_2240,N_696);
or U3260 (N_3260,N_1712,N_1947);
or U3261 (N_3261,N_766,N_2082);
xor U3262 (N_3262,N_1173,N_2281);
or U3263 (N_3263,N_454,N_1786);
nand U3264 (N_3264,N_1421,N_1179);
nor U3265 (N_3265,N_348,N_647);
nor U3266 (N_3266,N_403,N_2045);
nor U3267 (N_3267,N_835,N_2077);
or U3268 (N_3268,N_1442,N_241);
nor U3269 (N_3269,N_92,N_1242);
and U3270 (N_3270,N_2243,N_1783);
and U3271 (N_3271,N_1283,N_151);
nand U3272 (N_3272,N_1302,N_1818);
nand U3273 (N_3273,N_989,N_2295);
nor U3274 (N_3274,N_2499,N_2336);
or U3275 (N_3275,N_60,N_347);
and U3276 (N_3276,N_1752,N_1922);
nor U3277 (N_3277,N_1853,N_1002);
and U3278 (N_3278,N_2329,N_561);
and U3279 (N_3279,N_1864,N_1224);
nand U3280 (N_3280,N_1923,N_1915);
and U3281 (N_3281,N_2270,N_2361);
and U3282 (N_3282,N_825,N_922);
nor U3283 (N_3283,N_559,N_1766);
and U3284 (N_3284,N_295,N_1106);
nor U3285 (N_3285,N_963,N_1287);
and U3286 (N_3286,N_294,N_1813);
nor U3287 (N_3287,N_2292,N_592);
and U3288 (N_3288,N_1134,N_1229);
nand U3289 (N_3289,N_502,N_752);
nand U3290 (N_3290,N_1231,N_1836);
or U3291 (N_3291,N_1631,N_889);
nand U3292 (N_3292,N_1028,N_1016);
xor U3293 (N_3293,N_1298,N_693);
nor U3294 (N_3294,N_2311,N_740);
and U3295 (N_3295,N_2202,N_2090);
and U3296 (N_3296,N_2020,N_1887);
and U3297 (N_3297,N_2058,N_2109);
or U3298 (N_3298,N_253,N_2285);
nand U3299 (N_3299,N_1264,N_652);
nand U3300 (N_3300,N_337,N_162);
and U3301 (N_3301,N_851,N_2307);
and U3302 (N_3302,N_636,N_2151);
nor U3303 (N_3303,N_672,N_847);
and U3304 (N_3304,N_1654,N_2261);
nand U3305 (N_3305,N_958,N_844);
nand U3306 (N_3306,N_2449,N_1479);
nor U3307 (N_3307,N_1249,N_2001);
nand U3308 (N_3308,N_1196,N_328);
and U3309 (N_3309,N_810,N_2168);
or U3310 (N_3310,N_965,N_272);
or U3311 (N_3311,N_1810,N_1129);
and U3312 (N_3312,N_189,N_1273);
and U3313 (N_3313,N_2353,N_1742);
and U3314 (N_3314,N_2421,N_2111);
xnor U3315 (N_3315,N_542,N_317);
and U3316 (N_3316,N_178,N_824);
nor U3317 (N_3317,N_2153,N_1775);
or U3318 (N_3318,N_953,N_88);
nand U3319 (N_3319,N_1465,N_1077);
xor U3320 (N_3320,N_992,N_2464);
and U3321 (N_3321,N_1514,N_1534);
or U3322 (N_3322,N_1246,N_1841);
nand U3323 (N_3323,N_709,N_2429);
and U3324 (N_3324,N_48,N_2171);
nand U3325 (N_3325,N_176,N_197);
and U3326 (N_3326,N_29,N_990);
or U3327 (N_3327,N_406,N_204);
and U3328 (N_3328,N_750,N_1271);
and U3329 (N_3329,N_1176,N_1958);
nand U3330 (N_3330,N_445,N_893);
and U3331 (N_3331,N_2161,N_1807);
and U3332 (N_3332,N_1967,N_2348);
and U3333 (N_3333,N_2446,N_1023);
nor U3334 (N_3334,N_1137,N_1684);
and U3335 (N_3335,N_663,N_899);
nor U3336 (N_3336,N_2283,N_604);
nand U3337 (N_3337,N_867,N_2105);
nand U3338 (N_3338,N_817,N_122);
and U3339 (N_3339,N_1280,N_1820);
nor U3340 (N_3340,N_270,N_1872);
nor U3341 (N_3341,N_603,N_377);
and U3342 (N_3342,N_2173,N_53);
nor U3343 (N_3343,N_2475,N_2050);
and U3344 (N_3344,N_1197,N_419);
nand U3345 (N_3345,N_538,N_1186);
nor U3346 (N_3346,N_150,N_2472);
nor U3347 (N_3347,N_1683,N_2117);
nand U3348 (N_3348,N_539,N_806);
and U3349 (N_3349,N_526,N_157);
and U3350 (N_3350,N_852,N_1215);
nand U3351 (N_3351,N_108,N_1349);
nand U3352 (N_3352,N_2029,N_2234);
nor U3353 (N_3353,N_515,N_2158);
xnor U3354 (N_3354,N_326,N_1208);
or U3355 (N_3355,N_1780,N_2415);
and U3356 (N_3356,N_2070,N_2005);
and U3357 (N_3357,N_2288,N_121);
nor U3358 (N_3358,N_1954,N_1746);
nand U3359 (N_3359,N_754,N_1618);
nor U3360 (N_3360,N_342,N_421);
nand U3361 (N_3361,N_1525,N_919);
nor U3362 (N_3362,N_715,N_2121);
nor U3363 (N_3363,N_1511,N_1761);
and U3364 (N_3364,N_1921,N_1432);
or U3365 (N_3365,N_2489,N_681);
nor U3366 (N_3366,N_86,N_2354);
and U3367 (N_3367,N_1765,N_2260);
nor U3368 (N_3368,N_2417,N_2172);
nor U3369 (N_3369,N_720,N_639);
nand U3370 (N_3370,N_198,N_2049);
nand U3371 (N_3371,N_2196,N_455);
and U3372 (N_3372,N_1027,N_726);
and U3373 (N_3373,N_237,N_10);
and U3374 (N_3374,N_1548,N_1101);
nand U3375 (N_3375,N_874,N_111);
nand U3376 (N_3376,N_1781,N_2027);
and U3377 (N_3377,N_995,N_1171);
nor U3378 (N_3378,N_967,N_2419);
nand U3379 (N_3379,N_1140,N_267);
and U3380 (N_3380,N_540,N_710);
nand U3381 (N_3381,N_1159,N_468);
nor U3382 (N_3382,N_1558,N_13);
and U3383 (N_3383,N_2252,N_2193);
nand U3384 (N_3384,N_1686,N_714);
and U3385 (N_3385,N_931,N_475);
nand U3386 (N_3386,N_1409,N_830);
and U3387 (N_3387,N_1531,N_1025);
nand U3388 (N_3388,N_276,N_1132);
or U3389 (N_3389,N_1117,N_718);
and U3390 (N_3390,N_102,N_2326);
and U3391 (N_3391,N_1616,N_1109);
or U3392 (N_3392,N_200,N_658);
nand U3393 (N_3393,N_947,N_2239);
nor U3394 (N_3394,N_1717,N_64);
or U3395 (N_3395,N_1127,N_914);
and U3396 (N_3396,N_1856,N_649);
nor U3397 (N_3397,N_306,N_415);
or U3398 (N_3398,N_607,N_39);
nor U3399 (N_3399,N_996,N_2180);
nand U3400 (N_3400,N_1136,N_1095);
nand U3401 (N_3401,N_126,N_1407);
nand U3402 (N_3402,N_1652,N_1185);
and U3403 (N_3403,N_582,N_247);
and U3404 (N_3404,N_2207,N_634);
or U3405 (N_3405,N_1487,N_349);
nor U3406 (N_3406,N_760,N_688);
or U3407 (N_3407,N_1891,N_2486);
nand U3408 (N_3408,N_2275,N_81);
nand U3409 (N_3409,N_1330,N_1362);
and U3410 (N_3410,N_1513,N_2052);
or U3411 (N_3411,N_1649,N_1);
and U3412 (N_3412,N_2132,N_494);
nor U3413 (N_3413,N_2032,N_1091);
nand U3414 (N_3414,N_30,N_346);
and U3415 (N_3415,N_388,N_1809);
and U3416 (N_3416,N_2179,N_2140);
nor U3417 (N_3417,N_429,N_1611);
xnor U3418 (N_3418,N_1304,N_1942);
or U3419 (N_3419,N_1647,N_1195);
nor U3420 (N_3420,N_78,N_2385);
or U3421 (N_3421,N_2175,N_2112);
nor U3422 (N_3422,N_129,N_284);
nor U3423 (N_3423,N_2223,N_586);
nand U3424 (N_3424,N_2363,N_2386);
nor U3425 (N_3425,N_1019,N_1484);
or U3426 (N_3426,N_2356,N_2286);
and U3427 (N_3427,N_593,N_190);
nand U3428 (N_3428,N_1767,N_1985);
and U3429 (N_3429,N_712,N_2484);
nand U3430 (N_3430,N_1827,N_1541);
and U3431 (N_3431,N_637,N_2118);
nor U3432 (N_3432,N_1062,N_1056);
nand U3433 (N_3433,N_301,N_642);
and U3434 (N_3434,N_2448,N_1341);
and U3435 (N_3435,N_1564,N_1405);
nor U3436 (N_3436,N_1356,N_1857);
and U3437 (N_3437,N_112,N_2078);
or U3438 (N_3438,N_2087,N_1147);
nand U3439 (N_3439,N_605,N_669);
or U3440 (N_3440,N_881,N_1912);
and U3441 (N_3441,N_1588,N_2422);
and U3442 (N_3442,N_2395,N_1288);
nand U3443 (N_3443,N_1068,N_516);
and U3444 (N_3444,N_1580,N_621);
and U3445 (N_3445,N_2131,N_4);
and U3446 (N_3446,N_2124,N_1461);
nor U3447 (N_3447,N_452,N_1448);
and U3448 (N_3448,N_2255,N_214);
and U3449 (N_3449,N_1612,N_1963);
nor U3450 (N_3450,N_1785,N_2341);
or U3451 (N_3451,N_589,N_2081);
nor U3452 (N_3452,N_2183,N_2136);
nand U3453 (N_3453,N_2287,N_1444);
nor U3454 (N_3454,N_1478,N_668);
or U3455 (N_3455,N_1552,N_2375);
and U3456 (N_3456,N_587,N_2250);
and U3457 (N_3457,N_115,N_518);
nor U3458 (N_3458,N_1973,N_993);
or U3459 (N_3459,N_1402,N_1022);
nor U3460 (N_3460,N_314,N_2301);
nor U3461 (N_3461,N_832,N_1337);
nand U3462 (N_3462,N_2425,N_854);
nor U3463 (N_3463,N_1424,N_793);
nor U3464 (N_3464,N_2467,N_883);
or U3465 (N_3465,N_813,N_467);
nor U3466 (N_3466,N_164,N_1114);
nand U3467 (N_3467,N_572,N_1428);
xnor U3468 (N_3468,N_2229,N_2059);
nor U3469 (N_3469,N_434,N_1464);
and U3470 (N_3470,N_385,N_599);
and U3471 (N_3471,N_409,N_1943);
or U3472 (N_3472,N_1643,N_2267);
nor U3473 (N_3473,N_43,N_2376);
or U3474 (N_3474,N_1373,N_1122);
and U3475 (N_3475,N_2319,N_2258);
and U3476 (N_3476,N_17,N_193);
and U3477 (N_3477,N_2269,N_1008);
or U3478 (N_3478,N_2216,N_802);
nor U3479 (N_3479,N_616,N_1756);
nor U3480 (N_3480,N_1728,N_402);
or U3481 (N_3481,N_901,N_2246);
nor U3482 (N_3482,N_1486,N_242);
nand U3483 (N_3483,N_1567,N_845);
nor U3484 (N_3484,N_1321,N_1085);
and U3485 (N_3485,N_1734,N_1591);
and U3486 (N_3486,N_1310,N_2076);
nand U3487 (N_3487,N_1945,N_2414);
nand U3488 (N_3488,N_1987,N_1536);
and U3489 (N_3489,N_1795,N_394);
and U3490 (N_3490,N_2492,N_451);
nand U3491 (N_3491,N_161,N_2003);
or U3492 (N_3492,N_156,N_978);
nor U3493 (N_3493,N_840,N_2114);
or U3494 (N_3494,N_1284,N_2037);
and U3495 (N_3495,N_1870,N_562);
nor U3496 (N_3496,N_63,N_1714);
or U3497 (N_3497,N_585,N_1193);
or U3498 (N_3498,N_1169,N_1623);
nor U3499 (N_3499,N_228,N_1269);
nand U3500 (N_3500,N_1183,N_902);
nor U3501 (N_3501,N_2225,N_869);
nand U3502 (N_3502,N_1331,N_1274);
or U3503 (N_3503,N_759,N_1477);
nor U3504 (N_3504,N_1678,N_1075);
nor U3505 (N_3505,N_2487,N_128);
and U3506 (N_3506,N_1572,N_1380);
or U3507 (N_3507,N_1939,N_1620);
nand U3508 (N_3508,N_1641,N_697);
or U3509 (N_3509,N_1961,N_1971);
nor U3510 (N_3510,N_575,N_239);
or U3511 (N_3511,N_2338,N_1549);
or U3512 (N_3512,N_1723,N_1182);
nor U3513 (N_3513,N_1060,N_488);
nor U3514 (N_3514,N_106,N_1543);
and U3515 (N_3515,N_358,N_1143);
and U3516 (N_3516,N_1307,N_263);
xor U3517 (N_3517,N_2238,N_1662);
and U3518 (N_3518,N_1164,N_1375);
or U3519 (N_3519,N_2382,N_2167);
nor U3520 (N_3520,N_432,N_1875);
xor U3521 (N_3521,N_1757,N_805);
and U3522 (N_3522,N_2083,N_763);
nand U3523 (N_3523,N_1547,N_1944);
nand U3524 (N_3524,N_1646,N_1893);
and U3525 (N_3525,N_1211,N_890);
nand U3526 (N_3526,N_339,N_2342);
nand U3527 (N_3527,N_498,N_2099);
and U3528 (N_3528,N_1979,N_1079);
and U3529 (N_3529,N_753,N_660);
nor U3530 (N_3530,N_2405,N_1112);
or U3531 (N_3531,N_1387,N_1533);
or U3532 (N_3532,N_1076,N_684);
xnor U3533 (N_3533,N_1426,N_2445);
and U3534 (N_3534,N_351,N_152);
or U3535 (N_3535,N_1952,N_297);
or U3536 (N_3536,N_1082,N_365);
nor U3537 (N_3537,N_702,N_2182);
or U3538 (N_3538,N_682,N_1277);
and U3539 (N_3539,N_1244,N_1682);
nand U3540 (N_3540,N_725,N_196);
nor U3541 (N_3541,N_1791,N_1936);
nor U3542 (N_3542,N_1092,N_1268);
or U3543 (N_3543,N_925,N_234);
and U3544 (N_3544,N_428,N_1575);
or U3545 (N_3545,N_686,N_1420);
nand U3546 (N_3546,N_1590,N_1323);
and U3547 (N_3547,N_619,N_410);
nand U3548 (N_3548,N_831,N_273);
nand U3549 (N_3549,N_2447,N_961);
nand U3550 (N_3550,N_1721,N_1485);
and U3551 (N_3551,N_2200,N_1175);
or U3552 (N_3552,N_923,N_1440);
and U3553 (N_3553,N_1139,N_2145);
or U3554 (N_3554,N_401,N_928);
nand U3555 (N_3555,N_2400,N_1613);
and U3556 (N_3556,N_1333,N_1703);
nand U3557 (N_3557,N_34,N_1406);
and U3558 (N_3558,N_1747,N_1842);
and U3559 (N_3559,N_293,N_861);
and U3560 (N_3560,N_2160,N_588);
or U3561 (N_3561,N_770,N_1151);
nor U3562 (N_3562,N_2245,N_2035);
nor U3563 (N_3563,N_721,N_1343);
nor U3564 (N_3564,N_1245,N_1624);
and U3565 (N_3565,N_1472,N_1740);
and U3566 (N_3566,N_727,N_1993);
nor U3567 (N_3567,N_2462,N_2274);
and U3568 (N_3568,N_233,N_1729);
nand U3569 (N_3569,N_778,N_180);
nand U3570 (N_3570,N_2144,N_1551);
and U3571 (N_3571,N_1168,N_1895);
and U3572 (N_3572,N_1584,N_1956);
or U3573 (N_3573,N_1152,N_340);
and U3574 (N_3574,N_1061,N_553);
and U3575 (N_3575,N_1366,N_1617);
nor U3576 (N_3576,N_2384,N_2368);
nand U3577 (N_3577,N_2128,N_1184);
nand U3578 (N_3578,N_1578,N_898);
and U3579 (N_3579,N_2364,N_1965);
and U3580 (N_3580,N_2185,N_1735);
or U3581 (N_3581,N_1659,N_2438);
and U3582 (N_3582,N_2135,N_783);
or U3583 (N_3583,N_391,N_299);
nand U3584 (N_3584,N_2458,N_320);
or U3585 (N_3585,N_2011,N_2025);
or U3586 (N_3586,N_285,N_2166);
nor U3587 (N_3587,N_970,N_1194);
or U3588 (N_3588,N_386,N_1950);
nand U3589 (N_3589,N_2367,N_858);
or U3590 (N_3590,N_361,N_1855);
or U3591 (N_3591,N_1914,N_1052);
or U3592 (N_3592,N_248,N_628);
nor U3593 (N_3593,N_1314,N_2396);
nor U3594 (N_3594,N_1651,N_1745);
and U3595 (N_3595,N_2327,N_1566);
nand U3596 (N_3596,N_1365,N_380);
xnor U3597 (N_3597,N_1457,N_1636);
and U3598 (N_3598,N_773,N_2236);
and U3599 (N_3599,N_264,N_2330);
nor U3600 (N_3600,N_692,N_1938);
xnor U3601 (N_3601,N_1840,N_229);
nand U3602 (N_3602,N_626,N_384);
or U3603 (N_3603,N_945,N_1198);
nand U3604 (N_3604,N_473,N_1527);
nor U3605 (N_3605,N_2248,N_444);
nand U3606 (N_3606,N_1805,N_2280);
or U3607 (N_3607,N_2154,N_608);
and U3608 (N_3608,N_1322,N_1422);
nor U3609 (N_3609,N_1223,N_1351);
or U3610 (N_3610,N_1353,N_2147);
or U3611 (N_3611,N_985,N_2069);
and U3612 (N_3612,N_571,N_1237);
or U3613 (N_3613,N_1702,N_1520);
or U3614 (N_3614,N_368,N_123);
or U3615 (N_3615,N_609,N_1762);
and U3616 (N_3616,N_1257,N_1788);
nand U3617 (N_3617,N_942,N_2139);
or U3618 (N_3618,N_1670,N_555);
nor U3619 (N_3619,N_1203,N_1430);
nor U3620 (N_3620,N_54,N_2404);
nand U3621 (N_3621,N_1929,N_1784);
and U3622 (N_3622,N_1166,N_240);
nand U3623 (N_3623,N_2046,N_1475);
or U3624 (N_3624,N_1876,N_1202);
nor U3625 (N_3625,N_1861,N_907);
nand U3626 (N_3626,N_1904,N_2335);
xor U3627 (N_3627,N_382,N_1595);
nand U3628 (N_3628,N_789,N_137);
and U3629 (N_3629,N_183,N_948);
nand U3630 (N_3630,N_1796,N_738);
or U3631 (N_3631,N_1332,N_1209);
nand U3632 (N_3632,N_1553,N_85);
nor U3633 (N_3633,N_836,N_517);
nor U3634 (N_3634,N_732,N_2030);
or U3635 (N_3635,N_1898,N_165);
nor U3636 (N_3636,N_2169,N_1074);
and U3637 (N_3637,N_1227,N_1318);
nand U3638 (N_3638,N_130,N_1880);
nand U3639 (N_3639,N_1191,N_2101);
nor U3640 (N_3640,N_596,N_566);
nand U3641 (N_3641,N_1874,N_2350);
nor U3642 (N_3642,N_2496,N_1849);
nor U3643 (N_3643,N_2451,N_1305);
nor U3644 (N_3644,N_667,N_1905);
nor U3645 (N_3645,N_2435,N_2265);
xnor U3646 (N_3646,N_1941,N_1727);
or U3647 (N_3647,N_786,N_1946);
and U3648 (N_3648,N_977,N_1782);
nand U3649 (N_3649,N_855,N_1296);
nand U3650 (N_3650,N_1630,N_89);
nor U3651 (N_3651,N_453,N_1295);
and U3652 (N_3652,N_1517,N_2023);
and U3653 (N_3653,N_261,N_1669);
and U3654 (N_3654,N_181,N_569);
and U3655 (N_3655,N_345,N_633);
or U3656 (N_3656,N_2043,N_704);
nor U3657 (N_3657,N_744,N_304);
nor U3658 (N_3658,N_2096,N_2370);
or U3659 (N_3659,N_74,N_2141);
nor U3660 (N_3660,N_1634,N_458);
and U3661 (N_3661,N_997,N_2343);
nor U3662 (N_3662,N_1290,N_959);
or U3663 (N_3663,N_1754,N_275);
nand U3664 (N_3664,N_2345,N_2393);
nor U3665 (N_3665,N_2004,N_95);
nand U3666 (N_3666,N_859,N_1816);
nor U3667 (N_3667,N_1711,N_1903);
and U3668 (N_3668,N_2291,N_2296);
or U3669 (N_3669,N_746,N_496);
and U3670 (N_3670,N_383,N_2344);
nor U3671 (N_3671,N_423,N_231);
and U3672 (N_3672,N_2304,N_489);
nand U3673 (N_3673,N_250,N_788);
nor U3674 (N_3674,N_879,N_334);
nand U3675 (N_3675,N_991,N_2394);
nand U3676 (N_3676,N_1162,N_822);
or U3677 (N_3677,N_307,N_973);
or U3678 (N_3678,N_872,N_731);
or U3679 (N_3679,N_472,N_1748);
or U3680 (N_3680,N_2044,N_2093);
nand U3681 (N_3681,N_541,N_1565);
nand U3682 (N_3682,N_791,N_2119);
or U3683 (N_3683,N_1787,N_405);
or U3684 (N_3684,N_15,N_2010);
nand U3685 (N_3685,N_950,N_504);
nand U3686 (N_3686,N_20,N_2293);
nand U3687 (N_3687,N_939,N_944);
or U3688 (N_3688,N_659,N_1258);
and U3689 (N_3689,N_2156,N_820);
or U3690 (N_3690,N_2184,N_576);
or U3691 (N_3691,N_2205,N_565);
and U3692 (N_3692,N_1884,N_656);
xnor U3693 (N_3693,N_1837,N_1868);
nor U3694 (N_3694,N_12,N_665);
or U3695 (N_3695,N_905,N_503);
nand U3696 (N_3696,N_916,N_138);
and U3697 (N_3697,N_209,N_127);
nand U3698 (N_3698,N_580,N_826);
nor U3699 (N_3699,N_145,N_1317);
nand U3700 (N_3700,N_1338,N_318);
nor U3701 (N_3701,N_2436,N_698);
or U3702 (N_3702,N_8,N_2024);
nor U3703 (N_3703,N_26,N_1504);
nand U3704 (N_3704,N_2125,N_407);
nor U3705 (N_3705,N_2473,N_120);
nor U3706 (N_3706,N_838,N_1232);
nand U3707 (N_3707,N_1672,N_2227);
nor U3708 (N_3708,N_875,N_1459);
and U3709 (N_3709,N_436,N_212);
or U3710 (N_3710,N_177,N_981);
xnor U3711 (N_3711,N_871,N_1769);
nor U3712 (N_3712,N_1924,N_404);
or U3713 (N_3713,N_2164,N_943);
and U3714 (N_3714,N_1550,N_876);
and U3715 (N_3715,N_1364,N_1299);
and U3716 (N_3716,N_2284,N_1663);
and U3717 (N_3717,N_969,N_719);
nand U3718 (N_3718,N_775,N_676);
nor U3719 (N_3719,N_459,N_1982);
nor U3720 (N_3720,N_2218,N_2060);
xor U3721 (N_3721,N_2413,N_1394);
nor U3722 (N_3722,N_255,N_1251);
nor U3723 (N_3723,N_2308,N_1741);
and U3724 (N_3724,N_1704,N_1041);
nor U3725 (N_3725,N_2186,N_1228);
nand U3726 (N_3726,N_581,N_2146);
and U3727 (N_3727,N_528,N_1346);
nand U3728 (N_3728,N_570,N_935);
and U3729 (N_3729,N_1925,N_425);
nand U3730 (N_3730,N_1568,N_2228);
and U3731 (N_3731,N_479,N_2162);
nor U3732 (N_3732,N_2432,N_2403);
nor U3733 (N_3733,N_1576,N_260);
and U3734 (N_3734,N_1790,N_1348);
nand U3735 (N_3735,N_972,N_708);
nor U3736 (N_3736,N_1881,N_1571);
or U3737 (N_3737,N_1920,N_1498);
nor U3738 (N_3738,N_827,N_325);
and U3739 (N_3739,N_780,N_1640);
or U3740 (N_3740,N_761,N_866);
or U3741 (N_3741,N_2289,N_1596);
and U3742 (N_3742,N_1395,N_356);
and U3743 (N_3743,N_2247,N_1154);
nand U3744 (N_3744,N_2476,N_1070);
and U3745 (N_3745,N_1758,N_2450);
or U3746 (N_3746,N_1374,N_2065);
or U3747 (N_3747,N_536,N_1451);
nand U3748 (N_3748,N_2084,N_1976);
nor U3749 (N_3749,N_1047,N_1706);
nor U3750 (N_3750,N_1392,N_2310);
nor U3751 (N_3751,N_1736,N_2272);
and U3752 (N_3752,N_2305,N_2181);
or U3753 (N_3753,N_69,N_2457);
or U3754 (N_3754,N_918,N_1118);
and U3755 (N_3755,N_2128,N_2103);
nand U3756 (N_3756,N_1649,N_519);
or U3757 (N_3757,N_1755,N_887);
nand U3758 (N_3758,N_538,N_1308);
nand U3759 (N_3759,N_1602,N_2165);
and U3760 (N_3760,N_90,N_1191);
nor U3761 (N_3761,N_364,N_1624);
nand U3762 (N_3762,N_130,N_1776);
nand U3763 (N_3763,N_2372,N_1700);
or U3764 (N_3764,N_835,N_774);
nor U3765 (N_3765,N_606,N_1380);
or U3766 (N_3766,N_2489,N_116);
nand U3767 (N_3767,N_669,N_729);
or U3768 (N_3768,N_1873,N_804);
and U3769 (N_3769,N_1623,N_919);
nand U3770 (N_3770,N_409,N_2496);
nand U3771 (N_3771,N_1062,N_950);
or U3772 (N_3772,N_1681,N_1641);
nand U3773 (N_3773,N_1381,N_843);
nand U3774 (N_3774,N_2103,N_535);
xnor U3775 (N_3775,N_440,N_1916);
and U3776 (N_3776,N_1643,N_1574);
nand U3777 (N_3777,N_1398,N_2293);
or U3778 (N_3778,N_2465,N_700);
nand U3779 (N_3779,N_1078,N_593);
nand U3780 (N_3780,N_2215,N_1382);
nor U3781 (N_3781,N_1040,N_1706);
and U3782 (N_3782,N_110,N_536);
or U3783 (N_3783,N_1390,N_1438);
nand U3784 (N_3784,N_876,N_917);
nor U3785 (N_3785,N_69,N_2408);
and U3786 (N_3786,N_2286,N_929);
nand U3787 (N_3787,N_1084,N_1701);
and U3788 (N_3788,N_2362,N_708);
or U3789 (N_3789,N_244,N_1995);
nand U3790 (N_3790,N_538,N_1837);
nand U3791 (N_3791,N_2425,N_443);
or U3792 (N_3792,N_1678,N_492);
and U3793 (N_3793,N_418,N_1807);
nand U3794 (N_3794,N_529,N_115);
and U3795 (N_3795,N_1243,N_1178);
or U3796 (N_3796,N_276,N_705);
and U3797 (N_3797,N_1801,N_2247);
or U3798 (N_3798,N_1149,N_141);
or U3799 (N_3799,N_1017,N_714);
nand U3800 (N_3800,N_2045,N_1348);
and U3801 (N_3801,N_1155,N_902);
nand U3802 (N_3802,N_2296,N_2380);
nor U3803 (N_3803,N_1612,N_1031);
nand U3804 (N_3804,N_216,N_1908);
or U3805 (N_3805,N_618,N_424);
or U3806 (N_3806,N_1931,N_807);
nand U3807 (N_3807,N_2231,N_48);
nand U3808 (N_3808,N_1234,N_11);
and U3809 (N_3809,N_122,N_1089);
and U3810 (N_3810,N_2160,N_982);
nor U3811 (N_3811,N_1587,N_2256);
nor U3812 (N_3812,N_2243,N_2344);
and U3813 (N_3813,N_257,N_146);
nor U3814 (N_3814,N_1371,N_346);
nor U3815 (N_3815,N_1582,N_970);
or U3816 (N_3816,N_1191,N_2342);
or U3817 (N_3817,N_68,N_1904);
nor U3818 (N_3818,N_514,N_2336);
and U3819 (N_3819,N_2406,N_1143);
or U3820 (N_3820,N_1112,N_602);
nor U3821 (N_3821,N_288,N_318);
nor U3822 (N_3822,N_846,N_1090);
nand U3823 (N_3823,N_2338,N_1143);
nor U3824 (N_3824,N_1672,N_2287);
or U3825 (N_3825,N_1978,N_1868);
and U3826 (N_3826,N_1432,N_241);
and U3827 (N_3827,N_799,N_1347);
nand U3828 (N_3828,N_1504,N_1603);
nand U3829 (N_3829,N_420,N_647);
and U3830 (N_3830,N_271,N_60);
and U3831 (N_3831,N_516,N_421);
or U3832 (N_3832,N_1830,N_43);
nor U3833 (N_3833,N_1405,N_1199);
and U3834 (N_3834,N_612,N_1753);
nand U3835 (N_3835,N_719,N_980);
xor U3836 (N_3836,N_1773,N_1853);
nor U3837 (N_3837,N_1115,N_1455);
or U3838 (N_3838,N_2483,N_1112);
xnor U3839 (N_3839,N_1067,N_739);
or U3840 (N_3840,N_741,N_434);
nor U3841 (N_3841,N_903,N_987);
nand U3842 (N_3842,N_2328,N_2146);
or U3843 (N_3843,N_339,N_773);
nor U3844 (N_3844,N_1830,N_915);
nand U3845 (N_3845,N_1012,N_721);
nor U3846 (N_3846,N_853,N_2353);
nand U3847 (N_3847,N_1803,N_1626);
nor U3848 (N_3848,N_618,N_1268);
nand U3849 (N_3849,N_264,N_1834);
nor U3850 (N_3850,N_299,N_1312);
or U3851 (N_3851,N_2291,N_155);
nand U3852 (N_3852,N_4,N_1839);
nor U3853 (N_3853,N_2458,N_1936);
and U3854 (N_3854,N_1979,N_692);
nand U3855 (N_3855,N_856,N_1251);
nor U3856 (N_3856,N_1650,N_2239);
nand U3857 (N_3857,N_748,N_2460);
nand U3858 (N_3858,N_115,N_905);
and U3859 (N_3859,N_383,N_362);
or U3860 (N_3860,N_395,N_2359);
or U3861 (N_3861,N_2475,N_1292);
nor U3862 (N_3862,N_1496,N_411);
or U3863 (N_3863,N_847,N_1824);
or U3864 (N_3864,N_262,N_2496);
nand U3865 (N_3865,N_1398,N_1083);
nor U3866 (N_3866,N_1436,N_2465);
or U3867 (N_3867,N_1,N_994);
nor U3868 (N_3868,N_95,N_2449);
nand U3869 (N_3869,N_1843,N_1579);
or U3870 (N_3870,N_2183,N_799);
nand U3871 (N_3871,N_147,N_824);
nor U3872 (N_3872,N_247,N_936);
nor U3873 (N_3873,N_1831,N_1676);
and U3874 (N_3874,N_1670,N_916);
and U3875 (N_3875,N_1056,N_1799);
and U3876 (N_3876,N_2106,N_755);
nand U3877 (N_3877,N_787,N_527);
or U3878 (N_3878,N_2093,N_2417);
nand U3879 (N_3879,N_1264,N_1471);
nand U3880 (N_3880,N_881,N_1714);
nand U3881 (N_3881,N_1207,N_584);
xnor U3882 (N_3882,N_1844,N_1115);
or U3883 (N_3883,N_359,N_2178);
or U3884 (N_3884,N_608,N_936);
nand U3885 (N_3885,N_236,N_882);
and U3886 (N_3886,N_1993,N_149);
or U3887 (N_3887,N_2073,N_1499);
and U3888 (N_3888,N_1961,N_322);
nor U3889 (N_3889,N_1836,N_877);
and U3890 (N_3890,N_1575,N_424);
nor U3891 (N_3891,N_931,N_2226);
nand U3892 (N_3892,N_1050,N_714);
nor U3893 (N_3893,N_806,N_260);
nand U3894 (N_3894,N_611,N_1839);
nor U3895 (N_3895,N_1352,N_1290);
nor U3896 (N_3896,N_1952,N_1107);
or U3897 (N_3897,N_1925,N_851);
nand U3898 (N_3898,N_1193,N_707);
or U3899 (N_3899,N_1277,N_2026);
and U3900 (N_3900,N_1400,N_2132);
and U3901 (N_3901,N_2112,N_1976);
or U3902 (N_3902,N_370,N_896);
and U3903 (N_3903,N_430,N_1253);
nor U3904 (N_3904,N_2017,N_1620);
nand U3905 (N_3905,N_877,N_837);
nor U3906 (N_3906,N_2385,N_1500);
nand U3907 (N_3907,N_2200,N_258);
nor U3908 (N_3908,N_911,N_335);
nand U3909 (N_3909,N_870,N_2296);
xor U3910 (N_3910,N_1241,N_1630);
nor U3911 (N_3911,N_2053,N_1241);
xor U3912 (N_3912,N_444,N_1880);
or U3913 (N_3913,N_2025,N_639);
and U3914 (N_3914,N_1710,N_868);
or U3915 (N_3915,N_1873,N_2205);
and U3916 (N_3916,N_216,N_2120);
xnor U3917 (N_3917,N_1356,N_777);
nor U3918 (N_3918,N_1893,N_135);
and U3919 (N_3919,N_98,N_623);
nor U3920 (N_3920,N_615,N_1959);
and U3921 (N_3921,N_376,N_1567);
nor U3922 (N_3922,N_118,N_956);
nand U3923 (N_3923,N_646,N_1979);
nor U3924 (N_3924,N_1186,N_909);
nand U3925 (N_3925,N_1920,N_1443);
nand U3926 (N_3926,N_873,N_1163);
and U3927 (N_3927,N_973,N_1185);
or U3928 (N_3928,N_754,N_418);
nor U3929 (N_3929,N_2028,N_2362);
nand U3930 (N_3930,N_2257,N_192);
and U3931 (N_3931,N_2273,N_975);
or U3932 (N_3932,N_728,N_522);
nand U3933 (N_3933,N_1974,N_1417);
or U3934 (N_3934,N_789,N_874);
nor U3935 (N_3935,N_2336,N_1476);
or U3936 (N_3936,N_1716,N_1400);
nand U3937 (N_3937,N_2041,N_1064);
nand U3938 (N_3938,N_1868,N_990);
xor U3939 (N_3939,N_2121,N_535);
nand U3940 (N_3940,N_1847,N_38);
nor U3941 (N_3941,N_1072,N_1147);
or U3942 (N_3942,N_469,N_1793);
and U3943 (N_3943,N_1099,N_1754);
nand U3944 (N_3944,N_1876,N_1334);
nor U3945 (N_3945,N_1718,N_674);
and U3946 (N_3946,N_1453,N_832);
or U3947 (N_3947,N_1620,N_2131);
and U3948 (N_3948,N_2068,N_1654);
nor U3949 (N_3949,N_587,N_660);
nor U3950 (N_3950,N_2187,N_1520);
or U3951 (N_3951,N_1185,N_370);
nand U3952 (N_3952,N_576,N_2103);
nand U3953 (N_3953,N_2057,N_1052);
nand U3954 (N_3954,N_918,N_1535);
nand U3955 (N_3955,N_1758,N_1854);
nand U3956 (N_3956,N_990,N_527);
nor U3957 (N_3957,N_1092,N_588);
xor U3958 (N_3958,N_992,N_2378);
nand U3959 (N_3959,N_1058,N_772);
and U3960 (N_3960,N_472,N_13);
nand U3961 (N_3961,N_1891,N_363);
and U3962 (N_3962,N_1623,N_33);
nor U3963 (N_3963,N_1722,N_265);
or U3964 (N_3964,N_1436,N_1164);
nand U3965 (N_3965,N_1889,N_2122);
or U3966 (N_3966,N_16,N_1995);
nand U3967 (N_3967,N_2038,N_1483);
nor U3968 (N_3968,N_895,N_86);
or U3969 (N_3969,N_1723,N_234);
and U3970 (N_3970,N_1494,N_96);
nor U3971 (N_3971,N_952,N_137);
nand U3972 (N_3972,N_864,N_2051);
nor U3973 (N_3973,N_878,N_466);
nand U3974 (N_3974,N_1577,N_1061);
and U3975 (N_3975,N_542,N_1168);
nor U3976 (N_3976,N_2192,N_679);
nor U3977 (N_3977,N_13,N_2035);
and U3978 (N_3978,N_2174,N_1800);
nand U3979 (N_3979,N_12,N_198);
nor U3980 (N_3980,N_1474,N_453);
nor U3981 (N_3981,N_1262,N_70);
or U3982 (N_3982,N_938,N_690);
nor U3983 (N_3983,N_962,N_94);
and U3984 (N_3984,N_2181,N_2097);
nand U3985 (N_3985,N_1113,N_2028);
nor U3986 (N_3986,N_1395,N_1100);
and U3987 (N_3987,N_391,N_884);
or U3988 (N_3988,N_646,N_890);
or U3989 (N_3989,N_1144,N_800);
nor U3990 (N_3990,N_2152,N_16);
nor U3991 (N_3991,N_2020,N_2205);
nor U3992 (N_3992,N_1452,N_723);
nand U3993 (N_3993,N_1382,N_1576);
nor U3994 (N_3994,N_795,N_266);
nand U3995 (N_3995,N_2002,N_1002);
and U3996 (N_3996,N_349,N_1425);
nand U3997 (N_3997,N_2222,N_479);
and U3998 (N_3998,N_1880,N_1205);
or U3999 (N_3999,N_2126,N_2295);
nand U4000 (N_4000,N_1341,N_2212);
and U4001 (N_4001,N_915,N_1776);
nor U4002 (N_4002,N_916,N_2129);
nor U4003 (N_4003,N_384,N_1321);
nor U4004 (N_4004,N_1022,N_756);
nand U4005 (N_4005,N_297,N_267);
nor U4006 (N_4006,N_619,N_14);
and U4007 (N_4007,N_690,N_45);
or U4008 (N_4008,N_1454,N_627);
nand U4009 (N_4009,N_815,N_150);
nand U4010 (N_4010,N_1207,N_660);
or U4011 (N_4011,N_2099,N_1083);
nor U4012 (N_4012,N_1504,N_1751);
or U4013 (N_4013,N_1586,N_436);
xor U4014 (N_4014,N_1772,N_674);
xnor U4015 (N_4015,N_1386,N_2347);
nand U4016 (N_4016,N_1646,N_1293);
nor U4017 (N_4017,N_819,N_549);
or U4018 (N_4018,N_18,N_413);
nor U4019 (N_4019,N_968,N_2329);
or U4020 (N_4020,N_860,N_1976);
nor U4021 (N_4021,N_2310,N_944);
and U4022 (N_4022,N_1024,N_55);
nand U4023 (N_4023,N_1140,N_47);
or U4024 (N_4024,N_710,N_106);
xor U4025 (N_4025,N_2197,N_1981);
and U4026 (N_4026,N_139,N_1555);
nand U4027 (N_4027,N_213,N_2210);
xor U4028 (N_4028,N_64,N_250);
and U4029 (N_4029,N_481,N_1952);
or U4030 (N_4030,N_501,N_2226);
nor U4031 (N_4031,N_1730,N_997);
and U4032 (N_4032,N_731,N_0);
nand U4033 (N_4033,N_4,N_2465);
or U4034 (N_4034,N_1818,N_998);
or U4035 (N_4035,N_2312,N_1384);
nand U4036 (N_4036,N_594,N_1967);
and U4037 (N_4037,N_2155,N_278);
and U4038 (N_4038,N_1981,N_176);
nor U4039 (N_4039,N_937,N_828);
nand U4040 (N_4040,N_1391,N_2411);
and U4041 (N_4041,N_1300,N_1160);
or U4042 (N_4042,N_356,N_1133);
nand U4043 (N_4043,N_922,N_959);
and U4044 (N_4044,N_1950,N_1746);
nand U4045 (N_4045,N_2487,N_660);
nand U4046 (N_4046,N_1465,N_1638);
and U4047 (N_4047,N_1326,N_2328);
and U4048 (N_4048,N_2013,N_2481);
nor U4049 (N_4049,N_1324,N_878);
and U4050 (N_4050,N_726,N_2446);
or U4051 (N_4051,N_2460,N_1690);
and U4052 (N_4052,N_628,N_782);
and U4053 (N_4053,N_2225,N_377);
nor U4054 (N_4054,N_764,N_1733);
and U4055 (N_4055,N_762,N_103);
nor U4056 (N_4056,N_2272,N_2409);
and U4057 (N_4057,N_690,N_406);
nand U4058 (N_4058,N_2069,N_639);
nand U4059 (N_4059,N_519,N_2257);
nor U4060 (N_4060,N_1449,N_2230);
nor U4061 (N_4061,N_366,N_790);
nor U4062 (N_4062,N_756,N_2425);
or U4063 (N_4063,N_1648,N_772);
nor U4064 (N_4064,N_235,N_2116);
or U4065 (N_4065,N_27,N_559);
nand U4066 (N_4066,N_667,N_1327);
nor U4067 (N_4067,N_1539,N_1279);
nand U4068 (N_4068,N_632,N_270);
and U4069 (N_4069,N_1806,N_1882);
nand U4070 (N_4070,N_1715,N_1392);
and U4071 (N_4071,N_1496,N_90);
nor U4072 (N_4072,N_655,N_16);
or U4073 (N_4073,N_531,N_274);
nand U4074 (N_4074,N_154,N_2485);
nor U4075 (N_4075,N_2184,N_167);
nor U4076 (N_4076,N_2341,N_2074);
or U4077 (N_4077,N_1213,N_1687);
nand U4078 (N_4078,N_1518,N_2283);
nand U4079 (N_4079,N_1054,N_1359);
and U4080 (N_4080,N_1346,N_1423);
and U4081 (N_4081,N_1221,N_215);
and U4082 (N_4082,N_1486,N_2114);
nand U4083 (N_4083,N_2036,N_1394);
nand U4084 (N_4084,N_2158,N_1476);
nor U4085 (N_4085,N_2071,N_547);
or U4086 (N_4086,N_679,N_57);
and U4087 (N_4087,N_1885,N_1611);
nand U4088 (N_4088,N_635,N_32);
and U4089 (N_4089,N_2306,N_245);
or U4090 (N_4090,N_2496,N_1076);
nand U4091 (N_4091,N_2109,N_1172);
and U4092 (N_4092,N_1184,N_1904);
nand U4093 (N_4093,N_1489,N_927);
nand U4094 (N_4094,N_1615,N_1849);
nor U4095 (N_4095,N_1661,N_1827);
and U4096 (N_4096,N_808,N_1125);
nor U4097 (N_4097,N_1355,N_1031);
or U4098 (N_4098,N_990,N_1716);
and U4099 (N_4099,N_1362,N_1651);
and U4100 (N_4100,N_892,N_117);
or U4101 (N_4101,N_1225,N_2405);
or U4102 (N_4102,N_813,N_327);
and U4103 (N_4103,N_1108,N_2479);
xor U4104 (N_4104,N_2165,N_1286);
or U4105 (N_4105,N_2343,N_1970);
and U4106 (N_4106,N_1937,N_2386);
nor U4107 (N_4107,N_2222,N_912);
nor U4108 (N_4108,N_2332,N_1575);
or U4109 (N_4109,N_425,N_1602);
xor U4110 (N_4110,N_1025,N_2380);
xnor U4111 (N_4111,N_824,N_1736);
nor U4112 (N_4112,N_518,N_2406);
or U4113 (N_4113,N_915,N_204);
nand U4114 (N_4114,N_2452,N_927);
nor U4115 (N_4115,N_50,N_2046);
or U4116 (N_4116,N_570,N_82);
or U4117 (N_4117,N_831,N_2409);
and U4118 (N_4118,N_13,N_2216);
or U4119 (N_4119,N_2359,N_657);
and U4120 (N_4120,N_2300,N_2448);
nor U4121 (N_4121,N_1470,N_279);
and U4122 (N_4122,N_172,N_1467);
or U4123 (N_4123,N_229,N_1522);
nand U4124 (N_4124,N_799,N_1584);
nand U4125 (N_4125,N_1677,N_1235);
nand U4126 (N_4126,N_1639,N_1140);
nand U4127 (N_4127,N_1238,N_340);
and U4128 (N_4128,N_83,N_1764);
xnor U4129 (N_4129,N_2176,N_1602);
and U4130 (N_4130,N_775,N_823);
nand U4131 (N_4131,N_2185,N_1955);
or U4132 (N_4132,N_1289,N_697);
and U4133 (N_4133,N_1984,N_966);
nor U4134 (N_4134,N_530,N_568);
or U4135 (N_4135,N_2485,N_1236);
or U4136 (N_4136,N_2079,N_301);
and U4137 (N_4137,N_1522,N_217);
or U4138 (N_4138,N_1017,N_764);
nand U4139 (N_4139,N_2224,N_525);
nor U4140 (N_4140,N_539,N_618);
nor U4141 (N_4141,N_659,N_2343);
and U4142 (N_4142,N_1013,N_66);
nor U4143 (N_4143,N_1593,N_1751);
or U4144 (N_4144,N_2446,N_280);
nor U4145 (N_4145,N_1140,N_533);
or U4146 (N_4146,N_1223,N_999);
or U4147 (N_4147,N_1514,N_1771);
nand U4148 (N_4148,N_247,N_2136);
or U4149 (N_4149,N_63,N_1222);
and U4150 (N_4150,N_817,N_1899);
nand U4151 (N_4151,N_1809,N_907);
and U4152 (N_4152,N_1751,N_1373);
nand U4153 (N_4153,N_1414,N_561);
nand U4154 (N_4154,N_1995,N_2185);
xor U4155 (N_4155,N_1583,N_521);
or U4156 (N_4156,N_2362,N_1966);
nand U4157 (N_4157,N_1262,N_1541);
nand U4158 (N_4158,N_362,N_647);
and U4159 (N_4159,N_2031,N_74);
nor U4160 (N_4160,N_879,N_1152);
nand U4161 (N_4161,N_471,N_2453);
nor U4162 (N_4162,N_1609,N_2121);
nor U4163 (N_4163,N_579,N_1508);
nand U4164 (N_4164,N_1062,N_1643);
nand U4165 (N_4165,N_2267,N_585);
nand U4166 (N_4166,N_897,N_1969);
nor U4167 (N_4167,N_1360,N_873);
nor U4168 (N_4168,N_668,N_2429);
and U4169 (N_4169,N_1858,N_957);
or U4170 (N_4170,N_1302,N_2117);
and U4171 (N_4171,N_2122,N_2204);
nor U4172 (N_4172,N_523,N_725);
and U4173 (N_4173,N_1795,N_1223);
nand U4174 (N_4174,N_1198,N_616);
nand U4175 (N_4175,N_103,N_1232);
nand U4176 (N_4176,N_153,N_1084);
and U4177 (N_4177,N_303,N_1691);
or U4178 (N_4178,N_540,N_1573);
nand U4179 (N_4179,N_2141,N_1828);
nor U4180 (N_4180,N_1990,N_1366);
nor U4181 (N_4181,N_2015,N_2476);
nor U4182 (N_4182,N_2304,N_723);
and U4183 (N_4183,N_1918,N_1158);
and U4184 (N_4184,N_1804,N_2201);
nor U4185 (N_4185,N_136,N_1377);
and U4186 (N_4186,N_722,N_112);
nor U4187 (N_4187,N_2089,N_1118);
nor U4188 (N_4188,N_796,N_255);
or U4189 (N_4189,N_1762,N_1537);
or U4190 (N_4190,N_674,N_2256);
or U4191 (N_4191,N_284,N_346);
nor U4192 (N_4192,N_532,N_639);
and U4193 (N_4193,N_1147,N_827);
xnor U4194 (N_4194,N_2105,N_186);
and U4195 (N_4195,N_1089,N_236);
or U4196 (N_4196,N_1146,N_41);
nand U4197 (N_4197,N_1802,N_853);
and U4198 (N_4198,N_1236,N_1423);
or U4199 (N_4199,N_1054,N_2358);
nand U4200 (N_4200,N_1156,N_112);
nor U4201 (N_4201,N_718,N_1727);
nor U4202 (N_4202,N_2202,N_898);
nand U4203 (N_4203,N_1603,N_1186);
nand U4204 (N_4204,N_478,N_347);
or U4205 (N_4205,N_648,N_1966);
nand U4206 (N_4206,N_2491,N_1311);
nor U4207 (N_4207,N_2010,N_559);
and U4208 (N_4208,N_420,N_851);
or U4209 (N_4209,N_204,N_776);
or U4210 (N_4210,N_1410,N_414);
nor U4211 (N_4211,N_1733,N_335);
nor U4212 (N_4212,N_1071,N_671);
and U4213 (N_4213,N_2459,N_387);
and U4214 (N_4214,N_1873,N_218);
nor U4215 (N_4215,N_1620,N_959);
xnor U4216 (N_4216,N_316,N_1824);
nand U4217 (N_4217,N_1661,N_1793);
nor U4218 (N_4218,N_1392,N_2254);
nand U4219 (N_4219,N_2070,N_1556);
nand U4220 (N_4220,N_1857,N_133);
or U4221 (N_4221,N_1985,N_366);
nor U4222 (N_4222,N_1525,N_695);
and U4223 (N_4223,N_827,N_816);
and U4224 (N_4224,N_737,N_1324);
and U4225 (N_4225,N_2196,N_408);
nor U4226 (N_4226,N_905,N_316);
nand U4227 (N_4227,N_974,N_1393);
or U4228 (N_4228,N_383,N_256);
xor U4229 (N_4229,N_1247,N_888);
nand U4230 (N_4230,N_152,N_58);
nor U4231 (N_4231,N_1754,N_1082);
and U4232 (N_4232,N_1549,N_1254);
nand U4233 (N_4233,N_2235,N_431);
nor U4234 (N_4234,N_2317,N_472);
and U4235 (N_4235,N_119,N_236);
nor U4236 (N_4236,N_1439,N_1342);
or U4237 (N_4237,N_2103,N_2093);
nand U4238 (N_4238,N_1473,N_627);
or U4239 (N_4239,N_1186,N_384);
or U4240 (N_4240,N_1101,N_688);
or U4241 (N_4241,N_860,N_2339);
xor U4242 (N_4242,N_2145,N_2231);
nand U4243 (N_4243,N_1895,N_17);
or U4244 (N_4244,N_224,N_1087);
nand U4245 (N_4245,N_1712,N_1227);
or U4246 (N_4246,N_1607,N_606);
nor U4247 (N_4247,N_1236,N_2162);
or U4248 (N_4248,N_378,N_1181);
nor U4249 (N_4249,N_2450,N_1458);
or U4250 (N_4250,N_1991,N_777);
and U4251 (N_4251,N_864,N_2441);
nor U4252 (N_4252,N_1217,N_1929);
and U4253 (N_4253,N_1878,N_1866);
nand U4254 (N_4254,N_1996,N_1915);
nand U4255 (N_4255,N_1376,N_1572);
nor U4256 (N_4256,N_40,N_1314);
and U4257 (N_4257,N_411,N_47);
or U4258 (N_4258,N_1779,N_1349);
nand U4259 (N_4259,N_254,N_2334);
nand U4260 (N_4260,N_1714,N_2016);
and U4261 (N_4261,N_1315,N_2365);
or U4262 (N_4262,N_2153,N_2485);
nand U4263 (N_4263,N_592,N_1528);
nor U4264 (N_4264,N_1059,N_1986);
and U4265 (N_4265,N_2344,N_985);
nand U4266 (N_4266,N_458,N_432);
and U4267 (N_4267,N_1314,N_12);
xor U4268 (N_4268,N_2417,N_2481);
or U4269 (N_4269,N_1960,N_939);
or U4270 (N_4270,N_1998,N_1184);
nand U4271 (N_4271,N_1872,N_1161);
nand U4272 (N_4272,N_97,N_558);
nand U4273 (N_4273,N_115,N_1434);
nand U4274 (N_4274,N_1542,N_1125);
and U4275 (N_4275,N_2443,N_850);
or U4276 (N_4276,N_308,N_102);
or U4277 (N_4277,N_120,N_907);
or U4278 (N_4278,N_1470,N_2425);
and U4279 (N_4279,N_1486,N_56);
nor U4280 (N_4280,N_530,N_1135);
or U4281 (N_4281,N_863,N_2065);
nor U4282 (N_4282,N_1088,N_1320);
and U4283 (N_4283,N_2423,N_496);
nand U4284 (N_4284,N_323,N_2139);
or U4285 (N_4285,N_1473,N_1288);
and U4286 (N_4286,N_514,N_799);
nor U4287 (N_4287,N_154,N_259);
or U4288 (N_4288,N_1571,N_2334);
or U4289 (N_4289,N_2133,N_1727);
nand U4290 (N_4290,N_507,N_555);
nor U4291 (N_4291,N_1174,N_1300);
nand U4292 (N_4292,N_1031,N_1425);
nand U4293 (N_4293,N_1416,N_1470);
nand U4294 (N_4294,N_2081,N_1962);
and U4295 (N_4295,N_112,N_1142);
nor U4296 (N_4296,N_944,N_161);
and U4297 (N_4297,N_1632,N_1864);
or U4298 (N_4298,N_1197,N_2239);
nand U4299 (N_4299,N_1608,N_608);
and U4300 (N_4300,N_2292,N_1916);
nor U4301 (N_4301,N_2062,N_1897);
or U4302 (N_4302,N_1852,N_979);
nor U4303 (N_4303,N_577,N_1120);
nand U4304 (N_4304,N_864,N_1491);
and U4305 (N_4305,N_195,N_2135);
nand U4306 (N_4306,N_2396,N_564);
nor U4307 (N_4307,N_553,N_358);
and U4308 (N_4308,N_1209,N_1206);
and U4309 (N_4309,N_1777,N_213);
and U4310 (N_4310,N_2498,N_2142);
and U4311 (N_4311,N_1580,N_1725);
or U4312 (N_4312,N_853,N_77);
nor U4313 (N_4313,N_1385,N_871);
nor U4314 (N_4314,N_502,N_2460);
nand U4315 (N_4315,N_2441,N_334);
or U4316 (N_4316,N_225,N_1931);
or U4317 (N_4317,N_2031,N_30);
nand U4318 (N_4318,N_1702,N_1943);
and U4319 (N_4319,N_885,N_53);
nand U4320 (N_4320,N_2137,N_336);
nor U4321 (N_4321,N_1708,N_269);
nand U4322 (N_4322,N_588,N_1694);
or U4323 (N_4323,N_1915,N_1544);
xor U4324 (N_4324,N_2222,N_1540);
and U4325 (N_4325,N_1470,N_1650);
nor U4326 (N_4326,N_2282,N_186);
nor U4327 (N_4327,N_345,N_2484);
xnor U4328 (N_4328,N_1207,N_1101);
nor U4329 (N_4329,N_844,N_2220);
and U4330 (N_4330,N_2077,N_2319);
nor U4331 (N_4331,N_1442,N_130);
nor U4332 (N_4332,N_2401,N_19);
nand U4333 (N_4333,N_1772,N_632);
nand U4334 (N_4334,N_731,N_1254);
nand U4335 (N_4335,N_933,N_2113);
or U4336 (N_4336,N_2392,N_2076);
nand U4337 (N_4337,N_1821,N_2454);
nand U4338 (N_4338,N_29,N_2026);
nand U4339 (N_4339,N_219,N_267);
nor U4340 (N_4340,N_398,N_1606);
nor U4341 (N_4341,N_306,N_418);
and U4342 (N_4342,N_1917,N_64);
xor U4343 (N_4343,N_1026,N_376);
and U4344 (N_4344,N_2163,N_344);
or U4345 (N_4345,N_548,N_204);
nand U4346 (N_4346,N_1193,N_2179);
nor U4347 (N_4347,N_411,N_2260);
nand U4348 (N_4348,N_1586,N_2073);
or U4349 (N_4349,N_1965,N_2097);
nor U4350 (N_4350,N_2362,N_1731);
nor U4351 (N_4351,N_675,N_1177);
nand U4352 (N_4352,N_157,N_1472);
nor U4353 (N_4353,N_1672,N_1932);
nor U4354 (N_4354,N_1193,N_2001);
nor U4355 (N_4355,N_2433,N_2148);
nor U4356 (N_4356,N_828,N_1318);
nor U4357 (N_4357,N_2370,N_2421);
and U4358 (N_4358,N_2009,N_1739);
and U4359 (N_4359,N_87,N_2056);
and U4360 (N_4360,N_1686,N_2153);
xor U4361 (N_4361,N_1821,N_1277);
and U4362 (N_4362,N_1453,N_1227);
xnor U4363 (N_4363,N_983,N_1573);
nor U4364 (N_4364,N_1968,N_1120);
or U4365 (N_4365,N_1619,N_355);
nand U4366 (N_4366,N_1001,N_2395);
nand U4367 (N_4367,N_548,N_1696);
nand U4368 (N_4368,N_922,N_1354);
nand U4369 (N_4369,N_1816,N_10);
nor U4370 (N_4370,N_114,N_372);
or U4371 (N_4371,N_838,N_1407);
or U4372 (N_4372,N_965,N_1935);
nor U4373 (N_4373,N_2335,N_2196);
or U4374 (N_4374,N_1996,N_1655);
or U4375 (N_4375,N_558,N_2365);
nor U4376 (N_4376,N_1613,N_227);
nor U4377 (N_4377,N_1714,N_94);
and U4378 (N_4378,N_268,N_2393);
nand U4379 (N_4379,N_198,N_1246);
nand U4380 (N_4380,N_46,N_1809);
and U4381 (N_4381,N_1117,N_428);
nor U4382 (N_4382,N_238,N_17);
or U4383 (N_4383,N_490,N_1872);
xnor U4384 (N_4384,N_1587,N_431);
nor U4385 (N_4385,N_1190,N_381);
nand U4386 (N_4386,N_2208,N_1307);
or U4387 (N_4387,N_1102,N_2271);
nand U4388 (N_4388,N_2003,N_1205);
and U4389 (N_4389,N_620,N_1663);
and U4390 (N_4390,N_308,N_2216);
nor U4391 (N_4391,N_233,N_1954);
nand U4392 (N_4392,N_320,N_412);
nand U4393 (N_4393,N_2297,N_2196);
nor U4394 (N_4394,N_436,N_1654);
or U4395 (N_4395,N_584,N_976);
and U4396 (N_4396,N_1073,N_815);
or U4397 (N_4397,N_1481,N_363);
or U4398 (N_4398,N_1933,N_1205);
nor U4399 (N_4399,N_1074,N_1289);
nor U4400 (N_4400,N_1124,N_147);
nor U4401 (N_4401,N_817,N_2227);
nand U4402 (N_4402,N_2249,N_79);
and U4403 (N_4403,N_1164,N_1556);
nand U4404 (N_4404,N_1514,N_1726);
nor U4405 (N_4405,N_1795,N_385);
nand U4406 (N_4406,N_984,N_835);
nor U4407 (N_4407,N_828,N_1669);
nand U4408 (N_4408,N_1504,N_2076);
nand U4409 (N_4409,N_1094,N_1879);
nor U4410 (N_4410,N_103,N_413);
and U4411 (N_4411,N_1047,N_1457);
and U4412 (N_4412,N_1452,N_34);
or U4413 (N_4413,N_2356,N_633);
and U4414 (N_4414,N_416,N_1280);
nor U4415 (N_4415,N_1031,N_1341);
nor U4416 (N_4416,N_2317,N_1874);
and U4417 (N_4417,N_1778,N_1476);
nand U4418 (N_4418,N_1470,N_1406);
or U4419 (N_4419,N_718,N_711);
nor U4420 (N_4420,N_2451,N_2366);
nor U4421 (N_4421,N_690,N_1654);
and U4422 (N_4422,N_1504,N_659);
nand U4423 (N_4423,N_293,N_1237);
nand U4424 (N_4424,N_1275,N_1143);
or U4425 (N_4425,N_1193,N_298);
or U4426 (N_4426,N_1248,N_80);
and U4427 (N_4427,N_802,N_68);
and U4428 (N_4428,N_2240,N_1160);
and U4429 (N_4429,N_2016,N_1920);
nand U4430 (N_4430,N_2058,N_1066);
and U4431 (N_4431,N_1250,N_394);
and U4432 (N_4432,N_2236,N_29);
or U4433 (N_4433,N_1301,N_1068);
nor U4434 (N_4434,N_1800,N_1981);
and U4435 (N_4435,N_1563,N_1683);
nand U4436 (N_4436,N_1248,N_781);
nand U4437 (N_4437,N_2006,N_524);
and U4438 (N_4438,N_2397,N_820);
or U4439 (N_4439,N_636,N_2446);
nor U4440 (N_4440,N_2428,N_831);
nand U4441 (N_4441,N_2287,N_1047);
nand U4442 (N_4442,N_660,N_1863);
and U4443 (N_4443,N_1434,N_2155);
nand U4444 (N_4444,N_2446,N_2225);
and U4445 (N_4445,N_2434,N_2476);
nor U4446 (N_4446,N_1161,N_1382);
nor U4447 (N_4447,N_102,N_2448);
nand U4448 (N_4448,N_1905,N_711);
and U4449 (N_4449,N_2085,N_415);
and U4450 (N_4450,N_2314,N_2213);
or U4451 (N_4451,N_493,N_314);
and U4452 (N_4452,N_203,N_1709);
xnor U4453 (N_4453,N_510,N_1274);
xor U4454 (N_4454,N_2353,N_1005);
nand U4455 (N_4455,N_963,N_2221);
and U4456 (N_4456,N_2467,N_2487);
and U4457 (N_4457,N_2302,N_162);
or U4458 (N_4458,N_1425,N_632);
or U4459 (N_4459,N_1180,N_397);
and U4460 (N_4460,N_661,N_74);
xnor U4461 (N_4461,N_1420,N_163);
nor U4462 (N_4462,N_831,N_2189);
nand U4463 (N_4463,N_193,N_2247);
and U4464 (N_4464,N_2207,N_800);
or U4465 (N_4465,N_853,N_890);
and U4466 (N_4466,N_780,N_1680);
nor U4467 (N_4467,N_1735,N_1066);
and U4468 (N_4468,N_1853,N_1560);
nor U4469 (N_4469,N_965,N_2052);
or U4470 (N_4470,N_1375,N_1354);
and U4471 (N_4471,N_2280,N_10);
and U4472 (N_4472,N_1863,N_1918);
nand U4473 (N_4473,N_2481,N_2193);
nand U4474 (N_4474,N_259,N_29);
and U4475 (N_4475,N_1808,N_563);
xnor U4476 (N_4476,N_2123,N_160);
and U4477 (N_4477,N_1972,N_123);
nand U4478 (N_4478,N_2484,N_1772);
xnor U4479 (N_4479,N_974,N_1223);
and U4480 (N_4480,N_791,N_513);
and U4481 (N_4481,N_1155,N_740);
nor U4482 (N_4482,N_890,N_2477);
and U4483 (N_4483,N_1726,N_1521);
and U4484 (N_4484,N_1316,N_1404);
xnor U4485 (N_4485,N_1131,N_1187);
and U4486 (N_4486,N_1615,N_1586);
nor U4487 (N_4487,N_2191,N_119);
or U4488 (N_4488,N_2048,N_512);
nor U4489 (N_4489,N_2092,N_1789);
nand U4490 (N_4490,N_273,N_568);
nand U4491 (N_4491,N_147,N_1231);
nor U4492 (N_4492,N_1159,N_323);
nand U4493 (N_4493,N_1410,N_2440);
or U4494 (N_4494,N_377,N_300);
nor U4495 (N_4495,N_951,N_2058);
or U4496 (N_4496,N_310,N_2189);
xnor U4497 (N_4497,N_1441,N_2487);
or U4498 (N_4498,N_1029,N_562);
nor U4499 (N_4499,N_399,N_959);
nand U4500 (N_4500,N_1944,N_2484);
and U4501 (N_4501,N_709,N_1937);
or U4502 (N_4502,N_84,N_733);
nor U4503 (N_4503,N_1781,N_2042);
nor U4504 (N_4504,N_1946,N_648);
or U4505 (N_4505,N_81,N_266);
nor U4506 (N_4506,N_1873,N_2440);
nand U4507 (N_4507,N_906,N_926);
and U4508 (N_4508,N_92,N_1370);
xnor U4509 (N_4509,N_2328,N_1642);
and U4510 (N_4510,N_1479,N_1588);
xnor U4511 (N_4511,N_2397,N_1917);
and U4512 (N_4512,N_2286,N_2120);
or U4513 (N_4513,N_700,N_2333);
nor U4514 (N_4514,N_542,N_1856);
nand U4515 (N_4515,N_1288,N_2487);
and U4516 (N_4516,N_2296,N_2371);
or U4517 (N_4517,N_1320,N_2374);
or U4518 (N_4518,N_607,N_1081);
and U4519 (N_4519,N_62,N_60);
and U4520 (N_4520,N_227,N_1944);
and U4521 (N_4521,N_1776,N_162);
xor U4522 (N_4522,N_211,N_1322);
or U4523 (N_4523,N_1364,N_1670);
nand U4524 (N_4524,N_1450,N_1512);
and U4525 (N_4525,N_1368,N_2249);
and U4526 (N_4526,N_2267,N_1260);
nor U4527 (N_4527,N_1261,N_1232);
or U4528 (N_4528,N_519,N_1369);
nand U4529 (N_4529,N_2226,N_2033);
nand U4530 (N_4530,N_109,N_2375);
or U4531 (N_4531,N_425,N_422);
or U4532 (N_4532,N_1227,N_374);
or U4533 (N_4533,N_1415,N_622);
nor U4534 (N_4534,N_1864,N_2037);
nor U4535 (N_4535,N_1422,N_881);
and U4536 (N_4536,N_1762,N_1707);
or U4537 (N_4537,N_728,N_2200);
nor U4538 (N_4538,N_626,N_1553);
and U4539 (N_4539,N_402,N_2192);
nor U4540 (N_4540,N_103,N_792);
nand U4541 (N_4541,N_790,N_1688);
or U4542 (N_4542,N_7,N_456);
nor U4543 (N_4543,N_1562,N_807);
nor U4544 (N_4544,N_867,N_648);
or U4545 (N_4545,N_1106,N_986);
nor U4546 (N_4546,N_1656,N_1738);
nand U4547 (N_4547,N_1729,N_34);
nor U4548 (N_4548,N_1645,N_1094);
and U4549 (N_4549,N_2284,N_607);
or U4550 (N_4550,N_1901,N_2324);
nor U4551 (N_4551,N_1938,N_365);
nand U4552 (N_4552,N_563,N_2199);
nand U4553 (N_4553,N_262,N_2094);
and U4554 (N_4554,N_488,N_1045);
or U4555 (N_4555,N_1653,N_1387);
and U4556 (N_4556,N_407,N_50);
and U4557 (N_4557,N_2391,N_459);
nor U4558 (N_4558,N_157,N_445);
nand U4559 (N_4559,N_1763,N_2071);
or U4560 (N_4560,N_908,N_1196);
and U4561 (N_4561,N_1899,N_656);
or U4562 (N_4562,N_251,N_691);
nand U4563 (N_4563,N_1267,N_2192);
or U4564 (N_4564,N_477,N_1849);
or U4565 (N_4565,N_10,N_1690);
nor U4566 (N_4566,N_1721,N_645);
nand U4567 (N_4567,N_1995,N_300);
nand U4568 (N_4568,N_1289,N_1741);
and U4569 (N_4569,N_1989,N_159);
nand U4570 (N_4570,N_1217,N_469);
or U4571 (N_4571,N_866,N_1819);
and U4572 (N_4572,N_1769,N_1437);
or U4573 (N_4573,N_693,N_2226);
nor U4574 (N_4574,N_1366,N_2299);
nand U4575 (N_4575,N_1729,N_732);
xnor U4576 (N_4576,N_1618,N_365);
and U4577 (N_4577,N_657,N_2190);
nand U4578 (N_4578,N_1080,N_653);
nor U4579 (N_4579,N_72,N_449);
xnor U4580 (N_4580,N_2213,N_321);
nor U4581 (N_4581,N_2302,N_2230);
nand U4582 (N_4582,N_1414,N_85);
nand U4583 (N_4583,N_1785,N_1869);
or U4584 (N_4584,N_1935,N_2158);
xor U4585 (N_4585,N_1114,N_533);
or U4586 (N_4586,N_1895,N_1626);
nand U4587 (N_4587,N_1508,N_1568);
nand U4588 (N_4588,N_28,N_1431);
or U4589 (N_4589,N_535,N_1625);
nor U4590 (N_4590,N_2292,N_2014);
nor U4591 (N_4591,N_878,N_1100);
nand U4592 (N_4592,N_1382,N_1285);
xor U4593 (N_4593,N_1023,N_898);
nand U4594 (N_4594,N_1280,N_1658);
nand U4595 (N_4595,N_1223,N_2340);
and U4596 (N_4596,N_191,N_677);
xor U4597 (N_4597,N_339,N_1025);
and U4598 (N_4598,N_607,N_1493);
nor U4599 (N_4599,N_256,N_2364);
and U4600 (N_4600,N_980,N_1785);
nand U4601 (N_4601,N_2348,N_1782);
xor U4602 (N_4602,N_65,N_1625);
and U4603 (N_4603,N_2050,N_695);
and U4604 (N_4604,N_509,N_1778);
and U4605 (N_4605,N_1200,N_1239);
nand U4606 (N_4606,N_185,N_1169);
xnor U4607 (N_4607,N_595,N_868);
or U4608 (N_4608,N_2341,N_2335);
and U4609 (N_4609,N_1918,N_615);
and U4610 (N_4610,N_545,N_2112);
nor U4611 (N_4611,N_1335,N_1224);
nor U4612 (N_4612,N_1440,N_90);
and U4613 (N_4613,N_42,N_250);
nand U4614 (N_4614,N_2240,N_1805);
nand U4615 (N_4615,N_2322,N_1598);
or U4616 (N_4616,N_502,N_1984);
or U4617 (N_4617,N_578,N_1709);
or U4618 (N_4618,N_396,N_407);
or U4619 (N_4619,N_1055,N_2068);
and U4620 (N_4620,N_654,N_1505);
nor U4621 (N_4621,N_1670,N_1942);
nor U4622 (N_4622,N_833,N_262);
or U4623 (N_4623,N_1697,N_1373);
xnor U4624 (N_4624,N_440,N_2324);
or U4625 (N_4625,N_861,N_342);
or U4626 (N_4626,N_1332,N_2171);
nand U4627 (N_4627,N_2306,N_1626);
and U4628 (N_4628,N_1856,N_340);
or U4629 (N_4629,N_1636,N_1129);
and U4630 (N_4630,N_753,N_971);
nand U4631 (N_4631,N_2420,N_2282);
nand U4632 (N_4632,N_1442,N_1515);
or U4633 (N_4633,N_1032,N_1133);
nand U4634 (N_4634,N_613,N_80);
nor U4635 (N_4635,N_1010,N_1733);
or U4636 (N_4636,N_1982,N_743);
or U4637 (N_4637,N_356,N_430);
nor U4638 (N_4638,N_1400,N_1118);
nor U4639 (N_4639,N_316,N_780);
and U4640 (N_4640,N_1917,N_1596);
nor U4641 (N_4641,N_39,N_2370);
nor U4642 (N_4642,N_944,N_376);
or U4643 (N_4643,N_1861,N_1075);
nand U4644 (N_4644,N_641,N_1494);
nand U4645 (N_4645,N_543,N_947);
or U4646 (N_4646,N_180,N_1435);
and U4647 (N_4647,N_1852,N_504);
nor U4648 (N_4648,N_917,N_1583);
and U4649 (N_4649,N_911,N_1106);
or U4650 (N_4650,N_139,N_635);
nor U4651 (N_4651,N_435,N_160);
and U4652 (N_4652,N_152,N_2385);
nor U4653 (N_4653,N_2157,N_1016);
and U4654 (N_4654,N_1804,N_452);
nand U4655 (N_4655,N_2099,N_670);
nand U4656 (N_4656,N_1953,N_2165);
nand U4657 (N_4657,N_627,N_1672);
or U4658 (N_4658,N_169,N_585);
and U4659 (N_4659,N_1486,N_1470);
or U4660 (N_4660,N_1643,N_1268);
nand U4661 (N_4661,N_556,N_2435);
nor U4662 (N_4662,N_2216,N_1237);
and U4663 (N_4663,N_1454,N_2297);
nand U4664 (N_4664,N_1551,N_691);
nor U4665 (N_4665,N_1896,N_1825);
nand U4666 (N_4666,N_2372,N_1900);
nand U4667 (N_4667,N_1941,N_998);
or U4668 (N_4668,N_2282,N_263);
or U4669 (N_4669,N_2451,N_1922);
nor U4670 (N_4670,N_717,N_1380);
nor U4671 (N_4671,N_1253,N_1597);
nand U4672 (N_4672,N_99,N_738);
and U4673 (N_4673,N_2413,N_1864);
or U4674 (N_4674,N_1686,N_1297);
and U4675 (N_4675,N_354,N_884);
nand U4676 (N_4676,N_2114,N_2161);
or U4677 (N_4677,N_1787,N_309);
or U4678 (N_4678,N_1354,N_1395);
nand U4679 (N_4679,N_1785,N_217);
nand U4680 (N_4680,N_463,N_313);
nand U4681 (N_4681,N_1721,N_811);
nand U4682 (N_4682,N_1877,N_2467);
nor U4683 (N_4683,N_2126,N_2268);
nand U4684 (N_4684,N_1341,N_818);
nor U4685 (N_4685,N_2177,N_975);
or U4686 (N_4686,N_499,N_891);
nand U4687 (N_4687,N_1354,N_2048);
nor U4688 (N_4688,N_2372,N_2486);
nor U4689 (N_4689,N_1747,N_2388);
nor U4690 (N_4690,N_1491,N_1024);
xor U4691 (N_4691,N_1280,N_843);
nand U4692 (N_4692,N_900,N_1416);
and U4693 (N_4693,N_1018,N_1870);
nor U4694 (N_4694,N_1866,N_2203);
or U4695 (N_4695,N_362,N_1512);
or U4696 (N_4696,N_965,N_76);
nand U4697 (N_4697,N_109,N_608);
nand U4698 (N_4698,N_241,N_2393);
nand U4699 (N_4699,N_788,N_2396);
nor U4700 (N_4700,N_331,N_1545);
nand U4701 (N_4701,N_217,N_973);
nor U4702 (N_4702,N_646,N_682);
and U4703 (N_4703,N_215,N_2099);
and U4704 (N_4704,N_1894,N_1829);
or U4705 (N_4705,N_675,N_1528);
nand U4706 (N_4706,N_967,N_37);
or U4707 (N_4707,N_850,N_2336);
or U4708 (N_4708,N_17,N_797);
nor U4709 (N_4709,N_1276,N_1399);
nor U4710 (N_4710,N_484,N_2489);
or U4711 (N_4711,N_64,N_1956);
nor U4712 (N_4712,N_2141,N_2381);
nand U4713 (N_4713,N_696,N_1170);
and U4714 (N_4714,N_1244,N_1566);
and U4715 (N_4715,N_462,N_1289);
or U4716 (N_4716,N_1913,N_840);
and U4717 (N_4717,N_2318,N_359);
nand U4718 (N_4718,N_841,N_1577);
xnor U4719 (N_4719,N_1501,N_989);
or U4720 (N_4720,N_2454,N_104);
nand U4721 (N_4721,N_951,N_31);
or U4722 (N_4722,N_585,N_137);
xnor U4723 (N_4723,N_1558,N_1917);
nand U4724 (N_4724,N_143,N_1379);
nand U4725 (N_4725,N_1746,N_1996);
and U4726 (N_4726,N_1396,N_1556);
nand U4727 (N_4727,N_2377,N_1991);
xnor U4728 (N_4728,N_158,N_1795);
nor U4729 (N_4729,N_2084,N_931);
nand U4730 (N_4730,N_699,N_1005);
nand U4731 (N_4731,N_2042,N_768);
and U4732 (N_4732,N_1289,N_1641);
nand U4733 (N_4733,N_2229,N_2241);
nand U4734 (N_4734,N_1812,N_1142);
nand U4735 (N_4735,N_1225,N_1024);
or U4736 (N_4736,N_2029,N_918);
nand U4737 (N_4737,N_946,N_2416);
or U4738 (N_4738,N_317,N_1627);
or U4739 (N_4739,N_337,N_1937);
nand U4740 (N_4740,N_1785,N_1503);
or U4741 (N_4741,N_759,N_1053);
nand U4742 (N_4742,N_968,N_1582);
and U4743 (N_4743,N_369,N_11);
nand U4744 (N_4744,N_403,N_56);
nand U4745 (N_4745,N_2190,N_1530);
nor U4746 (N_4746,N_133,N_949);
nor U4747 (N_4747,N_1860,N_405);
or U4748 (N_4748,N_1379,N_1490);
nand U4749 (N_4749,N_1149,N_759);
and U4750 (N_4750,N_2401,N_1986);
and U4751 (N_4751,N_165,N_1793);
nor U4752 (N_4752,N_1820,N_288);
and U4753 (N_4753,N_1552,N_531);
nor U4754 (N_4754,N_1438,N_2087);
or U4755 (N_4755,N_889,N_1300);
and U4756 (N_4756,N_2435,N_2176);
or U4757 (N_4757,N_1534,N_334);
or U4758 (N_4758,N_1716,N_187);
and U4759 (N_4759,N_783,N_2222);
and U4760 (N_4760,N_1938,N_1464);
and U4761 (N_4761,N_1837,N_1958);
nand U4762 (N_4762,N_762,N_702);
and U4763 (N_4763,N_267,N_718);
nand U4764 (N_4764,N_229,N_1411);
nand U4765 (N_4765,N_2405,N_260);
nor U4766 (N_4766,N_2197,N_96);
nand U4767 (N_4767,N_2170,N_1508);
and U4768 (N_4768,N_2484,N_2210);
and U4769 (N_4769,N_2379,N_978);
or U4770 (N_4770,N_1367,N_282);
or U4771 (N_4771,N_1578,N_2304);
and U4772 (N_4772,N_400,N_993);
and U4773 (N_4773,N_77,N_2056);
nor U4774 (N_4774,N_1276,N_1325);
and U4775 (N_4775,N_1628,N_2204);
and U4776 (N_4776,N_1238,N_1836);
and U4777 (N_4777,N_1789,N_2009);
and U4778 (N_4778,N_79,N_1444);
nand U4779 (N_4779,N_1526,N_1120);
or U4780 (N_4780,N_550,N_2292);
nand U4781 (N_4781,N_1726,N_1909);
nand U4782 (N_4782,N_1682,N_481);
and U4783 (N_4783,N_1010,N_2297);
nor U4784 (N_4784,N_752,N_1695);
nor U4785 (N_4785,N_662,N_1787);
and U4786 (N_4786,N_930,N_101);
or U4787 (N_4787,N_1111,N_1133);
and U4788 (N_4788,N_2272,N_1734);
nand U4789 (N_4789,N_2339,N_2001);
nand U4790 (N_4790,N_1060,N_1489);
nand U4791 (N_4791,N_995,N_854);
nor U4792 (N_4792,N_1708,N_1856);
or U4793 (N_4793,N_2211,N_1978);
nand U4794 (N_4794,N_628,N_175);
nand U4795 (N_4795,N_6,N_656);
nor U4796 (N_4796,N_2023,N_200);
nand U4797 (N_4797,N_1502,N_2167);
nand U4798 (N_4798,N_2497,N_934);
nor U4799 (N_4799,N_1290,N_1562);
and U4800 (N_4800,N_1443,N_683);
nand U4801 (N_4801,N_2069,N_1709);
and U4802 (N_4802,N_1501,N_1241);
nand U4803 (N_4803,N_2430,N_945);
nand U4804 (N_4804,N_745,N_1859);
or U4805 (N_4805,N_1123,N_2418);
or U4806 (N_4806,N_2222,N_241);
nand U4807 (N_4807,N_1322,N_2017);
nor U4808 (N_4808,N_2454,N_416);
nor U4809 (N_4809,N_1656,N_1279);
or U4810 (N_4810,N_2186,N_796);
and U4811 (N_4811,N_1886,N_2448);
and U4812 (N_4812,N_1538,N_1309);
nand U4813 (N_4813,N_1448,N_2063);
nand U4814 (N_4814,N_2151,N_428);
xnor U4815 (N_4815,N_881,N_2003);
or U4816 (N_4816,N_2115,N_541);
or U4817 (N_4817,N_150,N_1164);
or U4818 (N_4818,N_469,N_2100);
or U4819 (N_4819,N_2042,N_1974);
or U4820 (N_4820,N_1299,N_1180);
nand U4821 (N_4821,N_1288,N_447);
nand U4822 (N_4822,N_249,N_157);
and U4823 (N_4823,N_2410,N_548);
nor U4824 (N_4824,N_36,N_702);
xor U4825 (N_4825,N_759,N_38);
or U4826 (N_4826,N_538,N_1946);
nor U4827 (N_4827,N_1911,N_853);
or U4828 (N_4828,N_1740,N_598);
or U4829 (N_4829,N_1205,N_932);
nor U4830 (N_4830,N_1969,N_1730);
and U4831 (N_4831,N_215,N_1879);
xor U4832 (N_4832,N_1076,N_2485);
nand U4833 (N_4833,N_1342,N_1778);
nor U4834 (N_4834,N_2305,N_262);
nand U4835 (N_4835,N_2380,N_700);
nand U4836 (N_4836,N_1352,N_2046);
and U4837 (N_4837,N_1598,N_2197);
and U4838 (N_4838,N_1951,N_2223);
nand U4839 (N_4839,N_365,N_2032);
xnor U4840 (N_4840,N_2054,N_923);
and U4841 (N_4841,N_1851,N_990);
or U4842 (N_4842,N_2119,N_717);
and U4843 (N_4843,N_696,N_2269);
nand U4844 (N_4844,N_618,N_1054);
nand U4845 (N_4845,N_2314,N_535);
and U4846 (N_4846,N_253,N_1225);
nand U4847 (N_4847,N_718,N_1981);
xnor U4848 (N_4848,N_1132,N_2425);
xnor U4849 (N_4849,N_928,N_478);
or U4850 (N_4850,N_133,N_1954);
and U4851 (N_4851,N_100,N_1032);
nand U4852 (N_4852,N_499,N_2320);
and U4853 (N_4853,N_316,N_370);
nand U4854 (N_4854,N_2211,N_1623);
nand U4855 (N_4855,N_743,N_893);
nor U4856 (N_4856,N_2107,N_883);
and U4857 (N_4857,N_235,N_2476);
and U4858 (N_4858,N_1435,N_1237);
and U4859 (N_4859,N_721,N_789);
and U4860 (N_4860,N_2360,N_496);
or U4861 (N_4861,N_2045,N_1985);
nand U4862 (N_4862,N_1356,N_2150);
nor U4863 (N_4863,N_2344,N_970);
or U4864 (N_4864,N_1171,N_1875);
nand U4865 (N_4865,N_1630,N_2254);
nor U4866 (N_4866,N_1898,N_1249);
nor U4867 (N_4867,N_2310,N_514);
xnor U4868 (N_4868,N_1061,N_1096);
or U4869 (N_4869,N_1849,N_1641);
nor U4870 (N_4870,N_1076,N_1481);
nor U4871 (N_4871,N_421,N_368);
and U4872 (N_4872,N_460,N_2492);
nor U4873 (N_4873,N_119,N_1717);
nand U4874 (N_4874,N_2073,N_870);
and U4875 (N_4875,N_1624,N_1794);
or U4876 (N_4876,N_613,N_2350);
and U4877 (N_4877,N_402,N_513);
or U4878 (N_4878,N_2140,N_1899);
and U4879 (N_4879,N_1485,N_2164);
nand U4880 (N_4880,N_993,N_2164);
xor U4881 (N_4881,N_2461,N_2459);
nand U4882 (N_4882,N_1209,N_1450);
nand U4883 (N_4883,N_2309,N_265);
and U4884 (N_4884,N_1874,N_1148);
nor U4885 (N_4885,N_1537,N_1562);
and U4886 (N_4886,N_2043,N_2252);
nor U4887 (N_4887,N_2121,N_1115);
nor U4888 (N_4888,N_206,N_1290);
and U4889 (N_4889,N_1925,N_1172);
and U4890 (N_4890,N_1816,N_78);
and U4891 (N_4891,N_2215,N_2464);
and U4892 (N_4892,N_678,N_1072);
nor U4893 (N_4893,N_910,N_532);
and U4894 (N_4894,N_1650,N_1906);
nor U4895 (N_4895,N_224,N_174);
nor U4896 (N_4896,N_557,N_535);
and U4897 (N_4897,N_758,N_184);
and U4898 (N_4898,N_2050,N_2127);
or U4899 (N_4899,N_2042,N_1446);
or U4900 (N_4900,N_1916,N_1131);
or U4901 (N_4901,N_1260,N_2436);
or U4902 (N_4902,N_1011,N_1402);
and U4903 (N_4903,N_2220,N_2399);
nor U4904 (N_4904,N_2394,N_1159);
and U4905 (N_4905,N_1438,N_1683);
nand U4906 (N_4906,N_1991,N_322);
nor U4907 (N_4907,N_1639,N_1446);
or U4908 (N_4908,N_2245,N_621);
nor U4909 (N_4909,N_2416,N_112);
nand U4910 (N_4910,N_2055,N_1995);
or U4911 (N_4911,N_1369,N_679);
nand U4912 (N_4912,N_1975,N_567);
and U4913 (N_4913,N_2157,N_1004);
and U4914 (N_4914,N_384,N_1683);
nor U4915 (N_4915,N_1134,N_125);
nand U4916 (N_4916,N_1838,N_108);
nand U4917 (N_4917,N_2454,N_1443);
and U4918 (N_4918,N_2149,N_603);
and U4919 (N_4919,N_973,N_783);
or U4920 (N_4920,N_1414,N_1007);
or U4921 (N_4921,N_830,N_1704);
and U4922 (N_4922,N_301,N_1331);
and U4923 (N_4923,N_1290,N_817);
or U4924 (N_4924,N_58,N_1872);
xnor U4925 (N_4925,N_1373,N_297);
nor U4926 (N_4926,N_170,N_1439);
nand U4927 (N_4927,N_1589,N_455);
or U4928 (N_4928,N_248,N_172);
or U4929 (N_4929,N_1440,N_1478);
nand U4930 (N_4930,N_1201,N_512);
and U4931 (N_4931,N_2163,N_1181);
and U4932 (N_4932,N_1403,N_2320);
nand U4933 (N_4933,N_1866,N_1507);
nor U4934 (N_4934,N_1447,N_1934);
nor U4935 (N_4935,N_1908,N_791);
or U4936 (N_4936,N_1782,N_2474);
xor U4937 (N_4937,N_1356,N_1700);
or U4938 (N_4938,N_2410,N_513);
nor U4939 (N_4939,N_1579,N_1343);
nand U4940 (N_4940,N_463,N_1892);
nor U4941 (N_4941,N_2084,N_1452);
or U4942 (N_4942,N_473,N_458);
nor U4943 (N_4943,N_1492,N_145);
or U4944 (N_4944,N_1232,N_418);
or U4945 (N_4945,N_2499,N_1308);
or U4946 (N_4946,N_541,N_154);
nor U4947 (N_4947,N_580,N_274);
xor U4948 (N_4948,N_648,N_576);
nand U4949 (N_4949,N_971,N_520);
and U4950 (N_4950,N_1025,N_2096);
or U4951 (N_4951,N_311,N_829);
nand U4952 (N_4952,N_2485,N_2429);
nor U4953 (N_4953,N_1749,N_219);
or U4954 (N_4954,N_1424,N_2358);
nand U4955 (N_4955,N_594,N_1804);
nand U4956 (N_4956,N_1395,N_672);
or U4957 (N_4957,N_2112,N_914);
or U4958 (N_4958,N_218,N_1590);
and U4959 (N_4959,N_165,N_1790);
and U4960 (N_4960,N_231,N_2100);
nand U4961 (N_4961,N_2042,N_2082);
and U4962 (N_4962,N_2297,N_708);
or U4963 (N_4963,N_751,N_845);
and U4964 (N_4964,N_487,N_1204);
and U4965 (N_4965,N_747,N_198);
nand U4966 (N_4966,N_239,N_920);
and U4967 (N_4967,N_2418,N_1283);
nor U4968 (N_4968,N_1426,N_2096);
nand U4969 (N_4969,N_752,N_935);
nand U4970 (N_4970,N_2431,N_347);
and U4971 (N_4971,N_1923,N_1220);
and U4972 (N_4972,N_2233,N_2491);
and U4973 (N_4973,N_2225,N_149);
nor U4974 (N_4974,N_2444,N_493);
nor U4975 (N_4975,N_889,N_988);
and U4976 (N_4976,N_447,N_254);
nor U4977 (N_4977,N_1410,N_1752);
or U4978 (N_4978,N_2189,N_373);
and U4979 (N_4979,N_1859,N_1749);
nand U4980 (N_4980,N_30,N_1963);
and U4981 (N_4981,N_88,N_1546);
nand U4982 (N_4982,N_134,N_2085);
xor U4983 (N_4983,N_542,N_282);
nor U4984 (N_4984,N_731,N_1047);
nand U4985 (N_4985,N_619,N_2257);
nor U4986 (N_4986,N_1508,N_2369);
nand U4987 (N_4987,N_1910,N_347);
nor U4988 (N_4988,N_1482,N_95);
nor U4989 (N_4989,N_1919,N_1799);
or U4990 (N_4990,N_1205,N_2324);
nand U4991 (N_4991,N_513,N_1182);
nor U4992 (N_4992,N_106,N_223);
and U4993 (N_4993,N_964,N_1160);
and U4994 (N_4994,N_1749,N_1200);
nand U4995 (N_4995,N_1793,N_53);
nor U4996 (N_4996,N_2162,N_1449);
or U4997 (N_4997,N_69,N_1889);
and U4998 (N_4998,N_2298,N_927);
and U4999 (N_4999,N_1636,N_728);
nor U5000 (N_5000,N_3590,N_2893);
nand U5001 (N_5001,N_2716,N_3110);
or U5002 (N_5002,N_4737,N_4046);
nor U5003 (N_5003,N_2715,N_3073);
nand U5004 (N_5004,N_4901,N_4178);
or U5005 (N_5005,N_2759,N_4564);
and U5006 (N_5006,N_3000,N_4187);
and U5007 (N_5007,N_4048,N_2573);
or U5008 (N_5008,N_4994,N_3809);
xor U5009 (N_5009,N_4806,N_4256);
xor U5010 (N_5010,N_4955,N_4555);
nand U5011 (N_5011,N_4462,N_3556);
nand U5012 (N_5012,N_4613,N_2500);
nand U5013 (N_5013,N_3818,N_3813);
or U5014 (N_5014,N_4467,N_4637);
nand U5015 (N_5015,N_3393,N_4371);
and U5016 (N_5016,N_2965,N_2852);
nor U5017 (N_5017,N_2723,N_2648);
nand U5018 (N_5018,N_2751,N_3721);
and U5019 (N_5019,N_2773,N_4592);
nand U5020 (N_5020,N_4952,N_4612);
and U5021 (N_5021,N_4846,N_3288);
or U5022 (N_5022,N_4760,N_3681);
nand U5023 (N_5023,N_3678,N_4535);
nor U5024 (N_5024,N_2941,N_3289);
nor U5025 (N_5025,N_3299,N_3364);
nor U5026 (N_5026,N_3359,N_4464);
or U5027 (N_5027,N_4608,N_4271);
nor U5028 (N_5028,N_3282,N_3932);
and U5029 (N_5029,N_3210,N_2671);
nand U5030 (N_5030,N_4505,N_2692);
nor U5031 (N_5031,N_2607,N_2824);
or U5032 (N_5032,N_4799,N_2653);
nor U5033 (N_5033,N_4215,N_2915);
or U5034 (N_5034,N_4122,N_4146);
or U5035 (N_5035,N_2705,N_4288);
and U5036 (N_5036,N_3736,N_4330);
and U5037 (N_5037,N_2986,N_4527);
nand U5038 (N_5038,N_4301,N_3400);
or U5039 (N_5039,N_3326,N_3330);
nand U5040 (N_5040,N_2518,N_2679);
or U5041 (N_5041,N_3455,N_2509);
nor U5042 (N_5042,N_4919,N_4318);
or U5043 (N_5043,N_3254,N_3952);
and U5044 (N_5044,N_4282,N_2588);
nand U5045 (N_5045,N_3841,N_4896);
and U5046 (N_5046,N_3948,N_3217);
and U5047 (N_5047,N_3941,N_3019);
nand U5048 (N_5048,N_3921,N_3543);
and U5049 (N_5049,N_4653,N_4925);
nand U5050 (N_5050,N_3443,N_3670);
or U5051 (N_5051,N_3188,N_4480);
and U5052 (N_5052,N_2961,N_4228);
nand U5053 (N_5053,N_4735,N_3204);
or U5054 (N_5054,N_4396,N_4913);
and U5055 (N_5055,N_4611,N_4320);
or U5056 (N_5056,N_2842,N_4112);
and U5057 (N_5057,N_3585,N_3270);
nand U5058 (N_5058,N_3738,N_3478);
or U5059 (N_5059,N_2718,N_4699);
nand U5060 (N_5060,N_3854,N_3870);
or U5061 (N_5061,N_2882,N_2950);
or U5062 (N_5062,N_3387,N_4574);
and U5063 (N_5063,N_4410,N_2779);
or U5064 (N_5064,N_3769,N_4807);
and U5065 (N_5065,N_4559,N_3296);
nor U5066 (N_5066,N_4784,N_4606);
and U5067 (N_5067,N_4314,N_3576);
or U5068 (N_5068,N_2974,N_3397);
nand U5069 (N_5069,N_3316,N_2778);
nor U5070 (N_5070,N_4227,N_3349);
or U5071 (N_5071,N_4299,N_4429);
nor U5072 (N_5072,N_4563,N_3242);
and U5073 (N_5073,N_4268,N_3713);
or U5074 (N_5074,N_3343,N_3466);
nor U5075 (N_5075,N_3682,N_4289);
nand U5076 (N_5076,N_2546,N_4625);
or U5077 (N_5077,N_4496,N_3194);
and U5078 (N_5078,N_4249,N_2649);
nand U5079 (N_5079,N_4181,N_3418);
and U5080 (N_5080,N_3355,N_4375);
and U5081 (N_5081,N_4381,N_3415);
nand U5082 (N_5082,N_2504,N_4786);
nor U5083 (N_5083,N_4999,N_3863);
nor U5084 (N_5084,N_4109,N_2939);
nand U5085 (N_5085,N_2952,N_4114);
nor U5086 (N_5086,N_4879,N_3532);
nor U5087 (N_5087,N_2642,N_4595);
nand U5088 (N_5088,N_4241,N_4804);
nor U5089 (N_5089,N_4317,N_4695);
nor U5090 (N_5090,N_3022,N_3832);
and U5091 (N_5091,N_2739,N_4300);
and U5092 (N_5092,N_4648,N_3431);
nor U5093 (N_5093,N_3665,N_2897);
nor U5094 (N_5094,N_4024,N_2665);
nand U5095 (N_5095,N_3584,N_3061);
or U5096 (N_5096,N_3561,N_4027);
and U5097 (N_5097,N_3843,N_4588);
or U5098 (N_5098,N_4091,N_4295);
and U5099 (N_5099,N_3929,N_3926);
or U5100 (N_5100,N_3512,N_3928);
nand U5101 (N_5101,N_3118,N_2514);
nor U5102 (N_5102,N_3341,N_2569);
and U5103 (N_5103,N_4344,N_3554);
or U5104 (N_5104,N_4622,N_4504);
nor U5105 (N_5105,N_3141,N_4517);
nor U5106 (N_5106,N_4058,N_2922);
nor U5107 (N_5107,N_4556,N_2972);
nand U5108 (N_5108,N_2626,N_4845);
nor U5109 (N_5109,N_3967,N_2964);
or U5110 (N_5110,N_3396,N_4746);
nand U5111 (N_5111,N_4508,N_3291);
or U5112 (N_5112,N_4500,N_3087);
nor U5113 (N_5113,N_3571,N_2937);
or U5114 (N_5114,N_4147,N_4275);
or U5115 (N_5115,N_4800,N_2808);
or U5116 (N_5116,N_4547,N_4190);
nor U5117 (N_5117,N_4420,N_3138);
nor U5118 (N_5118,N_4685,N_3889);
and U5119 (N_5119,N_2877,N_3435);
nand U5120 (N_5120,N_4149,N_2785);
and U5121 (N_5121,N_3862,N_3465);
nor U5122 (N_5122,N_3759,N_4053);
and U5123 (N_5123,N_4507,N_3773);
or U5124 (N_5124,N_3222,N_3143);
and U5125 (N_5125,N_4236,N_2566);
and U5126 (N_5126,N_3156,N_3895);
or U5127 (N_5127,N_4298,N_4473);
nor U5128 (N_5128,N_2823,N_4322);
or U5129 (N_5129,N_4132,N_2874);
or U5130 (N_5130,N_4033,N_2536);
and U5131 (N_5131,N_2782,N_4932);
nand U5132 (N_5132,N_3412,N_4356);
nor U5133 (N_5133,N_4198,N_3329);
nand U5134 (N_5134,N_4022,N_4051);
and U5135 (N_5135,N_2859,N_2756);
xnor U5136 (N_5136,N_3859,N_3972);
nor U5137 (N_5137,N_2737,N_3109);
nor U5138 (N_5138,N_4663,N_3399);
and U5139 (N_5139,N_4970,N_4544);
or U5140 (N_5140,N_4392,N_3882);
or U5141 (N_5141,N_4321,N_4394);
and U5142 (N_5142,N_3142,N_4003);
nand U5143 (N_5143,N_3215,N_2887);
xor U5144 (N_5144,N_3055,N_3710);
or U5145 (N_5145,N_3758,N_3059);
nor U5146 (N_5146,N_4414,N_2867);
or U5147 (N_5147,N_4313,N_4922);
and U5148 (N_5148,N_4627,N_2530);
and U5149 (N_5149,N_4454,N_4738);
xor U5150 (N_5150,N_4117,N_3776);
nor U5151 (N_5151,N_3559,N_4883);
nand U5152 (N_5152,N_4080,N_4002);
and U5153 (N_5153,N_2892,N_3408);
nor U5154 (N_5154,N_2969,N_3674);
nor U5155 (N_5155,N_3265,N_4809);
xor U5156 (N_5156,N_3508,N_3409);
nor U5157 (N_5157,N_3896,N_3957);
or U5158 (N_5158,N_2763,N_3199);
and U5159 (N_5159,N_3865,N_3629);
or U5160 (N_5160,N_3595,N_2647);
nor U5161 (N_5161,N_4078,N_3542);
nand U5162 (N_5162,N_2562,N_3735);
and U5163 (N_5163,N_3078,N_3521);
or U5164 (N_5164,N_3149,N_2931);
and U5165 (N_5165,N_3233,N_3088);
nand U5166 (N_5166,N_3120,N_3175);
nand U5167 (N_5167,N_4283,N_3891);
or U5168 (N_5168,N_4459,N_2698);
and U5169 (N_5169,N_4635,N_4667);
nor U5170 (N_5170,N_3371,N_4756);
and U5171 (N_5171,N_3636,N_3017);
nand U5172 (N_5172,N_3523,N_4810);
or U5173 (N_5173,N_3258,N_2899);
and U5174 (N_5174,N_3018,N_3557);
and U5175 (N_5175,N_3534,N_2989);
or U5176 (N_5176,N_4841,N_2829);
nor U5177 (N_5177,N_4927,N_3781);
nand U5178 (N_5178,N_3107,N_4175);
nand U5179 (N_5179,N_4533,N_4662);
or U5180 (N_5180,N_4520,N_3519);
nor U5181 (N_5181,N_3652,N_2855);
xnor U5182 (N_5182,N_3385,N_3866);
or U5183 (N_5183,N_4714,N_4052);
nor U5184 (N_5184,N_3626,N_4619);
xnor U5185 (N_5185,N_3915,N_4453);
nand U5186 (N_5186,N_3894,N_3111);
nand U5187 (N_5187,N_3064,N_4793);
and U5188 (N_5188,N_4775,N_3838);
or U5189 (N_5189,N_3367,N_4866);
and U5190 (N_5190,N_3406,N_4539);
and U5191 (N_5191,N_3731,N_3038);
nand U5192 (N_5192,N_4794,N_3795);
nor U5193 (N_5193,N_4551,N_3755);
nor U5194 (N_5194,N_4250,N_4047);
xnor U5195 (N_5195,N_3098,N_4749);
and U5196 (N_5196,N_3885,N_3427);
nand U5197 (N_5197,N_2582,N_2645);
nand U5198 (N_5198,N_4863,N_3065);
nand U5199 (N_5199,N_3789,N_4200);
or U5200 (N_5200,N_3322,N_3819);
and U5201 (N_5201,N_4808,N_4119);
nor U5202 (N_5202,N_4221,N_2979);
or U5203 (N_5203,N_4006,N_2574);
and U5204 (N_5204,N_4857,N_2564);
or U5205 (N_5205,N_4718,N_3995);
nor U5206 (N_5206,N_3839,N_3126);
or U5207 (N_5207,N_2553,N_3220);
or U5208 (N_5208,N_2538,N_3012);
nor U5209 (N_5209,N_2809,N_4944);
nand U5210 (N_5210,N_3504,N_4858);
and U5211 (N_5211,N_3032,N_3499);
nand U5212 (N_5212,N_4580,N_2516);
or U5213 (N_5213,N_4378,N_4797);
and U5214 (N_5214,N_2749,N_4696);
nor U5215 (N_5215,N_3628,N_4272);
or U5216 (N_5216,N_4329,N_2900);
and U5217 (N_5217,N_2620,N_3043);
and U5218 (N_5218,N_4722,N_2799);
and U5219 (N_5219,N_2924,N_3704);
and U5220 (N_5220,N_3760,N_3572);
and U5221 (N_5221,N_2643,N_3328);
nor U5222 (N_5222,N_2858,N_3606);
and U5223 (N_5223,N_4554,N_4031);
and U5224 (N_5224,N_3497,N_4964);
or U5225 (N_5225,N_4805,N_3315);
nor U5226 (N_5226,N_2850,N_4018);
nand U5227 (N_5227,N_4016,N_3487);
nand U5228 (N_5228,N_3570,N_3121);
and U5229 (N_5229,N_2521,N_4975);
and U5230 (N_5230,N_3583,N_3845);
and U5231 (N_5231,N_4099,N_3679);
and U5232 (N_5232,N_4801,N_3351);
or U5233 (N_5233,N_3611,N_4310);
nand U5234 (N_5234,N_2890,N_3276);
nand U5235 (N_5235,N_4391,N_2847);
nand U5236 (N_5236,N_3148,N_3671);
or U5237 (N_5237,N_3072,N_3688);
or U5238 (N_5238,N_3428,N_4812);
nor U5239 (N_5239,N_3568,N_4816);
nand U5240 (N_5240,N_4401,N_4363);
and U5241 (N_5241,N_4012,N_3963);
or U5242 (N_5242,N_3327,N_4292);
and U5243 (N_5243,N_2680,N_3546);
and U5244 (N_5244,N_4617,N_2810);
nor U5245 (N_5245,N_2513,N_3339);
or U5246 (N_5246,N_4055,N_4361);
or U5247 (N_5247,N_4509,N_4706);
or U5248 (N_5248,N_4946,N_4614);
nand U5249 (N_5249,N_3469,N_4357);
and U5250 (N_5250,N_2701,N_2519);
nor U5251 (N_5251,N_2896,N_4890);
and U5252 (N_5252,N_2730,N_4790);
or U5253 (N_5253,N_4302,N_4503);
nand U5254 (N_5254,N_2948,N_4803);
nand U5255 (N_5255,N_2868,N_4729);
nor U5256 (N_5256,N_4972,N_2787);
nor U5257 (N_5257,N_3998,N_4094);
or U5258 (N_5258,N_2529,N_3003);
nand U5259 (N_5259,N_4118,N_3638);
and U5260 (N_5260,N_4636,N_4102);
nand U5261 (N_5261,N_4001,N_4629);
nor U5262 (N_5262,N_2828,N_4213);
or U5263 (N_5263,N_4789,N_4083);
nand U5264 (N_5264,N_4713,N_2789);
and U5265 (N_5265,N_4628,N_3205);
nor U5266 (N_5266,N_4023,N_2605);
nand U5267 (N_5267,N_3659,N_4871);
and U5268 (N_5268,N_3305,N_2638);
and U5269 (N_5269,N_4561,N_4129);
nor U5270 (N_5270,N_4212,N_4367);
nor U5271 (N_5271,N_4202,N_4924);
or U5272 (N_5272,N_4416,N_2758);
nor U5273 (N_5273,N_4502,N_4769);
nor U5274 (N_5274,N_3284,N_4582);
or U5275 (N_5275,N_3268,N_3810);
or U5276 (N_5276,N_4290,N_4049);
nor U5277 (N_5277,N_4693,N_2794);
nor U5278 (N_5278,N_4189,N_3293);
or U5279 (N_5279,N_2693,N_3261);
nor U5280 (N_5280,N_2619,N_2780);
and U5281 (N_5281,N_2838,N_4264);
or U5282 (N_5282,N_4079,N_4604);
nand U5283 (N_5283,N_2677,N_2517);
or U5284 (N_5284,N_2926,N_4216);
nand U5285 (N_5285,N_2681,N_3058);
or U5286 (N_5286,N_4907,N_2938);
nor U5287 (N_5287,N_4751,N_4069);
or U5288 (N_5288,N_4222,N_2689);
nand U5289 (N_5289,N_3358,N_3023);
and U5290 (N_5290,N_2754,N_3250);
nand U5291 (N_5291,N_2916,N_3286);
or U5292 (N_5292,N_4245,N_3493);
or U5293 (N_5293,N_4203,N_2770);
nand U5294 (N_5294,N_4350,N_3514);
and U5295 (N_5295,N_3986,N_3698);
and U5296 (N_5296,N_4899,N_3575);
and U5297 (N_5297,N_2951,N_2578);
nor U5298 (N_5298,N_3770,N_4225);
or U5299 (N_5299,N_3026,N_2929);
nand U5300 (N_5300,N_4585,N_3647);
nand U5301 (N_5301,N_3165,N_4352);
or U5302 (N_5302,N_2658,N_4926);
or U5303 (N_5303,N_3962,N_3039);
nor U5304 (N_5304,N_3566,N_3475);
and U5305 (N_5305,N_3861,N_4020);
and U5306 (N_5306,N_4851,N_3388);
or U5307 (N_5307,N_2609,N_3005);
or U5308 (N_5308,N_3161,N_3008);
or U5309 (N_5309,N_3878,N_3052);
or U5310 (N_5310,N_4827,N_2728);
or U5311 (N_5311,N_3742,N_4639);
nor U5312 (N_5312,N_3977,N_4427);
nor U5313 (N_5313,N_4757,N_4597);
and U5314 (N_5314,N_3310,N_2800);
nor U5315 (N_5315,N_3906,N_2719);
nor U5316 (N_5316,N_3510,N_3833);
nand U5317 (N_5317,N_3452,N_4340);
or U5318 (N_5318,N_4432,N_3756);
nor U5319 (N_5319,N_3827,N_2703);
and U5320 (N_5320,N_2657,N_4712);
or U5321 (N_5321,N_3613,N_4631);
nor U5322 (N_5322,N_4446,N_4742);
nor U5323 (N_5323,N_4358,N_3164);
or U5324 (N_5324,N_2866,N_2676);
nand U5325 (N_5325,N_2793,N_4188);
nand U5326 (N_5326,N_3292,N_4743);
or U5327 (N_5327,N_3389,N_2735);
nor U5328 (N_5328,N_2981,N_3274);
or U5329 (N_5329,N_3476,N_3916);
and U5330 (N_5330,N_2709,N_4235);
xor U5331 (N_5331,N_4238,N_4115);
nor U5332 (N_5332,N_3528,N_2565);
nor U5333 (N_5333,N_4305,N_3498);
or U5334 (N_5334,N_4121,N_4103);
or U5335 (N_5335,N_2568,N_2544);
nand U5336 (N_5336,N_3004,N_4763);
nand U5337 (N_5337,N_4536,N_4353);
nor U5338 (N_5338,N_4828,N_4686);
or U5339 (N_5339,N_4296,N_4206);
nor U5340 (N_5340,N_3245,N_3836);
or U5341 (N_5341,N_2505,N_3070);
nor U5342 (N_5342,N_4711,N_4834);
nand U5343 (N_5343,N_3700,N_3190);
nand U5344 (N_5344,N_3035,N_4707);
nor U5345 (N_5345,N_4728,N_4398);
xor U5346 (N_5346,N_3486,N_4887);
nor U5347 (N_5347,N_2590,N_2987);
nor U5348 (N_5348,N_4985,N_4566);
nor U5349 (N_5349,N_4408,N_4258);
nand U5350 (N_5350,N_2559,N_3746);
nand U5351 (N_5351,N_4484,N_4874);
xor U5352 (N_5352,N_3162,N_4077);
or U5353 (N_5353,N_4573,N_3259);
nand U5354 (N_5354,N_3122,N_4439);
xor U5355 (N_5355,N_3708,N_2611);
nand U5356 (N_5356,N_3066,N_2833);
nor U5357 (N_5357,N_4720,N_4873);
nand U5358 (N_5358,N_3483,N_4948);
and U5359 (N_5359,N_3037,N_3015);
and U5360 (N_5360,N_3979,N_3170);
nor U5361 (N_5361,N_4204,N_3273);
or U5362 (N_5362,N_3285,N_4577);
nand U5363 (N_5363,N_2966,N_3256);
nand U5364 (N_5364,N_3235,N_3287);
or U5365 (N_5365,N_3548,N_4560);
nand U5366 (N_5366,N_3944,N_3201);
nor U5367 (N_5367,N_4602,N_3640);
nor U5368 (N_5368,N_4997,N_2869);
nand U5369 (N_5369,N_3530,N_2819);
or U5370 (N_5370,N_4589,N_2666);
nor U5371 (N_5371,N_4953,N_3732);
or U5372 (N_5372,N_3971,N_2876);
nor U5373 (N_5373,N_4687,N_2912);
nand U5374 (N_5374,N_4716,N_2683);
nor U5375 (N_5375,N_3232,N_4095);
nor U5376 (N_5376,N_3216,N_3612);
xor U5377 (N_5377,N_3042,N_3381);
nor U5378 (N_5378,N_4645,N_3077);
or U5379 (N_5379,N_3306,N_2860);
nor U5380 (N_5380,N_3701,N_3593);
and U5381 (N_5381,N_3344,N_4587);
nand U5382 (N_5382,N_3390,N_4962);
or U5383 (N_5383,N_4165,N_3227);
nand U5384 (N_5384,N_2772,N_3272);
and U5385 (N_5385,N_3459,N_4253);
and U5386 (N_5386,N_3696,N_4092);
xor U5387 (N_5387,N_4159,N_3569);
or U5388 (N_5388,N_4116,N_4898);
nor U5389 (N_5389,N_4017,N_4355);
and U5390 (N_5390,N_4174,N_4428);
or U5391 (N_5391,N_4399,N_3453);
nand U5392 (N_5392,N_3106,N_3127);
or U5393 (N_5393,N_4123,N_3646);
or U5394 (N_5394,N_2743,N_3822);
and U5395 (N_5395,N_4704,N_4261);
or U5396 (N_5396,N_3900,N_3423);
nor U5397 (N_5397,N_3604,N_4939);
nor U5398 (N_5398,N_4486,N_2904);
nor U5399 (N_5399,N_3890,N_4552);
nor U5400 (N_5400,N_4232,N_4549);
nand U5401 (N_5401,N_3847,N_3625);
or U5402 (N_5402,N_4059,N_3404);
or U5403 (N_5403,N_4967,N_2978);
nor U5404 (N_5404,N_3262,N_4651);
and U5405 (N_5405,N_4008,N_4374);
nand U5406 (N_5406,N_4067,N_2747);
nand U5407 (N_5407,N_2732,N_3560);
nor U5408 (N_5408,N_3353,N_2790);
nand U5409 (N_5409,N_3226,N_3132);
xor U5410 (N_5410,N_4700,N_4475);
nor U5411 (N_5411,N_4385,N_2925);
or U5412 (N_5412,N_3672,N_4279);
nor U5413 (N_5413,N_3115,N_3153);
nand U5414 (N_5414,N_3936,N_4445);
or U5415 (N_5415,N_2707,N_3183);
nand U5416 (N_5416,N_3438,N_3980);
nand U5417 (N_5417,N_3771,N_3211);
and U5418 (N_5418,N_4324,N_4902);
and U5419 (N_5419,N_2627,N_3814);
nand U5420 (N_5420,N_3231,N_4598);
nor U5421 (N_5421,N_3361,N_4194);
and U5422 (N_5422,N_4242,N_3757);
nor U5423 (N_5423,N_4425,N_3807);
nand U5424 (N_5424,N_3808,N_4940);
and U5425 (N_5425,N_4753,N_2587);
or U5426 (N_5426,N_4262,N_4669);
or U5427 (N_5427,N_3744,N_3166);
and U5428 (N_5428,N_3457,N_2555);
nor U5429 (N_5429,N_3405,N_3494);
nor U5430 (N_5430,N_3102,N_2920);
or U5431 (N_5431,N_4491,N_4167);
nor U5432 (N_5432,N_3860,N_3045);
or U5433 (N_5433,N_2910,N_4196);
nor U5434 (N_5434,N_3145,N_3116);
or U5435 (N_5435,N_4652,N_3100);
or U5436 (N_5436,N_3869,N_4820);
nor U5437 (N_5437,N_2724,N_4412);
and U5438 (N_5438,N_4528,N_3761);
nor U5439 (N_5439,N_4331,N_4442);
nand U5440 (N_5440,N_2746,N_2632);
and U5441 (N_5441,N_4770,N_4377);
or U5442 (N_5442,N_3345,N_4297);
and U5443 (N_5443,N_3252,N_2977);
or U5444 (N_5444,N_3527,N_4831);
nor U5445 (N_5445,N_4444,N_2767);
nor U5446 (N_5446,N_2820,N_4584);
and U5447 (N_5447,N_3937,N_4506);
nand U5448 (N_5448,N_4973,N_2963);
or U5449 (N_5449,N_4019,N_2599);
nand U5450 (N_5450,N_4307,N_4014);
or U5451 (N_5451,N_4021,N_3420);
or U5452 (N_5452,N_3634,N_3034);
nor U5453 (N_5453,N_4393,N_2710);
and U5454 (N_5454,N_3551,N_2523);
and U5455 (N_5455,N_4862,N_4701);
or U5456 (N_5456,N_4191,N_4068);
nand U5457 (N_5457,N_3752,N_2615);
and U5458 (N_5458,N_3942,N_4237);
or U5459 (N_5459,N_2670,N_4193);
and U5460 (N_5460,N_4802,N_3867);
nand U5461 (N_5461,N_4510,N_3692);
or U5462 (N_5462,N_4060,N_4255);
or U5463 (N_5463,N_3723,N_4692);
or U5464 (N_5464,N_3144,N_4007);
and U5465 (N_5465,N_4452,N_3223);
and U5466 (N_5466,N_3357,N_2750);
nand U5467 (N_5467,N_3354,N_3655);
and U5468 (N_5468,N_4097,N_2903);
nor U5469 (N_5469,N_3207,N_3275);
and U5470 (N_5470,N_3991,N_2621);
nor U5471 (N_5471,N_3642,N_2713);
and U5472 (N_5472,N_4918,N_4140);
nand U5473 (N_5473,N_4572,N_4882);
nor U5474 (N_5474,N_4265,N_3996);
or U5475 (N_5475,N_3880,N_3582);
or U5476 (N_5476,N_4571,N_4347);
nor U5477 (N_5477,N_2932,N_3128);
xor U5478 (N_5478,N_3380,N_2947);
or U5479 (N_5479,N_3464,N_3374);
and U5480 (N_5480,N_3535,N_3950);
or U5481 (N_5481,N_4942,N_3366);
nand U5482 (N_5482,N_2909,N_3976);
nand U5483 (N_5483,N_4826,N_4404);
and U5484 (N_5484,N_4610,N_4649);
or U5485 (N_5485,N_4618,N_3439);
nor U5486 (N_5486,N_2629,N_4817);
nor U5487 (N_5487,N_2945,N_4487);
xor U5488 (N_5488,N_4661,N_4673);
nand U5489 (N_5489,N_4721,N_3208);
nand U5490 (N_5490,N_4715,N_3373);
nor U5491 (N_5491,N_3150,N_4773);
nand U5492 (N_5492,N_4740,N_3785);
or U5493 (N_5493,N_3002,N_3981);
and U5494 (N_5494,N_4727,N_4133);
nor U5495 (N_5495,N_3167,N_4678);
nor U5496 (N_5496,N_3383,N_4380);
nor U5497 (N_5497,N_4426,N_3080);
nand U5498 (N_5498,N_3741,N_3522);
nor U5499 (N_5499,N_4087,N_4821);
nor U5500 (N_5500,N_4872,N_2875);
or U5501 (N_5501,N_4935,N_4739);
or U5502 (N_5502,N_3482,N_3021);
nand U5503 (N_5503,N_4304,N_2864);
or U5504 (N_5504,N_4066,N_4818);
or U5505 (N_5505,N_2744,N_4254);
nor U5506 (N_5506,N_2843,N_3685);
nor U5507 (N_5507,N_3084,N_2879);
nand U5508 (N_5508,N_3821,N_3083);
or U5509 (N_5509,N_2851,N_2672);
or U5510 (N_5510,N_3804,N_3673);
nand U5511 (N_5511,N_3421,N_2944);
or U5512 (N_5512,N_4867,N_3269);
nor U5513 (N_5513,N_3488,N_3563);
or U5514 (N_5514,N_4176,N_2745);
nor U5515 (N_5515,N_3520,N_3597);
nor U5516 (N_5516,N_4463,N_3099);
nand U5517 (N_5517,N_2606,N_3680);
or U5518 (N_5518,N_2918,N_3537);
or U5519 (N_5519,N_4759,N_4379);
nand U5520 (N_5520,N_4912,N_3044);
nand U5521 (N_5521,N_4941,N_2613);
nor U5522 (N_5522,N_4885,N_3263);
or U5523 (N_5523,N_3711,N_3683);
nand U5524 (N_5524,N_4346,N_4220);
nor U5525 (N_5525,N_4880,N_2596);
or U5526 (N_5526,N_3441,N_2992);
nand U5527 (N_5527,N_4151,N_4516);
and U5528 (N_5528,N_3662,N_2610);
or U5529 (N_5529,N_3539,N_3239);
nand U5530 (N_5530,N_4633,N_3684);
nand U5531 (N_5531,N_3172,N_2662);
nor U5532 (N_5532,N_4734,N_2848);
or U5533 (N_5533,N_3872,N_2857);
or U5534 (N_5534,N_2543,N_4842);
and U5535 (N_5535,N_3323,N_3069);
nand U5536 (N_5536,N_3879,N_3525);
or U5537 (N_5537,N_4397,N_2795);
nand U5538 (N_5538,N_3858,N_3857);
or U5539 (N_5539,N_4224,N_4998);
and U5540 (N_5540,N_4766,N_4311);
nor U5541 (N_5541,N_2881,N_4037);
or U5542 (N_5542,N_3787,N_2936);
xor U5543 (N_5543,N_2862,N_4195);
and U5544 (N_5544,N_2940,N_4388);
or U5545 (N_5545,N_3547,N_2872);
or U5546 (N_5546,N_3793,N_2933);
nand U5547 (N_5547,N_4415,N_3873);
and U5548 (N_5548,N_4177,N_4865);
nor U5549 (N_5549,N_4565,N_3724);
nor U5550 (N_5550,N_4869,N_4489);
nor U5551 (N_5551,N_3362,N_2934);
and U5552 (N_5552,N_3425,N_2817);
nor U5553 (N_5553,N_4986,N_3277);
and U5554 (N_5554,N_4145,N_4996);
or U5555 (N_5555,N_3063,N_4682);
or U5556 (N_5556,N_2551,N_3740);
nor U5557 (N_5557,N_4498,N_4034);
nor U5558 (N_5558,N_3001,N_4957);
or U5559 (N_5559,N_2576,N_4596);
and U5560 (N_5560,N_2526,N_4365);
or U5561 (N_5561,N_4657,N_3997);
nor U5562 (N_5562,N_2930,N_2949);
and U5563 (N_5563,N_3030,N_3632);
nand U5564 (N_5564,N_4339,N_3090);
nand U5565 (N_5565,N_4093,N_4035);
or U5566 (N_5566,N_3191,N_4768);
and U5567 (N_5567,N_4659,N_2664);
nor U5568 (N_5568,N_4169,N_2508);
nor U5569 (N_5569,N_3541,N_3918);
or U5570 (N_5570,N_4822,N_4073);
nor U5571 (N_5571,N_3766,N_3502);
nand U5572 (N_5572,N_3656,N_3955);
nor U5573 (N_5573,N_3219,N_2502);
or U5574 (N_5574,N_3562,N_4070);
nand U5575 (N_5575,N_4026,N_4954);
nor U5576 (N_5576,N_4492,N_3479);
or U5577 (N_5577,N_2639,N_3471);
nor U5578 (N_5578,N_2871,N_3317);
nor U5579 (N_5579,N_4974,N_4226);
or U5580 (N_5580,N_3320,N_2976);
or U5581 (N_5581,N_4601,N_3633);
or U5582 (N_5582,N_4931,N_4105);
or U5583 (N_5583,N_2831,N_2667);
or U5584 (N_5584,N_4231,N_4252);
nor U5585 (N_5585,N_3968,N_4640);
or U5586 (N_5586,N_2766,N_3308);
nor U5587 (N_5587,N_4660,N_2510);
or U5588 (N_5588,N_4684,N_3772);
xnor U5589 (N_5589,N_3422,N_3203);
and U5590 (N_5590,N_3725,N_3053);
nor U5591 (N_5591,N_2840,N_4752);
nand U5592 (N_5592,N_4409,N_3930);
nand U5593 (N_5593,N_4030,N_3762);
nand U5594 (N_5594,N_3864,N_2815);
nand U5595 (N_5595,N_2803,N_4041);
xnor U5596 (N_5596,N_3472,N_3850);
and U5597 (N_5597,N_3970,N_4744);
nand U5598 (N_5598,N_3432,N_4207);
nand U5599 (N_5599,N_2660,N_2712);
nand U5600 (N_5600,N_4832,N_3266);
nand U5601 (N_5601,N_4531,N_2579);
or U5602 (N_5602,N_3690,N_3726);
or U5603 (N_5603,N_3844,N_3648);
and U5604 (N_5604,N_4164,N_4458);
and U5605 (N_5605,N_4098,N_3325);
and U5606 (N_5606,N_3823,N_3007);
or U5607 (N_5607,N_4829,N_3414);
and U5608 (N_5608,N_3763,N_2729);
nand U5609 (N_5609,N_2540,N_4624);
nor U5610 (N_5610,N_3754,N_4141);
nor U5611 (N_5611,N_3301,N_4787);
or U5612 (N_5612,N_4230,N_2942);
and U5613 (N_5613,N_3531,N_2585);
nor U5614 (N_5614,N_3964,N_4326);
nor U5615 (N_5615,N_4772,N_4966);
nand U5616 (N_5616,N_3391,N_3218);
nor U5617 (N_5617,N_4780,N_2554);
xor U5618 (N_5618,N_4451,N_2996);
or U5619 (N_5619,N_3402,N_4855);
or U5620 (N_5620,N_4434,N_4777);
and U5621 (N_5621,N_4723,N_4915);
nor U5622 (N_5622,N_4825,N_3509);
and U5623 (N_5623,N_3447,N_2614);
nand U5624 (N_5624,N_4368,N_4166);
nor U5625 (N_5625,N_2591,N_4578);
nor U5626 (N_5626,N_2725,N_4950);
and U5627 (N_5627,N_3883,N_4124);
nand U5628 (N_5628,N_4303,N_4205);
or U5629 (N_5629,N_3020,N_4370);
and U5630 (N_5630,N_3706,N_4603);
or U5631 (N_5631,N_4266,N_4991);
nor U5632 (N_5632,N_4040,N_3480);
or U5633 (N_5633,N_3429,N_4813);
nand U5634 (N_5634,N_4372,N_4004);
or U5635 (N_5635,N_4341,N_4620);
and U5636 (N_5636,N_3503,N_2602);
nor U5637 (N_5637,N_3694,N_2631);
nand U5638 (N_5638,N_4168,N_3413);
nand U5639 (N_5639,N_2740,N_4889);
nand U5640 (N_5640,N_3013,N_4011);
nor U5641 (N_5641,N_3321,N_3105);
nand U5642 (N_5642,N_3664,N_3119);
nor U5643 (N_5643,N_2640,N_3516);
and U5644 (N_5644,N_3905,N_2777);
or U5645 (N_5645,N_4259,N_3623);
nand U5646 (N_5646,N_4977,N_2595);
nor U5647 (N_5647,N_4495,N_4483);
nor U5648 (N_5648,N_4032,N_4891);
and U5649 (N_5649,N_3825,N_3834);
or U5650 (N_5650,N_4210,N_3985);
or U5651 (N_5651,N_4774,N_3939);
and U5652 (N_5652,N_3605,N_4562);
nor U5653 (N_5653,N_3177,N_3187);
and U5654 (N_5654,N_4852,N_2764);
nor U5655 (N_5655,N_4519,N_4894);
nor U5656 (N_5656,N_4591,N_2550);
nand U5657 (N_5657,N_3722,N_4724);
nand U5658 (N_5658,N_4513,N_4490);
or U5659 (N_5659,N_4469,N_3369);
or U5660 (N_5660,N_4538,N_4934);
nand U5661 (N_5661,N_3686,N_4214);
nand U5662 (N_5662,N_3009,N_3951);
and U5663 (N_5663,N_4481,N_4748);
or U5664 (N_5664,N_4514,N_2533);
or U5665 (N_5665,N_3146,N_4148);
and U5666 (N_5666,N_4745,N_4668);
or U5667 (N_5667,N_3186,N_4111);
nor U5668 (N_5668,N_4930,N_4689);
or U5669 (N_5669,N_3999,N_4125);
nor U5670 (N_5670,N_2560,N_4945);
and U5671 (N_5671,N_3635,N_3377);
nor U5672 (N_5672,N_3993,N_3033);
and U5673 (N_5673,N_2532,N_3281);
and U5674 (N_5674,N_2906,N_3666);
nand U5675 (N_5675,N_3800,N_2846);
or U5676 (N_5676,N_3871,N_3468);
nand U5677 (N_5677,N_4570,N_3596);
nand U5678 (N_5678,N_2733,N_3372);
or U5679 (N_5679,N_4783,N_3049);
or U5680 (N_5680,N_4702,N_3136);
and U5681 (N_5681,N_3324,N_4664);
nor U5682 (N_5682,N_4518,N_3178);
nand U5683 (N_5683,N_4758,N_3511);
and U5684 (N_5684,N_3451,N_4269);
nor U5685 (N_5685,N_4497,N_2827);
and U5686 (N_5686,N_4750,N_2598);
nand U5687 (N_5687,N_3797,N_4448);
and U5688 (N_5688,N_2959,N_4085);
or U5689 (N_5689,N_3587,N_3574);
nand U5690 (N_5690,N_4390,N_3168);
and U5691 (N_5691,N_3174,N_4550);
or U5692 (N_5692,N_2894,N_4179);
or U5693 (N_5693,N_3564,N_4690);
nor U5694 (N_5694,N_3515,N_3375);
nor U5695 (N_5695,N_3079,N_4383);
nand U5696 (N_5696,N_2570,N_3485);
or U5697 (N_5697,N_2622,N_3947);
or U5698 (N_5698,N_2541,N_3767);
nand U5699 (N_5699,N_4792,N_3477);
nor U5700 (N_5700,N_3796,N_3173);
or U5701 (N_5701,N_4128,N_3303);
and U5702 (N_5702,N_3745,N_4246);
and U5703 (N_5703,N_4705,N_4100);
and U5704 (N_5704,N_2727,N_3820);
and U5705 (N_5705,N_3933,N_4084);
or U5706 (N_5706,N_4990,N_4009);
or U5707 (N_5707,N_2971,N_3319);
and U5708 (N_5708,N_2612,N_2522);
and U5709 (N_5709,N_4134,N_3778);
and U5710 (N_5710,N_4063,N_3619);
xnor U5711 (N_5711,N_4949,N_4848);
and U5712 (N_5712,N_4308,N_3816);
nor U5713 (N_5713,N_3992,N_4658);
nor U5714 (N_5714,N_2753,N_3176);
nor U5715 (N_5715,N_4836,N_4062);
nor U5716 (N_5716,N_4270,N_4529);
or U5717 (N_5717,N_4992,N_3689);
xor U5718 (N_5718,N_4910,N_2678);
and U5719 (N_5719,N_3553,N_3011);
nor U5720 (N_5720,N_4074,N_4075);
xor U5721 (N_5721,N_4569,N_4457);
nand U5722 (N_5722,N_4963,N_3831);
nor U5723 (N_5723,N_3333,N_3244);
and U5724 (N_5724,N_3765,N_3849);
nand U5725 (N_5725,N_4267,N_4281);
nor U5726 (N_5726,N_4015,N_2762);
or U5727 (N_5727,N_2581,N_4892);
nor U5728 (N_5728,N_2854,N_3040);
and U5729 (N_5729,N_2856,N_2980);
or U5730 (N_5730,N_3124,N_3644);
nor U5731 (N_5731,N_4138,N_4413);
nand U5732 (N_5732,N_2577,N_4732);
and U5733 (N_5733,N_3271,N_4201);
nand U5734 (N_5734,N_4218,N_4993);
or U5735 (N_5735,N_4131,N_3616);
nand U5736 (N_5736,N_4013,N_2586);
or U5737 (N_5737,N_4798,N_4819);
or U5738 (N_5738,N_3500,N_4568);
and U5739 (N_5739,N_3363,N_4512);
and U5740 (N_5740,N_3649,N_2968);
nor U5741 (N_5741,N_2515,N_2547);
nand U5742 (N_5742,N_4039,N_2935);
and U5743 (N_5743,N_4683,N_3715);
and U5744 (N_5744,N_3394,N_3189);
or U5745 (N_5745,N_2714,N_4104);
and U5746 (N_5746,N_3565,N_3987);
and U5747 (N_5747,N_4586,N_3193);
or U5748 (N_5748,N_4239,N_3302);
or U5749 (N_5749,N_2618,N_2520);
nor U5750 (N_5750,N_3501,N_3716);
and U5751 (N_5751,N_4360,N_2567);
nand U5752 (N_5752,N_3598,N_2913);
nor U5753 (N_5753,N_2633,N_4523);
nor U5754 (N_5754,N_3783,N_3990);
nand U5755 (N_5755,N_4600,N_4461);
nor U5756 (N_5756,N_3579,N_3835);
nor U5757 (N_5757,N_3331,N_4406);
and U5758 (N_5758,N_3376,N_4435);
or U5759 (N_5759,N_3602,N_3573);
nand U5760 (N_5760,N_2674,N_2511);
and U5761 (N_5761,N_2603,N_4152);
nand U5762 (N_5762,N_3255,N_4460);
nor U5763 (N_5763,N_4482,N_4843);
nor U5764 (N_5764,N_3600,N_2973);
and U5765 (N_5765,N_4325,N_4135);
nand U5766 (N_5766,N_4044,N_3016);
or U5767 (N_5767,N_4697,N_3886);
and U5768 (N_5768,N_4431,N_2742);
or U5769 (N_5769,N_4553,N_4359);
nand U5770 (N_5770,N_2919,N_4897);
or U5771 (N_5771,N_4319,N_4096);
nor U5772 (N_5772,N_4530,N_4710);
and U5773 (N_5773,N_4916,N_3904);
nor U5774 (N_5774,N_2928,N_3829);
nor U5775 (N_5775,N_2806,N_3892);
nand U5776 (N_5776,N_2634,N_4108);
xor U5777 (N_5777,N_2726,N_3076);
and U5778 (N_5778,N_4679,N_4864);
or U5779 (N_5779,N_3544,N_4691);
nor U5780 (N_5780,N_3473,N_3416);
nor U5781 (N_5781,N_3601,N_4395);
or U5782 (N_5782,N_3902,N_3764);
nor U5783 (N_5783,N_2625,N_4136);
nor U5784 (N_5784,N_3454,N_3702);
and U5785 (N_5785,N_3945,N_3267);
or U5786 (N_5786,N_3112,N_4436);
or U5787 (N_5787,N_4791,N_4348);
nand U5788 (N_5788,N_4987,N_4709);
or U5789 (N_5789,N_4666,N_3352);
or U5790 (N_5790,N_4795,N_3347);
and U5791 (N_5791,N_2531,N_4868);
and U5792 (N_5792,N_3667,N_3057);
and U5793 (N_5793,N_3828,N_3699);
nand U5794 (N_5794,N_4837,N_2801);
or U5795 (N_5795,N_4680,N_4884);
nand U5796 (N_5796,N_3974,N_4623);
nor U5797 (N_5797,N_3856,N_3641);
and U5798 (N_5798,N_3728,N_4676);
or U5799 (N_5799,N_3313,N_2503);
nand U5800 (N_5800,N_3297,N_2927);
and U5801 (N_5801,N_2826,N_3495);
nor U5802 (N_5802,N_2738,N_3360);
or U5803 (N_5803,N_4609,N_4731);
nand U5804 (N_5804,N_2883,N_3938);
nor U5805 (N_5805,N_4632,N_3481);
or U5806 (N_5806,N_2525,N_4782);
or U5807 (N_5807,N_4130,N_2623);
or U5808 (N_5808,N_3137,N_3739);
or U5809 (N_5809,N_2849,N_3888);
and U5810 (N_5810,N_3919,N_3378);
xnor U5811 (N_5811,N_3379,N_3350);
or U5812 (N_5812,N_3650,N_2807);
or U5813 (N_5813,N_3089,N_3129);
nor U5814 (N_5814,N_3676,N_3185);
nor U5815 (N_5815,N_2624,N_3749);
nor U5816 (N_5816,N_3586,N_3096);
or U5817 (N_5817,N_2923,N_4764);
nand U5818 (N_5818,N_4881,N_3050);
or U5819 (N_5819,N_4456,N_3086);
nand U5820 (N_5820,N_3460,N_2822);
and U5821 (N_5821,N_4219,N_2902);
xor U5822 (N_5822,N_4969,N_2982);
nor U5823 (N_5823,N_3290,N_3436);
or U5824 (N_5824,N_2818,N_2535);
nor U5825 (N_5825,N_3163,N_3123);
or U5826 (N_5826,N_3897,N_2873);
and U5827 (N_5827,N_4182,N_3748);
nand U5828 (N_5828,N_2994,N_2956);
and U5829 (N_5829,N_4558,N_2954);
xnor U5830 (N_5830,N_4675,N_3526);
or U5831 (N_5831,N_4708,N_3751);
xor U5832 (N_5832,N_4594,N_4430);
and U5833 (N_5833,N_4437,N_3085);
or U5834 (N_5834,N_4180,N_3707);
or U5835 (N_5835,N_3703,N_2528);
xnor U5836 (N_5836,N_2775,N_3811);
nor U5837 (N_5837,N_4421,N_3907);
or U5838 (N_5838,N_2636,N_3171);
nor U5839 (N_5839,N_3152,N_3335);
nor U5840 (N_5840,N_4933,N_3714);
xnor U5841 (N_5841,N_3609,N_3484);
nand U5842 (N_5842,N_2507,N_3914);
or U5843 (N_5843,N_3081,N_2686);
nand U5844 (N_5844,N_4833,N_3855);
nand U5845 (N_5845,N_4815,N_4575);
and U5846 (N_5846,N_3093,N_4466);
nand U5847 (N_5847,N_3221,N_4028);
nor U5848 (N_5848,N_3631,N_4243);
nand U5849 (N_5849,N_4438,N_3840);
nor U5850 (N_5850,N_4615,N_3507);
or U5851 (N_5851,N_3737,N_4251);
and U5852 (N_5852,N_4419,N_3368);
and U5853 (N_5853,N_2830,N_4638);
or U5854 (N_5854,N_2769,N_3837);
or U5855 (N_5855,N_4335,N_3901);
nor U5856 (N_5856,N_4788,N_3924);
xor U5857 (N_5857,N_2545,N_2663);
or U5858 (N_5858,N_3238,N_3663);
nand U5859 (N_5859,N_3912,N_4315);
and U5860 (N_5860,N_4155,N_2717);
and U5861 (N_5861,N_4796,N_4499);
nor U5862 (N_5862,N_4511,N_3474);
and U5863 (N_5863,N_3312,N_3654);
or U5864 (N_5864,N_3846,N_4754);
or U5865 (N_5865,N_3131,N_3790);
nor U5866 (N_5866,N_3264,N_3155);
nor U5867 (N_5867,N_4521,N_2617);
nand U5868 (N_5868,N_2955,N_2580);
nor U5869 (N_5869,N_4386,N_4154);
or U5870 (N_5870,N_2998,N_2953);
nor U5871 (N_5871,N_4650,N_3348);
and U5872 (N_5872,N_4472,N_3140);
nand U5873 (N_5873,N_3456,N_3134);
and U5874 (N_5874,N_3687,N_3720);
or U5875 (N_5875,N_4376,N_4199);
and U5876 (N_5876,N_2616,N_3960);
nand U5877 (N_5877,N_4838,N_3782);
nand U5878 (N_5878,N_4576,N_2752);
or U5879 (N_5879,N_3496,N_3524);
and U5880 (N_5880,N_4978,N_3294);
or U5881 (N_5881,N_4309,N_4965);
or U5882 (N_5882,N_3931,N_4605);
nand U5883 (N_5883,N_4655,N_4233);
nor U5884 (N_5884,N_3719,N_4057);
nand U5885 (N_5885,N_4208,N_3969);
and U5886 (N_5886,N_4677,N_3424);
nand U5887 (N_5887,N_2921,N_3382);
nor U5888 (N_5888,N_2748,N_4343);
nor U5889 (N_5889,N_4725,N_3529);
nand U5890 (N_5890,N_3295,N_3014);
or U5891 (N_5891,N_4471,N_3103);
nand U5892 (N_5892,N_4327,N_3848);
xnor U5893 (N_5893,N_4908,N_3961);
and U5894 (N_5894,N_4830,N_4823);
or U5895 (N_5895,N_4076,N_3450);
and U5896 (N_5896,N_3506,N_3734);
xnor U5897 (N_5897,N_3307,N_2991);
or U5898 (N_5898,N_2970,N_3946);
nand U5899 (N_5899,N_4762,N_3792);
or U5900 (N_5900,N_3433,N_3956);
nor U5901 (N_5901,N_4888,N_2889);
nand U5902 (N_5902,N_4373,N_4342);
nor U5903 (N_5903,N_2985,N_2891);
nor U5904 (N_5904,N_3607,N_4936);
or U5905 (N_5905,N_2975,N_3139);
nor U5906 (N_5906,N_3228,N_4217);
nand U5907 (N_5907,N_3419,N_4137);
or U5908 (N_5908,N_3594,N_4000);
nand U5909 (N_5909,N_2865,N_4672);
nor U5910 (N_5910,N_3989,N_3338);
nand U5911 (N_5911,N_3036,N_4403);
nand U5912 (N_5912,N_4029,N_2524);
or U5913 (N_5913,N_4323,N_4470);
nand U5914 (N_5914,N_3984,N_4054);
nand U5915 (N_5915,N_3812,N_3908);
nor U5916 (N_5916,N_2628,N_2700);
or U5917 (N_5917,N_2690,N_2583);
nor U5918 (N_5918,N_3817,N_3283);
or U5919 (N_5919,N_2552,N_2630);
nand U5920 (N_5920,N_2835,N_3444);
and U5921 (N_5921,N_3505,N_4719);
and U5922 (N_5922,N_4071,N_3028);
nand U5923 (N_5923,N_2549,N_2699);
and U5924 (N_5924,N_3518,N_2802);
nor U5925 (N_5925,N_3592,N_4501);
nor U5926 (N_5926,N_4532,N_4042);
nand U5927 (N_5927,N_3750,N_3899);
nand U5928 (N_5928,N_3108,N_3824);
or U5929 (N_5929,N_2604,N_2837);
nand U5930 (N_5930,N_4876,N_3558);
and U5931 (N_5931,N_4306,N_2957);
or U5932 (N_5932,N_3180,N_3801);
and U5933 (N_5933,N_4928,N_4334);
or U5934 (N_5934,N_4741,N_2836);
nor U5935 (N_5935,N_3730,N_4450);
xor U5936 (N_5936,N_2637,N_3160);
nor U5937 (N_5937,N_4186,N_4407);
and U5938 (N_5938,N_3630,N_3743);
nor U5939 (N_5939,N_3340,N_2557);
nand U5940 (N_5940,N_2805,N_3449);
nand U5941 (N_5941,N_2537,N_3463);
or U5942 (N_5942,N_2804,N_3615);
nand U5943 (N_5943,N_4293,N_3791);
or U5944 (N_5944,N_4917,N_3910);
or U5945 (N_5945,N_4839,N_3513);
nor U5946 (N_5946,N_3041,N_4670);
nand U5947 (N_5947,N_3922,N_2656);
nor U5948 (N_5948,N_4229,N_3851);
or U5949 (N_5949,N_3356,N_4056);
and U5950 (N_5950,N_2993,N_3799);
and U5951 (N_5951,N_3212,N_3940);
or U5952 (N_5952,N_2722,N_3591);
xnor U5953 (N_5953,N_2781,N_4440);
nand U5954 (N_5954,N_4477,N_4522);
and U5955 (N_5955,N_4654,N_4593);
and U5956 (N_5956,N_2644,N_4465);
or U5957 (N_5957,N_2834,N_4276);
or U5958 (N_5958,N_3620,N_3184);
nor U5959 (N_5959,N_3893,N_4493);
or U5960 (N_5960,N_3780,N_4607);
nor U5961 (N_5961,N_4853,N_2761);
nor U5962 (N_5962,N_4183,N_4981);
nand U5963 (N_5963,N_2608,N_3336);
or U5964 (N_5964,N_3334,N_2962);
and U5965 (N_5965,N_4938,N_4086);
or U5966 (N_5966,N_4844,N_3913);
or U5967 (N_5967,N_4337,N_4364);
nand U5968 (N_5968,N_3179,N_4153);
and U5969 (N_5969,N_3877,N_3975);
or U5970 (N_5970,N_4634,N_4171);
xnor U5971 (N_5971,N_4943,N_4455);
or U5972 (N_5972,N_3949,N_4982);
nor U5973 (N_5973,N_3577,N_4170);
nand U5974 (N_5974,N_4010,N_4278);
nor U5975 (N_5975,N_3280,N_4139);
and U5976 (N_5976,N_2853,N_4110);
or U5977 (N_5977,N_4681,N_2702);
or U5978 (N_5978,N_2651,N_3784);
nand U5979 (N_5979,N_4835,N_2736);
xor U5980 (N_5980,N_3225,N_4583);
nor U5981 (N_5981,N_2512,N_3881);
nor U5982 (N_5982,N_3392,N_2788);
or U5983 (N_5983,N_4274,N_3693);
nand U5984 (N_5984,N_3712,N_4411);
and U5985 (N_5985,N_4143,N_4285);
or U5986 (N_5986,N_3552,N_4860);
nor U5987 (N_5987,N_2685,N_4160);
nor U5988 (N_5988,N_3169,N_4674);
and U5989 (N_5989,N_3151,N_2765);
or U5990 (N_5990,N_3802,N_4273);
and U5991 (N_5991,N_2784,N_2593);
and U5992 (N_5992,N_4980,N_3094);
or U5993 (N_5993,N_3243,N_2506);
nor U5994 (N_5994,N_4476,N_3442);
nand U5995 (N_5995,N_2786,N_3113);
xnor U5996 (N_5996,N_4877,N_4106);
nor U5997 (N_5997,N_2888,N_4485);
or U5998 (N_5998,N_2534,N_3006);
or U5999 (N_5999,N_3230,N_3206);
nand U6000 (N_6000,N_3417,N_2907);
and U6001 (N_6001,N_3545,N_3653);
xor U6002 (N_6002,N_3603,N_4778);
nor U6003 (N_6003,N_4630,N_3082);
or U6004 (N_6004,N_3549,N_3815);
or U6005 (N_6005,N_2650,N_3240);
and U6006 (N_6006,N_3697,N_4911);
nand U6007 (N_6007,N_4263,N_4671);
or U6008 (N_6008,N_2898,N_2601);
or U6009 (N_6009,N_3925,N_3842);
nand U6010 (N_6010,N_2659,N_3954);
nor U6011 (N_6011,N_3047,N_3071);
nor U6012 (N_6012,N_3876,N_4088);
nand U6013 (N_6013,N_2697,N_3917);
and U6014 (N_6014,N_3779,N_2797);
nand U6015 (N_6015,N_3154,N_2734);
nor U6016 (N_6016,N_2821,N_4698);
and U6017 (N_6017,N_4976,N_4209);
nor U6018 (N_6018,N_3589,N_2584);
and U6019 (N_6019,N_2654,N_4101);
and U6020 (N_6020,N_4656,N_4644);
and U6021 (N_6021,N_4694,N_3794);
and U6022 (N_6022,N_3934,N_4402);
or U6023 (N_6023,N_2600,N_4156);
and U6024 (N_6024,N_3826,N_4968);
nor U6025 (N_6025,N_3852,N_3627);
nand U6026 (N_6026,N_3875,N_4861);
or U6027 (N_6027,N_3314,N_3470);
or U6028 (N_6028,N_4338,N_2641);
nor U6029 (N_6029,N_3538,N_2990);
nand U6030 (N_6030,N_2675,N_3580);
and U6031 (N_6031,N_3401,N_2870);
or U6032 (N_6032,N_4443,N_4328);
and U6033 (N_6033,N_3973,N_3246);
nand U6034 (N_6034,N_4280,N_2988);
nand U6035 (N_6035,N_3135,N_4937);
nand U6036 (N_6036,N_4113,N_4389);
nand U6037 (N_6037,N_3198,N_4447);
and U6038 (N_6038,N_4951,N_3651);
nand U6039 (N_6039,N_3774,N_3279);
nand U6040 (N_6040,N_2886,N_4244);
and U6041 (N_6041,N_4240,N_2796);
nor U6042 (N_6042,N_4626,N_4895);
nor U6043 (N_6043,N_4333,N_3445);
and U6044 (N_6044,N_3031,N_3965);
and U6045 (N_6045,N_3581,N_4064);
nand U6046 (N_6046,N_3959,N_3555);
and U6047 (N_6047,N_4349,N_3786);
nor U6048 (N_6048,N_3709,N_2825);
or U6049 (N_6049,N_3430,N_3982);
nand U6050 (N_6050,N_3610,N_2563);
nand U6051 (N_6051,N_4878,N_4184);
nand U6052 (N_6052,N_2548,N_3236);
nor U6053 (N_6053,N_2908,N_4286);
nand U6054 (N_6054,N_3311,N_4959);
nand U6055 (N_6055,N_3729,N_2694);
nor U6056 (N_6056,N_3994,N_3298);
and U6057 (N_6057,N_3213,N_4038);
nor U6058 (N_6058,N_4548,N_3874);
xnor U6059 (N_6059,N_4173,N_4441);
xor U6060 (N_6060,N_2501,N_2589);
nor U6061 (N_6061,N_4736,N_4036);
nand U6062 (N_6062,N_4870,N_4387);
and U6063 (N_6063,N_2755,N_3705);
and U6064 (N_6064,N_3958,N_3027);
and U6065 (N_6065,N_2885,N_4287);
or U6066 (N_6066,N_2741,N_4717);
and U6067 (N_6067,N_3068,N_2943);
nand U6068 (N_6068,N_4983,N_3966);
and U6069 (N_6069,N_2880,N_4172);
and U6070 (N_6070,N_2841,N_2696);
or U6071 (N_6071,N_4947,N_2844);
nor U6072 (N_6072,N_4433,N_4534);
or U6073 (N_6073,N_3257,N_3158);
nand U6074 (N_6074,N_3318,N_3304);
nand U6075 (N_6075,N_4366,N_4161);
and U6076 (N_6076,N_3095,N_3978);
xor U6077 (N_6077,N_4567,N_4291);
and U6078 (N_6078,N_2652,N_4479);
nand U6079 (N_6079,N_2895,N_2757);
nand U6080 (N_6080,N_4921,N_3209);
and U6081 (N_6081,N_4089,N_4260);
nand U6082 (N_6082,N_4557,N_2901);
and U6083 (N_6083,N_2706,N_3182);
nand U6084 (N_6084,N_4400,N_3370);
nor U6085 (N_6085,N_2597,N_3117);
or U6086 (N_6086,N_4923,N_4616);
nor U6087 (N_6087,N_4294,N_4418);
or U6088 (N_6088,N_2691,N_3202);
or U6089 (N_6089,N_2914,N_2592);
nor U6090 (N_6090,N_4886,N_3657);
nor U6091 (N_6091,N_4665,N_4541);
and U6092 (N_6092,N_4248,N_4405);
nor U6093 (N_6093,N_2771,N_4524);
or U6094 (N_6094,N_3868,N_2561);
and U6095 (N_6095,N_4537,N_4893);
nor U6096 (N_6096,N_3157,N_4157);
nor U6097 (N_6097,N_3309,N_2594);
nand U6098 (N_6098,N_3920,N_4336);
and U6099 (N_6099,N_2571,N_4185);
and U6100 (N_6100,N_4312,N_4747);
or U6101 (N_6101,N_3675,N_4579);
nor U6102 (N_6102,N_3788,N_4988);
or U6103 (N_6103,N_2731,N_3278);
or U6104 (N_6104,N_3025,N_2884);
or U6105 (N_6105,N_3775,N_3645);
nand U6106 (N_6106,N_3365,N_3753);
or U6107 (N_6107,N_2542,N_4726);
nor U6108 (N_6108,N_3200,N_4192);
nand U6109 (N_6109,N_4257,N_3249);
and U6110 (N_6110,N_4688,N_4449);
or U6111 (N_6111,N_2558,N_3060);
and U6112 (N_6112,N_4515,N_4920);
or U6113 (N_6113,N_3695,N_3803);
nor U6114 (N_6114,N_4045,N_3909);
nor U6115 (N_6115,N_3051,N_4050);
and U6116 (N_6116,N_2967,N_4351);
or U6117 (N_6117,N_4382,N_4468);
or U6118 (N_6118,N_4641,N_3062);
nor U6119 (N_6119,N_4903,N_2669);
nor U6120 (N_6120,N_4958,N_2861);
nand U6121 (N_6121,N_3599,N_3691);
or U6122 (N_6122,N_4474,N_4277);
nand U6123 (N_6123,N_4005,N_4761);
or U6124 (N_6124,N_4971,N_3491);
nand U6125 (N_6125,N_4642,N_3410);
and U6126 (N_6126,N_2839,N_3798);
and U6127 (N_6127,N_2911,N_4647);
and U6128 (N_6128,N_4081,N_4590);
or U6129 (N_6129,N_3434,N_4646);
nor U6130 (N_6130,N_4526,N_4840);
and U6131 (N_6131,N_2704,N_2816);
nor U6132 (N_6132,N_4875,N_2905);
and U6133 (N_6133,N_3853,N_3953);
nor U6134 (N_6134,N_3130,N_3718);
or U6135 (N_6135,N_2995,N_3492);
and U6136 (N_6136,N_3395,N_4223);
nor U6137 (N_6137,N_3550,N_2768);
nor U6138 (N_6138,N_3446,N_4163);
or U6139 (N_6139,N_3747,N_4107);
and U6140 (N_6140,N_2811,N_3125);
nor U6141 (N_6141,N_3458,N_4424);
and U6142 (N_6142,N_3669,N_3467);
and U6143 (N_6143,N_4090,N_3181);
nor U6144 (N_6144,N_4061,N_3300);
or U6145 (N_6145,N_4540,N_4730);
nand U6146 (N_6146,N_2999,N_3067);
nand U6147 (N_6147,N_4849,N_2776);
nand U6148 (N_6148,N_4354,N_3229);
and U6149 (N_6149,N_2711,N_3567);
nand U6150 (N_6150,N_2688,N_3342);
and U6151 (N_6151,N_4316,N_3097);
nor U6152 (N_6152,N_2539,N_4995);
nand U6153 (N_6153,N_3805,N_2878);
or U6154 (N_6154,N_2997,N_4814);
or U6155 (N_6155,N_3988,N_3224);
nor U6156 (N_6156,N_4332,N_4120);
and U6157 (N_6157,N_3622,N_2760);
nand U6158 (N_6158,N_3114,N_2708);
and U6159 (N_6159,N_3024,N_3621);
and U6160 (N_6160,N_2720,N_3237);
nand U6161 (N_6161,N_4345,N_2812);
nor U6162 (N_6162,N_3462,N_2813);
nand U6163 (N_6163,N_2572,N_3332);
nor U6164 (N_6164,N_3578,N_3935);
or U6165 (N_6165,N_4423,N_4776);
or U6166 (N_6166,N_4733,N_4643);
nand U6167 (N_6167,N_4779,N_4929);
nor U6168 (N_6168,N_4900,N_3660);
nor U6169 (N_6169,N_3658,N_3260);
and U6170 (N_6170,N_4859,N_4767);
nor U6171 (N_6171,N_3056,N_3643);
and U6172 (N_6172,N_2673,N_2983);
and U6173 (N_6173,N_3983,N_3624);
nand U6174 (N_6174,N_3195,N_2774);
nor U6175 (N_6175,N_3898,N_2917);
and U6176 (N_6176,N_3806,N_4781);
nand U6177 (N_6177,N_4904,N_4765);
nor U6178 (N_6178,N_3214,N_2684);
nand U6179 (N_6179,N_4621,N_3540);
and U6180 (N_6180,N_3923,N_4065);
or U6181 (N_6181,N_4247,N_4127);
and U6182 (N_6182,N_2635,N_4525);
and U6183 (N_6183,N_4422,N_3104);
or U6184 (N_6184,N_4979,N_3346);
nand U6185 (N_6185,N_3384,N_3196);
or U6186 (N_6186,N_4856,N_4850);
or U6187 (N_6187,N_3147,N_2682);
nor U6188 (N_6188,N_3101,N_3490);
and U6189 (N_6189,N_4703,N_4234);
or U6190 (N_6190,N_4984,N_2556);
and U6191 (N_6191,N_3884,N_3248);
nor U6192 (N_6192,N_3253,N_4854);
nor U6193 (N_6193,N_3717,N_3159);
or U6194 (N_6194,N_4043,N_4543);
nor U6195 (N_6195,N_3637,N_2783);
nor U6196 (N_6196,N_3091,N_3092);
and U6197 (N_6197,N_2695,N_4811);
nand U6198 (N_6198,N_4494,N_4771);
and U6199 (N_6199,N_4197,N_3677);
nor U6200 (N_6200,N_3777,N_4478);
nand U6201 (N_6201,N_3074,N_3448);
nor U6202 (N_6202,N_3403,N_3830);
and U6203 (N_6203,N_3234,N_2984);
nor U6204 (N_6204,N_4025,N_2575);
and U6205 (N_6205,N_3661,N_4158);
or U6206 (N_6206,N_4162,N_3903);
xor U6207 (N_6207,N_4488,N_2655);
nand U6208 (N_6208,N_2798,N_3241);
and U6209 (N_6209,N_3887,N_3927);
or U6210 (N_6210,N_4126,N_3618);
nor U6211 (N_6211,N_3617,N_3075);
or U6212 (N_6212,N_4542,N_4961);
and U6213 (N_6213,N_3727,N_4755);
or U6214 (N_6214,N_4599,N_4989);
or U6215 (N_6215,N_3247,N_3029);
nor U6216 (N_6216,N_3251,N_4909);
or U6217 (N_6217,N_3768,N_2946);
and U6218 (N_6218,N_4417,N_4914);
and U6219 (N_6219,N_2668,N_4284);
nand U6220 (N_6220,N_4546,N_3192);
or U6221 (N_6221,N_4956,N_4082);
nand U6222 (N_6222,N_4142,N_4072);
nand U6223 (N_6223,N_3733,N_4144);
or U6224 (N_6224,N_3639,N_2687);
nand U6225 (N_6225,N_2863,N_2721);
and U6226 (N_6226,N_4384,N_3533);
and U6227 (N_6227,N_3440,N_3437);
and U6228 (N_6228,N_3010,N_3197);
and U6229 (N_6229,N_3608,N_2527);
and U6230 (N_6230,N_4906,N_3461);
or U6231 (N_6231,N_4545,N_3411);
or U6232 (N_6232,N_3407,N_4362);
nor U6233 (N_6233,N_4824,N_2845);
and U6234 (N_6234,N_4905,N_3517);
nand U6235 (N_6235,N_3386,N_3054);
and U6236 (N_6236,N_4960,N_4369);
and U6237 (N_6237,N_2791,N_3398);
and U6238 (N_6238,N_3133,N_2832);
and U6239 (N_6239,N_2661,N_3048);
and U6240 (N_6240,N_4150,N_3943);
or U6241 (N_6241,N_4211,N_3489);
nor U6242 (N_6242,N_3426,N_2792);
and U6243 (N_6243,N_3337,N_2958);
xnor U6244 (N_6244,N_2646,N_3588);
nor U6245 (N_6245,N_3536,N_4847);
and U6246 (N_6246,N_2960,N_3911);
nand U6247 (N_6247,N_4785,N_3614);
nor U6248 (N_6248,N_4581,N_3046);
nand U6249 (N_6249,N_3668,N_2814);
nor U6250 (N_6250,N_4203,N_4430);
nor U6251 (N_6251,N_2905,N_3345);
nor U6252 (N_6252,N_4023,N_4526);
nor U6253 (N_6253,N_2918,N_4386);
or U6254 (N_6254,N_4506,N_4929);
and U6255 (N_6255,N_4975,N_4450);
nand U6256 (N_6256,N_3123,N_3792);
nand U6257 (N_6257,N_4226,N_3438);
nor U6258 (N_6258,N_4825,N_3952);
or U6259 (N_6259,N_3749,N_4038);
or U6260 (N_6260,N_4020,N_2525);
or U6261 (N_6261,N_4572,N_2560);
and U6262 (N_6262,N_2621,N_4121);
or U6263 (N_6263,N_4956,N_4288);
nor U6264 (N_6264,N_4983,N_3066);
or U6265 (N_6265,N_4726,N_4959);
or U6266 (N_6266,N_3884,N_3962);
nor U6267 (N_6267,N_3505,N_3693);
or U6268 (N_6268,N_4865,N_4744);
nand U6269 (N_6269,N_4901,N_3108);
or U6270 (N_6270,N_3519,N_2950);
and U6271 (N_6271,N_3931,N_3573);
and U6272 (N_6272,N_4727,N_4524);
xor U6273 (N_6273,N_4088,N_3125);
nand U6274 (N_6274,N_4508,N_4884);
and U6275 (N_6275,N_3299,N_4164);
and U6276 (N_6276,N_3057,N_4508);
nor U6277 (N_6277,N_4551,N_3535);
nand U6278 (N_6278,N_4200,N_3455);
or U6279 (N_6279,N_3219,N_4127);
and U6280 (N_6280,N_4482,N_3542);
nor U6281 (N_6281,N_4110,N_3714);
or U6282 (N_6282,N_3587,N_3278);
nor U6283 (N_6283,N_3921,N_4395);
or U6284 (N_6284,N_3875,N_2602);
nor U6285 (N_6285,N_2738,N_4182);
or U6286 (N_6286,N_3971,N_4363);
and U6287 (N_6287,N_4874,N_3402);
and U6288 (N_6288,N_4745,N_3171);
and U6289 (N_6289,N_4433,N_4359);
nand U6290 (N_6290,N_4282,N_3152);
nand U6291 (N_6291,N_3457,N_3114);
nor U6292 (N_6292,N_3826,N_3190);
nor U6293 (N_6293,N_4504,N_3227);
nor U6294 (N_6294,N_3609,N_4568);
or U6295 (N_6295,N_3556,N_4976);
or U6296 (N_6296,N_3774,N_3766);
or U6297 (N_6297,N_4755,N_4542);
nand U6298 (N_6298,N_4360,N_3501);
or U6299 (N_6299,N_3816,N_2514);
nor U6300 (N_6300,N_4561,N_4537);
nor U6301 (N_6301,N_3231,N_4391);
nor U6302 (N_6302,N_3707,N_2859);
xor U6303 (N_6303,N_3900,N_2591);
nand U6304 (N_6304,N_4236,N_2966);
nor U6305 (N_6305,N_2896,N_4978);
or U6306 (N_6306,N_4776,N_2534);
or U6307 (N_6307,N_3210,N_4339);
and U6308 (N_6308,N_2625,N_4525);
nand U6309 (N_6309,N_3698,N_4255);
nand U6310 (N_6310,N_4032,N_2844);
nor U6311 (N_6311,N_4833,N_4306);
or U6312 (N_6312,N_4815,N_3345);
nand U6313 (N_6313,N_2764,N_3378);
xnor U6314 (N_6314,N_3259,N_4063);
nand U6315 (N_6315,N_2760,N_3870);
nand U6316 (N_6316,N_3840,N_4967);
or U6317 (N_6317,N_4369,N_4585);
or U6318 (N_6318,N_3332,N_3598);
nor U6319 (N_6319,N_3576,N_4387);
nand U6320 (N_6320,N_2567,N_2726);
or U6321 (N_6321,N_3589,N_4089);
and U6322 (N_6322,N_2691,N_3862);
or U6323 (N_6323,N_3306,N_3810);
or U6324 (N_6324,N_2750,N_4117);
nand U6325 (N_6325,N_2999,N_2727);
and U6326 (N_6326,N_3847,N_4020);
nor U6327 (N_6327,N_3479,N_2582);
and U6328 (N_6328,N_3910,N_3246);
or U6329 (N_6329,N_4373,N_3811);
and U6330 (N_6330,N_2946,N_3158);
nand U6331 (N_6331,N_3062,N_2696);
or U6332 (N_6332,N_4898,N_3562);
nand U6333 (N_6333,N_4264,N_4954);
nand U6334 (N_6334,N_3619,N_4987);
nor U6335 (N_6335,N_2790,N_3100);
nand U6336 (N_6336,N_4149,N_3139);
nand U6337 (N_6337,N_4053,N_3443);
or U6338 (N_6338,N_4598,N_4580);
nor U6339 (N_6339,N_4993,N_4110);
and U6340 (N_6340,N_3980,N_4882);
and U6341 (N_6341,N_4665,N_4028);
nand U6342 (N_6342,N_2702,N_3877);
nand U6343 (N_6343,N_4993,N_3118);
nand U6344 (N_6344,N_2559,N_3505);
nor U6345 (N_6345,N_4801,N_3952);
or U6346 (N_6346,N_2694,N_4812);
nor U6347 (N_6347,N_3782,N_4043);
or U6348 (N_6348,N_4359,N_2635);
and U6349 (N_6349,N_2524,N_2648);
nand U6350 (N_6350,N_4166,N_4283);
and U6351 (N_6351,N_3277,N_3284);
nand U6352 (N_6352,N_2539,N_3766);
nor U6353 (N_6353,N_4041,N_4384);
nand U6354 (N_6354,N_2753,N_2684);
and U6355 (N_6355,N_2633,N_4219);
and U6356 (N_6356,N_2703,N_3454);
nand U6357 (N_6357,N_4577,N_2636);
or U6358 (N_6358,N_2657,N_4537);
and U6359 (N_6359,N_3216,N_3078);
or U6360 (N_6360,N_3668,N_2737);
and U6361 (N_6361,N_3753,N_4932);
xnor U6362 (N_6362,N_3129,N_4527);
or U6363 (N_6363,N_4765,N_4285);
nor U6364 (N_6364,N_4579,N_3966);
and U6365 (N_6365,N_3948,N_4729);
nand U6366 (N_6366,N_4404,N_2603);
and U6367 (N_6367,N_3420,N_4361);
nor U6368 (N_6368,N_2785,N_4392);
nor U6369 (N_6369,N_2772,N_4385);
and U6370 (N_6370,N_2957,N_4503);
nand U6371 (N_6371,N_2724,N_2897);
xnor U6372 (N_6372,N_2741,N_3712);
nand U6373 (N_6373,N_3175,N_3659);
nand U6374 (N_6374,N_3840,N_4614);
and U6375 (N_6375,N_2831,N_4530);
or U6376 (N_6376,N_2772,N_4541);
nor U6377 (N_6377,N_2879,N_4109);
nand U6378 (N_6378,N_3886,N_4195);
nand U6379 (N_6379,N_3557,N_3124);
or U6380 (N_6380,N_4397,N_3112);
nor U6381 (N_6381,N_4507,N_3768);
nand U6382 (N_6382,N_4041,N_4159);
nand U6383 (N_6383,N_4507,N_4985);
or U6384 (N_6384,N_4552,N_3632);
nor U6385 (N_6385,N_2539,N_3844);
nand U6386 (N_6386,N_3000,N_4804);
and U6387 (N_6387,N_2547,N_3129);
nand U6388 (N_6388,N_3155,N_4161);
or U6389 (N_6389,N_4355,N_2900);
nand U6390 (N_6390,N_3409,N_3125);
or U6391 (N_6391,N_3931,N_2696);
xor U6392 (N_6392,N_2904,N_3400);
and U6393 (N_6393,N_3332,N_4360);
xor U6394 (N_6394,N_3083,N_4527);
nor U6395 (N_6395,N_3713,N_3728);
and U6396 (N_6396,N_2513,N_4628);
or U6397 (N_6397,N_2598,N_3799);
or U6398 (N_6398,N_4652,N_2548);
or U6399 (N_6399,N_4236,N_4933);
or U6400 (N_6400,N_3696,N_3925);
nor U6401 (N_6401,N_2880,N_3267);
or U6402 (N_6402,N_4964,N_4101);
xnor U6403 (N_6403,N_2647,N_3562);
nand U6404 (N_6404,N_4834,N_2781);
or U6405 (N_6405,N_4100,N_3335);
and U6406 (N_6406,N_2756,N_2662);
nand U6407 (N_6407,N_3700,N_4292);
nand U6408 (N_6408,N_2575,N_4006);
and U6409 (N_6409,N_4832,N_2823);
nor U6410 (N_6410,N_4887,N_4481);
nor U6411 (N_6411,N_3338,N_3104);
and U6412 (N_6412,N_4223,N_4523);
nor U6413 (N_6413,N_3676,N_3075);
or U6414 (N_6414,N_3679,N_2849);
or U6415 (N_6415,N_3622,N_2873);
nand U6416 (N_6416,N_4445,N_3752);
nor U6417 (N_6417,N_3298,N_3356);
xnor U6418 (N_6418,N_4981,N_3109);
and U6419 (N_6419,N_3871,N_4804);
and U6420 (N_6420,N_2660,N_3142);
nand U6421 (N_6421,N_2811,N_2513);
xnor U6422 (N_6422,N_2915,N_3331);
nand U6423 (N_6423,N_3745,N_2664);
or U6424 (N_6424,N_3205,N_2673);
or U6425 (N_6425,N_4355,N_4900);
nor U6426 (N_6426,N_2635,N_3043);
nand U6427 (N_6427,N_4958,N_2929);
nor U6428 (N_6428,N_3243,N_4229);
nor U6429 (N_6429,N_4577,N_4970);
or U6430 (N_6430,N_3139,N_2817);
nor U6431 (N_6431,N_3438,N_2796);
and U6432 (N_6432,N_3555,N_3168);
or U6433 (N_6433,N_2788,N_3035);
and U6434 (N_6434,N_4445,N_4605);
nor U6435 (N_6435,N_2792,N_4621);
nand U6436 (N_6436,N_3072,N_2597);
xor U6437 (N_6437,N_4439,N_3884);
nand U6438 (N_6438,N_2501,N_3653);
nor U6439 (N_6439,N_2648,N_4255);
nand U6440 (N_6440,N_3322,N_3042);
nand U6441 (N_6441,N_4206,N_2912);
nor U6442 (N_6442,N_3784,N_3327);
xor U6443 (N_6443,N_3508,N_2966);
nor U6444 (N_6444,N_3240,N_3481);
or U6445 (N_6445,N_2970,N_3423);
or U6446 (N_6446,N_3920,N_4478);
or U6447 (N_6447,N_4236,N_4150);
nor U6448 (N_6448,N_3252,N_2675);
nand U6449 (N_6449,N_2780,N_3689);
and U6450 (N_6450,N_4721,N_3558);
and U6451 (N_6451,N_3896,N_4191);
nor U6452 (N_6452,N_4961,N_2837);
nand U6453 (N_6453,N_4456,N_4735);
nand U6454 (N_6454,N_2699,N_4247);
and U6455 (N_6455,N_2665,N_4296);
nand U6456 (N_6456,N_2637,N_4983);
or U6457 (N_6457,N_3645,N_2725);
nand U6458 (N_6458,N_4599,N_4791);
or U6459 (N_6459,N_2929,N_4004);
nand U6460 (N_6460,N_2520,N_3359);
and U6461 (N_6461,N_4499,N_4366);
nor U6462 (N_6462,N_3871,N_2890);
or U6463 (N_6463,N_3440,N_3376);
nand U6464 (N_6464,N_2690,N_4793);
nand U6465 (N_6465,N_4466,N_2981);
or U6466 (N_6466,N_3108,N_2819);
nand U6467 (N_6467,N_4814,N_3055);
and U6468 (N_6468,N_4623,N_2848);
and U6469 (N_6469,N_4407,N_3740);
nor U6470 (N_6470,N_3616,N_2694);
or U6471 (N_6471,N_4929,N_3402);
or U6472 (N_6472,N_4771,N_2848);
nor U6473 (N_6473,N_2900,N_4260);
nor U6474 (N_6474,N_4057,N_3907);
nor U6475 (N_6475,N_4403,N_3955);
and U6476 (N_6476,N_4903,N_2748);
or U6477 (N_6477,N_3271,N_4455);
nand U6478 (N_6478,N_4136,N_3539);
nor U6479 (N_6479,N_3380,N_4394);
and U6480 (N_6480,N_4242,N_4594);
nor U6481 (N_6481,N_3226,N_4420);
nand U6482 (N_6482,N_4816,N_4655);
nor U6483 (N_6483,N_4775,N_2558);
xnor U6484 (N_6484,N_4812,N_4259);
nand U6485 (N_6485,N_2672,N_4358);
or U6486 (N_6486,N_3960,N_4840);
nor U6487 (N_6487,N_3144,N_3340);
nand U6488 (N_6488,N_3451,N_2892);
and U6489 (N_6489,N_3080,N_4079);
nand U6490 (N_6490,N_3430,N_4297);
and U6491 (N_6491,N_4918,N_3594);
or U6492 (N_6492,N_4313,N_3683);
xor U6493 (N_6493,N_4289,N_4372);
or U6494 (N_6494,N_3430,N_3308);
and U6495 (N_6495,N_4809,N_2607);
and U6496 (N_6496,N_4074,N_4040);
or U6497 (N_6497,N_4992,N_2701);
nor U6498 (N_6498,N_3618,N_4326);
nand U6499 (N_6499,N_3135,N_3802);
nor U6500 (N_6500,N_3868,N_2526);
and U6501 (N_6501,N_4992,N_3421);
and U6502 (N_6502,N_4891,N_4284);
nand U6503 (N_6503,N_2739,N_3330);
nand U6504 (N_6504,N_3218,N_3146);
xor U6505 (N_6505,N_4031,N_3806);
or U6506 (N_6506,N_4457,N_4775);
and U6507 (N_6507,N_4254,N_3199);
nor U6508 (N_6508,N_2587,N_4436);
or U6509 (N_6509,N_2784,N_4272);
or U6510 (N_6510,N_4790,N_2944);
or U6511 (N_6511,N_3568,N_4008);
nand U6512 (N_6512,N_3768,N_3044);
or U6513 (N_6513,N_3759,N_3454);
nor U6514 (N_6514,N_4474,N_2780);
nand U6515 (N_6515,N_2525,N_3717);
nand U6516 (N_6516,N_3908,N_3167);
and U6517 (N_6517,N_3701,N_4673);
and U6518 (N_6518,N_3217,N_4002);
nor U6519 (N_6519,N_3700,N_3901);
nor U6520 (N_6520,N_4033,N_4304);
nand U6521 (N_6521,N_4859,N_4502);
and U6522 (N_6522,N_2879,N_4979);
and U6523 (N_6523,N_4920,N_4092);
and U6524 (N_6524,N_2557,N_4228);
and U6525 (N_6525,N_4037,N_2844);
or U6526 (N_6526,N_2782,N_2647);
or U6527 (N_6527,N_3320,N_2907);
nand U6528 (N_6528,N_3058,N_3417);
nor U6529 (N_6529,N_3901,N_2879);
or U6530 (N_6530,N_3560,N_3365);
nand U6531 (N_6531,N_2684,N_4178);
nand U6532 (N_6532,N_2702,N_3346);
and U6533 (N_6533,N_3078,N_4320);
and U6534 (N_6534,N_3581,N_4440);
and U6535 (N_6535,N_2521,N_3745);
or U6536 (N_6536,N_4253,N_4914);
and U6537 (N_6537,N_3143,N_4467);
nor U6538 (N_6538,N_4406,N_3800);
or U6539 (N_6539,N_3387,N_3267);
nor U6540 (N_6540,N_3774,N_2509);
and U6541 (N_6541,N_2861,N_3252);
and U6542 (N_6542,N_4628,N_3995);
or U6543 (N_6543,N_4382,N_4637);
nand U6544 (N_6544,N_3174,N_3938);
nor U6545 (N_6545,N_2602,N_4563);
and U6546 (N_6546,N_3655,N_3076);
or U6547 (N_6547,N_3703,N_4075);
or U6548 (N_6548,N_3782,N_2671);
or U6549 (N_6549,N_3010,N_2976);
nor U6550 (N_6550,N_4798,N_4289);
nand U6551 (N_6551,N_3416,N_4731);
nor U6552 (N_6552,N_3970,N_3810);
and U6553 (N_6553,N_2564,N_3234);
nor U6554 (N_6554,N_4589,N_4535);
nor U6555 (N_6555,N_3612,N_3965);
nand U6556 (N_6556,N_4465,N_3576);
nand U6557 (N_6557,N_4139,N_3287);
nand U6558 (N_6558,N_4287,N_4078);
xnor U6559 (N_6559,N_4427,N_4581);
or U6560 (N_6560,N_4322,N_3247);
nor U6561 (N_6561,N_3332,N_3608);
nand U6562 (N_6562,N_4069,N_3178);
and U6563 (N_6563,N_3329,N_4225);
nor U6564 (N_6564,N_4069,N_3319);
or U6565 (N_6565,N_3392,N_3687);
xor U6566 (N_6566,N_4784,N_3805);
nor U6567 (N_6567,N_3931,N_3937);
or U6568 (N_6568,N_4961,N_2976);
or U6569 (N_6569,N_4528,N_2824);
nand U6570 (N_6570,N_3825,N_3656);
nand U6571 (N_6571,N_2746,N_4997);
and U6572 (N_6572,N_3689,N_4908);
nand U6573 (N_6573,N_2783,N_3277);
or U6574 (N_6574,N_3231,N_4733);
nor U6575 (N_6575,N_3134,N_3163);
or U6576 (N_6576,N_4339,N_3118);
xor U6577 (N_6577,N_4166,N_3300);
nor U6578 (N_6578,N_3017,N_3769);
or U6579 (N_6579,N_3804,N_3471);
nand U6580 (N_6580,N_3568,N_3819);
nor U6581 (N_6581,N_3451,N_4862);
and U6582 (N_6582,N_4913,N_3568);
nand U6583 (N_6583,N_4941,N_2544);
nand U6584 (N_6584,N_3991,N_3044);
nor U6585 (N_6585,N_3406,N_2797);
nand U6586 (N_6586,N_3233,N_4656);
or U6587 (N_6587,N_4332,N_3731);
nor U6588 (N_6588,N_4662,N_3606);
and U6589 (N_6589,N_2721,N_4644);
nand U6590 (N_6590,N_4326,N_3966);
nand U6591 (N_6591,N_4598,N_4468);
nor U6592 (N_6592,N_3508,N_4816);
or U6593 (N_6593,N_4143,N_3792);
nand U6594 (N_6594,N_3712,N_4799);
nand U6595 (N_6595,N_4372,N_3867);
nand U6596 (N_6596,N_4624,N_3990);
nor U6597 (N_6597,N_2759,N_3031);
nand U6598 (N_6598,N_4806,N_4018);
and U6599 (N_6599,N_3444,N_3440);
and U6600 (N_6600,N_4442,N_2664);
nand U6601 (N_6601,N_4950,N_3030);
nand U6602 (N_6602,N_4997,N_4907);
or U6603 (N_6603,N_3986,N_2528);
nand U6604 (N_6604,N_3845,N_3612);
and U6605 (N_6605,N_3891,N_4181);
and U6606 (N_6606,N_4652,N_4137);
and U6607 (N_6607,N_3896,N_4171);
nor U6608 (N_6608,N_3269,N_3709);
nand U6609 (N_6609,N_3880,N_3981);
or U6610 (N_6610,N_4888,N_3452);
nor U6611 (N_6611,N_2635,N_2884);
nand U6612 (N_6612,N_4789,N_4457);
nand U6613 (N_6613,N_3424,N_2931);
or U6614 (N_6614,N_4663,N_3905);
and U6615 (N_6615,N_2880,N_2861);
nor U6616 (N_6616,N_2521,N_3845);
or U6617 (N_6617,N_4107,N_3933);
nor U6618 (N_6618,N_4293,N_2568);
nand U6619 (N_6619,N_3339,N_3860);
and U6620 (N_6620,N_3196,N_3347);
nand U6621 (N_6621,N_3070,N_2640);
or U6622 (N_6622,N_2750,N_4804);
or U6623 (N_6623,N_3208,N_3125);
nor U6624 (N_6624,N_3418,N_2727);
nand U6625 (N_6625,N_3112,N_3070);
nand U6626 (N_6626,N_2926,N_3785);
and U6627 (N_6627,N_4989,N_3038);
nand U6628 (N_6628,N_4072,N_3416);
nand U6629 (N_6629,N_4006,N_2764);
nor U6630 (N_6630,N_4450,N_4358);
or U6631 (N_6631,N_4699,N_2753);
and U6632 (N_6632,N_3834,N_3305);
and U6633 (N_6633,N_3607,N_3622);
nor U6634 (N_6634,N_4285,N_4165);
nand U6635 (N_6635,N_4110,N_4494);
nor U6636 (N_6636,N_2876,N_3872);
and U6637 (N_6637,N_3974,N_4987);
nand U6638 (N_6638,N_4351,N_3735);
or U6639 (N_6639,N_3038,N_3589);
and U6640 (N_6640,N_4237,N_4710);
or U6641 (N_6641,N_4198,N_3699);
and U6642 (N_6642,N_3021,N_4455);
nor U6643 (N_6643,N_3769,N_2968);
nor U6644 (N_6644,N_3420,N_3762);
xnor U6645 (N_6645,N_2915,N_3805);
or U6646 (N_6646,N_4704,N_3473);
nand U6647 (N_6647,N_2668,N_3942);
or U6648 (N_6648,N_4778,N_4313);
nand U6649 (N_6649,N_3831,N_4509);
or U6650 (N_6650,N_4601,N_4287);
or U6651 (N_6651,N_3881,N_4257);
or U6652 (N_6652,N_3380,N_2840);
and U6653 (N_6653,N_4391,N_4710);
nand U6654 (N_6654,N_3564,N_3172);
or U6655 (N_6655,N_4101,N_4086);
nand U6656 (N_6656,N_4919,N_2847);
or U6657 (N_6657,N_4744,N_4916);
nand U6658 (N_6658,N_2584,N_3643);
and U6659 (N_6659,N_4841,N_3657);
nand U6660 (N_6660,N_2918,N_3840);
nand U6661 (N_6661,N_4392,N_2876);
nor U6662 (N_6662,N_4960,N_3709);
nor U6663 (N_6663,N_3822,N_3944);
nor U6664 (N_6664,N_2919,N_4002);
nand U6665 (N_6665,N_3236,N_3038);
nor U6666 (N_6666,N_4815,N_4888);
and U6667 (N_6667,N_4807,N_3575);
or U6668 (N_6668,N_2697,N_3306);
and U6669 (N_6669,N_2852,N_3444);
and U6670 (N_6670,N_4818,N_4170);
or U6671 (N_6671,N_3191,N_4166);
nor U6672 (N_6672,N_3646,N_3243);
or U6673 (N_6673,N_4650,N_3620);
xnor U6674 (N_6674,N_3560,N_2850);
nand U6675 (N_6675,N_3456,N_3750);
or U6676 (N_6676,N_2668,N_2770);
nand U6677 (N_6677,N_4524,N_4083);
or U6678 (N_6678,N_3819,N_3227);
and U6679 (N_6679,N_3122,N_4314);
and U6680 (N_6680,N_4883,N_4323);
nand U6681 (N_6681,N_2723,N_3692);
nand U6682 (N_6682,N_2510,N_4548);
or U6683 (N_6683,N_3174,N_3549);
nor U6684 (N_6684,N_3051,N_4406);
or U6685 (N_6685,N_4365,N_3337);
xor U6686 (N_6686,N_4587,N_4205);
or U6687 (N_6687,N_4469,N_3807);
nand U6688 (N_6688,N_3127,N_3941);
or U6689 (N_6689,N_3517,N_4983);
nand U6690 (N_6690,N_2518,N_4100);
or U6691 (N_6691,N_3276,N_4994);
xnor U6692 (N_6692,N_3765,N_3745);
or U6693 (N_6693,N_4621,N_2862);
or U6694 (N_6694,N_3893,N_2985);
and U6695 (N_6695,N_3774,N_3680);
nor U6696 (N_6696,N_3038,N_4232);
nor U6697 (N_6697,N_4856,N_4517);
nand U6698 (N_6698,N_4701,N_2668);
nand U6699 (N_6699,N_3949,N_3082);
nand U6700 (N_6700,N_4489,N_4230);
or U6701 (N_6701,N_2967,N_2811);
nand U6702 (N_6702,N_4757,N_3619);
nand U6703 (N_6703,N_4474,N_4229);
nor U6704 (N_6704,N_4207,N_3986);
nand U6705 (N_6705,N_4784,N_3724);
and U6706 (N_6706,N_3101,N_2929);
xnor U6707 (N_6707,N_3921,N_3911);
nand U6708 (N_6708,N_3964,N_3247);
nand U6709 (N_6709,N_3271,N_3897);
or U6710 (N_6710,N_2974,N_3009);
and U6711 (N_6711,N_2850,N_3170);
and U6712 (N_6712,N_3883,N_3285);
nand U6713 (N_6713,N_4504,N_3710);
and U6714 (N_6714,N_3957,N_3856);
nand U6715 (N_6715,N_4722,N_4806);
nand U6716 (N_6716,N_4933,N_2903);
or U6717 (N_6717,N_2858,N_3573);
nand U6718 (N_6718,N_3855,N_2617);
nand U6719 (N_6719,N_4912,N_2918);
nor U6720 (N_6720,N_2919,N_4873);
xor U6721 (N_6721,N_2743,N_3984);
or U6722 (N_6722,N_2590,N_3726);
nor U6723 (N_6723,N_2954,N_4694);
or U6724 (N_6724,N_4126,N_3646);
or U6725 (N_6725,N_3762,N_3830);
or U6726 (N_6726,N_4528,N_3431);
xnor U6727 (N_6727,N_3722,N_3682);
xnor U6728 (N_6728,N_2693,N_3279);
nor U6729 (N_6729,N_4489,N_4558);
or U6730 (N_6730,N_4190,N_3600);
and U6731 (N_6731,N_3334,N_4006);
and U6732 (N_6732,N_4030,N_4559);
nand U6733 (N_6733,N_4027,N_3199);
nor U6734 (N_6734,N_4489,N_4353);
nor U6735 (N_6735,N_4044,N_3241);
nor U6736 (N_6736,N_2579,N_4436);
and U6737 (N_6737,N_3182,N_4844);
or U6738 (N_6738,N_4012,N_3447);
or U6739 (N_6739,N_3511,N_4245);
or U6740 (N_6740,N_4625,N_2917);
nor U6741 (N_6741,N_3848,N_3066);
xnor U6742 (N_6742,N_4720,N_4327);
nand U6743 (N_6743,N_2921,N_4894);
nor U6744 (N_6744,N_3450,N_3329);
or U6745 (N_6745,N_3818,N_2931);
and U6746 (N_6746,N_4101,N_3188);
nand U6747 (N_6747,N_3684,N_4414);
and U6748 (N_6748,N_4506,N_3598);
and U6749 (N_6749,N_2651,N_3942);
nand U6750 (N_6750,N_3893,N_4498);
nor U6751 (N_6751,N_4155,N_4513);
nor U6752 (N_6752,N_4712,N_4121);
nand U6753 (N_6753,N_3577,N_2514);
or U6754 (N_6754,N_4486,N_4818);
nor U6755 (N_6755,N_2863,N_2517);
and U6756 (N_6756,N_4185,N_3807);
or U6757 (N_6757,N_3488,N_2745);
and U6758 (N_6758,N_4218,N_3054);
and U6759 (N_6759,N_3489,N_3801);
and U6760 (N_6760,N_3588,N_3625);
nand U6761 (N_6761,N_3537,N_3955);
and U6762 (N_6762,N_3469,N_4323);
nor U6763 (N_6763,N_4023,N_4509);
and U6764 (N_6764,N_3081,N_3402);
nor U6765 (N_6765,N_3901,N_3935);
or U6766 (N_6766,N_2908,N_2525);
and U6767 (N_6767,N_4697,N_3921);
nand U6768 (N_6768,N_4754,N_2779);
or U6769 (N_6769,N_3278,N_4932);
nand U6770 (N_6770,N_2564,N_3765);
nand U6771 (N_6771,N_3110,N_4111);
or U6772 (N_6772,N_4032,N_2821);
nor U6773 (N_6773,N_3989,N_3744);
nor U6774 (N_6774,N_3162,N_4039);
or U6775 (N_6775,N_3782,N_2780);
and U6776 (N_6776,N_4072,N_4928);
or U6777 (N_6777,N_4816,N_4600);
and U6778 (N_6778,N_3699,N_4202);
nor U6779 (N_6779,N_2831,N_3405);
nor U6780 (N_6780,N_4641,N_4007);
or U6781 (N_6781,N_2651,N_2890);
or U6782 (N_6782,N_4577,N_4474);
nand U6783 (N_6783,N_4473,N_4938);
nor U6784 (N_6784,N_2776,N_2782);
or U6785 (N_6785,N_4062,N_4549);
nand U6786 (N_6786,N_4709,N_3572);
or U6787 (N_6787,N_4771,N_3258);
and U6788 (N_6788,N_2593,N_3237);
nand U6789 (N_6789,N_2921,N_4055);
or U6790 (N_6790,N_3320,N_3855);
and U6791 (N_6791,N_4380,N_4362);
nor U6792 (N_6792,N_4063,N_3272);
nand U6793 (N_6793,N_2500,N_2841);
nor U6794 (N_6794,N_4976,N_3677);
and U6795 (N_6795,N_3137,N_2780);
nand U6796 (N_6796,N_2836,N_3369);
and U6797 (N_6797,N_3968,N_3901);
or U6798 (N_6798,N_4895,N_2796);
xnor U6799 (N_6799,N_3085,N_4084);
xor U6800 (N_6800,N_4072,N_4426);
nor U6801 (N_6801,N_2856,N_3925);
or U6802 (N_6802,N_4670,N_4727);
xnor U6803 (N_6803,N_3050,N_4828);
nor U6804 (N_6804,N_3555,N_3518);
nand U6805 (N_6805,N_3370,N_3493);
or U6806 (N_6806,N_3895,N_2724);
nor U6807 (N_6807,N_4138,N_4862);
nor U6808 (N_6808,N_3423,N_3085);
nor U6809 (N_6809,N_4518,N_4782);
nor U6810 (N_6810,N_3878,N_3792);
nand U6811 (N_6811,N_3216,N_3949);
or U6812 (N_6812,N_4257,N_2517);
and U6813 (N_6813,N_3387,N_2605);
and U6814 (N_6814,N_2798,N_3443);
nor U6815 (N_6815,N_3338,N_4661);
and U6816 (N_6816,N_2643,N_4771);
or U6817 (N_6817,N_4100,N_3537);
or U6818 (N_6818,N_4092,N_3637);
or U6819 (N_6819,N_4293,N_2644);
and U6820 (N_6820,N_4076,N_4323);
xor U6821 (N_6821,N_3879,N_4351);
nor U6822 (N_6822,N_3268,N_2705);
nor U6823 (N_6823,N_4550,N_3153);
or U6824 (N_6824,N_4433,N_3417);
nand U6825 (N_6825,N_4488,N_2518);
nand U6826 (N_6826,N_4934,N_4499);
and U6827 (N_6827,N_4341,N_4959);
and U6828 (N_6828,N_2853,N_3167);
and U6829 (N_6829,N_3535,N_4579);
and U6830 (N_6830,N_2906,N_4244);
nor U6831 (N_6831,N_4366,N_4467);
nand U6832 (N_6832,N_3773,N_3808);
or U6833 (N_6833,N_4267,N_4673);
nor U6834 (N_6834,N_4535,N_4775);
nand U6835 (N_6835,N_3767,N_4609);
nand U6836 (N_6836,N_4691,N_4113);
nand U6837 (N_6837,N_2756,N_3029);
nand U6838 (N_6838,N_4046,N_3416);
nor U6839 (N_6839,N_3675,N_4004);
or U6840 (N_6840,N_4079,N_4989);
nor U6841 (N_6841,N_4263,N_4662);
nand U6842 (N_6842,N_4427,N_4453);
nor U6843 (N_6843,N_3345,N_3118);
nor U6844 (N_6844,N_3480,N_2826);
or U6845 (N_6845,N_2802,N_4804);
or U6846 (N_6846,N_2615,N_3092);
and U6847 (N_6847,N_3947,N_3576);
nor U6848 (N_6848,N_4957,N_3252);
or U6849 (N_6849,N_4984,N_2697);
and U6850 (N_6850,N_4596,N_4540);
and U6851 (N_6851,N_3705,N_3700);
nand U6852 (N_6852,N_4884,N_3914);
or U6853 (N_6853,N_4749,N_2881);
and U6854 (N_6854,N_2630,N_2860);
nand U6855 (N_6855,N_3370,N_4271);
nor U6856 (N_6856,N_3838,N_2810);
nand U6857 (N_6857,N_3990,N_2941);
nand U6858 (N_6858,N_3045,N_4040);
or U6859 (N_6859,N_4193,N_4832);
and U6860 (N_6860,N_3975,N_3038);
or U6861 (N_6861,N_4037,N_3288);
nand U6862 (N_6862,N_4925,N_2640);
nand U6863 (N_6863,N_4816,N_3137);
nand U6864 (N_6864,N_4659,N_3325);
or U6865 (N_6865,N_2597,N_4006);
nand U6866 (N_6866,N_4003,N_4498);
nand U6867 (N_6867,N_4911,N_3731);
and U6868 (N_6868,N_3598,N_3993);
or U6869 (N_6869,N_3710,N_4403);
or U6870 (N_6870,N_4728,N_3094);
or U6871 (N_6871,N_4858,N_4354);
nand U6872 (N_6872,N_2644,N_3386);
and U6873 (N_6873,N_4768,N_4549);
and U6874 (N_6874,N_4735,N_4622);
or U6875 (N_6875,N_4367,N_2847);
or U6876 (N_6876,N_2603,N_2652);
nor U6877 (N_6877,N_3918,N_3727);
and U6878 (N_6878,N_4095,N_3594);
nor U6879 (N_6879,N_2675,N_3231);
and U6880 (N_6880,N_4342,N_4672);
nand U6881 (N_6881,N_2649,N_3299);
and U6882 (N_6882,N_4374,N_2777);
nor U6883 (N_6883,N_2661,N_3275);
nor U6884 (N_6884,N_3591,N_4401);
or U6885 (N_6885,N_4499,N_2507);
and U6886 (N_6886,N_3756,N_3778);
nand U6887 (N_6887,N_3558,N_3711);
and U6888 (N_6888,N_2987,N_4008);
nand U6889 (N_6889,N_3621,N_3560);
or U6890 (N_6890,N_3538,N_4501);
nor U6891 (N_6891,N_4389,N_4031);
or U6892 (N_6892,N_4644,N_2754);
nand U6893 (N_6893,N_2792,N_3351);
and U6894 (N_6894,N_4441,N_3868);
nand U6895 (N_6895,N_4423,N_4845);
nand U6896 (N_6896,N_3712,N_4713);
nor U6897 (N_6897,N_4563,N_3136);
or U6898 (N_6898,N_4304,N_4413);
xnor U6899 (N_6899,N_3877,N_2507);
nand U6900 (N_6900,N_3818,N_2915);
nor U6901 (N_6901,N_2842,N_2655);
nor U6902 (N_6902,N_4906,N_3625);
nand U6903 (N_6903,N_3222,N_4539);
nor U6904 (N_6904,N_2594,N_4537);
or U6905 (N_6905,N_3046,N_3267);
nor U6906 (N_6906,N_2922,N_4673);
and U6907 (N_6907,N_4095,N_4474);
nand U6908 (N_6908,N_4587,N_3815);
and U6909 (N_6909,N_4367,N_3192);
or U6910 (N_6910,N_2540,N_2752);
and U6911 (N_6911,N_4802,N_4575);
nand U6912 (N_6912,N_3613,N_4345);
nand U6913 (N_6913,N_4800,N_3815);
nand U6914 (N_6914,N_4008,N_4490);
and U6915 (N_6915,N_2574,N_3521);
nor U6916 (N_6916,N_4588,N_3551);
or U6917 (N_6917,N_4323,N_3960);
nand U6918 (N_6918,N_3205,N_4893);
and U6919 (N_6919,N_4266,N_4346);
or U6920 (N_6920,N_3790,N_3602);
nand U6921 (N_6921,N_4600,N_4755);
or U6922 (N_6922,N_4331,N_2872);
or U6923 (N_6923,N_3083,N_4926);
or U6924 (N_6924,N_2604,N_3829);
nor U6925 (N_6925,N_3304,N_4738);
nand U6926 (N_6926,N_3590,N_4168);
nand U6927 (N_6927,N_2570,N_4435);
nor U6928 (N_6928,N_3202,N_3474);
or U6929 (N_6929,N_4228,N_2539);
and U6930 (N_6930,N_4926,N_4855);
nor U6931 (N_6931,N_4624,N_3370);
and U6932 (N_6932,N_4269,N_3896);
or U6933 (N_6933,N_4609,N_4498);
nor U6934 (N_6934,N_4334,N_3604);
and U6935 (N_6935,N_3981,N_2803);
nand U6936 (N_6936,N_2686,N_4967);
nor U6937 (N_6937,N_3100,N_3346);
or U6938 (N_6938,N_3696,N_4501);
or U6939 (N_6939,N_4873,N_2532);
and U6940 (N_6940,N_3252,N_2785);
nor U6941 (N_6941,N_4646,N_3989);
xnor U6942 (N_6942,N_4617,N_4831);
nand U6943 (N_6943,N_3196,N_3336);
nor U6944 (N_6944,N_4890,N_4812);
or U6945 (N_6945,N_4119,N_3317);
nor U6946 (N_6946,N_3269,N_2650);
nor U6947 (N_6947,N_3802,N_4021);
and U6948 (N_6948,N_2674,N_3326);
and U6949 (N_6949,N_2618,N_2926);
or U6950 (N_6950,N_2622,N_4072);
or U6951 (N_6951,N_3822,N_2998);
and U6952 (N_6952,N_2756,N_4643);
and U6953 (N_6953,N_3343,N_4790);
or U6954 (N_6954,N_3256,N_2918);
nor U6955 (N_6955,N_2846,N_4907);
nand U6956 (N_6956,N_3453,N_4154);
and U6957 (N_6957,N_4479,N_2614);
nor U6958 (N_6958,N_4177,N_3941);
or U6959 (N_6959,N_4724,N_3773);
or U6960 (N_6960,N_4102,N_2537);
nand U6961 (N_6961,N_3559,N_3202);
and U6962 (N_6962,N_4287,N_3307);
nand U6963 (N_6963,N_2565,N_4949);
and U6964 (N_6964,N_3468,N_2703);
nor U6965 (N_6965,N_4868,N_3166);
and U6966 (N_6966,N_4797,N_3328);
nand U6967 (N_6967,N_4221,N_2513);
nor U6968 (N_6968,N_4557,N_3814);
xor U6969 (N_6969,N_3078,N_3551);
or U6970 (N_6970,N_3674,N_3184);
and U6971 (N_6971,N_3401,N_4162);
and U6972 (N_6972,N_4800,N_4566);
and U6973 (N_6973,N_3004,N_4979);
nor U6974 (N_6974,N_4460,N_4324);
xor U6975 (N_6975,N_4928,N_2605);
or U6976 (N_6976,N_2978,N_2654);
nor U6977 (N_6977,N_4632,N_3395);
nand U6978 (N_6978,N_4516,N_3609);
or U6979 (N_6979,N_4384,N_4017);
and U6980 (N_6980,N_4460,N_3169);
and U6981 (N_6981,N_4962,N_4258);
nand U6982 (N_6982,N_4532,N_4642);
nand U6983 (N_6983,N_4575,N_3517);
or U6984 (N_6984,N_3098,N_3484);
xnor U6985 (N_6985,N_4422,N_3581);
and U6986 (N_6986,N_3952,N_4750);
or U6987 (N_6987,N_3750,N_4441);
and U6988 (N_6988,N_4967,N_4330);
and U6989 (N_6989,N_4676,N_3116);
and U6990 (N_6990,N_3404,N_2744);
nand U6991 (N_6991,N_3998,N_3702);
or U6992 (N_6992,N_3918,N_3531);
nor U6993 (N_6993,N_4333,N_2658);
nand U6994 (N_6994,N_4387,N_3893);
and U6995 (N_6995,N_4236,N_3625);
and U6996 (N_6996,N_4239,N_4023);
and U6997 (N_6997,N_4037,N_3000);
and U6998 (N_6998,N_2648,N_3574);
nand U6999 (N_6999,N_2749,N_3367);
nor U7000 (N_7000,N_3908,N_3632);
nor U7001 (N_7001,N_3442,N_3781);
nand U7002 (N_7002,N_2838,N_3188);
nand U7003 (N_7003,N_3593,N_3313);
and U7004 (N_7004,N_4923,N_4363);
and U7005 (N_7005,N_2824,N_2935);
or U7006 (N_7006,N_3007,N_2640);
nand U7007 (N_7007,N_4350,N_3942);
nor U7008 (N_7008,N_3984,N_2706);
xnor U7009 (N_7009,N_4338,N_3292);
or U7010 (N_7010,N_3142,N_3050);
or U7011 (N_7011,N_3381,N_3312);
nor U7012 (N_7012,N_4001,N_2653);
xor U7013 (N_7013,N_4988,N_2889);
and U7014 (N_7014,N_3978,N_4842);
nor U7015 (N_7015,N_2513,N_4297);
or U7016 (N_7016,N_3227,N_4957);
and U7017 (N_7017,N_2892,N_3775);
or U7018 (N_7018,N_3326,N_3724);
xor U7019 (N_7019,N_3865,N_2527);
and U7020 (N_7020,N_3781,N_3760);
nor U7021 (N_7021,N_2509,N_3949);
nand U7022 (N_7022,N_4857,N_3851);
and U7023 (N_7023,N_3307,N_2769);
and U7024 (N_7024,N_3625,N_4058);
nor U7025 (N_7025,N_3102,N_2829);
or U7026 (N_7026,N_4136,N_3800);
or U7027 (N_7027,N_3198,N_3555);
nor U7028 (N_7028,N_4346,N_2904);
and U7029 (N_7029,N_4719,N_4408);
or U7030 (N_7030,N_4417,N_4299);
nor U7031 (N_7031,N_2925,N_3836);
and U7032 (N_7032,N_2932,N_3486);
and U7033 (N_7033,N_3758,N_4274);
nor U7034 (N_7034,N_4114,N_2557);
nor U7035 (N_7035,N_4933,N_4213);
or U7036 (N_7036,N_3749,N_4465);
nand U7037 (N_7037,N_3463,N_3116);
or U7038 (N_7038,N_4339,N_2783);
and U7039 (N_7039,N_4945,N_3850);
or U7040 (N_7040,N_3075,N_4417);
xnor U7041 (N_7041,N_4345,N_3930);
nor U7042 (N_7042,N_4773,N_3520);
nor U7043 (N_7043,N_3554,N_4510);
nor U7044 (N_7044,N_4885,N_2844);
nor U7045 (N_7045,N_3273,N_4431);
or U7046 (N_7046,N_3416,N_3494);
nor U7047 (N_7047,N_3770,N_4373);
nand U7048 (N_7048,N_4912,N_3544);
and U7049 (N_7049,N_4474,N_4426);
nand U7050 (N_7050,N_3326,N_4539);
xnor U7051 (N_7051,N_2966,N_3562);
or U7052 (N_7052,N_3516,N_3553);
or U7053 (N_7053,N_2778,N_4652);
or U7054 (N_7054,N_4205,N_4882);
and U7055 (N_7055,N_3625,N_3350);
nor U7056 (N_7056,N_4389,N_3308);
and U7057 (N_7057,N_3796,N_3060);
nand U7058 (N_7058,N_3962,N_2736);
nand U7059 (N_7059,N_4922,N_4028);
or U7060 (N_7060,N_4171,N_4348);
nand U7061 (N_7061,N_4140,N_3490);
nor U7062 (N_7062,N_4205,N_3456);
nand U7063 (N_7063,N_4485,N_3506);
nor U7064 (N_7064,N_4461,N_3797);
xnor U7065 (N_7065,N_4908,N_2558);
nand U7066 (N_7066,N_2802,N_3472);
or U7067 (N_7067,N_4786,N_2940);
and U7068 (N_7068,N_2733,N_2578);
and U7069 (N_7069,N_4601,N_4980);
nor U7070 (N_7070,N_3525,N_2991);
or U7071 (N_7071,N_4083,N_3364);
and U7072 (N_7072,N_4227,N_4969);
nand U7073 (N_7073,N_2911,N_3029);
and U7074 (N_7074,N_3713,N_4554);
xnor U7075 (N_7075,N_3732,N_2989);
and U7076 (N_7076,N_4996,N_4027);
xor U7077 (N_7077,N_4910,N_4414);
or U7078 (N_7078,N_4335,N_4627);
nor U7079 (N_7079,N_3330,N_4285);
or U7080 (N_7080,N_3456,N_3021);
or U7081 (N_7081,N_3577,N_4496);
nor U7082 (N_7082,N_3013,N_3662);
nand U7083 (N_7083,N_4449,N_3358);
nand U7084 (N_7084,N_4946,N_4620);
nor U7085 (N_7085,N_4301,N_3548);
or U7086 (N_7086,N_4552,N_3009);
nor U7087 (N_7087,N_2917,N_3756);
nor U7088 (N_7088,N_3669,N_4844);
nand U7089 (N_7089,N_4675,N_4475);
or U7090 (N_7090,N_3440,N_2872);
nor U7091 (N_7091,N_4882,N_4022);
xor U7092 (N_7092,N_3008,N_4598);
and U7093 (N_7093,N_4718,N_3011);
nor U7094 (N_7094,N_3384,N_4001);
and U7095 (N_7095,N_4875,N_3095);
nor U7096 (N_7096,N_3447,N_2984);
nand U7097 (N_7097,N_3180,N_3012);
nand U7098 (N_7098,N_3139,N_3421);
and U7099 (N_7099,N_4632,N_4717);
or U7100 (N_7100,N_2590,N_3288);
xnor U7101 (N_7101,N_3708,N_3620);
or U7102 (N_7102,N_3230,N_3158);
or U7103 (N_7103,N_2936,N_3789);
nor U7104 (N_7104,N_3115,N_2701);
nor U7105 (N_7105,N_4443,N_4275);
or U7106 (N_7106,N_2990,N_4999);
xnor U7107 (N_7107,N_2669,N_3865);
xnor U7108 (N_7108,N_3329,N_4879);
or U7109 (N_7109,N_2784,N_4456);
nor U7110 (N_7110,N_2726,N_4862);
nor U7111 (N_7111,N_4448,N_2514);
nand U7112 (N_7112,N_4783,N_2616);
nor U7113 (N_7113,N_3896,N_4928);
and U7114 (N_7114,N_2594,N_4873);
and U7115 (N_7115,N_4435,N_3753);
and U7116 (N_7116,N_2857,N_2962);
nor U7117 (N_7117,N_2725,N_3884);
nand U7118 (N_7118,N_3339,N_3910);
or U7119 (N_7119,N_2809,N_4466);
nor U7120 (N_7120,N_4360,N_4797);
and U7121 (N_7121,N_4352,N_2629);
and U7122 (N_7122,N_2546,N_4943);
or U7123 (N_7123,N_4733,N_3956);
nor U7124 (N_7124,N_4356,N_4926);
or U7125 (N_7125,N_3118,N_4810);
nand U7126 (N_7126,N_4604,N_4192);
and U7127 (N_7127,N_2762,N_4785);
and U7128 (N_7128,N_4123,N_4045);
nor U7129 (N_7129,N_3784,N_3772);
nor U7130 (N_7130,N_3697,N_4916);
nor U7131 (N_7131,N_3142,N_3028);
nand U7132 (N_7132,N_4111,N_2577);
and U7133 (N_7133,N_4305,N_3899);
nand U7134 (N_7134,N_2800,N_3721);
and U7135 (N_7135,N_3652,N_4849);
or U7136 (N_7136,N_2547,N_4226);
nand U7137 (N_7137,N_3535,N_3281);
and U7138 (N_7138,N_3603,N_4472);
and U7139 (N_7139,N_4368,N_2726);
and U7140 (N_7140,N_4180,N_3008);
or U7141 (N_7141,N_3271,N_4393);
nand U7142 (N_7142,N_2592,N_2751);
nor U7143 (N_7143,N_4832,N_3557);
or U7144 (N_7144,N_2879,N_3082);
and U7145 (N_7145,N_3035,N_4673);
nor U7146 (N_7146,N_4221,N_3910);
and U7147 (N_7147,N_4008,N_4412);
xor U7148 (N_7148,N_3243,N_4935);
nand U7149 (N_7149,N_3334,N_3390);
and U7150 (N_7150,N_4519,N_3693);
and U7151 (N_7151,N_3596,N_4521);
or U7152 (N_7152,N_4608,N_4347);
nand U7153 (N_7153,N_3883,N_3641);
nor U7154 (N_7154,N_3694,N_4882);
or U7155 (N_7155,N_2592,N_4912);
nand U7156 (N_7156,N_2551,N_4537);
or U7157 (N_7157,N_4151,N_3460);
and U7158 (N_7158,N_4043,N_4240);
nand U7159 (N_7159,N_4007,N_4947);
nand U7160 (N_7160,N_4632,N_2512);
and U7161 (N_7161,N_4091,N_4438);
nor U7162 (N_7162,N_3524,N_3193);
nor U7163 (N_7163,N_2588,N_3352);
xor U7164 (N_7164,N_4590,N_4632);
and U7165 (N_7165,N_4094,N_4504);
nor U7166 (N_7166,N_2615,N_3156);
nand U7167 (N_7167,N_4565,N_3625);
nand U7168 (N_7168,N_3819,N_4823);
nand U7169 (N_7169,N_4825,N_4341);
and U7170 (N_7170,N_3845,N_2560);
nand U7171 (N_7171,N_4843,N_3459);
nor U7172 (N_7172,N_4109,N_4872);
nand U7173 (N_7173,N_3553,N_3833);
nor U7174 (N_7174,N_2870,N_4451);
and U7175 (N_7175,N_3638,N_4580);
nand U7176 (N_7176,N_2917,N_2619);
and U7177 (N_7177,N_2504,N_3786);
nor U7178 (N_7178,N_4517,N_3791);
nor U7179 (N_7179,N_2587,N_3697);
nand U7180 (N_7180,N_2779,N_3546);
nand U7181 (N_7181,N_4753,N_4267);
nor U7182 (N_7182,N_2565,N_3778);
and U7183 (N_7183,N_4769,N_4281);
and U7184 (N_7184,N_4115,N_2533);
and U7185 (N_7185,N_3455,N_3219);
and U7186 (N_7186,N_4161,N_4004);
nand U7187 (N_7187,N_4604,N_4758);
nand U7188 (N_7188,N_3861,N_4257);
or U7189 (N_7189,N_2974,N_2621);
nor U7190 (N_7190,N_4483,N_3947);
and U7191 (N_7191,N_3741,N_4404);
nand U7192 (N_7192,N_4443,N_2523);
nor U7193 (N_7193,N_4639,N_2699);
and U7194 (N_7194,N_3607,N_3343);
nand U7195 (N_7195,N_2617,N_4703);
nor U7196 (N_7196,N_4086,N_2610);
nor U7197 (N_7197,N_3544,N_3780);
or U7198 (N_7198,N_2722,N_4879);
and U7199 (N_7199,N_3449,N_4184);
nor U7200 (N_7200,N_3440,N_4466);
and U7201 (N_7201,N_4967,N_4841);
or U7202 (N_7202,N_4817,N_3143);
or U7203 (N_7203,N_2748,N_3539);
or U7204 (N_7204,N_3025,N_4754);
nand U7205 (N_7205,N_3178,N_2637);
nor U7206 (N_7206,N_4346,N_3247);
nor U7207 (N_7207,N_2761,N_2860);
xnor U7208 (N_7208,N_3957,N_4884);
or U7209 (N_7209,N_4968,N_4020);
or U7210 (N_7210,N_3894,N_3606);
and U7211 (N_7211,N_4683,N_3724);
nor U7212 (N_7212,N_3953,N_3931);
nand U7213 (N_7213,N_4635,N_3180);
nor U7214 (N_7214,N_2833,N_3037);
xnor U7215 (N_7215,N_3684,N_3747);
or U7216 (N_7216,N_4725,N_4997);
or U7217 (N_7217,N_4009,N_3714);
or U7218 (N_7218,N_4240,N_3175);
or U7219 (N_7219,N_2508,N_3531);
or U7220 (N_7220,N_3873,N_3336);
or U7221 (N_7221,N_4505,N_4453);
nand U7222 (N_7222,N_2746,N_4323);
or U7223 (N_7223,N_2537,N_2673);
nor U7224 (N_7224,N_4035,N_4775);
nand U7225 (N_7225,N_4181,N_4401);
nor U7226 (N_7226,N_4078,N_4108);
and U7227 (N_7227,N_3038,N_3410);
nor U7228 (N_7228,N_4216,N_4538);
or U7229 (N_7229,N_3118,N_4510);
and U7230 (N_7230,N_3631,N_4295);
or U7231 (N_7231,N_3279,N_4702);
nor U7232 (N_7232,N_4785,N_3270);
nor U7233 (N_7233,N_3405,N_2629);
nand U7234 (N_7234,N_3972,N_4183);
and U7235 (N_7235,N_3013,N_3443);
or U7236 (N_7236,N_3937,N_4705);
nand U7237 (N_7237,N_4653,N_3843);
or U7238 (N_7238,N_3779,N_3305);
or U7239 (N_7239,N_4428,N_4829);
nor U7240 (N_7240,N_3620,N_3381);
nor U7241 (N_7241,N_4344,N_3968);
and U7242 (N_7242,N_2853,N_3289);
nor U7243 (N_7243,N_4000,N_4350);
and U7244 (N_7244,N_2670,N_4205);
and U7245 (N_7245,N_3917,N_3710);
nand U7246 (N_7246,N_3008,N_3206);
nand U7247 (N_7247,N_2981,N_3034);
and U7248 (N_7248,N_4478,N_3167);
nand U7249 (N_7249,N_3077,N_2753);
and U7250 (N_7250,N_3962,N_4859);
xor U7251 (N_7251,N_3941,N_4342);
nor U7252 (N_7252,N_4648,N_3951);
and U7253 (N_7253,N_4366,N_3090);
and U7254 (N_7254,N_3041,N_2856);
nand U7255 (N_7255,N_4819,N_4004);
and U7256 (N_7256,N_4056,N_4361);
nand U7257 (N_7257,N_3550,N_4445);
nand U7258 (N_7258,N_3291,N_4794);
and U7259 (N_7259,N_3366,N_2574);
and U7260 (N_7260,N_3007,N_4990);
nand U7261 (N_7261,N_2953,N_3217);
and U7262 (N_7262,N_3928,N_4711);
nor U7263 (N_7263,N_4586,N_2670);
nor U7264 (N_7264,N_3258,N_4677);
or U7265 (N_7265,N_2527,N_4767);
nand U7266 (N_7266,N_3712,N_3236);
or U7267 (N_7267,N_2714,N_3185);
nor U7268 (N_7268,N_4693,N_4979);
nand U7269 (N_7269,N_3819,N_3240);
and U7270 (N_7270,N_4883,N_2526);
or U7271 (N_7271,N_3962,N_4752);
xor U7272 (N_7272,N_3858,N_3168);
nor U7273 (N_7273,N_2568,N_3947);
nor U7274 (N_7274,N_4499,N_4275);
nor U7275 (N_7275,N_2554,N_2555);
or U7276 (N_7276,N_2841,N_4695);
nor U7277 (N_7277,N_4186,N_4712);
and U7278 (N_7278,N_2699,N_2526);
nand U7279 (N_7279,N_3837,N_2906);
and U7280 (N_7280,N_4930,N_2841);
and U7281 (N_7281,N_4579,N_3903);
nor U7282 (N_7282,N_4259,N_3303);
nor U7283 (N_7283,N_4933,N_3351);
nand U7284 (N_7284,N_4525,N_2533);
nor U7285 (N_7285,N_3986,N_3978);
and U7286 (N_7286,N_2787,N_2688);
and U7287 (N_7287,N_2748,N_4562);
xnor U7288 (N_7288,N_4488,N_2801);
or U7289 (N_7289,N_2916,N_3917);
nor U7290 (N_7290,N_4518,N_3186);
and U7291 (N_7291,N_3176,N_3784);
nand U7292 (N_7292,N_3854,N_4976);
and U7293 (N_7293,N_3995,N_2959);
or U7294 (N_7294,N_4981,N_3745);
or U7295 (N_7295,N_4699,N_3695);
nand U7296 (N_7296,N_3707,N_4635);
nand U7297 (N_7297,N_2718,N_4470);
nor U7298 (N_7298,N_3793,N_2907);
and U7299 (N_7299,N_4409,N_4065);
and U7300 (N_7300,N_2730,N_3743);
nor U7301 (N_7301,N_4774,N_4875);
and U7302 (N_7302,N_4046,N_3510);
and U7303 (N_7303,N_4646,N_4700);
and U7304 (N_7304,N_4907,N_4008);
or U7305 (N_7305,N_3320,N_3164);
nor U7306 (N_7306,N_3470,N_4054);
or U7307 (N_7307,N_4481,N_3557);
and U7308 (N_7308,N_2866,N_2509);
or U7309 (N_7309,N_3672,N_2651);
nand U7310 (N_7310,N_4205,N_3684);
nor U7311 (N_7311,N_4096,N_2948);
nand U7312 (N_7312,N_4718,N_4552);
or U7313 (N_7313,N_4455,N_3564);
and U7314 (N_7314,N_3594,N_3604);
nor U7315 (N_7315,N_3029,N_4245);
xor U7316 (N_7316,N_3924,N_3486);
and U7317 (N_7317,N_4281,N_4758);
nand U7318 (N_7318,N_3990,N_4967);
nor U7319 (N_7319,N_3456,N_2921);
or U7320 (N_7320,N_4941,N_2744);
nor U7321 (N_7321,N_3782,N_3140);
and U7322 (N_7322,N_4775,N_3836);
nor U7323 (N_7323,N_3255,N_2703);
nand U7324 (N_7324,N_3421,N_4930);
and U7325 (N_7325,N_2652,N_4612);
or U7326 (N_7326,N_4098,N_4477);
or U7327 (N_7327,N_4102,N_3066);
and U7328 (N_7328,N_3782,N_4628);
and U7329 (N_7329,N_4857,N_3026);
nor U7330 (N_7330,N_3624,N_4385);
nor U7331 (N_7331,N_2835,N_4006);
nor U7332 (N_7332,N_3913,N_4761);
or U7333 (N_7333,N_3742,N_2846);
nor U7334 (N_7334,N_4751,N_3559);
and U7335 (N_7335,N_4333,N_4632);
and U7336 (N_7336,N_4316,N_4888);
nor U7337 (N_7337,N_4657,N_2748);
nand U7338 (N_7338,N_2963,N_4192);
or U7339 (N_7339,N_4730,N_4981);
xnor U7340 (N_7340,N_2628,N_3332);
nor U7341 (N_7341,N_3528,N_3909);
or U7342 (N_7342,N_4250,N_4527);
nand U7343 (N_7343,N_3616,N_3250);
nand U7344 (N_7344,N_4828,N_4070);
or U7345 (N_7345,N_3843,N_2890);
and U7346 (N_7346,N_3996,N_3007);
nand U7347 (N_7347,N_3702,N_3347);
nor U7348 (N_7348,N_4685,N_3751);
or U7349 (N_7349,N_4704,N_3625);
nor U7350 (N_7350,N_4710,N_4106);
nor U7351 (N_7351,N_2586,N_4833);
and U7352 (N_7352,N_3012,N_4941);
nand U7353 (N_7353,N_3140,N_4287);
nand U7354 (N_7354,N_3820,N_2668);
nand U7355 (N_7355,N_4104,N_2670);
xor U7356 (N_7356,N_3546,N_3320);
and U7357 (N_7357,N_4606,N_4078);
or U7358 (N_7358,N_3992,N_4261);
and U7359 (N_7359,N_4339,N_4394);
or U7360 (N_7360,N_2570,N_3272);
or U7361 (N_7361,N_3254,N_3193);
xnor U7362 (N_7362,N_4812,N_2756);
nor U7363 (N_7363,N_4522,N_3090);
and U7364 (N_7364,N_4671,N_3675);
and U7365 (N_7365,N_4665,N_3327);
and U7366 (N_7366,N_4952,N_4049);
nor U7367 (N_7367,N_2958,N_3412);
and U7368 (N_7368,N_4888,N_4488);
or U7369 (N_7369,N_2674,N_2759);
nand U7370 (N_7370,N_4239,N_3082);
and U7371 (N_7371,N_3384,N_2828);
or U7372 (N_7372,N_3978,N_3247);
or U7373 (N_7373,N_4928,N_2708);
nand U7374 (N_7374,N_4544,N_3819);
nand U7375 (N_7375,N_4189,N_4377);
or U7376 (N_7376,N_4940,N_3705);
or U7377 (N_7377,N_2691,N_2554);
and U7378 (N_7378,N_3919,N_2657);
and U7379 (N_7379,N_4909,N_3654);
nand U7380 (N_7380,N_3736,N_4504);
nand U7381 (N_7381,N_3563,N_3855);
nand U7382 (N_7382,N_3976,N_3799);
nand U7383 (N_7383,N_2969,N_4976);
and U7384 (N_7384,N_3786,N_4377);
nand U7385 (N_7385,N_4643,N_3548);
nand U7386 (N_7386,N_3475,N_4728);
and U7387 (N_7387,N_3097,N_4808);
and U7388 (N_7388,N_4288,N_3857);
and U7389 (N_7389,N_3383,N_4597);
or U7390 (N_7390,N_2587,N_3224);
nor U7391 (N_7391,N_2575,N_3573);
nor U7392 (N_7392,N_3134,N_3525);
or U7393 (N_7393,N_4795,N_2957);
nor U7394 (N_7394,N_4536,N_3237);
and U7395 (N_7395,N_2553,N_3102);
nor U7396 (N_7396,N_3980,N_4577);
or U7397 (N_7397,N_3278,N_4493);
nor U7398 (N_7398,N_2542,N_3923);
and U7399 (N_7399,N_3283,N_3264);
nand U7400 (N_7400,N_3954,N_2735);
nor U7401 (N_7401,N_3364,N_2911);
and U7402 (N_7402,N_3989,N_4015);
nor U7403 (N_7403,N_4060,N_4528);
nand U7404 (N_7404,N_4126,N_3554);
or U7405 (N_7405,N_4084,N_3097);
nand U7406 (N_7406,N_2739,N_3433);
and U7407 (N_7407,N_3287,N_4891);
or U7408 (N_7408,N_2830,N_3315);
and U7409 (N_7409,N_3330,N_4721);
nand U7410 (N_7410,N_2566,N_4707);
and U7411 (N_7411,N_3807,N_3184);
nand U7412 (N_7412,N_2605,N_4211);
nor U7413 (N_7413,N_3178,N_3934);
nor U7414 (N_7414,N_4666,N_3567);
or U7415 (N_7415,N_3882,N_3030);
or U7416 (N_7416,N_3735,N_3810);
nand U7417 (N_7417,N_3397,N_3519);
and U7418 (N_7418,N_4665,N_4758);
nor U7419 (N_7419,N_4108,N_4974);
nand U7420 (N_7420,N_4378,N_3525);
or U7421 (N_7421,N_4652,N_4599);
and U7422 (N_7422,N_2782,N_3095);
nor U7423 (N_7423,N_3161,N_3650);
nor U7424 (N_7424,N_2951,N_3665);
and U7425 (N_7425,N_4424,N_4842);
nor U7426 (N_7426,N_3673,N_3017);
nor U7427 (N_7427,N_3814,N_2520);
nor U7428 (N_7428,N_4949,N_4427);
and U7429 (N_7429,N_3943,N_4042);
or U7430 (N_7430,N_3120,N_3745);
nand U7431 (N_7431,N_4581,N_2589);
and U7432 (N_7432,N_3481,N_3892);
nor U7433 (N_7433,N_2583,N_3398);
and U7434 (N_7434,N_3005,N_3981);
nand U7435 (N_7435,N_3411,N_4877);
nand U7436 (N_7436,N_2683,N_4240);
or U7437 (N_7437,N_4452,N_3023);
and U7438 (N_7438,N_4095,N_4604);
nor U7439 (N_7439,N_3468,N_3243);
nor U7440 (N_7440,N_3068,N_3747);
and U7441 (N_7441,N_3721,N_2868);
and U7442 (N_7442,N_3401,N_3406);
or U7443 (N_7443,N_3623,N_4995);
or U7444 (N_7444,N_4574,N_3609);
xor U7445 (N_7445,N_4318,N_3850);
or U7446 (N_7446,N_3768,N_4765);
nor U7447 (N_7447,N_4985,N_3108);
nor U7448 (N_7448,N_4030,N_3022);
nand U7449 (N_7449,N_4488,N_2609);
and U7450 (N_7450,N_2957,N_3650);
or U7451 (N_7451,N_4931,N_4690);
nor U7452 (N_7452,N_2693,N_4355);
or U7453 (N_7453,N_4283,N_3938);
or U7454 (N_7454,N_2911,N_3217);
nor U7455 (N_7455,N_2790,N_3459);
or U7456 (N_7456,N_3430,N_3635);
or U7457 (N_7457,N_3523,N_3078);
nor U7458 (N_7458,N_4342,N_2797);
and U7459 (N_7459,N_4913,N_3831);
nor U7460 (N_7460,N_4046,N_3190);
or U7461 (N_7461,N_4533,N_3349);
and U7462 (N_7462,N_3253,N_3604);
or U7463 (N_7463,N_4234,N_4413);
nor U7464 (N_7464,N_4964,N_3476);
nand U7465 (N_7465,N_3420,N_4247);
nor U7466 (N_7466,N_3833,N_3708);
or U7467 (N_7467,N_2831,N_3861);
or U7468 (N_7468,N_4691,N_3985);
nor U7469 (N_7469,N_3692,N_2931);
or U7470 (N_7470,N_4736,N_3250);
or U7471 (N_7471,N_4224,N_4389);
nand U7472 (N_7472,N_3298,N_3806);
nor U7473 (N_7473,N_4816,N_3254);
and U7474 (N_7474,N_3450,N_3727);
xor U7475 (N_7475,N_4678,N_4716);
nand U7476 (N_7476,N_3887,N_4435);
and U7477 (N_7477,N_2937,N_4189);
nor U7478 (N_7478,N_3275,N_3897);
nand U7479 (N_7479,N_3169,N_2512);
or U7480 (N_7480,N_3561,N_3929);
or U7481 (N_7481,N_3105,N_2693);
and U7482 (N_7482,N_3408,N_3929);
nor U7483 (N_7483,N_3253,N_4140);
xor U7484 (N_7484,N_4610,N_2614);
or U7485 (N_7485,N_2954,N_3961);
or U7486 (N_7486,N_4821,N_3835);
or U7487 (N_7487,N_4167,N_2976);
and U7488 (N_7488,N_3997,N_2662);
nor U7489 (N_7489,N_4559,N_4004);
nand U7490 (N_7490,N_3392,N_3804);
nor U7491 (N_7491,N_4830,N_3456);
nor U7492 (N_7492,N_3231,N_2702);
or U7493 (N_7493,N_3277,N_3533);
nor U7494 (N_7494,N_3151,N_4956);
nor U7495 (N_7495,N_3897,N_3065);
and U7496 (N_7496,N_3120,N_3806);
nor U7497 (N_7497,N_4676,N_2831);
and U7498 (N_7498,N_2630,N_2588);
or U7499 (N_7499,N_4821,N_4629);
nand U7500 (N_7500,N_5487,N_5693);
nand U7501 (N_7501,N_5203,N_6611);
nor U7502 (N_7502,N_5520,N_6499);
or U7503 (N_7503,N_5426,N_5638);
nor U7504 (N_7504,N_5287,N_5876);
nand U7505 (N_7505,N_7407,N_7422);
and U7506 (N_7506,N_6606,N_5022);
xnor U7507 (N_7507,N_6101,N_5476);
nor U7508 (N_7508,N_7111,N_5659);
or U7509 (N_7509,N_6698,N_5236);
and U7510 (N_7510,N_6182,N_5888);
or U7511 (N_7511,N_6954,N_6386);
nor U7512 (N_7512,N_5951,N_6543);
xnor U7513 (N_7513,N_7132,N_5217);
and U7514 (N_7514,N_6517,N_7210);
and U7515 (N_7515,N_6950,N_5967);
and U7516 (N_7516,N_6081,N_7247);
and U7517 (N_7517,N_5878,N_6258);
or U7518 (N_7518,N_5529,N_6332);
nand U7519 (N_7519,N_5899,N_5056);
and U7520 (N_7520,N_5050,N_5858);
or U7521 (N_7521,N_6043,N_5434);
and U7522 (N_7522,N_7203,N_5710);
nand U7523 (N_7523,N_6012,N_6335);
or U7524 (N_7524,N_6170,N_6888);
or U7525 (N_7525,N_6647,N_6524);
and U7526 (N_7526,N_5215,N_5936);
nand U7527 (N_7527,N_5684,N_5625);
and U7528 (N_7528,N_5871,N_6457);
and U7529 (N_7529,N_6481,N_5163);
nand U7530 (N_7530,N_7103,N_5782);
nor U7531 (N_7531,N_5692,N_5610);
nor U7532 (N_7532,N_6164,N_5963);
nor U7533 (N_7533,N_6917,N_6935);
and U7534 (N_7534,N_6575,N_5147);
or U7535 (N_7535,N_7094,N_6760);
nand U7536 (N_7536,N_7029,N_7163);
or U7537 (N_7537,N_5616,N_7200);
nor U7538 (N_7538,N_5517,N_5035);
nor U7539 (N_7539,N_5094,N_6480);
nor U7540 (N_7540,N_6713,N_5618);
or U7541 (N_7541,N_6069,N_7009);
nand U7542 (N_7542,N_5764,N_5802);
and U7543 (N_7543,N_6261,N_5869);
nor U7544 (N_7544,N_5142,N_6431);
nor U7545 (N_7545,N_5188,N_6951);
and U7546 (N_7546,N_6648,N_5703);
and U7547 (N_7547,N_5250,N_7388);
nand U7548 (N_7548,N_6465,N_7327);
or U7549 (N_7549,N_6024,N_5283);
and U7550 (N_7550,N_7320,N_7489);
nand U7551 (N_7551,N_6336,N_6135);
or U7552 (N_7552,N_7336,N_6508);
nor U7553 (N_7553,N_6856,N_7175);
nor U7554 (N_7554,N_5093,N_5536);
nor U7555 (N_7555,N_5401,N_5446);
or U7556 (N_7556,N_7410,N_6512);
nand U7557 (N_7557,N_7182,N_7346);
and U7558 (N_7558,N_7118,N_6551);
nor U7559 (N_7559,N_5687,N_5999);
xor U7560 (N_7560,N_6102,N_6692);
nand U7561 (N_7561,N_5443,N_5230);
and U7562 (N_7562,N_6781,N_5008);
nand U7563 (N_7563,N_6639,N_6836);
and U7564 (N_7564,N_6117,N_6263);
nand U7565 (N_7565,N_7147,N_7167);
nor U7566 (N_7566,N_7433,N_5809);
nand U7567 (N_7567,N_5467,N_6239);
or U7568 (N_7568,N_6688,N_6138);
and U7569 (N_7569,N_6425,N_7142);
nand U7570 (N_7570,N_6742,N_7217);
nand U7571 (N_7571,N_5512,N_7183);
nand U7572 (N_7572,N_5136,N_7380);
nand U7573 (N_7573,N_6221,N_5202);
nor U7574 (N_7574,N_5277,N_5767);
or U7575 (N_7575,N_5732,N_5130);
nand U7576 (N_7576,N_6734,N_6326);
and U7577 (N_7577,N_5053,N_5745);
nand U7578 (N_7578,N_5198,N_5168);
nand U7579 (N_7579,N_6708,N_6806);
or U7580 (N_7580,N_5375,N_6889);
or U7581 (N_7581,N_6721,N_6343);
nand U7582 (N_7582,N_6977,N_7364);
nor U7583 (N_7583,N_5281,N_5252);
nor U7584 (N_7584,N_5227,N_7330);
nor U7585 (N_7585,N_5909,N_6382);
nor U7586 (N_7586,N_6354,N_7243);
nand U7587 (N_7587,N_7076,N_7214);
nand U7588 (N_7588,N_6001,N_6016);
nand U7589 (N_7589,N_5741,N_6829);
or U7590 (N_7590,N_6469,N_5826);
xor U7591 (N_7591,N_5892,N_7257);
and U7592 (N_7592,N_6541,N_7098);
and U7593 (N_7593,N_6381,N_6372);
nand U7594 (N_7594,N_6034,N_5962);
nand U7595 (N_7595,N_7000,N_7493);
nor U7596 (N_7596,N_6274,N_6448);
xnor U7597 (N_7597,N_5643,N_6180);
or U7598 (N_7598,N_6696,N_7169);
and U7599 (N_7599,N_5814,N_7265);
nor U7600 (N_7600,N_6632,N_5792);
nand U7601 (N_7601,N_5313,N_5724);
or U7602 (N_7602,N_6724,N_6233);
nand U7603 (N_7603,N_5066,N_5112);
nand U7604 (N_7604,N_7351,N_6881);
and U7605 (N_7605,N_5355,N_6675);
or U7606 (N_7606,N_6376,N_5354);
xnor U7607 (N_7607,N_5074,N_5451);
nand U7608 (N_7608,N_7357,N_6694);
or U7609 (N_7609,N_7019,N_7415);
nor U7610 (N_7610,N_5275,N_5413);
nor U7611 (N_7611,N_6341,N_7476);
and U7612 (N_7612,N_5437,N_7144);
nor U7613 (N_7613,N_7358,N_5279);
nor U7614 (N_7614,N_6729,N_7323);
or U7615 (N_7615,N_5042,N_5020);
and U7616 (N_7616,N_6362,N_5730);
nand U7617 (N_7617,N_5399,N_5356);
nand U7618 (N_7618,N_6402,N_5417);
nor U7619 (N_7619,N_6825,N_6582);
nand U7620 (N_7620,N_6364,N_5073);
and U7621 (N_7621,N_5243,N_6350);
nor U7622 (N_7622,N_7171,N_5928);
nor U7623 (N_7623,N_5182,N_5611);
nand U7624 (N_7624,N_7461,N_5551);
or U7625 (N_7625,N_6559,N_5652);
or U7626 (N_7626,N_7091,N_6861);
nor U7627 (N_7627,N_5783,N_5903);
and U7628 (N_7628,N_6454,N_6941);
or U7629 (N_7629,N_6897,N_5263);
and U7630 (N_7630,N_5360,N_6505);
and U7631 (N_7631,N_7438,N_6610);
and U7632 (N_7632,N_5108,N_7035);
nor U7633 (N_7633,N_7048,N_5205);
and U7634 (N_7634,N_6224,N_5258);
or U7635 (N_7635,N_7256,N_5219);
or U7636 (N_7636,N_6331,N_6145);
nand U7637 (N_7637,N_6419,N_5160);
nor U7638 (N_7638,N_5118,N_7063);
or U7639 (N_7639,N_7016,N_5850);
or U7640 (N_7640,N_6305,N_5456);
or U7641 (N_7641,N_5155,N_7213);
nor U7642 (N_7642,N_5877,N_6065);
or U7643 (N_7643,N_7208,N_6777);
or U7644 (N_7644,N_6723,N_5726);
nand U7645 (N_7645,N_6474,N_7225);
or U7646 (N_7646,N_6568,N_7109);
and U7647 (N_7647,N_6616,N_5332);
nor U7648 (N_7648,N_5237,N_6835);
nor U7649 (N_7649,N_7081,N_5922);
nor U7650 (N_7650,N_5851,N_6496);
nor U7651 (N_7651,N_5369,N_6363);
nand U7652 (N_7652,N_5221,N_7240);
or U7653 (N_7653,N_5123,N_6473);
and U7654 (N_7654,N_6468,N_5766);
or U7655 (N_7655,N_6566,N_6097);
nand U7656 (N_7656,N_5240,N_7499);
or U7657 (N_7657,N_5546,N_5116);
nand U7658 (N_7658,N_6895,N_6338);
or U7659 (N_7659,N_6106,N_5880);
and U7660 (N_7660,N_7367,N_5212);
nand U7661 (N_7661,N_7231,N_6818);
nand U7662 (N_7662,N_7047,N_5996);
nor U7663 (N_7663,N_6112,N_7356);
nor U7664 (N_7664,N_7316,N_7153);
or U7665 (N_7665,N_6380,N_5075);
nor U7666 (N_7666,N_5830,N_6007);
and U7667 (N_7667,N_5786,N_5907);
or U7668 (N_7668,N_6183,N_6203);
or U7669 (N_7669,N_7404,N_5971);
nor U7670 (N_7670,N_5402,N_6803);
nand U7671 (N_7671,N_7282,N_6942);
nand U7672 (N_7672,N_6902,N_5498);
nor U7673 (N_7673,N_6535,N_6032);
and U7674 (N_7674,N_5007,N_6218);
and U7675 (N_7675,N_6492,N_6743);
and U7676 (N_7676,N_5040,N_5622);
nand U7677 (N_7677,N_6680,N_5658);
and U7678 (N_7678,N_6281,N_7391);
nor U7679 (N_7679,N_5651,N_7424);
nor U7680 (N_7680,N_6288,N_7400);
and U7681 (N_7681,N_5389,N_7409);
nand U7682 (N_7682,N_5098,N_5382);
nor U7683 (N_7683,N_5746,N_5091);
nor U7684 (N_7684,N_6022,N_5743);
nand U7685 (N_7685,N_5571,N_6719);
or U7686 (N_7686,N_6973,N_5010);
and U7687 (N_7687,N_6831,N_5583);
and U7688 (N_7688,N_6152,N_5699);
and U7689 (N_7689,N_5863,N_7307);
nand U7690 (N_7690,N_5896,N_5438);
or U7691 (N_7691,N_5348,N_7450);
nand U7692 (N_7692,N_5044,N_5597);
nand U7693 (N_7693,N_6588,N_5819);
nor U7694 (N_7694,N_6325,N_5852);
nor U7695 (N_7695,N_6494,N_6731);
nor U7696 (N_7696,N_5410,N_6545);
and U7697 (N_7697,N_5895,N_5196);
or U7698 (N_7698,N_5980,N_5028);
nor U7699 (N_7699,N_5078,N_7412);
nand U7700 (N_7700,N_5445,N_6245);
xor U7701 (N_7701,N_7227,N_7129);
xnor U7702 (N_7702,N_7224,N_6660);
or U7703 (N_7703,N_6303,N_7013);
or U7704 (N_7704,N_7432,N_5935);
and U7705 (N_7705,N_6714,N_7151);
nand U7706 (N_7706,N_6893,N_5841);
nand U7707 (N_7707,N_5343,N_5043);
and U7708 (N_7708,N_7290,N_6177);
nand U7709 (N_7709,N_6634,N_7181);
nand U7710 (N_7710,N_5139,N_5333);
and U7711 (N_7711,N_5486,N_6870);
and U7712 (N_7712,N_6046,N_7014);
xor U7713 (N_7713,N_5728,N_7492);
nor U7714 (N_7714,N_6828,N_7219);
or U7715 (N_7715,N_6383,N_5114);
and U7716 (N_7716,N_5729,N_7015);
or U7717 (N_7717,N_6324,N_5034);
xnor U7718 (N_7718,N_5801,N_6479);
and U7719 (N_7719,N_6763,N_6287);
nor U7720 (N_7720,N_6518,N_5273);
nor U7721 (N_7721,N_6079,N_7365);
or U7722 (N_7722,N_6732,N_5550);
nand U7723 (N_7723,N_5596,N_7377);
nand U7724 (N_7724,N_6433,N_6072);
or U7725 (N_7725,N_7350,N_6410);
and U7726 (N_7726,N_6008,N_5499);
nor U7727 (N_7727,N_6397,N_5158);
and U7728 (N_7728,N_5985,N_5945);
and U7729 (N_7729,N_5183,N_6925);
nand U7730 (N_7730,N_6948,N_6513);
or U7731 (N_7731,N_6432,N_5779);
or U7732 (N_7732,N_5146,N_5843);
and U7733 (N_7733,N_7223,N_7315);
nor U7734 (N_7734,N_6979,N_5342);
or U7735 (N_7735,N_6173,N_5119);
or U7736 (N_7736,N_7392,N_6238);
and U7737 (N_7737,N_6875,N_5798);
nor U7738 (N_7738,N_6579,N_6330);
and U7739 (N_7739,N_6059,N_6876);
or U7740 (N_7740,N_7102,N_5524);
nor U7741 (N_7741,N_5599,N_5302);
nor U7742 (N_7742,N_7027,N_7309);
nor U7743 (N_7743,N_5379,N_5968);
or U7744 (N_7744,N_7185,N_6544);
nor U7745 (N_7745,N_6569,N_6067);
or U7746 (N_7746,N_7294,N_7335);
nand U7747 (N_7747,N_5126,N_5308);
or U7748 (N_7748,N_5910,N_5521);
or U7749 (N_7749,N_6538,N_7259);
or U7750 (N_7750,N_6993,N_6100);
xor U7751 (N_7751,N_6787,N_7340);
or U7752 (N_7752,N_5105,N_5969);
or U7753 (N_7753,N_6796,N_6528);
nor U7754 (N_7754,N_6564,N_6042);
or U7755 (N_7755,N_6428,N_7475);
nor U7756 (N_7756,N_7332,N_5757);
nor U7757 (N_7757,N_7230,N_6879);
and U7758 (N_7758,N_7434,N_5689);
or U7759 (N_7759,N_5986,N_5548);
and U7760 (N_7760,N_6843,N_5898);
or U7761 (N_7761,N_6549,N_5489);
or U7762 (N_7762,N_5916,N_6241);
and U7763 (N_7763,N_5371,N_5660);
and U7764 (N_7764,N_5580,N_6178);
or U7765 (N_7765,N_5266,N_5452);
xor U7766 (N_7766,N_5061,N_6655);
nand U7767 (N_7767,N_5813,N_5566);
nor U7768 (N_7768,N_5937,N_5657);
and U7769 (N_7769,N_6312,N_5519);
nor U7770 (N_7770,N_6792,N_5787);
nand U7771 (N_7771,N_5125,N_6720);
and U7772 (N_7772,N_6726,N_5948);
and U7773 (N_7773,N_7361,N_6027);
or U7774 (N_7774,N_6758,N_7157);
nor U7775 (N_7775,N_5224,N_7397);
nand U7776 (N_7776,N_7337,N_6411);
nand U7777 (N_7777,N_7239,N_6366);
nand U7778 (N_7778,N_7473,N_5682);
and U7779 (N_7779,N_6011,N_7269);
or U7780 (N_7780,N_5997,N_5531);
nand U7781 (N_7781,N_6445,N_5785);
or U7782 (N_7782,N_5448,N_5908);
and U7783 (N_7783,N_5923,N_6936);
nor U7784 (N_7784,N_7135,N_6478);
nor U7785 (N_7785,N_6915,N_6650);
xor U7786 (N_7786,N_5799,N_7176);
nor U7787 (N_7787,N_7403,N_6797);
nand U7788 (N_7788,N_5469,N_6812);
nor U7789 (N_7789,N_7284,N_5432);
or U7790 (N_7790,N_7498,N_6980);
nand U7791 (N_7791,N_7241,N_5268);
and U7792 (N_7792,N_5323,N_6292);
and U7793 (N_7793,N_7453,N_5530);
nand U7794 (N_7794,N_5412,N_6130);
nand U7795 (N_7795,N_5733,N_5423);
nor U7796 (N_7796,N_5930,N_6681);
and U7797 (N_7797,N_7326,N_7348);
nand U7798 (N_7798,N_6399,N_6764);
or U7799 (N_7799,N_6127,N_7347);
nand U7800 (N_7800,N_5036,N_6458);
and U7801 (N_7801,N_6665,N_6147);
xnor U7802 (N_7802,N_6852,N_7460);
nand U7803 (N_7803,N_5686,N_5806);
or U7804 (N_7804,N_6028,N_5700);
and U7805 (N_7805,N_6710,N_7373);
nand U7806 (N_7806,N_6859,N_6486);
nor U7807 (N_7807,N_6430,N_5515);
nand U7808 (N_7808,N_7341,N_5336);
and U7809 (N_7809,N_6004,N_7168);
nor U7810 (N_7810,N_5192,N_5015);
or U7811 (N_7811,N_7463,N_5906);
or U7812 (N_7812,N_6208,N_5481);
or U7813 (N_7813,N_5305,N_6311);
or U7814 (N_7814,N_6377,N_5902);
nor U7815 (N_7815,N_7068,N_6896);
nor U7816 (N_7816,N_6594,N_5345);
and U7817 (N_7817,N_5848,N_5052);
or U7818 (N_7818,N_5140,N_6006);
nor U7819 (N_7819,N_6497,N_5939);
and U7820 (N_7820,N_6808,N_5178);
nor U7821 (N_7821,N_6601,N_5002);
or U7822 (N_7822,N_6157,N_6659);
nand U7823 (N_7823,N_7104,N_5321);
or U7824 (N_7824,N_7079,N_7108);
or U7825 (N_7825,N_6089,N_7023);
nand U7826 (N_7826,N_6176,N_6622);
and U7827 (N_7827,N_6965,N_5655);
nand U7828 (N_7828,N_6276,N_6563);
nor U7829 (N_7829,N_5561,N_6706);
nor U7830 (N_7830,N_7051,N_5001);
or U7831 (N_7831,N_5817,N_5009);
or U7832 (N_7832,N_5316,N_6817);
nor U7833 (N_7833,N_7296,N_6572);
and U7834 (N_7834,N_6320,N_6196);
nand U7835 (N_7835,N_5479,N_7036);
nor U7836 (N_7836,N_6237,N_6301);
or U7837 (N_7837,N_6009,N_7084);
nand U7838 (N_7838,N_5269,N_6142);
nand U7839 (N_7839,N_5491,N_5823);
nand U7840 (N_7840,N_7288,N_6277);
and U7841 (N_7841,N_6995,N_6539);
or U7842 (N_7842,N_6119,N_5918);
or U7843 (N_7843,N_5995,N_6969);
or U7844 (N_7844,N_6631,N_5404);
xor U7845 (N_7845,N_5246,N_6751);
nand U7846 (N_7846,N_5027,N_7369);
nand U7847 (N_7847,N_6395,N_6375);
and U7848 (N_7848,N_6037,N_6598);
nand U7849 (N_7849,N_5496,N_5712);
or U7850 (N_7850,N_7095,N_7008);
or U7851 (N_7851,N_5037,N_6854);
nor U7852 (N_7852,N_6991,N_6349);
and U7853 (N_7853,N_6798,N_5656);
and U7854 (N_7854,N_5185,N_7056);
nand U7855 (N_7855,N_7179,N_5478);
nor U7856 (N_7856,N_6235,N_6580);
or U7857 (N_7857,N_6839,N_6450);
nor U7858 (N_7858,N_5339,N_6511);
xnor U7859 (N_7859,N_7331,N_5966);
xnor U7860 (N_7860,N_6819,N_6901);
and U7861 (N_7861,N_6133,N_7101);
or U7862 (N_7862,N_6063,N_7310);
xor U7863 (N_7863,N_5816,N_5849);
nand U7864 (N_7864,N_6911,N_7413);
nor U7865 (N_7865,N_6023,N_5088);
or U7866 (N_7866,N_5528,N_7110);
nand U7867 (N_7867,N_7207,N_5483);
nor U7868 (N_7868,N_5606,N_6691);
and U7869 (N_7869,N_7186,N_6964);
or U7870 (N_7870,N_6955,N_5420);
nand U7871 (N_7871,N_7226,N_6298);
nor U7872 (N_7872,N_5705,N_6629);
and U7873 (N_7873,N_7164,N_6273);
nand U7874 (N_7874,N_7308,N_7021);
and U7875 (N_7875,N_7170,N_7339);
nand U7876 (N_7876,N_5623,N_5152);
nand U7877 (N_7877,N_5172,N_7467);
xor U7878 (N_7878,N_7464,N_5954);
and U7879 (N_7879,N_6414,N_6617);
nor U7880 (N_7880,N_6248,N_6213);
or U7881 (N_7881,N_5400,N_7345);
nor U7882 (N_7882,N_7086,N_5422);
nand U7883 (N_7883,N_5701,N_5847);
nand U7884 (N_7884,N_6701,N_6068);
or U7885 (N_7885,N_5698,N_6833);
nor U7886 (N_7886,N_7483,N_6830);
or U7887 (N_7887,N_6938,N_5326);
or U7888 (N_7888,N_7234,N_5681);
nor U7889 (N_7889,N_6978,N_7298);
or U7890 (N_7890,N_6999,N_5029);
nor U7891 (N_7891,N_6318,N_5790);
xnor U7892 (N_7892,N_6577,N_5854);
nor U7893 (N_7893,N_7177,N_6014);
or U7894 (N_7894,N_6765,N_6307);
nor U7895 (N_7895,N_5299,N_5291);
xor U7896 (N_7896,N_6773,N_6667);
or U7897 (N_7897,N_5145,N_6086);
or U7898 (N_7898,N_5624,N_5444);
or U7899 (N_7899,N_5385,N_5613);
or U7900 (N_7900,N_6933,N_5493);
nand U7901 (N_7901,N_5941,N_6618);
or U7902 (N_7902,N_6429,N_5708);
nand U7903 (N_7903,N_6250,N_6845);
and U7904 (N_7904,N_7488,N_6385);
or U7905 (N_7905,N_5472,N_5235);
or U7906 (N_7906,N_6927,N_5862);
and U7907 (N_7907,N_6744,N_5170);
or U7908 (N_7908,N_6913,N_7299);
nor U7909 (N_7909,N_6960,N_6874);
xnor U7910 (N_7910,N_5984,N_5855);
and U7911 (N_7911,N_5381,N_5516);
nand U7912 (N_7912,N_5663,N_5748);
nand U7913 (N_7913,N_5455,N_5654);
nor U7914 (N_7914,N_7055,N_7353);
or U7915 (N_7915,N_7359,N_6739);
or U7916 (N_7916,N_5386,N_5238);
and U7917 (N_7917,N_6489,N_5407);
nor U7918 (N_7918,N_6416,N_5859);
or U7919 (N_7919,N_7093,N_7437);
xor U7920 (N_7920,N_7440,N_5406);
and U7921 (N_7921,N_5179,N_6842);
and U7922 (N_7922,N_5820,N_5347);
and U7923 (N_7923,N_5359,N_7466);
nand U7924 (N_7924,N_5092,N_7130);
nor U7925 (N_7925,N_5264,N_5337);
and U7926 (N_7926,N_5331,N_5510);
nor U7927 (N_7927,N_5294,N_6256);
nor U7928 (N_7928,N_6459,N_6220);
nand U7929 (N_7929,N_5608,N_5041);
or U7930 (N_7930,N_7018,N_6207);
nor U7931 (N_7931,N_7007,N_7459);
nor U7932 (N_7932,N_6053,N_6405);
and U7933 (N_7933,N_6365,N_6158);
nand U7934 (N_7934,N_5867,N_7212);
nor U7935 (N_7935,N_6045,N_6730);
nor U7936 (N_7936,N_5208,N_5584);
nand U7937 (N_7937,N_6054,N_6871);
and U7938 (N_7938,N_6339,N_5206);
nand U7939 (N_7939,N_5436,N_5523);
or U7940 (N_7940,N_5211,N_5846);
nor U7941 (N_7941,N_6916,N_7199);
and U7942 (N_7942,N_5535,N_5893);
nand U7943 (N_7943,N_6384,N_7303);
nor U7944 (N_7944,N_6216,N_6484);
or U7945 (N_7945,N_5141,N_6304);
nand U7946 (N_7946,N_5070,N_6867);
and U7947 (N_7947,N_7100,N_6986);
nand U7948 (N_7948,N_5242,N_6774);
and U7949 (N_7949,N_6727,N_6426);
or U7950 (N_7950,N_5482,N_6961);
or U7951 (N_7951,N_5973,N_5419);
or U7952 (N_7952,N_6653,N_7285);
nor U7953 (N_7953,N_7074,N_6056);
or U7954 (N_7954,N_7220,N_6175);
and U7955 (N_7955,N_5772,N_7423);
nand U7956 (N_7956,N_6576,N_6776);
nand U7957 (N_7957,N_5319,N_6026);
nand U7958 (N_7958,N_5931,N_7280);
and U7959 (N_7959,N_6715,N_7117);
and U7960 (N_7960,N_5260,N_5718);
xor U7961 (N_7961,N_7266,N_5788);
nand U7962 (N_7962,N_5598,N_5947);
nor U7963 (N_7963,N_6025,N_5166);
or U7964 (N_7964,N_7494,N_6793);
and U7965 (N_7965,N_5870,N_5961);
and U7966 (N_7966,N_5679,N_6905);
nor U7967 (N_7967,N_6850,N_7472);
and U7968 (N_7968,N_6111,N_6868);
and U7969 (N_7969,N_6515,N_6699);
or U7970 (N_7970,N_5097,N_6533);
or U7971 (N_7971,N_6785,N_5731);
nor U7972 (N_7972,N_5307,N_5991);
and U7973 (N_7973,N_7158,N_7448);
nand U7974 (N_7974,N_5480,N_5573);
nand U7975 (N_7975,N_5396,N_6373);
nand U7976 (N_7976,N_7062,N_7362);
and U7977 (N_7977,N_5591,N_5460);
nor U7978 (N_7978,N_5740,N_6075);
nor U7979 (N_7979,N_6612,N_6171);
or U7980 (N_7980,N_5917,N_7270);
or U7981 (N_7981,N_7378,N_5513);
nand U7982 (N_7982,N_6930,N_6998);
or U7983 (N_7983,N_6306,N_5167);
and U7984 (N_7984,N_5349,N_7428);
or U7985 (N_7985,N_5769,N_6323);
and U7986 (N_7986,N_6663,N_5494);
or U7987 (N_7987,N_5579,N_6128);
or U7988 (N_7988,N_6195,N_6849);
or U7989 (N_7989,N_7318,N_6947);
nor U7990 (N_7990,N_5156,N_7190);
or U7991 (N_7991,N_6167,N_5645);
nor U7992 (N_7992,N_6010,N_6623);
nand U7993 (N_7993,N_5322,N_6529);
and U7994 (N_7994,N_5462,N_6020);
and U7995 (N_7995,N_6125,N_6226);
nor U7996 (N_7996,N_5318,N_5879);
or U7997 (N_7997,N_5542,N_6487);
nor U7998 (N_7998,N_5742,N_5831);
or U7999 (N_7999,N_6581,N_7305);
or U8000 (N_8000,N_6662,N_6262);
nand U8001 (N_8001,N_6123,N_6666);
or U8002 (N_8002,N_6636,N_7154);
or U8003 (N_8003,N_5233,N_6073);
nand U8004 (N_8004,N_5926,N_5134);
or U8005 (N_8005,N_6219,N_6705);
or U8006 (N_8006,N_6567,N_6589);
nor U8007 (N_8007,N_6752,N_6702);
and U8008 (N_8008,N_5750,N_6420);
xor U8009 (N_8009,N_5840,N_6738);
nand U8010 (N_8010,N_5934,N_6943);
nand U8011 (N_8011,N_6987,N_5811);
or U8012 (N_8012,N_6619,N_6573);
or U8013 (N_8013,N_5884,N_5887);
nor U8014 (N_8014,N_5065,N_6982);
and U8015 (N_8015,N_7037,N_6676);
or U8016 (N_8016,N_6712,N_5062);
nor U8017 (N_8017,N_7321,N_5175);
nand U8018 (N_8018,N_7405,N_5013);
or U8019 (N_8019,N_5590,N_5974);
nor U8020 (N_8020,N_6613,N_6558);
or U8021 (N_8021,N_6439,N_6635);
xor U8022 (N_8022,N_5048,N_6295);
or U8023 (N_8023,N_6590,N_5159);
nor U8024 (N_8024,N_5586,N_7024);
and U8025 (N_8025,N_7012,N_7237);
nand U8026 (N_8026,N_7491,N_6811);
nand U8027 (N_8027,N_7033,N_6268);
or U8028 (N_8028,N_6092,N_7444);
and U8029 (N_8029,N_5758,N_5285);
or U8030 (N_8030,N_6456,N_6932);
and U8031 (N_8031,N_5970,N_6161);
and U8032 (N_8032,N_7470,N_6766);
and U8033 (N_8033,N_6887,N_7289);
or U8034 (N_8034,N_6309,N_6252);
or U8035 (N_8035,N_7443,N_5711);
or U8036 (N_8036,N_7449,N_7401);
nor U8037 (N_8037,N_5755,N_6506);
nand U8038 (N_8038,N_5644,N_6525);
nor U8039 (N_8039,N_5232,N_6424);
nand U8040 (N_8040,N_6369,N_6593);
and U8041 (N_8041,N_6899,N_6614);
or U8042 (N_8042,N_7090,N_6215);
xnor U8043 (N_8043,N_7291,N_6584);
nor U8044 (N_8044,N_6404,N_5556);
nor U8045 (N_8045,N_5665,N_5680);
nor U8046 (N_8046,N_7139,N_5953);
and U8047 (N_8047,N_6784,N_5949);
nand U8048 (N_8048,N_6407,N_5087);
nor U8049 (N_8049,N_7194,N_6646);
nor U8050 (N_8050,N_6387,N_7136);
and U8051 (N_8051,N_7205,N_7149);
and U8052 (N_8052,N_6093,N_6786);
nand U8053 (N_8053,N_6482,N_7211);
or U8054 (N_8054,N_6374,N_5418);
nand U8055 (N_8055,N_6583,N_5567);
and U8056 (N_8056,N_5329,N_7381);
and U8057 (N_8057,N_6968,N_6039);
and U8058 (N_8058,N_5518,N_5957);
nor U8059 (N_8059,N_7342,N_5722);
xnor U8060 (N_8060,N_6750,N_7115);
or U8061 (N_8061,N_5587,N_7319);
and U8062 (N_8062,N_6150,N_6231);
nor U8063 (N_8063,N_7134,N_6735);
or U8064 (N_8064,N_7481,N_6199);
nor U8065 (N_8065,N_5671,N_6084);
nor U8066 (N_8066,N_5857,N_6695);
or U8067 (N_8067,N_7274,N_5920);
nand U8068 (N_8068,N_6661,N_5405);
nand U8069 (N_8069,N_6052,N_6963);
nor U8070 (N_8070,N_7099,N_5789);
nor U8071 (N_8071,N_6741,N_5912);
nand U8072 (N_8072,N_7174,N_6556);
nor U8073 (N_8073,N_6126,N_6447);
and U8074 (N_8074,N_6070,N_5129);
and U8075 (N_8075,N_6624,N_7411);
or U8076 (N_8076,N_5099,N_5593);
or U8077 (N_8077,N_6604,N_5216);
or U8078 (N_8078,N_6683,N_6342);
and U8079 (N_8079,N_6488,N_7487);
nor U8080 (N_8080,N_5505,N_5780);
nor U8081 (N_8081,N_6453,N_7173);
xnor U8082 (N_8082,N_5293,N_6700);
nand U8083 (N_8083,N_6082,N_7471);
nor U8084 (N_8084,N_5468,N_7271);
and U8085 (N_8085,N_6483,N_7128);
nand U8086 (N_8086,N_5194,N_6223);
nor U8087 (N_8087,N_5558,N_5330);
and U8088 (N_8088,N_5344,N_5719);
nor U8089 (N_8089,N_5180,N_6230);
and U8090 (N_8090,N_5128,N_5803);
and U8091 (N_8091,N_5540,N_5568);
nor U8092 (N_8092,N_5633,N_6674);
nand U8093 (N_8093,N_6547,N_7408);
nor U8094 (N_8094,N_7034,N_5955);
nor U8095 (N_8095,N_5670,N_6837);
and U8096 (N_8096,N_7420,N_5214);
or U8097 (N_8097,N_7087,N_5621);
and U8098 (N_8098,N_5944,N_6418);
nor U8099 (N_8099,N_6200,N_5807);
nor U8100 (N_8100,N_5666,N_5176);
nor U8101 (N_8101,N_6504,N_5781);
nand U8102 (N_8102,N_6560,N_6021);
nor U8103 (N_8103,N_6058,N_7040);
or U8104 (N_8104,N_5562,N_6278);
and U8105 (N_8105,N_5033,N_5324);
nand U8106 (N_8106,N_6031,N_7389);
nor U8107 (N_8107,N_5805,N_6664);
xnor U8108 (N_8108,N_5637,N_6865);
nor U8109 (N_8109,N_6253,N_6189);
or U8110 (N_8110,N_5415,N_5289);
nand U8111 (N_8111,N_6795,N_7001);
xnor U8112 (N_8112,N_6427,N_5527);
or U8113 (N_8113,N_6869,N_7486);
nand U8114 (N_8114,N_7417,N_5539);
or U8115 (N_8115,N_5340,N_7107);
nor U8116 (N_8116,N_6972,N_6555);
and U8117 (N_8117,N_5458,N_7071);
or U8118 (N_8118,N_6988,N_6452);
or U8119 (N_8119,N_6975,N_6754);
and U8120 (N_8120,N_7083,N_7229);
or U8121 (N_8121,N_7382,N_6953);
and U8122 (N_8122,N_6514,N_5200);
nand U8123 (N_8123,N_6678,N_7414);
or U8124 (N_8124,N_6652,N_6313);
nand U8125 (N_8125,N_7122,N_6587);
and U8126 (N_8126,N_5885,N_6912);
nand U8127 (N_8127,N_5122,N_5694);
and U8128 (N_8128,N_7328,N_5084);
nand U8129 (N_8129,N_7131,N_6534);
nand U8130 (N_8130,N_7060,N_5071);
and U8131 (N_8131,N_5244,N_5601);
nand U8132 (N_8132,N_6821,N_7322);
xor U8133 (N_8133,N_6160,N_7272);
and U8134 (N_8134,N_5605,N_6668);
nor U8135 (N_8135,N_5101,N_6047);
nand U8136 (N_8136,N_7141,N_5127);
nand U8137 (N_8137,N_6838,N_5791);
and U8138 (N_8138,N_5133,N_5760);
or U8139 (N_8139,N_7092,N_6148);
or U8140 (N_8140,N_5284,N_6585);
nand U8141 (N_8141,N_5303,N_6841);
or U8142 (N_8142,N_6327,N_5470);
and U8143 (N_8143,N_5998,N_6351);
nor U8144 (N_8144,N_5353,N_6222);
nand U8145 (N_8145,N_7393,N_7172);
nor U8146 (N_8146,N_5150,N_5187);
nand U8147 (N_8147,N_5821,N_7236);
nand U8148 (N_8148,N_7371,N_6926);
nand U8149 (N_8149,N_6300,N_5526);
nor U8150 (N_8150,N_5853,N_6813);
nand U8151 (N_8151,N_5504,N_7264);
xnor U8152 (N_8152,N_5164,N_6185);
or U8153 (N_8153,N_7260,N_6872);
nor U8154 (N_8154,N_5435,N_7191);
and U8155 (N_8155,N_6401,N_6378);
or U8156 (N_8156,N_5592,N_7155);
nand U8157 (N_8157,N_6194,N_6257);
and U8158 (N_8158,N_7072,N_5575);
nor U8159 (N_8159,N_6139,N_6791);
or U8160 (N_8160,N_7049,N_7416);
nand U8161 (N_8161,N_5677,N_5257);
or U8162 (N_8162,N_6608,N_7297);
or U8163 (N_8163,N_6168,N_5439);
and U8164 (N_8164,N_6149,N_7248);
nand U8165 (N_8165,N_5121,N_5314);
nand U8166 (N_8166,N_5829,N_7287);
nand U8167 (N_8167,N_6884,N_6209);
nor U8168 (N_8168,N_6061,N_5144);
nand U8169 (N_8169,N_7273,N_5943);
nand U8170 (N_8170,N_5749,N_7436);
nand U8171 (N_8171,N_5372,N_6451);
nand U8172 (N_8172,N_6711,N_5576);
nor U8173 (N_8173,N_5021,N_6562);
or U8174 (N_8174,N_6851,N_5664);
or U8175 (N_8175,N_6421,N_6759);
or U8176 (N_8176,N_5860,N_6266);
and U8177 (N_8177,N_6609,N_7043);
and U8178 (N_8178,N_5473,N_5398);
and U8179 (N_8179,N_6903,N_6319);
or U8180 (N_8180,N_5177,N_5977);
nor U8181 (N_8181,N_6244,N_7125);
nand U8182 (N_8182,N_6790,N_6788);
nand U8183 (N_8183,N_5311,N_6907);
nor U8184 (N_8184,N_5025,N_5085);
or U8185 (N_8185,N_6403,N_6285);
or U8186 (N_8186,N_5921,N_5032);
nor U8187 (N_8187,N_5102,N_7031);
nand U8188 (N_8188,N_5441,N_5634);
or U8189 (N_8189,N_5153,N_6190);
nand U8190 (N_8190,N_5570,N_5600);
and U8191 (N_8191,N_6055,N_5428);
nand U8192 (N_8192,N_5775,N_6463);
nand U8193 (N_8193,N_6314,N_7458);
nor U8194 (N_8194,N_6002,N_5804);
xor U8195 (N_8195,N_5442,N_6898);
nand U8196 (N_8196,N_5054,N_6212);
or U8197 (N_8197,N_5274,N_5304);
and U8198 (N_8198,N_6749,N_7425);
nor U8199 (N_8199,N_6883,N_6471);
nor U8200 (N_8200,N_6087,N_5721);
and U8201 (N_8201,N_5228,N_5770);
and U8202 (N_8202,N_6246,N_5296);
nor U8203 (N_8203,N_6400,N_7325);
nor U8204 (N_8204,N_5866,N_6800);
and U8205 (N_8205,N_6918,N_6491);
or U8206 (N_8206,N_5904,N_6206);
nor U8207 (N_8207,N_6360,N_5392);
nor U8208 (N_8208,N_5315,N_5604);
and U8209 (N_8209,N_5818,N_5195);
and U8210 (N_8210,N_5393,N_7252);
nor U8211 (N_8211,N_5557,N_6810);
nand U8212 (N_8212,N_5614,N_5842);
nand U8213 (N_8213,N_6141,N_5430);
xor U8214 (N_8214,N_6962,N_5254);
nand U8215 (N_8215,N_5014,N_7166);
and U8216 (N_8216,N_5068,N_5245);
or U8217 (N_8217,N_5776,N_7069);
and U8218 (N_8218,N_5016,N_5595);
and U8219 (N_8219,N_6503,N_5502);
or U8220 (N_8220,N_5023,N_6049);
and U8221 (N_8221,N_5295,N_5628);
nor U8222 (N_8222,N_6163,N_5373);
and U8223 (N_8223,N_7278,N_6099);
nand U8224 (N_8224,N_5143,N_5777);
or U8225 (N_8225,N_6641,N_5697);
and U8226 (N_8226,N_6789,N_5218);
and U8227 (N_8227,N_5762,N_5495);
nand U8228 (N_8228,N_6283,N_5383);
or U8229 (N_8229,N_6733,N_6193);
or U8230 (N_8230,N_7061,N_6957);
and U8231 (N_8231,N_6050,N_5873);
and U8232 (N_8232,N_5204,N_5135);
nand U8233 (N_8233,N_6931,N_7242);
and U8234 (N_8234,N_7004,N_6550);
nand U8235 (N_8235,N_7300,N_6297);
and U8236 (N_8236,N_6029,N_7374);
or U8237 (N_8237,N_5365,N_5282);
or U8238 (N_8238,N_5734,N_5110);
and U8239 (N_8239,N_6210,N_5358);
xnor U8240 (N_8240,N_5090,N_6827);
or U8241 (N_8241,N_6371,N_5874);
nor U8242 (N_8242,N_7159,N_7429);
or U8243 (N_8243,N_6956,N_6921);
and U8244 (N_8244,N_7344,N_7233);
and U8245 (N_8245,N_7070,N_5541);
and U8246 (N_8246,N_6967,N_6140);
or U8247 (N_8247,N_5889,N_6689);
nor U8248 (N_8248,N_6855,N_7442);
or U8249 (N_8249,N_7343,N_5325);
and U8250 (N_8250,N_5683,N_6466);
and U8251 (N_8251,N_5543,N_5485);
nand U8252 (N_8252,N_5626,N_7120);
nand U8253 (N_8253,N_6783,N_5149);
nand U8254 (N_8254,N_5411,N_5261);
or U8255 (N_8255,N_5301,N_5226);
and U8256 (N_8256,N_7313,N_6090);
xor U8257 (N_8257,N_7372,N_5267);
and U8258 (N_8258,N_5673,N_5038);
xor U8259 (N_8259,N_7202,N_5248);
nand U8260 (N_8260,N_6561,N_6527);
nor U8261 (N_8261,N_6094,N_6107);
or U8262 (N_8262,N_5572,N_5209);
and U8263 (N_8263,N_6151,N_6782);
nor U8264 (N_8264,N_5678,N_5832);
nor U8265 (N_8265,N_6018,N_6772);
nand U8266 (N_8266,N_6275,N_5662);
nor U8267 (N_8267,N_6415,N_5181);
nor U8268 (N_8268,N_5754,N_7418);
and U8269 (N_8269,N_7379,N_7253);
nor U8270 (N_8270,N_5454,N_6187);
nand U8271 (N_8271,N_7140,N_7195);
and U8272 (N_8272,N_6470,N_6908);
and U8273 (N_8273,N_6687,N_5171);
or U8274 (N_8274,N_6361,N_5736);
nor U8275 (N_8275,N_7126,N_5585);
or U8276 (N_8276,N_5501,N_7406);
and U8277 (N_8277,N_7368,N_5064);
or U8278 (N_8278,N_6048,N_6085);
nand U8279 (N_8279,N_5753,N_6906);
or U8280 (N_8280,N_7431,N_5229);
nor U8281 (N_8281,N_6853,N_7127);
nand U8282 (N_8282,N_6934,N_7469);
or U8283 (N_8283,N_6779,N_5650);
nand U8284 (N_8284,N_6542,N_7304);
nor U8285 (N_8285,N_5950,N_6051);
or U8286 (N_8286,N_7333,N_7390);
nor U8287 (N_8287,N_5271,N_7306);
or U8288 (N_8288,N_5207,N_7376);
nand U8289 (N_8289,N_6642,N_6367);
or U8290 (N_8290,N_6740,N_5100);
nand U8291 (N_8291,N_6103,N_5881);
and U8292 (N_8292,N_5901,N_5278);
nor U8293 (N_8293,N_6625,N_7192);
or U8294 (N_8294,N_5328,N_7113);
nor U8295 (N_8295,N_5076,N_5612);
or U8296 (N_8296,N_6165,N_5751);
or U8297 (N_8297,N_5565,N_7038);
or U8298 (N_8298,N_5836,N_6626);
nor U8299 (N_8299,N_7254,N_7352);
nor U8300 (N_8300,N_6078,N_5005);
and U8301 (N_8301,N_6502,N_6162);
or U8302 (N_8302,N_5197,N_5828);
and U8303 (N_8303,N_5704,N_5350);
and U8304 (N_8304,N_5773,N_5765);
nor U8305 (N_8305,N_6770,N_7238);
nand U8306 (N_8306,N_7066,N_6461);
nand U8307 (N_8307,N_5306,N_6657);
or U8308 (N_8308,N_6423,N_6816);
or U8309 (N_8309,N_6467,N_7067);
and U8310 (N_8310,N_6985,N_6229);
nand U8311 (N_8311,N_6270,N_5844);
or U8312 (N_8312,N_6638,N_5431);
nor U8313 (N_8313,N_7032,N_6820);
or U8314 (N_8314,N_5364,N_5104);
or U8315 (N_8315,N_6509,N_5376);
or U8316 (N_8316,N_7427,N_5707);
nand U8317 (N_8317,N_5560,N_7312);
nand U8318 (N_8318,N_5827,N_5544);
and U8319 (N_8319,N_6118,N_5225);
nand U8320 (N_8320,N_5559,N_5461);
nor U8321 (N_8321,N_6929,N_6690);
nor U8322 (N_8322,N_6279,N_5290);
nand U8323 (N_8323,N_6745,N_5978);
or U8324 (N_8324,N_7387,N_7146);
xnor U8325 (N_8325,N_5905,N_6799);
and U8326 (N_8326,N_7187,N_5900);
nand U8327 (N_8327,N_6442,N_5011);
nand U8328 (N_8328,N_5484,N_5894);
nor U8329 (N_8329,N_6413,N_5771);
nand U8330 (N_8330,N_6914,N_5627);
and U8331 (N_8331,N_6847,N_5312);
or U8332 (N_8332,N_7184,N_6994);
and U8333 (N_8333,N_6844,N_6408);
or U8334 (N_8334,N_6462,N_7292);
xnor U8335 (N_8335,N_7215,N_7073);
nand U8336 (N_8336,N_7042,N_6684);
and U8337 (N_8337,N_6264,N_7468);
and U8338 (N_8338,N_6296,N_6108);
and U8339 (N_8339,N_6062,N_6409);
or U8340 (N_8340,N_5334,N_7006);
nand U8341 (N_8341,N_5737,N_5635);
or U8342 (N_8342,N_5631,N_6794);
and U8343 (N_8343,N_7329,N_6615);
or U8344 (N_8344,N_6291,N_5026);
nor U8345 (N_8345,N_5174,N_7386);
and U8346 (N_8346,N_5629,N_6345);
nand U8347 (N_8347,N_5309,N_6254);
nand U8348 (N_8348,N_7088,N_6670);
nor U8349 (N_8349,N_6591,N_7020);
and U8350 (N_8350,N_6271,N_5547);
and U8351 (N_8351,N_7053,N_7311);
xor U8352 (N_8352,N_6095,N_6113);
or U8353 (N_8353,N_5822,N_5004);
nand U8354 (N_8354,N_6600,N_5131);
or U8355 (N_8355,N_6885,N_7178);
or U8356 (N_8356,N_6643,N_5380);
and U8357 (N_8357,N_5808,N_6390);
nor U8358 (N_8358,N_5045,N_5241);
nor U8359 (N_8359,N_7314,N_5691);
or U8360 (N_8360,N_7058,N_5825);
or U8361 (N_8361,N_7421,N_6443);
nor U8362 (N_8362,N_5838,N_6728);
or U8363 (N_8363,N_6546,N_6227);
nand U8364 (N_8364,N_7106,N_6000);
and U8365 (N_8365,N_6198,N_6894);
nor U8366 (N_8366,N_5675,N_7267);
nand U8367 (N_8367,N_7198,N_7465);
nand U8368 (N_8368,N_6121,N_6098);
and U8369 (N_8369,N_6074,N_5983);
nand U8370 (N_8370,N_6919,N_6599);
nor U8371 (N_8371,N_5933,N_5378);
and U8372 (N_8372,N_5739,N_7003);
or U8373 (N_8373,N_5793,N_5103);
nand U8374 (N_8374,N_6693,N_6769);
or U8375 (N_8375,N_7383,N_6472);
and U8376 (N_8376,N_7030,N_6682);
nor U8377 (N_8377,N_5554,N_5222);
and U8378 (N_8378,N_6060,N_6446);
or U8379 (N_8379,N_6204,N_7085);
and U8380 (N_8380,N_7446,N_6909);
nand U8381 (N_8381,N_5976,N_6398);
nand U8382 (N_8382,N_5500,N_7057);
and U8383 (N_8383,N_5837,N_6071);
or U8384 (N_8384,N_6565,N_6333);
and U8385 (N_8385,N_7148,N_7145);
or U8386 (N_8386,N_5946,N_7162);
and U8387 (N_8387,N_7165,N_5553);
or U8388 (N_8388,N_5956,N_6672);
nand U8389 (N_8389,N_5609,N_6249);
nand U8390 (N_8390,N_6526,N_5958);
nor U8391 (N_8391,N_5942,N_5377);
or U8392 (N_8392,N_7011,N_7349);
nor U8393 (N_8393,N_5702,N_5988);
nand U8394 (N_8394,N_5414,N_5063);
or U8395 (N_8395,N_6485,N_6234);
xor U8396 (N_8396,N_5619,N_5569);
nor U8397 (N_8397,N_5545,N_6586);
nand U8398 (N_8398,N_5839,N_7375);
nor U8399 (N_8399,N_6191,N_5690);
or U8400 (N_8400,N_6282,N_6976);
nand U8401 (N_8401,N_6396,N_5642);
nor U8402 (N_8402,N_5409,N_6357);
nor U8403 (N_8403,N_6348,N_5059);
nand U8404 (N_8404,N_6153,N_6144);
nand U8405 (N_8405,N_5298,N_7281);
and U8406 (N_8406,N_5477,N_5096);
and U8407 (N_8407,N_6937,N_6316);
nor U8408 (N_8408,N_5169,N_5695);
nor U8409 (N_8409,N_6044,N_5317);
nand U8410 (N_8410,N_7121,N_5723);
or U8411 (N_8411,N_5184,N_7258);
nor U8412 (N_8412,N_7457,N_6181);
and U8413 (N_8413,N_5148,N_6703);
nor U8414 (N_8414,N_5982,N_5812);
and U8415 (N_8415,N_6038,N_6814);
or U8416 (N_8416,N_5759,N_5617);
xnor U8417 (N_8417,N_7078,N_6076);
and U8418 (N_8418,N_5362,N_6970);
nor U8419 (N_8419,N_5151,N_6557);
xor U8420 (N_8420,N_5492,N_5833);
and U8421 (N_8421,N_6088,N_6860);
nand U8422 (N_8422,N_5856,N_6904);
or U8423 (N_8423,N_6352,N_6412);
nor U8424 (N_8424,N_6406,N_6620);
nor U8425 (N_8425,N_5162,N_6866);
nor U8426 (N_8426,N_6602,N_6597);
and U8427 (N_8427,N_7080,N_6946);
nor U8428 (N_8428,N_5810,N_5173);
and U8429 (N_8429,N_5897,N_6293);
or U8430 (N_8430,N_5199,N_5157);
and U8431 (N_8431,N_5602,N_5213);
nor U8432 (N_8432,N_6928,N_7046);
xor U8433 (N_8433,N_7123,N_5030);
and U8434 (N_8434,N_7119,N_7152);
nand U8435 (N_8435,N_5017,N_6255);
and U8436 (N_8436,N_6110,N_7354);
and U8437 (N_8437,N_6716,N_5095);
or U8438 (N_8438,N_7116,N_6201);
nor U8439 (N_8439,N_5989,N_6188);
or U8440 (N_8440,N_5834,N_5265);
or U8441 (N_8441,N_5727,N_7150);
nor U8442 (N_8442,N_6355,N_5276);
and U8443 (N_8443,N_5891,N_5138);
or U8444 (N_8444,N_6379,N_5716);
nor U8445 (N_8445,N_6757,N_6057);
nand U8446 (N_8446,N_5113,N_5057);
and U8447 (N_8447,N_7399,N_5338);
nor U8448 (N_8448,N_5051,N_6628);
nor U8449 (N_8449,N_5055,N_5459);
nand U8450 (N_8450,N_6358,N_5649);
xnor U8451 (N_8451,N_5661,N_6753);
or U8452 (N_8452,N_6272,N_6507);
or U8453 (N_8453,N_5457,N_6137);
or U8454 (N_8454,N_5351,N_6476);
or U8455 (N_8455,N_6801,N_5620);
and U8456 (N_8456,N_6780,N_6778);
and U8457 (N_8457,N_6033,N_7124);
nor U8458 (N_8458,N_5574,N_5993);
nor U8459 (N_8459,N_6725,N_5653);
or U8460 (N_8460,N_6356,N_5925);
nor U8461 (N_8461,N_7143,N_7324);
and U8462 (N_8462,N_6630,N_5286);
and U8463 (N_8463,N_7160,N_5083);
or U8464 (N_8464,N_5427,N_6251);
or U8465 (N_8465,N_5262,N_6391);
nor U8466 (N_8466,N_5511,N_5919);
nor U8467 (N_8467,N_5464,N_6832);
or U8468 (N_8468,N_5341,N_6718);
nand U8469 (N_8469,N_7275,N_6516);
or U8470 (N_8470,N_5959,N_6464);
or U8471 (N_8471,N_5534,N_6120);
nand U8472 (N_8472,N_5752,N_5768);
or U8473 (N_8473,N_5384,N_6992);
or U8474 (N_8474,N_5735,N_6321);
and U8475 (N_8475,N_6041,N_5555);
or U8476 (N_8476,N_5929,N_5990);
nor U8477 (N_8477,N_7114,N_6302);
and U8478 (N_8478,N_6434,N_6146);
and U8479 (N_8479,N_6329,N_6910);
nor U8480 (N_8480,N_7279,N_6388);
and U8481 (N_8481,N_7338,N_6621);
xnor U8482 (N_8482,N_5672,N_6958);
nand U8483 (N_8483,N_5506,N_5514);
nor U8484 (N_8484,N_6521,N_5253);
xnor U8485 (N_8485,N_7044,N_6981);
nor U8486 (N_8486,N_6804,N_5538);
and U8487 (N_8487,N_7495,N_7218);
xor U8488 (N_8488,N_5024,N_6578);
nor U8489 (N_8489,N_6334,N_6669);
nand U8490 (N_8490,N_6826,N_5738);
nand U8491 (N_8491,N_6105,N_7482);
nor U8492 (N_8492,N_5784,N_5747);
or U8493 (N_8493,N_5449,N_6704);
or U8494 (N_8494,N_6864,N_5165);
or U8495 (N_8495,N_6877,N_5234);
nand U8496 (N_8496,N_5465,N_5861);
nand U8497 (N_8497,N_6807,N_5882);
nor U8498 (N_8498,N_5987,N_6923);
nor U8499 (N_8499,N_7005,N_5111);
or U8500 (N_8500,N_5582,N_5994);
and U8501 (N_8501,N_5564,N_7041);
or U8502 (N_8502,N_5471,N_6815);
and U8503 (N_8503,N_7396,N_6134);
xor U8504 (N_8504,N_7283,N_5915);
nand U8505 (N_8505,N_6761,N_6202);
and U8506 (N_8506,N_6131,N_7050);
nand U8507 (N_8507,N_5421,N_6755);
and U8508 (N_8508,N_5031,N_6520);
or U8509 (N_8509,N_6846,N_6500);
nand U8510 (N_8510,N_7456,N_7188);
nor U8511 (N_8511,N_5676,N_5320);
or U8512 (N_8512,N_6924,N_6289);
and U8513 (N_8513,N_5154,N_7244);
and U8514 (N_8514,N_5077,N_5352);
nand U8515 (N_8515,N_7002,N_5280);
nand U8516 (N_8516,N_6322,N_5835);
nor U8517 (N_8517,N_5674,N_7221);
and U8518 (N_8518,N_6959,N_5081);
nand U8519 (N_8519,N_5532,N_5522);
nor U8520 (N_8520,N_5507,N_7366);
nor U8521 (N_8521,N_7197,N_5952);
and U8522 (N_8522,N_5335,N_7384);
or U8523 (N_8523,N_5646,N_6136);
nor U8524 (N_8524,N_6124,N_6003);
or U8525 (N_8525,N_5475,N_6205);
and U8526 (N_8526,N_7133,N_5450);
or U8527 (N_8527,N_6824,N_7263);
nor U8528 (N_8528,N_6554,N_5577);
nand U8529 (N_8529,N_6192,N_7077);
and U8530 (N_8530,N_6114,N_6104);
or U8531 (N_8531,N_5824,N_6552);
or U8532 (N_8532,N_6736,N_5395);
and U8533 (N_8533,N_7370,N_6834);
and U8534 (N_8534,N_6574,N_6592);
or U8535 (N_8535,N_7277,N_6156);
nor U8536 (N_8536,N_5357,N_6495);
and U8537 (N_8537,N_5641,N_6886);
nor U8538 (N_8538,N_5914,N_6603);
nand U8539 (N_8539,N_7455,N_6155);
nand U8540 (N_8540,N_7268,N_5992);
nand U8541 (N_8541,N_5089,N_6184);
or U8542 (N_8542,N_5006,N_6417);
nor U8543 (N_8543,N_7065,N_6166);
and U8544 (N_8544,N_5012,N_5797);
nor U8545 (N_8545,N_7452,N_5688);
xor U8546 (N_8546,N_6997,N_6242);
or U8547 (N_8547,N_6717,N_6438);
nor U8548 (N_8548,N_5778,N_5272);
and U8549 (N_8549,N_6232,N_6091);
nor U8550 (N_8550,N_5709,N_5669);
nand U8551 (N_8551,N_5363,N_7189);
nand U8552 (N_8552,N_6640,N_6083);
or U8553 (N_8553,N_7052,N_7222);
and U8554 (N_8554,N_7276,N_6159);
nor U8555 (N_8555,N_6989,N_7045);
or U8556 (N_8556,N_6290,N_6109);
and U8557 (N_8557,N_6858,N_7096);
or U8558 (N_8558,N_6654,N_5049);
nor U8559 (N_8559,N_6873,N_5490);
or U8560 (N_8560,N_5106,N_5047);
and U8561 (N_8561,N_5964,N_6344);
and U8562 (N_8562,N_6966,N_5408);
xor U8563 (N_8563,N_6882,N_5120);
xor U8564 (N_8564,N_6548,N_7426);
nand U8565 (N_8565,N_5239,N_6891);
and U8566 (N_8566,N_5361,N_6337);
nand U8567 (N_8567,N_6746,N_7232);
nor U8568 (N_8568,N_6064,N_6762);
nand U8569 (N_8569,N_6493,N_5080);
nor U8570 (N_8570,N_6359,N_5424);
or U8571 (N_8571,N_5761,N_6519);
or U8572 (N_8572,N_5890,N_6530);
and U8573 (N_8573,N_5774,N_5845);
and U8574 (N_8574,N_5715,N_7156);
and U8575 (N_8575,N_5189,N_7228);
or U8576 (N_8576,N_5115,N_5965);
or U8577 (N_8577,N_5815,N_6096);
nor U8578 (N_8578,N_6179,N_6677);
xor U8579 (N_8579,N_6671,N_6080);
nand U8580 (N_8580,N_5018,N_6225);
nand U8581 (N_8581,N_6477,N_6984);
nand U8582 (N_8582,N_6570,N_5981);
and U8583 (N_8583,N_5685,N_6214);
nor U8584 (N_8584,N_6510,N_7075);
and U8585 (N_8585,N_5795,N_6658);
and U8586 (N_8586,N_5132,N_5589);
nand U8587 (N_8587,N_5137,N_5794);
nand U8588 (N_8588,N_7302,N_6537);
nand U8589 (N_8589,N_5488,N_6922);
nor U8590 (N_8590,N_5639,N_6651);
nand U8591 (N_8591,N_7089,N_5706);
nand U8592 (N_8592,N_7485,N_6015);
and U8593 (N_8593,N_6531,N_6596);
and U8594 (N_8594,N_5394,N_7201);
nand U8595 (N_8595,N_6892,N_6679);
nor U8596 (N_8596,N_6983,N_5509);
and U8597 (N_8597,N_5578,N_6940);
nor U8598 (N_8598,N_5297,N_6017);
or U8599 (N_8599,N_6260,N_7039);
nor U8600 (N_8600,N_6686,N_6900);
nand U8601 (N_8601,N_7054,N_7454);
nand U8602 (N_8602,N_6685,N_6143);
nor U8603 (N_8603,N_7360,N_7445);
nor U8604 (N_8604,N_6522,N_5440);
nor U8605 (N_8605,N_5800,N_6862);
or U8606 (N_8606,N_7490,N_6217);
and U8607 (N_8607,N_6422,N_6243);
and U8608 (N_8608,N_6974,N_6269);
and U8609 (N_8609,N_6247,N_6637);
nor U8610 (N_8610,N_7477,N_6186);
nand U8611 (N_8611,N_6005,N_6267);
nor U8612 (N_8612,N_5193,N_6536);
nand U8613 (N_8613,N_7480,N_5503);
or U8614 (N_8614,N_6310,N_7251);
and U8615 (N_8615,N_5191,N_6294);
xnor U8616 (N_8616,N_6174,N_7193);
nor U8617 (N_8617,N_5391,N_7204);
or U8618 (N_8618,N_5210,N_5497);
and U8619 (N_8619,N_7250,N_7497);
or U8620 (N_8620,N_5453,N_5292);
or U8621 (N_8621,N_6013,N_5046);
or U8622 (N_8622,N_6532,N_5346);
nand U8623 (N_8623,N_5429,N_5367);
nand U8624 (N_8624,N_6490,N_6498);
and U8625 (N_8625,N_7059,N_5960);
nand U8626 (N_8626,N_7484,N_7209);
nand U8627 (N_8627,N_6649,N_5508);
nor U8628 (N_8628,N_6722,N_7447);
nand U8629 (N_8629,N_5067,N_7026);
nor U8630 (N_8630,N_6228,N_6644);
nand U8631 (N_8631,N_5387,N_6444);
nand U8632 (N_8632,N_6939,N_6299);
nor U8633 (N_8633,N_6540,N_6347);
and U8634 (N_8634,N_5255,N_5924);
or U8635 (N_8635,N_5249,N_5433);
nand U8636 (N_8636,N_6328,N_6315);
nor U8637 (N_8637,N_6996,N_7394);
nand U8638 (N_8638,N_5886,N_5251);
nor U8639 (N_8639,N_7395,N_7478);
and U8640 (N_8640,N_6627,N_5533);
nand U8641 (N_8641,N_7161,N_5927);
nand U8642 (N_8642,N_6848,N_7334);
nor U8643 (N_8643,N_6265,N_7474);
nand U8644 (N_8644,N_6449,N_6353);
nand U8645 (N_8645,N_5003,N_7022);
nand U8646 (N_8646,N_5186,N_6595);
nand U8647 (N_8647,N_7439,N_5327);
nand U8648 (N_8648,N_5865,N_5366);
nand U8649 (N_8649,N_7301,N_5696);
nand U8650 (N_8650,N_7245,N_6019);
nor U8651 (N_8651,N_5310,N_5220);
nand U8652 (N_8652,N_6697,N_6435);
nand U8653 (N_8653,N_6768,N_7286);
and U8654 (N_8654,N_6460,N_6809);
or U8655 (N_8655,N_6040,N_5632);
nand U8656 (N_8656,N_7138,N_5975);
nor U8657 (N_8657,N_6441,N_7255);
nand U8658 (N_8658,N_6805,N_6370);
nor U8659 (N_8659,N_7317,N_6392);
or U8660 (N_8660,N_5717,N_6284);
or U8661 (N_8661,N_5072,N_6605);
nor U8662 (N_8662,N_7010,N_6475);
or U8663 (N_8663,N_6129,N_6822);
and U8664 (N_8664,N_6132,N_5603);
or U8665 (N_8665,N_5911,N_5124);
or U8666 (N_8666,N_6878,N_7025);
or U8667 (N_8667,N_5416,N_5630);
or U8668 (N_8668,N_5872,N_7112);
and U8669 (N_8669,N_5913,N_6890);
nor U8670 (N_8670,N_5474,N_6036);
and U8671 (N_8671,N_5300,N_6035);
nor U8672 (N_8672,N_7206,N_7295);
nand U8673 (N_8673,N_5368,N_7441);
and U8674 (N_8674,N_5932,N_6553);
nor U8675 (N_8675,N_5374,N_5069);
and U8676 (N_8676,N_5231,N_7262);
nor U8677 (N_8677,N_5563,N_7246);
nor U8678 (N_8678,N_6122,N_6971);
nand U8679 (N_8679,N_6863,N_6707);
nand U8680 (N_8680,N_5000,N_6747);
nand U8681 (N_8681,N_5288,N_7419);
nand U8682 (N_8682,N_7017,N_7137);
nor U8683 (N_8683,N_5714,N_5079);
or U8684 (N_8684,N_6673,N_6440);
or U8685 (N_8685,N_6066,N_5972);
nor U8686 (N_8686,N_5058,N_7496);
nand U8687 (N_8687,N_5875,N_6920);
nor U8688 (N_8688,N_5594,N_5744);
and U8689 (N_8689,N_6115,N_5763);
and U8690 (N_8690,N_6756,N_5247);
nand U8691 (N_8691,N_5190,N_7028);
nand U8692 (N_8692,N_6455,N_6211);
and U8693 (N_8693,N_6880,N_7216);
or U8694 (N_8694,N_5588,N_7385);
or U8695 (N_8695,N_6393,N_6645);
and U8696 (N_8696,N_6116,N_5537);
and U8697 (N_8697,N_7249,N_6437);
and U8698 (N_8698,N_6571,N_6656);
nand U8699 (N_8699,N_6286,N_5082);
nand U8700 (N_8700,N_5636,N_6197);
and U8701 (N_8701,N_6154,N_7451);
and U8702 (N_8702,N_5201,N_5109);
nor U8703 (N_8703,N_5397,N_7430);
nor U8704 (N_8704,N_6840,N_6523);
nand U8705 (N_8705,N_5581,N_5607);
or U8706 (N_8706,N_6236,N_6172);
or U8707 (N_8707,N_6394,N_5615);
or U8708 (N_8708,N_7479,N_5019);
and U8709 (N_8709,N_7293,N_5060);
and U8710 (N_8710,N_5883,N_5713);
nor U8711 (N_8711,N_5647,N_6990);
nand U8712 (N_8712,N_5938,N_7196);
and U8713 (N_8713,N_5425,N_5117);
and U8714 (N_8714,N_6633,N_5525);
or U8715 (N_8715,N_7261,N_6857);
nand U8716 (N_8716,N_5370,N_5390);
and U8717 (N_8717,N_6077,N_5403);
or U8718 (N_8718,N_5463,N_5256);
and U8719 (N_8719,N_5466,N_6259);
and U8720 (N_8720,N_6737,N_5796);
or U8721 (N_8721,N_5086,N_7180);
or U8722 (N_8722,N_6368,N_6771);
and U8723 (N_8723,N_6030,N_7064);
nand U8724 (N_8724,N_5107,N_6436);
or U8725 (N_8725,N_5039,N_6709);
nand U8726 (N_8726,N_7435,N_6317);
and U8727 (N_8727,N_6501,N_5668);
nor U8728 (N_8728,N_6607,N_5270);
and U8729 (N_8729,N_5667,N_5640);
and U8730 (N_8730,N_5756,N_5979);
nand U8731 (N_8731,N_6802,N_6346);
and U8732 (N_8732,N_6748,N_5720);
nor U8733 (N_8733,N_7097,N_5161);
nand U8734 (N_8734,N_5223,N_5259);
and U8735 (N_8735,N_6389,N_5864);
and U8736 (N_8736,N_5725,N_7462);
nor U8737 (N_8737,N_5549,N_6945);
or U8738 (N_8738,N_5388,N_7363);
and U8739 (N_8739,N_5648,N_7105);
nor U8740 (N_8740,N_6767,N_6308);
nand U8741 (N_8741,N_5868,N_6949);
or U8742 (N_8742,N_7235,N_6952);
and U8743 (N_8743,N_7398,N_6823);
nand U8744 (N_8744,N_6280,N_6169);
and U8745 (N_8745,N_6340,N_6775);
or U8746 (N_8746,N_7402,N_5552);
and U8747 (N_8747,N_5940,N_5447);
and U8748 (N_8748,N_6944,N_7082);
or U8749 (N_8749,N_7355,N_6240);
or U8750 (N_8750,N_7340,N_7173);
nand U8751 (N_8751,N_6217,N_5870);
nand U8752 (N_8752,N_6186,N_6116);
nor U8753 (N_8753,N_6874,N_7128);
or U8754 (N_8754,N_5221,N_6573);
nand U8755 (N_8755,N_7419,N_5038);
or U8756 (N_8756,N_5163,N_6042);
nand U8757 (N_8757,N_7214,N_6065);
or U8758 (N_8758,N_5855,N_5860);
and U8759 (N_8759,N_5783,N_6695);
nand U8760 (N_8760,N_6310,N_6120);
nand U8761 (N_8761,N_7254,N_6349);
or U8762 (N_8762,N_5901,N_7194);
nand U8763 (N_8763,N_6915,N_6055);
nand U8764 (N_8764,N_6194,N_6541);
and U8765 (N_8765,N_5254,N_7309);
and U8766 (N_8766,N_7347,N_6866);
xor U8767 (N_8767,N_5152,N_6093);
and U8768 (N_8768,N_6955,N_5329);
nand U8769 (N_8769,N_7476,N_6735);
or U8770 (N_8770,N_7423,N_6225);
nand U8771 (N_8771,N_5877,N_6388);
nand U8772 (N_8772,N_5355,N_7020);
nor U8773 (N_8773,N_6272,N_6121);
nand U8774 (N_8774,N_6767,N_6778);
and U8775 (N_8775,N_5301,N_6874);
and U8776 (N_8776,N_5435,N_6302);
and U8777 (N_8777,N_7192,N_6111);
and U8778 (N_8778,N_7191,N_6058);
and U8779 (N_8779,N_6688,N_5536);
or U8780 (N_8780,N_5155,N_7394);
and U8781 (N_8781,N_5681,N_5659);
nand U8782 (N_8782,N_7078,N_6560);
nor U8783 (N_8783,N_6998,N_7391);
and U8784 (N_8784,N_6599,N_7177);
or U8785 (N_8785,N_7366,N_7066);
or U8786 (N_8786,N_6643,N_5218);
or U8787 (N_8787,N_7432,N_6870);
or U8788 (N_8788,N_5756,N_6622);
and U8789 (N_8789,N_6363,N_5940);
and U8790 (N_8790,N_5256,N_6152);
and U8791 (N_8791,N_6081,N_7031);
nor U8792 (N_8792,N_6584,N_5643);
and U8793 (N_8793,N_6751,N_5512);
and U8794 (N_8794,N_5171,N_5464);
nand U8795 (N_8795,N_5765,N_6862);
and U8796 (N_8796,N_6871,N_6608);
and U8797 (N_8797,N_5292,N_6056);
nand U8798 (N_8798,N_7059,N_6902);
nand U8799 (N_8799,N_6168,N_5636);
and U8800 (N_8800,N_5221,N_6723);
nand U8801 (N_8801,N_5091,N_5241);
nor U8802 (N_8802,N_6201,N_5666);
and U8803 (N_8803,N_5484,N_7157);
and U8804 (N_8804,N_7326,N_5598);
or U8805 (N_8805,N_7206,N_5992);
and U8806 (N_8806,N_5665,N_5632);
and U8807 (N_8807,N_6366,N_6625);
nor U8808 (N_8808,N_5487,N_6977);
nand U8809 (N_8809,N_7314,N_6275);
nand U8810 (N_8810,N_6417,N_6721);
nor U8811 (N_8811,N_6246,N_5797);
nor U8812 (N_8812,N_6842,N_6210);
nand U8813 (N_8813,N_5597,N_7151);
or U8814 (N_8814,N_6105,N_6523);
nor U8815 (N_8815,N_5935,N_5130);
nand U8816 (N_8816,N_7051,N_6724);
and U8817 (N_8817,N_5779,N_7494);
and U8818 (N_8818,N_5199,N_5201);
or U8819 (N_8819,N_5738,N_5043);
and U8820 (N_8820,N_5538,N_5105);
or U8821 (N_8821,N_5897,N_5417);
and U8822 (N_8822,N_6994,N_6065);
nand U8823 (N_8823,N_5141,N_6935);
nor U8824 (N_8824,N_6712,N_5306);
nor U8825 (N_8825,N_6325,N_5733);
or U8826 (N_8826,N_5617,N_6059);
or U8827 (N_8827,N_6826,N_7499);
or U8828 (N_8828,N_6504,N_7492);
nand U8829 (N_8829,N_6059,N_7231);
nand U8830 (N_8830,N_7433,N_6455);
and U8831 (N_8831,N_6937,N_5161);
and U8832 (N_8832,N_5271,N_5340);
or U8833 (N_8833,N_7287,N_7135);
nor U8834 (N_8834,N_6881,N_5496);
nor U8835 (N_8835,N_6851,N_5138);
nand U8836 (N_8836,N_6780,N_7096);
and U8837 (N_8837,N_6355,N_6302);
nand U8838 (N_8838,N_5791,N_6957);
and U8839 (N_8839,N_6199,N_6237);
or U8840 (N_8840,N_7438,N_7363);
and U8841 (N_8841,N_7269,N_6353);
nand U8842 (N_8842,N_6585,N_5591);
nand U8843 (N_8843,N_7017,N_5986);
nand U8844 (N_8844,N_6293,N_6682);
nand U8845 (N_8845,N_6425,N_6854);
or U8846 (N_8846,N_6686,N_7035);
and U8847 (N_8847,N_7195,N_6691);
and U8848 (N_8848,N_7053,N_6858);
or U8849 (N_8849,N_5499,N_6436);
and U8850 (N_8850,N_5228,N_5133);
nand U8851 (N_8851,N_5238,N_7012);
and U8852 (N_8852,N_6672,N_5410);
nand U8853 (N_8853,N_6495,N_7124);
nand U8854 (N_8854,N_6081,N_5306);
or U8855 (N_8855,N_6086,N_5685);
nand U8856 (N_8856,N_6097,N_5755);
or U8857 (N_8857,N_7242,N_7319);
and U8858 (N_8858,N_5865,N_5635);
nor U8859 (N_8859,N_5316,N_7081);
and U8860 (N_8860,N_7147,N_6475);
or U8861 (N_8861,N_6750,N_6925);
nand U8862 (N_8862,N_5787,N_7449);
xor U8863 (N_8863,N_6678,N_6438);
or U8864 (N_8864,N_5000,N_5165);
or U8865 (N_8865,N_5870,N_5868);
or U8866 (N_8866,N_5255,N_5145);
or U8867 (N_8867,N_6980,N_7457);
nand U8868 (N_8868,N_6590,N_5189);
xor U8869 (N_8869,N_7378,N_5360);
nor U8870 (N_8870,N_6237,N_5612);
or U8871 (N_8871,N_5881,N_5844);
nor U8872 (N_8872,N_6140,N_5423);
nand U8873 (N_8873,N_6688,N_6791);
or U8874 (N_8874,N_6722,N_5064);
nand U8875 (N_8875,N_6662,N_7043);
nor U8876 (N_8876,N_5720,N_5845);
xnor U8877 (N_8877,N_6135,N_6129);
nand U8878 (N_8878,N_6344,N_6611);
or U8879 (N_8879,N_5976,N_7309);
and U8880 (N_8880,N_5495,N_6491);
or U8881 (N_8881,N_6549,N_6590);
nand U8882 (N_8882,N_5279,N_6628);
or U8883 (N_8883,N_5710,N_6723);
nor U8884 (N_8884,N_6038,N_6716);
and U8885 (N_8885,N_6993,N_6291);
nor U8886 (N_8886,N_6577,N_5568);
and U8887 (N_8887,N_7096,N_5907);
nor U8888 (N_8888,N_5903,N_5453);
and U8889 (N_8889,N_5026,N_5562);
or U8890 (N_8890,N_5287,N_6512);
or U8891 (N_8891,N_6588,N_5166);
and U8892 (N_8892,N_7032,N_7472);
and U8893 (N_8893,N_6799,N_7414);
nand U8894 (N_8894,N_6756,N_5804);
nand U8895 (N_8895,N_5076,N_5965);
nand U8896 (N_8896,N_7241,N_6202);
and U8897 (N_8897,N_5555,N_6377);
nand U8898 (N_8898,N_6515,N_7297);
nor U8899 (N_8899,N_6586,N_7229);
and U8900 (N_8900,N_5897,N_6881);
and U8901 (N_8901,N_6371,N_5812);
and U8902 (N_8902,N_5277,N_6927);
nand U8903 (N_8903,N_6513,N_7201);
xor U8904 (N_8904,N_7134,N_5098);
or U8905 (N_8905,N_5679,N_7464);
nor U8906 (N_8906,N_7418,N_6556);
and U8907 (N_8907,N_6574,N_5127);
and U8908 (N_8908,N_6406,N_5523);
and U8909 (N_8909,N_5069,N_6830);
nor U8910 (N_8910,N_5449,N_5431);
nand U8911 (N_8911,N_6248,N_7224);
or U8912 (N_8912,N_5147,N_5527);
or U8913 (N_8913,N_5262,N_6926);
nand U8914 (N_8914,N_5130,N_6596);
xor U8915 (N_8915,N_7270,N_6280);
or U8916 (N_8916,N_6045,N_7006);
and U8917 (N_8917,N_5909,N_7139);
nand U8918 (N_8918,N_5386,N_5134);
nand U8919 (N_8919,N_5808,N_5246);
xor U8920 (N_8920,N_5424,N_5521);
nand U8921 (N_8921,N_6809,N_6433);
nor U8922 (N_8922,N_7149,N_5567);
nor U8923 (N_8923,N_7474,N_6461);
or U8924 (N_8924,N_5881,N_5883);
nor U8925 (N_8925,N_5543,N_6515);
and U8926 (N_8926,N_6778,N_6277);
and U8927 (N_8927,N_7264,N_5254);
nand U8928 (N_8928,N_5488,N_6476);
nor U8929 (N_8929,N_5670,N_6254);
nor U8930 (N_8930,N_5909,N_5487);
nand U8931 (N_8931,N_6597,N_7278);
and U8932 (N_8932,N_5447,N_5209);
or U8933 (N_8933,N_7184,N_6500);
and U8934 (N_8934,N_6151,N_5916);
nor U8935 (N_8935,N_7379,N_7488);
and U8936 (N_8936,N_6143,N_6579);
nand U8937 (N_8937,N_5960,N_7081);
and U8938 (N_8938,N_7394,N_5097);
nor U8939 (N_8939,N_6788,N_5998);
nor U8940 (N_8940,N_6755,N_5536);
and U8941 (N_8941,N_6234,N_7089);
nand U8942 (N_8942,N_7340,N_5862);
nand U8943 (N_8943,N_6084,N_6169);
and U8944 (N_8944,N_6513,N_6376);
nand U8945 (N_8945,N_5780,N_7205);
nand U8946 (N_8946,N_5709,N_5595);
nand U8947 (N_8947,N_7385,N_6577);
and U8948 (N_8948,N_7209,N_6202);
xor U8949 (N_8949,N_5265,N_5103);
and U8950 (N_8950,N_5612,N_7142);
and U8951 (N_8951,N_5718,N_5285);
xnor U8952 (N_8952,N_6392,N_6314);
or U8953 (N_8953,N_7056,N_7218);
or U8954 (N_8954,N_5687,N_6243);
or U8955 (N_8955,N_6422,N_6498);
nand U8956 (N_8956,N_5622,N_6487);
nand U8957 (N_8957,N_5475,N_6552);
or U8958 (N_8958,N_5938,N_5069);
xor U8959 (N_8959,N_6376,N_6976);
nor U8960 (N_8960,N_6315,N_6112);
or U8961 (N_8961,N_5637,N_7210);
nand U8962 (N_8962,N_6299,N_5940);
nand U8963 (N_8963,N_5109,N_6514);
nand U8964 (N_8964,N_6272,N_5129);
or U8965 (N_8965,N_6269,N_5116);
or U8966 (N_8966,N_5817,N_5066);
nand U8967 (N_8967,N_6249,N_5620);
and U8968 (N_8968,N_6891,N_7193);
or U8969 (N_8969,N_5240,N_5927);
nand U8970 (N_8970,N_5284,N_5430);
or U8971 (N_8971,N_6300,N_6172);
and U8972 (N_8972,N_6683,N_6146);
nand U8973 (N_8973,N_5883,N_6564);
xor U8974 (N_8974,N_5680,N_5966);
or U8975 (N_8975,N_6761,N_7211);
nor U8976 (N_8976,N_6616,N_6215);
nand U8977 (N_8977,N_7494,N_5164);
nor U8978 (N_8978,N_6024,N_5590);
nor U8979 (N_8979,N_6618,N_5386);
nor U8980 (N_8980,N_5368,N_5697);
or U8981 (N_8981,N_7421,N_6113);
and U8982 (N_8982,N_7246,N_6444);
nor U8983 (N_8983,N_7156,N_6709);
nand U8984 (N_8984,N_5571,N_5253);
and U8985 (N_8985,N_5871,N_6108);
and U8986 (N_8986,N_7038,N_5614);
or U8987 (N_8987,N_6600,N_5858);
and U8988 (N_8988,N_6112,N_6030);
nor U8989 (N_8989,N_6880,N_6224);
nand U8990 (N_8990,N_6107,N_7126);
nand U8991 (N_8991,N_5367,N_6716);
nor U8992 (N_8992,N_7372,N_6981);
nand U8993 (N_8993,N_6947,N_7413);
xor U8994 (N_8994,N_5322,N_7318);
and U8995 (N_8995,N_7251,N_5837);
or U8996 (N_8996,N_5067,N_7438);
xnor U8997 (N_8997,N_6465,N_7266);
nand U8998 (N_8998,N_5049,N_7206);
or U8999 (N_8999,N_7184,N_7428);
xor U9000 (N_9000,N_7115,N_7420);
nor U9001 (N_9001,N_6986,N_6299);
xor U9002 (N_9002,N_7089,N_6321);
nand U9003 (N_9003,N_6087,N_7453);
and U9004 (N_9004,N_5875,N_6888);
nand U9005 (N_9005,N_6345,N_6548);
nand U9006 (N_9006,N_5207,N_5369);
or U9007 (N_9007,N_5191,N_7208);
nand U9008 (N_9008,N_6010,N_5413);
or U9009 (N_9009,N_6274,N_7116);
nor U9010 (N_9010,N_6529,N_5093);
nand U9011 (N_9011,N_7238,N_6026);
nand U9012 (N_9012,N_6829,N_6112);
and U9013 (N_9013,N_6942,N_6459);
and U9014 (N_9014,N_5774,N_5856);
or U9015 (N_9015,N_5832,N_6644);
nand U9016 (N_9016,N_5823,N_6148);
or U9017 (N_9017,N_6609,N_7442);
and U9018 (N_9018,N_6019,N_5167);
or U9019 (N_9019,N_7356,N_7451);
nor U9020 (N_9020,N_5631,N_7308);
nor U9021 (N_9021,N_5135,N_5241);
or U9022 (N_9022,N_7221,N_5928);
and U9023 (N_9023,N_5072,N_5257);
or U9024 (N_9024,N_6125,N_7166);
or U9025 (N_9025,N_6635,N_6012);
or U9026 (N_9026,N_5433,N_6093);
nand U9027 (N_9027,N_7352,N_7048);
and U9028 (N_9028,N_7256,N_6526);
or U9029 (N_9029,N_6546,N_7154);
or U9030 (N_9030,N_6492,N_7438);
and U9031 (N_9031,N_6839,N_5637);
and U9032 (N_9032,N_6741,N_5493);
or U9033 (N_9033,N_7013,N_5062);
xnor U9034 (N_9034,N_6233,N_5208);
xor U9035 (N_9035,N_7211,N_5561);
and U9036 (N_9036,N_5658,N_6621);
and U9037 (N_9037,N_6377,N_5614);
or U9038 (N_9038,N_6867,N_7201);
nand U9039 (N_9039,N_5148,N_5693);
or U9040 (N_9040,N_7398,N_5785);
or U9041 (N_9041,N_5859,N_5611);
nor U9042 (N_9042,N_7372,N_7201);
nand U9043 (N_9043,N_6798,N_7232);
xor U9044 (N_9044,N_5798,N_7389);
nor U9045 (N_9045,N_6587,N_6945);
nor U9046 (N_9046,N_5444,N_5947);
nand U9047 (N_9047,N_6952,N_7028);
or U9048 (N_9048,N_6769,N_6050);
and U9049 (N_9049,N_5548,N_7280);
and U9050 (N_9050,N_5653,N_6186);
nand U9051 (N_9051,N_7332,N_7193);
or U9052 (N_9052,N_6945,N_7348);
or U9053 (N_9053,N_5070,N_6589);
and U9054 (N_9054,N_5508,N_5447);
nand U9055 (N_9055,N_5828,N_6944);
or U9056 (N_9056,N_7040,N_7222);
or U9057 (N_9057,N_6196,N_6526);
xor U9058 (N_9058,N_7488,N_6113);
or U9059 (N_9059,N_6232,N_6167);
or U9060 (N_9060,N_5555,N_7076);
and U9061 (N_9061,N_5759,N_5125);
nor U9062 (N_9062,N_5311,N_5155);
nor U9063 (N_9063,N_7480,N_5668);
or U9064 (N_9064,N_5753,N_7347);
or U9065 (N_9065,N_6569,N_5495);
nor U9066 (N_9066,N_7035,N_6245);
or U9067 (N_9067,N_7246,N_6956);
nor U9068 (N_9068,N_6092,N_5091);
nand U9069 (N_9069,N_6442,N_5164);
or U9070 (N_9070,N_5705,N_5787);
nand U9071 (N_9071,N_6439,N_6036);
and U9072 (N_9072,N_5024,N_6059);
nor U9073 (N_9073,N_6953,N_7100);
or U9074 (N_9074,N_6999,N_6412);
and U9075 (N_9075,N_6185,N_5293);
nor U9076 (N_9076,N_6456,N_5459);
and U9077 (N_9077,N_6412,N_5058);
nor U9078 (N_9078,N_6260,N_6306);
or U9079 (N_9079,N_7309,N_5291);
nor U9080 (N_9080,N_6342,N_6611);
nand U9081 (N_9081,N_7047,N_7002);
nand U9082 (N_9082,N_6215,N_5945);
and U9083 (N_9083,N_5289,N_5933);
nand U9084 (N_9084,N_6111,N_5891);
nor U9085 (N_9085,N_6692,N_6226);
nand U9086 (N_9086,N_5662,N_5476);
or U9087 (N_9087,N_5380,N_6884);
or U9088 (N_9088,N_5781,N_5015);
and U9089 (N_9089,N_6909,N_5331);
nor U9090 (N_9090,N_7174,N_7162);
and U9091 (N_9091,N_6230,N_6179);
and U9092 (N_9092,N_7358,N_7466);
xor U9093 (N_9093,N_7347,N_5143);
nor U9094 (N_9094,N_6991,N_5716);
nand U9095 (N_9095,N_7104,N_6633);
nand U9096 (N_9096,N_7206,N_5795);
and U9097 (N_9097,N_6068,N_7207);
nand U9098 (N_9098,N_5305,N_6877);
and U9099 (N_9099,N_6360,N_6171);
nand U9100 (N_9100,N_5917,N_6640);
nand U9101 (N_9101,N_6015,N_5704);
or U9102 (N_9102,N_7388,N_6052);
xnor U9103 (N_9103,N_6502,N_5049);
nand U9104 (N_9104,N_7378,N_5114);
nand U9105 (N_9105,N_5647,N_6053);
nand U9106 (N_9106,N_6999,N_6282);
nand U9107 (N_9107,N_5831,N_6386);
nor U9108 (N_9108,N_5110,N_7358);
nor U9109 (N_9109,N_7024,N_5531);
and U9110 (N_9110,N_7186,N_5035);
nand U9111 (N_9111,N_6379,N_6135);
and U9112 (N_9112,N_6107,N_5384);
and U9113 (N_9113,N_7404,N_6208);
or U9114 (N_9114,N_6390,N_5059);
nor U9115 (N_9115,N_6231,N_6074);
or U9116 (N_9116,N_5361,N_6265);
or U9117 (N_9117,N_5881,N_5662);
and U9118 (N_9118,N_5997,N_6662);
nor U9119 (N_9119,N_7037,N_7014);
nor U9120 (N_9120,N_6858,N_5641);
nor U9121 (N_9121,N_5099,N_5388);
or U9122 (N_9122,N_5906,N_6465);
or U9123 (N_9123,N_6197,N_5821);
nand U9124 (N_9124,N_6734,N_7442);
nor U9125 (N_9125,N_5618,N_5126);
nand U9126 (N_9126,N_6914,N_7254);
or U9127 (N_9127,N_5911,N_5722);
nor U9128 (N_9128,N_6447,N_5933);
nor U9129 (N_9129,N_7425,N_6035);
or U9130 (N_9130,N_6782,N_6801);
nand U9131 (N_9131,N_6093,N_5150);
or U9132 (N_9132,N_6601,N_6290);
nor U9133 (N_9133,N_5247,N_7230);
nand U9134 (N_9134,N_5779,N_6278);
nand U9135 (N_9135,N_7049,N_5747);
nor U9136 (N_9136,N_5573,N_7326);
and U9137 (N_9137,N_5746,N_7140);
or U9138 (N_9138,N_5520,N_5732);
and U9139 (N_9139,N_7480,N_7484);
nor U9140 (N_9140,N_6383,N_6004);
and U9141 (N_9141,N_7215,N_6294);
xnor U9142 (N_9142,N_5375,N_5711);
nand U9143 (N_9143,N_6023,N_7118);
nand U9144 (N_9144,N_5664,N_6298);
nor U9145 (N_9145,N_5789,N_5952);
and U9146 (N_9146,N_5330,N_5897);
and U9147 (N_9147,N_5804,N_6330);
nand U9148 (N_9148,N_6275,N_7165);
and U9149 (N_9149,N_6152,N_6284);
xor U9150 (N_9150,N_7019,N_7199);
and U9151 (N_9151,N_6685,N_5800);
and U9152 (N_9152,N_7041,N_5060);
and U9153 (N_9153,N_5141,N_6293);
or U9154 (N_9154,N_5259,N_5587);
and U9155 (N_9155,N_5319,N_6796);
nand U9156 (N_9156,N_6329,N_7056);
or U9157 (N_9157,N_5944,N_6344);
or U9158 (N_9158,N_6781,N_6570);
nor U9159 (N_9159,N_6433,N_6462);
or U9160 (N_9160,N_6417,N_6949);
or U9161 (N_9161,N_7190,N_7367);
nand U9162 (N_9162,N_6563,N_5757);
and U9163 (N_9163,N_5214,N_5257);
nor U9164 (N_9164,N_6861,N_6686);
nand U9165 (N_9165,N_6294,N_6100);
nor U9166 (N_9166,N_6496,N_5491);
nor U9167 (N_9167,N_6130,N_6015);
nand U9168 (N_9168,N_5282,N_5812);
or U9169 (N_9169,N_6953,N_6427);
and U9170 (N_9170,N_5041,N_6989);
nand U9171 (N_9171,N_6028,N_5276);
and U9172 (N_9172,N_5649,N_5430);
and U9173 (N_9173,N_7128,N_6261);
nor U9174 (N_9174,N_5322,N_5558);
nor U9175 (N_9175,N_5017,N_5242);
nor U9176 (N_9176,N_7261,N_5809);
nand U9177 (N_9177,N_6304,N_6580);
nand U9178 (N_9178,N_5241,N_5337);
or U9179 (N_9179,N_7054,N_5093);
nor U9180 (N_9180,N_5719,N_5548);
and U9181 (N_9181,N_5894,N_5165);
or U9182 (N_9182,N_6636,N_7367);
nand U9183 (N_9183,N_6447,N_5571);
nor U9184 (N_9184,N_7102,N_7045);
nand U9185 (N_9185,N_5789,N_7362);
and U9186 (N_9186,N_6127,N_5257);
and U9187 (N_9187,N_7126,N_5787);
nand U9188 (N_9188,N_7495,N_6347);
and U9189 (N_9189,N_6799,N_5736);
nand U9190 (N_9190,N_5345,N_6653);
nand U9191 (N_9191,N_5666,N_7402);
nor U9192 (N_9192,N_6352,N_6435);
nand U9193 (N_9193,N_6398,N_7166);
nand U9194 (N_9194,N_5234,N_6709);
nand U9195 (N_9195,N_6818,N_5624);
nor U9196 (N_9196,N_6705,N_6043);
or U9197 (N_9197,N_7024,N_7107);
or U9198 (N_9198,N_6915,N_6183);
and U9199 (N_9199,N_6592,N_6430);
nand U9200 (N_9200,N_5401,N_6119);
and U9201 (N_9201,N_7145,N_5725);
or U9202 (N_9202,N_5368,N_5112);
or U9203 (N_9203,N_6244,N_6275);
nor U9204 (N_9204,N_6340,N_6494);
and U9205 (N_9205,N_5265,N_7406);
nor U9206 (N_9206,N_6640,N_5644);
or U9207 (N_9207,N_6720,N_7038);
and U9208 (N_9208,N_5057,N_6555);
nand U9209 (N_9209,N_5855,N_7229);
nand U9210 (N_9210,N_5596,N_6738);
and U9211 (N_9211,N_6191,N_6128);
and U9212 (N_9212,N_6171,N_6177);
and U9213 (N_9213,N_6024,N_6935);
and U9214 (N_9214,N_5480,N_5914);
nand U9215 (N_9215,N_7033,N_5817);
nand U9216 (N_9216,N_5267,N_5739);
or U9217 (N_9217,N_6555,N_7087);
nor U9218 (N_9218,N_7020,N_6646);
nor U9219 (N_9219,N_5811,N_6927);
and U9220 (N_9220,N_5790,N_5308);
nor U9221 (N_9221,N_6095,N_6164);
or U9222 (N_9222,N_5180,N_5358);
and U9223 (N_9223,N_5255,N_6178);
or U9224 (N_9224,N_6975,N_6455);
nor U9225 (N_9225,N_5566,N_6501);
nor U9226 (N_9226,N_6325,N_5477);
nor U9227 (N_9227,N_7286,N_7383);
or U9228 (N_9228,N_7102,N_6724);
nor U9229 (N_9229,N_5228,N_6193);
and U9230 (N_9230,N_7316,N_7269);
and U9231 (N_9231,N_6841,N_7251);
or U9232 (N_9232,N_5829,N_6370);
or U9233 (N_9233,N_7126,N_6998);
nor U9234 (N_9234,N_7274,N_6380);
nor U9235 (N_9235,N_5498,N_5023);
nor U9236 (N_9236,N_5708,N_5812);
nand U9237 (N_9237,N_6756,N_6107);
nand U9238 (N_9238,N_6100,N_7108);
nand U9239 (N_9239,N_6213,N_5738);
or U9240 (N_9240,N_7001,N_5830);
nand U9241 (N_9241,N_5441,N_5192);
nand U9242 (N_9242,N_5726,N_7383);
or U9243 (N_9243,N_6993,N_5262);
nor U9244 (N_9244,N_6240,N_6261);
nand U9245 (N_9245,N_5778,N_7241);
nor U9246 (N_9246,N_6786,N_5283);
nor U9247 (N_9247,N_6694,N_6794);
nor U9248 (N_9248,N_6230,N_6995);
nand U9249 (N_9249,N_6547,N_6487);
or U9250 (N_9250,N_7461,N_5132);
and U9251 (N_9251,N_7141,N_6267);
or U9252 (N_9252,N_6273,N_6165);
or U9253 (N_9253,N_6413,N_6288);
or U9254 (N_9254,N_6660,N_7435);
nor U9255 (N_9255,N_5655,N_6462);
and U9256 (N_9256,N_5983,N_6642);
nand U9257 (N_9257,N_5706,N_6940);
or U9258 (N_9258,N_7435,N_7254);
and U9259 (N_9259,N_5067,N_5949);
nand U9260 (N_9260,N_6132,N_6401);
nor U9261 (N_9261,N_6238,N_6264);
nand U9262 (N_9262,N_6915,N_6378);
or U9263 (N_9263,N_5729,N_5871);
or U9264 (N_9264,N_6248,N_6171);
and U9265 (N_9265,N_7278,N_7327);
or U9266 (N_9266,N_7139,N_5313);
nor U9267 (N_9267,N_5946,N_5994);
nor U9268 (N_9268,N_5834,N_6266);
nand U9269 (N_9269,N_6747,N_7346);
and U9270 (N_9270,N_5227,N_7280);
nand U9271 (N_9271,N_5628,N_6093);
and U9272 (N_9272,N_5450,N_6970);
nor U9273 (N_9273,N_6194,N_5812);
and U9274 (N_9274,N_6068,N_5519);
nand U9275 (N_9275,N_6118,N_5729);
nor U9276 (N_9276,N_5917,N_7479);
or U9277 (N_9277,N_5275,N_7400);
nor U9278 (N_9278,N_7371,N_5557);
nand U9279 (N_9279,N_5270,N_5451);
and U9280 (N_9280,N_7362,N_5360);
nor U9281 (N_9281,N_6472,N_5078);
nand U9282 (N_9282,N_5410,N_7096);
nor U9283 (N_9283,N_5518,N_7327);
nor U9284 (N_9284,N_5784,N_6517);
and U9285 (N_9285,N_7107,N_7051);
nand U9286 (N_9286,N_7088,N_5150);
or U9287 (N_9287,N_5950,N_5945);
or U9288 (N_9288,N_5855,N_6153);
and U9289 (N_9289,N_5792,N_7074);
or U9290 (N_9290,N_5649,N_6816);
nand U9291 (N_9291,N_6803,N_6255);
or U9292 (N_9292,N_5559,N_6827);
and U9293 (N_9293,N_5863,N_6861);
nand U9294 (N_9294,N_6093,N_5251);
or U9295 (N_9295,N_5308,N_6560);
or U9296 (N_9296,N_6308,N_7281);
and U9297 (N_9297,N_6558,N_6408);
and U9298 (N_9298,N_5434,N_6673);
or U9299 (N_9299,N_6652,N_5522);
and U9300 (N_9300,N_7059,N_7407);
and U9301 (N_9301,N_6579,N_6603);
and U9302 (N_9302,N_7036,N_6237);
nor U9303 (N_9303,N_5808,N_5356);
and U9304 (N_9304,N_7078,N_6680);
nand U9305 (N_9305,N_6062,N_6520);
or U9306 (N_9306,N_7388,N_6531);
and U9307 (N_9307,N_6354,N_6313);
or U9308 (N_9308,N_7368,N_6885);
nor U9309 (N_9309,N_7330,N_7469);
nor U9310 (N_9310,N_7478,N_6536);
and U9311 (N_9311,N_5478,N_5421);
or U9312 (N_9312,N_6423,N_6446);
or U9313 (N_9313,N_5402,N_5273);
nor U9314 (N_9314,N_7203,N_6200);
or U9315 (N_9315,N_6639,N_6151);
and U9316 (N_9316,N_6747,N_7061);
nand U9317 (N_9317,N_5267,N_5784);
nand U9318 (N_9318,N_6691,N_7350);
or U9319 (N_9319,N_6007,N_6717);
nor U9320 (N_9320,N_6024,N_6064);
and U9321 (N_9321,N_5376,N_6361);
nor U9322 (N_9322,N_6416,N_6835);
and U9323 (N_9323,N_7287,N_7464);
and U9324 (N_9324,N_7137,N_7490);
nor U9325 (N_9325,N_5871,N_5245);
or U9326 (N_9326,N_7331,N_5609);
or U9327 (N_9327,N_5927,N_5938);
or U9328 (N_9328,N_5585,N_7420);
and U9329 (N_9329,N_5002,N_6262);
nor U9330 (N_9330,N_5377,N_6652);
nand U9331 (N_9331,N_6282,N_6249);
nor U9332 (N_9332,N_6660,N_5765);
or U9333 (N_9333,N_5488,N_6935);
nor U9334 (N_9334,N_6344,N_6996);
and U9335 (N_9335,N_6202,N_5200);
nand U9336 (N_9336,N_5831,N_7404);
or U9337 (N_9337,N_5256,N_5450);
nand U9338 (N_9338,N_5209,N_6474);
nand U9339 (N_9339,N_6456,N_5192);
and U9340 (N_9340,N_5091,N_5787);
nand U9341 (N_9341,N_5753,N_6379);
nor U9342 (N_9342,N_6420,N_7151);
and U9343 (N_9343,N_5574,N_7202);
nor U9344 (N_9344,N_5422,N_5786);
nand U9345 (N_9345,N_5785,N_5576);
or U9346 (N_9346,N_6159,N_5290);
or U9347 (N_9347,N_5784,N_6540);
and U9348 (N_9348,N_5833,N_5637);
or U9349 (N_9349,N_5308,N_5502);
or U9350 (N_9350,N_6990,N_5870);
nand U9351 (N_9351,N_6256,N_6876);
or U9352 (N_9352,N_7464,N_6518);
or U9353 (N_9353,N_7253,N_7292);
and U9354 (N_9354,N_6069,N_7265);
nor U9355 (N_9355,N_5847,N_6695);
and U9356 (N_9356,N_6433,N_5559);
nor U9357 (N_9357,N_6635,N_7385);
nand U9358 (N_9358,N_6536,N_6807);
nor U9359 (N_9359,N_7166,N_7291);
or U9360 (N_9360,N_5156,N_5418);
nand U9361 (N_9361,N_6266,N_5673);
nand U9362 (N_9362,N_5839,N_7158);
nand U9363 (N_9363,N_6211,N_5250);
or U9364 (N_9364,N_6570,N_7492);
and U9365 (N_9365,N_5177,N_6495);
or U9366 (N_9366,N_7134,N_6496);
or U9367 (N_9367,N_6572,N_5707);
nand U9368 (N_9368,N_5759,N_6236);
and U9369 (N_9369,N_6370,N_6858);
nor U9370 (N_9370,N_5943,N_6017);
nor U9371 (N_9371,N_6642,N_6311);
nand U9372 (N_9372,N_6965,N_6556);
nand U9373 (N_9373,N_6313,N_5586);
nand U9374 (N_9374,N_7041,N_7127);
nor U9375 (N_9375,N_5003,N_5321);
nand U9376 (N_9376,N_6946,N_5907);
or U9377 (N_9377,N_5279,N_6147);
or U9378 (N_9378,N_7491,N_7104);
nor U9379 (N_9379,N_5633,N_6375);
and U9380 (N_9380,N_6048,N_5567);
nor U9381 (N_9381,N_5562,N_5446);
or U9382 (N_9382,N_6280,N_6391);
nand U9383 (N_9383,N_6168,N_5332);
and U9384 (N_9384,N_6601,N_5740);
nand U9385 (N_9385,N_5555,N_6964);
or U9386 (N_9386,N_5035,N_6489);
and U9387 (N_9387,N_5042,N_7183);
or U9388 (N_9388,N_5037,N_5678);
nor U9389 (N_9389,N_6847,N_6376);
nand U9390 (N_9390,N_6739,N_6369);
and U9391 (N_9391,N_6950,N_7124);
nor U9392 (N_9392,N_6120,N_5518);
nor U9393 (N_9393,N_7406,N_5628);
and U9394 (N_9394,N_7463,N_6397);
xor U9395 (N_9395,N_7339,N_5370);
and U9396 (N_9396,N_6295,N_7398);
nand U9397 (N_9397,N_5284,N_5429);
nor U9398 (N_9398,N_5983,N_6208);
nand U9399 (N_9399,N_7491,N_7355);
nor U9400 (N_9400,N_5339,N_7122);
xnor U9401 (N_9401,N_5299,N_6856);
nand U9402 (N_9402,N_6539,N_6201);
and U9403 (N_9403,N_6709,N_6249);
and U9404 (N_9404,N_5216,N_6562);
and U9405 (N_9405,N_5490,N_7393);
or U9406 (N_9406,N_7056,N_6537);
nand U9407 (N_9407,N_7015,N_6380);
or U9408 (N_9408,N_5796,N_7275);
and U9409 (N_9409,N_5284,N_7097);
nand U9410 (N_9410,N_6707,N_5946);
or U9411 (N_9411,N_6413,N_5462);
nand U9412 (N_9412,N_5712,N_6410);
or U9413 (N_9413,N_6863,N_7439);
or U9414 (N_9414,N_5289,N_5195);
and U9415 (N_9415,N_5060,N_6269);
nor U9416 (N_9416,N_5198,N_7251);
and U9417 (N_9417,N_6325,N_6058);
and U9418 (N_9418,N_6217,N_5500);
or U9419 (N_9419,N_7439,N_6107);
nand U9420 (N_9420,N_6747,N_6509);
or U9421 (N_9421,N_5231,N_6362);
and U9422 (N_9422,N_7123,N_5297);
xor U9423 (N_9423,N_6440,N_6832);
nand U9424 (N_9424,N_5071,N_5062);
nor U9425 (N_9425,N_6985,N_7401);
nand U9426 (N_9426,N_7397,N_6321);
or U9427 (N_9427,N_5807,N_6601);
nor U9428 (N_9428,N_6889,N_6266);
or U9429 (N_9429,N_6757,N_6678);
and U9430 (N_9430,N_5661,N_7334);
nor U9431 (N_9431,N_7256,N_7285);
nor U9432 (N_9432,N_7372,N_6050);
and U9433 (N_9433,N_7409,N_5001);
or U9434 (N_9434,N_7283,N_6806);
and U9435 (N_9435,N_6220,N_5711);
and U9436 (N_9436,N_5276,N_7253);
and U9437 (N_9437,N_6463,N_6556);
nand U9438 (N_9438,N_5202,N_7226);
or U9439 (N_9439,N_5356,N_6149);
and U9440 (N_9440,N_6831,N_5427);
and U9441 (N_9441,N_5303,N_6345);
and U9442 (N_9442,N_6553,N_7048);
nand U9443 (N_9443,N_6122,N_5459);
nor U9444 (N_9444,N_5704,N_5670);
nor U9445 (N_9445,N_6253,N_5083);
or U9446 (N_9446,N_6402,N_5608);
or U9447 (N_9447,N_7155,N_6629);
nand U9448 (N_9448,N_5037,N_5460);
or U9449 (N_9449,N_6455,N_6863);
nor U9450 (N_9450,N_5366,N_5405);
nor U9451 (N_9451,N_5264,N_7276);
or U9452 (N_9452,N_5289,N_5028);
nand U9453 (N_9453,N_5495,N_6823);
and U9454 (N_9454,N_6862,N_6866);
nand U9455 (N_9455,N_6752,N_5681);
nand U9456 (N_9456,N_6973,N_6404);
xnor U9457 (N_9457,N_6780,N_6150);
nand U9458 (N_9458,N_5290,N_6346);
nand U9459 (N_9459,N_7452,N_6536);
nand U9460 (N_9460,N_6598,N_5704);
nor U9461 (N_9461,N_7124,N_7167);
and U9462 (N_9462,N_6363,N_7499);
or U9463 (N_9463,N_5501,N_6747);
and U9464 (N_9464,N_6347,N_7068);
and U9465 (N_9465,N_5367,N_5080);
nor U9466 (N_9466,N_6923,N_5947);
nor U9467 (N_9467,N_5875,N_7376);
nor U9468 (N_9468,N_6806,N_5596);
nand U9469 (N_9469,N_5221,N_7046);
or U9470 (N_9470,N_5022,N_5383);
or U9471 (N_9471,N_5843,N_6799);
xnor U9472 (N_9472,N_6434,N_5895);
and U9473 (N_9473,N_7118,N_5165);
or U9474 (N_9474,N_7296,N_5377);
nand U9475 (N_9475,N_6380,N_6495);
nand U9476 (N_9476,N_6380,N_5824);
or U9477 (N_9477,N_6785,N_7108);
nand U9478 (N_9478,N_5341,N_5238);
and U9479 (N_9479,N_6350,N_7038);
and U9480 (N_9480,N_6299,N_6650);
nor U9481 (N_9481,N_5422,N_6722);
xor U9482 (N_9482,N_5285,N_6687);
nor U9483 (N_9483,N_6163,N_5036);
or U9484 (N_9484,N_5143,N_6459);
nand U9485 (N_9485,N_7269,N_7085);
or U9486 (N_9486,N_5744,N_5101);
or U9487 (N_9487,N_7286,N_5236);
or U9488 (N_9488,N_7364,N_6855);
nand U9489 (N_9489,N_5163,N_6414);
or U9490 (N_9490,N_6913,N_6139);
or U9491 (N_9491,N_5676,N_5811);
or U9492 (N_9492,N_6915,N_6970);
xnor U9493 (N_9493,N_5430,N_5220);
and U9494 (N_9494,N_7202,N_5594);
nor U9495 (N_9495,N_7452,N_5282);
or U9496 (N_9496,N_6888,N_5879);
and U9497 (N_9497,N_7126,N_5746);
or U9498 (N_9498,N_6099,N_6775);
and U9499 (N_9499,N_6282,N_5730);
and U9500 (N_9500,N_6900,N_7457);
nand U9501 (N_9501,N_5461,N_5533);
or U9502 (N_9502,N_6319,N_5790);
and U9503 (N_9503,N_6912,N_6962);
nand U9504 (N_9504,N_6713,N_5269);
and U9505 (N_9505,N_6791,N_5312);
nand U9506 (N_9506,N_6079,N_5857);
or U9507 (N_9507,N_5333,N_5943);
and U9508 (N_9508,N_7374,N_5203);
and U9509 (N_9509,N_5626,N_6156);
nor U9510 (N_9510,N_7294,N_7045);
and U9511 (N_9511,N_5469,N_5850);
and U9512 (N_9512,N_7293,N_5587);
xnor U9513 (N_9513,N_7193,N_5663);
or U9514 (N_9514,N_6350,N_5967);
or U9515 (N_9515,N_6025,N_6316);
and U9516 (N_9516,N_6342,N_5052);
nand U9517 (N_9517,N_5778,N_6320);
nor U9518 (N_9518,N_5820,N_5175);
and U9519 (N_9519,N_6802,N_6578);
nand U9520 (N_9520,N_6598,N_7170);
and U9521 (N_9521,N_5352,N_5229);
nand U9522 (N_9522,N_6517,N_7169);
nand U9523 (N_9523,N_6857,N_5033);
nand U9524 (N_9524,N_5350,N_6379);
and U9525 (N_9525,N_6685,N_5883);
xor U9526 (N_9526,N_7146,N_6418);
and U9527 (N_9527,N_7335,N_6942);
nand U9528 (N_9528,N_6168,N_5228);
and U9529 (N_9529,N_5393,N_5118);
nand U9530 (N_9530,N_6310,N_6955);
or U9531 (N_9531,N_5578,N_6357);
nand U9532 (N_9532,N_5568,N_5091);
nand U9533 (N_9533,N_7494,N_7117);
xor U9534 (N_9534,N_5550,N_5425);
nand U9535 (N_9535,N_7249,N_6098);
or U9536 (N_9536,N_5823,N_7269);
and U9537 (N_9537,N_5358,N_5192);
or U9538 (N_9538,N_7161,N_5677);
nor U9539 (N_9539,N_7361,N_5370);
or U9540 (N_9540,N_6627,N_5228);
and U9541 (N_9541,N_6132,N_6583);
nor U9542 (N_9542,N_6694,N_5770);
or U9543 (N_9543,N_5341,N_6756);
xnor U9544 (N_9544,N_6137,N_5293);
nor U9545 (N_9545,N_6952,N_7101);
nor U9546 (N_9546,N_5831,N_7480);
or U9547 (N_9547,N_6117,N_5039);
or U9548 (N_9548,N_5293,N_6193);
nor U9549 (N_9549,N_7049,N_7406);
and U9550 (N_9550,N_6648,N_7464);
nand U9551 (N_9551,N_6303,N_6359);
or U9552 (N_9552,N_7102,N_5760);
nor U9553 (N_9553,N_5809,N_6698);
nand U9554 (N_9554,N_6436,N_6840);
and U9555 (N_9555,N_6076,N_6029);
and U9556 (N_9556,N_6577,N_7077);
xor U9557 (N_9557,N_7279,N_5707);
nor U9558 (N_9558,N_5195,N_6335);
and U9559 (N_9559,N_6578,N_5188);
and U9560 (N_9560,N_7305,N_5631);
nor U9561 (N_9561,N_6430,N_6209);
or U9562 (N_9562,N_7439,N_7220);
and U9563 (N_9563,N_5496,N_6171);
nor U9564 (N_9564,N_5364,N_5621);
nand U9565 (N_9565,N_6241,N_6785);
or U9566 (N_9566,N_5242,N_5635);
nand U9567 (N_9567,N_7248,N_5243);
and U9568 (N_9568,N_5539,N_6427);
nor U9569 (N_9569,N_6948,N_7259);
nor U9570 (N_9570,N_6497,N_7040);
xnor U9571 (N_9571,N_7159,N_5850);
nor U9572 (N_9572,N_6935,N_5772);
or U9573 (N_9573,N_5569,N_6079);
and U9574 (N_9574,N_5497,N_5041);
nand U9575 (N_9575,N_6013,N_6713);
and U9576 (N_9576,N_6778,N_6929);
nand U9577 (N_9577,N_5587,N_5809);
and U9578 (N_9578,N_5184,N_7472);
nand U9579 (N_9579,N_7220,N_6559);
nor U9580 (N_9580,N_6933,N_5585);
nand U9581 (N_9581,N_7404,N_6665);
nor U9582 (N_9582,N_5879,N_7083);
nor U9583 (N_9583,N_5487,N_7210);
and U9584 (N_9584,N_7251,N_6917);
or U9585 (N_9585,N_6489,N_7076);
or U9586 (N_9586,N_5320,N_6332);
xnor U9587 (N_9587,N_6300,N_5580);
nor U9588 (N_9588,N_6507,N_6461);
nor U9589 (N_9589,N_5564,N_6520);
or U9590 (N_9590,N_6067,N_6925);
nor U9591 (N_9591,N_6976,N_5284);
nand U9592 (N_9592,N_6299,N_5603);
or U9593 (N_9593,N_6604,N_6542);
nor U9594 (N_9594,N_5440,N_5980);
nor U9595 (N_9595,N_7000,N_6058);
nand U9596 (N_9596,N_7053,N_5757);
nand U9597 (N_9597,N_5332,N_7191);
xnor U9598 (N_9598,N_7351,N_7327);
or U9599 (N_9599,N_6558,N_5805);
and U9600 (N_9600,N_7213,N_5701);
nand U9601 (N_9601,N_7237,N_6583);
nand U9602 (N_9602,N_5162,N_7399);
and U9603 (N_9603,N_6969,N_6372);
nor U9604 (N_9604,N_6519,N_6994);
and U9605 (N_9605,N_5349,N_5695);
nand U9606 (N_9606,N_5017,N_6010);
and U9607 (N_9607,N_5664,N_5079);
or U9608 (N_9608,N_7303,N_7275);
nand U9609 (N_9609,N_5015,N_5535);
and U9610 (N_9610,N_5726,N_7253);
nand U9611 (N_9611,N_7187,N_7029);
nor U9612 (N_9612,N_5769,N_6144);
or U9613 (N_9613,N_6675,N_7099);
and U9614 (N_9614,N_6669,N_5667);
nand U9615 (N_9615,N_7423,N_7064);
nor U9616 (N_9616,N_5500,N_5663);
and U9617 (N_9617,N_5768,N_5591);
nor U9618 (N_9618,N_6860,N_7161);
nor U9619 (N_9619,N_6702,N_6041);
or U9620 (N_9620,N_7156,N_5510);
or U9621 (N_9621,N_5400,N_6050);
or U9622 (N_9622,N_5658,N_5716);
nor U9623 (N_9623,N_5078,N_5493);
and U9624 (N_9624,N_6185,N_6790);
nand U9625 (N_9625,N_7340,N_7270);
and U9626 (N_9626,N_6638,N_5273);
or U9627 (N_9627,N_7119,N_6884);
or U9628 (N_9628,N_5982,N_6653);
nor U9629 (N_9629,N_5250,N_7028);
nor U9630 (N_9630,N_6044,N_6990);
or U9631 (N_9631,N_5382,N_7246);
nor U9632 (N_9632,N_6073,N_6306);
or U9633 (N_9633,N_5859,N_5507);
nor U9634 (N_9634,N_7356,N_7392);
or U9635 (N_9635,N_7380,N_6040);
nand U9636 (N_9636,N_7443,N_6324);
xnor U9637 (N_9637,N_6305,N_5880);
and U9638 (N_9638,N_7256,N_6237);
nand U9639 (N_9639,N_6931,N_6772);
or U9640 (N_9640,N_6103,N_5823);
nor U9641 (N_9641,N_7122,N_6252);
nor U9642 (N_9642,N_6018,N_6109);
nand U9643 (N_9643,N_7199,N_6789);
or U9644 (N_9644,N_6684,N_6408);
nand U9645 (N_9645,N_6737,N_7192);
nand U9646 (N_9646,N_5968,N_5049);
and U9647 (N_9647,N_6494,N_5224);
or U9648 (N_9648,N_7026,N_5206);
or U9649 (N_9649,N_7385,N_5936);
nor U9650 (N_9650,N_6471,N_5345);
or U9651 (N_9651,N_5087,N_6497);
nand U9652 (N_9652,N_7316,N_6099);
or U9653 (N_9653,N_5241,N_7111);
nor U9654 (N_9654,N_5644,N_7009);
or U9655 (N_9655,N_6264,N_5212);
nand U9656 (N_9656,N_6815,N_6759);
nand U9657 (N_9657,N_7424,N_6380);
nor U9658 (N_9658,N_5417,N_6620);
nor U9659 (N_9659,N_6082,N_5819);
and U9660 (N_9660,N_6441,N_5738);
and U9661 (N_9661,N_5625,N_5199);
nand U9662 (N_9662,N_5577,N_5224);
nand U9663 (N_9663,N_7101,N_5193);
or U9664 (N_9664,N_5479,N_7136);
nor U9665 (N_9665,N_6822,N_5183);
or U9666 (N_9666,N_7267,N_7357);
nor U9667 (N_9667,N_6738,N_5980);
or U9668 (N_9668,N_6626,N_7051);
nand U9669 (N_9669,N_6871,N_6611);
nor U9670 (N_9670,N_5287,N_5861);
or U9671 (N_9671,N_6237,N_5369);
nor U9672 (N_9672,N_7481,N_5785);
and U9673 (N_9673,N_5055,N_5285);
nand U9674 (N_9674,N_5745,N_5036);
or U9675 (N_9675,N_5842,N_5445);
nor U9676 (N_9676,N_6445,N_6951);
and U9677 (N_9677,N_5462,N_7244);
and U9678 (N_9678,N_5386,N_5763);
nand U9679 (N_9679,N_7267,N_7332);
nor U9680 (N_9680,N_6156,N_6076);
nor U9681 (N_9681,N_5673,N_5321);
and U9682 (N_9682,N_5924,N_5402);
nand U9683 (N_9683,N_6474,N_5265);
nor U9684 (N_9684,N_5549,N_5708);
and U9685 (N_9685,N_5424,N_6390);
nand U9686 (N_9686,N_5857,N_5793);
nand U9687 (N_9687,N_5555,N_5580);
and U9688 (N_9688,N_5926,N_5999);
nor U9689 (N_9689,N_6983,N_5029);
nor U9690 (N_9690,N_5134,N_6912);
nor U9691 (N_9691,N_5923,N_5746);
and U9692 (N_9692,N_5508,N_7238);
or U9693 (N_9693,N_6526,N_5282);
nor U9694 (N_9694,N_6597,N_6911);
nor U9695 (N_9695,N_6263,N_6644);
nor U9696 (N_9696,N_5225,N_7399);
or U9697 (N_9697,N_5105,N_5250);
and U9698 (N_9698,N_5460,N_6033);
nor U9699 (N_9699,N_5146,N_6906);
and U9700 (N_9700,N_6846,N_6579);
or U9701 (N_9701,N_5691,N_6959);
nand U9702 (N_9702,N_6027,N_6076);
or U9703 (N_9703,N_6058,N_5199);
and U9704 (N_9704,N_5706,N_5801);
or U9705 (N_9705,N_6735,N_6436);
nor U9706 (N_9706,N_6830,N_6666);
or U9707 (N_9707,N_5678,N_6985);
nand U9708 (N_9708,N_6027,N_7485);
nor U9709 (N_9709,N_7118,N_5034);
nor U9710 (N_9710,N_5668,N_7428);
or U9711 (N_9711,N_5124,N_5903);
xor U9712 (N_9712,N_6464,N_7016);
or U9713 (N_9713,N_5352,N_6146);
xor U9714 (N_9714,N_5608,N_5362);
nand U9715 (N_9715,N_6775,N_6529);
nand U9716 (N_9716,N_5474,N_6999);
or U9717 (N_9717,N_7217,N_5653);
and U9718 (N_9718,N_5139,N_7001);
xor U9719 (N_9719,N_6903,N_5227);
and U9720 (N_9720,N_6919,N_6930);
and U9721 (N_9721,N_6399,N_5680);
or U9722 (N_9722,N_5487,N_5879);
nand U9723 (N_9723,N_5326,N_5844);
or U9724 (N_9724,N_5787,N_6109);
and U9725 (N_9725,N_5723,N_7263);
nand U9726 (N_9726,N_6803,N_5940);
nor U9727 (N_9727,N_5899,N_6842);
nand U9728 (N_9728,N_6317,N_6679);
and U9729 (N_9729,N_6995,N_6907);
nand U9730 (N_9730,N_5816,N_5515);
nand U9731 (N_9731,N_5856,N_6985);
and U9732 (N_9732,N_5413,N_5354);
nand U9733 (N_9733,N_7242,N_5916);
and U9734 (N_9734,N_5277,N_5951);
nand U9735 (N_9735,N_6393,N_5574);
nand U9736 (N_9736,N_5881,N_7038);
or U9737 (N_9737,N_5698,N_7039);
nand U9738 (N_9738,N_6337,N_6044);
or U9739 (N_9739,N_6938,N_7414);
and U9740 (N_9740,N_5728,N_6136);
xnor U9741 (N_9741,N_7237,N_7138);
and U9742 (N_9742,N_6148,N_6999);
and U9743 (N_9743,N_6179,N_6682);
and U9744 (N_9744,N_6013,N_5324);
and U9745 (N_9745,N_5236,N_6479);
or U9746 (N_9746,N_5044,N_7472);
nor U9747 (N_9747,N_5968,N_7118);
nor U9748 (N_9748,N_5176,N_7028);
nor U9749 (N_9749,N_5516,N_5526);
or U9750 (N_9750,N_6802,N_5909);
nor U9751 (N_9751,N_5694,N_6167);
nand U9752 (N_9752,N_5877,N_5252);
and U9753 (N_9753,N_5332,N_5794);
nand U9754 (N_9754,N_6108,N_5464);
nor U9755 (N_9755,N_7465,N_7295);
nor U9756 (N_9756,N_7307,N_5948);
or U9757 (N_9757,N_7075,N_6948);
and U9758 (N_9758,N_7162,N_5980);
or U9759 (N_9759,N_6068,N_6445);
nor U9760 (N_9760,N_6282,N_7044);
nand U9761 (N_9761,N_5344,N_7052);
nand U9762 (N_9762,N_5518,N_5884);
or U9763 (N_9763,N_6511,N_5505);
nor U9764 (N_9764,N_6497,N_5186);
and U9765 (N_9765,N_7023,N_5057);
nand U9766 (N_9766,N_6347,N_6508);
nor U9767 (N_9767,N_6839,N_6489);
nand U9768 (N_9768,N_7400,N_5949);
nand U9769 (N_9769,N_5490,N_6250);
and U9770 (N_9770,N_5813,N_5029);
nor U9771 (N_9771,N_7133,N_6157);
and U9772 (N_9772,N_5750,N_7325);
nor U9773 (N_9773,N_5255,N_5411);
or U9774 (N_9774,N_5060,N_5302);
nand U9775 (N_9775,N_7115,N_6168);
nand U9776 (N_9776,N_7409,N_6680);
or U9777 (N_9777,N_6228,N_7105);
nand U9778 (N_9778,N_7222,N_6129);
nor U9779 (N_9779,N_5177,N_5626);
nand U9780 (N_9780,N_7480,N_5022);
nand U9781 (N_9781,N_6282,N_5067);
nor U9782 (N_9782,N_6110,N_6506);
or U9783 (N_9783,N_7085,N_6465);
nand U9784 (N_9784,N_5259,N_5098);
xor U9785 (N_9785,N_6533,N_5579);
nand U9786 (N_9786,N_7484,N_7355);
or U9787 (N_9787,N_7375,N_6181);
nor U9788 (N_9788,N_5985,N_6776);
or U9789 (N_9789,N_5168,N_6729);
and U9790 (N_9790,N_6491,N_5926);
and U9791 (N_9791,N_6904,N_5870);
nand U9792 (N_9792,N_5505,N_6025);
nand U9793 (N_9793,N_6088,N_6316);
and U9794 (N_9794,N_5848,N_7183);
or U9795 (N_9795,N_5855,N_5075);
or U9796 (N_9796,N_5640,N_6669);
nor U9797 (N_9797,N_5547,N_7146);
or U9798 (N_9798,N_6281,N_7468);
or U9799 (N_9799,N_6712,N_5783);
nand U9800 (N_9800,N_5243,N_6131);
or U9801 (N_9801,N_6041,N_6856);
nor U9802 (N_9802,N_6993,N_6213);
nor U9803 (N_9803,N_7332,N_6311);
and U9804 (N_9804,N_6329,N_6916);
nor U9805 (N_9805,N_6845,N_6785);
nand U9806 (N_9806,N_6055,N_5824);
nand U9807 (N_9807,N_6317,N_6799);
xor U9808 (N_9808,N_5069,N_6938);
or U9809 (N_9809,N_6461,N_7108);
and U9810 (N_9810,N_5700,N_6513);
and U9811 (N_9811,N_6003,N_6014);
or U9812 (N_9812,N_5153,N_5215);
nor U9813 (N_9813,N_5835,N_7089);
nand U9814 (N_9814,N_5563,N_7140);
and U9815 (N_9815,N_6852,N_7286);
nand U9816 (N_9816,N_5833,N_5234);
or U9817 (N_9817,N_6101,N_5774);
or U9818 (N_9818,N_5895,N_5812);
or U9819 (N_9819,N_5922,N_6388);
or U9820 (N_9820,N_7413,N_7031);
or U9821 (N_9821,N_6284,N_6186);
nand U9822 (N_9822,N_6782,N_5751);
or U9823 (N_9823,N_6664,N_6558);
nor U9824 (N_9824,N_6471,N_5383);
nand U9825 (N_9825,N_5084,N_7286);
or U9826 (N_9826,N_5163,N_5234);
and U9827 (N_9827,N_6143,N_5271);
nand U9828 (N_9828,N_6665,N_6360);
and U9829 (N_9829,N_6755,N_5220);
or U9830 (N_9830,N_7339,N_7158);
nand U9831 (N_9831,N_6593,N_5354);
xnor U9832 (N_9832,N_5147,N_6349);
nand U9833 (N_9833,N_5654,N_5540);
nand U9834 (N_9834,N_6320,N_6292);
or U9835 (N_9835,N_5207,N_6982);
nand U9836 (N_9836,N_6660,N_5608);
nor U9837 (N_9837,N_7239,N_5931);
nand U9838 (N_9838,N_6403,N_7377);
or U9839 (N_9839,N_5729,N_6430);
nor U9840 (N_9840,N_5198,N_6013);
nor U9841 (N_9841,N_5452,N_6217);
nor U9842 (N_9842,N_5495,N_7373);
and U9843 (N_9843,N_5487,N_7086);
or U9844 (N_9844,N_6316,N_7070);
nor U9845 (N_9845,N_5268,N_6724);
nor U9846 (N_9846,N_6251,N_7035);
or U9847 (N_9847,N_5379,N_6952);
nor U9848 (N_9848,N_6547,N_5574);
nor U9849 (N_9849,N_5408,N_6056);
or U9850 (N_9850,N_5857,N_6613);
nand U9851 (N_9851,N_7328,N_7065);
nand U9852 (N_9852,N_7206,N_5395);
and U9853 (N_9853,N_7418,N_5870);
or U9854 (N_9854,N_6486,N_5404);
and U9855 (N_9855,N_7220,N_5495);
or U9856 (N_9856,N_5592,N_6519);
or U9857 (N_9857,N_7361,N_7023);
and U9858 (N_9858,N_6614,N_6556);
nand U9859 (N_9859,N_5543,N_5440);
nor U9860 (N_9860,N_6553,N_6439);
nand U9861 (N_9861,N_5422,N_5618);
and U9862 (N_9862,N_6195,N_7415);
xnor U9863 (N_9863,N_6721,N_7300);
or U9864 (N_9864,N_5821,N_7122);
nand U9865 (N_9865,N_6475,N_7434);
and U9866 (N_9866,N_5628,N_6695);
and U9867 (N_9867,N_6704,N_7075);
nand U9868 (N_9868,N_6956,N_5237);
or U9869 (N_9869,N_5410,N_6204);
and U9870 (N_9870,N_6620,N_6542);
or U9871 (N_9871,N_6892,N_5918);
nor U9872 (N_9872,N_6080,N_5594);
or U9873 (N_9873,N_7067,N_5932);
nor U9874 (N_9874,N_6156,N_6207);
or U9875 (N_9875,N_5851,N_6326);
or U9876 (N_9876,N_5784,N_5989);
or U9877 (N_9877,N_6185,N_7420);
nand U9878 (N_9878,N_6900,N_6814);
nor U9879 (N_9879,N_6946,N_7055);
or U9880 (N_9880,N_6462,N_5944);
nand U9881 (N_9881,N_5177,N_6311);
nor U9882 (N_9882,N_5698,N_6421);
or U9883 (N_9883,N_7146,N_6683);
and U9884 (N_9884,N_5906,N_6987);
and U9885 (N_9885,N_5318,N_5621);
nand U9886 (N_9886,N_5327,N_5650);
nand U9887 (N_9887,N_6115,N_6797);
xor U9888 (N_9888,N_5832,N_5151);
or U9889 (N_9889,N_5009,N_7112);
nand U9890 (N_9890,N_6604,N_7170);
nand U9891 (N_9891,N_7403,N_5911);
nand U9892 (N_9892,N_7451,N_5042);
nand U9893 (N_9893,N_6636,N_5485);
nand U9894 (N_9894,N_5119,N_6449);
and U9895 (N_9895,N_5090,N_6790);
and U9896 (N_9896,N_7182,N_6266);
nand U9897 (N_9897,N_5711,N_6110);
or U9898 (N_9898,N_5042,N_5755);
or U9899 (N_9899,N_6060,N_5595);
and U9900 (N_9900,N_5864,N_7295);
nand U9901 (N_9901,N_6041,N_6332);
nor U9902 (N_9902,N_5003,N_6009);
nor U9903 (N_9903,N_5942,N_6753);
nand U9904 (N_9904,N_6727,N_7474);
nor U9905 (N_9905,N_7080,N_6958);
or U9906 (N_9906,N_5945,N_6541);
or U9907 (N_9907,N_5127,N_6495);
and U9908 (N_9908,N_7199,N_7392);
nand U9909 (N_9909,N_6626,N_6539);
nor U9910 (N_9910,N_5198,N_6964);
or U9911 (N_9911,N_6948,N_6557);
or U9912 (N_9912,N_7332,N_7004);
or U9913 (N_9913,N_6303,N_6554);
and U9914 (N_9914,N_7298,N_5683);
or U9915 (N_9915,N_6143,N_5715);
nor U9916 (N_9916,N_7141,N_6819);
and U9917 (N_9917,N_6745,N_6097);
nand U9918 (N_9918,N_6759,N_6972);
nor U9919 (N_9919,N_6649,N_6551);
nand U9920 (N_9920,N_5170,N_6568);
and U9921 (N_9921,N_6856,N_5834);
and U9922 (N_9922,N_5419,N_6591);
or U9923 (N_9923,N_6621,N_6350);
and U9924 (N_9924,N_5662,N_7322);
and U9925 (N_9925,N_5933,N_5595);
nor U9926 (N_9926,N_5069,N_6857);
and U9927 (N_9927,N_5189,N_6280);
and U9928 (N_9928,N_6453,N_6751);
or U9929 (N_9929,N_6107,N_6269);
nor U9930 (N_9930,N_5998,N_5248);
and U9931 (N_9931,N_5411,N_5923);
and U9932 (N_9932,N_7072,N_6825);
and U9933 (N_9933,N_6540,N_6663);
nor U9934 (N_9934,N_7027,N_5790);
nor U9935 (N_9935,N_6742,N_7029);
nor U9936 (N_9936,N_5154,N_7368);
or U9937 (N_9937,N_5015,N_5072);
nand U9938 (N_9938,N_6666,N_6816);
or U9939 (N_9939,N_6565,N_5492);
nor U9940 (N_9940,N_5025,N_7202);
nor U9941 (N_9941,N_6737,N_5163);
and U9942 (N_9942,N_6871,N_7300);
nor U9943 (N_9943,N_6795,N_6423);
and U9944 (N_9944,N_7244,N_7076);
and U9945 (N_9945,N_6734,N_7078);
nand U9946 (N_9946,N_5203,N_6438);
and U9947 (N_9947,N_6184,N_5209);
nor U9948 (N_9948,N_5390,N_5218);
nand U9949 (N_9949,N_6528,N_6208);
or U9950 (N_9950,N_5850,N_6832);
nand U9951 (N_9951,N_5081,N_6659);
nand U9952 (N_9952,N_6111,N_7389);
nand U9953 (N_9953,N_6383,N_6196);
nand U9954 (N_9954,N_5083,N_6292);
and U9955 (N_9955,N_5877,N_5130);
xnor U9956 (N_9956,N_6020,N_6988);
and U9957 (N_9957,N_7367,N_7472);
and U9958 (N_9958,N_6218,N_6289);
nand U9959 (N_9959,N_5225,N_7138);
nand U9960 (N_9960,N_6210,N_6882);
nor U9961 (N_9961,N_6320,N_6728);
nor U9962 (N_9962,N_6967,N_5772);
and U9963 (N_9963,N_6611,N_5086);
or U9964 (N_9964,N_5061,N_5236);
or U9965 (N_9965,N_6934,N_5805);
and U9966 (N_9966,N_6415,N_7262);
nor U9967 (N_9967,N_5608,N_6803);
or U9968 (N_9968,N_7377,N_5943);
or U9969 (N_9969,N_5559,N_7092);
and U9970 (N_9970,N_5000,N_6238);
or U9971 (N_9971,N_5848,N_5003);
and U9972 (N_9972,N_5902,N_6096);
xnor U9973 (N_9973,N_7395,N_5919);
nand U9974 (N_9974,N_7479,N_6594);
or U9975 (N_9975,N_7439,N_6969);
or U9976 (N_9976,N_5582,N_5611);
and U9977 (N_9977,N_5722,N_7208);
and U9978 (N_9978,N_6389,N_6434);
or U9979 (N_9979,N_7425,N_7316);
and U9980 (N_9980,N_6079,N_5753);
nor U9981 (N_9981,N_6824,N_6451);
nand U9982 (N_9982,N_6964,N_5140);
nand U9983 (N_9983,N_5270,N_7081);
or U9984 (N_9984,N_5439,N_6242);
and U9985 (N_9985,N_5384,N_5339);
nor U9986 (N_9986,N_7127,N_7370);
nand U9987 (N_9987,N_5918,N_6564);
nor U9988 (N_9988,N_5611,N_7122);
nor U9989 (N_9989,N_6642,N_7105);
and U9990 (N_9990,N_6156,N_7184);
nor U9991 (N_9991,N_5999,N_6096);
xor U9992 (N_9992,N_6152,N_7079);
and U9993 (N_9993,N_6819,N_6382);
or U9994 (N_9994,N_7150,N_6223);
or U9995 (N_9995,N_7023,N_7228);
and U9996 (N_9996,N_5378,N_5238);
or U9997 (N_9997,N_5511,N_5762);
nor U9998 (N_9998,N_6358,N_6605);
nor U9999 (N_9999,N_5041,N_5487);
nor UO_0 (O_0,N_8564,N_9401);
and UO_1 (O_1,N_8392,N_7511);
nand UO_2 (O_2,N_7783,N_7991);
or UO_3 (O_3,N_7774,N_8165);
and UO_4 (O_4,N_9266,N_8590);
and UO_5 (O_5,N_9173,N_8602);
or UO_6 (O_6,N_8479,N_8049);
nand UO_7 (O_7,N_8523,N_9952);
nand UO_8 (O_8,N_8976,N_9199);
or UO_9 (O_9,N_8474,N_8865);
or UO_10 (O_10,N_9544,N_9295);
nand UO_11 (O_11,N_8438,N_8414);
or UO_12 (O_12,N_9884,N_9965);
nor UO_13 (O_13,N_9851,N_9862);
nand UO_14 (O_14,N_9506,N_8265);
nor UO_15 (O_15,N_9435,N_7943);
and UO_16 (O_16,N_9793,N_8686);
nand UO_17 (O_17,N_8561,N_7916);
nor UO_18 (O_18,N_8021,N_8399);
nor UO_19 (O_19,N_7917,N_9584);
and UO_20 (O_20,N_7900,N_9445);
and UO_21 (O_21,N_7575,N_8897);
or UO_22 (O_22,N_8596,N_9852);
and UO_23 (O_23,N_7849,N_7524);
nor UO_24 (O_24,N_9135,N_8948);
nor UO_25 (O_25,N_8762,N_9707);
and UO_26 (O_26,N_8396,N_7997);
and UO_27 (O_27,N_9321,N_8237);
xnor UO_28 (O_28,N_9896,N_8988);
or UO_29 (O_29,N_7519,N_7821);
nor UO_30 (O_30,N_9616,N_8943);
or UO_31 (O_31,N_8017,N_9123);
or UO_32 (O_32,N_8133,N_9557);
and UO_33 (O_33,N_8428,N_7859);
or UO_34 (O_34,N_9715,N_8725);
or UO_35 (O_35,N_8683,N_9479);
or UO_36 (O_36,N_8589,N_9861);
and UO_37 (O_37,N_9450,N_8741);
and UO_38 (O_38,N_9685,N_9904);
xor UO_39 (O_39,N_9358,N_7583);
nor UO_40 (O_40,N_8199,N_8455);
nor UO_41 (O_41,N_9976,N_7853);
or UO_42 (O_42,N_8168,N_9193);
nand UO_43 (O_43,N_8170,N_9430);
nor UO_44 (O_44,N_7970,N_9386);
and UO_45 (O_45,N_9697,N_8851);
and UO_46 (O_46,N_7792,N_8166);
nand UO_47 (O_47,N_9877,N_9227);
or UO_48 (O_48,N_8158,N_7995);
or UO_49 (O_49,N_9624,N_9818);
nor UO_50 (O_50,N_9836,N_8185);
nor UO_51 (O_51,N_8978,N_8633);
nor UO_52 (O_52,N_7981,N_9819);
nand UO_53 (O_53,N_8912,N_9252);
nand UO_54 (O_54,N_8294,N_9675);
and UO_55 (O_55,N_8664,N_7504);
nor UO_56 (O_56,N_9301,N_9639);
and UO_57 (O_57,N_9421,N_7617);
nand UO_58 (O_58,N_9592,N_8124);
nand UO_59 (O_59,N_9567,N_9731);
or UO_60 (O_60,N_8630,N_8097);
nand UO_61 (O_61,N_8003,N_9935);
nand UO_62 (O_62,N_9413,N_9814);
nand UO_63 (O_63,N_8347,N_9628);
and UO_64 (O_64,N_9765,N_7579);
nand UO_65 (O_65,N_9171,N_9408);
nand UO_66 (O_66,N_9810,N_9000);
and UO_67 (O_67,N_8586,N_8763);
or UO_68 (O_68,N_8526,N_8736);
or UO_69 (O_69,N_9328,N_8768);
nor UO_70 (O_70,N_8844,N_8252);
and UO_71 (O_71,N_9237,N_8351);
and UO_72 (O_72,N_9929,N_7702);
and UO_73 (O_73,N_8814,N_9642);
nor UO_74 (O_74,N_9327,N_8323);
nor UO_75 (O_75,N_7542,N_9322);
and UO_76 (O_76,N_8301,N_8466);
or UO_77 (O_77,N_9342,N_7957);
or UO_78 (O_78,N_7962,N_7503);
xnor UO_79 (O_79,N_9086,N_7666);
and UO_80 (O_80,N_8211,N_9293);
nand UO_81 (O_81,N_9615,N_9687);
nand UO_82 (O_82,N_8179,N_9478);
nand UO_83 (O_83,N_8924,N_7967);
nor UO_84 (O_84,N_8416,N_8288);
nand UO_85 (O_85,N_8436,N_7982);
nor UO_86 (O_86,N_8385,N_8061);
nand UO_87 (O_87,N_7836,N_9238);
nand UO_88 (O_88,N_8092,N_8950);
nor UO_89 (O_89,N_8853,N_9329);
and UO_90 (O_90,N_8813,N_9243);
and UO_91 (O_91,N_8189,N_8531);
nand UO_92 (O_92,N_9739,N_8108);
or UO_93 (O_93,N_9525,N_8473);
nand UO_94 (O_94,N_7866,N_7825);
nand UO_95 (O_95,N_7685,N_7614);
or UO_96 (O_96,N_8908,N_7551);
nand UO_97 (O_97,N_9411,N_9370);
nor UO_98 (O_98,N_9859,N_8171);
and UO_99 (O_99,N_8841,N_8256);
or UO_100 (O_100,N_8666,N_8553);
nand UO_101 (O_101,N_8462,N_8842);
and UO_102 (O_102,N_9931,N_7518);
and UO_103 (O_103,N_9597,N_8148);
or UO_104 (O_104,N_8742,N_7740);
and UO_105 (O_105,N_9688,N_9234);
nor UO_106 (O_106,N_8577,N_9829);
xnor UO_107 (O_107,N_9847,N_9082);
nand UO_108 (O_108,N_9735,N_9283);
and UO_109 (O_109,N_8552,N_7779);
nor UO_110 (O_110,N_9728,N_9477);
and UO_111 (O_111,N_9330,N_9660);
nor UO_112 (O_112,N_9442,N_8492);
and UO_113 (O_113,N_9871,N_9941);
and UO_114 (O_114,N_8491,N_9451);
or UO_115 (O_115,N_9088,N_7677);
nand UO_116 (O_116,N_8270,N_9657);
and UO_117 (O_117,N_8753,N_9311);
or UO_118 (O_118,N_8793,N_8091);
or UO_119 (O_119,N_7892,N_8063);
nand UO_120 (O_120,N_7985,N_8386);
or UO_121 (O_121,N_8443,N_9111);
and UO_122 (O_122,N_7976,N_8595);
nor UO_123 (O_123,N_9602,N_9343);
nor UO_124 (O_124,N_8981,N_9133);
and UO_125 (O_125,N_8556,N_9956);
or UO_126 (O_126,N_8891,N_7824);
or UO_127 (O_127,N_9107,N_8144);
or UO_128 (O_128,N_9629,N_9215);
nand UO_129 (O_129,N_8638,N_7840);
or UO_130 (O_130,N_8790,N_8373);
nand UO_131 (O_131,N_7545,N_8919);
nor UO_132 (O_132,N_9394,N_9800);
nor UO_133 (O_133,N_9940,N_9932);
nor UO_134 (O_134,N_8224,N_9471);
or UO_135 (O_135,N_7506,N_8073);
or UO_136 (O_136,N_9744,N_8041);
nand UO_137 (O_137,N_8248,N_9348);
nor UO_138 (O_138,N_9963,N_7777);
nand UO_139 (O_139,N_8990,N_7785);
nand UO_140 (O_140,N_9975,N_8051);
nand UO_141 (O_141,N_8212,N_8974);
or UO_142 (O_142,N_9103,N_8751);
nand UO_143 (O_143,N_9604,N_8054);
or UO_144 (O_144,N_8606,N_9038);
nand UO_145 (O_145,N_9794,N_7746);
nand UO_146 (O_146,N_7901,N_8783);
nand UO_147 (O_147,N_7771,N_9520);
nand UO_148 (O_148,N_9574,N_7915);
and UO_149 (O_149,N_7910,N_9019);
and UO_150 (O_150,N_7532,N_9489);
nand UO_151 (O_151,N_9369,N_8805);
or UO_152 (O_152,N_8951,N_8567);
and UO_153 (O_153,N_7974,N_9811);
or UO_154 (O_154,N_8952,N_7797);
and UO_155 (O_155,N_9446,N_9198);
nor UO_156 (O_156,N_8264,N_8417);
nor UO_157 (O_157,N_9864,N_8314);
nor UO_158 (O_158,N_8501,N_8230);
nand UO_159 (O_159,N_8758,N_9101);
and UO_160 (O_160,N_7730,N_9955);
nand UO_161 (O_161,N_8057,N_9580);
nand UO_162 (O_162,N_9326,N_8512);
xor UO_163 (O_163,N_9878,N_8111);
nor UO_164 (O_164,N_8784,N_9235);
or UO_165 (O_165,N_9049,N_8617);
nor UO_166 (O_166,N_9319,N_9143);
nor UO_167 (O_167,N_9412,N_8538);
or UO_168 (O_168,N_9880,N_8184);
and UO_169 (O_169,N_9159,N_9933);
nor UO_170 (O_170,N_8127,N_9732);
and UO_171 (O_171,N_8076,N_9384);
or UO_172 (O_172,N_9536,N_9080);
nand UO_173 (O_173,N_8773,N_7869);
and UO_174 (O_174,N_9559,N_8801);
nand UO_175 (O_175,N_9516,N_7927);
xnor UO_176 (O_176,N_9959,N_9913);
nand UO_177 (O_177,N_8706,N_9673);
nand UO_178 (O_178,N_8651,N_8328);
or UO_179 (O_179,N_9434,N_9346);
or UO_180 (O_180,N_8223,N_8113);
or UO_181 (O_181,N_8046,N_8478);
and UO_182 (O_182,N_8828,N_8957);
and UO_183 (O_183,N_9226,N_7599);
nor UO_184 (O_184,N_9149,N_9946);
and UO_185 (O_185,N_8870,N_7500);
nor UO_186 (O_186,N_8695,N_8746);
and UO_187 (O_187,N_9883,N_9265);
nand UO_188 (O_188,N_9296,N_9930);
and UO_189 (O_189,N_9891,N_7736);
nand UO_190 (O_190,N_9982,N_9014);
xnor UO_191 (O_191,N_8283,N_8599);
nor UO_192 (O_192,N_9449,N_8321);
nor UO_193 (O_193,N_9182,N_9834);
nand UO_194 (O_194,N_8818,N_8662);
and UO_195 (O_195,N_8581,N_9591);
and UO_196 (O_196,N_8145,N_9908);
and UO_197 (O_197,N_7589,N_8542);
xnor UO_198 (O_198,N_8447,N_8835);
nor UO_199 (O_199,N_7906,N_8259);
and UO_200 (O_200,N_7793,N_7944);
or UO_201 (O_201,N_9514,N_7939);
and UO_202 (O_202,N_8527,N_9548);
nor UO_203 (O_203,N_8900,N_8286);
nor UO_204 (O_204,N_9254,N_9417);
and UO_205 (O_205,N_8667,N_7674);
nand UO_206 (O_206,N_8302,N_9665);
nand UO_207 (O_207,N_7555,N_8047);
or UO_208 (O_208,N_7582,N_8193);
or UO_209 (O_209,N_9705,N_8937);
nor UO_210 (O_210,N_9826,N_9132);
xor UO_211 (O_211,N_7585,N_8500);
nand UO_212 (O_212,N_8739,N_9773);
and UO_213 (O_213,N_9058,N_7652);
and UO_214 (O_214,N_8954,N_8597);
and UO_215 (O_215,N_9969,N_8487);
nor UO_216 (O_216,N_7822,N_8713);
nand UO_217 (O_217,N_8050,N_7856);
and UO_218 (O_218,N_7880,N_7592);
nor UO_219 (O_219,N_9331,N_8499);
nor UO_220 (O_220,N_9183,N_8112);
or UO_221 (O_221,N_8128,N_9870);
and UO_222 (O_222,N_8454,N_8044);
and UO_223 (O_223,N_8291,N_8456);
or UO_224 (O_224,N_8559,N_9024);
nand UO_225 (O_225,N_7665,N_8820);
and UO_226 (O_226,N_8761,N_8536);
nand UO_227 (O_227,N_8665,N_9611);
or UO_228 (O_228,N_8977,N_7828);
or UO_229 (O_229,N_8293,N_8955);
nor UO_230 (O_230,N_7660,N_9169);
nand UO_231 (O_231,N_7854,N_8240);
and UO_232 (O_232,N_9483,N_8135);
or UO_233 (O_233,N_8378,N_8837);
nand UO_234 (O_234,N_8432,N_8513);
nand UO_235 (O_235,N_9512,N_8102);
nor UO_236 (O_236,N_8635,N_7903);
xor UO_237 (O_237,N_7933,N_9120);
or UO_238 (O_238,N_9919,N_7775);
or UO_239 (O_239,N_9422,N_8172);
or UO_240 (O_240,N_8023,N_7725);
and UO_241 (O_241,N_7656,N_9906);
and UO_242 (O_242,N_7514,N_9363);
xnor UO_243 (O_243,N_8752,N_9129);
and UO_244 (O_244,N_9733,N_8772);
and UO_245 (O_245,N_8922,N_9162);
or UO_246 (O_246,N_7929,N_9555);
and UO_247 (O_247,N_9911,N_8352);
or UO_248 (O_248,N_9991,N_7923);
nand UO_249 (O_249,N_8575,N_8963);
nand UO_250 (O_250,N_9569,N_7513);
or UO_251 (O_251,N_9798,N_9703);
and UO_252 (O_252,N_9858,N_7966);
and UO_253 (O_253,N_7651,N_9889);
or UO_254 (O_254,N_9094,N_9978);
nand UO_255 (O_255,N_9897,N_9997);
and UO_256 (O_256,N_9637,N_9473);
or UO_257 (O_257,N_7881,N_7734);
nand UO_258 (O_258,N_7516,N_9281);
or UO_259 (O_259,N_9158,N_8383);
or UO_260 (O_260,N_9304,N_9404);
nor UO_261 (O_261,N_9313,N_8368);
nor UO_262 (O_262,N_8118,N_8181);
nand UO_263 (O_263,N_7826,N_8770);
nand UO_264 (O_264,N_9620,N_7591);
nand UO_265 (O_265,N_8251,N_7701);
and UO_266 (O_266,N_9560,N_7650);
xor UO_267 (O_267,N_9153,N_7558);
and UO_268 (O_268,N_9119,N_7567);
and UO_269 (O_269,N_8268,N_8940);
nor UO_270 (O_270,N_8945,N_8962);
and UO_271 (O_271,N_8439,N_7969);
nor UO_272 (O_272,N_8472,N_9087);
and UO_273 (O_273,N_9361,N_9267);
and UO_274 (O_274,N_9064,N_7517);
and UO_275 (O_275,N_7726,N_7930);
and UO_276 (O_276,N_8360,N_7619);
nand UO_277 (O_277,N_9314,N_8074);
or UO_278 (O_278,N_8696,N_9092);
and UO_279 (O_279,N_8515,N_9797);
or UO_280 (O_280,N_9831,N_8344);
and UO_281 (O_281,N_9568,N_8804);
nor UO_282 (O_282,N_8134,N_9270);
nand UO_283 (O_283,N_9184,N_9730);
or UO_284 (O_284,N_9924,N_7705);
nor UO_285 (O_285,N_8882,N_9779);
xnor UO_286 (O_286,N_8271,N_9833);
or UO_287 (O_287,N_8588,N_7681);
nor UO_288 (O_288,N_9035,N_8260);
nor UO_289 (O_289,N_9505,N_9855);
nand UO_290 (O_290,N_9306,N_8210);
or UO_291 (O_291,N_7597,N_8780);
nand UO_292 (O_292,N_8038,N_8403);
and UO_293 (O_293,N_9280,N_8522);
nor UO_294 (O_294,N_9549,N_8488);
nand UO_295 (O_295,N_9324,N_9274);
nor UO_296 (O_296,N_7834,N_8637);
and UO_297 (O_297,N_8121,N_8088);
and UO_298 (O_298,N_9668,N_8206);
or UO_299 (O_299,N_7622,N_9632);
and UO_300 (O_300,N_9890,N_9072);
and UO_301 (O_301,N_8099,N_7913);
nor UO_302 (O_302,N_7601,N_9294);
nor UO_303 (O_303,N_9144,N_9219);
and UO_304 (O_304,N_8649,N_9258);
xnor UO_305 (O_305,N_9579,N_8704);
and UO_306 (O_306,N_9200,N_9392);
or UO_307 (O_307,N_7918,N_9607);
or UO_308 (O_308,N_8546,N_8519);
and UO_309 (O_309,N_7909,N_9013);
and UO_310 (O_310,N_7898,N_7907);
and UO_311 (O_311,N_7722,N_8470);
nand UO_312 (O_312,N_9095,N_7757);
and UO_313 (O_313,N_8973,N_8390);
and UO_314 (O_314,N_7895,N_7946);
and UO_315 (O_315,N_8072,N_8678);
nand UO_316 (O_316,N_9110,N_8899);
or UO_317 (O_317,N_7507,N_8201);
nor UO_318 (O_318,N_8255,N_7573);
and UO_319 (O_319,N_8316,N_7754);
or UO_320 (O_320,N_9461,N_8530);
nor UO_321 (O_321,N_9915,N_8895);
nor UO_322 (O_322,N_8587,N_9677);
or UO_323 (O_323,N_7745,N_8132);
and UO_324 (O_324,N_9888,N_9659);
nor UO_325 (O_325,N_8312,N_7934);
or UO_326 (O_326,N_8720,N_9522);
nand UO_327 (O_327,N_8468,N_9766);
or UO_328 (O_328,N_9105,N_9106);
and UO_329 (O_329,N_9065,N_8320);
nand UO_330 (O_330,N_9586,N_7949);
nor UO_331 (O_331,N_9954,N_9601);
xor UO_332 (O_332,N_8708,N_8938);
or UO_333 (O_333,N_7586,N_9165);
nand UO_334 (O_334,N_8953,N_9373);
nand UO_335 (O_335,N_9042,N_8239);
or UO_336 (O_336,N_8202,N_7902);
nor UO_337 (O_337,N_9951,N_8180);
and UO_338 (O_338,N_8615,N_9315);
nand UO_339 (O_339,N_7543,N_8880);
nand UO_340 (O_340,N_8892,N_7813);
or UO_341 (O_341,N_8246,N_7735);
or UO_342 (O_342,N_8387,N_8009);
nor UO_343 (O_343,N_8916,N_9511);
and UO_344 (O_344,N_8430,N_8888);
nand UO_345 (O_345,N_8534,N_9748);
nor UO_346 (O_346,N_9172,N_9290);
and UO_347 (O_347,N_8086,N_9720);
nor UO_348 (O_348,N_9104,N_9509);
or UO_349 (O_349,N_8528,N_8242);
and UO_350 (O_350,N_8701,N_7887);
nand UO_351 (O_351,N_7690,N_8384);
nor UO_352 (O_352,N_9857,N_7788);
or UO_353 (O_353,N_9071,N_9581);
and UO_354 (O_354,N_8755,N_9981);
xor UO_355 (O_355,N_8100,N_7897);
and UO_356 (O_356,N_7696,N_8415);
and UO_357 (O_357,N_8004,N_9902);
nor UO_358 (O_358,N_7747,N_8558);
and UO_359 (O_359,N_8660,N_9467);
xnor UO_360 (O_360,N_8254,N_9115);
and UO_361 (O_361,N_8020,N_8109);
nor UO_362 (O_362,N_8845,N_8093);
nand UO_363 (O_363,N_7986,N_9136);
or UO_364 (O_364,N_9879,N_9070);
nor UO_365 (O_365,N_9006,N_9351);
or UO_366 (O_366,N_7875,N_9519);
nand UO_367 (O_367,N_8732,N_7996);
nor UO_368 (O_368,N_8547,N_7649);
nor UO_369 (O_369,N_9947,N_9223);
and UO_370 (O_370,N_7661,N_8327);
nand UO_371 (O_371,N_8276,N_9093);
or UO_372 (O_372,N_7721,N_9460);
and UO_373 (O_373,N_9518,N_9073);
or UO_374 (O_374,N_8213,N_9098);
or UO_375 (O_375,N_8766,N_8485);
nand UO_376 (O_376,N_7805,N_9517);
and UO_377 (O_377,N_7807,N_8715);
nor UO_378 (O_378,N_8508,N_8346);
nor UO_379 (O_379,N_8453,N_9218);
or UO_380 (O_380,N_7676,N_9145);
xor UO_381 (O_381,N_8925,N_8815);
nor UO_382 (O_382,N_7803,N_8411);
nor UO_383 (O_383,N_8568,N_7819);
nor UO_384 (O_384,N_8391,N_8656);
nor UO_385 (O_385,N_9125,N_8860);
nor UO_386 (O_386,N_8873,N_8484);
or UO_387 (O_387,N_7955,N_7609);
nand UO_388 (O_388,N_8257,N_9613);
nor UO_389 (O_389,N_9850,N_9986);
nand UO_390 (O_390,N_8449,N_8641);
and UO_391 (O_391,N_9967,N_7978);
nand UO_392 (O_392,N_8698,N_9211);
nor UO_393 (O_393,N_8303,N_8130);
nand UO_394 (O_394,N_8469,N_9026);
xnor UO_395 (O_395,N_8707,N_8410);
nand UO_396 (O_396,N_8016,N_8744);
and UO_397 (O_397,N_8819,N_8620);
and UO_398 (O_398,N_8369,N_9214);
nand UO_399 (O_399,N_9783,N_8156);
and UO_400 (O_400,N_9583,N_9843);
nor UO_401 (O_401,N_8594,N_9605);
nand UO_402 (O_402,N_8196,N_9807);
or UO_403 (O_403,N_9454,N_8238);
or UO_404 (O_404,N_8161,N_7693);
and UO_405 (O_405,N_8426,N_8343);
xnor UO_406 (O_406,N_9337,N_9790);
nor UO_407 (O_407,N_8983,N_8584);
or UO_408 (O_408,N_9029,N_8167);
nand UO_409 (O_409,N_9117,N_7637);
nand UO_410 (O_410,N_9695,N_8728);
nor UO_411 (O_411,N_9684,N_7574);
nor UO_412 (O_412,N_7863,N_8769);
and UO_413 (O_413,N_8848,N_8794);
and UO_414 (O_414,N_9085,N_8292);
and UO_415 (O_415,N_9918,N_7546);
nand UO_416 (O_416,N_8944,N_8195);
and UO_417 (O_417,N_9740,N_8674);
nor UO_418 (O_418,N_7624,N_9063);
and UO_419 (O_419,N_8176,N_8094);
and UO_420 (O_420,N_8404,N_8183);
or UO_421 (O_421,N_8636,N_8480);
nand UO_422 (O_422,N_9154,N_9815);
nand UO_423 (O_423,N_8274,N_9641);
nand UO_424 (O_424,N_7595,N_9423);
and UO_425 (O_425,N_7741,N_7928);
and UO_426 (O_426,N_9285,N_7911);
nor UO_427 (O_427,N_7889,N_9551);
xnor UO_428 (O_428,N_8947,N_9468);
xnor UO_429 (O_429,N_8825,N_8277);
nand UO_430 (O_430,N_9187,N_9067);
nand UO_431 (O_431,N_8122,N_8205);
nand UO_432 (O_432,N_8685,N_8192);
or UO_433 (O_433,N_8318,N_9868);
nand UO_434 (O_434,N_8011,N_9257);
nor UO_435 (O_435,N_8015,N_9802);
and UO_436 (O_436,N_7795,N_8863);
nand UO_437 (O_437,N_9979,N_8996);
or UO_438 (O_438,N_7936,N_9875);
nand UO_439 (O_439,N_8743,N_7862);
nand UO_440 (O_440,N_7646,N_9916);
nand UO_441 (O_441,N_8361,N_9114);
nor UO_442 (O_442,N_7522,N_8893);
or UO_443 (O_443,N_7508,N_7525);
nand UO_444 (O_444,N_8754,N_9150);
or UO_445 (O_445,N_8243,N_7694);
and UO_446 (O_446,N_8653,N_8774);
nor UO_447 (O_447,N_9163,N_8543);
nor UO_448 (O_448,N_8215,N_9335);
nand UO_449 (O_449,N_8131,N_9431);
nand UO_450 (O_450,N_8370,N_9535);
and UO_451 (O_451,N_8826,N_8616);
nand UO_452 (O_452,N_8796,N_9709);
nor UO_453 (O_453,N_7753,N_9622);
nand UO_454 (O_454,N_9533,N_7993);
xnor UO_455 (O_455,N_7852,N_9221);
nand UO_456 (O_456,N_9960,N_8476);
and UO_457 (O_457,N_9977,N_9139);
or UO_458 (O_458,N_9465,N_9312);
or UO_459 (O_459,N_8861,N_8569);
nor UO_460 (O_460,N_8281,N_9920);
and UO_461 (O_461,N_9061,N_8781);
nor UO_462 (O_462,N_8740,N_9081);
or UO_463 (O_463,N_8084,N_9475);
or UO_464 (O_464,N_9022,N_9841);
nor UO_465 (O_465,N_8961,N_7891);
and UO_466 (O_466,N_9573,N_9690);
or UO_467 (O_467,N_8997,N_9490);
nor UO_468 (O_468,N_9357,N_8855);
nor UO_469 (O_469,N_7724,N_8789);
and UO_470 (O_470,N_7844,N_9378);
or UO_471 (O_471,N_9409,N_8482);
nor UO_472 (O_472,N_7587,N_9714);
nand UO_473 (O_473,N_8363,N_9228);
or UO_474 (O_474,N_7645,N_7553);
nand UO_475 (O_475,N_8125,N_8490);
and UO_476 (O_476,N_9069,N_7748);
nor UO_477 (O_477,N_8942,N_8505);
nor UO_478 (O_478,N_9926,N_9538);
or UO_479 (O_479,N_9985,N_9962);
nor UO_480 (O_480,N_8823,N_7535);
or UO_481 (O_481,N_9663,N_9040);
and UO_482 (O_482,N_8078,N_9344);
or UO_483 (O_483,N_8450,N_9127);
nor UO_484 (O_484,N_9076,N_9900);
and UO_485 (O_485,N_9774,N_8562);
nor UO_486 (O_486,N_8064,N_8750);
or UO_487 (O_487,N_9231,N_9134);
or UO_488 (O_488,N_8854,N_9565);
or UO_489 (O_489,N_8504,N_9524);
nor UO_490 (O_490,N_9371,N_9618);
nor UO_491 (O_491,N_7893,N_9664);
or UO_492 (O_492,N_8053,N_8267);
or UO_493 (O_493,N_8036,N_9174);
or UO_494 (O_494,N_9308,N_8349);
and UO_495 (O_495,N_9131,N_7706);
nor UO_496 (O_496,N_9255,N_9742);
and UO_497 (O_497,N_8198,N_7794);
nand UO_498 (O_498,N_9694,N_9288);
nand UO_499 (O_499,N_8747,N_8779);
and UO_500 (O_500,N_9617,N_9097);
nor UO_501 (O_501,N_9661,N_8910);
and UO_502 (O_502,N_9722,N_7580);
nor UO_503 (O_503,N_7987,N_7602);
or UO_504 (O_504,N_9844,N_7615);
or UO_505 (O_505,N_7572,N_7835);
nand UO_506 (O_506,N_9074,N_7989);
nor UO_507 (O_507,N_9990,N_9575);
or UO_508 (O_508,N_9813,N_8147);
and UO_509 (O_509,N_7905,N_8310);
and UO_510 (O_510,N_8580,N_9096);
nand UO_511 (O_511,N_9746,N_8110);
or UO_512 (O_512,N_9262,N_9441);
nand UO_513 (O_513,N_9682,N_8059);
and UO_514 (O_514,N_8593,N_8164);
nand UO_515 (O_515,N_8115,N_8712);
nor UO_516 (O_516,N_7733,N_7679);
and UO_517 (O_517,N_8991,N_8724);
nor UO_518 (O_518,N_9176,N_8507);
nor UO_519 (O_519,N_8757,N_7768);
nor UO_520 (O_520,N_9151,N_9571);
or UO_521 (O_521,N_8231,N_7979);
nor UO_522 (O_522,N_7971,N_7964);
nand UO_523 (O_523,N_8668,N_7505);
nor UO_524 (O_524,N_8304,N_7922);
or UO_525 (O_525,N_9124,N_9667);
or UO_526 (O_526,N_8611,N_8759);
xor UO_527 (O_527,N_8463,N_8669);
nand UO_528 (O_528,N_9658,N_8300);
or UO_529 (O_529,N_9041,N_7699);
or UO_530 (O_530,N_9084,N_9300);
nor UO_531 (O_531,N_8871,N_7743);
or UO_532 (O_532,N_9492,N_8075);
xor UO_533 (O_533,N_8833,N_8080);
or UO_534 (O_534,N_8266,N_8337);
and UO_535 (O_535,N_9636,N_8623);
or UO_536 (O_536,N_9588,N_8000);
and UO_537 (O_537,N_8726,N_9068);
nor UO_538 (O_538,N_8603,N_7556);
or UO_539 (O_539,N_9164,N_8776);
nor UO_540 (O_540,N_8735,N_9222);
nor UO_541 (O_541,N_9273,N_8037);
nor UO_542 (O_542,N_9246,N_9768);
nand UO_543 (O_543,N_9718,N_8083);
and UO_544 (O_544,N_7596,N_7628);
and UO_545 (O_545,N_9700,N_9398);
nand UO_546 (O_546,N_7564,N_9502);
nor UO_547 (O_547,N_7620,N_9083);
nor UO_548 (O_548,N_8245,N_7719);
xor UO_549 (O_549,N_8077,N_8809);
or UO_550 (O_550,N_8889,N_7621);
nor UO_551 (O_551,N_9034,N_9470);
nor UO_552 (O_552,N_8186,N_8433);
nand UO_553 (O_553,N_8290,N_9118);
or UO_554 (O_554,N_9100,N_8035);
nor UO_555 (O_555,N_7631,N_9152);
or UO_556 (O_556,N_8070,N_9747);
or UO_557 (O_557,N_7780,N_7626);
or UO_558 (O_558,N_8672,N_8029);
and UO_559 (O_559,N_8413,N_8688);
xor UO_560 (O_560,N_9830,N_9835);
nor UO_561 (O_561,N_8297,N_7695);
nand UO_562 (O_562,N_9554,N_9474);
and UO_563 (O_563,N_7765,N_9874);
or UO_564 (O_564,N_8548,N_8631);
or UO_565 (O_565,N_8901,N_9113);
or UO_566 (O_566,N_9380,N_8217);
nand UO_567 (O_567,N_8442,N_9418);
nand UO_568 (O_568,N_7501,N_9448);
nand UO_569 (O_569,N_8503,N_9846);
or UO_570 (O_570,N_9432,N_7715);
nand UO_571 (O_571,N_9692,N_9156);
nor UO_572 (O_572,N_8225,N_9427);
or UO_573 (O_573,N_8541,N_7636);
or UO_574 (O_574,N_9599,N_7827);
or UO_575 (O_575,N_9276,N_9775);
xor UO_576 (O_576,N_8279,N_7616);
nand UO_577 (O_577,N_9012,N_8493);
nor UO_578 (O_578,N_8560,N_7940);
or UO_579 (O_579,N_9680,N_8516);
nand UO_580 (O_580,N_8307,N_8169);
or UO_581 (O_581,N_8388,N_7723);
nand UO_582 (O_582,N_7576,N_7712);
nand UO_583 (O_583,N_8345,N_8788);
nor UO_584 (O_584,N_8014,N_7919);
or UO_585 (O_585,N_8218,N_8898);
nand UO_586 (O_586,N_9403,N_9712);
or UO_587 (O_587,N_8545,N_9181);
nand UO_588 (O_588,N_9318,N_9876);
and UO_589 (O_589,N_9625,N_9056);
or UO_590 (O_590,N_9202,N_7557);
nand UO_591 (O_591,N_9698,N_9964);
nand UO_592 (O_592,N_7662,N_9501);
nor UO_593 (O_593,N_7659,N_9832);
nand UO_594 (O_594,N_8601,N_7547);
or UO_595 (O_595,N_9972,N_8068);
nor UO_596 (O_596,N_8608,N_9443);
nand UO_597 (O_597,N_7876,N_8859);
nor UO_598 (O_598,N_9291,N_9786);
nand UO_599 (O_599,N_7578,N_8032);
or UO_600 (O_600,N_8458,N_8085);
or UO_601 (O_601,N_9395,N_8355);
and UO_602 (O_602,N_8065,N_9282);
nand UO_603 (O_603,N_9078,N_8339);
and UO_604 (O_604,N_8654,N_9770);
nand UO_605 (O_605,N_7851,N_8721);
nor UO_606 (O_606,N_8262,N_9825);
nand UO_607 (O_607,N_8807,N_8887);
and UO_608 (O_608,N_9157,N_8055);
or UO_609 (O_609,N_8716,N_9260);
nor UO_610 (O_610,N_9928,N_7784);
or UO_611 (O_611,N_8821,N_8614);
nor UO_612 (O_612,N_9333,N_9699);
and UO_613 (O_613,N_8096,N_7510);
nor UO_614 (O_614,N_9542,N_8795);
xor UO_615 (O_615,N_9648,N_8315);
nor UO_616 (O_616,N_8684,N_7625);
and UO_617 (O_617,N_9047,N_8573);
and UO_618 (O_618,N_7937,N_8718);
nor UO_619 (O_619,N_8460,N_8714);
and UO_620 (O_620,N_7588,N_8572);
or UO_621 (O_621,N_8612,N_8282);
and UO_622 (O_622,N_8353,N_9205);
nand UO_623 (O_623,N_8409,N_7800);
nand UO_624 (O_624,N_9914,N_9971);
or UO_625 (O_625,N_8993,N_9004);
nor UO_626 (O_626,N_7810,N_9726);
and UO_627 (O_627,N_8979,N_9400);
or UO_628 (O_628,N_7843,N_8467);
and UO_629 (O_629,N_8338,N_7932);
or UO_630 (O_630,N_9585,N_8272);
nand UO_631 (O_631,N_9057,N_9749);
and UO_632 (O_632,N_9796,N_7766);
nor UO_633 (O_633,N_9966,N_9498);
xnor UO_634 (O_634,N_9323,N_9689);
nand UO_635 (O_635,N_7896,N_9046);
nor UO_636 (O_636,N_9647,N_8022);
and UO_637 (O_637,N_7814,N_9241);
and UO_638 (O_638,N_8551,N_9993);
xnor UO_639 (O_639,N_8295,N_9736);
and UO_640 (O_640,N_9466,N_9741);
and UO_641 (O_641,N_9230,N_9008);
and UO_642 (O_642,N_9532,N_9232);
and UO_643 (O_643,N_8932,N_8968);
or UO_644 (O_644,N_8178,N_7984);
nand UO_645 (O_645,N_8906,N_9892);
and UO_646 (O_646,N_9507,N_8284);
nand UO_647 (O_647,N_8475,N_8673);
or UO_648 (O_648,N_8849,N_8421);
or UO_649 (O_649,N_9556,N_9578);
or UO_650 (O_650,N_8244,N_7945);
nor UO_651 (O_651,N_8778,N_8812);
nor UO_652 (O_652,N_9805,N_9486);
xnor UO_653 (O_653,N_7926,N_9936);
nor UO_654 (O_654,N_7714,N_8650);
and UO_655 (O_655,N_9112,N_7847);
and UO_656 (O_656,N_9547,N_9052);
nor UO_657 (O_657,N_8026,N_8729);
or UO_658 (O_658,N_8142,N_9649);
nand UO_659 (O_659,N_9030,N_7769);
or UO_660 (O_660,N_9789,N_7832);
and UO_661 (O_661,N_8400,N_9005);
and UO_662 (O_662,N_9681,N_9912);
nand UO_663 (O_663,N_8236,N_8334);
nor UO_664 (O_664,N_8843,N_8129);
nor UO_665 (O_665,N_9869,N_8095);
nor UO_666 (O_666,N_9973,N_9801);
nand UO_667 (O_667,N_9406,N_9349);
nor UO_668 (O_668,N_7635,N_9643);
or UO_669 (O_669,N_8705,N_9894);
and UO_670 (O_670,N_9679,N_9706);
and UO_671 (O_671,N_8019,N_9051);
or UO_672 (O_672,N_8465,N_7890);
or UO_673 (O_673,N_9416,N_8874);
nand UO_674 (O_674,N_9848,N_9970);
or UO_675 (O_675,N_8362,N_9822);
and UO_676 (O_676,N_9651,N_8582);
nor UO_677 (O_677,N_9382,N_7749);
nor UO_678 (O_678,N_8106,N_9727);
nand UO_679 (O_679,N_7776,N_9860);
and UO_680 (O_680,N_8232,N_7570);
or UO_681 (O_681,N_9824,N_9186);
nand UO_682 (O_682,N_9755,N_8253);
or UO_683 (O_683,N_8151,N_7687);
xnor UO_684 (O_684,N_9045,N_8680);
or UO_685 (O_685,N_9102,N_9350);
and UO_686 (O_686,N_8250,N_8424);
nand UO_687 (O_687,N_9764,N_8048);
and UO_688 (O_688,N_9179,N_7842);
nor UO_689 (O_689,N_9310,N_8356);
nor UO_690 (O_690,N_8040,N_8535);
and UO_691 (O_691,N_7772,N_8771);
and UO_692 (O_692,N_7942,N_8502);
and UO_693 (O_693,N_8446,N_9272);
nand UO_694 (O_694,N_8878,N_8497);
or UO_695 (O_695,N_8579,N_9155);
or UO_696 (O_696,N_7633,N_8071);
nand UO_697 (O_697,N_8811,N_9397);
or UO_698 (O_698,N_8836,N_7550);
or UO_699 (O_699,N_8143,N_9244);
nor UO_700 (O_700,N_8734,N_9208);
and UO_701 (O_701,N_9504,N_8975);
nand UO_702 (O_702,N_8749,N_9570);
nor UO_703 (O_703,N_9701,N_9017);
or UO_704 (O_704,N_7860,N_8427);
nand UO_705 (O_705,N_8985,N_9368);
or UO_706 (O_706,N_9138,N_7885);
and UO_707 (O_707,N_7538,N_8359);
nand UO_708 (O_708,N_8367,N_7764);
nor UO_709 (O_709,N_8921,N_8831);
nand UO_710 (O_710,N_9160,N_9758);
and UO_711 (O_711,N_9909,N_8642);
nor UO_712 (O_712,N_9503,N_8645);
nor UO_713 (O_713,N_7565,N_9180);
and UO_714 (O_714,N_8477,N_8305);
or UO_715 (O_715,N_9020,N_8220);
nand UO_716 (O_716,N_7716,N_7611);
nor UO_717 (O_717,N_9091,N_8797);
and UO_718 (O_718,N_9195,N_9148);
or UO_719 (O_719,N_9872,N_8640);
nand UO_720 (O_720,N_9016,N_7998);
and UO_721 (O_721,N_9271,N_9481);
nor UO_722 (O_722,N_8087,N_9839);
and UO_723 (O_723,N_7924,N_8219);
nand UO_724 (O_724,N_8856,N_8911);
and UO_725 (O_725,N_9059,N_7830);
and UO_726 (O_726,N_9899,N_8155);
and UO_727 (O_727,N_9545,N_9332);
or UO_728 (O_728,N_9405,N_9541);
or UO_729 (O_729,N_9015,N_8737);
nor UO_730 (O_730,N_8625,N_8857);
or UO_731 (O_731,N_8431,N_9756);
or UO_732 (O_732,N_9044,N_8452);
and UO_733 (O_733,N_9734,N_8119);
nand UO_734 (O_734,N_8233,N_9721);
nand UO_735 (O_735,N_9320,N_8730);
nor UO_736 (O_736,N_9630,N_8226);
and UO_737 (O_737,N_9079,N_7593);
and UO_738 (O_738,N_9887,N_8936);
nand UO_739 (O_739,N_8489,N_7672);
nor UO_740 (O_740,N_8506,N_8958);
nor UO_741 (O_741,N_9754,N_9196);
xor UO_742 (O_742,N_7629,N_7763);
xor UO_743 (O_743,N_9170,N_9785);
or UO_744 (O_744,N_8149,N_9961);
nor UO_745 (O_745,N_8946,N_8786);
nand UO_746 (O_746,N_9949,N_8792);
and UO_747 (O_747,N_7798,N_9393);
and UO_748 (O_748,N_8643,N_9485);
or UO_749 (O_749,N_9167,N_9619);
or UO_750 (O_750,N_8408,N_9958);
nor UO_751 (O_751,N_9109,N_8263);
nand UO_752 (O_752,N_8883,N_8298);
nand UO_753 (O_753,N_9669,N_8959);
and UO_754 (O_754,N_7751,N_8838);
and UO_755 (O_755,N_8971,N_7639);
or UO_756 (O_756,N_9229,N_7908);
and UO_757 (O_757,N_9488,N_7874);
or UO_758 (O_758,N_9564,N_8311);
nor UO_759 (O_759,N_9903,N_8690);
and UO_760 (O_760,N_9191,N_8554);
and UO_761 (O_761,N_8033,N_9299);
nand UO_762 (O_762,N_7950,N_8394);
xor UO_763 (O_763,N_8309,N_9806);
or UO_764 (O_764,N_8357,N_9251);
nand UO_765 (O_765,N_9175,N_7728);
and UO_766 (O_766,N_9823,N_8208);
nor UO_767 (O_767,N_8024,N_7686);
nand UO_768 (O_768,N_8549,N_7938);
nand UO_769 (O_769,N_7804,N_7787);
or UO_770 (O_770,N_8872,N_7873);
nor UO_771 (O_771,N_9686,N_9011);
nor UO_772 (O_772,N_9944,N_9204);
nor UO_773 (O_773,N_9444,N_8313);
and UO_774 (O_774,N_7948,N_8647);
nand UO_775 (O_775,N_9691,N_8082);
xnor UO_776 (O_776,N_8802,N_9761);
and UO_777 (O_777,N_8222,N_9166);
and UO_778 (O_778,N_9645,N_9213);
nand UO_779 (O_779,N_9898,N_8628);
nor UO_780 (O_780,N_7675,N_9339);
or UO_781 (O_781,N_8691,N_7529);
or UO_782 (O_782,N_9713,N_8459);
and UO_783 (O_783,N_7640,N_7526);
and UO_784 (O_784,N_9760,N_7818);
or UO_785 (O_785,N_8808,N_9609);
nor UO_786 (O_786,N_9635,N_9537);
nand UO_787 (O_787,N_7738,N_8661);
or UO_788 (O_788,N_9122,N_8434);
nand UO_789 (O_789,N_7604,N_8114);
or UO_790 (O_790,N_9905,N_9539);
nand UO_791 (O_791,N_7590,N_7758);
nand UO_792 (O_792,N_8194,N_8956);
and UO_793 (O_793,N_8867,N_8495);
and UO_794 (O_794,N_8565,N_9753);
nand UO_795 (O_795,N_8986,N_9347);
and UO_796 (O_796,N_9224,N_9048);
nor UO_797 (O_797,N_9279,N_9572);
or UO_798 (O_798,N_7806,N_8123);
and UO_799 (O_799,N_9763,N_7756);
or UO_800 (O_800,N_7855,N_8663);
nor UO_801 (O_801,N_7654,N_9676);
or UO_802 (O_802,N_8935,N_9010);
or UO_803 (O_803,N_8188,N_9927);
or UO_804 (O_804,N_8733,N_9385);
or UO_805 (O_805,N_7698,N_7947);
and UO_806 (O_806,N_7571,N_8969);
and UO_807 (O_807,N_7727,N_9192);
nand UO_808 (O_808,N_9895,N_9496);
nor UO_809 (O_809,N_7644,N_8079);
and UO_810 (O_810,N_7850,N_7697);
or UO_811 (O_811,N_9399,N_7867);
nor UO_812 (O_812,N_9002,N_9595);
or UO_813 (O_813,N_8655,N_9816);
and UO_814 (O_814,N_8419,N_9529);
nor UO_815 (O_815,N_8229,N_8141);
and UO_816 (O_816,N_7914,N_9389);
nor UO_817 (O_817,N_7707,N_7789);
and UO_818 (O_818,N_8850,N_9220);
nand UO_819 (O_819,N_8437,N_8209);
nand UO_820 (O_820,N_8731,N_7953);
nor UO_821 (O_821,N_9633,N_7638);
or UO_822 (O_822,N_7549,N_7817);
or UO_823 (O_823,N_8366,N_9495);
or UO_824 (O_824,N_7531,N_9608);
nand UO_825 (O_825,N_9039,N_7523);
or UO_826 (O_826,N_8389,N_7678);
nand UO_827 (O_827,N_8425,N_8719);
nor UO_828 (O_828,N_9245,N_7963);
nor UO_829 (O_829,N_7912,N_8299);
nand UO_830 (O_830,N_7759,N_9838);
or UO_831 (O_831,N_8407,N_8001);
or UO_832 (O_832,N_8393,N_9603);
and UO_833 (O_833,N_8350,N_8510);
and UO_834 (O_834,N_8153,N_8081);
nor UO_835 (O_835,N_9256,N_8090);
nor UO_836 (O_836,N_7972,N_8177);
and UO_837 (O_837,N_9236,N_8107);
xnor UO_838 (O_838,N_8570,N_9396);
nor UO_839 (O_839,N_8967,N_7755);
and UO_840 (O_840,N_8089,N_7871);
nor UO_841 (O_841,N_8375,N_8886);
nor UO_842 (O_842,N_9021,N_9778);
nor UO_843 (O_843,N_7670,N_8738);
and UO_844 (O_844,N_9053,N_8700);
and UO_845 (O_845,N_9576,N_7801);
or UO_846 (O_846,N_9414,N_9459);
nor UO_847 (O_847,N_9108,N_9729);
nand UO_848 (O_848,N_9447,N_8025);
nor UO_849 (O_849,N_9938,N_8694);
nor UO_850 (O_850,N_8273,N_9606);
nand UO_851 (O_851,N_9031,N_8261);
and UO_852 (O_852,N_8395,N_8162);
nand UO_853 (O_853,N_9589,N_8994);
or UO_854 (O_854,N_8471,N_9225);
nor UO_855 (O_855,N_9777,N_8175);
and UO_856 (O_856,N_8532,N_9762);
nor UO_857 (O_857,N_9840,N_8152);
nand UO_858 (O_858,N_9027,N_8333);
and UO_859 (O_859,N_8116,N_8555);
nand UO_860 (O_860,N_8782,N_9757);
nand UO_861 (O_861,N_9194,N_9745);
and UO_862 (O_862,N_7509,N_7739);
nor UO_863 (O_863,N_8928,N_8540);
and UO_864 (O_864,N_9999,N_7692);
or UO_865 (O_865,N_8010,N_9820);
xnor UO_866 (O_866,N_8340,N_9670);
nand UO_867 (O_867,N_9240,N_8884);
nor UO_868 (O_868,N_8646,N_8634);
or UO_869 (O_869,N_7581,N_7566);
or UO_870 (O_870,N_7534,N_9582);
and UO_871 (O_871,N_8566,N_9808);
and UO_872 (O_872,N_7641,N_7634);
or UO_873 (O_873,N_7858,N_9433);
nor UO_874 (O_874,N_9640,N_8557);
or UO_875 (O_875,N_8371,N_8609);
nand UO_876 (O_876,N_8406,N_8418);
nor UO_877 (O_877,N_9210,N_9530);
and UO_878 (O_878,N_8420,N_8626);
or UO_879 (O_879,N_9804,N_8330);
or UO_880 (O_880,N_9948,N_7833);
and UO_881 (O_881,N_8126,N_9782);
or UO_882 (O_882,N_9372,N_8798);
nor UO_883 (O_883,N_8457,N_8764);
xnor UO_884 (O_884,N_8140,N_9161);
and UO_885 (O_885,N_9674,N_9562);
or UO_886 (O_886,N_9638,N_7839);
and UO_887 (O_887,N_9352,N_9360);
and UO_888 (O_888,N_7790,N_8380);
or UO_889 (O_889,N_8159,N_8600);
and UO_890 (O_890,N_8160,N_8970);
and UO_891 (O_891,N_8034,N_9436);
nand UO_892 (O_892,N_7977,N_8875);
and UO_893 (O_893,N_9217,N_8287);
nand UO_894 (O_894,N_8514,N_9716);
and UO_895 (O_895,N_8972,N_7657);
nand UO_896 (O_896,N_8657,N_8042);
and UO_897 (O_897,N_7664,N_7594);
and UO_898 (O_898,N_8204,N_8806);
and UO_899 (O_899,N_9499,N_9402);
nand UO_900 (O_900,N_8060,N_7512);
nor UO_901 (O_901,N_7729,N_8285);
and UO_902 (O_902,N_7954,N_9286);
xnor UO_903 (O_903,N_7618,N_9821);
or UO_904 (O_904,N_8852,N_9410);
xor UO_905 (O_905,N_9717,N_9419);
nor UO_906 (O_906,N_9452,N_7630);
or UO_907 (O_907,N_8829,N_7961);
nor UO_908 (O_908,N_8377,N_9696);
and UO_909 (O_909,N_8296,N_8621);
or UO_910 (O_910,N_7886,N_8914);
or UO_911 (O_911,N_8681,N_9885);
or UO_912 (O_912,N_8675,N_7965);
and UO_913 (O_913,N_9863,N_9866);
nor UO_914 (O_914,N_9381,N_8216);
nand UO_915 (O_915,N_9767,N_8289);
nor UO_916 (O_916,N_7920,N_9001);
nand UO_917 (O_917,N_7781,N_9292);
nor UO_918 (O_918,N_9702,N_8800);
nand UO_919 (O_919,N_9626,N_8043);
nor UO_920 (O_920,N_7959,N_9463);
nand UO_921 (O_921,N_9425,N_8571);
nor UO_922 (O_922,N_8917,N_8348);
nor UO_923 (O_923,N_9216,N_7812);
or UO_924 (O_924,N_9429,N_7809);
xnor UO_925 (O_925,N_9242,N_9634);
or UO_926 (O_926,N_8799,N_7663);
and UO_927 (O_927,N_9003,N_9203);
or UO_928 (O_928,N_8539,N_8905);
nand UO_929 (O_929,N_9922,N_9247);
nor UO_930 (O_930,N_8982,N_9546);
or UO_931 (O_931,N_9212,N_7682);
or UO_932 (O_932,N_8939,N_8098);
nor UO_933 (O_933,N_8441,N_8687);
nor UO_934 (O_934,N_7848,N_8173);
or UO_935 (O_935,N_7643,N_9845);
and UO_936 (O_936,N_9552,N_7536);
and UO_937 (O_937,N_9995,N_9881);
nand UO_938 (O_938,N_7539,N_7782);
and UO_939 (O_939,N_9263,N_8822);
and UO_940 (O_940,N_8521,N_8903);
nand UO_941 (O_941,N_9743,N_8365);
nand UO_942 (O_942,N_9853,N_9189);
or UO_943 (O_943,N_9652,N_8676);
and UO_944 (O_944,N_8235,N_8918);
and UO_945 (O_945,N_9998,N_9037);
nand UO_946 (O_946,N_8702,N_9099);
and UO_947 (O_947,N_9341,N_9988);
nand UO_948 (O_948,N_9996,N_7975);
nand UO_949 (O_949,N_7872,N_9772);
and UO_950 (O_950,N_7968,N_9374);
or UO_951 (O_951,N_8866,N_9316);
nand UO_952 (O_952,N_8598,N_8278);
or UO_953 (O_953,N_8894,N_9116);
nand UO_954 (O_954,N_8550,N_8066);
or UO_955 (O_955,N_9842,N_8652);
and UO_956 (O_956,N_9594,N_8398);
nor UO_957 (O_957,N_8103,N_8941);
and UO_958 (O_958,N_9515,N_8045);
and UO_959 (O_959,N_9391,N_8028);
nor UO_960 (O_960,N_7605,N_8832);
and UO_961 (O_961,N_8354,N_8325);
and UO_962 (O_962,N_9610,N_8931);
nor UO_963 (O_963,N_7708,N_8563);
nor UO_964 (O_964,N_7870,N_9462);
nand UO_965 (O_965,N_9942,N_8885);
or UO_966 (O_966,N_8039,N_9140);
or UO_967 (O_967,N_8486,N_8317);
and UO_968 (O_968,N_7994,N_9704);
and UO_969 (O_969,N_8607,N_8632);
nor UO_970 (O_970,N_7673,N_9303);
nand UO_971 (O_971,N_8322,N_8275);
or UO_972 (O_972,N_7767,N_8342);
nor UO_973 (O_973,N_9787,N_8163);
nand UO_974 (O_974,N_7815,N_7808);
nor UO_975 (O_975,N_7552,N_8902);
and UO_976 (O_976,N_8374,N_9992);
and UO_977 (O_977,N_9656,N_7750);
and UO_978 (O_978,N_8904,N_8241);
nor UO_979 (O_979,N_9075,N_9527);
nand UO_980 (O_980,N_8138,N_9759);
or UO_981 (O_981,N_8765,N_7680);
and UO_982 (O_982,N_8249,N_9141);
nand UO_983 (O_983,N_7811,N_9424);
and UO_984 (O_984,N_8998,N_9510);
nor UO_985 (O_985,N_9945,N_7515);
nand UO_986 (O_986,N_9197,N_8723);
nand UO_987 (O_987,N_8464,N_8445);
or UO_988 (O_988,N_8926,N_9130);
nor UO_989 (O_989,N_9923,N_9865);
nand UO_990 (O_990,N_9275,N_7648);
nor UO_991 (O_991,N_8816,N_9356);
nand UO_992 (O_992,N_9521,N_9233);
nand UO_993 (O_993,N_9627,N_7647);
xor UO_994 (O_994,N_7671,N_7845);
nand UO_995 (O_995,N_8005,N_8692);
or UO_996 (O_996,N_9309,N_8927);
nand UO_997 (O_997,N_8397,N_7612);
or UO_998 (O_998,N_9873,N_7865);
or UO_999 (O_999,N_9974,N_9937);
nand UO_1000 (O_1000,N_8405,N_7973);
nor UO_1001 (O_1001,N_9837,N_8767);
nand UO_1002 (O_1002,N_9018,N_8306);
xor UO_1003 (O_1003,N_7530,N_9428);
nand UO_1004 (O_1004,N_9284,N_9943);
or UO_1005 (O_1005,N_9827,N_8989);
and UO_1006 (O_1006,N_8258,N_8335);
nor UO_1007 (O_1007,N_8364,N_9359);
or UO_1008 (O_1008,N_9596,N_9666);
or UO_1009 (O_1009,N_7704,N_9882);
nor UO_1010 (O_1010,N_8610,N_9209);
nor UO_1011 (O_1011,N_8137,N_7632);
and UO_1012 (O_1012,N_9910,N_8592);
and UO_1013 (O_1013,N_8139,N_9593);
and UO_1014 (O_1014,N_7703,N_9631);
and UO_1015 (O_1015,N_9201,N_9738);
nor UO_1016 (O_1016,N_9365,N_7778);
nor UO_1017 (O_1017,N_8174,N_8992);
and UO_1018 (O_1018,N_9769,N_8960);
and UO_1019 (O_1019,N_9340,N_9497);
nor UO_1020 (O_1020,N_8444,N_8907);
nand UO_1021 (O_1021,N_7642,N_9957);
and UO_1022 (O_1022,N_7537,N_8341);
nand UO_1023 (O_1023,N_9458,N_9803);
or UO_1024 (O_1024,N_9493,N_9540);
nand UO_1025 (O_1025,N_9476,N_7527);
nor UO_1026 (O_1026,N_7731,N_9776);
or UO_1027 (O_1027,N_7838,N_9355);
or UO_1028 (O_1028,N_8326,N_8379);
or UO_1029 (O_1029,N_9487,N_9711);
or UO_1030 (O_1030,N_9177,N_9307);
or UO_1031 (O_1031,N_9375,N_8402);
nand UO_1032 (O_1032,N_9253,N_9438);
nor UO_1033 (O_1033,N_9090,N_9983);
or UO_1034 (O_1034,N_7829,N_8697);
nand UO_1035 (O_1035,N_7689,N_8710);
nor UO_1036 (O_1036,N_9207,N_8525);
and UO_1037 (O_1037,N_8896,N_9650);
nand UO_1038 (O_1038,N_8964,N_9178);
and UO_1039 (O_1039,N_9867,N_7837);
or UO_1040 (O_1040,N_8913,N_9484);
nand UO_1041 (O_1041,N_9723,N_8929);
nand UO_1042 (O_1042,N_9353,N_8930);
nor UO_1043 (O_1043,N_8966,N_7613);
or UO_1044 (O_1044,N_9379,N_9456);
nand UO_1045 (O_1045,N_8677,N_9269);
and UO_1046 (O_1046,N_9671,N_9032);
or UO_1047 (O_1047,N_7941,N_8791);
and UO_1048 (O_1048,N_7718,N_9653);
or UO_1049 (O_1049,N_8644,N_8329);
and UO_1050 (O_1050,N_9121,N_7925);
nor UO_1051 (O_1051,N_8481,N_9953);
nand UO_1052 (O_1052,N_8756,N_7737);
and UO_1053 (O_1053,N_9854,N_9543);
nor UO_1054 (O_1054,N_9917,N_9791);
and UO_1055 (O_1055,N_8187,N_8117);
or UO_1056 (O_1056,N_9033,N_8830);
nor UO_1057 (O_1057,N_8461,N_7668);
or UO_1058 (O_1058,N_9060,N_7603);
and UO_1059 (O_1059,N_8544,N_9482);
or UO_1060 (O_1060,N_8693,N_9239);
nor UO_1061 (O_1061,N_8711,N_8007);
nand UO_1062 (O_1062,N_7713,N_9590);
nand UO_1063 (O_1063,N_9907,N_9261);
and UO_1064 (O_1064,N_7732,N_9420);
or UO_1065 (O_1065,N_8827,N_9377);
nand UO_1066 (O_1066,N_7883,N_8629);
or UO_1067 (O_1067,N_9050,N_9440);
nor UO_1068 (O_1068,N_8105,N_8622);
nand UO_1069 (O_1069,N_9464,N_8627);
nand UO_1070 (O_1070,N_8336,N_7921);
or UO_1071 (O_1071,N_9469,N_9407);
and UO_1072 (O_1072,N_7846,N_9925);
nand UO_1073 (O_1073,N_8824,N_9248);
xnor UO_1074 (O_1074,N_9750,N_8965);
or UO_1075 (O_1075,N_8618,N_8868);
nor UO_1076 (O_1076,N_8533,N_9142);
or UO_1077 (O_1077,N_8451,N_7791);
nor UO_1078 (O_1078,N_8376,N_9453);
nand UO_1079 (O_1079,N_8817,N_7988);
nor UO_1080 (O_1080,N_9491,N_9939);
or UO_1081 (O_1081,N_8146,N_8056);
or UO_1082 (O_1082,N_8984,N_8722);
nand UO_1083 (O_1083,N_8923,N_9480);
nor UO_1084 (O_1084,N_8067,N_9563);
and UO_1085 (O_1085,N_9921,N_7569);
and UO_1086 (O_1086,N_7877,N_7868);
or UO_1087 (O_1087,N_9062,N_8777);
and UO_1088 (O_1088,N_7864,N_8529);
nand UO_1089 (O_1089,N_8518,N_9550);
and UO_1090 (O_1090,N_8682,N_8810);
and UO_1091 (O_1091,N_9302,N_9250);
or UO_1092 (O_1092,N_9345,N_8120);
nor UO_1093 (O_1093,N_9325,N_9989);
nor UO_1094 (O_1094,N_9598,N_9513);
nor UO_1095 (O_1095,N_8062,N_8498);
nand UO_1096 (O_1096,N_9644,N_8839);
nor UO_1097 (O_1097,N_9387,N_9561);
nand UO_1098 (O_1098,N_8331,N_9249);
nand UO_1099 (O_1099,N_7541,N_9724);
nand UO_1100 (O_1100,N_9278,N_9526);
or UO_1101 (O_1101,N_9066,N_8104);
nand UO_1102 (O_1102,N_7888,N_9886);
nor UO_1103 (O_1103,N_9577,N_9383);
or UO_1104 (O_1104,N_8760,N_9780);
nand UO_1105 (O_1105,N_8200,N_9508);
or UO_1106 (O_1106,N_7882,N_8002);
and UO_1107 (O_1107,N_9828,N_8018);
and UO_1108 (O_1108,N_7554,N_8013);
and UO_1109 (O_1109,N_9893,N_7528);
and UO_1110 (O_1110,N_8157,N_9693);
nor UO_1111 (O_1111,N_7980,N_9390);
and UO_1112 (O_1112,N_9259,N_8670);
nand UO_1113 (O_1113,N_8412,N_9980);
nand UO_1114 (O_1114,N_8517,N_9362);
nand UO_1115 (O_1115,N_8006,N_7990);
nor UO_1116 (O_1116,N_8679,N_8717);
nor UO_1117 (O_1117,N_8027,N_9055);
nand UO_1118 (O_1118,N_7983,N_9455);
or UO_1119 (O_1119,N_9752,N_9987);
and UO_1120 (O_1120,N_7878,N_8269);
nor UO_1121 (O_1121,N_9089,N_7623);
or UO_1122 (O_1122,N_8448,N_7960);
and UO_1123 (O_1123,N_9137,N_9268);
nor UO_1124 (O_1124,N_9338,N_8574);
and UO_1125 (O_1125,N_8101,N_8847);
or UO_1126 (O_1126,N_8494,N_7561);
or UO_1127 (O_1127,N_9600,N_9528);
nor UO_1128 (O_1128,N_9289,N_7598);
nand UO_1129 (O_1129,N_8197,N_8576);
nor UO_1130 (O_1130,N_7658,N_8987);
or UO_1131 (O_1131,N_9531,N_9054);
or UO_1132 (O_1132,N_7931,N_7884);
or UO_1133 (O_1133,N_9128,N_8934);
nand UO_1134 (O_1134,N_8069,N_7502);
nand UO_1135 (O_1135,N_8381,N_8332);
nor UO_1136 (O_1136,N_8052,N_9367);
nor UO_1137 (O_1137,N_8358,N_9500);
or UO_1138 (O_1138,N_8834,N_9566);
and UO_1139 (O_1139,N_9719,N_7958);
and UO_1140 (O_1140,N_7894,N_9305);
nand UO_1141 (O_1141,N_9799,N_7548);
nand UO_1142 (O_1142,N_9457,N_8190);
and UO_1143 (O_1143,N_8496,N_7816);
or UO_1144 (O_1144,N_9994,N_7752);
and UO_1145 (O_1145,N_8846,N_9426);
nand UO_1146 (O_1146,N_9025,N_9028);
and UO_1147 (O_1147,N_9984,N_7560);
and UO_1148 (O_1148,N_8648,N_9587);
nand UO_1149 (O_1149,N_7691,N_7823);
nand UO_1150 (O_1150,N_9376,N_8308);
or UO_1151 (O_1151,N_9553,N_9849);
nor UO_1152 (O_1152,N_7568,N_9950);
nand UO_1153 (O_1153,N_9336,N_9614);
xor UO_1154 (O_1154,N_8524,N_7904);
nand UO_1155 (O_1155,N_9534,N_7655);
or UO_1156 (O_1156,N_8234,N_9437);
or UO_1157 (O_1157,N_8639,N_8031);
nand UO_1158 (O_1158,N_8909,N_7711);
or UO_1159 (O_1159,N_8227,N_8435);
xor UO_1160 (O_1160,N_7992,N_7533);
nor UO_1161 (O_1161,N_9147,N_8803);
and UO_1162 (O_1162,N_8423,N_9298);
and UO_1163 (O_1163,N_7709,N_9751);
or UO_1164 (O_1164,N_8191,N_7669);
and UO_1165 (O_1165,N_7627,N_8787);
nand UO_1166 (O_1166,N_9817,N_9672);
or UO_1167 (O_1167,N_8920,N_7559);
and UO_1168 (O_1168,N_8214,N_8591);
nor UO_1169 (O_1169,N_8890,N_8671);
and UO_1170 (O_1170,N_7584,N_9077);
or UO_1171 (O_1171,N_7600,N_9277);
and UO_1172 (O_1172,N_7520,N_7717);
and UO_1173 (O_1173,N_9621,N_7799);
nand UO_1174 (O_1174,N_9678,N_8422);
nor UO_1175 (O_1175,N_8881,N_9009);
nand UO_1176 (O_1176,N_8154,N_8689);
nor UO_1177 (O_1177,N_8012,N_9126);
and UO_1178 (O_1178,N_7710,N_7802);
nand UO_1179 (O_1179,N_8980,N_9968);
nand UO_1180 (O_1180,N_7540,N_9472);
nor UO_1181 (O_1181,N_8136,N_7951);
and UO_1182 (O_1182,N_8247,N_7684);
nor UO_1183 (O_1183,N_8658,N_8862);
nand UO_1184 (O_1184,N_9494,N_9809);
nand UO_1185 (O_1185,N_8876,N_8915);
and UO_1186 (O_1186,N_8382,N_9654);
nor UO_1187 (O_1187,N_8221,N_8624);
xor UO_1188 (O_1188,N_8228,N_8511);
or UO_1189 (O_1189,N_9146,N_8869);
xor UO_1190 (O_1190,N_9388,N_7956);
and UO_1191 (O_1191,N_8748,N_9366);
nand UO_1192 (O_1192,N_7796,N_8949);
and UO_1193 (O_1193,N_9297,N_8537);
and UO_1194 (O_1194,N_8864,N_8324);
nor UO_1195 (O_1195,N_9934,N_7562);
or UO_1196 (O_1196,N_8509,N_8401);
and UO_1197 (O_1197,N_9781,N_7760);
nand UO_1198 (O_1198,N_9792,N_9023);
and UO_1199 (O_1199,N_9264,N_9334);
nor UO_1200 (O_1200,N_7563,N_8585);
nand UO_1201 (O_1201,N_7744,N_9646);
nor UO_1202 (O_1202,N_7683,N_9036);
or UO_1203 (O_1203,N_7786,N_8613);
and UO_1204 (O_1204,N_8372,N_9168);
nand UO_1205 (O_1205,N_9364,N_9725);
or UO_1206 (O_1206,N_7667,N_7899);
or UO_1207 (O_1207,N_9415,N_7831);
nor UO_1208 (O_1208,N_7610,N_9655);
or UO_1209 (O_1209,N_7688,N_7521);
and UO_1210 (O_1210,N_9206,N_9612);
xnor UO_1211 (O_1211,N_9558,N_9788);
and UO_1212 (O_1212,N_8207,N_8703);
and UO_1213 (O_1213,N_9771,N_8879);
or UO_1214 (O_1214,N_7841,N_7742);
nand UO_1215 (O_1215,N_8583,N_8182);
or UO_1216 (O_1216,N_7607,N_7861);
nand UO_1217 (O_1217,N_9737,N_7762);
and UO_1218 (O_1218,N_9901,N_8727);
or UO_1219 (O_1219,N_8858,N_9007);
and UO_1220 (O_1220,N_9710,N_7879);
or UO_1221 (O_1221,N_8203,N_7952);
xor UO_1222 (O_1222,N_8150,N_8604);
nand UO_1223 (O_1223,N_8008,N_9287);
and UO_1224 (O_1224,N_8578,N_8709);
xnor UO_1225 (O_1225,N_9523,N_9795);
nor UO_1226 (O_1226,N_8319,N_9043);
nand UO_1227 (O_1227,N_7577,N_9784);
nor UO_1228 (O_1228,N_8605,N_9439);
nor UO_1229 (O_1229,N_8877,N_7653);
or UO_1230 (O_1230,N_7820,N_7935);
nor UO_1231 (O_1231,N_8030,N_8775);
nand UO_1232 (O_1232,N_7606,N_8699);
or UO_1233 (O_1233,N_9185,N_8933);
or UO_1234 (O_1234,N_9812,N_8440);
nor UO_1235 (O_1235,N_7720,N_9317);
xor UO_1236 (O_1236,N_8483,N_9354);
nand UO_1237 (O_1237,N_9662,N_8058);
nand UO_1238 (O_1238,N_9190,N_8840);
or UO_1239 (O_1239,N_8429,N_9856);
nor UO_1240 (O_1240,N_8785,N_8619);
and UO_1241 (O_1241,N_9683,N_7544);
and UO_1242 (O_1242,N_8995,N_7770);
nor UO_1243 (O_1243,N_8280,N_7857);
nand UO_1244 (O_1244,N_7773,N_8745);
nand UO_1245 (O_1245,N_7608,N_9188);
nor UO_1246 (O_1246,N_9708,N_8659);
nor UO_1247 (O_1247,N_9623,N_8520);
and UO_1248 (O_1248,N_7999,N_8999);
xnor UO_1249 (O_1249,N_7700,N_7761);
and UO_1250 (O_1250,N_8511,N_8838);
and UO_1251 (O_1251,N_9764,N_9088);
or UO_1252 (O_1252,N_8694,N_9540);
nand UO_1253 (O_1253,N_7678,N_7516);
or UO_1254 (O_1254,N_8838,N_7758);
xnor UO_1255 (O_1255,N_9942,N_7515);
or UO_1256 (O_1256,N_9527,N_9735);
nand UO_1257 (O_1257,N_7883,N_7863);
nand UO_1258 (O_1258,N_8887,N_9574);
and UO_1259 (O_1259,N_9491,N_8774);
or UO_1260 (O_1260,N_8460,N_9411);
and UO_1261 (O_1261,N_8558,N_9082);
and UO_1262 (O_1262,N_9493,N_9868);
and UO_1263 (O_1263,N_8526,N_8731);
and UO_1264 (O_1264,N_7627,N_8192);
nor UO_1265 (O_1265,N_9776,N_9858);
and UO_1266 (O_1266,N_8363,N_9038);
and UO_1267 (O_1267,N_8400,N_8382);
nor UO_1268 (O_1268,N_8749,N_9718);
or UO_1269 (O_1269,N_9298,N_8610);
nor UO_1270 (O_1270,N_9062,N_7796);
and UO_1271 (O_1271,N_9874,N_7861);
or UO_1272 (O_1272,N_8025,N_9848);
xnor UO_1273 (O_1273,N_8120,N_9461);
or UO_1274 (O_1274,N_7714,N_7585);
nand UO_1275 (O_1275,N_8014,N_9490);
nand UO_1276 (O_1276,N_9098,N_8921);
nor UO_1277 (O_1277,N_8850,N_9225);
and UO_1278 (O_1278,N_9030,N_8184);
nor UO_1279 (O_1279,N_7914,N_7651);
or UO_1280 (O_1280,N_9543,N_7937);
nand UO_1281 (O_1281,N_8739,N_8649);
nor UO_1282 (O_1282,N_9386,N_7959);
nand UO_1283 (O_1283,N_8879,N_9395);
nand UO_1284 (O_1284,N_8744,N_9646);
nand UO_1285 (O_1285,N_7770,N_9151);
nand UO_1286 (O_1286,N_9503,N_9787);
nand UO_1287 (O_1287,N_7708,N_7911);
and UO_1288 (O_1288,N_7510,N_8616);
or UO_1289 (O_1289,N_8533,N_7840);
or UO_1290 (O_1290,N_9992,N_7957);
nor UO_1291 (O_1291,N_8582,N_9619);
or UO_1292 (O_1292,N_9157,N_9935);
and UO_1293 (O_1293,N_7922,N_8834);
nand UO_1294 (O_1294,N_8516,N_8680);
xnor UO_1295 (O_1295,N_9965,N_8306);
nor UO_1296 (O_1296,N_7906,N_7623);
and UO_1297 (O_1297,N_7998,N_9592);
xor UO_1298 (O_1298,N_8305,N_7953);
nand UO_1299 (O_1299,N_9604,N_8651);
or UO_1300 (O_1300,N_8772,N_9248);
nor UO_1301 (O_1301,N_7725,N_8802);
and UO_1302 (O_1302,N_9065,N_9435);
and UO_1303 (O_1303,N_7734,N_7614);
nor UO_1304 (O_1304,N_8775,N_8361);
xor UO_1305 (O_1305,N_9653,N_8697);
or UO_1306 (O_1306,N_9188,N_8911);
or UO_1307 (O_1307,N_9583,N_8652);
or UO_1308 (O_1308,N_7928,N_8656);
nand UO_1309 (O_1309,N_9343,N_8468);
nand UO_1310 (O_1310,N_9365,N_9897);
and UO_1311 (O_1311,N_9238,N_8070);
nor UO_1312 (O_1312,N_9831,N_8769);
or UO_1313 (O_1313,N_9577,N_7965);
or UO_1314 (O_1314,N_9957,N_8718);
and UO_1315 (O_1315,N_7755,N_8297);
or UO_1316 (O_1316,N_7819,N_9059);
nor UO_1317 (O_1317,N_8247,N_7990);
and UO_1318 (O_1318,N_7940,N_9056);
or UO_1319 (O_1319,N_8088,N_9592);
nand UO_1320 (O_1320,N_8412,N_8989);
and UO_1321 (O_1321,N_8623,N_8207);
or UO_1322 (O_1322,N_9279,N_7919);
and UO_1323 (O_1323,N_9343,N_8671);
nor UO_1324 (O_1324,N_9338,N_8026);
or UO_1325 (O_1325,N_9125,N_7651);
or UO_1326 (O_1326,N_9566,N_7964);
xnor UO_1327 (O_1327,N_8326,N_9053);
nand UO_1328 (O_1328,N_9905,N_7529);
nand UO_1329 (O_1329,N_7903,N_8300);
and UO_1330 (O_1330,N_9612,N_9644);
or UO_1331 (O_1331,N_7921,N_9836);
and UO_1332 (O_1332,N_8972,N_8289);
and UO_1333 (O_1333,N_7670,N_8433);
or UO_1334 (O_1334,N_7892,N_8701);
nand UO_1335 (O_1335,N_9628,N_9235);
or UO_1336 (O_1336,N_7972,N_9118);
or UO_1337 (O_1337,N_9338,N_9012);
or UO_1338 (O_1338,N_8202,N_7770);
and UO_1339 (O_1339,N_8372,N_8923);
nand UO_1340 (O_1340,N_8483,N_8277);
or UO_1341 (O_1341,N_8590,N_8442);
nor UO_1342 (O_1342,N_8995,N_9231);
and UO_1343 (O_1343,N_9902,N_8474);
and UO_1344 (O_1344,N_9257,N_8041);
nand UO_1345 (O_1345,N_9914,N_9666);
or UO_1346 (O_1346,N_8271,N_7642);
or UO_1347 (O_1347,N_9444,N_8550);
and UO_1348 (O_1348,N_8886,N_8376);
nor UO_1349 (O_1349,N_8465,N_9242);
and UO_1350 (O_1350,N_8471,N_9073);
nor UO_1351 (O_1351,N_8087,N_9213);
nor UO_1352 (O_1352,N_7791,N_9234);
and UO_1353 (O_1353,N_8720,N_8105);
or UO_1354 (O_1354,N_9860,N_9186);
or UO_1355 (O_1355,N_8398,N_7614);
or UO_1356 (O_1356,N_9328,N_8835);
or UO_1357 (O_1357,N_9594,N_9863);
and UO_1358 (O_1358,N_7774,N_7734);
nand UO_1359 (O_1359,N_7931,N_9781);
and UO_1360 (O_1360,N_7598,N_7723);
and UO_1361 (O_1361,N_7792,N_9433);
nand UO_1362 (O_1362,N_8238,N_8047);
or UO_1363 (O_1363,N_9482,N_9633);
nand UO_1364 (O_1364,N_8954,N_9070);
nor UO_1365 (O_1365,N_8331,N_8606);
nand UO_1366 (O_1366,N_7872,N_9352);
nand UO_1367 (O_1367,N_9972,N_9479);
xor UO_1368 (O_1368,N_9693,N_8628);
and UO_1369 (O_1369,N_9019,N_8540);
nor UO_1370 (O_1370,N_9464,N_8785);
nor UO_1371 (O_1371,N_7767,N_8149);
or UO_1372 (O_1372,N_8951,N_9337);
or UO_1373 (O_1373,N_9746,N_8892);
nor UO_1374 (O_1374,N_9201,N_9359);
and UO_1375 (O_1375,N_8150,N_8251);
or UO_1376 (O_1376,N_9534,N_7651);
nand UO_1377 (O_1377,N_7507,N_7516);
or UO_1378 (O_1378,N_7970,N_8196);
nor UO_1379 (O_1379,N_8616,N_9490);
or UO_1380 (O_1380,N_8098,N_9787);
nor UO_1381 (O_1381,N_8277,N_9296);
or UO_1382 (O_1382,N_9061,N_7753);
or UO_1383 (O_1383,N_9614,N_9951);
and UO_1384 (O_1384,N_8648,N_7665);
or UO_1385 (O_1385,N_8218,N_8027);
nor UO_1386 (O_1386,N_8763,N_9607);
nor UO_1387 (O_1387,N_9077,N_8816);
and UO_1388 (O_1388,N_8794,N_9838);
nor UO_1389 (O_1389,N_8154,N_9359);
or UO_1390 (O_1390,N_9224,N_8681);
nor UO_1391 (O_1391,N_7564,N_8156);
and UO_1392 (O_1392,N_9866,N_8170);
nand UO_1393 (O_1393,N_7985,N_9680);
nand UO_1394 (O_1394,N_8815,N_8399);
nand UO_1395 (O_1395,N_9486,N_8546);
nand UO_1396 (O_1396,N_7827,N_7531);
or UO_1397 (O_1397,N_7793,N_7957);
and UO_1398 (O_1398,N_8221,N_8254);
and UO_1399 (O_1399,N_9982,N_7606);
nand UO_1400 (O_1400,N_9830,N_7527);
or UO_1401 (O_1401,N_8398,N_9486);
nand UO_1402 (O_1402,N_9402,N_8036);
nand UO_1403 (O_1403,N_8274,N_9864);
nor UO_1404 (O_1404,N_9583,N_9802);
and UO_1405 (O_1405,N_9000,N_8671);
and UO_1406 (O_1406,N_8003,N_8524);
or UO_1407 (O_1407,N_9313,N_9181);
and UO_1408 (O_1408,N_7562,N_8532);
and UO_1409 (O_1409,N_8007,N_7914);
or UO_1410 (O_1410,N_7780,N_9521);
xor UO_1411 (O_1411,N_8881,N_7910);
or UO_1412 (O_1412,N_9057,N_8287);
and UO_1413 (O_1413,N_9417,N_9820);
nor UO_1414 (O_1414,N_8836,N_8692);
nand UO_1415 (O_1415,N_8124,N_7962);
nand UO_1416 (O_1416,N_9308,N_8273);
and UO_1417 (O_1417,N_8788,N_8403);
and UO_1418 (O_1418,N_9063,N_7507);
or UO_1419 (O_1419,N_7886,N_8613);
and UO_1420 (O_1420,N_8461,N_9152);
and UO_1421 (O_1421,N_8186,N_9333);
nor UO_1422 (O_1422,N_8170,N_9224);
and UO_1423 (O_1423,N_8746,N_9377);
nand UO_1424 (O_1424,N_8735,N_8403);
nor UO_1425 (O_1425,N_8256,N_7944);
nor UO_1426 (O_1426,N_8768,N_7834);
or UO_1427 (O_1427,N_7664,N_9220);
and UO_1428 (O_1428,N_9336,N_9093);
nand UO_1429 (O_1429,N_9144,N_8255);
nor UO_1430 (O_1430,N_8249,N_8691);
nand UO_1431 (O_1431,N_7784,N_8822);
nor UO_1432 (O_1432,N_8183,N_9743);
nand UO_1433 (O_1433,N_9241,N_8725);
and UO_1434 (O_1434,N_9766,N_8188);
and UO_1435 (O_1435,N_8394,N_8995);
and UO_1436 (O_1436,N_7792,N_9372);
nor UO_1437 (O_1437,N_9452,N_9275);
or UO_1438 (O_1438,N_8296,N_9681);
and UO_1439 (O_1439,N_7952,N_8431);
and UO_1440 (O_1440,N_7539,N_8751);
nor UO_1441 (O_1441,N_7605,N_9137);
nand UO_1442 (O_1442,N_9613,N_8253);
nand UO_1443 (O_1443,N_8851,N_7530);
nand UO_1444 (O_1444,N_9812,N_8438);
and UO_1445 (O_1445,N_7810,N_8425);
and UO_1446 (O_1446,N_7746,N_9165);
nor UO_1447 (O_1447,N_9455,N_8876);
or UO_1448 (O_1448,N_7612,N_9991);
nor UO_1449 (O_1449,N_8405,N_8742);
nor UO_1450 (O_1450,N_7966,N_7751);
nor UO_1451 (O_1451,N_9876,N_9270);
nand UO_1452 (O_1452,N_8871,N_8636);
or UO_1453 (O_1453,N_9175,N_8058);
nor UO_1454 (O_1454,N_8062,N_7774);
or UO_1455 (O_1455,N_7927,N_9425);
or UO_1456 (O_1456,N_8521,N_9366);
nand UO_1457 (O_1457,N_8828,N_9717);
and UO_1458 (O_1458,N_7693,N_7577);
or UO_1459 (O_1459,N_7962,N_8548);
and UO_1460 (O_1460,N_7594,N_8440);
or UO_1461 (O_1461,N_9372,N_9549);
or UO_1462 (O_1462,N_9496,N_9129);
or UO_1463 (O_1463,N_8259,N_8818);
and UO_1464 (O_1464,N_9075,N_9771);
nor UO_1465 (O_1465,N_8360,N_7845);
nand UO_1466 (O_1466,N_8058,N_8597);
or UO_1467 (O_1467,N_7638,N_9754);
or UO_1468 (O_1468,N_9495,N_9207);
and UO_1469 (O_1469,N_7653,N_9168);
nor UO_1470 (O_1470,N_7505,N_8859);
nor UO_1471 (O_1471,N_9543,N_9101);
and UO_1472 (O_1472,N_9828,N_9299);
and UO_1473 (O_1473,N_8919,N_9672);
nand UO_1474 (O_1474,N_7694,N_7547);
nand UO_1475 (O_1475,N_9440,N_7631);
or UO_1476 (O_1476,N_7540,N_9049);
or UO_1477 (O_1477,N_8579,N_9839);
nand UO_1478 (O_1478,N_8397,N_8894);
nand UO_1479 (O_1479,N_7741,N_9968);
or UO_1480 (O_1480,N_8099,N_8086);
nand UO_1481 (O_1481,N_9980,N_9390);
nand UO_1482 (O_1482,N_8184,N_8004);
nor UO_1483 (O_1483,N_8769,N_8309);
nor UO_1484 (O_1484,N_8967,N_7965);
nand UO_1485 (O_1485,N_8897,N_9947);
or UO_1486 (O_1486,N_7579,N_8976);
or UO_1487 (O_1487,N_9122,N_9776);
or UO_1488 (O_1488,N_8849,N_8590);
or UO_1489 (O_1489,N_9910,N_8118);
nand UO_1490 (O_1490,N_8624,N_8587);
nor UO_1491 (O_1491,N_8332,N_9007);
or UO_1492 (O_1492,N_9468,N_8513);
or UO_1493 (O_1493,N_9221,N_9614);
nand UO_1494 (O_1494,N_9481,N_8898);
and UO_1495 (O_1495,N_9879,N_9365);
or UO_1496 (O_1496,N_8266,N_8974);
nand UO_1497 (O_1497,N_9046,N_9690);
nor UO_1498 (O_1498,N_9907,N_9075);
and UO_1499 (O_1499,N_7576,N_7998);
endmodule