module basic_1000_10000_1500_4_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_374,In_987);
xnor U1 (N_1,In_567,In_269);
xor U2 (N_2,In_105,In_586);
xor U3 (N_3,In_430,In_727);
nor U4 (N_4,In_553,In_541);
and U5 (N_5,In_484,In_194);
nand U6 (N_6,In_888,In_692);
xnor U7 (N_7,In_811,In_342);
xor U8 (N_8,In_635,In_436);
and U9 (N_9,In_290,In_603);
xor U10 (N_10,In_524,In_85);
nand U11 (N_11,In_417,In_206);
xnor U12 (N_12,In_594,In_490);
nand U13 (N_13,In_893,In_877);
or U14 (N_14,In_247,In_869);
xnor U15 (N_15,In_992,In_701);
nand U16 (N_16,In_421,In_610);
nand U17 (N_17,In_584,In_273);
nor U18 (N_18,In_264,In_621);
and U19 (N_19,In_95,In_467);
nor U20 (N_20,In_11,In_321);
or U21 (N_21,In_155,In_416);
xor U22 (N_22,In_932,In_378);
and U23 (N_23,In_108,In_56);
nor U24 (N_24,In_5,In_402);
nor U25 (N_25,In_880,In_600);
nor U26 (N_26,In_423,In_845);
nand U27 (N_27,In_156,In_400);
and U28 (N_28,In_233,In_881);
or U29 (N_29,In_122,In_179);
and U30 (N_30,In_134,In_32);
xnor U31 (N_31,In_736,In_839);
nor U32 (N_32,In_446,In_577);
nor U33 (N_33,In_817,In_547);
nor U34 (N_34,In_459,In_825);
nand U35 (N_35,In_466,In_98);
xor U36 (N_36,In_173,In_268);
or U37 (N_37,In_746,In_4);
nand U38 (N_38,In_424,In_931);
xnor U39 (N_39,In_818,In_997);
or U40 (N_40,In_868,In_199);
nor U41 (N_41,In_969,In_797);
and U42 (N_42,In_558,In_878);
xor U43 (N_43,In_795,In_219);
or U44 (N_44,In_352,In_734);
or U45 (N_45,In_464,In_136);
xnor U46 (N_46,In_544,In_668);
nor U47 (N_47,In_67,In_760);
and U48 (N_48,In_14,In_562);
nor U49 (N_49,In_961,In_425);
xnor U50 (N_50,In_504,In_815);
and U51 (N_51,In_559,In_10);
nand U52 (N_52,In_353,In_389);
nor U53 (N_53,In_683,In_367);
and U54 (N_54,In_791,In_114);
nand U55 (N_55,In_862,In_226);
nand U56 (N_56,In_783,In_404);
nand U57 (N_57,In_472,In_474);
nor U58 (N_58,In_285,In_415);
or U59 (N_59,In_399,In_560);
or U60 (N_60,In_99,In_958);
and U61 (N_61,In_595,In_437);
nand U62 (N_62,In_677,In_312);
nor U63 (N_63,In_820,In_757);
xnor U64 (N_64,In_836,In_326);
nand U65 (N_65,In_686,In_176);
and U66 (N_66,In_337,In_328);
nor U67 (N_67,In_241,In_171);
xnor U68 (N_68,In_412,In_77);
nand U69 (N_69,In_450,In_742);
nand U70 (N_70,In_261,In_24);
nor U71 (N_71,In_808,In_23);
nor U72 (N_72,In_955,In_468);
or U73 (N_73,In_407,In_934);
nand U74 (N_74,In_491,In_956);
nand U75 (N_75,In_566,In_401);
nand U76 (N_76,In_42,In_609);
nand U77 (N_77,In_385,In_840);
or U78 (N_78,In_585,In_807);
or U79 (N_79,In_605,In_302);
and U80 (N_80,In_952,In_364);
or U81 (N_81,In_715,In_498);
xnor U82 (N_82,In_645,In_118);
xor U83 (N_83,In_887,In_912);
xnor U84 (N_84,In_455,In_111);
and U85 (N_85,In_920,In_202);
and U86 (N_86,In_964,In_422);
nor U87 (N_87,In_255,In_804);
xor U88 (N_88,In_59,In_444);
or U89 (N_89,In_227,In_790);
or U90 (N_90,In_813,In_231);
and U91 (N_91,In_565,In_771);
or U92 (N_92,In_942,In_244);
nand U93 (N_93,In_914,In_348);
xor U94 (N_94,In_475,In_222);
and U95 (N_95,In_922,In_120);
or U96 (N_96,In_165,In_154);
xnor U97 (N_97,In_483,In_220);
or U98 (N_98,In_245,In_403);
xor U99 (N_99,In_162,In_338);
or U100 (N_100,In_230,In_678);
nand U101 (N_101,In_396,In_477);
xnor U102 (N_102,In_188,In_428);
xnor U103 (N_103,In_427,In_236);
or U104 (N_104,In_469,In_993);
nand U105 (N_105,In_274,In_612);
and U106 (N_106,In_270,In_954);
nor U107 (N_107,In_478,In_482);
nor U108 (N_108,In_718,In_685);
and U109 (N_109,In_671,In_83);
nor U110 (N_110,In_267,In_824);
nor U111 (N_111,In_237,In_172);
or U112 (N_112,In_913,In_539);
and U113 (N_113,In_68,In_394);
and U114 (N_114,In_131,In_20);
nor U115 (N_115,In_885,In_616);
and U116 (N_116,In_345,In_849);
nand U117 (N_117,In_251,In_691);
and U118 (N_118,In_370,In_919);
or U119 (N_119,In_725,In_755);
nand U120 (N_120,In_281,In_806);
xor U121 (N_121,In_829,In_960);
nand U122 (N_122,In_810,In_841);
or U123 (N_123,In_842,In_925);
xor U124 (N_124,In_777,In_723);
nor U125 (N_125,In_253,In_679);
nor U126 (N_126,In_589,In_170);
nand U127 (N_127,In_75,In_381);
and U128 (N_128,In_871,In_145);
xor U129 (N_129,In_301,In_709);
or U130 (N_130,In_962,In_340);
and U131 (N_131,In_773,In_69);
nor U132 (N_132,In_397,In_15);
nor U133 (N_133,In_994,In_796);
and U134 (N_134,In_512,In_212);
and U135 (N_135,In_426,In_33);
or U136 (N_136,In_531,In_895);
or U137 (N_137,In_283,In_185);
nand U138 (N_138,In_117,In_58);
or U139 (N_139,In_943,In_159);
xor U140 (N_140,In_722,In_648);
nor U141 (N_141,In_471,In_908);
or U142 (N_142,In_271,In_661);
and U143 (N_143,In_456,In_485);
nor U144 (N_144,In_667,In_789);
and U145 (N_145,In_6,In_707);
xor U146 (N_146,In_322,In_814);
or U147 (N_147,In_545,In_664);
xnor U148 (N_148,In_753,In_160);
and U149 (N_149,In_659,In_666);
nor U150 (N_150,In_240,In_657);
or U151 (N_151,In_758,In_107);
or U152 (N_152,In_699,In_304);
or U153 (N_153,In_1,In_386);
nor U154 (N_154,In_833,In_508);
nor U155 (N_155,In_313,In_556);
or U156 (N_156,In_7,In_537);
and U157 (N_157,In_535,In_182);
nor U158 (N_158,In_163,In_630);
and U159 (N_159,In_435,In_158);
xor U160 (N_160,In_191,In_60);
and U161 (N_161,In_618,In_947);
nand U162 (N_162,In_307,In_63);
xor U163 (N_163,In_768,In_31);
nand U164 (N_164,In_979,In_985);
or U165 (N_165,In_112,In_362);
and U166 (N_166,In_706,In_688);
nor U167 (N_167,In_902,In_133);
xnor U168 (N_168,In_991,In_81);
or U169 (N_169,In_644,In_533);
or U170 (N_170,In_724,In_195);
or U171 (N_171,In_517,In_640);
nand U172 (N_172,In_257,In_26);
xor U173 (N_173,In_384,In_106);
nand U174 (N_174,In_729,In_708);
nand U175 (N_175,In_260,In_147);
and U176 (N_176,In_127,In_897);
nand U177 (N_177,In_102,In_470);
and U178 (N_178,In_637,In_882);
nand U179 (N_179,In_827,In_168);
nor U180 (N_180,In_44,In_324);
nor U181 (N_181,In_792,In_333);
or U182 (N_182,In_900,In_598);
xnor U183 (N_183,In_3,In_363);
nand U184 (N_184,In_971,In_883);
and U185 (N_185,In_809,In_216);
nor U186 (N_186,In_731,In_287);
nor U187 (N_187,In_572,In_816);
nand U188 (N_188,In_583,In_948);
xnor U189 (N_189,In_911,In_702);
or U190 (N_190,In_523,In_295);
xor U191 (N_191,In_988,In_234);
and U192 (N_192,In_534,In_628);
and U193 (N_193,In_905,In_890);
or U194 (N_194,In_607,In_113);
nand U195 (N_195,In_898,In_497);
nand U196 (N_196,In_291,In_747);
nor U197 (N_197,In_892,In_924);
and U198 (N_198,In_970,In_936);
nor U199 (N_199,In_844,In_21);
and U200 (N_200,In_696,In_510);
nand U201 (N_201,In_857,In_332);
and U202 (N_202,In_899,In_999);
nand U203 (N_203,In_513,In_432);
nor U204 (N_204,In_441,In_439);
xnor U205 (N_205,In_479,In_506);
xnor U206 (N_206,In_953,In_292);
and U207 (N_207,In_30,In_61);
or U208 (N_208,In_27,In_97);
or U209 (N_209,In_49,In_681);
nor U210 (N_210,In_55,In_794);
nor U211 (N_211,In_380,In_996);
nand U212 (N_212,In_778,In_859);
nor U213 (N_213,In_488,In_740);
xor U214 (N_214,In_726,In_821);
and U215 (N_215,In_235,In_409);
nand U216 (N_216,In_383,In_779);
nor U217 (N_217,In_481,In_838);
xnor U218 (N_218,In_650,In_100);
nand U219 (N_219,In_769,In_434);
or U220 (N_220,In_141,In_937);
nand U221 (N_221,In_643,In_84);
nand U222 (N_222,In_855,In_655);
and U223 (N_223,In_339,In_476);
nor U224 (N_224,In_354,In_848);
nand U225 (N_225,In_410,In_239);
and U226 (N_226,In_92,In_308);
and U227 (N_227,In_34,In_135);
nand U228 (N_228,In_390,In_80);
nor U229 (N_229,In_907,In_633);
or U230 (N_230,In_774,In_527);
nand U231 (N_231,In_629,In_263);
xor U232 (N_232,In_972,In_940);
or U233 (N_233,In_846,In_798);
and U234 (N_234,In_801,In_528);
nor U235 (N_235,In_288,In_732);
nand U236 (N_236,In_186,In_148);
and U237 (N_237,In_944,In_837);
or U238 (N_238,In_623,In_945);
xnor U239 (N_239,In_254,In_414);
and U240 (N_240,In_502,In_152);
or U241 (N_241,In_453,In_716);
or U242 (N_242,In_359,In_110);
or U243 (N_243,In_178,In_48);
nor U244 (N_244,In_66,In_627);
nand U245 (N_245,In_634,In_856);
and U246 (N_246,In_311,In_826);
nor U247 (N_247,In_300,In_793);
nand U248 (N_248,In_142,In_124);
or U249 (N_249,In_509,In_418);
xor U250 (N_250,In_323,In_754);
or U251 (N_251,In_19,In_903);
nand U252 (N_252,In_876,In_36);
nor U253 (N_253,In_144,In_909);
nor U254 (N_254,In_358,In_90);
or U255 (N_255,In_540,In_543);
xor U256 (N_256,In_64,In_977);
xor U257 (N_257,In_78,In_749);
and U258 (N_258,In_398,In_371);
and U259 (N_259,In_596,In_129);
and U260 (N_260,In_293,In_183);
nand U261 (N_261,In_207,In_554);
or U262 (N_262,In_198,In_73);
nand U263 (N_263,In_587,In_896);
xor U264 (N_264,In_720,In_519);
nor U265 (N_265,In_568,In_721);
xor U266 (N_266,In_344,In_615);
xnor U267 (N_267,In_196,In_756);
and U268 (N_268,In_458,In_43);
nor U269 (N_269,In_980,In_489);
nor U270 (N_270,In_772,In_599);
nand U271 (N_271,In_828,In_682);
and U272 (N_272,In_733,In_50);
and U273 (N_273,In_164,In_984);
or U274 (N_274,In_665,In_486);
and U275 (N_275,In_608,In_652);
xnor U276 (N_276,In_926,In_847);
or U277 (N_277,In_822,In_916);
or U278 (N_278,In_886,In_710);
xor U279 (N_279,In_606,In_590);
xnor U280 (N_280,In_8,In_552);
nor U281 (N_281,In_571,In_939);
nand U282 (N_282,In_904,In_126);
and U283 (N_283,In_711,In_901);
or U284 (N_284,In_576,In_128);
nand U285 (N_285,In_387,In_146);
nor U286 (N_286,In_39,In_713);
nor U287 (N_287,In_581,In_2);
nand U288 (N_288,In_649,In_373);
nor U289 (N_289,In_743,In_306);
or U290 (N_290,In_151,In_800);
and U291 (N_291,In_569,In_918);
or U292 (N_292,In_592,In_325);
nand U293 (N_293,In_203,In_712);
nand U294 (N_294,In_530,In_35);
xor U295 (N_295,In_96,In_157);
xnor U296 (N_296,In_588,In_161);
xnor U297 (N_297,In_787,In_823);
nor U298 (N_298,In_449,In_86);
or U299 (N_299,In_694,In_310);
or U300 (N_300,In_448,In_121);
or U301 (N_301,In_957,In_891);
and U302 (N_302,In_210,In_246);
xnor U303 (N_303,In_275,In_990);
and U304 (N_304,In_770,In_983);
nand U305 (N_305,In_282,In_391);
or U306 (N_306,In_54,In_279);
nor U307 (N_307,In_632,In_884);
xnor U308 (N_308,In_550,In_87);
nor U309 (N_309,In_863,In_376);
or U310 (N_310,In_499,In_580);
nand U311 (N_311,In_631,In_104);
and U312 (N_312,In_366,In_284);
or U313 (N_313,In_115,In_289);
nand U314 (N_314,In_388,In_16);
and U315 (N_315,In_445,In_299);
nor U316 (N_316,In_197,In_45);
nor U317 (N_317,In_548,In_91);
nand U318 (N_318,In_835,In_698);
xnor U319 (N_319,In_213,In_297);
and U320 (N_320,In_329,In_256);
nand U321 (N_321,In_761,In_921);
or U322 (N_322,In_494,In_894);
xor U323 (N_323,In_143,In_174);
xnor U324 (N_324,In_579,In_703);
xnor U325 (N_325,In_258,In_687);
and U326 (N_326,In_201,In_546);
nand U327 (N_327,In_819,In_37);
xor U328 (N_328,In_870,In_465);
nand U329 (N_329,In_38,In_536);
xnor U330 (N_330,In_866,In_315);
xor U331 (N_331,In_763,In_314);
or U332 (N_332,In_626,In_180);
and U333 (N_333,In_433,In_834);
and U334 (N_334,In_693,In_927);
nand U335 (N_335,In_538,In_785);
or U336 (N_336,In_419,In_675);
xnor U337 (N_337,In_343,In_211);
nand U338 (N_338,In_762,In_495);
or U339 (N_339,In_860,In_689);
nor U340 (N_340,In_116,In_70);
nand U341 (N_341,In_356,In_719);
and U342 (N_342,In_831,In_351);
or U343 (N_343,In_94,In_867);
nand U344 (N_344,In_123,In_728);
or U345 (N_345,In_204,In_591);
or U346 (N_346,In_319,In_745);
or U347 (N_347,In_684,In_169);
or U348 (N_348,In_973,In_408);
nor U349 (N_349,In_17,In_9);
nand U350 (N_350,In_874,In_167);
and U351 (N_351,In_741,In_593);
or U352 (N_352,In_420,In_153);
nor U353 (N_353,In_850,In_89);
xor U354 (N_354,In_967,In_624);
and U355 (N_355,In_208,In_906);
nand U356 (N_356,In_974,In_51);
xnor U357 (N_357,In_252,In_109);
nand U358 (N_358,In_177,In_457);
and U359 (N_359,In_872,In_582);
and U360 (N_360,In_636,In_493);
or U361 (N_361,In_74,In_651);
nor U362 (N_362,In_638,In_296);
nand U363 (N_363,In_641,In_205);
nor U364 (N_364,In_654,In_963);
and U365 (N_365,In_413,In_473);
nand U366 (N_366,In_674,In_557);
and U367 (N_367,In_280,In_336);
or U368 (N_368,In_551,In_563);
nand U369 (N_369,In_187,In_959);
or U370 (N_370,In_946,In_786);
xor U371 (N_371,In_656,In_346);
nor U372 (N_372,In_601,In_639);
nand U373 (N_373,In_928,In_739);
xnor U374 (N_374,In_18,In_125);
xnor U375 (N_375,In_697,In_520);
nand U376 (N_376,In_805,In_614);
xor U377 (N_377,In_442,In_132);
nand U378 (N_378,In_975,In_272);
or U379 (N_379,In_864,In_989);
nor U380 (N_380,In_765,In_249);
and U381 (N_381,In_873,In_357);
and U382 (N_382,In_392,In_215);
nand U383 (N_383,In_361,In_46);
or U384 (N_384,In_865,In_737);
nor U385 (N_385,In_752,In_217);
xnor U386 (N_386,In_695,In_47);
nor U387 (N_387,In_347,In_851);
nand U388 (N_388,In_672,In_406);
nor U389 (N_389,In_12,In_889);
nand U390 (N_390,In_65,In_852);
or U391 (N_391,In_330,In_669);
or U392 (N_392,In_748,In_574);
and U393 (N_393,In_209,In_915);
nor U394 (N_394,In_518,In_298);
xor U395 (N_395,In_780,In_149);
nor U396 (N_396,In_830,In_184);
and U397 (N_397,In_611,In_248);
and U398 (N_398,In_526,In_341);
xor U399 (N_399,In_776,In_395);
and U400 (N_400,In_622,In_119);
nand U401 (N_401,In_71,In_318);
and U402 (N_402,In_130,In_62);
and U403 (N_403,In_447,In_788);
xor U404 (N_404,In_57,In_532);
or U405 (N_405,In_923,In_705);
xor U406 (N_406,In_573,In_561);
nor U407 (N_407,In_137,In_744);
nor U408 (N_408,In_79,In_784);
and U409 (N_409,In_294,In_738);
or U410 (N_410,In_843,In_0);
nand U411 (N_411,In_853,In_646);
and U412 (N_412,In_981,In_305);
nor U413 (N_413,In_438,In_858);
nor U414 (N_414,In_735,In_879);
and U415 (N_415,In_138,In_405);
or U416 (N_416,In_714,In_262);
or U417 (N_417,In_181,In_730);
xor U418 (N_418,In_965,In_225);
or U419 (N_419,In_101,In_53);
nor U420 (N_420,In_454,In_515);
or U421 (N_421,In_597,In_750);
and U422 (N_422,In_286,In_501);
and U423 (N_423,In_349,In_369);
and U424 (N_424,In_647,In_620);
nand U425 (N_425,In_982,In_28);
nor U426 (N_426,In_480,In_22);
and U427 (N_427,In_662,In_511);
and U428 (N_428,In_670,In_452);
and U429 (N_429,In_917,In_492);
nand U430 (N_430,In_335,In_461);
xnor U431 (N_431,In_998,In_832);
or U432 (N_432,In_372,In_193);
or U433 (N_433,In_375,In_625);
nand U434 (N_434,In_500,In_229);
nor U435 (N_435,In_379,In_224);
or U436 (N_436,In_575,In_463);
xnor U437 (N_437,In_764,In_52);
and U438 (N_438,In_250,In_976);
nand U439 (N_439,In_192,In_658);
nor U440 (N_440,In_767,In_929);
nand U441 (N_441,In_910,In_411);
nor U442 (N_442,In_516,In_334);
or U443 (N_443,In_242,In_232);
nor U444 (N_444,In_443,In_542);
and U445 (N_445,In_503,In_570);
and U446 (N_446,In_189,In_941);
or U447 (N_447,In_175,In_303);
xnor U448 (N_448,In_995,In_496);
nand U449 (N_449,In_41,In_660);
nor U450 (N_450,In_700,In_803);
and U451 (N_451,In_781,In_653);
nand U452 (N_452,In_13,In_949);
xor U453 (N_453,In_214,In_619);
nor U454 (N_454,In_799,In_29);
nand U455 (N_455,In_525,In_522);
nand U456 (N_456,In_440,In_382);
xor U457 (N_457,In_166,In_316);
and U458 (N_458,In_40,In_968);
nand U459 (N_459,In_564,In_951);
nor U460 (N_460,In_393,In_320);
xnor U461 (N_461,In_72,In_266);
xnor U462 (N_462,In_875,In_317);
and U463 (N_463,In_854,In_529);
or U464 (N_464,In_617,In_676);
nand U465 (N_465,In_223,In_429);
or U466 (N_466,In_150,In_82);
nor U467 (N_467,In_704,In_986);
nand U468 (N_468,In_613,In_680);
nor U469 (N_469,In_930,In_238);
xnor U470 (N_470,In_978,In_451);
nor U471 (N_471,In_782,In_462);
and U472 (N_472,In_690,In_139);
or U473 (N_473,In_766,In_368);
and U474 (N_474,In_331,In_276);
and U475 (N_475,In_861,In_717);
or U476 (N_476,In_938,In_140);
nand U477 (N_477,In_812,In_759);
nor U478 (N_478,In_243,In_365);
or U479 (N_479,In_218,In_103);
and U480 (N_480,In_505,In_76);
xnor U481 (N_481,In_93,In_350);
and U482 (N_482,In_309,In_514);
or U483 (N_483,In_460,In_935);
or U484 (N_484,In_487,In_933);
xnor U485 (N_485,In_377,In_25);
nand U486 (N_486,In_555,In_604);
nand U487 (N_487,In_578,In_549);
or U488 (N_488,In_966,In_88);
nand U489 (N_489,In_360,In_950);
or U490 (N_490,In_259,In_228);
and U491 (N_491,In_663,In_507);
and U492 (N_492,In_642,In_278);
and U493 (N_493,In_327,In_775);
or U494 (N_494,In_431,In_200);
nand U495 (N_495,In_277,In_190);
xor U496 (N_496,In_265,In_602);
or U497 (N_497,In_521,In_751);
xnor U498 (N_498,In_802,In_221);
or U499 (N_499,In_355,In_673);
xor U500 (N_500,In_102,In_153);
or U501 (N_501,In_608,In_600);
xor U502 (N_502,In_507,In_615);
or U503 (N_503,In_344,In_802);
nand U504 (N_504,In_662,In_319);
nand U505 (N_505,In_353,In_899);
xnor U506 (N_506,In_968,In_627);
nor U507 (N_507,In_879,In_555);
xor U508 (N_508,In_939,In_735);
nand U509 (N_509,In_370,In_994);
nor U510 (N_510,In_487,In_988);
xor U511 (N_511,In_967,In_731);
xnor U512 (N_512,In_710,In_543);
xor U513 (N_513,In_59,In_65);
nor U514 (N_514,In_528,In_256);
or U515 (N_515,In_957,In_784);
nand U516 (N_516,In_524,In_727);
nor U517 (N_517,In_26,In_66);
and U518 (N_518,In_258,In_900);
or U519 (N_519,In_635,In_546);
and U520 (N_520,In_988,In_118);
and U521 (N_521,In_232,In_297);
and U522 (N_522,In_394,In_635);
and U523 (N_523,In_72,In_198);
nand U524 (N_524,In_343,In_697);
and U525 (N_525,In_175,In_592);
nor U526 (N_526,In_719,In_477);
nand U527 (N_527,In_927,In_801);
or U528 (N_528,In_550,In_257);
xor U529 (N_529,In_694,In_18);
or U530 (N_530,In_193,In_899);
and U531 (N_531,In_54,In_924);
or U532 (N_532,In_611,In_550);
nand U533 (N_533,In_866,In_743);
nor U534 (N_534,In_570,In_349);
nand U535 (N_535,In_509,In_974);
or U536 (N_536,In_856,In_619);
nand U537 (N_537,In_93,In_689);
xnor U538 (N_538,In_150,In_775);
or U539 (N_539,In_714,In_954);
and U540 (N_540,In_495,In_882);
or U541 (N_541,In_605,In_731);
and U542 (N_542,In_594,In_310);
nand U543 (N_543,In_824,In_272);
and U544 (N_544,In_286,In_203);
and U545 (N_545,In_338,In_703);
and U546 (N_546,In_873,In_442);
xor U547 (N_547,In_93,In_409);
or U548 (N_548,In_871,In_296);
or U549 (N_549,In_907,In_143);
nand U550 (N_550,In_186,In_281);
nand U551 (N_551,In_860,In_920);
xor U552 (N_552,In_463,In_935);
nor U553 (N_553,In_814,In_58);
nor U554 (N_554,In_139,In_456);
xnor U555 (N_555,In_256,In_356);
nand U556 (N_556,In_835,In_934);
xor U557 (N_557,In_198,In_217);
and U558 (N_558,In_431,In_179);
xor U559 (N_559,In_681,In_823);
nor U560 (N_560,In_749,In_14);
or U561 (N_561,In_896,In_726);
and U562 (N_562,In_264,In_210);
and U563 (N_563,In_612,In_736);
or U564 (N_564,In_564,In_11);
nand U565 (N_565,In_568,In_167);
xor U566 (N_566,In_863,In_48);
xor U567 (N_567,In_431,In_880);
nand U568 (N_568,In_455,In_586);
nand U569 (N_569,In_909,In_140);
or U570 (N_570,In_810,In_507);
xor U571 (N_571,In_290,In_218);
nor U572 (N_572,In_261,In_631);
xor U573 (N_573,In_771,In_396);
nand U574 (N_574,In_745,In_482);
and U575 (N_575,In_550,In_337);
nor U576 (N_576,In_76,In_981);
xnor U577 (N_577,In_56,In_684);
nor U578 (N_578,In_221,In_363);
nand U579 (N_579,In_677,In_799);
or U580 (N_580,In_19,In_392);
nand U581 (N_581,In_659,In_203);
xor U582 (N_582,In_803,In_201);
nor U583 (N_583,In_904,In_10);
or U584 (N_584,In_313,In_269);
nand U585 (N_585,In_922,In_763);
or U586 (N_586,In_157,In_899);
nor U587 (N_587,In_990,In_852);
nor U588 (N_588,In_732,In_186);
xor U589 (N_589,In_169,In_465);
nand U590 (N_590,In_63,In_944);
and U591 (N_591,In_996,In_254);
and U592 (N_592,In_519,In_935);
and U593 (N_593,In_558,In_673);
xor U594 (N_594,In_365,In_236);
nand U595 (N_595,In_689,In_409);
xor U596 (N_596,In_584,In_39);
nor U597 (N_597,In_537,In_792);
nand U598 (N_598,In_442,In_623);
nor U599 (N_599,In_658,In_450);
nand U600 (N_600,In_382,In_413);
nor U601 (N_601,In_24,In_23);
or U602 (N_602,In_916,In_629);
xor U603 (N_603,In_202,In_790);
xnor U604 (N_604,In_602,In_354);
xor U605 (N_605,In_848,In_536);
and U606 (N_606,In_197,In_904);
xnor U607 (N_607,In_373,In_451);
xnor U608 (N_608,In_676,In_540);
or U609 (N_609,In_399,In_863);
nand U610 (N_610,In_675,In_30);
and U611 (N_611,In_532,In_756);
or U612 (N_612,In_593,In_988);
xnor U613 (N_613,In_711,In_410);
nand U614 (N_614,In_8,In_324);
xnor U615 (N_615,In_884,In_10);
nor U616 (N_616,In_438,In_167);
or U617 (N_617,In_847,In_277);
or U618 (N_618,In_246,In_376);
or U619 (N_619,In_744,In_43);
xnor U620 (N_620,In_407,In_586);
xor U621 (N_621,In_133,In_844);
xor U622 (N_622,In_491,In_278);
nand U623 (N_623,In_722,In_401);
nor U624 (N_624,In_195,In_934);
and U625 (N_625,In_45,In_750);
nor U626 (N_626,In_132,In_59);
nor U627 (N_627,In_88,In_381);
and U628 (N_628,In_512,In_787);
nand U629 (N_629,In_705,In_70);
or U630 (N_630,In_501,In_536);
or U631 (N_631,In_425,In_84);
xnor U632 (N_632,In_746,In_121);
xnor U633 (N_633,In_170,In_494);
nor U634 (N_634,In_297,In_573);
or U635 (N_635,In_539,In_715);
nand U636 (N_636,In_755,In_153);
and U637 (N_637,In_250,In_477);
xnor U638 (N_638,In_235,In_698);
nand U639 (N_639,In_316,In_985);
nor U640 (N_640,In_298,In_65);
nor U641 (N_641,In_482,In_729);
nand U642 (N_642,In_250,In_639);
nand U643 (N_643,In_166,In_368);
and U644 (N_644,In_1,In_681);
nand U645 (N_645,In_776,In_55);
or U646 (N_646,In_860,In_598);
or U647 (N_647,In_285,In_526);
nor U648 (N_648,In_659,In_518);
nor U649 (N_649,In_764,In_187);
nand U650 (N_650,In_773,In_18);
or U651 (N_651,In_522,In_169);
nand U652 (N_652,In_216,In_737);
nor U653 (N_653,In_744,In_118);
nor U654 (N_654,In_411,In_395);
or U655 (N_655,In_30,In_557);
nor U656 (N_656,In_25,In_407);
nor U657 (N_657,In_992,In_653);
or U658 (N_658,In_772,In_487);
nand U659 (N_659,In_517,In_243);
nand U660 (N_660,In_581,In_485);
xnor U661 (N_661,In_126,In_729);
or U662 (N_662,In_875,In_737);
and U663 (N_663,In_686,In_474);
xor U664 (N_664,In_619,In_395);
and U665 (N_665,In_410,In_138);
or U666 (N_666,In_466,In_196);
xnor U667 (N_667,In_150,In_275);
or U668 (N_668,In_545,In_575);
nand U669 (N_669,In_406,In_549);
or U670 (N_670,In_732,In_242);
xor U671 (N_671,In_711,In_274);
nor U672 (N_672,In_620,In_503);
nor U673 (N_673,In_133,In_976);
xor U674 (N_674,In_214,In_150);
or U675 (N_675,In_742,In_311);
nor U676 (N_676,In_764,In_299);
nor U677 (N_677,In_373,In_208);
xnor U678 (N_678,In_51,In_539);
and U679 (N_679,In_111,In_936);
nor U680 (N_680,In_633,In_776);
nor U681 (N_681,In_663,In_349);
nor U682 (N_682,In_852,In_576);
and U683 (N_683,In_940,In_401);
nand U684 (N_684,In_259,In_982);
xnor U685 (N_685,In_325,In_438);
nor U686 (N_686,In_823,In_330);
xnor U687 (N_687,In_449,In_649);
nand U688 (N_688,In_946,In_609);
xnor U689 (N_689,In_225,In_856);
or U690 (N_690,In_362,In_285);
xnor U691 (N_691,In_773,In_64);
nor U692 (N_692,In_107,In_197);
or U693 (N_693,In_586,In_707);
nand U694 (N_694,In_731,In_134);
nand U695 (N_695,In_212,In_504);
and U696 (N_696,In_121,In_713);
nand U697 (N_697,In_153,In_509);
or U698 (N_698,In_776,In_763);
or U699 (N_699,In_231,In_654);
nand U700 (N_700,In_697,In_47);
nand U701 (N_701,In_836,In_458);
nand U702 (N_702,In_140,In_521);
or U703 (N_703,In_423,In_45);
nor U704 (N_704,In_154,In_357);
nor U705 (N_705,In_645,In_828);
nor U706 (N_706,In_891,In_505);
xnor U707 (N_707,In_357,In_801);
or U708 (N_708,In_278,In_254);
xnor U709 (N_709,In_644,In_128);
and U710 (N_710,In_664,In_202);
and U711 (N_711,In_717,In_767);
nand U712 (N_712,In_912,In_144);
xnor U713 (N_713,In_941,In_656);
xnor U714 (N_714,In_344,In_287);
or U715 (N_715,In_326,In_708);
or U716 (N_716,In_505,In_773);
nand U717 (N_717,In_91,In_985);
and U718 (N_718,In_600,In_227);
or U719 (N_719,In_213,In_964);
nand U720 (N_720,In_339,In_918);
nand U721 (N_721,In_460,In_828);
or U722 (N_722,In_445,In_74);
and U723 (N_723,In_547,In_695);
xor U724 (N_724,In_99,In_241);
xor U725 (N_725,In_175,In_634);
xor U726 (N_726,In_990,In_346);
xor U727 (N_727,In_998,In_133);
xor U728 (N_728,In_423,In_279);
nor U729 (N_729,In_413,In_742);
nor U730 (N_730,In_441,In_528);
and U731 (N_731,In_167,In_921);
or U732 (N_732,In_30,In_332);
nand U733 (N_733,In_652,In_590);
nand U734 (N_734,In_604,In_230);
and U735 (N_735,In_786,In_825);
xor U736 (N_736,In_217,In_243);
and U737 (N_737,In_763,In_176);
nor U738 (N_738,In_426,In_600);
xnor U739 (N_739,In_815,In_844);
xor U740 (N_740,In_183,In_754);
xnor U741 (N_741,In_771,In_213);
xor U742 (N_742,In_456,In_428);
nand U743 (N_743,In_796,In_661);
nand U744 (N_744,In_629,In_368);
and U745 (N_745,In_631,In_470);
nor U746 (N_746,In_787,In_963);
or U747 (N_747,In_862,In_1);
nand U748 (N_748,In_820,In_956);
nand U749 (N_749,In_273,In_355);
or U750 (N_750,In_539,In_367);
or U751 (N_751,In_893,In_704);
or U752 (N_752,In_355,In_917);
and U753 (N_753,In_856,In_764);
xor U754 (N_754,In_53,In_166);
and U755 (N_755,In_31,In_154);
nand U756 (N_756,In_443,In_576);
nor U757 (N_757,In_832,In_608);
xnor U758 (N_758,In_739,In_449);
nand U759 (N_759,In_256,In_574);
or U760 (N_760,In_978,In_962);
or U761 (N_761,In_26,In_642);
nand U762 (N_762,In_681,In_730);
and U763 (N_763,In_120,In_711);
nand U764 (N_764,In_135,In_741);
xnor U765 (N_765,In_230,In_528);
or U766 (N_766,In_880,In_553);
and U767 (N_767,In_892,In_18);
or U768 (N_768,In_273,In_271);
nor U769 (N_769,In_838,In_669);
and U770 (N_770,In_626,In_592);
nor U771 (N_771,In_834,In_644);
xor U772 (N_772,In_652,In_494);
and U773 (N_773,In_735,In_297);
xor U774 (N_774,In_984,In_669);
or U775 (N_775,In_168,In_467);
nor U776 (N_776,In_462,In_515);
nor U777 (N_777,In_430,In_758);
nand U778 (N_778,In_53,In_340);
xnor U779 (N_779,In_557,In_996);
and U780 (N_780,In_24,In_758);
or U781 (N_781,In_344,In_259);
and U782 (N_782,In_622,In_86);
nor U783 (N_783,In_161,In_174);
nor U784 (N_784,In_255,In_407);
or U785 (N_785,In_618,In_314);
and U786 (N_786,In_985,In_532);
nor U787 (N_787,In_610,In_575);
nand U788 (N_788,In_212,In_309);
nand U789 (N_789,In_387,In_759);
and U790 (N_790,In_428,In_646);
or U791 (N_791,In_115,In_357);
nand U792 (N_792,In_529,In_766);
and U793 (N_793,In_144,In_123);
and U794 (N_794,In_611,In_115);
nand U795 (N_795,In_129,In_689);
nor U796 (N_796,In_339,In_252);
and U797 (N_797,In_855,In_615);
xor U798 (N_798,In_450,In_775);
nand U799 (N_799,In_158,In_961);
or U800 (N_800,In_435,In_346);
xnor U801 (N_801,In_875,In_739);
xor U802 (N_802,In_194,In_336);
xnor U803 (N_803,In_460,In_674);
or U804 (N_804,In_535,In_775);
nor U805 (N_805,In_15,In_33);
nor U806 (N_806,In_960,In_473);
nor U807 (N_807,In_32,In_18);
and U808 (N_808,In_424,In_975);
xor U809 (N_809,In_115,In_808);
nor U810 (N_810,In_381,In_816);
or U811 (N_811,In_499,In_303);
or U812 (N_812,In_895,In_313);
nor U813 (N_813,In_760,In_521);
xnor U814 (N_814,In_266,In_436);
xnor U815 (N_815,In_876,In_661);
or U816 (N_816,In_618,In_193);
or U817 (N_817,In_409,In_695);
nor U818 (N_818,In_466,In_24);
xnor U819 (N_819,In_682,In_46);
xor U820 (N_820,In_535,In_713);
nor U821 (N_821,In_749,In_411);
or U822 (N_822,In_121,In_895);
or U823 (N_823,In_542,In_824);
nand U824 (N_824,In_789,In_244);
nor U825 (N_825,In_181,In_632);
nand U826 (N_826,In_728,In_997);
nand U827 (N_827,In_848,In_835);
and U828 (N_828,In_629,In_488);
xor U829 (N_829,In_668,In_343);
nand U830 (N_830,In_896,In_452);
and U831 (N_831,In_331,In_159);
and U832 (N_832,In_277,In_544);
nor U833 (N_833,In_560,In_839);
nand U834 (N_834,In_515,In_851);
and U835 (N_835,In_136,In_623);
xnor U836 (N_836,In_351,In_821);
xnor U837 (N_837,In_475,In_105);
xnor U838 (N_838,In_581,In_818);
and U839 (N_839,In_851,In_462);
nand U840 (N_840,In_88,In_871);
and U841 (N_841,In_49,In_383);
nor U842 (N_842,In_143,In_583);
and U843 (N_843,In_519,In_659);
xnor U844 (N_844,In_833,In_981);
xnor U845 (N_845,In_452,In_435);
and U846 (N_846,In_806,In_282);
and U847 (N_847,In_865,In_26);
nand U848 (N_848,In_504,In_164);
xnor U849 (N_849,In_302,In_357);
nand U850 (N_850,In_809,In_631);
nand U851 (N_851,In_69,In_636);
xnor U852 (N_852,In_957,In_824);
xnor U853 (N_853,In_753,In_881);
nand U854 (N_854,In_550,In_763);
xor U855 (N_855,In_326,In_465);
or U856 (N_856,In_351,In_827);
and U857 (N_857,In_668,In_391);
nand U858 (N_858,In_660,In_366);
xnor U859 (N_859,In_824,In_606);
and U860 (N_860,In_794,In_829);
and U861 (N_861,In_766,In_98);
nand U862 (N_862,In_84,In_971);
and U863 (N_863,In_973,In_804);
nor U864 (N_864,In_990,In_687);
and U865 (N_865,In_636,In_316);
nand U866 (N_866,In_587,In_376);
xnor U867 (N_867,In_134,In_926);
nand U868 (N_868,In_251,In_470);
xnor U869 (N_869,In_881,In_721);
xnor U870 (N_870,In_3,In_905);
xnor U871 (N_871,In_369,In_449);
nor U872 (N_872,In_380,In_313);
and U873 (N_873,In_791,In_635);
and U874 (N_874,In_144,In_141);
xor U875 (N_875,In_79,In_729);
xor U876 (N_876,In_429,In_250);
nor U877 (N_877,In_556,In_426);
and U878 (N_878,In_677,In_654);
xor U879 (N_879,In_146,In_807);
nand U880 (N_880,In_561,In_668);
nand U881 (N_881,In_376,In_332);
and U882 (N_882,In_140,In_686);
nor U883 (N_883,In_560,In_585);
nor U884 (N_884,In_8,In_275);
or U885 (N_885,In_362,In_341);
or U886 (N_886,In_195,In_558);
nor U887 (N_887,In_879,In_240);
xnor U888 (N_888,In_453,In_353);
or U889 (N_889,In_804,In_894);
or U890 (N_890,In_904,In_327);
and U891 (N_891,In_589,In_640);
nor U892 (N_892,In_285,In_887);
xnor U893 (N_893,In_193,In_726);
and U894 (N_894,In_14,In_781);
nand U895 (N_895,In_767,In_299);
nand U896 (N_896,In_933,In_979);
xnor U897 (N_897,In_376,In_700);
and U898 (N_898,In_499,In_892);
nand U899 (N_899,In_833,In_990);
nand U900 (N_900,In_640,In_408);
nand U901 (N_901,In_306,In_151);
nand U902 (N_902,In_884,In_871);
xor U903 (N_903,In_285,In_407);
or U904 (N_904,In_636,In_73);
or U905 (N_905,In_965,In_351);
or U906 (N_906,In_128,In_351);
and U907 (N_907,In_4,In_348);
xor U908 (N_908,In_949,In_90);
nand U909 (N_909,In_429,In_987);
or U910 (N_910,In_542,In_483);
and U911 (N_911,In_388,In_877);
nand U912 (N_912,In_227,In_570);
nand U913 (N_913,In_928,In_22);
or U914 (N_914,In_465,In_7);
and U915 (N_915,In_251,In_310);
nor U916 (N_916,In_723,In_895);
nand U917 (N_917,In_952,In_663);
nand U918 (N_918,In_933,In_907);
and U919 (N_919,In_551,In_585);
nand U920 (N_920,In_800,In_237);
and U921 (N_921,In_840,In_209);
xor U922 (N_922,In_190,In_426);
nor U923 (N_923,In_870,In_929);
xor U924 (N_924,In_613,In_268);
xor U925 (N_925,In_619,In_206);
and U926 (N_926,In_648,In_229);
nor U927 (N_927,In_766,In_911);
nand U928 (N_928,In_872,In_427);
and U929 (N_929,In_138,In_968);
nor U930 (N_930,In_249,In_91);
xor U931 (N_931,In_895,In_463);
or U932 (N_932,In_790,In_759);
nor U933 (N_933,In_149,In_335);
and U934 (N_934,In_427,In_474);
and U935 (N_935,In_622,In_3);
xnor U936 (N_936,In_201,In_687);
xor U937 (N_937,In_589,In_519);
xor U938 (N_938,In_519,In_549);
or U939 (N_939,In_498,In_380);
nor U940 (N_940,In_908,In_219);
or U941 (N_941,In_683,In_719);
and U942 (N_942,In_689,In_707);
nor U943 (N_943,In_127,In_752);
nand U944 (N_944,In_947,In_511);
and U945 (N_945,In_150,In_862);
nor U946 (N_946,In_69,In_776);
nand U947 (N_947,In_334,In_195);
xor U948 (N_948,In_84,In_481);
xor U949 (N_949,In_400,In_174);
and U950 (N_950,In_684,In_706);
nor U951 (N_951,In_454,In_248);
nand U952 (N_952,In_131,In_296);
xnor U953 (N_953,In_970,In_815);
or U954 (N_954,In_455,In_251);
and U955 (N_955,In_448,In_870);
and U956 (N_956,In_309,In_49);
xor U957 (N_957,In_831,In_528);
and U958 (N_958,In_176,In_768);
nor U959 (N_959,In_664,In_58);
nor U960 (N_960,In_792,In_796);
and U961 (N_961,In_475,In_179);
nor U962 (N_962,In_59,In_307);
or U963 (N_963,In_956,In_895);
xnor U964 (N_964,In_522,In_916);
nand U965 (N_965,In_383,In_885);
nand U966 (N_966,In_506,In_694);
and U967 (N_967,In_726,In_231);
xor U968 (N_968,In_564,In_775);
or U969 (N_969,In_778,In_554);
xnor U970 (N_970,In_189,In_753);
xor U971 (N_971,In_379,In_969);
nand U972 (N_972,In_280,In_115);
xor U973 (N_973,In_886,In_308);
xnor U974 (N_974,In_407,In_534);
nor U975 (N_975,In_968,In_444);
nor U976 (N_976,In_425,In_679);
and U977 (N_977,In_491,In_365);
and U978 (N_978,In_608,In_34);
or U979 (N_979,In_475,In_967);
nand U980 (N_980,In_42,In_611);
or U981 (N_981,In_566,In_104);
and U982 (N_982,In_542,In_444);
nor U983 (N_983,In_135,In_403);
and U984 (N_984,In_359,In_980);
nand U985 (N_985,In_847,In_563);
xor U986 (N_986,In_877,In_635);
nand U987 (N_987,In_700,In_544);
nand U988 (N_988,In_477,In_294);
xor U989 (N_989,In_312,In_787);
xor U990 (N_990,In_44,In_353);
or U991 (N_991,In_28,In_537);
or U992 (N_992,In_617,In_784);
and U993 (N_993,In_25,In_231);
xor U994 (N_994,In_62,In_540);
nor U995 (N_995,In_370,In_75);
nor U996 (N_996,In_320,In_719);
or U997 (N_997,In_184,In_436);
nor U998 (N_998,In_213,In_188);
nor U999 (N_999,In_813,In_884);
nand U1000 (N_1000,In_99,In_360);
or U1001 (N_1001,In_342,In_326);
and U1002 (N_1002,In_606,In_46);
or U1003 (N_1003,In_555,In_421);
nand U1004 (N_1004,In_200,In_671);
or U1005 (N_1005,In_985,In_577);
xor U1006 (N_1006,In_202,In_417);
xnor U1007 (N_1007,In_248,In_469);
and U1008 (N_1008,In_813,In_213);
and U1009 (N_1009,In_529,In_830);
or U1010 (N_1010,In_377,In_162);
xor U1011 (N_1011,In_523,In_831);
nor U1012 (N_1012,In_924,In_55);
and U1013 (N_1013,In_347,In_81);
or U1014 (N_1014,In_632,In_670);
and U1015 (N_1015,In_612,In_921);
nand U1016 (N_1016,In_525,In_765);
or U1017 (N_1017,In_920,In_276);
nand U1018 (N_1018,In_858,In_667);
xnor U1019 (N_1019,In_6,In_726);
xor U1020 (N_1020,In_899,In_29);
nor U1021 (N_1021,In_489,In_458);
or U1022 (N_1022,In_399,In_638);
xnor U1023 (N_1023,In_523,In_909);
xnor U1024 (N_1024,In_427,In_490);
nand U1025 (N_1025,In_482,In_231);
nor U1026 (N_1026,In_232,In_445);
nor U1027 (N_1027,In_419,In_240);
or U1028 (N_1028,In_272,In_803);
xor U1029 (N_1029,In_886,In_443);
and U1030 (N_1030,In_353,In_331);
or U1031 (N_1031,In_632,In_826);
nand U1032 (N_1032,In_491,In_685);
nor U1033 (N_1033,In_915,In_681);
nor U1034 (N_1034,In_872,In_79);
or U1035 (N_1035,In_883,In_291);
and U1036 (N_1036,In_412,In_575);
nand U1037 (N_1037,In_587,In_207);
xor U1038 (N_1038,In_721,In_175);
and U1039 (N_1039,In_349,In_49);
nor U1040 (N_1040,In_928,In_931);
nor U1041 (N_1041,In_614,In_809);
nor U1042 (N_1042,In_507,In_759);
and U1043 (N_1043,In_681,In_624);
or U1044 (N_1044,In_239,In_193);
nand U1045 (N_1045,In_605,In_308);
or U1046 (N_1046,In_369,In_674);
xor U1047 (N_1047,In_190,In_998);
xor U1048 (N_1048,In_362,In_173);
nor U1049 (N_1049,In_278,In_124);
and U1050 (N_1050,In_970,In_120);
and U1051 (N_1051,In_881,In_202);
nor U1052 (N_1052,In_448,In_69);
xor U1053 (N_1053,In_509,In_401);
xor U1054 (N_1054,In_519,In_407);
and U1055 (N_1055,In_676,In_306);
nand U1056 (N_1056,In_495,In_554);
or U1057 (N_1057,In_300,In_916);
nor U1058 (N_1058,In_369,In_203);
nand U1059 (N_1059,In_947,In_835);
and U1060 (N_1060,In_821,In_755);
xor U1061 (N_1061,In_90,In_271);
nand U1062 (N_1062,In_973,In_306);
nor U1063 (N_1063,In_316,In_216);
or U1064 (N_1064,In_128,In_317);
nand U1065 (N_1065,In_910,In_844);
or U1066 (N_1066,In_339,In_197);
nand U1067 (N_1067,In_261,In_433);
and U1068 (N_1068,In_593,In_882);
nand U1069 (N_1069,In_460,In_549);
or U1070 (N_1070,In_660,In_32);
and U1071 (N_1071,In_521,In_900);
or U1072 (N_1072,In_491,In_306);
nor U1073 (N_1073,In_129,In_671);
nor U1074 (N_1074,In_814,In_826);
xor U1075 (N_1075,In_767,In_127);
nand U1076 (N_1076,In_732,In_96);
nor U1077 (N_1077,In_969,In_527);
xor U1078 (N_1078,In_926,In_999);
or U1079 (N_1079,In_898,In_936);
xnor U1080 (N_1080,In_566,In_377);
or U1081 (N_1081,In_960,In_983);
or U1082 (N_1082,In_496,In_121);
xnor U1083 (N_1083,In_370,In_449);
or U1084 (N_1084,In_335,In_563);
xnor U1085 (N_1085,In_216,In_666);
and U1086 (N_1086,In_807,In_168);
and U1087 (N_1087,In_968,In_972);
xor U1088 (N_1088,In_343,In_371);
nand U1089 (N_1089,In_414,In_130);
nor U1090 (N_1090,In_572,In_240);
and U1091 (N_1091,In_514,In_278);
and U1092 (N_1092,In_400,In_534);
nand U1093 (N_1093,In_59,In_971);
nand U1094 (N_1094,In_784,In_763);
nor U1095 (N_1095,In_29,In_525);
and U1096 (N_1096,In_428,In_759);
xor U1097 (N_1097,In_1,In_599);
xnor U1098 (N_1098,In_345,In_325);
nand U1099 (N_1099,In_289,In_615);
and U1100 (N_1100,In_888,In_158);
or U1101 (N_1101,In_42,In_404);
or U1102 (N_1102,In_883,In_393);
or U1103 (N_1103,In_46,In_698);
nor U1104 (N_1104,In_271,In_84);
xor U1105 (N_1105,In_59,In_695);
and U1106 (N_1106,In_830,In_163);
or U1107 (N_1107,In_567,In_412);
and U1108 (N_1108,In_72,In_975);
and U1109 (N_1109,In_248,In_766);
nor U1110 (N_1110,In_652,In_100);
or U1111 (N_1111,In_105,In_55);
xnor U1112 (N_1112,In_418,In_192);
nand U1113 (N_1113,In_403,In_163);
or U1114 (N_1114,In_951,In_852);
nor U1115 (N_1115,In_143,In_294);
nor U1116 (N_1116,In_371,In_884);
or U1117 (N_1117,In_102,In_206);
nor U1118 (N_1118,In_806,In_38);
nand U1119 (N_1119,In_56,In_382);
nand U1120 (N_1120,In_722,In_113);
nor U1121 (N_1121,In_731,In_40);
or U1122 (N_1122,In_903,In_368);
or U1123 (N_1123,In_74,In_841);
xor U1124 (N_1124,In_395,In_326);
nand U1125 (N_1125,In_846,In_145);
nor U1126 (N_1126,In_18,In_522);
and U1127 (N_1127,In_976,In_525);
xnor U1128 (N_1128,In_205,In_450);
nand U1129 (N_1129,In_940,In_81);
xor U1130 (N_1130,In_204,In_289);
and U1131 (N_1131,In_917,In_51);
xnor U1132 (N_1132,In_149,In_281);
nand U1133 (N_1133,In_657,In_355);
xor U1134 (N_1134,In_433,In_508);
nand U1135 (N_1135,In_267,In_810);
nand U1136 (N_1136,In_150,In_743);
xnor U1137 (N_1137,In_399,In_641);
nand U1138 (N_1138,In_279,In_593);
nor U1139 (N_1139,In_69,In_21);
nand U1140 (N_1140,In_909,In_373);
xnor U1141 (N_1141,In_203,In_478);
and U1142 (N_1142,In_477,In_160);
nor U1143 (N_1143,In_761,In_109);
and U1144 (N_1144,In_923,In_697);
xnor U1145 (N_1145,In_772,In_471);
nor U1146 (N_1146,In_689,In_612);
nand U1147 (N_1147,In_495,In_672);
xor U1148 (N_1148,In_393,In_151);
xor U1149 (N_1149,In_833,In_634);
nand U1150 (N_1150,In_495,In_492);
or U1151 (N_1151,In_561,In_438);
or U1152 (N_1152,In_287,In_622);
and U1153 (N_1153,In_411,In_350);
and U1154 (N_1154,In_656,In_561);
nor U1155 (N_1155,In_416,In_448);
xor U1156 (N_1156,In_429,In_999);
or U1157 (N_1157,In_295,In_537);
or U1158 (N_1158,In_767,In_345);
nand U1159 (N_1159,In_60,In_91);
nand U1160 (N_1160,In_79,In_54);
nor U1161 (N_1161,In_737,In_412);
nand U1162 (N_1162,In_591,In_273);
nand U1163 (N_1163,In_654,In_341);
nor U1164 (N_1164,In_286,In_204);
or U1165 (N_1165,In_394,In_288);
and U1166 (N_1166,In_650,In_505);
xor U1167 (N_1167,In_498,In_930);
or U1168 (N_1168,In_888,In_402);
nor U1169 (N_1169,In_747,In_878);
and U1170 (N_1170,In_851,In_633);
or U1171 (N_1171,In_992,In_47);
xnor U1172 (N_1172,In_86,In_933);
nor U1173 (N_1173,In_531,In_653);
nand U1174 (N_1174,In_846,In_94);
nor U1175 (N_1175,In_921,In_770);
or U1176 (N_1176,In_387,In_807);
or U1177 (N_1177,In_721,In_111);
or U1178 (N_1178,In_708,In_222);
nor U1179 (N_1179,In_350,In_321);
nand U1180 (N_1180,In_64,In_897);
nor U1181 (N_1181,In_157,In_537);
xor U1182 (N_1182,In_105,In_340);
and U1183 (N_1183,In_167,In_474);
or U1184 (N_1184,In_774,In_458);
nor U1185 (N_1185,In_261,In_412);
nand U1186 (N_1186,In_249,In_894);
nand U1187 (N_1187,In_131,In_78);
nor U1188 (N_1188,In_102,In_676);
and U1189 (N_1189,In_788,In_551);
and U1190 (N_1190,In_341,In_477);
or U1191 (N_1191,In_994,In_530);
and U1192 (N_1192,In_77,In_723);
and U1193 (N_1193,In_953,In_117);
or U1194 (N_1194,In_912,In_889);
nor U1195 (N_1195,In_410,In_700);
nor U1196 (N_1196,In_132,In_149);
nand U1197 (N_1197,In_706,In_306);
nand U1198 (N_1198,In_336,In_721);
xnor U1199 (N_1199,In_347,In_441);
or U1200 (N_1200,In_913,In_376);
xor U1201 (N_1201,In_453,In_572);
and U1202 (N_1202,In_857,In_605);
or U1203 (N_1203,In_67,In_538);
nor U1204 (N_1204,In_211,In_418);
nor U1205 (N_1205,In_902,In_826);
xnor U1206 (N_1206,In_799,In_299);
xor U1207 (N_1207,In_553,In_815);
xor U1208 (N_1208,In_111,In_590);
or U1209 (N_1209,In_362,In_652);
xnor U1210 (N_1210,In_720,In_153);
xor U1211 (N_1211,In_723,In_403);
xor U1212 (N_1212,In_783,In_332);
nor U1213 (N_1213,In_965,In_199);
and U1214 (N_1214,In_743,In_457);
and U1215 (N_1215,In_660,In_523);
nand U1216 (N_1216,In_321,In_662);
or U1217 (N_1217,In_887,In_411);
nand U1218 (N_1218,In_535,In_303);
nand U1219 (N_1219,In_881,In_411);
xor U1220 (N_1220,In_904,In_670);
nand U1221 (N_1221,In_161,In_710);
nand U1222 (N_1222,In_265,In_528);
nor U1223 (N_1223,In_803,In_256);
nor U1224 (N_1224,In_364,In_981);
nor U1225 (N_1225,In_555,In_131);
or U1226 (N_1226,In_781,In_722);
and U1227 (N_1227,In_858,In_14);
nand U1228 (N_1228,In_902,In_312);
or U1229 (N_1229,In_475,In_549);
nor U1230 (N_1230,In_17,In_367);
xor U1231 (N_1231,In_108,In_388);
nand U1232 (N_1232,In_795,In_966);
and U1233 (N_1233,In_87,In_397);
xnor U1234 (N_1234,In_476,In_901);
xor U1235 (N_1235,In_47,In_258);
xor U1236 (N_1236,In_52,In_358);
xnor U1237 (N_1237,In_87,In_50);
nand U1238 (N_1238,In_624,In_330);
nor U1239 (N_1239,In_763,In_283);
xor U1240 (N_1240,In_630,In_977);
and U1241 (N_1241,In_386,In_278);
nand U1242 (N_1242,In_802,In_196);
nor U1243 (N_1243,In_945,In_827);
xor U1244 (N_1244,In_872,In_130);
nand U1245 (N_1245,In_365,In_405);
and U1246 (N_1246,In_560,In_442);
xor U1247 (N_1247,In_477,In_347);
and U1248 (N_1248,In_509,In_680);
nor U1249 (N_1249,In_865,In_3);
nand U1250 (N_1250,In_547,In_938);
or U1251 (N_1251,In_950,In_366);
or U1252 (N_1252,In_804,In_199);
nor U1253 (N_1253,In_710,In_900);
xnor U1254 (N_1254,In_125,In_930);
nor U1255 (N_1255,In_391,In_421);
nor U1256 (N_1256,In_342,In_115);
nor U1257 (N_1257,In_706,In_39);
and U1258 (N_1258,In_602,In_9);
xnor U1259 (N_1259,In_608,In_435);
or U1260 (N_1260,In_403,In_259);
xor U1261 (N_1261,In_465,In_526);
nand U1262 (N_1262,In_958,In_676);
or U1263 (N_1263,In_831,In_71);
nand U1264 (N_1264,In_822,In_55);
xor U1265 (N_1265,In_851,In_936);
and U1266 (N_1266,In_418,In_144);
xnor U1267 (N_1267,In_968,In_542);
nor U1268 (N_1268,In_47,In_428);
xnor U1269 (N_1269,In_173,In_298);
xnor U1270 (N_1270,In_325,In_817);
and U1271 (N_1271,In_552,In_163);
xor U1272 (N_1272,In_209,In_215);
nand U1273 (N_1273,In_255,In_827);
nand U1274 (N_1274,In_330,In_634);
xnor U1275 (N_1275,In_761,In_484);
xor U1276 (N_1276,In_140,In_295);
xor U1277 (N_1277,In_443,In_845);
and U1278 (N_1278,In_568,In_197);
and U1279 (N_1279,In_533,In_507);
nand U1280 (N_1280,In_306,In_33);
or U1281 (N_1281,In_711,In_278);
or U1282 (N_1282,In_490,In_321);
xnor U1283 (N_1283,In_826,In_122);
nor U1284 (N_1284,In_960,In_707);
nor U1285 (N_1285,In_863,In_715);
or U1286 (N_1286,In_896,In_607);
xor U1287 (N_1287,In_121,In_956);
and U1288 (N_1288,In_286,In_540);
or U1289 (N_1289,In_104,In_93);
and U1290 (N_1290,In_761,In_987);
nand U1291 (N_1291,In_352,In_788);
nand U1292 (N_1292,In_298,In_778);
and U1293 (N_1293,In_568,In_264);
nand U1294 (N_1294,In_361,In_549);
xnor U1295 (N_1295,In_859,In_242);
xor U1296 (N_1296,In_895,In_483);
xnor U1297 (N_1297,In_794,In_880);
nor U1298 (N_1298,In_67,In_660);
xnor U1299 (N_1299,In_270,In_766);
or U1300 (N_1300,In_601,In_385);
xnor U1301 (N_1301,In_625,In_148);
nor U1302 (N_1302,In_808,In_637);
nor U1303 (N_1303,In_185,In_476);
xor U1304 (N_1304,In_268,In_345);
nand U1305 (N_1305,In_814,In_118);
or U1306 (N_1306,In_97,In_551);
xor U1307 (N_1307,In_98,In_281);
xnor U1308 (N_1308,In_724,In_326);
nor U1309 (N_1309,In_71,In_81);
and U1310 (N_1310,In_771,In_412);
nor U1311 (N_1311,In_278,In_406);
and U1312 (N_1312,In_33,In_987);
xnor U1313 (N_1313,In_93,In_680);
nand U1314 (N_1314,In_231,In_7);
nor U1315 (N_1315,In_968,In_524);
nand U1316 (N_1316,In_707,In_445);
and U1317 (N_1317,In_395,In_485);
nor U1318 (N_1318,In_242,In_946);
xnor U1319 (N_1319,In_580,In_814);
xnor U1320 (N_1320,In_934,In_531);
nand U1321 (N_1321,In_694,In_497);
and U1322 (N_1322,In_559,In_73);
xor U1323 (N_1323,In_548,In_785);
or U1324 (N_1324,In_949,In_397);
nor U1325 (N_1325,In_328,In_685);
and U1326 (N_1326,In_305,In_367);
nand U1327 (N_1327,In_640,In_455);
or U1328 (N_1328,In_545,In_231);
nor U1329 (N_1329,In_251,In_461);
nand U1330 (N_1330,In_901,In_328);
nand U1331 (N_1331,In_157,In_30);
or U1332 (N_1332,In_137,In_115);
xnor U1333 (N_1333,In_374,In_65);
xnor U1334 (N_1334,In_379,In_981);
and U1335 (N_1335,In_995,In_869);
xnor U1336 (N_1336,In_367,In_479);
and U1337 (N_1337,In_776,In_735);
nor U1338 (N_1338,In_498,In_868);
nand U1339 (N_1339,In_509,In_740);
nor U1340 (N_1340,In_850,In_870);
nand U1341 (N_1341,In_131,In_804);
nand U1342 (N_1342,In_807,In_192);
nand U1343 (N_1343,In_82,In_262);
nand U1344 (N_1344,In_760,In_491);
nor U1345 (N_1345,In_435,In_108);
and U1346 (N_1346,In_106,In_7);
xnor U1347 (N_1347,In_65,In_398);
or U1348 (N_1348,In_124,In_831);
xnor U1349 (N_1349,In_891,In_286);
and U1350 (N_1350,In_622,In_429);
or U1351 (N_1351,In_997,In_60);
and U1352 (N_1352,In_185,In_249);
or U1353 (N_1353,In_163,In_682);
and U1354 (N_1354,In_187,In_747);
or U1355 (N_1355,In_261,In_943);
nand U1356 (N_1356,In_468,In_429);
and U1357 (N_1357,In_293,In_989);
and U1358 (N_1358,In_215,In_658);
xor U1359 (N_1359,In_495,In_394);
and U1360 (N_1360,In_167,In_858);
and U1361 (N_1361,In_702,In_745);
nand U1362 (N_1362,In_571,In_527);
and U1363 (N_1363,In_823,In_874);
nor U1364 (N_1364,In_676,In_731);
nand U1365 (N_1365,In_784,In_253);
or U1366 (N_1366,In_704,In_920);
xnor U1367 (N_1367,In_460,In_366);
xor U1368 (N_1368,In_141,In_134);
and U1369 (N_1369,In_724,In_74);
or U1370 (N_1370,In_300,In_778);
or U1371 (N_1371,In_438,In_949);
or U1372 (N_1372,In_640,In_995);
and U1373 (N_1373,In_718,In_704);
and U1374 (N_1374,In_814,In_109);
or U1375 (N_1375,In_964,In_511);
nand U1376 (N_1376,In_851,In_495);
xor U1377 (N_1377,In_187,In_326);
xnor U1378 (N_1378,In_348,In_585);
nand U1379 (N_1379,In_631,In_732);
or U1380 (N_1380,In_552,In_16);
and U1381 (N_1381,In_452,In_758);
and U1382 (N_1382,In_134,In_871);
or U1383 (N_1383,In_137,In_465);
nor U1384 (N_1384,In_267,In_435);
nand U1385 (N_1385,In_708,In_126);
nand U1386 (N_1386,In_61,In_279);
or U1387 (N_1387,In_32,In_553);
or U1388 (N_1388,In_468,In_547);
and U1389 (N_1389,In_791,In_917);
or U1390 (N_1390,In_953,In_296);
or U1391 (N_1391,In_324,In_828);
or U1392 (N_1392,In_531,In_925);
nand U1393 (N_1393,In_386,In_222);
nand U1394 (N_1394,In_533,In_217);
nand U1395 (N_1395,In_691,In_816);
nor U1396 (N_1396,In_567,In_767);
nor U1397 (N_1397,In_896,In_782);
and U1398 (N_1398,In_517,In_599);
nor U1399 (N_1399,In_892,In_891);
or U1400 (N_1400,In_773,In_51);
nand U1401 (N_1401,In_858,In_430);
or U1402 (N_1402,In_128,In_253);
and U1403 (N_1403,In_993,In_253);
and U1404 (N_1404,In_182,In_251);
xor U1405 (N_1405,In_597,In_765);
nor U1406 (N_1406,In_512,In_490);
xnor U1407 (N_1407,In_772,In_731);
xor U1408 (N_1408,In_426,In_320);
xor U1409 (N_1409,In_691,In_15);
xnor U1410 (N_1410,In_437,In_411);
and U1411 (N_1411,In_965,In_854);
and U1412 (N_1412,In_196,In_233);
and U1413 (N_1413,In_705,In_345);
and U1414 (N_1414,In_440,In_744);
nand U1415 (N_1415,In_973,In_407);
xor U1416 (N_1416,In_503,In_925);
or U1417 (N_1417,In_62,In_137);
xnor U1418 (N_1418,In_344,In_233);
xnor U1419 (N_1419,In_566,In_99);
nand U1420 (N_1420,In_136,In_340);
nand U1421 (N_1421,In_191,In_364);
or U1422 (N_1422,In_429,In_800);
nand U1423 (N_1423,In_830,In_585);
or U1424 (N_1424,In_834,In_324);
xnor U1425 (N_1425,In_7,In_149);
nand U1426 (N_1426,In_313,In_962);
nor U1427 (N_1427,In_127,In_735);
or U1428 (N_1428,In_431,In_416);
and U1429 (N_1429,In_888,In_17);
or U1430 (N_1430,In_175,In_285);
nand U1431 (N_1431,In_901,In_452);
xnor U1432 (N_1432,In_679,In_166);
or U1433 (N_1433,In_251,In_610);
and U1434 (N_1434,In_870,In_344);
and U1435 (N_1435,In_278,In_440);
xor U1436 (N_1436,In_530,In_37);
or U1437 (N_1437,In_992,In_77);
and U1438 (N_1438,In_758,In_442);
xor U1439 (N_1439,In_282,In_691);
nand U1440 (N_1440,In_672,In_676);
nand U1441 (N_1441,In_872,In_567);
xor U1442 (N_1442,In_801,In_872);
nand U1443 (N_1443,In_304,In_433);
nand U1444 (N_1444,In_874,In_918);
or U1445 (N_1445,In_254,In_30);
or U1446 (N_1446,In_354,In_423);
or U1447 (N_1447,In_109,In_427);
nor U1448 (N_1448,In_272,In_795);
or U1449 (N_1449,In_297,In_154);
or U1450 (N_1450,In_853,In_402);
and U1451 (N_1451,In_141,In_146);
or U1452 (N_1452,In_289,In_999);
nor U1453 (N_1453,In_604,In_899);
nor U1454 (N_1454,In_473,In_957);
nand U1455 (N_1455,In_490,In_291);
xor U1456 (N_1456,In_810,In_115);
or U1457 (N_1457,In_370,In_6);
and U1458 (N_1458,In_56,In_742);
nor U1459 (N_1459,In_733,In_102);
nor U1460 (N_1460,In_720,In_575);
xnor U1461 (N_1461,In_492,In_614);
nand U1462 (N_1462,In_340,In_449);
and U1463 (N_1463,In_628,In_188);
or U1464 (N_1464,In_276,In_796);
nor U1465 (N_1465,In_767,In_34);
or U1466 (N_1466,In_751,In_724);
nor U1467 (N_1467,In_211,In_677);
nor U1468 (N_1468,In_542,In_656);
nand U1469 (N_1469,In_489,In_826);
and U1470 (N_1470,In_892,In_960);
nand U1471 (N_1471,In_737,In_914);
xnor U1472 (N_1472,In_457,In_436);
xor U1473 (N_1473,In_130,In_293);
or U1474 (N_1474,In_353,In_593);
and U1475 (N_1475,In_463,In_402);
nand U1476 (N_1476,In_259,In_973);
or U1477 (N_1477,In_73,In_20);
xnor U1478 (N_1478,In_127,In_377);
xnor U1479 (N_1479,In_565,In_324);
and U1480 (N_1480,In_841,In_417);
and U1481 (N_1481,In_296,In_796);
nor U1482 (N_1482,In_88,In_452);
and U1483 (N_1483,In_274,In_200);
and U1484 (N_1484,In_462,In_879);
and U1485 (N_1485,In_514,In_393);
and U1486 (N_1486,In_826,In_979);
nor U1487 (N_1487,In_332,In_349);
or U1488 (N_1488,In_153,In_323);
xor U1489 (N_1489,In_497,In_23);
xor U1490 (N_1490,In_224,In_570);
or U1491 (N_1491,In_465,In_858);
or U1492 (N_1492,In_137,In_574);
or U1493 (N_1493,In_790,In_673);
and U1494 (N_1494,In_719,In_419);
nand U1495 (N_1495,In_396,In_917);
nor U1496 (N_1496,In_798,In_811);
and U1497 (N_1497,In_614,In_838);
xnor U1498 (N_1498,In_257,In_453);
or U1499 (N_1499,In_609,In_676);
and U1500 (N_1500,In_850,In_295);
or U1501 (N_1501,In_127,In_373);
xor U1502 (N_1502,In_733,In_984);
xor U1503 (N_1503,In_531,In_605);
or U1504 (N_1504,In_135,In_391);
xnor U1505 (N_1505,In_335,In_840);
or U1506 (N_1506,In_370,In_154);
or U1507 (N_1507,In_734,In_369);
xor U1508 (N_1508,In_595,In_575);
or U1509 (N_1509,In_204,In_884);
nand U1510 (N_1510,In_68,In_69);
or U1511 (N_1511,In_595,In_828);
or U1512 (N_1512,In_149,In_16);
nand U1513 (N_1513,In_171,In_950);
or U1514 (N_1514,In_162,In_156);
nor U1515 (N_1515,In_837,In_607);
and U1516 (N_1516,In_132,In_231);
xor U1517 (N_1517,In_363,In_514);
nor U1518 (N_1518,In_990,In_197);
xnor U1519 (N_1519,In_28,In_48);
and U1520 (N_1520,In_293,In_182);
nand U1521 (N_1521,In_853,In_125);
nor U1522 (N_1522,In_376,In_900);
nor U1523 (N_1523,In_735,In_405);
nor U1524 (N_1524,In_51,In_722);
and U1525 (N_1525,In_982,In_435);
or U1526 (N_1526,In_994,In_44);
and U1527 (N_1527,In_617,In_135);
nor U1528 (N_1528,In_230,In_254);
or U1529 (N_1529,In_669,In_419);
and U1530 (N_1530,In_750,In_530);
nor U1531 (N_1531,In_729,In_169);
and U1532 (N_1532,In_625,In_895);
and U1533 (N_1533,In_72,In_42);
nand U1534 (N_1534,In_595,In_179);
and U1535 (N_1535,In_722,In_504);
xnor U1536 (N_1536,In_464,In_130);
and U1537 (N_1537,In_830,In_117);
nor U1538 (N_1538,In_67,In_912);
or U1539 (N_1539,In_872,In_959);
nand U1540 (N_1540,In_641,In_541);
nor U1541 (N_1541,In_562,In_878);
nand U1542 (N_1542,In_863,In_619);
and U1543 (N_1543,In_503,In_572);
or U1544 (N_1544,In_173,In_336);
nor U1545 (N_1545,In_658,In_458);
or U1546 (N_1546,In_702,In_436);
or U1547 (N_1547,In_934,In_871);
nand U1548 (N_1548,In_18,In_388);
xnor U1549 (N_1549,In_581,In_796);
xor U1550 (N_1550,In_333,In_353);
or U1551 (N_1551,In_72,In_532);
nand U1552 (N_1552,In_603,In_351);
nand U1553 (N_1553,In_756,In_453);
xor U1554 (N_1554,In_540,In_188);
xor U1555 (N_1555,In_968,In_25);
nor U1556 (N_1556,In_201,In_804);
nor U1557 (N_1557,In_563,In_221);
or U1558 (N_1558,In_57,In_20);
nor U1559 (N_1559,In_505,In_35);
nand U1560 (N_1560,In_790,In_557);
or U1561 (N_1561,In_823,In_44);
nor U1562 (N_1562,In_403,In_366);
and U1563 (N_1563,In_934,In_994);
or U1564 (N_1564,In_907,In_403);
and U1565 (N_1565,In_455,In_562);
nor U1566 (N_1566,In_579,In_365);
and U1567 (N_1567,In_317,In_198);
and U1568 (N_1568,In_201,In_411);
nor U1569 (N_1569,In_62,In_803);
xnor U1570 (N_1570,In_696,In_964);
xor U1571 (N_1571,In_155,In_685);
and U1572 (N_1572,In_642,In_244);
and U1573 (N_1573,In_683,In_899);
or U1574 (N_1574,In_717,In_150);
nand U1575 (N_1575,In_28,In_98);
nor U1576 (N_1576,In_865,In_555);
nor U1577 (N_1577,In_140,In_262);
nand U1578 (N_1578,In_619,In_792);
nor U1579 (N_1579,In_595,In_671);
and U1580 (N_1580,In_936,In_858);
and U1581 (N_1581,In_300,In_355);
nor U1582 (N_1582,In_665,In_739);
xnor U1583 (N_1583,In_583,In_613);
nand U1584 (N_1584,In_689,In_859);
nor U1585 (N_1585,In_123,In_883);
and U1586 (N_1586,In_874,In_771);
xor U1587 (N_1587,In_35,In_118);
and U1588 (N_1588,In_431,In_975);
nor U1589 (N_1589,In_555,In_40);
xor U1590 (N_1590,In_836,In_956);
and U1591 (N_1591,In_775,In_437);
nand U1592 (N_1592,In_218,In_332);
or U1593 (N_1593,In_94,In_726);
nand U1594 (N_1594,In_828,In_49);
nand U1595 (N_1595,In_865,In_450);
nand U1596 (N_1596,In_207,In_664);
xnor U1597 (N_1597,In_779,In_46);
xor U1598 (N_1598,In_370,In_106);
nand U1599 (N_1599,In_93,In_175);
nand U1600 (N_1600,In_887,In_844);
nand U1601 (N_1601,In_222,In_749);
and U1602 (N_1602,In_803,In_788);
or U1603 (N_1603,In_377,In_225);
nand U1604 (N_1604,In_762,In_116);
and U1605 (N_1605,In_275,In_518);
nor U1606 (N_1606,In_832,In_598);
nand U1607 (N_1607,In_614,In_362);
xor U1608 (N_1608,In_80,In_431);
nor U1609 (N_1609,In_798,In_491);
or U1610 (N_1610,In_50,In_618);
and U1611 (N_1611,In_612,In_498);
and U1612 (N_1612,In_49,In_371);
and U1613 (N_1613,In_982,In_690);
and U1614 (N_1614,In_32,In_290);
nand U1615 (N_1615,In_675,In_493);
and U1616 (N_1616,In_645,In_905);
nand U1617 (N_1617,In_855,In_831);
nand U1618 (N_1618,In_609,In_619);
nand U1619 (N_1619,In_198,In_24);
or U1620 (N_1620,In_307,In_676);
nor U1621 (N_1621,In_311,In_551);
nor U1622 (N_1622,In_207,In_331);
or U1623 (N_1623,In_864,In_37);
nor U1624 (N_1624,In_411,In_855);
xor U1625 (N_1625,In_735,In_328);
nand U1626 (N_1626,In_245,In_910);
or U1627 (N_1627,In_393,In_25);
or U1628 (N_1628,In_629,In_360);
nor U1629 (N_1629,In_471,In_505);
nor U1630 (N_1630,In_828,In_4);
nand U1631 (N_1631,In_330,In_257);
and U1632 (N_1632,In_820,In_242);
nor U1633 (N_1633,In_908,In_13);
and U1634 (N_1634,In_705,In_274);
and U1635 (N_1635,In_56,In_261);
nor U1636 (N_1636,In_976,In_313);
nand U1637 (N_1637,In_938,In_630);
xor U1638 (N_1638,In_885,In_210);
and U1639 (N_1639,In_195,In_21);
or U1640 (N_1640,In_206,In_376);
or U1641 (N_1641,In_793,In_155);
xor U1642 (N_1642,In_662,In_644);
or U1643 (N_1643,In_537,In_441);
or U1644 (N_1644,In_429,In_271);
xnor U1645 (N_1645,In_882,In_53);
nand U1646 (N_1646,In_269,In_814);
nor U1647 (N_1647,In_61,In_177);
xnor U1648 (N_1648,In_22,In_833);
nand U1649 (N_1649,In_707,In_743);
and U1650 (N_1650,In_837,In_86);
and U1651 (N_1651,In_425,In_393);
nand U1652 (N_1652,In_924,In_637);
nor U1653 (N_1653,In_347,In_211);
nand U1654 (N_1654,In_679,In_656);
or U1655 (N_1655,In_570,In_247);
nor U1656 (N_1656,In_468,In_22);
and U1657 (N_1657,In_578,In_849);
or U1658 (N_1658,In_545,In_557);
xnor U1659 (N_1659,In_202,In_190);
nor U1660 (N_1660,In_12,In_265);
or U1661 (N_1661,In_578,In_54);
or U1662 (N_1662,In_25,In_45);
nor U1663 (N_1663,In_102,In_593);
xnor U1664 (N_1664,In_177,In_133);
nor U1665 (N_1665,In_977,In_233);
and U1666 (N_1666,In_345,In_826);
nand U1667 (N_1667,In_144,In_615);
xor U1668 (N_1668,In_222,In_971);
and U1669 (N_1669,In_167,In_461);
and U1670 (N_1670,In_283,In_738);
nor U1671 (N_1671,In_907,In_542);
nand U1672 (N_1672,In_113,In_961);
xor U1673 (N_1673,In_598,In_758);
nand U1674 (N_1674,In_192,In_99);
nand U1675 (N_1675,In_788,In_314);
nor U1676 (N_1676,In_702,In_763);
and U1677 (N_1677,In_338,In_582);
nor U1678 (N_1678,In_387,In_105);
nor U1679 (N_1679,In_289,In_843);
nand U1680 (N_1680,In_405,In_66);
and U1681 (N_1681,In_531,In_12);
nand U1682 (N_1682,In_827,In_603);
nand U1683 (N_1683,In_142,In_433);
nor U1684 (N_1684,In_251,In_732);
nor U1685 (N_1685,In_23,In_193);
or U1686 (N_1686,In_606,In_6);
nor U1687 (N_1687,In_213,In_459);
or U1688 (N_1688,In_786,In_110);
or U1689 (N_1689,In_386,In_195);
or U1690 (N_1690,In_883,In_523);
xor U1691 (N_1691,In_157,In_251);
nor U1692 (N_1692,In_563,In_960);
or U1693 (N_1693,In_458,In_860);
nor U1694 (N_1694,In_463,In_585);
nand U1695 (N_1695,In_733,In_146);
xor U1696 (N_1696,In_813,In_710);
nand U1697 (N_1697,In_722,In_68);
nor U1698 (N_1698,In_490,In_45);
nand U1699 (N_1699,In_355,In_662);
xnor U1700 (N_1700,In_908,In_478);
or U1701 (N_1701,In_640,In_535);
nor U1702 (N_1702,In_161,In_946);
and U1703 (N_1703,In_41,In_922);
xor U1704 (N_1704,In_322,In_654);
nand U1705 (N_1705,In_480,In_169);
and U1706 (N_1706,In_650,In_752);
nor U1707 (N_1707,In_650,In_696);
and U1708 (N_1708,In_44,In_867);
or U1709 (N_1709,In_743,In_226);
xor U1710 (N_1710,In_862,In_923);
nand U1711 (N_1711,In_890,In_101);
xnor U1712 (N_1712,In_824,In_121);
and U1713 (N_1713,In_601,In_363);
and U1714 (N_1714,In_448,In_198);
and U1715 (N_1715,In_741,In_617);
and U1716 (N_1716,In_204,In_624);
nand U1717 (N_1717,In_915,In_849);
nor U1718 (N_1718,In_384,In_917);
nand U1719 (N_1719,In_439,In_6);
nand U1720 (N_1720,In_518,In_895);
and U1721 (N_1721,In_12,In_948);
xor U1722 (N_1722,In_651,In_718);
or U1723 (N_1723,In_4,In_52);
or U1724 (N_1724,In_367,In_268);
nand U1725 (N_1725,In_759,In_214);
xnor U1726 (N_1726,In_428,In_170);
nand U1727 (N_1727,In_213,In_970);
nand U1728 (N_1728,In_370,In_710);
nand U1729 (N_1729,In_690,In_355);
nor U1730 (N_1730,In_614,In_354);
and U1731 (N_1731,In_213,In_245);
xor U1732 (N_1732,In_184,In_744);
nand U1733 (N_1733,In_575,In_876);
or U1734 (N_1734,In_119,In_353);
and U1735 (N_1735,In_249,In_308);
xnor U1736 (N_1736,In_900,In_323);
xor U1737 (N_1737,In_563,In_520);
and U1738 (N_1738,In_89,In_482);
and U1739 (N_1739,In_68,In_688);
or U1740 (N_1740,In_444,In_372);
or U1741 (N_1741,In_532,In_167);
nor U1742 (N_1742,In_194,In_797);
or U1743 (N_1743,In_360,In_775);
xor U1744 (N_1744,In_382,In_285);
nand U1745 (N_1745,In_185,In_281);
nor U1746 (N_1746,In_222,In_459);
or U1747 (N_1747,In_68,In_554);
nor U1748 (N_1748,In_905,In_302);
nand U1749 (N_1749,In_384,In_130);
and U1750 (N_1750,In_666,In_843);
xnor U1751 (N_1751,In_288,In_902);
and U1752 (N_1752,In_225,In_261);
nor U1753 (N_1753,In_497,In_328);
xor U1754 (N_1754,In_477,In_413);
and U1755 (N_1755,In_998,In_374);
nor U1756 (N_1756,In_321,In_93);
nor U1757 (N_1757,In_885,In_96);
or U1758 (N_1758,In_88,In_185);
nor U1759 (N_1759,In_74,In_149);
nand U1760 (N_1760,In_649,In_27);
nor U1761 (N_1761,In_306,In_90);
nand U1762 (N_1762,In_865,In_561);
nor U1763 (N_1763,In_845,In_442);
nor U1764 (N_1764,In_714,In_827);
nor U1765 (N_1765,In_577,In_784);
nand U1766 (N_1766,In_492,In_407);
nand U1767 (N_1767,In_187,In_208);
or U1768 (N_1768,In_136,In_823);
nand U1769 (N_1769,In_124,In_86);
nor U1770 (N_1770,In_629,In_342);
nor U1771 (N_1771,In_380,In_365);
nor U1772 (N_1772,In_530,In_275);
nand U1773 (N_1773,In_569,In_889);
nor U1774 (N_1774,In_506,In_110);
nor U1775 (N_1775,In_85,In_271);
nand U1776 (N_1776,In_4,In_26);
nor U1777 (N_1777,In_625,In_76);
xnor U1778 (N_1778,In_728,In_436);
nor U1779 (N_1779,In_387,In_155);
or U1780 (N_1780,In_455,In_479);
and U1781 (N_1781,In_848,In_363);
and U1782 (N_1782,In_338,In_469);
or U1783 (N_1783,In_516,In_105);
xnor U1784 (N_1784,In_949,In_910);
or U1785 (N_1785,In_238,In_332);
and U1786 (N_1786,In_420,In_658);
nor U1787 (N_1787,In_869,In_74);
xnor U1788 (N_1788,In_967,In_577);
and U1789 (N_1789,In_376,In_74);
nor U1790 (N_1790,In_739,In_584);
or U1791 (N_1791,In_192,In_548);
and U1792 (N_1792,In_484,In_631);
and U1793 (N_1793,In_493,In_317);
xnor U1794 (N_1794,In_152,In_545);
xor U1795 (N_1795,In_429,In_247);
nand U1796 (N_1796,In_550,In_937);
and U1797 (N_1797,In_313,In_891);
nor U1798 (N_1798,In_996,In_871);
nand U1799 (N_1799,In_154,In_851);
or U1800 (N_1800,In_688,In_146);
nand U1801 (N_1801,In_138,In_702);
xnor U1802 (N_1802,In_992,In_556);
or U1803 (N_1803,In_898,In_132);
nor U1804 (N_1804,In_915,In_747);
nand U1805 (N_1805,In_726,In_785);
or U1806 (N_1806,In_304,In_379);
and U1807 (N_1807,In_255,In_570);
or U1808 (N_1808,In_871,In_318);
nand U1809 (N_1809,In_115,In_559);
nand U1810 (N_1810,In_586,In_627);
and U1811 (N_1811,In_126,In_523);
xnor U1812 (N_1812,In_128,In_552);
and U1813 (N_1813,In_361,In_81);
nor U1814 (N_1814,In_57,In_79);
nor U1815 (N_1815,In_379,In_201);
or U1816 (N_1816,In_498,In_142);
nand U1817 (N_1817,In_935,In_45);
or U1818 (N_1818,In_754,In_258);
nor U1819 (N_1819,In_124,In_981);
nand U1820 (N_1820,In_310,In_73);
nor U1821 (N_1821,In_615,In_542);
and U1822 (N_1822,In_222,In_25);
nand U1823 (N_1823,In_642,In_128);
and U1824 (N_1824,In_764,In_225);
nand U1825 (N_1825,In_804,In_279);
or U1826 (N_1826,In_941,In_987);
nand U1827 (N_1827,In_676,In_9);
xnor U1828 (N_1828,In_51,In_543);
nand U1829 (N_1829,In_978,In_585);
xnor U1830 (N_1830,In_778,In_952);
and U1831 (N_1831,In_140,In_267);
nand U1832 (N_1832,In_242,In_32);
nand U1833 (N_1833,In_239,In_493);
and U1834 (N_1834,In_555,In_239);
or U1835 (N_1835,In_885,In_91);
and U1836 (N_1836,In_837,In_409);
xor U1837 (N_1837,In_745,In_127);
nor U1838 (N_1838,In_381,In_49);
and U1839 (N_1839,In_790,In_133);
nand U1840 (N_1840,In_299,In_687);
xor U1841 (N_1841,In_193,In_298);
nor U1842 (N_1842,In_875,In_266);
xnor U1843 (N_1843,In_701,In_635);
and U1844 (N_1844,In_662,In_590);
and U1845 (N_1845,In_398,In_228);
or U1846 (N_1846,In_454,In_268);
xnor U1847 (N_1847,In_559,In_859);
xnor U1848 (N_1848,In_895,In_470);
and U1849 (N_1849,In_869,In_970);
nor U1850 (N_1850,In_252,In_405);
or U1851 (N_1851,In_463,In_454);
and U1852 (N_1852,In_128,In_25);
or U1853 (N_1853,In_201,In_673);
and U1854 (N_1854,In_52,In_490);
nand U1855 (N_1855,In_169,In_687);
xor U1856 (N_1856,In_413,In_0);
nand U1857 (N_1857,In_918,In_117);
xor U1858 (N_1858,In_162,In_147);
or U1859 (N_1859,In_780,In_248);
and U1860 (N_1860,In_461,In_872);
nor U1861 (N_1861,In_45,In_696);
nor U1862 (N_1862,In_150,In_604);
nand U1863 (N_1863,In_296,In_118);
or U1864 (N_1864,In_959,In_327);
xnor U1865 (N_1865,In_649,In_998);
nand U1866 (N_1866,In_591,In_611);
nand U1867 (N_1867,In_565,In_310);
xnor U1868 (N_1868,In_768,In_537);
nor U1869 (N_1869,In_28,In_989);
nor U1870 (N_1870,In_419,In_704);
xnor U1871 (N_1871,In_960,In_995);
and U1872 (N_1872,In_371,In_292);
nor U1873 (N_1873,In_721,In_377);
or U1874 (N_1874,In_662,In_383);
nand U1875 (N_1875,In_538,In_271);
or U1876 (N_1876,In_805,In_734);
or U1877 (N_1877,In_365,In_876);
or U1878 (N_1878,In_509,In_38);
nor U1879 (N_1879,In_704,In_324);
nand U1880 (N_1880,In_563,In_142);
and U1881 (N_1881,In_445,In_120);
nand U1882 (N_1882,In_862,In_284);
nor U1883 (N_1883,In_244,In_89);
nand U1884 (N_1884,In_599,In_486);
or U1885 (N_1885,In_325,In_620);
or U1886 (N_1886,In_289,In_589);
or U1887 (N_1887,In_189,In_590);
nor U1888 (N_1888,In_591,In_248);
nand U1889 (N_1889,In_467,In_334);
xor U1890 (N_1890,In_706,In_717);
nor U1891 (N_1891,In_112,In_874);
or U1892 (N_1892,In_127,In_136);
nor U1893 (N_1893,In_692,In_929);
or U1894 (N_1894,In_472,In_383);
nand U1895 (N_1895,In_517,In_958);
nor U1896 (N_1896,In_685,In_779);
nor U1897 (N_1897,In_515,In_898);
nand U1898 (N_1898,In_93,In_727);
and U1899 (N_1899,In_36,In_4);
or U1900 (N_1900,In_36,In_864);
xnor U1901 (N_1901,In_224,In_734);
xnor U1902 (N_1902,In_912,In_60);
nand U1903 (N_1903,In_403,In_606);
and U1904 (N_1904,In_997,In_843);
and U1905 (N_1905,In_58,In_940);
and U1906 (N_1906,In_179,In_215);
nand U1907 (N_1907,In_69,In_76);
nor U1908 (N_1908,In_880,In_25);
xor U1909 (N_1909,In_427,In_241);
nand U1910 (N_1910,In_803,In_0);
and U1911 (N_1911,In_480,In_919);
and U1912 (N_1912,In_20,In_499);
and U1913 (N_1913,In_141,In_142);
nand U1914 (N_1914,In_951,In_132);
nand U1915 (N_1915,In_25,In_142);
nor U1916 (N_1916,In_625,In_130);
xor U1917 (N_1917,In_218,In_945);
and U1918 (N_1918,In_71,In_176);
or U1919 (N_1919,In_356,In_189);
xor U1920 (N_1920,In_856,In_77);
and U1921 (N_1921,In_940,In_18);
xnor U1922 (N_1922,In_312,In_108);
or U1923 (N_1923,In_411,In_85);
xnor U1924 (N_1924,In_998,In_946);
and U1925 (N_1925,In_284,In_713);
or U1926 (N_1926,In_255,In_675);
or U1927 (N_1927,In_994,In_616);
nor U1928 (N_1928,In_564,In_86);
or U1929 (N_1929,In_742,In_383);
or U1930 (N_1930,In_106,In_368);
nor U1931 (N_1931,In_303,In_547);
xor U1932 (N_1932,In_160,In_863);
or U1933 (N_1933,In_680,In_960);
and U1934 (N_1934,In_325,In_692);
or U1935 (N_1935,In_258,In_287);
xor U1936 (N_1936,In_991,In_160);
or U1937 (N_1937,In_432,In_450);
and U1938 (N_1938,In_58,In_887);
and U1939 (N_1939,In_914,In_19);
and U1940 (N_1940,In_922,In_177);
nor U1941 (N_1941,In_233,In_778);
and U1942 (N_1942,In_365,In_799);
nor U1943 (N_1943,In_526,In_36);
or U1944 (N_1944,In_169,In_651);
or U1945 (N_1945,In_301,In_128);
nor U1946 (N_1946,In_64,In_19);
nand U1947 (N_1947,In_130,In_913);
nor U1948 (N_1948,In_563,In_350);
nor U1949 (N_1949,In_532,In_646);
xnor U1950 (N_1950,In_2,In_248);
xnor U1951 (N_1951,In_169,In_455);
nor U1952 (N_1952,In_95,In_765);
nor U1953 (N_1953,In_450,In_414);
xor U1954 (N_1954,In_929,In_157);
nand U1955 (N_1955,In_399,In_869);
nand U1956 (N_1956,In_433,In_819);
and U1957 (N_1957,In_572,In_741);
and U1958 (N_1958,In_333,In_285);
nand U1959 (N_1959,In_752,In_300);
nor U1960 (N_1960,In_268,In_628);
nor U1961 (N_1961,In_8,In_373);
nor U1962 (N_1962,In_631,In_896);
or U1963 (N_1963,In_861,In_241);
xor U1964 (N_1964,In_176,In_584);
or U1965 (N_1965,In_548,In_675);
or U1966 (N_1966,In_739,In_641);
nor U1967 (N_1967,In_6,In_652);
xor U1968 (N_1968,In_89,In_895);
xor U1969 (N_1969,In_462,In_456);
nand U1970 (N_1970,In_406,In_185);
nor U1971 (N_1971,In_197,In_457);
and U1972 (N_1972,In_652,In_864);
xnor U1973 (N_1973,In_20,In_646);
nand U1974 (N_1974,In_485,In_768);
and U1975 (N_1975,In_556,In_729);
or U1976 (N_1976,In_400,In_691);
nor U1977 (N_1977,In_930,In_908);
xor U1978 (N_1978,In_757,In_863);
nand U1979 (N_1979,In_342,In_281);
nand U1980 (N_1980,In_356,In_157);
or U1981 (N_1981,In_960,In_709);
or U1982 (N_1982,In_734,In_798);
xor U1983 (N_1983,In_677,In_391);
xnor U1984 (N_1984,In_309,In_821);
xnor U1985 (N_1985,In_909,In_633);
or U1986 (N_1986,In_226,In_153);
nand U1987 (N_1987,In_223,In_281);
xnor U1988 (N_1988,In_601,In_490);
and U1989 (N_1989,In_10,In_658);
xor U1990 (N_1990,In_838,In_247);
or U1991 (N_1991,In_111,In_639);
xnor U1992 (N_1992,In_978,In_194);
or U1993 (N_1993,In_159,In_820);
or U1994 (N_1994,In_635,In_558);
nor U1995 (N_1995,In_556,In_424);
or U1996 (N_1996,In_87,In_139);
nor U1997 (N_1997,In_858,In_87);
xor U1998 (N_1998,In_624,In_773);
xnor U1999 (N_1999,In_385,In_873);
nor U2000 (N_2000,In_443,In_232);
nor U2001 (N_2001,In_479,In_175);
nand U2002 (N_2002,In_220,In_689);
nand U2003 (N_2003,In_748,In_381);
nor U2004 (N_2004,In_174,In_609);
nor U2005 (N_2005,In_907,In_253);
nor U2006 (N_2006,In_536,In_538);
nand U2007 (N_2007,In_823,In_779);
nand U2008 (N_2008,In_388,In_977);
or U2009 (N_2009,In_810,In_511);
nand U2010 (N_2010,In_495,In_981);
and U2011 (N_2011,In_785,In_440);
or U2012 (N_2012,In_482,In_864);
xor U2013 (N_2013,In_286,In_34);
nor U2014 (N_2014,In_74,In_287);
or U2015 (N_2015,In_325,In_163);
and U2016 (N_2016,In_269,In_345);
nor U2017 (N_2017,In_955,In_445);
or U2018 (N_2018,In_596,In_582);
nor U2019 (N_2019,In_971,In_985);
or U2020 (N_2020,In_956,In_168);
and U2021 (N_2021,In_475,In_538);
and U2022 (N_2022,In_943,In_458);
or U2023 (N_2023,In_286,In_962);
nand U2024 (N_2024,In_487,In_465);
nand U2025 (N_2025,In_781,In_590);
xor U2026 (N_2026,In_867,In_870);
nor U2027 (N_2027,In_741,In_180);
or U2028 (N_2028,In_447,In_778);
xnor U2029 (N_2029,In_135,In_867);
and U2030 (N_2030,In_823,In_746);
xor U2031 (N_2031,In_333,In_247);
nor U2032 (N_2032,In_911,In_852);
nor U2033 (N_2033,In_799,In_150);
xnor U2034 (N_2034,In_928,In_84);
or U2035 (N_2035,In_187,In_454);
and U2036 (N_2036,In_208,In_352);
and U2037 (N_2037,In_974,In_711);
and U2038 (N_2038,In_19,In_47);
xor U2039 (N_2039,In_998,In_550);
or U2040 (N_2040,In_888,In_304);
and U2041 (N_2041,In_175,In_497);
nor U2042 (N_2042,In_981,In_469);
or U2043 (N_2043,In_547,In_721);
xnor U2044 (N_2044,In_133,In_808);
or U2045 (N_2045,In_821,In_643);
nor U2046 (N_2046,In_906,In_814);
nand U2047 (N_2047,In_952,In_424);
xnor U2048 (N_2048,In_182,In_781);
xnor U2049 (N_2049,In_964,In_557);
or U2050 (N_2050,In_328,In_637);
xor U2051 (N_2051,In_68,In_868);
xor U2052 (N_2052,In_58,In_116);
or U2053 (N_2053,In_512,In_747);
nor U2054 (N_2054,In_20,In_476);
or U2055 (N_2055,In_11,In_887);
nand U2056 (N_2056,In_558,In_125);
and U2057 (N_2057,In_496,In_806);
and U2058 (N_2058,In_287,In_474);
and U2059 (N_2059,In_104,In_155);
nand U2060 (N_2060,In_234,In_620);
xnor U2061 (N_2061,In_876,In_113);
nor U2062 (N_2062,In_15,In_614);
or U2063 (N_2063,In_143,In_911);
xnor U2064 (N_2064,In_287,In_742);
nor U2065 (N_2065,In_500,In_926);
or U2066 (N_2066,In_387,In_119);
or U2067 (N_2067,In_88,In_160);
xor U2068 (N_2068,In_228,In_913);
and U2069 (N_2069,In_84,In_754);
nor U2070 (N_2070,In_835,In_72);
and U2071 (N_2071,In_704,In_481);
xor U2072 (N_2072,In_742,In_706);
xor U2073 (N_2073,In_55,In_850);
nand U2074 (N_2074,In_916,In_823);
nor U2075 (N_2075,In_866,In_359);
or U2076 (N_2076,In_835,In_421);
and U2077 (N_2077,In_861,In_309);
or U2078 (N_2078,In_33,In_62);
or U2079 (N_2079,In_458,In_276);
xor U2080 (N_2080,In_352,In_36);
nor U2081 (N_2081,In_822,In_682);
nor U2082 (N_2082,In_460,In_186);
nand U2083 (N_2083,In_636,In_608);
and U2084 (N_2084,In_446,In_101);
nor U2085 (N_2085,In_312,In_676);
nor U2086 (N_2086,In_227,In_873);
and U2087 (N_2087,In_504,In_275);
xor U2088 (N_2088,In_868,In_599);
nand U2089 (N_2089,In_290,In_877);
or U2090 (N_2090,In_215,In_134);
xnor U2091 (N_2091,In_465,In_590);
nand U2092 (N_2092,In_548,In_839);
or U2093 (N_2093,In_550,In_391);
or U2094 (N_2094,In_456,In_111);
or U2095 (N_2095,In_329,In_651);
or U2096 (N_2096,In_829,In_760);
or U2097 (N_2097,In_172,In_629);
nor U2098 (N_2098,In_635,In_493);
or U2099 (N_2099,In_541,In_786);
nor U2100 (N_2100,In_89,In_658);
xor U2101 (N_2101,In_727,In_971);
xnor U2102 (N_2102,In_686,In_955);
nor U2103 (N_2103,In_658,In_91);
nand U2104 (N_2104,In_31,In_647);
or U2105 (N_2105,In_422,In_691);
nor U2106 (N_2106,In_394,In_425);
or U2107 (N_2107,In_997,In_529);
nor U2108 (N_2108,In_125,In_134);
or U2109 (N_2109,In_731,In_656);
nor U2110 (N_2110,In_688,In_248);
nand U2111 (N_2111,In_52,In_728);
and U2112 (N_2112,In_877,In_830);
nand U2113 (N_2113,In_807,In_889);
and U2114 (N_2114,In_614,In_539);
or U2115 (N_2115,In_268,In_673);
xor U2116 (N_2116,In_390,In_965);
or U2117 (N_2117,In_412,In_591);
or U2118 (N_2118,In_294,In_819);
and U2119 (N_2119,In_692,In_95);
nor U2120 (N_2120,In_897,In_972);
nor U2121 (N_2121,In_914,In_754);
xnor U2122 (N_2122,In_891,In_861);
nor U2123 (N_2123,In_285,In_773);
or U2124 (N_2124,In_348,In_833);
nor U2125 (N_2125,In_551,In_186);
nand U2126 (N_2126,In_561,In_678);
nand U2127 (N_2127,In_551,In_119);
nand U2128 (N_2128,In_814,In_904);
xor U2129 (N_2129,In_687,In_440);
and U2130 (N_2130,In_449,In_824);
or U2131 (N_2131,In_763,In_473);
nand U2132 (N_2132,In_738,In_97);
xnor U2133 (N_2133,In_335,In_718);
or U2134 (N_2134,In_723,In_862);
or U2135 (N_2135,In_880,In_926);
or U2136 (N_2136,In_763,In_699);
or U2137 (N_2137,In_777,In_835);
xor U2138 (N_2138,In_771,In_890);
and U2139 (N_2139,In_624,In_573);
nand U2140 (N_2140,In_780,In_334);
nor U2141 (N_2141,In_936,In_179);
or U2142 (N_2142,In_173,In_530);
xnor U2143 (N_2143,In_876,In_263);
nor U2144 (N_2144,In_936,In_984);
xor U2145 (N_2145,In_762,In_850);
and U2146 (N_2146,In_320,In_867);
nor U2147 (N_2147,In_104,In_936);
xor U2148 (N_2148,In_344,In_413);
and U2149 (N_2149,In_937,In_387);
nor U2150 (N_2150,In_274,In_795);
and U2151 (N_2151,In_422,In_785);
or U2152 (N_2152,In_7,In_996);
or U2153 (N_2153,In_713,In_275);
xor U2154 (N_2154,In_430,In_241);
nor U2155 (N_2155,In_50,In_261);
or U2156 (N_2156,In_84,In_354);
nand U2157 (N_2157,In_784,In_769);
nor U2158 (N_2158,In_916,In_795);
or U2159 (N_2159,In_970,In_463);
or U2160 (N_2160,In_7,In_127);
nand U2161 (N_2161,In_725,In_588);
and U2162 (N_2162,In_641,In_217);
and U2163 (N_2163,In_321,In_911);
or U2164 (N_2164,In_160,In_467);
nand U2165 (N_2165,In_496,In_62);
or U2166 (N_2166,In_696,In_954);
xnor U2167 (N_2167,In_326,In_905);
nor U2168 (N_2168,In_146,In_456);
or U2169 (N_2169,In_876,In_456);
and U2170 (N_2170,In_307,In_540);
and U2171 (N_2171,In_552,In_494);
nand U2172 (N_2172,In_460,In_882);
nand U2173 (N_2173,In_35,In_554);
or U2174 (N_2174,In_224,In_291);
and U2175 (N_2175,In_704,In_790);
nand U2176 (N_2176,In_366,In_537);
nor U2177 (N_2177,In_200,In_638);
nor U2178 (N_2178,In_438,In_564);
and U2179 (N_2179,In_581,In_68);
nor U2180 (N_2180,In_891,In_636);
xor U2181 (N_2181,In_497,In_49);
and U2182 (N_2182,In_746,In_642);
or U2183 (N_2183,In_645,In_950);
xor U2184 (N_2184,In_990,In_108);
xnor U2185 (N_2185,In_307,In_998);
and U2186 (N_2186,In_705,In_715);
nor U2187 (N_2187,In_719,In_199);
and U2188 (N_2188,In_247,In_686);
or U2189 (N_2189,In_504,In_478);
nor U2190 (N_2190,In_744,In_606);
nand U2191 (N_2191,In_506,In_715);
nor U2192 (N_2192,In_886,In_541);
xnor U2193 (N_2193,In_860,In_41);
nand U2194 (N_2194,In_725,In_581);
or U2195 (N_2195,In_421,In_654);
nand U2196 (N_2196,In_86,In_413);
xnor U2197 (N_2197,In_238,In_386);
xor U2198 (N_2198,In_536,In_657);
nand U2199 (N_2199,In_21,In_750);
nand U2200 (N_2200,In_492,In_25);
or U2201 (N_2201,In_6,In_504);
and U2202 (N_2202,In_313,In_101);
xnor U2203 (N_2203,In_915,In_174);
xnor U2204 (N_2204,In_763,In_777);
and U2205 (N_2205,In_1,In_490);
nand U2206 (N_2206,In_458,In_375);
xor U2207 (N_2207,In_0,In_819);
and U2208 (N_2208,In_873,In_101);
and U2209 (N_2209,In_491,In_977);
or U2210 (N_2210,In_150,In_870);
or U2211 (N_2211,In_379,In_535);
xor U2212 (N_2212,In_680,In_916);
nor U2213 (N_2213,In_957,In_310);
or U2214 (N_2214,In_338,In_834);
and U2215 (N_2215,In_668,In_110);
xor U2216 (N_2216,In_919,In_567);
nand U2217 (N_2217,In_867,In_883);
nand U2218 (N_2218,In_81,In_553);
and U2219 (N_2219,In_123,In_750);
nor U2220 (N_2220,In_963,In_488);
and U2221 (N_2221,In_2,In_552);
and U2222 (N_2222,In_41,In_326);
nor U2223 (N_2223,In_435,In_677);
nand U2224 (N_2224,In_809,In_262);
nor U2225 (N_2225,In_940,In_442);
nand U2226 (N_2226,In_569,In_927);
xor U2227 (N_2227,In_821,In_926);
and U2228 (N_2228,In_224,In_965);
nor U2229 (N_2229,In_889,In_776);
nor U2230 (N_2230,In_267,In_170);
and U2231 (N_2231,In_246,In_137);
or U2232 (N_2232,In_390,In_680);
or U2233 (N_2233,In_78,In_421);
nand U2234 (N_2234,In_688,In_310);
nand U2235 (N_2235,In_888,In_810);
and U2236 (N_2236,In_280,In_419);
nand U2237 (N_2237,In_737,In_107);
nor U2238 (N_2238,In_272,In_649);
or U2239 (N_2239,In_368,In_273);
nor U2240 (N_2240,In_453,In_28);
xor U2241 (N_2241,In_673,In_464);
or U2242 (N_2242,In_995,In_889);
xnor U2243 (N_2243,In_923,In_860);
nor U2244 (N_2244,In_261,In_549);
xnor U2245 (N_2245,In_891,In_622);
xnor U2246 (N_2246,In_726,In_277);
nor U2247 (N_2247,In_635,In_518);
xor U2248 (N_2248,In_394,In_256);
nand U2249 (N_2249,In_990,In_666);
and U2250 (N_2250,In_184,In_25);
nand U2251 (N_2251,In_573,In_217);
xnor U2252 (N_2252,In_14,In_44);
xnor U2253 (N_2253,In_117,In_869);
nor U2254 (N_2254,In_982,In_232);
and U2255 (N_2255,In_627,In_221);
nand U2256 (N_2256,In_284,In_36);
xor U2257 (N_2257,In_329,In_555);
xnor U2258 (N_2258,In_703,In_518);
nor U2259 (N_2259,In_864,In_696);
nor U2260 (N_2260,In_959,In_209);
nor U2261 (N_2261,In_440,In_8);
and U2262 (N_2262,In_448,In_517);
or U2263 (N_2263,In_818,In_105);
nor U2264 (N_2264,In_852,In_767);
xnor U2265 (N_2265,In_18,In_60);
nand U2266 (N_2266,In_646,In_809);
nor U2267 (N_2267,In_569,In_30);
and U2268 (N_2268,In_203,In_258);
or U2269 (N_2269,In_371,In_714);
or U2270 (N_2270,In_798,In_743);
nand U2271 (N_2271,In_482,In_298);
nand U2272 (N_2272,In_677,In_156);
and U2273 (N_2273,In_906,In_237);
nand U2274 (N_2274,In_39,In_947);
and U2275 (N_2275,In_420,In_68);
and U2276 (N_2276,In_762,In_922);
nor U2277 (N_2277,In_575,In_263);
nor U2278 (N_2278,In_257,In_46);
nand U2279 (N_2279,In_313,In_73);
and U2280 (N_2280,In_36,In_261);
nand U2281 (N_2281,In_57,In_150);
or U2282 (N_2282,In_301,In_96);
and U2283 (N_2283,In_336,In_199);
nand U2284 (N_2284,In_723,In_853);
or U2285 (N_2285,In_655,In_436);
nor U2286 (N_2286,In_926,In_679);
nand U2287 (N_2287,In_851,In_865);
and U2288 (N_2288,In_987,In_803);
or U2289 (N_2289,In_581,In_180);
nor U2290 (N_2290,In_670,In_749);
or U2291 (N_2291,In_598,In_421);
nand U2292 (N_2292,In_369,In_994);
xnor U2293 (N_2293,In_677,In_64);
xor U2294 (N_2294,In_285,In_311);
nand U2295 (N_2295,In_471,In_272);
nor U2296 (N_2296,In_681,In_539);
nand U2297 (N_2297,In_601,In_367);
nand U2298 (N_2298,In_529,In_581);
nor U2299 (N_2299,In_7,In_519);
nand U2300 (N_2300,In_754,In_854);
xor U2301 (N_2301,In_552,In_313);
xor U2302 (N_2302,In_677,In_796);
nand U2303 (N_2303,In_718,In_460);
xnor U2304 (N_2304,In_798,In_113);
or U2305 (N_2305,In_299,In_327);
nand U2306 (N_2306,In_207,In_831);
nor U2307 (N_2307,In_522,In_907);
or U2308 (N_2308,In_556,In_273);
nand U2309 (N_2309,In_736,In_452);
nor U2310 (N_2310,In_981,In_751);
or U2311 (N_2311,In_611,In_659);
nand U2312 (N_2312,In_410,In_618);
xnor U2313 (N_2313,In_786,In_611);
xnor U2314 (N_2314,In_469,In_252);
or U2315 (N_2315,In_736,In_517);
xor U2316 (N_2316,In_877,In_790);
nor U2317 (N_2317,In_305,In_629);
and U2318 (N_2318,In_666,In_752);
or U2319 (N_2319,In_142,In_961);
or U2320 (N_2320,In_798,In_14);
or U2321 (N_2321,In_950,In_820);
xor U2322 (N_2322,In_924,In_884);
xor U2323 (N_2323,In_160,In_171);
xnor U2324 (N_2324,In_7,In_38);
nand U2325 (N_2325,In_32,In_943);
or U2326 (N_2326,In_36,In_701);
xor U2327 (N_2327,In_520,In_950);
nor U2328 (N_2328,In_409,In_344);
or U2329 (N_2329,In_925,In_77);
nor U2330 (N_2330,In_455,In_240);
and U2331 (N_2331,In_108,In_597);
and U2332 (N_2332,In_134,In_175);
nor U2333 (N_2333,In_580,In_287);
nor U2334 (N_2334,In_268,In_176);
nor U2335 (N_2335,In_328,In_694);
xor U2336 (N_2336,In_469,In_467);
nand U2337 (N_2337,In_986,In_868);
or U2338 (N_2338,In_446,In_625);
nor U2339 (N_2339,In_748,In_51);
nand U2340 (N_2340,In_730,In_975);
nand U2341 (N_2341,In_505,In_175);
nor U2342 (N_2342,In_488,In_470);
or U2343 (N_2343,In_123,In_860);
nor U2344 (N_2344,In_488,In_153);
and U2345 (N_2345,In_725,In_936);
nand U2346 (N_2346,In_512,In_892);
or U2347 (N_2347,In_436,In_45);
or U2348 (N_2348,In_465,In_162);
and U2349 (N_2349,In_370,In_263);
xor U2350 (N_2350,In_426,In_513);
and U2351 (N_2351,In_902,In_465);
xor U2352 (N_2352,In_291,In_569);
nand U2353 (N_2353,In_388,In_435);
or U2354 (N_2354,In_196,In_156);
and U2355 (N_2355,In_974,In_191);
or U2356 (N_2356,In_657,In_334);
nor U2357 (N_2357,In_663,In_103);
nand U2358 (N_2358,In_356,In_573);
nor U2359 (N_2359,In_238,In_286);
or U2360 (N_2360,In_427,In_661);
or U2361 (N_2361,In_222,In_117);
nand U2362 (N_2362,In_381,In_896);
or U2363 (N_2363,In_582,In_785);
xnor U2364 (N_2364,In_713,In_914);
nand U2365 (N_2365,In_175,In_680);
xnor U2366 (N_2366,In_137,In_578);
and U2367 (N_2367,In_26,In_570);
nand U2368 (N_2368,In_167,In_567);
nand U2369 (N_2369,In_487,In_168);
or U2370 (N_2370,In_631,In_786);
xnor U2371 (N_2371,In_983,In_263);
xnor U2372 (N_2372,In_47,In_820);
nor U2373 (N_2373,In_136,In_939);
or U2374 (N_2374,In_780,In_291);
and U2375 (N_2375,In_526,In_360);
or U2376 (N_2376,In_416,In_235);
and U2377 (N_2377,In_804,In_293);
and U2378 (N_2378,In_717,In_391);
or U2379 (N_2379,In_171,In_817);
xnor U2380 (N_2380,In_593,In_505);
nand U2381 (N_2381,In_266,In_307);
nand U2382 (N_2382,In_842,In_771);
xor U2383 (N_2383,In_527,In_311);
and U2384 (N_2384,In_464,In_665);
nor U2385 (N_2385,In_192,In_596);
and U2386 (N_2386,In_997,In_964);
xor U2387 (N_2387,In_308,In_862);
nor U2388 (N_2388,In_847,In_542);
xnor U2389 (N_2389,In_362,In_843);
nor U2390 (N_2390,In_604,In_330);
and U2391 (N_2391,In_69,In_690);
or U2392 (N_2392,In_831,In_881);
nand U2393 (N_2393,In_982,In_603);
xnor U2394 (N_2394,In_956,In_569);
nand U2395 (N_2395,In_434,In_875);
nor U2396 (N_2396,In_552,In_580);
or U2397 (N_2397,In_285,In_535);
nand U2398 (N_2398,In_679,In_454);
xor U2399 (N_2399,In_838,In_651);
nand U2400 (N_2400,In_167,In_249);
xor U2401 (N_2401,In_574,In_681);
nor U2402 (N_2402,In_465,In_75);
or U2403 (N_2403,In_257,In_743);
xnor U2404 (N_2404,In_140,In_540);
nor U2405 (N_2405,In_879,In_688);
nand U2406 (N_2406,In_131,In_595);
xnor U2407 (N_2407,In_152,In_92);
xor U2408 (N_2408,In_354,In_321);
or U2409 (N_2409,In_220,In_110);
nor U2410 (N_2410,In_149,In_146);
nand U2411 (N_2411,In_949,In_683);
or U2412 (N_2412,In_742,In_146);
xnor U2413 (N_2413,In_736,In_160);
nand U2414 (N_2414,In_610,In_233);
nor U2415 (N_2415,In_665,In_409);
or U2416 (N_2416,In_431,In_563);
nand U2417 (N_2417,In_60,In_546);
and U2418 (N_2418,In_842,In_69);
nor U2419 (N_2419,In_832,In_65);
nor U2420 (N_2420,In_559,In_761);
or U2421 (N_2421,In_125,In_461);
xnor U2422 (N_2422,In_315,In_506);
or U2423 (N_2423,In_822,In_37);
nor U2424 (N_2424,In_169,In_39);
or U2425 (N_2425,In_265,In_924);
and U2426 (N_2426,In_137,In_603);
or U2427 (N_2427,In_31,In_547);
nor U2428 (N_2428,In_733,In_104);
nor U2429 (N_2429,In_144,In_966);
xor U2430 (N_2430,In_529,In_453);
nand U2431 (N_2431,In_257,In_638);
nand U2432 (N_2432,In_225,In_423);
and U2433 (N_2433,In_154,In_316);
or U2434 (N_2434,In_2,In_20);
xnor U2435 (N_2435,In_961,In_899);
xnor U2436 (N_2436,In_167,In_951);
and U2437 (N_2437,In_433,In_438);
xnor U2438 (N_2438,In_840,In_488);
or U2439 (N_2439,In_908,In_418);
xor U2440 (N_2440,In_131,In_231);
nand U2441 (N_2441,In_665,In_250);
xnor U2442 (N_2442,In_45,In_541);
nand U2443 (N_2443,In_396,In_173);
and U2444 (N_2444,In_716,In_939);
nand U2445 (N_2445,In_730,In_99);
or U2446 (N_2446,In_730,In_256);
and U2447 (N_2447,In_952,In_268);
nor U2448 (N_2448,In_996,In_176);
nand U2449 (N_2449,In_138,In_11);
nor U2450 (N_2450,In_404,In_794);
or U2451 (N_2451,In_100,In_704);
and U2452 (N_2452,In_214,In_9);
nor U2453 (N_2453,In_921,In_166);
xnor U2454 (N_2454,In_163,In_778);
nor U2455 (N_2455,In_891,In_651);
and U2456 (N_2456,In_135,In_300);
xnor U2457 (N_2457,In_85,In_933);
nand U2458 (N_2458,In_992,In_217);
and U2459 (N_2459,In_940,In_935);
xnor U2460 (N_2460,In_724,In_626);
or U2461 (N_2461,In_359,In_735);
xnor U2462 (N_2462,In_603,In_178);
nand U2463 (N_2463,In_193,In_248);
nor U2464 (N_2464,In_128,In_365);
or U2465 (N_2465,In_50,In_191);
xor U2466 (N_2466,In_205,In_856);
or U2467 (N_2467,In_776,In_25);
nand U2468 (N_2468,In_946,In_641);
nand U2469 (N_2469,In_547,In_422);
nor U2470 (N_2470,In_74,In_349);
nand U2471 (N_2471,In_946,In_495);
nor U2472 (N_2472,In_263,In_767);
nor U2473 (N_2473,In_196,In_783);
nand U2474 (N_2474,In_161,In_518);
nand U2475 (N_2475,In_317,In_352);
or U2476 (N_2476,In_82,In_525);
xor U2477 (N_2477,In_756,In_755);
nand U2478 (N_2478,In_455,In_643);
and U2479 (N_2479,In_682,In_16);
nor U2480 (N_2480,In_764,In_688);
xnor U2481 (N_2481,In_82,In_946);
xnor U2482 (N_2482,In_24,In_51);
and U2483 (N_2483,In_689,In_311);
and U2484 (N_2484,In_879,In_742);
nand U2485 (N_2485,In_154,In_87);
or U2486 (N_2486,In_485,In_531);
xnor U2487 (N_2487,In_778,In_377);
nand U2488 (N_2488,In_700,In_516);
nor U2489 (N_2489,In_212,In_151);
xnor U2490 (N_2490,In_203,In_494);
nor U2491 (N_2491,In_824,In_431);
or U2492 (N_2492,In_451,In_953);
xnor U2493 (N_2493,In_729,In_822);
nor U2494 (N_2494,In_682,In_755);
nand U2495 (N_2495,In_193,In_765);
and U2496 (N_2496,In_868,In_808);
or U2497 (N_2497,In_629,In_920);
or U2498 (N_2498,In_317,In_247);
nor U2499 (N_2499,In_860,In_686);
xnor U2500 (N_2500,N_1289,N_1736);
nor U2501 (N_2501,N_1896,N_1986);
and U2502 (N_2502,N_1365,N_1115);
and U2503 (N_2503,N_528,N_1313);
and U2504 (N_2504,N_1058,N_616);
nand U2505 (N_2505,N_1048,N_1708);
nor U2506 (N_2506,N_26,N_594);
and U2507 (N_2507,N_1245,N_1966);
and U2508 (N_2508,N_409,N_2091);
or U2509 (N_2509,N_1588,N_724);
nand U2510 (N_2510,N_1276,N_1807);
nor U2511 (N_2511,N_1603,N_1013);
or U2512 (N_2512,N_1952,N_2161);
nor U2513 (N_2513,N_1817,N_62);
xor U2514 (N_2514,N_890,N_778);
nand U2515 (N_2515,N_1546,N_2129);
and U2516 (N_2516,N_913,N_991);
and U2517 (N_2517,N_2344,N_767);
xor U2518 (N_2518,N_96,N_741);
or U2519 (N_2519,N_1785,N_1002);
nor U2520 (N_2520,N_153,N_898);
nand U2521 (N_2521,N_276,N_609);
and U2522 (N_2522,N_675,N_2094);
nand U2523 (N_2523,N_136,N_1090);
xor U2524 (N_2524,N_2496,N_2082);
nand U2525 (N_2525,N_1455,N_1052);
or U2526 (N_2526,N_1252,N_1995);
or U2527 (N_2527,N_444,N_975);
nand U2528 (N_2528,N_259,N_1357);
nand U2529 (N_2529,N_760,N_2202);
or U2530 (N_2530,N_1571,N_623);
or U2531 (N_2531,N_2440,N_1471);
nor U2532 (N_2532,N_2273,N_1403);
or U2533 (N_2533,N_173,N_1866);
xnor U2534 (N_2534,N_422,N_2302);
xnor U2535 (N_2535,N_1159,N_1776);
xnor U2536 (N_2536,N_1713,N_1521);
nand U2537 (N_2537,N_80,N_909);
xor U2538 (N_2538,N_2035,N_1229);
nand U2539 (N_2539,N_1574,N_1172);
and U2540 (N_2540,N_780,N_2461);
xor U2541 (N_2541,N_1110,N_994);
and U2542 (N_2542,N_1767,N_2016);
nor U2543 (N_2543,N_2296,N_227);
nor U2544 (N_2544,N_1270,N_2128);
and U2545 (N_2545,N_2348,N_2441);
nand U2546 (N_2546,N_1747,N_919);
and U2547 (N_2547,N_1044,N_556);
and U2548 (N_2548,N_1806,N_2414);
or U2549 (N_2549,N_2422,N_251);
xor U2550 (N_2550,N_4,N_1870);
or U2551 (N_2551,N_1724,N_1146);
or U2552 (N_2552,N_606,N_2474);
nand U2553 (N_2553,N_216,N_997);
xor U2554 (N_2554,N_639,N_1749);
nor U2555 (N_2555,N_1005,N_1491);
and U2556 (N_2556,N_580,N_375);
xor U2557 (N_2557,N_2339,N_1194);
nor U2558 (N_2558,N_228,N_1390);
and U2559 (N_2559,N_957,N_2485);
and U2560 (N_2560,N_1963,N_42);
and U2561 (N_2561,N_10,N_1371);
xnor U2562 (N_2562,N_1716,N_1913);
and U2563 (N_2563,N_236,N_2154);
xnor U2564 (N_2564,N_870,N_2290);
or U2565 (N_2565,N_396,N_2194);
nand U2566 (N_2566,N_1853,N_1445);
or U2567 (N_2567,N_1352,N_1812);
and U2568 (N_2568,N_1466,N_2173);
or U2569 (N_2569,N_186,N_1797);
and U2570 (N_2570,N_1225,N_1184);
nand U2571 (N_2571,N_2018,N_1326);
or U2572 (N_2572,N_1780,N_493);
xor U2573 (N_2573,N_813,N_1862);
nand U2574 (N_2574,N_550,N_497);
nor U2575 (N_2575,N_2151,N_1856);
and U2576 (N_2576,N_2253,N_821);
and U2577 (N_2577,N_1869,N_1486);
and U2578 (N_2578,N_1458,N_1338);
or U2579 (N_2579,N_2079,N_1965);
or U2580 (N_2580,N_1924,N_1155);
nor U2581 (N_2581,N_2355,N_1317);
nand U2582 (N_2582,N_2384,N_895);
nand U2583 (N_2583,N_822,N_1507);
xnor U2584 (N_2584,N_374,N_769);
nand U2585 (N_2585,N_2388,N_281);
xor U2586 (N_2586,N_637,N_103);
nand U2587 (N_2587,N_81,N_1782);
xnor U2588 (N_2588,N_52,N_1889);
and U2589 (N_2589,N_827,N_363);
nand U2590 (N_2590,N_1114,N_17);
nor U2591 (N_2591,N_1695,N_768);
and U2592 (N_2592,N_845,N_1787);
and U2593 (N_2593,N_1144,N_321);
and U2594 (N_2594,N_250,N_2421);
and U2595 (N_2595,N_783,N_1875);
and U2596 (N_2596,N_702,N_1982);
nand U2597 (N_2597,N_55,N_810);
xor U2598 (N_2598,N_917,N_735);
or U2599 (N_2599,N_2375,N_2434);
or U2600 (N_2600,N_1468,N_534);
nor U2601 (N_2601,N_428,N_607);
and U2602 (N_2602,N_2244,N_1926);
nor U2603 (N_2603,N_888,N_1474);
nand U2604 (N_2604,N_468,N_586);
and U2605 (N_2605,N_722,N_1582);
xor U2606 (N_2606,N_1720,N_2373);
nand U2607 (N_2607,N_1070,N_1441);
xnor U2608 (N_2608,N_1666,N_1388);
nor U2609 (N_2609,N_1062,N_1630);
nand U2610 (N_2610,N_535,N_345);
nand U2611 (N_2611,N_1904,N_327);
xor U2612 (N_2612,N_2424,N_1795);
nor U2613 (N_2613,N_1631,N_201);
or U2614 (N_2614,N_1948,N_48);
nand U2615 (N_2615,N_1804,N_2451);
and U2616 (N_2616,N_1580,N_1688);
nand U2617 (N_2617,N_430,N_2241);
nor U2618 (N_2618,N_1814,N_383);
or U2619 (N_2619,N_1949,N_1894);
or U2620 (N_2620,N_1000,N_825);
and U2621 (N_2621,N_817,N_2191);
nor U2622 (N_2622,N_588,N_1673);
and U2623 (N_2623,N_1855,N_2051);
or U2624 (N_2624,N_410,N_2398);
or U2625 (N_2625,N_2300,N_2317);
nand U2626 (N_2626,N_877,N_764);
nor U2627 (N_2627,N_1642,N_1009);
or U2628 (N_2628,N_356,N_501);
or U2629 (N_2629,N_464,N_1880);
or U2630 (N_2630,N_116,N_2392);
and U2631 (N_2631,N_1260,N_1698);
xnor U2632 (N_2632,N_57,N_656);
nand U2633 (N_2633,N_2370,N_1246);
and U2634 (N_2634,N_1548,N_1001);
or U2635 (N_2635,N_1811,N_297);
nand U2636 (N_2636,N_1101,N_1535);
xor U2637 (N_2637,N_1956,N_1779);
xor U2638 (N_2638,N_642,N_1784);
or U2639 (N_2639,N_1874,N_98);
or U2640 (N_2640,N_923,N_2040);
and U2641 (N_2641,N_1938,N_217);
or U2642 (N_2642,N_630,N_266);
or U2643 (N_2643,N_2219,N_2141);
nor U2644 (N_2644,N_645,N_482);
and U2645 (N_2645,N_102,N_1692);
or U2646 (N_2646,N_564,N_2104);
xnor U2647 (N_2647,N_1353,N_1653);
nand U2648 (N_2648,N_91,N_2420);
nor U2649 (N_2649,N_1136,N_1424);
or U2650 (N_2650,N_1450,N_2369);
nor U2651 (N_2651,N_536,N_322);
xor U2652 (N_2652,N_2307,N_1263);
nor U2653 (N_2653,N_2319,N_2447);
nand U2654 (N_2654,N_1061,N_1211);
xor U2655 (N_2655,N_912,N_1722);
nor U2656 (N_2656,N_222,N_1657);
or U2657 (N_2657,N_859,N_70);
and U2658 (N_2658,N_2301,N_474);
xnor U2659 (N_2659,N_1757,N_2119);
or U2660 (N_2660,N_1689,N_677);
or U2661 (N_2661,N_734,N_1074);
or U2662 (N_2662,N_940,N_1640);
nor U2663 (N_2663,N_53,N_242);
xnor U2664 (N_2664,N_2397,N_1867);
and U2665 (N_2665,N_1872,N_1564);
xnor U2666 (N_2666,N_2145,N_2257);
and U2667 (N_2667,N_2405,N_1930);
nor U2668 (N_2668,N_969,N_1342);
nor U2669 (N_2669,N_1515,N_1834);
and U2670 (N_2670,N_1555,N_584);
nor U2671 (N_2671,N_234,N_1557);
nor U2672 (N_2672,N_124,N_1402);
nand U2673 (N_2673,N_519,N_350);
nand U2674 (N_2674,N_690,N_2146);
nand U2675 (N_2675,N_589,N_1614);
nand U2676 (N_2676,N_868,N_1199);
or U2677 (N_2677,N_2395,N_2069);
and U2678 (N_2678,N_1361,N_1024);
or U2679 (N_2679,N_1764,N_1479);
xor U2680 (N_2680,N_43,N_665);
or U2681 (N_2681,N_1873,N_2499);
or U2682 (N_2682,N_2498,N_604);
and U2683 (N_2683,N_1607,N_527);
nand U2684 (N_2684,N_502,N_233);
or U2685 (N_2685,N_469,N_833);
nor U2686 (N_2686,N_158,N_567);
xor U2687 (N_2687,N_1054,N_971);
nand U2688 (N_2688,N_782,N_964);
nor U2689 (N_2689,N_111,N_1355);
xnor U2690 (N_2690,N_2366,N_432);
or U2691 (N_2691,N_1796,N_621);
nand U2692 (N_2692,N_1594,N_1824);
or U2693 (N_2693,N_654,N_1026);
or U2694 (N_2694,N_1432,N_988);
or U2695 (N_2695,N_2433,N_1368);
nand U2696 (N_2696,N_1803,N_1297);
and U2697 (N_2697,N_1818,N_230);
nand U2698 (N_2698,N_50,N_754);
xnor U2699 (N_2699,N_2013,N_2214);
nand U2700 (N_2700,N_277,N_808);
and U2701 (N_2701,N_1208,N_2014);
nand U2702 (N_2702,N_2134,N_1775);
and U2703 (N_2703,N_532,N_2256);
nor U2704 (N_2704,N_1156,N_379);
and U2705 (N_2705,N_1298,N_487);
or U2706 (N_2706,N_1623,N_2320);
xnor U2707 (N_2707,N_459,N_169);
nor U2708 (N_2708,N_1007,N_318);
nand U2709 (N_2709,N_662,N_245);
xnor U2710 (N_2710,N_800,N_424);
or U2711 (N_2711,N_1404,N_498);
nor U2712 (N_2712,N_2218,N_1228);
nor U2713 (N_2713,N_849,N_2403);
nand U2714 (N_2714,N_2316,N_548);
nor U2715 (N_2715,N_1016,N_1900);
nor U2716 (N_2716,N_1838,N_1373);
or U2717 (N_2717,N_1508,N_184);
nor U2718 (N_2718,N_613,N_147);
nor U2719 (N_2719,N_926,N_271);
nor U2720 (N_2720,N_1964,N_771);
nor U2721 (N_2721,N_161,N_1978);
xnor U2722 (N_2722,N_1127,N_2329);
or U2723 (N_2723,N_2185,N_1004);
nand U2724 (N_2724,N_1946,N_811);
nor U2725 (N_2725,N_2401,N_33);
xnor U2726 (N_2726,N_1847,N_466);
and U2727 (N_2727,N_1751,N_2205);
xor U2728 (N_2728,N_110,N_1358);
nor U2729 (N_2729,N_2153,N_602);
or U2730 (N_2730,N_2081,N_698);
or U2731 (N_2731,N_2155,N_1088);
or U2732 (N_2732,N_807,N_2111);
nand U2733 (N_2733,N_1791,N_2043);
and U2734 (N_2734,N_2342,N_1008);
nor U2735 (N_2735,N_457,N_2176);
nand U2736 (N_2736,N_775,N_1029);
nor U2737 (N_2737,N_992,N_1268);
nor U2738 (N_2738,N_23,N_191);
nand U2739 (N_2739,N_1844,N_1711);
nand U2740 (N_2740,N_1768,N_2026);
and U2741 (N_2741,N_911,N_2450);
or U2742 (N_2742,N_830,N_1379);
nand U2743 (N_2743,N_2105,N_1031);
nor U2744 (N_2744,N_2167,N_2462);
nand U2745 (N_2745,N_590,N_585);
or U2746 (N_2746,N_353,N_1370);
xor U2747 (N_2747,N_2318,N_265);
and U2748 (N_2748,N_2232,N_143);
xnor U2749 (N_2749,N_1858,N_1382);
nor U2750 (N_2750,N_842,N_720);
and U2751 (N_2751,N_303,N_2458);
or U2752 (N_2752,N_1735,N_24);
or U2753 (N_2753,N_2124,N_1124);
nor U2754 (N_2754,N_1163,N_1612);
or U2755 (N_2755,N_875,N_2243);
xnor U2756 (N_2756,N_1097,N_1089);
or U2757 (N_2757,N_47,N_1221);
and U2758 (N_2758,N_932,N_1798);
and U2759 (N_2759,N_1710,N_406);
nor U2760 (N_2760,N_1399,N_514);
nand U2761 (N_2761,N_2275,N_1160);
nor U2762 (N_2762,N_1686,N_2266);
nor U2763 (N_2763,N_13,N_533);
nor U2764 (N_2764,N_892,N_500);
or U2765 (N_2765,N_786,N_829);
and U2766 (N_2766,N_712,N_508);
nor U2767 (N_2767,N_1534,N_543);
or U2768 (N_2768,N_2,N_2295);
and U2769 (N_2769,N_641,N_1408);
xnor U2770 (N_2770,N_75,N_1635);
nand U2771 (N_2771,N_905,N_1);
nand U2772 (N_2772,N_2235,N_382);
xor U2773 (N_2773,N_2140,N_2431);
nor U2774 (N_2774,N_1075,N_688);
xnor U2775 (N_2775,N_1456,N_1602);
or U2776 (N_2776,N_1691,N_2123);
and U2777 (N_2777,N_1091,N_2265);
nand U2778 (N_2778,N_312,N_416);
or U2779 (N_2779,N_1674,N_2239);
or U2780 (N_2780,N_1381,N_1618);
nor U2781 (N_2781,N_2207,N_1893);
xnor U2782 (N_2782,N_1042,N_127);
or U2783 (N_2783,N_253,N_706);
nand U2784 (N_2784,N_5,N_2473);
nor U2785 (N_2785,N_206,N_388);
nand U2786 (N_2786,N_324,N_2263);
and U2787 (N_2787,N_581,N_935);
nor U2788 (N_2788,N_1319,N_1970);
or U2789 (N_2789,N_1516,N_1047);
nand U2790 (N_2790,N_1830,N_1422);
nand U2791 (N_2791,N_1218,N_1117);
and U2792 (N_2792,N_38,N_816);
and U2793 (N_2793,N_1011,N_343);
xnor U2794 (N_2794,N_790,N_1933);
and U2795 (N_2795,N_1559,N_572);
nand U2796 (N_2796,N_1286,N_105);
xor U2797 (N_2797,N_2228,N_1315);
xnor U2798 (N_2798,N_2245,N_1067);
and U2799 (N_2799,N_707,N_2330);
xnor U2800 (N_2800,N_2357,N_2116);
nand U2801 (N_2801,N_1200,N_1071);
or U2802 (N_2802,N_2197,N_294);
nor U2803 (N_2803,N_1230,N_1027);
nor U2804 (N_2804,N_1185,N_540);
xnor U2805 (N_2805,N_2053,N_2097);
xnor U2806 (N_2806,N_1277,N_58);
or U2807 (N_2807,N_1278,N_2314);
nor U2808 (N_2808,N_1821,N_1079);
xor U2809 (N_2809,N_1659,N_1620);
nand U2810 (N_2810,N_1741,N_319);
nor U2811 (N_2811,N_729,N_2101);
and U2812 (N_2812,N_126,N_1799);
and U2813 (N_2813,N_862,N_2432);
or U2814 (N_2814,N_974,N_595);
and U2815 (N_2815,N_339,N_2138);
xnor U2816 (N_2816,N_2203,N_652);
nand U2817 (N_2817,N_1738,N_2147);
and U2818 (N_2818,N_1261,N_1714);
and U2819 (N_2819,N_192,N_1754);
xnor U2820 (N_2820,N_561,N_2063);
nand U2821 (N_2821,N_1096,N_1119);
xnor U2822 (N_2822,N_1086,N_880);
nor U2823 (N_2823,N_1452,N_2379);
nand U2824 (N_2824,N_30,N_2274);
xnor U2825 (N_2825,N_743,N_274);
xor U2826 (N_2826,N_462,N_268);
nor U2827 (N_2827,N_505,N_1693);
or U2828 (N_2828,N_411,N_1411);
or U2829 (N_2829,N_162,N_1243);
nand U2830 (N_2830,N_1446,N_97);
and U2831 (N_2831,N_229,N_198);
or U2832 (N_2832,N_655,N_820);
and U2833 (N_2833,N_1364,N_826);
nor U2834 (N_2834,N_349,N_1248);
and U2835 (N_2835,N_824,N_195);
or U2836 (N_2836,N_134,N_60);
nand U2837 (N_2837,N_2287,N_1766);
nor U2838 (N_2838,N_1911,N_762);
nor U2839 (N_2839,N_1529,N_311);
xnor U2840 (N_2840,N_1310,N_865);
nor U2841 (N_2841,N_916,N_455);
and U2842 (N_2842,N_2168,N_755);
xnor U2843 (N_2843,N_215,N_1921);
nor U2844 (N_2844,N_2071,N_948);
xor U2845 (N_2845,N_9,N_939);
nand U2846 (N_2846,N_2072,N_333);
or U2847 (N_2847,N_579,N_732);
nor U2848 (N_2848,N_2048,N_1406);
and U2849 (N_2849,N_1863,N_335);
or U2850 (N_2850,N_618,N_360);
or U2851 (N_2851,N_1916,N_2312);
and U2852 (N_2852,N_273,N_1374);
or U2853 (N_2853,N_2471,N_1316);
nor U2854 (N_2854,N_1238,N_1461);
nor U2855 (N_2855,N_1250,N_1483);
and U2856 (N_2856,N_560,N_1519);
and U2857 (N_2857,N_2130,N_575);
nand U2858 (N_2858,N_1759,N_856);
nor U2859 (N_2859,N_750,N_1280);
xor U2860 (N_2860,N_2127,N_113);
or U2861 (N_2861,N_2327,N_1920);
and U2862 (N_2862,N_1457,N_78);
nor U2863 (N_2863,N_243,N_1919);
xor U2864 (N_2864,N_1178,N_366);
and U2865 (N_2865,N_2046,N_2261);
nand U2866 (N_2866,N_264,N_1849);
nor U2867 (N_2867,N_2436,N_114);
nand U2868 (N_2868,N_1961,N_1544);
xor U2869 (N_2869,N_1646,N_44);
nand U2870 (N_2870,N_7,N_1888);
xnor U2871 (N_2871,N_446,N_1223);
and U2872 (N_2872,N_1667,N_2064);
nor U2873 (N_2873,N_1709,N_1660);
xnor U2874 (N_2874,N_922,N_847);
nor U2875 (N_2875,N_1533,N_1652);
and U2876 (N_2876,N_302,N_1209);
nand U2877 (N_2877,N_1942,N_344);
nand U2878 (N_2878,N_1081,N_320);
nand U2879 (N_2879,N_672,N_612);
xor U2880 (N_2880,N_336,N_1421);
nor U2881 (N_2881,N_673,N_1624);
xnor U2882 (N_2882,N_270,N_2075);
nor U2883 (N_2883,N_1940,N_1416);
and U2884 (N_2884,N_1752,N_1760);
xnor U2885 (N_2885,N_568,N_2426);
nor U2886 (N_2886,N_473,N_1335);
or U2887 (N_2887,N_15,N_730);
nand U2888 (N_2888,N_1586,N_224);
nor U2889 (N_2889,N_983,N_305);
xnor U2890 (N_2890,N_1312,N_1613);
nand U2891 (N_2891,N_2021,N_152);
nand U2892 (N_2892,N_963,N_944);
nand U2893 (N_2893,N_516,N_1939);
nor U2894 (N_2894,N_1340,N_2238);
xnor U2895 (N_2895,N_2309,N_1046);
or U2896 (N_2896,N_1309,N_263);
nand U2897 (N_2897,N_1305,N_2445);
and U2898 (N_2898,N_1188,N_331);
nor U2899 (N_2899,N_1407,N_2449);
xor U2900 (N_2900,N_2490,N_232);
and U2901 (N_2901,N_1678,N_1082);
or U2902 (N_2902,N_1448,N_1655);
and U2903 (N_2903,N_758,N_1765);
nand U2904 (N_2904,N_1723,N_381);
xnor U2905 (N_2905,N_1572,N_1690);
nand U2906 (N_2906,N_848,N_2492);
nand U2907 (N_2907,N_194,N_421);
nand U2908 (N_2908,N_1242,N_1628);
nand U2909 (N_2909,N_279,N_565);
and U2910 (N_2910,N_471,N_1839);
or U2911 (N_2911,N_2341,N_1943);
or U2912 (N_2912,N_981,N_1592);
nor U2913 (N_2913,N_2179,N_2083);
or U2914 (N_2914,N_1541,N_1258);
or U2915 (N_2915,N_1384,N_1625);
or U2916 (N_2916,N_1366,N_141);
xor U2917 (N_2917,N_980,N_1427);
nor U2918 (N_2918,N_1816,N_1475);
or U2919 (N_2919,N_1142,N_503);
xnor U2920 (N_2920,N_1443,N_397);
or U2921 (N_2921,N_2269,N_465);
nor U2922 (N_2922,N_1396,N_2429);
nand U2923 (N_2923,N_1861,N_2353);
and U2924 (N_2924,N_2195,N_2484);
nand U2925 (N_2925,N_486,N_918);
nor U2926 (N_2926,N_2036,N_2345);
xnor U2927 (N_2927,N_1099,N_2497);
nor U2928 (N_2928,N_1901,N_1848);
xnor U2929 (N_2929,N_1012,N_1512);
xnor U2930 (N_2930,N_1264,N_2022);
nand U2931 (N_2931,N_2099,N_1526);
or U2932 (N_2932,N_1569,N_289);
or U2933 (N_2933,N_2443,N_2188);
or U2934 (N_2934,N_1189,N_982);
nor U2935 (N_2935,N_1165,N_338);
xor U2936 (N_2936,N_1810,N_2206);
and U2937 (N_2937,N_569,N_2407);
nand U2938 (N_2938,N_66,N_267);
and U2939 (N_2939,N_1898,N_747);
and U2940 (N_2940,N_1887,N_417);
nand U2941 (N_2941,N_2196,N_1173);
nor U2942 (N_2942,N_740,N_77);
and U2943 (N_2943,N_2285,N_2017);
or U2944 (N_2944,N_2204,N_1257);
xor U2945 (N_2945,N_1649,N_1287);
or U2946 (N_2946,N_622,N_2216);
nand U2947 (N_2947,N_1198,N_1739);
xor U2948 (N_2948,N_647,N_1700);
or U2949 (N_2949,N_1318,N_628);
xor U2950 (N_2950,N_524,N_1885);
xnor U2951 (N_2951,N_1573,N_2041);
nor U2952 (N_2952,N_1647,N_2313);
and U2953 (N_2953,N_598,N_235);
nand U2954 (N_2954,N_88,N_28);
xnor U2955 (N_2955,N_239,N_1589);
nand U2956 (N_2956,N_663,N_14);
nor U2957 (N_2957,N_1547,N_958);
nor U2958 (N_2958,N_1068,N_1701);
nand U2959 (N_2959,N_1464,N_391);
or U2960 (N_2960,N_1922,N_1339);
and U2961 (N_2961,N_1899,N_1410);
xor U2962 (N_2962,N_2180,N_1145);
nor U2963 (N_2963,N_342,N_513);
nand U2964 (N_2964,N_970,N_962);
and U2965 (N_2965,N_1356,N_1217);
nand U2966 (N_2966,N_71,N_262);
nand U2967 (N_2967,N_2004,N_1311);
or U2968 (N_2968,N_1324,N_832);
and U2969 (N_2969,N_1300,N_1671);
nand U2970 (N_2970,N_1294,N_34);
nand U2971 (N_2971,N_1419,N_1078);
nor U2972 (N_2972,N_1656,N_1503);
nand U2973 (N_2973,N_1442,N_1362);
nand U2974 (N_2974,N_176,N_171);
or U2975 (N_2975,N_1302,N_2411);
nor U2976 (N_2976,N_2215,N_1219);
xor U2977 (N_2977,N_857,N_678);
and U2978 (N_2978,N_2326,N_121);
xor U2979 (N_2979,N_1345,N_2482);
xnor U2980 (N_2980,N_840,N_838);
xor U2981 (N_2981,N_854,N_2463);
and U2982 (N_2982,N_1267,N_128);
nor U2983 (N_2983,N_700,N_1331);
nor U2984 (N_2984,N_2009,N_19);
xnor U2985 (N_2985,N_1397,N_1805);
or U2986 (N_2986,N_2323,N_633);
nor U2987 (N_2987,N_226,N_1212);
or U2988 (N_2988,N_2371,N_1846);
nand U2989 (N_2989,N_2349,N_853);
and U2990 (N_2990,N_361,N_2280);
or U2991 (N_2991,N_1215,N_65);
and U2992 (N_2992,N_2262,N_1420);
nor U2993 (N_2993,N_879,N_2117);
xor U2994 (N_2994,N_1241,N_313);
nand U2995 (N_2995,N_1262,N_530);
and U2996 (N_2996,N_788,N_139);
or U2997 (N_2997,N_1405,N_2107);
or U2998 (N_2998,N_617,N_325);
nand U2999 (N_2999,N_436,N_1577);
nand U3000 (N_3000,N_183,N_2377);
nor U3001 (N_3001,N_272,N_1850);
xnor U3002 (N_3002,N_546,N_2159);
nor U3003 (N_3003,N_2356,N_597);
and U3004 (N_3004,N_1825,N_2047);
xor U3005 (N_3005,N_2056,N_2058);
xor U3006 (N_3006,N_931,N_2057);
nor U3007 (N_3007,N_2080,N_1327);
nor U3008 (N_3008,N_2025,N_679);
or U3009 (N_3009,N_1727,N_1575);
nand U3010 (N_3010,N_2067,N_525);
nor U3011 (N_3011,N_828,N_300);
and U3012 (N_3012,N_1095,N_1291);
or U3013 (N_3013,N_681,N_1453);
xor U3014 (N_3014,N_1332,N_2142);
nor U3015 (N_3015,N_999,N_1412);
nand U3016 (N_3016,N_341,N_1538);
or U3017 (N_3017,N_987,N_252);
nand U3018 (N_3018,N_2225,N_1003);
nand U3019 (N_3019,N_674,N_1845);
and U3020 (N_3020,N_1354,N_2113);
and U3021 (N_3021,N_1234,N_1487);
nand U3022 (N_3022,N_408,N_18);
or U3023 (N_3023,N_1608,N_1206);
and U3024 (N_3024,N_545,N_1224);
xnor U3025 (N_3025,N_908,N_1932);
nor U3026 (N_3026,N_1186,N_1890);
nand U3027 (N_3027,N_1333,N_1851);
or U3028 (N_3028,N_1039,N_2281);
or U3029 (N_3029,N_1154,N_2231);
or U3030 (N_3030,N_1451,N_1111);
nor U3031 (N_3031,N_643,N_899);
nand U3032 (N_3032,N_275,N_792);
xor U3033 (N_3033,N_897,N_2272);
and U3034 (N_3034,N_2062,N_73);
nand U3035 (N_3035,N_851,N_512);
and U3036 (N_3036,N_1585,N_438);
and U3037 (N_3037,N_1367,N_1414);
nand U3038 (N_3038,N_1860,N_1344);
nand U3039 (N_3039,N_1321,N_1658);
xnor U3040 (N_3040,N_950,N_2054);
xor U3041 (N_3041,N_627,N_2282);
nor U3042 (N_3042,N_1522,N_537);
nor U3043 (N_3043,N_608,N_119);
xnor U3044 (N_3044,N_1231,N_1598);
and U3045 (N_3045,N_1105,N_1937);
or U3046 (N_3046,N_2387,N_2001);
nand U3047 (N_3047,N_518,N_329);
xor U3048 (N_3048,N_1207,N_659);
nor U3049 (N_3049,N_631,N_2045);
or U3050 (N_3050,N_1944,N_2220);
nand U3051 (N_3051,N_1122,N_1034);
or U3052 (N_3052,N_2031,N_779);
nand U3053 (N_3053,N_803,N_651);
nor U3054 (N_3054,N_1728,N_891);
or U3055 (N_3055,N_2166,N_910);
nand U3056 (N_3056,N_2133,N_667);
nand U3057 (N_3057,N_1721,N_2255);
or U3058 (N_3058,N_731,N_1014);
or U3059 (N_3059,N_1369,N_2034);
and U3060 (N_3060,N_442,N_1543);
or U3061 (N_3061,N_626,N_1663);
nand U3062 (N_3062,N_317,N_1259);
nand U3063 (N_3063,N_140,N_881);
and U3064 (N_3064,N_1501,N_2351);
or U3065 (N_3065,N_1152,N_2294);
nand U3066 (N_3066,N_2157,N_115);
or U3067 (N_3067,N_1587,N_959);
nand U3068 (N_3068,N_727,N_36);
nand U3069 (N_3069,N_1553,N_2270);
nand U3070 (N_3070,N_714,N_1702);
xnor U3071 (N_3071,N_1552,N_1743);
nor U3072 (N_3072,N_573,N_1545);
or U3073 (N_3073,N_1496,N_1195);
nand U3074 (N_3074,N_154,N_1057);
nor U3075 (N_3075,N_1925,N_2494);
or U3076 (N_3076,N_2288,N_2359);
nor U3077 (N_3077,N_2493,N_2334);
nand U3078 (N_3078,N_1567,N_299);
nor U3079 (N_3079,N_2131,N_1174);
xor U3080 (N_3080,N_1891,N_1472);
xnor U3081 (N_3081,N_2007,N_129);
nor U3082 (N_3082,N_814,N_791);
xnor U3083 (N_3083,N_2383,N_197);
nor U3084 (N_3084,N_1980,N_59);
nor U3085 (N_3085,N_2495,N_1147);
and U3086 (N_3086,N_1910,N_189);
xnor U3087 (N_3087,N_2102,N_2417);
and U3088 (N_3088,N_2089,N_1864);
nand U3089 (N_3089,N_701,N_1151);
xor U3090 (N_3090,N_2065,N_2439);
xnor U3091 (N_3091,N_348,N_203);
nor U3092 (N_3092,N_1629,N_1697);
and U3093 (N_3093,N_1109,N_1394);
nor U3094 (N_3094,N_109,N_310);
or U3095 (N_3095,N_2201,N_521);
or U3096 (N_3096,N_1328,N_247);
xnor U3097 (N_3097,N_1049,N_934);
and U3098 (N_3098,N_1755,N_1134);
nand U3099 (N_3099,N_570,N_288);
and U3100 (N_3100,N_2283,N_1684);
xnor U3101 (N_3101,N_223,N_2399);
or U3102 (N_3102,N_2110,N_1777);
or U3103 (N_3103,N_304,N_1597);
nor U3104 (N_3104,N_1123,N_1732);
or U3105 (N_3105,N_159,N_753);
nor U3106 (N_3106,N_795,N_1244);
nand U3107 (N_3107,N_2077,N_1072);
and U3108 (N_3108,N_924,N_1447);
nand U3109 (N_3109,N_1578,N_2435);
nand U3110 (N_3110,N_2049,N_238);
xnor U3111 (N_3111,N_1758,N_1974);
nor U3112 (N_3112,N_285,N_1917);
xnor U3113 (N_3113,N_1616,N_1051);
nand U3114 (N_3114,N_592,N_571);
nor U3115 (N_3115,N_2286,N_1950);
nor U3116 (N_3116,N_818,N_125);
xnor U3117 (N_3117,N_1112,N_1540);
and U3118 (N_3118,N_1030,N_1882);
nand U3119 (N_3119,N_46,N_2181);
xnor U3120 (N_3120,N_2000,N_488);
or U3121 (N_3121,N_1737,N_1554);
and U3122 (N_3122,N_1161,N_952);
nor U3123 (N_3123,N_1562,N_1934);
or U3124 (N_3124,N_2242,N_1772);
nand U3125 (N_3125,N_1528,N_1583);
and U3126 (N_3126,N_2310,N_2212);
or U3127 (N_3127,N_1984,N_1387);
nor U3128 (N_3128,N_1129,N_1897);
nand U3129 (N_3129,N_12,N_298);
or U3130 (N_3130,N_76,N_2158);
and U3131 (N_3131,N_373,N_2164);
or U3132 (N_3132,N_1744,N_399);
or U3133 (N_3133,N_472,N_649);
and U3134 (N_3134,N_257,N_67);
and U3135 (N_3135,N_772,N_2125);
nand U3136 (N_3136,N_1604,N_308);
nand U3137 (N_3137,N_330,N_1485);
xnor U3138 (N_3138,N_106,N_456);
and U3139 (N_3139,N_2306,N_1610);
xor U3140 (N_3140,N_490,N_2149);
and U3141 (N_3141,N_1638,N_90);
and U3142 (N_3142,N_200,N_405);
nor U3143 (N_3143,N_2086,N_435);
xor U3144 (N_3144,N_749,N_2044);
nor U3145 (N_3145,N_889,N_1376);
nand U3146 (N_3146,N_334,N_1108);
xor U3147 (N_3147,N_1290,N_2118);
or U3148 (N_3148,N_759,N_1835);
nand U3149 (N_3149,N_2224,N_291);
nor U3150 (N_3150,N_693,N_120);
nor U3151 (N_3151,N_1437,N_689);
xor U3152 (N_3152,N_1336,N_711);
and U3153 (N_3153,N_583,N_640);
and U3154 (N_3154,N_812,N_2246);
nor U3155 (N_3155,N_1255,N_1827);
or U3156 (N_3156,N_960,N_933);
or U3157 (N_3157,N_723,N_207);
or U3158 (N_3158,N_156,N_2236);
or U3159 (N_3159,N_669,N_781);
nand U3160 (N_3160,N_2413,N_737);
nand U3161 (N_3161,N_352,N_1304);
or U3162 (N_3162,N_506,N_188);
nor U3163 (N_3163,N_2006,N_1019);
xor U3164 (N_3164,N_458,N_1945);
nand U3165 (N_3165,N_489,N_1135);
or U3166 (N_3166,N_1202,N_2322);
and U3167 (N_3167,N_208,N_2470);
and U3168 (N_3168,N_2343,N_2279);
nand U3169 (N_3169,N_372,N_1531);
and U3170 (N_3170,N_682,N_1928);
and U3171 (N_3171,N_946,N_2475);
and U3172 (N_3172,N_1137,N_2015);
xnor U3173 (N_3173,N_1773,N_1083);
xor U3174 (N_3174,N_1494,N_440);
nand U3175 (N_3175,N_2396,N_1881);
or U3176 (N_3176,N_2175,N_2308);
nor U3177 (N_3177,N_704,N_295);
and U3178 (N_3178,N_2247,N_240);
nand U3179 (N_3179,N_746,N_1314);
nor U3180 (N_3180,N_1465,N_1063);
xnor U3181 (N_3181,N_1831,N_558);
xnor U3182 (N_3182,N_1429,N_2354);
or U3183 (N_3183,N_1823,N_25);
and U3184 (N_3184,N_386,N_2008);
xor U3185 (N_3185,N_2378,N_1975);
and U3186 (N_3186,N_1018,N_1323);
and U3187 (N_3187,N_685,N_151);
xor U3188 (N_3188,N_1505,N_475);
or U3189 (N_3189,N_316,N_713);
nor U3190 (N_3190,N_1842,N_2192);
and U3191 (N_3191,N_1473,N_286);
and U3192 (N_3192,N_2132,N_836);
nor U3193 (N_3193,N_2087,N_148);
nand U3194 (N_3194,N_2174,N_638);
or U3195 (N_3195,N_915,N_831);
xnor U3196 (N_3196,N_2331,N_511);
xor U3197 (N_3197,N_777,N_1232);
nor U3198 (N_3198,N_177,N_1840);
and U3199 (N_3199,N_2088,N_450);
xnor U3200 (N_3200,N_896,N_601);
nand U3201 (N_3201,N_789,N_739);
xnor U3202 (N_3202,N_1687,N_2233);
nor U3203 (N_3203,N_1668,N_929);
and U3204 (N_3204,N_3,N_404);
nor U3205 (N_3205,N_2020,N_549);
or U3206 (N_3206,N_387,N_1788);
nor U3207 (N_3207,N_1477,N_1017);
or U3208 (N_3208,N_1976,N_1010);
xor U3209 (N_3209,N_646,N_426);
or U3210 (N_3210,N_1495,N_85);
nand U3211 (N_3211,N_293,N_2222);
or U3212 (N_3212,N_1157,N_1994);
xor U3213 (N_3213,N_2410,N_582);
and U3214 (N_3214,N_1568,N_1959);
nand U3215 (N_3215,N_2409,N_858);
or U3216 (N_3216,N_1794,N_218);
nand U3217 (N_3217,N_721,N_1045);
nand U3218 (N_3218,N_2183,N_1166);
or U3219 (N_3219,N_2023,N_419);
and U3220 (N_3220,N_1902,N_961);
nor U3221 (N_3221,N_2374,N_1417);
nand U3222 (N_3222,N_2152,N_1783);
nor U3223 (N_3223,N_2213,N_170);
and U3224 (N_3224,N_2260,N_1819);
xnor U3225 (N_3225,N_984,N_531);
and U3226 (N_3226,N_2002,N_1563);
xor U3227 (N_3227,N_1990,N_2381);
xnor U3228 (N_3228,N_1611,N_615);
xor U3229 (N_3229,N_1532,N_146);
and U3230 (N_3230,N_2476,N_1334);
xor U3231 (N_3231,N_1476,N_1274);
nor U3232 (N_3232,N_1969,N_2106);
nor U3233 (N_3233,N_1415,N_1285);
xnor U3234 (N_3234,N_1053,N_1680);
and U3235 (N_3235,N_2284,N_1179);
nor U3236 (N_3236,N_2385,N_1064);
and U3237 (N_3237,N_2454,N_1398);
nand U3238 (N_3238,N_717,N_1036);
xnor U3239 (N_3239,N_2217,N_1346);
nand U3240 (N_3240,N_515,N_185);
nand U3241 (N_3241,N_168,N_2486);
or U3242 (N_3242,N_624,N_855);
or U3243 (N_3243,N_2479,N_256);
nand U3244 (N_3244,N_1833,N_1761);
or U3245 (N_3245,N_763,N_496);
xnor U3246 (N_3246,N_1549,N_1955);
or U3247 (N_3247,N_181,N_996);
and U3248 (N_3248,N_2394,N_979);
and U3249 (N_3249,N_99,N_2208);
nor U3250 (N_3250,N_653,N_1359);
and U3251 (N_3251,N_695,N_1272);
nor U3252 (N_3252,N_359,N_2171);
xor U3253 (N_3253,N_1181,N_2278);
nor U3254 (N_3254,N_1632,N_2361);
xnor U3255 (N_3255,N_668,N_951);
xnor U3256 (N_3256,N_1433,N_599);
and U3257 (N_3257,N_220,N_1028);
xnor U3258 (N_3258,N_412,N_930);
or U3259 (N_3259,N_1183,N_776);
or U3260 (N_3260,N_2199,N_902);
or U3261 (N_3261,N_296,N_365);
or U3262 (N_3262,N_2136,N_989);
xnor U3263 (N_3263,N_736,N_1929);
nor U3264 (N_3264,N_1706,N_846);
nand U3265 (N_3265,N_326,N_2052);
nor U3266 (N_3266,N_925,N_687);
nand U3267 (N_3267,N_2172,N_2416);
and U3268 (N_3268,N_1648,N_2122);
xor U3269 (N_3269,N_1469,N_1705);
or U3270 (N_3270,N_2221,N_2143);
xor U3271 (N_3271,N_1584,N_1085);
nor U3272 (N_3272,N_2019,N_1606);
and U3273 (N_3273,N_332,N_2182);
nor U3274 (N_3274,N_392,N_680);
nand U3275 (N_3275,N_1150,N_914);
and U3276 (N_3276,N_1400,N_1918);
and U3277 (N_3277,N_563,N_133);
and U3278 (N_3278,N_427,N_844);
or U3279 (N_3279,N_611,N_1999);
and U3280 (N_3280,N_2092,N_413);
and U3281 (N_3281,N_1233,N_2060);
and U3282 (N_3282,N_968,N_2325);
nand U3283 (N_3283,N_1214,N_2332);
xor U3284 (N_3284,N_703,N_1988);
or U3285 (N_3285,N_559,N_101);
nor U3286 (N_3286,N_1685,N_1763);
nand U3287 (N_3287,N_2120,N_258);
nand U3288 (N_3288,N_1789,N_144);
nor U3289 (N_3289,N_1985,N_2400);
and U3290 (N_3290,N_774,N_2249);
or U3291 (N_3291,N_79,N_784);
or U3292 (N_3292,N_2186,N_562);
xor U3293 (N_3293,N_873,N_625);
or U3294 (N_3294,N_449,N_977);
nor U3295 (N_3295,N_1193,N_1670);
xor U3296 (N_3296,N_84,N_2210);
or U3297 (N_3297,N_708,N_2271);
or U3298 (N_3298,N_1282,N_1240);
or U3299 (N_3299,N_671,N_1912);
and U3300 (N_3300,N_1717,N_2068);
nor U3301 (N_3301,N_1936,N_1470);
nor U3302 (N_3302,N_603,N_799);
and U3303 (N_3303,N_309,N_1162);
xnor U3304 (N_3304,N_928,N_255);
nand U3305 (N_3305,N_819,N_1401);
or U3306 (N_3306,N_1140,N_1800);
or U3307 (N_3307,N_1661,N_1871);
nor U3308 (N_3308,N_2466,N_2304);
nand U3309 (N_3309,N_2472,N_1149);
xnor U3310 (N_3310,N_2382,N_45);
nand U3311 (N_3311,N_1377,N_2084);
and U3312 (N_3312,N_32,N_1192);
nand U3313 (N_3313,N_1973,N_942);
nand U3314 (N_3314,N_1251,N_1941);
xnor U3315 (N_3315,N_943,N_1622);
or U3316 (N_3316,N_1694,N_429);
or U3317 (N_3317,N_2003,N_346);
nand U3318 (N_3318,N_1906,N_433);
nand U3319 (N_3319,N_2250,N_2070);
nor U3320 (N_3320,N_1914,N_112);
nor U3321 (N_3321,N_794,N_2139);
or U3322 (N_3322,N_2362,N_1383);
or U3323 (N_3323,N_448,N_691);
xor U3324 (N_3324,N_1813,N_2095);
or U3325 (N_3325,N_1459,N_871);
xnor U3326 (N_3326,N_1363,N_635);
nor U3327 (N_3327,N_481,N_1645);
nand U3328 (N_3328,N_2055,N_1762);
xor U3329 (N_3329,N_1550,N_415);
nor U3330 (N_3330,N_664,N_2448);
nand U3331 (N_3331,N_1141,N_254);
nor U3332 (N_3332,N_2226,N_591);
nor U3333 (N_3333,N_1015,N_2011);
and U3334 (N_3334,N_2193,N_1467);
or U3335 (N_3335,N_1636,N_1704);
or U3336 (N_3336,N_248,N_876);
nor U3337 (N_3337,N_2162,N_1391);
nand U3338 (N_3338,N_2457,N_1490);
or U3339 (N_3339,N_1627,N_1820);
and U3340 (N_3340,N_1740,N_2277);
nand U3341 (N_3341,N_577,N_1774);
and U3342 (N_3342,N_1118,N_2163);
nor U3343 (N_3343,N_213,N_1197);
xnor U3344 (N_3344,N_670,N_1478);
and U3345 (N_3345,N_2050,N_1092);
nand U3346 (N_3346,N_802,N_600);
and U3347 (N_3347,N_1841,N_1983);
nor U3348 (N_3348,N_709,N_1423);
nand U3349 (N_3349,N_956,N_1669);
nor U3350 (N_3350,N_418,N_1293);
nor U3351 (N_3351,N_1069,N_1525);
or U3352 (N_3352,N_2333,N_1664);
or U3353 (N_3353,N_149,N_1822);
nor U3354 (N_3354,N_400,N_938);
and U3355 (N_3355,N_1672,N_447);
or U3356 (N_3356,N_64,N_2030);
nor U3357 (N_3357,N_632,N_1915);
or U3358 (N_3358,N_823,N_2404);
nor U3359 (N_3359,N_804,N_2074);
and U3360 (N_3360,N_1271,N_1745);
or U3361 (N_3361,N_2419,N_553);
or U3362 (N_3362,N_504,N_715);
nor U3363 (N_3363,N_596,N_2418);
nor U3364 (N_3364,N_82,N_993);
or U3365 (N_3365,N_402,N_165);
nor U3366 (N_3366,N_2338,N_1537);
or U3367 (N_3367,N_941,N_1322);
or U3368 (N_3368,N_2364,N_1499);
xnor U3369 (N_3369,N_998,N_100);
nand U3370 (N_3370,N_439,N_2187);
and U3371 (N_3371,N_477,N_1284);
and U3372 (N_3372,N_2363,N_1056);
or U3373 (N_3373,N_1125,N_407);
xor U3374 (N_3374,N_1348,N_1484);
and U3375 (N_3375,N_2390,N_182);
nor U3376 (N_3376,N_131,N_1536);
xor U3377 (N_3377,N_1650,N_2352);
or U3378 (N_3378,N_122,N_882);
and U3379 (N_3379,N_2252,N_2478);
and U3380 (N_3380,N_209,N_2135);
or U3381 (N_3381,N_538,N_1038);
nand U3382 (N_3382,N_1527,N_22);
nand U3383 (N_3383,N_2459,N_878);
and U3384 (N_3384,N_976,N_1449);
nor U3385 (N_3385,N_437,N_11);
or U3386 (N_3386,N_2264,N_2427);
and U3387 (N_3387,N_290,N_2469);
nor U3388 (N_3388,N_973,N_2037);
nand U3389 (N_3389,N_2340,N_2229);
nand U3390 (N_3390,N_699,N_1033);
nand U3391 (N_3391,N_1132,N_21);
nand U3392 (N_3392,N_869,N_834);
and U3393 (N_3393,N_2465,N_1201);
nor U3394 (N_3394,N_936,N_557);
nand U3395 (N_3395,N_2438,N_2251);
nand U3396 (N_3396,N_2368,N_1247);
or U3397 (N_3397,N_1809,N_1094);
and U3398 (N_3398,N_1981,N_2032);
nor U3399 (N_3399,N_2085,N_692);
or U3400 (N_3400,N_2005,N_1249);
and U3401 (N_3401,N_990,N_1059);
or U3402 (N_3402,N_1107,N_2098);
nor U3403 (N_3403,N_1393,N_180);
xor U3404 (N_3404,N_2024,N_2358);
or U3405 (N_3405,N_644,N_1216);
or U3406 (N_3406,N_395,N_1596);
nand U3407 (N_3407,N_1210,N_850);
nor U3408 (N_3408,N_1164,N_1222);
xor U3409 (N_3409,N_966,N_340);
nor U3410 (N_3410,N_2305,N_1256);
or U3411 (N_3411,N_2169,N_451);
nor U3412 (N_3412,N_765,N_2428);
or U3413 (N_3413,N_1182,N_2012);
xnor U3414 (N_3414,N_460,N_554);
or U3415 (N_3415,N_1993,N_138);
and U3416 (N_3416,N_1865,N_864);
and U3417 (N_3417,N_1350,N_796);
nand U3418 (N_3418,N_1953,N_1380);
xor U3419 (N_3419,N_967,N_1227);
and U3420 (N_3420,N_118,N_108);
nor U3421 (N_3421,N_1177,N_1303);
nand U3422 (N_3422,N_86,N_403);
nor U3423 (N_3423,N_1619,N_470);
nor U3424 (N_3424,N_1205,N_20);
or U3425 (N_3425,N_2346,N_1022);
xor U3426 (N_3426,N_1121,N_1306);
nor U3427 (N_3427,N_199,N_752);
nand U3428 (N_3428,N_2078,N_246);
and U3429 (N_3429,N_1020,N_1876);
and U3430 (N_3430,N_269,N_541);
nand U3431 (N_3431,N_2491,N_1504);
and U3432 (N_3432,N_1637,N_526);
and U3433 (N_3433,N_1778,N_1428);
or U3434 (N_3434,N_797,N_378);
xnor U3435 (N_3435,N_1167,N_1372);
nor U3436 (N_3436,N_390,N_1947);
and U3437 (N_3437,N_716,N_2402);
and U3438 (N_3438,N_2189,N_1633);
or U3439 (N_3439,N_2464,N_2367);
and U3440 (N_3440,N_160,N_1093);
and U3441 (N_3441,N_900,N_1750);
nor U3442 (N_3442,N_1237,N_1593);
nand U3443 (N_3443,N_1131,N_1729);
nand U3444 (N_3444,N_280,N_2198);
nor U3445 (N_3445,N_314,N_886);
xnor U3446 (N_3446,N_1565,N_883);
nand U3447 (N_3447,N_1308,N_2039);
nand U3448 (N_3448,N_2456,N_787);
xor U3449 (N_3449,N_187,N_362);
nor U3450 (N_3450,N_1561,N_1826);
xnor U3451 (N_3451,N_507,N_1438);
nor U3452 (N_3452,N_1273,N_2480);
nor U3453 (N_3453,N_1998,N_551);
xnor U3454 (N_3454,N_1292,N_719);
and U3455 (N_3455,N_2437,N_174);
or U3456 (N_3456,N_887,N_860);
nand U3457 (N_3457,N_1444,N_906);
nor U3458 (N_3458,N_1489,N_69);
or U3459 (N_3459,N_2240,N_2254);
nand U3460 (N_3460,N_1643,N_587);
and U3461 (N_3461,N_423,N_552);
or U3462 (N_3462,N_37,N_190);
nor U3463 (N_3463,N_1641,N_676);
nand U3464 (N_3464,N_1269,N_1753);
and U3465 (N_3465,N_1979,N_1349);
and U3466 (N_3466,N_202,N_955);
and U3467 (N_3467,N_1719,N_94);
nor U3468 (N_3468,N_2115,N_1133);
nor U3469 (N_3469,N_2315,N_1279);
xnor U3470 (N_3470,N_1120,N_1098);
nor U3471 (N_3471,N_1126,N_1288);
nor U3472 (N_3472,N_1626,N_306);
and U3473 (N_3473,N_1236,N_357);
nor U3474 (N_3474,N_2170,N_2452);
xor U3475 (N_3475,N_1815,N_1566);
xor U3476 (N_3476,N_1253,N_523);
nor U3477 (N_3477,N_1879,N_1771);
or U3478 (N_3478,N_2259,N_1235);
or U3479 (N_3479,N_1852,N_380);
or U3480 (N_3480,N_292,N_1518);
and U3481 (N_3481,N_1502,N_2237);
nand U3482 (N_3482,N_1021,N_1175);
xor U3483 (N_3483,N_49,N_2109);
xnor U3484 (N_3484,N_393,N_872);
and U3485 (N_3485,N_725,N_547);
and U3486 (N_3486,N_1644,N_196);
nand U3487 (N_3487,N_1203,N_1730);
nand U3488 (N_3488,N_135,N_841);
and U3489 (N_3489,N_485,N_476);
nor U3490 (N_3490,N_1600,N_744);
nand U3491 (N_3491,N_244,N_937);
or U3492 (N_3492,N_1488,N_751);
xnor U3493 (N_3493,N_1106,N_2425);
and U3494 (N_3494,N_61,N_1859);
nor U3495 (N_3495,N_1073,N_1715);
or U3496 (N_3496,N_1590,N_1347);
or U3497 (N_3497,N_710,N_1430);
nand U3498 (N_3498,N_117,N_1409);
or U3499 (N_3499,N_2165,N_954);
nand U3500 (N_3500,N_1330,N_1576);
or U3501 (N_3501,N_347,N_1176);
xnor U3502 (N_3502,N_770,N_1725);
xor U3503 (N_3503,N_2073,N_2211);
nor U3504 (N_3504,N_661,N_2112);
or U3505 (N_3505,N_1843,N_1511);
and U3506 (N_3506,N_2467,N_1542);
nor U3507 (N_3507,N_1337,N_1100);
nand U3508 (N_3508,N_1968,N_748);
nand U3509 (N_3509,N_130,N_495);
nor U3510 (N_3510,N_1523,N_634);
nand U3511 (N_3511,N_1639,N_2415);
nor U3512 (N_3512,N_41,N_142);
nor U3513 (N_3513,N_733,N_2442);
or U3514 (N_3514,N_1731,N_1375);
nor U3515 (N_3515,N_29,N_927);
xnor U3516 (N_3516,N_726,N_2477);
nand U3517 (N_3517,N_1854,N_2380);
xor U3518 (N_3518,N_1651,N_2156);
nand U3519 (N_3519,N_284,N_1905);
nand U3520 (N_3520,N_921,N_1296);
and U3521 (N_3521,N_283,N_1204);
or U3522 (N_3522,N_1699,N_454);
or U3523 (N_3523,N_2444,N_1191);
xor U3524 (N_3524,N_157,N_1520);
or U3525 (N_3525,N_1801,N_2121);
nand U3526 (N_3526,N_377,N_2360);
or U3527 (N_3527,N_1703,N_39);
xor U3528 (N_3528,N_2028,N_368);
and U3529 (N_3529,N_1884,N_1187);
nand U3530 (N_3530,N_249,N_1892);
or U3531 (N_3531,N_1043,N_1513);
or U3532 (N_3532,N_123,N_463);
xnor U3533 (N_3533,N_2292,N_555);
and U3534 (N_3534,N_2489,N_1742);
nor U3535 (N_3535,N_1605,N_1556);
nor U3536 (N_3536,N_434,N_694);
xnor U3537 (N_3537,N_385,N_1239);
xnor U3538 (N_3538,N_2372,N_2177);
nand U3539 (N_3539,N_2376,N_995);
nand U3540 (N_3540,N_2289,N_1883);
or U3541 (N_3541,N_1426,N_1793);
nand U3542 (N_3542,N_95,N_2324);
nor U3543 (N_3543,N_441,N_16);
and U3544 (N_3544,N_2227,N_1493);
xor U3545 (N_3545,N_31,N_1770);
nor U3546 (N_3546,N_1967,N_2337);
or U3547 (N_3547,N_1802,N_301);
xor U3548 (N_3548,N_2190,N_337);
nor U3549 (N_3549,N_1265,N_544);
or U3550 (N_3550,N_1681,N_1040);
xor U3551 (N_3551,N_852,N_2276);
xnor U3552 (N_3552,N_93,N_484);
nand U3553 (N_3553,N_260,N_287);
nor U3554 (N_3554,N_1601,N_904);
or U3555 (N_3555,N_443,N_901);
xor U3556 (N_3556,N_1143,N_542);
or U3557 (N_3557,N_815,N_2230);
nand U3558 (N_3558,N_1180,N_221);
or U3559 (N_3559,N_389,N_2393);
xor U3560 (N_3560,N_1196,N_1972);
nor U3561 (N_3561,N_605,N_1909);
xnor U3562 (N_3562,N_1746,N_2350);
nand U3563 (N_3563,N_1836,N_1877);
or U3564 (N_3564,N_1168,N_431);
nand U3565 (N_3565,N_92,N_212);
nor U3566 (N_3566,N_1481,N_425);
or U3567 (N_3567,N_1707,N_2408);
or U3568 (N_3568,N_1378,N_2446);
and U3569 (N_3569,N_204,N_394);
and U3570 (N_3570,N_2029,N_757);
or U3571 (N_3571,N_219,N_1153);
nor U3572 (N_3572,N_74,N_985);
and U3573 (N_3573,N_2150,N_978);
and U3574 (N_3574,N_1329,N_467);
or U3575 (N_3575,N_839,N_972);
nor U3576 (N_3576,N_494,N_2468);
nor U3577 (N_3577,N_705,N_1275);
nor U3578 (N_3578,N_237,N_132);
and U3579 (N_3579,N_1463,N_167);
nor U3580 (N_3580,N_1769,N_1084);
nor U3581 (N_3581,N_1295,N_1595);
xnor U3582 (N_3582,N_2321,N_2200);
or U3583 (N_3583,N_1139,N_1509);
xor U3584 (N_3584,N_620,N_1439);
xor U3585 (N_3585,N_1037,N_517);
nand U3586 (N_3586,N_56,N_2406);
and U3587 (N_3587,N_354,N_1220);
or U3588 (N_3588,N_696,N_1454);
xnor U3589 (N_3589,N_509,N_1299);
xnor U3590 (N_3590,N_686,N_2453);
nand U3591 (N_3591,N_445,N_1351);
nand U3592 (N_3592,N_619,N_1418);
xor U3593 (N_3593,N_358,N_145);
nand U3594 (N_3594,N_2033,N_766);
and U3595 (N_3595,N_660,N_1957);
and U3596 (N_3596,N_837,N_461);
and U3597 (N_3597,N_793,N_1954);
xor U3598 (N_3598,N_761,N_54);
and U3599 (N_3599,N_756,N_1103);
xor U3600 (N_3600,N_666,N_1790);
and U3601 (N_3601,N_1104,N_785);
nor U3602 (N_3602,N_593,N_1480);
nor U3603 (N_3603,N_867,N_1991);
nor U3604 (N_3604,N_2299,N_2090);
nand U3605 (N_3605,N_1080,N_1169);
or U3606 (N_3606,N_163,N_1510);
xnor U3607 (N_3607,N_1931,N_742);
nor U3608 (N_3608,N_1551,N_1718);
xnor U3609 (N_3609,N_1971,N_2061);
and U3610 (N_3610,N_2114,N_920);
xor U3611 (N_3611,N_697,N_483);
nand U3612 (N_3612,N_1102,N_894);
nand U3613 (N_3613,N_323,N_2386);
or U3614 (N_3614,N_953,N_2335);
nor U3615 (N_3615,N_1266,N_1128);
nand U3616 (N_3616,N_1958,N_718);
xor U3617 (N_3617,N_1886,N_480);
nand U3618 (N_3618,N_63,N_2042);
and U3619 (N_3619,N_1634,N_104);
nand U3620 (N_3620,N_798,N_2137);
and U3621 (N_3621,N_1023,N_364);
and U3622 (N_3622,N_1436,N_1609);
or U3623 (N_3623,N_2293,N_1617);
or U3624 (N_3624,N_809,N_1076);
nand U3625 (N_3625,N_520,N_68);
and U3626 (N_3626,N_2336,N_1462);
nor U3627 (N_3627,N_861,N_1514);
and U3628 (N_3628,N_2423,N_1055);
nor U3629 (N_3629,N_1997,N_903);
nand U3630 (N_3630,N_1148,N_1923);
nor U3631 (N_3631,N_210,N_164);
nand U3632 (N_3632,N_1621,N_479);
nand U3633 (N_3633,N_1035,N_2391);
nor U3634 (N_3634,N_636,N_893);
nor U3635 (N_3635,N_491,N_1440);
nor U3636 (N_3636,N_205,N_1077);
nand U3637 (N_3637,N_1190,N_83);
nand U3638 (N_3638,N_1389,N_2291);
nor U3639 (N_3639,N_1558,N_1392);
nand U3640 (N_3640,N_1341,N_1832);
or U3641 (N_3641,N_2010,N_658);
or U3642 (N_3642,N_2223,N_1050);
nand U3643 (N_3643,N_1301,N_1060);
and U3644 (N_3644,N_801,N_315);
xnor U3645 (N_3645,N_1837,N_1492);
xor U3646 (N_3646,N_1786,N_805);
and U3647 (N_3647,N_1712,N_728);
nor U3648 (N_3648,N_2487,N_1828);
xor U3649 (N_3649,N_949,N_1662);
or U3650 (N_3650,N_1360,N_835);
or U3651 (N_3651,N_986,N_1682);
and U3652 (N_3652,N_1138,N_1654);
xnor U3653 (N_3653,N_214,N_2297);
and U3654 (N_3654,N_2126,N_539);
and U3655 (N_3655,N_1683,N_907);
nor U3656 (N_3656,N_1425,N_2076);
nand U3657 (N_3657,N_1677,N_1560);
and U3658 (N_3658,N_1734,N_1977);
xor U3659 (N_3659,N_684,N_420);
nand U3660 (N_3660,N_2488,N_1987);
nand U3661 (N_3661,N_1676,N_2258);
and U3662 (N_3662,N_2365,N_1895);
or U3663 (N_3663,N_6,N_648);
or U3664 (N_3664,N_241,N_2481);
and U3665 (N_3665,N_150,N_1992);
nor U3666 (N_3666,N_51,N_1158);
or U3667 (N_3667,N_2483,N_1591);
and U3668 (N_3668,N_1679,N_2108);
or U3669 (N_3669,N_371,N_657);
nand U3670 (N_3670,N_773,N_510);
or U3671 (N_3671,N_1581,N_884);
nand U3672 (N_3672,N_2311,N_398);
nor U3673 (N_3673,N_1343,N_1065);
nand U3674 (N_3674,N_2160,N_945);
or U3675 (N_3675,N_529,N_1281);
xor U3676 (N_3676,N_2460,N_2027);
and U3677 (N_3677,N_1951,N_1025);
or U3678 (N_3678,N_1996,N_384);
or U3679 (N_3679,N_282,N_1006);
or U3680 (N_3680,N_2248,N_1226);
and U3681 (N_3681,N_574,N_1395);
and U3682 (N_3682,N_1087,N_370);
nand U3683 (N_3683,N_1283,N_650);
and U3684 (N_3684,N_178,N_172);
and U3685 (N_3685,N_211,N_1307);
nor U3686 (N_3686,N_1170,N_1213);
and U3687 (N_3687,N_453,N_1524);
xor U3688 (N_3688,N_0,N_1615);
nand U3689 (N_3689,N_231,N_2328);
and U3690 (N_3690,N_947,N_307);
xor U3691 (N_3691,N_1497,N_1579);
nand U3692 (N_3692,N_367,N_1171);
or U3693 (N_3693,N_452,N_193);
nand U3694 (N_3694,N_179,N_107);
xnor U3695 (N_3695,N_2148,N_2234);
xor U3696 (N_3696,N_2412,N_1498);
nand U3697 (N_3697,N_369,N_2389);
xnor U3698 (N_3698,N_2267,N_566);
or U3699 (N_3699,N_1733,N_89);
and U3700 (N_3700,N_2298,N_225);
or U3701 (N_3701,N_1517,N_40);
nand U3702 (N_3702,N_2268,N_1500);
nand U3703 (N_3703,N_1116,N_1927);
nand U3704 (N_3704,N_1829,N_2093);
and U3705 (N_3705,N_738,N_1325);
or U3706 (N_3706,N_35,N_1726);
nor U3707 (N_3707,N_278,N_137);
or U3708 (N_3708,N_576,N_1665);
nor U3709 (N_3709,N_1868,N_2347);
or U3710 (N_3710,N_72,N_87);
or U3711 (N_3711,N_351,N_1530);
nand U3712 (N_3712,N_1989,N_376);
nand U3713 (N_3713,N_2184,N_843);
and U3714 (N_3714,N_1431,N_2038);
nor U3715 (N_3715,N_863,N_2096);
nor U3716 (N_3716,N_683,N_478);
xnor U3717 (N_3717,N_27,N_1908);
and U3718 (N_3718,N_355,N_806);
nand U3719 (N_3719,N_1066,N_1878);
or U3720 (N_3720,N_1960,N_1482);
and U3721 (N_3721,N_175,N_1675);
nand U3722 (N_3722,N_155,N_1506);
or U3723 (N_3723,N_1113,N_1539);
nor U3724 (N_3724,N_2066,N_2059);
or U3725 (N_3725,N_261,N_166);
xnor U3726 (N_3726,N_1696,N_629);
xor U3727 (N_3727,N_1041,N_1130);
nor U3728 (N_3728,N_401,N_1808);
nor U3729 (N_3729,N_414,N_1320);
nor U3730 (N_3730,N_2303,N_1907);
or U3731 (N_3731,N_1857,N_885);
nor U3732 (N_3732,N_2103,N_578);
nand U3733 (N_3733,N_1032,N_2144);
nor U3734 (N_3734,N_610,N_1254);
nand U3735 (N_3735,N_1435,N_965);
nor U3736 (N_3736,N_1413,N_492);
xnor U3737 (N_3737,N_1599,N_499);
nor U3738 (N_3738,N_745,N_2209);
and U3739 (N_3739,N_2100,N_2455);
nor U3740 (N_3740,N_866,N_1386);
or U3741 (N_3741,N_1460,N_1434);
nor U3742 (N_3742,N_2178,N_1570);
nor U3743 (N_3743,N_1748,N_2430);
nor U3744 (N_3744,N_1935,N_1385);
nand U3745 (N_3745,N_8,N_874);
xnor U3746 (N_3746,N_328,N_614);
and U3747 (N_3747,N_1792,N_1903);
nand U3748 (N_3748,N_1756,N_1962);
or U3749 (N_3749,N_522,N_1781);
nand U3750 (N_3750,N_1562,N_351);
nor U3751 (N_3751,N_614,N_2251);
and U3752 (N_3752,N_1746,N_749);
and U3753 (N_3753,N_1087,N_1716);
nand U3754 (N_3754,N_1960,N_2281);
nor U3755 (N_3755,N_1960,N_714);
nor U3756 (N_3756,N_1522,N_207);
nor U3757 (N_3757,N_760,N_1797);
xor U3758 (N_3758,N_737,N_1806);
nor U3759 (N_3759,N_508,N_1308);
nor U3760 (N_3760,N_253,N_1799);
and U3761 (N_3761,N_1040,N_194);
xor U3762 (N_3762,N_1612,N_418);
and U3763 (N_3763,N_2106,N_1220);
or U3764 (N_3764,N_2277,N_548);
nand U3765 (N_3765,N_1317,N_587);
nor U3766 (N_3766,N_21,N_656);
and U3767 (N_3767,N_1402,N_2140);
or U3768 (N_3768,N_1968,N_400);
nand U3769 (N_3769,N_2048,N_2391);
nor U3770 (N_3770,N_2184,N_1051);
nor U3771 (N_3771,N_1531,N_1163);
nand U3772 (N_3772,N_1436,N_1227);
xnor U3773 (N_3773,N_1177,N_1059);
nor U3774 (N_3774,N_1244,N_1397);
or U3775 (N_3775,N_1863,N_1394);
or U3776 (N_3776,N_1919,N_1201);
nand U3777 (N_3777,N_967,N_2215);
nand U3778 (N_3778,N_969,N_1556);
nor U3779 (N_3779,N_328,N_272);
nor U3780 (N_3780,N_445,N_500);
and U3781 (N_3781,N_2413,N_2399);
or U3782 (N_3782,N_1923,N_1843);
nand U3783 (N_3783,N_1882,N_525);
nand U3784 (N_3784,N_1921,N_721);
nand U3785 (N_3785,N_1438,N_111);
nand U3786 (N_3786,N_1237,N_2361);
or U3787 (N_3787,N_606,N_863);
nand U3788 (N_3788,N_105,N_657);
or U3789 (N_3789,N_836,N_949);
nor U3790 (N_3790,N_894,N_2487);
or U3791 (N_3791,N_185,N_2131);
and U3792 (N_3792,N_691,N_2253);
xnor U3793 (N_3793,N_1493,N_746);
nor U3794 (N_3794,N_378,N_299);
and U3795 (N_3795,N_2070,N_2420);
or U3796 (N_3796,N_187,N_2283);
or U3797 (N_3797,N_48,N_2318);
or U3798 (N_3798,N_1571,N_2461);
and U3799 (N_3799,N_1237,N_1242);
xor U3800 (N_3800,N_1625,N_1103);
and U3801 (N_3801,N_832,N_2423);
or U3802 (N_3802,N_730,N_1946);
nor U3803 (N_3803,N_1129,N_2473);
and U3804 (N_3804,N_2356,N_787);
nor U3805 (N_3805,N_83,N_542);
or U3806 (N_3806,N_694,N_937);
nor U3807 (N_3807,N_1088,N_172);
nand U3808 (N_3808,N_712,N_1189);
nor U3809 (N_3809,N_534,N_1045);
nor U3810 (N_3810,N_30,N_2158);
nand U3811 (N_3811,N_1793,N_1333);
nand U3812 (N_3812,N_2467,N_577);
nor U3813 (N_3813,N_1002,N_43);
or U3814 (N_3814,N_1531,N_1836);
or U3815 (N_3815,N_1195,N_1208);
nor U3816 (N_3816,N_20,N_1741);
or U3817 (N_3817,N_1140,N_1976);
or U3818 (N_3818,N_647,N_424);
nand U3819 (N_3819,N_1260,N_2293);
xor U3820 (N_3820,N_2255,N_925);
nor U3821 (N_3821,N_458,N_2494);
xnor U3822 (N_3822,N_1014,N_179);
xor U3823 (N_3823,N_1198,N_2188);
nor U3824 (N_3824,N_1984,N_1451);
xnor U3825 (N_3825,N_2017,N_1587);
nand U3826 (N_3826,N_1004,N_2391);
xor U3827 (N_3827,N_2237,N_1231);
or U3828 (N_3828,N_1765,N_793);
or U3829 (N_3829,N_943,N_1213);
or U3830 (N_3830,N_1170,N_1712);
xnor U3831 (N_3831,N_1285,N_974);
nor U3832 (N_3832,N_1581,N_660);
and U3833 (N_3833,N_2084,N_1757);
xor U3834 (N_3834,N_2142,N_350);
and U3835 (N_3835,N_699,N_1140);
nor U3836 (N_3836,N_2009,N_1077);
nand U3837 (N_3837,N_134,N_465);
nand U3838 (N_3838,N_907,N_688);
and U3839 (N_3839,N_917,N_978);
nand U3840 (N_3840,N_1090,N_1916);
or U3841 (N_3841,N_2054,N_1957);
xnor U3842 (N_3842,N_1208,N_1422);
nor U3843 (N_3843,N_937,N_1300);
nor U3844 (N_3844,N_142,N_901);
xor U3845 (N_3845,N_2383,N_1321);
xnor U3846 (N_3846,N_1418,N_1351);
xor U3847 (N_3847,N_1290,N_2094);
or U3848 (N_3848,N_796,N_1224);
nor U3849 (N_3849,N_1385,N_2126);
nor U3850 (N_3850,N_2285,N_144);
xnor U3851 (N_3851,N_653,N_302);
or U3852 (N_3852,N_2068,N_1417);
and U3853 (N_3853,N_483,N_1070);
nand U3854 (N_3854,N_1799,N_957);
or U3855 (N_3855,N_677,N_1214);
xnor U3856 (N_3856,N_580,N_1448);
and U3857 (N_3857,N_340,N_1670);
xor U3858 (N_3858,N_338,N_658);
nor U3859 (N_3859,N_1081,N_2173);
nand U3860 (N_3860,N_1080,N_1417);
nand U3861 (N_3861,N_2,N_1772);
or U3862 (N_3862,N_2106,N_1567);
or U3863 (N_3863,N_860,N_2255);
nor U3864 (N_3864,N_413,N_282);
or U3865 (N_3865,N_459,N_199);
and U3866 (N_3866,N_124,N_2477);
and U3867 (N_3867,N_1563,N_610);
nor U3868 (N_3868,N_1346,N_1792);
or U3869 (N_3869,N_233,N_1062);
or U3870 (N_3870,N_1677,N_2031);
or U3871 (N_3871,N_2288,N_13);
xor U3872 (N_3872,N_26,N_1668);
xnor U3873 (N_3873,N_1434,N_1405);
xnor U3874 (N_3874,N_776,N_726);
and U3875 (N_3875,N_1847,N_1172);
or U3876 (N_3876,N_2149,N_468);
and U3877 (N_3877,N_550,N_770);
and U3878 (N_3878,N_721,N_1122);
and U3879 (N_3879,N_1999,N_1402);
or U3880 (N_3880,N_46,N_1889);
nor U3881 (N_3881,N_154,N_1703);
xor U3882 (N_3882,N_464,N_427);
and U3883 (N_3883,N_550,N_1734);
xor U3884 (N_3884,N_1680,N_1898);
nand U3885 (N_3885,N_1369,N_1298);
and U3886 (N_3886,N_400,N_2453);
nor U3887 (N_3887,N_1315,N_715);
and U3888 (N_3888,N_1580,N_1566);
and U3889 (N_3889,N_2452,N_1177);
and U3890 (N_3890,N_2019,N_2316);
and U3891 (N_3891,N_666,N_1946);
or U3892 (N_3892,N_1232,N_456);
nand U3893 (N_3893,N_1155,N_2352);
and U3894 (N_3894,N_2176,N_1869);
or U3895 (N_3895,N_994,N_1989);
xnor U3896 (N_3896,N_1550,N_1707);
xor U3897 (N_3897,N_1934,N_1239);
nor U3898 (N_3898,N_162,N_2221);
nor U3899 (N_3899,N_1280,N_898);
xnor U3900 (N_3900,N_1358,N_246);
and U3901 (N_3901,N_1211,N_2211);
nand U3902 (N_3902,N_190,N_1194);
and U3903 (N_3903,N_1401,N_1577);
or U3904 (N_3904,N_549,N_503);
xnor U3905 (N_3905,N_2391,N_449);
or U3906 (N_3906,N_1069,N_2214);
or U3907 (N_3907,N_1670,N_1364);
nor U3908 (N_3908,N_2062,N_635);
xor U3909 (N_3909,N_2033,N_580);
nor U3910 (N_3910,N_2082,N_311);
xor U3911 (N_3911,N_357,N_560);
or U3912 (N_3912,N_2147,N_1350);
nor U3913 (N_3913,N_1475,N_1508);
nor U3914 (N_3914,N_1478,N_855);
xnor U3915 (N_3915,N_890,N_1564);
and U3916 (N_3916,N_2351,N_1521);
xnor U3917 (N_3917,N_2380,N_60);
nor U3918 (N_3918,N_1979,N_2037);
and U3919 (N_3919,N_1578,N_2024);
and U3920 (N_3920,N_120,N_239);
xor U3921 (N_3921,N_486,N_2416);
xor U3922 (N_3922,N_114,N_2426);
nor U3923 (N_3923,N_1804,N_819);
or U3924 (N_3924,N_1030,N_2017);
and U3925 (N_3925,N_725,N_1449);
nor U3926 (N_3926,N_430,N_2294);
nand U3927 (N_3927,N_1703,N_51);
nor U3928 (N_3928,N_1364,N_1190);
or U3929 (N_3929,N_1935,N_1723);
or U3930 (N_3930,N_1331,N_2093);
nor U3931 (N_3931,N_63,N_367);
xor U3932 (N_3932,N_600,N_1968);
nand U3933 (N_3933,N_1013,N_503);
nor U3934 (N_3934,N_1334,N_2461);
xnor U3935 (N_3935,N_1340,N_816);
nor U3936 (N_3936,N_866,N_65);
or U3937 (N_3937,N_707,N_881);
or U3938 (N_3938,N_1488,N_353);
or U3939 (N_3939,N_2250,N_2147);
and U3940 (N_3940,N_1762,N_1949);
nand U3941 (N_3941,N_1307,N_1203);
xor U3942 (N_3942,N_363,N_988);
nor U3943 (N_3943,N_844,N_2492);
or U3944 (N_3944,N_2211,N_1396);
nand U3945 (N_3945,N_2251,N_2483);
nor U3946 (N_3946,N_465,N_765);
and U3947 (N_3947,N_2275,N_1953);
and U3948 (N_3948,N_657,N_969);
or U3949 (N_3949,N_825,N_63);
nand U3950 (N_3950,N_1534,N_2192);
or U3951 (N_3951,N_1796,N_740);
nor U3952 (N_3952,N_2286,N_1919);
nor U3953 (N_3953,N_16,N_1965);
nand U3954 (N_3954,N_1798,N_1428);
nor U3955 (N_3955,N_833,N_2421);
nor U3956 (N_3956,N_1301,N_889);
xor U3957 (N_3957,N_2037,N_2401);
or U3958 (N_3958,N_1163,N_1793);
or U3959 (N_3959,N_2213,N_938);
nor U3960 (N_3960,N_896,N_2111);
nand U3961 (N_3961,N_454,N_153);
nor U3962 (N_3962,N_2269,N_207);
and U3963 (N_3963,N_1546,N_1854);
nor U3964 (N_3964,N_236,N_1158);
nor U3965 (N_3965,N_432,N_1629);
and U3966 (N_3966,N_740,N_615);
and U3967 (N_3967,N_603,N_2480);
nor U3968 (N_3968,N_1412,N_910);
nor U3969 (N_3969,N_1194,N_1722);
nand U3970 (N_3970,N_1670,N_514);
nor U3971 (N_3971,N_1827,N_824);
nand U3972 (N_3972,N_445,N_851);
nor U3973 (N_3973,N_2275,N_259);
nand U3974 (N_3974,N_2418,N_1466);
xnor U3975 (N_3975,N_1549,N_2320);
nand U3976 (N_3976,N_62,N_2456);
nand U3977 (N_3977,N_1740,N_818);
and U3978 (N_3978,N_2107,N_1282);
and U3979 (N_3979,N_787,N_676);
xor U3980 (N_3980,N_2450,N_1954);
and U3981 (N_3981,N_10,N_2280);
xnor U3982 (N_3982,N_2127,N_1355);
nand U3983 (N_3983,N_850,N_2447);
xnor U3984 (N_3984,N_417,N_159);
nand U3985 (N_3985,N_418,N_334);
or U3986 (N_3986,N_2072,N_882);
nand U3987 (N_3987,N_178,N_1939);
nor U3988 (N_3988,N_1423,N_421);
or U3989 (N_3989,N_1970,N_1606);
nand U3990 (N_3990,N_1644,N_1095);
or U3991 (N_3991,N_2242,N_285);
and U3992 (N_3992,N_2125,N_1482);
or U3993 (N_3993,N_320,N_2011);
nand U3994 (N_3994,N_1252,N_649);
nor U3995 (N_3995,N_1142,N_2048);
and U3996 (N_3996,N_1066,N_964);
and U3997 (N_3997,N_2032,N_1114);
nand U3998 (N_3998,N_603,N_625);
xor U3999 (N_3999,N_2189,N_2030);
and U4000 (N_4000,N_1051,N_374);
nand U4001 (N_4001,N_2077,N_1991);
and U4002 (N_4002,N_405,N_499);
nand U4003 (N_4003,N_1503,N_1817);
xor U4004 (N_4004,N_2179,N_1682);
nand U4005 (N_4005,N_2255,N_1068);
nor U4006 (N_4006,N_943,N_30);
or U4007 (N_4007,N_959,N_2124);
nor U4008 (N_4008,N_335,N_2475);
nor U4009 (N_4009,N_2173,N_1232);
nor U4010 (N_4010,N_1533,N_1993);
nor U4011 (N_4011,N_1270,N_2275);
or U4012 (N_4012,N_260,N_1971);
nor U4013 (N_4013,N_2124,N_1689);
and U4014 (N_4014,N_16,N_1174);
xor U4015 (N_4015,N_2356,N_551);
and U4016 (N_4016,N_1663,N_817);
or U4017 (N_4017,N_2098,N_1714);
nor U4018 (N_4018,N_2407,N_147);
xnor U4019 (N_4019,N_756,N_1316);
and U4020 (N_4020,N_1801,N_1624);
nor U4021 (N_4021,N_49,N_1271);
or U4022 (N_4022,N_394,N_2369);
and U4023 (N_4023,N_742,N_1646);
and U4024 (N_4024,N_1086,N_2112);
or U4025 (N_4025,N_1207,N_337);
nor U4026 (N_4026,N_1881,N_1563);
or U4027 (N_4027,N_1482,N_2383);
xor U4028 (N_4028,N_1278,N_1724);
and U4029 (N_4029,N_139,N_748);
nand U4030 (N_4030,N_861,N_364);
nand U4031 (N_4031,N_1926,N_15);
nor U4032 (N_4032,N_1581,N_815);
or U4033 (N_4033,N_2250,N_706);
nor U4034 (N_4034,N_40,N_1853);
xor U4035 (N_4035,N_1251,N_499);
nand U4036 (N_4036,N_987,N_2001);
or U4037 (N_4037,N_1258,N_1860);
nand U4038 (N_4038,N_544,N_1579);
nand U4039 (N_4039,N_326,N_1289);
nor U4040 (N_4040,N_100,N_2180);
nand U4041 (N_4041,N_2391,N_1419);
xnor U4042 (N_4042,N_1078,N_2267);
nand U4043 (N_4043,N_209,N_1996);
or U4044 (N_4044,N_2348,N_1638);
nand U4045 (N_4045,N_1851,N_877);
nor U4046 (N_4046,N_1911,N_2396);
nand U4047 (N_4047,N_1506,N_2272);
nand U4048 (N_4048,N_265,N_1777);
or U4049 (N_4049,N_32,N_806);
nor U4050 (N_4050,N_337,N_375);
xor U4051 (N_4051,N_2235,N_2444);
xor U4052 (N_4052,N_665,N_330);
xor U4053 (N_4053,N_749,N_1127);
and U4054 (N_4054,N_2383,N_1593);
nand U4055 (N_4055,N_133,N_669);
xnor U4056 (N_4056,N_1058,N_2048);
nand U4057 (N_4057,N_2122,N_709);
nor U4058 (N_4058,N_800,N_2135);
xor U4059 (N_4059,N_1420,N_2448);
nand U4060 (N_4060,N_628,N_1097);
nor U4061 (N_4061,N_1976,N_2114);
or U4062 (N_4062,N_1736,N_1020);
nand U4063 (N_4063,N_60,N_2155);
and U4064 (N_4064,N_637,N_1469);
nor U4065 (N_4065,N_991,N_354);
nand U4066 (N_4066,N_1611,N_971);
nand U4067 (N_4067,N_2226,N_498);
and U4068 (N_4068,N_1238,N_1844);
and U4069 (N_4069,N_859,N_1118);
nand U4070 (N_4070,N_1150,N_648);
or U4071 (N_4071,N_2283,N_363);
xnor U4072 (N_4072,N_712,N_880);
nand U4073 (N_4073,N_322,N_1665);
xor U4074 (N_4074,N_232,N_2088);
or U4075 (N_4075,N_1758,N_202);
nand U4076 (N_4076,N_399,N_456);
nor U4077 (N_4077,N_2274,N_694);
or U4078 (N_4078,N_2267,N_473);
nand U4079 (N_4079,N_221,N_326);
nor U4080 (N_4080,N_1448,N_133);
or U4081 (N_4081,N_391,N_2491);
and U4082 (N_4082,N_913,N_1239);
or U4083 (N_4083,N_306,N_286);
nand U4084 (N_4084,N_992,N_716);
xor U4085 (N_4085,N_2295,N_345);
xnor U4086 (N_4086,N_1088,N_2423);
and U4087 (N_4087,N_1838,N_1122);
or U4088 (N_4088,N_574,N_49);
or U4089 (N_4089,N_1233,N_2030);
xnor U4090 (N_4090,N_2230,N_2462);
nor U4091 (N_4091,N_2228,N_604);
xnor U4092 (N_4092,N_1845,N_150);
xor U4093 (N_4093,N_1756,N_589);
xnor U4094 (N_4094,N_2126,N_1065);
xor U4095 (N_4095,N_2104,N_400);
and U4096 (N_4096,N_972,N_462);
nor U4097 (N_4097,N_1893,N_2188);
and U4098 (N_4098,N_968,N_1487);
or U4099 (N_4099,N_934,N_1349);
and U4100 (N_4100,N_515,N_331);
nor U4101 (N_4101,N_2190,N_1692);
or U4102 (N_4102,N_1844,N_1768);
xor U4103 (N_4103,N_716,N_1104);
xnor U4104 (N_4104,N_1208,N_532);
xor U4105 (N_4105,N_1002,N_477);
and U4106 (N_4106,N_1898,N_360);
and U4107 (N_4107,N_67,N_1377);
xnor U4108 (N_4108,N_2116,N_37);
xor U4109 (N_4109,N_1086,N_450);
xor U4110 (N_4110,N_2271,N_866);
xnor U4111 (N_4111,N_1589,N_968);
nor U4112 (N_4112,N_868,N_1423);
xnor U4113 (N_4113,N_516,N_1208);
nor U4114 (N_4114,N_180,N_1527);
nand U4115 (N_4115,N_1744,N_669);
and U4116 (N_4116,N_1111,N_135);
nor U4117 (N_4117,N_1082,N_698);
nand U4118 (N_4118,N_140,N_1160);
nand U4119 (N_4119,N_896,N_331);
xnor U4120 (N_4120,N_823,N_795);
nand U4121 (N_4121,N_213,N_2014);
or U4122 (N_4122,N_809,N_2341);
and U4123 (N_4123,N_974,N_1226);
xor U4124 (N_4124,N_773,N_992);
nor U4125 (N_4125,N_333,N_2441);
nand U4126 (N_4126,N_2361,N_333);
and U4127 (N_4127,N_211,N_2361);
nand U4128 (N_4128,N_977,N_2167);
and U4129 (N_4129,N_2144,N_207);
nor U4130 (N_4130,N_1309,N_86);
and U4131 (N_4131,N_452,N_722);
xnor U4132 (N_4132,N_414,N_1411);
or U4133 (N_4133,N_1272,N_29);
nand U4134 (N_4134,N_2125,N_392);
and U4135 (N_4135,N_2491,N_404);
nand U4136 (N_4136,N_955,N_1192);
or U4137 (N_4137,N_1669,N_277);
and U4138 (N_4138,N_1357,N_1101);
and U4139 (N_4139,N_751,N_959);
nand U4140 (N_4140,N_1732,N_81);
or U4141 (N_4141,N_1777,N_1302);
and U4142 (N_4142,N_2139,N_1123);
xor U4143 (N_4143,N_112,N_1290);
or U4144 (N_4144,N_1117,N_149);
xor U4145 (N_4145,N_708,N_364);
or U4146 (N_4146,N_13,N_1765);
nand U4147 (N_4147,N_2180,N_2420);
or U4148 (N_4148,N_43,N_1115);
xnor U4149 (N_4149,N_2151,N_418);
and U4150 (N_4150,N_980,N_740);
nand U4151 (N_4151,N_3,N_1978);
nand U4152 (N_4152,N_1740,N_746);
nor U4153 (N_4153,N_2390,N_2251);
xnor U4154 (N_4154,N_150,N_2372);
or U4155 (N_4155,N_783,N_1738);
nor U4156 (N_4156,N_1608,N_348);
or U4157 (N_4157,N_543,N_1405);
nor U4158 (N_4158,N_2076,N_1017);
xor U4159 (N_4159,N_1485,N_1914);
or U4160 (N_4160,N_2219,N_1998);
nand U4161 (N_4161,N_2252,N_1472);
nor U4162 (N_4162,N_903,N_703);
nor U4163 (N_4163,N_2283,N_2097);
nand U4164 (N_4164,N_1343,N_274);
nor U4165 (N_4165,N_1186,N_396);
xor U4166 (N_4166,N_26,N_235);
or U4167 (N_4167,N_1553,N_2274);
nand U4168 (N_4168,N_760,N_700);
nor U4169 (N_4169,N_591,N_1537);
and U4170 (N_4170,N_1002,N_2185);
or U4171 (N_4171,N_1961,N_925);
xor U4172 (N_4172,N_1743,N_725);
and U4173 (N_4173,N_1902,N_1270);
or U4174 (N_4174,N_1933,N_1800);
nor U4175 (N_4175,N_1034,N_1131);
or U4176 (N_4176,N_107,N_1059);
xor U4177 (N_4177,N_934,N_593);
nand U4178 (N_4178,N_842,N_477);
nand U4179 (N_4179,N_2132,N_358);
or U4180 (N_4180,N_409,N_2045);
xnor U4181 (N_4181,N_2479,N_683);
nand U4182 (N_4182,N_323,N_1528);
and U4183 (N_4183,N_1366,N_1956);
or U4184 (N_4184,N_1887,N_2313);
or U4185 (N_4185,N_1376,N_1888);
nor U4186 (N_4186,N_1243,N_300);
nor U4187 (N_4187,N_1178,N_2247);
nor U4188 (N_4188,N_2087,N_1764);
xnor U4189 (N_4189,N_619,N_1662);
xor U4190 (N_4190,N_1838,N_2299);
and U4191 (N_4191,N_1702,N_800);
and U4192 (N_4192,N_2101,N_2478);
xnor U4193 (N_4193,N_2159,N_2002);
and U4194 (N_4194,N_780,N_404);
or U4195 (N_4195,N_79,N_1880);
and U4196 (N_4196,N_434,N_898);
and U4197 (N_4197,N_674,N_1545);
nand U4198 (N_4198,N_2444,N_1545);
or U4199 (N_4199,N_2022,N_235);
nand U4200 (N_4200,N_1576,N_1239);
nand U4201 (N_4201,N_294,N_1881);
nand U4202 (N_4202,N_159,N_1041);
and U4203 (N_4203,N_1341,N_1306);
and U4204 (N_4204,N_1141,N_251);
xnor U4205 (N_4205,N_762,N_699);
or U4206 (N_4206,N_1194,N_1197);
and U4207 (N_4207,N_202,N_2306);
nand U4208 (N_4208,N_1743,N_671);
or U4209 (N_4209,N_1182,N_981);
xnor U4210 (N_4210,N_646,N_1713);
and U4211 (N_4211,N_912,N_2350);
nand U4212 (N_4212,N_282,N_538);
nor U4213 (N_4213,N_1908,N_302);
nor U4214 (N_4214,N_447,N_1046);
xnor U4215 (N_4215,N_1994,N_1972);
or U4216 (N_4216,N_1487,N_206);
xnor U4217 (N_4217,N_580,N_2190);
nand U4218 (N_4218,N_2157,N_1027);
nand U4219 (N_4219,N_21,N_180);
or U4220 (N_4220,N_2476,N_2081);
nor U4221 (N_4221,N_1155,N_1463);
nand U4222 (N_4222,N_599,N_1784);
nor U4223 (N_4223,N_455,N_1441);
and U4224 (N_4224,N_643,N_1333);
and U4225 (N_4225,N_52,N_1753);
nand U4226 (N_4226,N_660,N_2076);
and U4227 (N_4227,N_178,N_2442);
or U4228 (N_4228,N_1886,N_1747);
nor U4229 (N_4229,N_2413,N_2118);
and U4230 (N_4230,N_2301,N_1947);
or U4231 (N_4231,N_1449,N_1990);
nand U4232 (N_4232,N_1522,N_1737);
xor U4233 (N_4233,N_2064,N_817);
nand U4234 (N_4234,N_821,N_1630);
or U4235 (N_4235,N_565,N_2096);
nand U4236 (N_4236,N_179,N_3);
or U4237 (N_4237,N_2393,N_2291);
nor U4238 (N_4238,N_1923,N_447);
nor U4239 (N_4239,N_2100,N_501);
xnor U4240 (N_4240,N_88,N_1782);
and U4241 (N_4241,N_594,N_850);
or U4242 (N_4242,N_67,N_1594);
nand U4243 (N_4243,N_634,N_713);
xor U4244 (N_4244,N_1769,N_2330);
nand U4245 (N_4245,N_1318,N_964);
or U4246 (N_4246,N_1744,N_847);
nor U4247 (N_4247,N_1408,N_1765);
or U4248 (N_4248,N_2238,N_2332);
or U4249 (N_4249,N_794,N_984);
nor U4250 (N_4250,N_1617,N_1968);
and U4251 (N_4251,N_1664,N_2465);
or U4252 (N_4252,N_2347,N_904);
nor U4253 (N_4253,N_2145,N_2085);
and U4254 (N_4254,N_1127,N_2065);
or U4255 (N_4255,N_2403,N_1250);
or U4256 (N_4256,N_1254,N_2278);
xor U4257 (N_4257,N_2119,N_1929);
or U4258 (N_4258,N_2449,N_369);
nor U4259 (N_4259,N_1370,N_1761);
xor U4260 (N_4260,N_1242,N_944);
or U4261 (N_4261,N_723,N_1163);
or U4262 (N_4262,N_2221,N_656);
nand U4263 (N_4263,N_471,N_141);
nor U4264 (N_4264,N_1428,N_1735);
xnor U4265 (N_4265,N_262,N_2033);
and U4266 (N_4266,N_1922,N_2456);
nor U4267 (N_4267,N_1693,N_378);
nand U4268 (N_4268,N_249,N_1645);
xnor U4269 (N_4269,N_1158,N_2244);
or U4270 (N_4270,N_1249,N_1678);
nand U4271 (N_4271,N_2097,N_2129);
xor U4272 (N_4272,N_690,N_325);
and U4273 (N_4273,N_1472,N_1832);
and U4274 (N_4274,N_506,N_1451);
nor U4275 (N_4275,N_1856,N_1891);
xnor U4276 (N_4276,N_1993,N_541);
nor U4277 (N_4277,N_1547,N_1895);
xnor U4278 (N_4278,N_981,N_881);
nor U4279 (N_4279,N_1953,N_341);
xor U4280 (N_4280,N_1330,N_1425);
nor U4281 (N_4281,N_1449,N_1607);
and U4282 (N_4282,N_477,N_16);
and U4283 (N_4283,N_920,N_1495);
or U4284 (N_4284,N_1200,N_756);
and U4285 (N_4285,N_1379,N_2184);
nand U4286 (N_4286,N_1698,N_1822);
nor U4287 (N_4287,N_711,N_1461);
xnor U4288 (N_4288,N_2317,N_1504);
xnor U4289 (N_4289,N_218,N_1807);
nand U4290 (N_4290,N_1387,N_1605);
nand U4291 (N_4291,N_115,N_1162);
or U4292 (N_4292,N_328,N_1249);
xor U4293 (N_4293,N_1511,N_1088);
nor U4294 (N_4294,N_1115,N_1450);
nand U4295 (N_4295,N_1863,N_1299);
and U4296 (N_4296,N_1615,N_1138);
nor U4297 (N_4297,N_721,N_1520);
or U4298 (N_4298,N_1535,N_1825);
nand U4299 (N_4299,N_1006,N_403);
and U4300 (N_4300,N_1258,N_2209);
xor U4301 (N_4301,N_804,N_675);
and U4302 (N_4302,N_2385,N_939);
or U4303 (N_4303,N_536,N_140);
nor U4304 (N_4304,N_967,N_1825);
and U4305 (N_4305,N_1338,N_119);
nand U4306 (N_4306,N_2460,N_747);
nor U4307 (N_4307,N_2261,N_1900);
and U4308 (N_4308,N_1539,N_1750);
xor U4309 (N_4309,N_698,N_496);
nand U4310 (N_4310,N_2325,N_2142);
nor U4311 (N_4311,N_2205,N_1761);
xor U4312 (N_4312,N_222,N_528);
xor U4313 (N_4313,N_1045,N_494);
xor U4314 (N_4314,N_530,N_679);
nor U4315 (N_4315,N_561,N_1463);
or U4316 (N_4316,N_135,N_1075);
nand U4317 (N_4317,N_1663,N_709);
xor U4318 (N_4318,N_418,N_1383);
nand U4319 (N_4319,N_477,N_469);
nor U4320 (N_4320,N_1099,N_1274);
and U4321 (N_4321,N_141,N_843);
and U4322 (N_4322,N_2364,N_759);
nor U4323 (N_4323,N_337,N_786);
and U4324 (N_4324,N_629,N_418);
xor U4325 (N_4325,N_66,N_2238);
nand U4326 (N_4326,N_2270,N_1822);
and U4327 (N_4327,N_35,N_667);
nand U4328 (N_4328,N_2239,N_128);
nor U4329 (N_4329,N_1180,N_414);
nand U4330 (N_4330,N_763,N_1241);
or U4331 (N_4331,N_424,N_1147);
and U4332 (N_4332,N_2151,N_789);
nor U4333 (N_4333,N_895,N_796);
nor U4334 (N_4334,N_93,N_1078);
nor U4335 (N_4335,N_2058,N_1480);
nand U4336 (N_4336,N_1875,N_1365);
xnor U4337 (N_4337,N_1027,N_578);
nand U4338 (N_4338,N_2056,N_1495);
or U4339 (N_4339,N_1213,N_345);
nor U4340 (N_4340,N_509,N_330);
xor U4341 (N_4341,N_1431,N_2431);
or U4342 (N_4342,N_374,N_2276);
and U4343 (N_4343,N_1031,N_1070);
or U4344 (N_4344,N_85,N_1067);
nor U4345 (N_4345,N_500,N_1215);
or U4346 (N_4346,N_1613,N_1760);
and U4347 (N_4347,N_1012,N_868);
and U4348 (N_4348,N_1311,N_883);
and U4349 (N_4349,N_828,N_60);
and U4350 (N_4350,N_893,N_1762);
nor U4351 (N_4351,N_310,N_2361);
nand U4352 (N_4352,N_2091,N_441);
or U4353 (N_4353,N_1624,N_159);
xor U4354 (N_4354,N_347,N_931);
or U4355 (N_4355,N_1443,N_2237);
or U4356 (N_4356,N_1056,N_1017);
nor U4357 (N_4357,N_1634,N_483);
xor U4358 (N_4358,N_1871,N_304);
xor U4359 (N_4359,N_1239,N_893);
nand U4360 (N_4360,N_48,N_251);
or U4361 (N_4361,N_2045,N_1383);
nor U4362 (N_4362,N_504,N_1451);
nor U4363 (N_4363,N_1206,N_2138);
nand U4364 (N_4364,N_429,N_1788);
and U4365 (N_4365,N_221,N_1217);
nand U4366 (N_4366,N_1091,N_1106);
or U4367 (N_4367,N_116,N_1893);
nand U4368 (N_4368,N_1265,N_622);
or U4369 (N_4369,N_286,N_2338);
and U4370 (N_4370,N_1830,N_1423);
and U4371 (N_4371,N_420,N_1917);
xor U4372 (N_4372,N_808,N_1414);
nor U4373 (N_4373,N_1619,N_459);
or U4374 (N_4374,N_1754,N_1318);
nand U4375 (N_4375,N_1712,N_271);
nor U4376 (N_4376,N_901,N_624);
xnor U4377 (N_4377,N_1029,N_357);
nor U4378 (N_4378,N_235,N_1880);
and U4379 (N_4379,N_549,N_1234);
and U4380 (N_4380,N_2181,N_1822);
nand U4381 (N_4381,N_1534,N_1761);
nor U4382 (N_4382,N_82,N_884);
xor U4383 (N_4383,N_1753,N_712);
or U4384 (N_4384,N_1843,N_1131);
nand U4385 (N_4385,N_1188,N_2193);
nor U4386 (N_4386,N_683,N_355);
nor U4387 (N_4387,N_472,N_755);
and U4388 (N_4388,N_745,N_1472);
or U4389 (N_4389,N_178,N_1595);
and U4390 (N_4390,N_1618,N_2241);
nand U4391 (N_4391,N_1506,N_2339);
nor U4392 (N_4392,N_832,N_2193);
or U4393 (N_4393,N_818,N_1028);
xor U4394 (N_4394,N_1619,N_1037);
and U4395 (N_4395,N_873,N_1970);
or U4396 (N_4396,N_502,N_1802);
nor U4397 (N_4397,N_189,N_2414);
nor U4398 (N_4398,N_2378,N_1353);
and U4399 (N_4399,N_384,N_370);
or U4400 (N_4400,N_1740,N_794);
and U4401 (N_4401,N_548,N_1410);
nand U4402 (N_4402,N_430,N_1573);
xnor U4403 (N_4403,N_2415,N_2177);
nand U4404 (N_4404,N_237,N_1630);
nand U4405 (N_4405,N_1204,N_2004);
nand U4406 (N_4406,N_1465,N_2454);
and U4407 (N_4407,N_1735,N_2254);
nor U4408 (N_4408,N_1756,N_1475);
or U4409 (N_4409,N_1032,N_795);
nor U4410 (N_4410,N_1260,N_1457);
and U4411 (N_4411,N_118,N_1694);
nor U4412 (N_4412,N_993,N_104);
nor U4413 (N_4413,N_1094,N_2414);
xnor U4414 (N_4414,N_661,N_1938);
nor U4415 (N_4415,N_1170,N_2151);
or U4416 (N_4416,N_1622,N_70);
or U4417 (N_4417,N_2264,N_1733);
and U4418 (N_4418,N_1743,N_155);
or U4419 (N_4419,N_505,N_638);
xor U4420 (N_4420,N_2334,N_1063);
or U4421 (N_4421,N_1561,N_2283);
and U4422 (N_4422,N_2020,N_503);
or U4423 (N_4423,N_496,N_2042);
nor U4424 (N_4424,N_502,N_1991);
nand U4425 (N_4425,N_1100,N_1186);
xnor U4426 (N_4426,N_2233,N_756);
nand U4427 (N_4427,N_554,N_1233);
nand U4428 (N_4428,N_580,N_244);
or U4429 (N_4429,N_662,N_2206);
nand U4430 (N_4430,N_155,N_87);
nand U4431 (N_4431,N_808,N_1773);
and U4432 (N_4432,N_2354,N_651);
xnor U4433 (N_4433,N_2358,N_1003);
or U4434 (N_4434,N_2062,N_1991);
or U4435 (N_4435,N_1322,N_108);
nor U4436 (N_4436,N_1657,N_1830);
nand U4437 (N_4437,N_1876,N_1586);
and U4438 (N_4438,N_654,N_2219);
or U4439 (N_4439,N_1439,N_551);
nand U4440 (N_4440,N_1331,N_18);
xnor U4441 (N_4441,N_2329,N_1657);
nand U4442 (N_4442,N_1203,N_1163);
nand U4443 (N_4443,N_146,N_1005);
nand U4444 (N_4444,N_1901,N_1856);
nor U4445 (N_4445,N_1971,N_2320);
or U4446 (N_4446,N_1732,N_364);
or U4447 (N_4447,N_236,N_1951);
nor U4448 (N_4448,N_172,N_2473);
nand U4449 (N_4449,N_1830,N_362);
nand U4450 (N_4450,N_1461,N_675);
and U4451 (N_4451,N_1671,N_526);
xor U4452 (N_4452,N_27,N_1524);
nor U4453 (N_4453,N_1737,N_21);
nor U4454 (N_4454,N_762,N_463);
nor U4455 (N_4455,N_606,N_1232);
or U4456 (N_4456,N_1451,N_284);
nand U4457 (N_4457,N_2168,N_1945);
or U4458 (N_4458,N_1242,N_1156);
and U4459 (N_4459,N_1404,N_490);
nor U4460 (N_4460,N_1278,N_572);
nor U4461 (N_4461,N_1259,N_880);
nand U4462 (N_4462,N_2115,N_330);
and U4463 (N_4463,N_2313,N_1435);
nor U4464 (N_4464,N_712,N_2038);
nor U4465 (N_4465,N_890,N_2093);
nor U4466 (N_4466,N_605,N_2432);
or U4467 (N_4467,N_1537,N_799);
nor U4468 (N_4468,N_137,N_271);
nand U4469 (N_4469,N_1413,N_301);
and U4470 (N_4470,N_2401,N_679);
xnor U4471 (N_4471,N_2380,N_481);
nor U4472 (N_4472,N_1512,N_1087);
and U4473 (N_4473,N_1917,N_581);
xnor U4474 (N_4474,N_506,N_2389);
xnor U4475 (N_4475,N_2366,N_1999);
nand U4476 (N_4476,N_2487,N_1064);
nand U4477 (N_4477,N_530,N_2205);
and U4478 (N_4478,N_2253,N_1291);
and U4479 (N_4479,N_213,N_1383);
and U4480 (N_4480,N_985,N_1665);
nor U4481 (N_4481,N_694,N_2434);
nor U4482 (N_4482,N_1261,N_1494);
nor U4483 (N_4483,N_1705,N_849);
and U4484 (N_4484,N_849,N_246);
and U4485 (N_4485,N_1773,N_817);
xor U4486 (N_4486,N_649,N_2064);
xor U4487 (N_4487,N_252,N_401);
or U4488 (N_4488,N_100,N_1297);
nor U4489 (N_4489,N_2165,N_1626);
nor U4490 (N_4490,N_2413,N_1124);
and U4491 (N_4491,N_14,N_946);
or U4492 (N_4492,N_753,N_690);
nor U4493 (N_4493,N_2227,N_1931);
nand U4494 (N_4494,N_1107,N_860);
nand U4495 (N_4495,N_1063,N_1612);
and U4496 (N_4496,N_1712,N_856);
xnor U4497 (N_4497,N_783,N_2029);
xor U4498 (N_4498,N_383,N_249);
and U4499 (N_4499,N_235,N_1265);
or U4500 (N_4500,N_723,N_356);
and U4501 (N_4501,N_2111,N_1695);
nand U4502 (N_4502,N_52,N_2007);
nor U4503 (N_4503,N_775,N_1387);
or U4504 (N_4504,N_418,N_1248);
xnor U4505 (N_4505,N_2486,N_2444);
or U4506 (N_4506,N_2496,N_840);
nor U4507 (N_4507,N_1553,N_1653);
nand U4508 (N_4508,N_1004,N_2003);
or U4509 (N_4509,N_1822,N_1041);
or U4510 (N_4510,N_1837,N_79);
or U4511 (N_4511,N_1148,N_193);
or U4512 (N_4512,N_2115,N_699);
or U4513 (N_4513,N_2476,N_1559);
or U4514 (N_4514,N_24,N_358);
or U4515 (N_4515,N_799,N_1842);
nand U4516 (N_4516,N_1199,N_1574);
and U4517 (N_4517,N_1143,N_2465);
or U4518 (N_4518,N_443,N_2023);
nand U4519 (N_4519,N_2332,N_797);
nand U4520 (N_4520,N_1322,N_1611);
nand U4521 (N_4521,N_1925,N_2408);
and U4522 (N_4522,N_611,N_783);
nand U4523 (N_4523,N_1971,N_1171);
or U4524 (N_4524,N_1700,N_372);
xnor U4525 (N_4525,N_2398,N_424);
or U4526 (N_4526,N_777,N_724);
xnor U4527 (N_4527,N_2463,N_2027);
or U4528 (N_4528,N_1435,N_2317);
nand U4529 (N_4529,N_2069,N_1336);
or U4530 (N_4530,N_1235,N_1289);
nand U4531 (N_4531,N_406,N_2401);
nor U4532 (N_4532,N_1439,N_204);
and U4533 (N_4533,N_536,N_2140);
xnor U4534 (N_4534,N_484,N_372);
or U4535 (N_4535,N_296,N_127);
or U4536 (N_4536,N_2090,N_138);
or U4537 (N_4537,N_818,N_1227);
and U4538 (N_4538,N_1039,N_1028);
or U4539 (N_4539,N_1924,N_1986);
xor U4540 (N_4540,N_800,N_1779);
nor U4541 (N_4541,N_2464,N_1213);
nand U4542 (N_4542,N_136,N_1220);
nand U4543 (N_4543,N_2453,N_112);
and U4544 (N_4544,N_2400,N_1577);
and U4545 (N_4545,N_940,N_1068);
nand U4546 (N_4546,N_1612,N_533);
or U4547 (N_4547,N_1417,N_2137);
or U4548 (N_4548,N_724,N_70);
and U4549 (N_4549,N_2338,N_873);
and U4550 (N_4550,N_2449,N_1084);
and U4551 (N_4551,N_1209,N_764);
or U4552 (N_4552,N_1419,N_1661);
or U4553 (N_4553,N_1478,N_1305);
or U4554 (N_4554,N_2065,N_428);
nand U4555 (N_4555,N_88,N_73);
or U4556 (N_4556,N_1362,N_558);
nand U4557 (N_4557,N_1450,N_1557);
nand U4558 (N_4558,N_182,N_998);
and U4559 (N_4559,N_466,N_2015);
nor U4560 (N_4560,N_1894,N_1304);
or U4561 (N_4561,N_750,N_1936);
nor U4562 (N_4562,N_701,N_1962);
or U4563 (N_4563,N_1859,N_78);
nand U4564 (N_4564,N_205,N_1581);
nor U4565 (N_4565,N_1896,N_2339);
nor U4566 (N_4566,N_2204,N_749);
and U4567 (N_4567,N_508,N_2448);
xor U4568 (N_4568,N_938,N_1164);
xor U4569 (N_4569,N_733,N_1228);
nand U4570 (N_4570,N_1424,N_1976);
nor U4571 (N_4571,N_59,N_1886);
xnor U4572 (N_4572,N_758,N_2381);
nor U4573 (N_4573,N_2133,N_2169);
nand U4574 (N_4574,N_439,N_2351);
and U4575 (N_4575,N_1974,N_114);
xor U4576 (N_4576,N_1130,N_301);
and U4577 (N_4577,N_1407,N_143);
nor U4578 (N_4578,N_1477,N_1116);
or U4579 (N_4579,N_198,N_873);
nor U4580 (N_4580,N_2263,N_584);
nor U4581 (N_4581,N_1206,N_705);
xnor U4582 (N_4582,N_617,N_889);
and U4583 (N_4583,N_271,N_1365);
xor U4584 (N_4584,N_2202,N_774);
nand U4585 (N_4585,N_771,N_280);
nand U4586 (N_4586,N_242,N_87);
xnor U4587 (N_4587,N_1026,N_1984);
nand U4588 (N_4588,N_1863,N_1251);
xor U4589 (N_4589,N_640,N_241);
nor U4590 (N_4590,N_1580,N_1592);
or U4591 (N_4591,N_2484,N_907);
or U4592 (N_4592,N_639,N_267);
nor U4593 (N_4593,N_719,N_923);
nand U4594 (N_4594,N_1469,N_750);
and U4595 (N_4595,N_1220,N_2);
nand U4596 (N_4596,N_1357,N_679);
nand U4597 (N_4597,N_2252,N_2287);
and U4598 (N_4598,N_1433,N_1603);
xor U4599 (N_4599,N_23,N_177);
and U4600 (N_4600,N_287,N_390);
xnor U4601 (N_4601,N_1959,N_712);
or U4602 (N_4602,N_2129,N_650);
and U4603 (N_4603,N_1247,N_1945);
or U4604 (N_4604,N_1184,N_2111);
xnor U4605 (N_4605,N_526,N_711);
nor U4606 (N_4606,N_1872,N_74);
and U4607 (N_4607,N_899,N_481);
and U4608 (N_4608,N_816,N_738);
xor U4609 (N_4609,N_1377,N_593);
and U4610 (N_4610,N_386,N_1597);
nand U4611 (N_4611,N_864,N_243);
or U4612 (N_4612,N_2341,N_540);
and U4613 (N_4613,N_1418,N_2280);
and U4614 (N_4614,N_995,N_988);
xor U4615 (N_4615,N_1575,N_1300);
nor U4616 (N_4616,N_402,N_1628);
nor U4617 (N_4617,N_1857,N_1934);
nand U4618 (N_4618,N_377,N_1275);
xnor U4619 (N_4619,N_219,N_749);
xor U4620 (N_4620,N_1030,N_1958);
nand U4621 (N_4621,N_990,N_2401);
nand U4622 (N_4622,N_1762,N_225);
or U4623 (N_4623,N_1299,N_696);
nor U4624 (N_4624,N_1372,N_650);
and U4625 (N_4625,N_1296,N_2459);
xnor U4626 (N_4626,N_49,N_2080);
nor U4627 (N_4627,N_2268,N_2257);
xnor U4628 (N_4628,N_1218,N_126);
nand U4629 (N_4629,N_730,N_1530);
xnor U4630 (N_4630,N_390,N_1800);
nor U4631 (N_4631,N_2170,N_82);
nor U4632 (N_4632,N_914,N_2218);
xor U4633 (N_4633,N_2044,N_590);
nor U4634 (N_4634,N_1,N_1741);
and U4635 (N_4635,N_615,N_1661);
xor U4636 (N_4636,N_1004,N_498);
and U4637 (N_4637,N_202,N_652);
and U4638 (N_4638,N_861,N_1924);
xnor U4639 (N_4639,N_1829,N_776);
and U4640 (N_4640,N_1714,N_1821);
nand U4641 (N_4641,N_888,N_462);
nor U4642 (N_4642,N_1323,N_2107);
nand U4643 (N_4643,N_1315,N_1806);
and U4644 (N_4644,N_820,N_1291);
nor U4645 (N_4645,N_1065,N_2470);
xnor U4646 (N_4646,N_2137,N_419);
nor U4647 (N_4647,N_361,N_20);
and U4648 (N_4648,N_1540,N_163);
and U4649 (N_4649,N_172,N_1322);
nor U4650 (N_4650,N_996,N_315);
and U4651 (N_4651,N_1132,N_1381);
or U4652 (N_4652,N_1254,N_1747);
nor U4653 (N_4653,N_1087,N_1942);
nand U4654 (N_4654,N_225,N_190);
nor U4655 (N_4655,N_1783,N_1486);
nand U4656 (N_4656,N_1393,N_530);
nor U4657 (N_4657,N_1709,N_1112);
and U4658 (N_4658,N_2085,N_1475);
nor U4659 (N_4659,N_204,N_2011);
nand U4660 (N_4660,N_2086,N_739);
or U4661 (N_4661,N_1007,N_2163);
xnor U4662 (N_4662,N_459,N_118);
nand U4663 (N_4663,N_588,N_850);
and U4664 (N_4664,N_2326,N_415);
and U4665 (N_4665,N_1034,N_1615);
xnor U4666 (N_4666,N_1347,N_1164);
and U4667 (N_4667,N_1244,N_1333);
or U4668 (N_4668,N_1192,N_5);
and U4669 (N_4669,N_1828,N_349);
nand U4670 (N_4670,N_522,N_1848);
or U4671 (N_4671,N_1119,N_1938);
nor U4672 (N_4672,N_2290,N_2170);
or U4673 (N_4673,N_497,N_1704);
or U4674 (N_4674,N_2269,N_239);
or U4675 (N_4675,N_1098,N_2151);
and U4676 (N_4676,N_2324,N_1971);
xnor U4677 (N_4677,N_2161,N_1607);
nand U4678 (N_4678,N_2062,N_1661);
xor U4679 (N_4679,N_140,N_2151);
nor U4680 (N_4680,N_1890,N_1332);
and U4681 (N_4681,N_917,N_107);
xor U4682 (N_4682,N_2294,N_892);
nor U4683 (N_4683,N_804,N_919);
nor U4684 (N_4684,N_784,N_696);
nand U4685 (N_4685,N_1140,N_1933);
nor U4686 (N_4686,N_851,N_1901);
nor U4687 (N_4687,N_679,N_1407);
nand U4688 (N_4688,N_1133,N_1974);
xnor U4689 (N_4689,N_12,N_516);
and U4690 (N_4690,N_2474,N_924);
or U4691 (N_4691,N_445,N_1291);
nand U4692 (N_4692,N_465,N_2109);
or U4693 (N_4693,N_1254,N_737);
nand U4694 (N_4694,N_2329,N_1478);
and U4695 (N_4695,N_365,N_569);
nand U4696 (N_4696,N_1114,N_996);
and U4697 (N_4697,N_1422,N_1461);
xor U4698 (N_4698,N_2497,N_947);
or U4699 (N_4699,N_2319,N_686);
nand U4700 (N_4700,N_2342,N_1377);
and U4701 (N_4701,N_599,N_350);
xnor U4702 (N_4702,N_2407,N_32);
nand U4703 (N_4703,N_96,N_1947);
xor U4704 (N_4704,N_986,N_1010);
and U4705 (N_4705,N_927,N_1485);
nor U4706 (N_4706,N_1392,N_2462);
nor U4707 (N_4707,N_2397,N_335);
nand U4708 (N_4708,N_855,N_2104);
nand U4709 (N_4709,N_1298,N_1932);
xnor U4710 (N_4710,N_1701,N_97);
nand U4711 (N_4711,N_843,N_1222);
nand U4712 (N_4712,N_998,N_848);
or U4713 (N_4713,N_2477,N_2409);
and U4714 (N_4714,N_813,N_1078);
or U4715 (N_4715,N_1772,N_675);
nand U4716 (N_4716,N_1954,N_180);
xor U4717 (N_4717,N_2054,N_1008);
or U4718 (N_4718,N_1682,N_2449);
nand U4719 (N_4719,N_1351,N_1950);
nor U4720 (N_4720,N_128,N_178);
xor U4721 (N_4721,N_753,N_543);
and U4722 (N_4722,N_1829,N_56);
nor U4723 (N_4723,N_1961,N_397);
or U4724 (N_4724,N_793,N_90);
nand U4725 (N_4725,N_140,N_2059);
or U4726 (N_4726,N_2016,N_2399);
and U4727 (N_4727,N_1067,N_1185);
xor U4728 (N_4728,N_1058,N_2364);
nor U4729 (N_4729,N_1446,N_1408);
nand U4730 (N_4730,N_1090,N_202);
xnor U4731 (N_4731,N_2420,N_193);
nor U4732 (N_4732,N_1701,N_500);
nor U4733 (N_4733,N_2314,N_391);
nand U4734 (N_4734,N_1740,N_9);
nand U4735 (N_4735,N_828,N_940);
or U4736 (N_4736,N_1054,N_2423);
nor U4737 (N_4737,N_2135,N_2109);
xnor U4738 (N_4738,N_1646,N_1304);
and U4739 (N_4739,N_1864,N_251);
nor U4740 (N_4740,N_660,N_1475);
xor U4741 (N_4741,N_1848,N_379);
nor U4742 (N_4742,N_1388,N_1040);
nand U4743 (N_4743,N_251,N_746);
and U4744 (N_4744,N_848,N_199);
xnor U4745 (N_4745,N_1169,N_1079);
nor U4746 (N_4746,N_1141,N_783);
and U4747 (N_4747,N_949,N_1994);
or U4748 (N_4748,N_2304,N_1091);
and U4749 (N_4749,N_1512,N_266);
nor U4750 (N_4750,N_1831,N_1483);
nand U4751 (N_4751,N_814,N_2140);
or U4752 (N_4752,N_2221,N_2396);
xnor U4753 (N_4753,N_677,N_160);
nand U4754 (N_4754,N_1185,N_660);
nand U4755 (N_4755,N_1135,N_1429);
nor U4756 (N_4756,N_2207,N_868);
nor U4757 (N_4757,N_1785,N_1576);
nand U4758 (N_4758,N_1692,N_2181);
and U4759 (N_4759,N_2031,N_86);
and U4760 (N_4760,N_232,N_2239);
xnor U4761 (N_4761,N_324,N_2383);
nor U4762 (N_4762,N_2423,N_302);
or U4763 (N_4763,N_836,N_2243);
or U4764 (N_4764,N_1466,N_851);
nor U4765 (N_4765,N_2373,N_2437);
nor U4766 (N_4766,N_521,N_1132);
or U4767 (N_4767,N_2163,N_1063);
and U4768 (N_4768,N_1286,N_55);
or U4769 (N_4769,N_1989,N_1021);
nand U4770 (N_4770,N_1494,N_2042);
nand U4771 (N_4771,N_373,N_169);
and U4772 (N_4772,N_327,N_2245);
or U4773 (N_4773,N_1003,N_2436);
or U4774 (N_4774,N_1390,N_160);
nor U4775 (N_4775,N_1523,N_77);
and U4776 (N_4776,N_1583,N_1527);
nand U4777 (N_4777,N_1078,N_1324);
nor U4778 (N_4778,N_143,N_1316);
or U4779 (N_4779,N_2335,N_1485);
nand U4780 (N_4780,N_237,N_213);
and U4781 (N_4781,N_1778,N_705);
nor U4782 (N_4782,N_922,N_1089);
nor U4783 (N_4783,N_639,N_1987);
xnor U4784 (N_4784,N_1518,N_114);
or U4785 (N_4785,N_579,N_645);
xor U4786 (N_4786,N_377,N_78);
nand U4787 (N_4787,N_443,N_1729);
and U4788 (N_4788,N_2141,N_2498);
xor U4789 (N_4789,N_1919,N_84);
or U4790 (N_4790,N_1336,N_835);
nor U4791 (N_4791,N_2455,N_790);
nand U4792 (N_4792,N_502,N_438);
and U4793 (N_4793,N_576,N_1904);
and U4794 (N_4794,N_1110,N_1643);
nand U4795 (N_4795,N_1869,N_2460);
nand U4796 (N_4796,N_613,N_858);
xnor U4797 (N_4797,N_327,N_2225);
and U4798 (N_4798,N_939,N_33);
nand U4799 (N_4799,N_302,N_235);
or U4800 (N_4800,N_1672,N_450);
or U4801 (N_4801,N_903,N_376);
or U4802 (N_4802,N_2469,N_340);
xor U4803 (N_4803,N_2020,N_2242);
nor U4804 (N_4804,N_812,N_170);
nand U4805 (N_4805,N_788,N_2173);
xnor U4806 (N_4806,N_2068,N_1564);
or U4807 (N_4807,N_239,N_63);
and U4808 (N_4808,N_2262,N_238);
nand U4809 (N_4809,N_1927,N_482);
nor U4810 (N_4810,N_431,N_29);
or U4811 (N_4811,N_0,N_941);
xnor U4812 (N_4812,N_1418,N_2233);
nor U4813 (N_4813,N_4,N_819);
nor U4814 (N_4814,N_150,N_1497);
nand U4815 (N_4815,N_1941,N_522);
xnor U4816 (N_4816,N_2085,N_1324);
or U4817 (N_4817,N_318,N_201);
nor U4818 (N_4818,N_2138,N_1615);
xnor U4819 (N_4819,N_1907,N_1182);
nor U4820 (N_4820,N_649,N_1401);
xor U4821 (N_4821,N_851,N_665);
nor U4822 (N_4822,N_619,N_383);
or U4823 (N_4823,N_84,N_396);
or U4824 (N_4824,N_2082,N_1725);
and U4825 (N_4825,N_1212,N_826);
nor U4826 (N_4826,N_903,N_2038);
and U4827 (N_4827,N_2041,N_275);
nand U4828 (N_4828,N_2425,N_1092);
nor U4829 (N_4829,N_2284,N_532);
or U4830 (N_4830,N_986,N_1703);
and U4831 (N_4831,N_1318,N_2137);
xor U4832 (N_4832,N_113,N_531);
or U4833 (N_4833,N_184,N_759);
nand U4834 (N_4834,N_887,N_1210);
and U4835 (N_4835,N_496,N_420);
and U4836 (N_4836,N_2028,N_673);
and U4837 (N_4837,N_1890,N_1618);
and U4838 (N_4838,N_2364,N_824);
xor U4839 (N_4839,N_1455,N_1295);
nand U4840 (N_4840,N_1914,N_6);
xnor U4841 (N_4841,N_318,N_177);
nand U4842 (N_4842,N_1999,N_718);
or U4843 (N_4843,N_2103,N_1727);
and U4844 (N_4844,N_2101,N_1143);
or U4845 (N_4845,N_1230,N_1841);
xnor U4846 (N_4846,N_364,N_49);
nor U4847 (N_4847,N_1336,N_2403);
or U4848 (N_4848,N_56,N_1960);
or U4849 (N_4849,N_1225,N_197);
or U4850 (N_4850,N_1661,N_389);
nand U4851 (N_4851,N_855,N_2323);
nand U4852 (N_4852,N_2463,N_1204);
nor U4853 (N_4853,N_1463,N_1533);
nor U4854 (N_4854,N_1079,N_1684);
nand U4855 (N_4855,N_551,N_1629);
xnor U4856 (N_4856,N_2492,N_1397);
and U4857 (N_4857,N_2090,N_1296);
nor U4858 (N_4858,N_110,N_260);
xnor U4859 (N_4859,N_1854,N_1324);
and U4860 (N_4860,N_1400,N_1267);
or U4861 (N_4861,N_2318,N_1596);
xor U4862 (N_4862,N_2052,N_961);
nor U4863 (N_4863,N_39,N_828);
nor U4864 (N_4864,N_1471,N_268);
or U4865 (N_4865,N_1768,N_1413);
nor U4866 (N_4866,N_1393,N_2202);
and U4867 (N_4867,N_1073,N_1618);
nand U4868 (N_4868,N_317,N_963);
nor U4869 (N_4869,N_1391,N_1526);
xor U4870 (N_4870,N_1921,N_578);
and U4871 (N_4871,N_2461,N_819);
xnor U4872 (N_4872,N_1095,N_1846);
nand U4873 (N_4873,N_1803,N_2017);
and U4874 (N_4874,N_1943,N_1891);
and U4875 (N_4875,N_2247,N_1752);
or U4876 (N_4876,N_2129,N_180);
xor U4877 (N_4877,N_799,N_1259);
or U4878 (N_4878,N_989,N_1798);
or U4879 (N_4879,N_582,N_2193);
nand U4880 (N_4880,N_1933,N_1255);
xor U4881 (N_4881,N_839,N_2110);
nor U4882 (N_4882,N_612,N_99);
xor U4883 (N_4883,N_1317,N_468);
xnor U4884 (N_4884,N_2208,N_2252);
nor U4885 (N_4885,N_644,N_653);
nor U4886 (N_4886,N_996,N_472);
or U4887 (N_4887,N_2069,N_767);
or U4888 (N_4888,N_1502,N_1665);
nand U4889 (N_4889,N_1911,N_595);
nor U4890 (N_4890,N_2356,N_2381);
and U4891 (N_4891,N_2050,N_2361);
and U4892 (N_4892,N_2426,N_2427);
nand U4893 (N_4893,N_332,N_2063);
nor U4894 (N_4894,N_695,N_1755);
nand U4895 (N_4895,N_1535,N_1151);
nand U4896 (N_4896,N_1206,N_1073);
xor U4897 (N_4897,N_1713,N_842);
and U4898 (N_4898,N_361,N_2174);
xor U4899 (N_4899,N_189,N_1481);
xnor U4900 (N_4900,N_894,N_644);
or U4901 (N_4901,N_132,N_910);
and U4902 (N_4902,N_966,N_2144);
nor U4903 (N_4903,N_829,N_2385);
xnor U4904 (N_4904,N_1107,N_807);
or U4905 (N_4905,N_438,N_656);
nor U4906 (N_4906,N_1746,N_511);
nor U4907 (N_4907,N_2072,N_1796);
or U4908 (N_4908,N_2306,N_1446);
nor U4909 (N_4909,N_2050,N_501);
or U4910 (N_4910,N_734,N_2298);
nand U4911 (N_4911,N_971,N_1287);
and U4912 (N_4912,N_2153,N_321);
and U4913 (N_4913,N_88,N_1823);
nand U4914 (N_4914,N_1802,N_2431);
and U4915 (N_4915,N_119,N_2225);
nand U4916 (N_4916,N_882,N_547);
and U4917 (N_4917,N_906,N_1010);
and U4918 (N_4918,N_1380,N_605);
or U4919 (N_4919,N_317,N_1002);
nand U4920 (N_4920,N_689,N_1120);
or U4921 (N_4921,N_1642,N_2475);
and U4922 (N_4922,N_1935,N_1693);
or U4923 (N_4923,N_1244,N_1595);
or U4924 (N_4924,N_1205,N_1242);
nand U4925 (N_4925,N_1791,N_1733);
xor U4926 (N_4926,N_1208,N_724);
xnor U4927 (N_4927,N_1306,N_476);
or U4928 (N_4928,N_925,N_1380);
nor U4929 (N_4929,N_1206,N_1369);
nor U4930 (N_4930,N_1430,N_388);
and U4931 (N_4931,N_881,N_1848);
xor U4932 (N_4932,N_1936,N_234);
nand U4933 (N_4933,N_2454,N_356);
xor U4934 (N_4934,N_220,N_1301);
and U4935 (N_4935,N_605,N_2245);
and U4936 (N_4936,N_2126,N_2165);
or U4937 (N_4937,N_2265,N_666);
or U4938 (N_4938,N_1147,N_1939);
xor U4939 (N_4939,N_72,N_1921);
xor U4940 (N_4940,N_987,N_1336);
or U4941 (N_4941,N_526,N_218);
nor U4942 (N_4942,N_319,N_1662);
nand U4943 (N_4943,N_1560,N_2207);
nor U4944 (N_4944,N_394,N_611);
xor U4945 (N_4945,N_2433,N_947);
nor U4946 (N_4946,N_63,N_869);
nor U4947 (N_4947,N_595,N_810);
xnor U4948 (N_4948,N_203,N_1451);
or U4949 (N_4949,N_2305,N_1618);
nor U4950 (N_4950,N_728,N_511);
or U4951 (N_4951,N_2124,N_1313);
nand U4952 (N_4952,N_1458,N_1758);
and U4953 (N_4953,N_2174,N_1306);
and U4954 (N_4954,N_2031,N_2446);
xnor U4955 (N_4955,N_847,N_1390);
or U4956 (N_4956,N_619,N_452);
xor U4957 (N_4957,N_1120,N_2043);
xnor U4958 (N_4958,N_2090,N_1597);
nand U4959 (N_4959,N_317,N_1650);
and U4960 (N_4960,N_86,N_157);
or U4961 (N_4961,N_1986,N_2423);
and U4962 (N_4962,N_1423,N_2452);
xor U4963 (N_4963,N_852,N_2061);
nand U4964 (N_4964,N_801,N_29);
or U4965 (N_4965,N_740,N_1206);
nor U4966 (N_4966,N_702,N_830);
nor U4967 (N_4967,N_1985,N_194);
nand U4968 (N_4968,N_879,N_302);
nor U4969 (N_4969,N_1396,N_122);
nor U4970 (N_4970,N_708,N_1715);
or U4971 (N_4971,N_1012,N_604);
nand U4972 (N_4972,N_2377,N_733);
xnor U4973 (N_4973,N_1563,N_2406);
xor U4974 (N_4974,N_1892,N_448);
and U4975 (N_4975,N_74,N_1228);
and U4976 (N_4976,N_2051,N_331);
nand U4977 (N_4977,N_1503,N_1904);
and U4978 (N_4978,N_1676,N_1738);
and U4979 (N_4979,N_390,N_596);
or U4980 (N_4980,N_102,N_1561);
and U4981 (N_4981,N_291,N_60);
or U4982 (N_4982,N_1651,N_479);
nand U4983 (N_4983,N_1079,N_827);
nor U4984 (N_4984,N_1620,N_1118);
and U4985 (N_4985,N_1992,N_2301);
or U4986 (N_4986,N_814,N_1017);
and U4987 (N_4987,N_1341,N_1914);
or U4988 (N_4988,N_1904,N_1181);
xnor U4989 (N_4989,N_508,N_716);
or U4990 (N_4990,N_816,N_1946);
xor U4991 (N_4991,N_13,N_316);
nor U4992 (N_4992,N_1378,N_575);
nor U4993 (N_4993,N_1343,N_808);
xor U4994 (N_4994,N_1015,N_1152);
nand U4995 (N_4995,N_1380,N_2012);
xor U4996 (N_4996,N_1198,N_2186);
xor U4997 (N_4997,N_1969,N_2438);
nor U4998 (N_4998,N_1846,N_142);
nor U4999 (N_4999,N_817,N_35);
and U5000 (N_5000,N_4296,N_3540);
nand U5001 (N_5001,N_3520,N_4547);
and U5002 (N_5002,N_4095,N_4026);
nor U5003 (N_5003,N_3419,N_3867);
and U5004 (N_5004,N_4705,N_4925);
nor U5005 (N_5005,N_2944,N_4678);
or U5006 (N_5006,N_4040,N_3715);
xnor U5007 (N_5007,N_3376,N_2604);
nand U5008 (N_5008,N_3707,N_3687);
and U5009 (N_5009,N_3193,N_2546);
or U5010 (N_5010,N_4598,N_3802);
and U5011 (N_5011,N_4195,N_3406);
nor U5012 (N_5012,N_4029,N_3442);
and U5013 (N_5013,N_2791,N_3990);
xnor U5014 (N_5014,N_4256,N_4315);
xnor U5015 (N_5015,N_4197,N_3784);
nor U5016 (N_5016,N_4438,N_4441);
nand U5017 (N_5017,N_2613,N_2807);
nand U5018 (N_5018,N_3674,N_2889);
nand U5019 (N_5019,N_4389,N_2759);
nand U5020 (N_5020,N_4929,N_3813);
and U5021 (N_5021,N_4071,N_4770);
or U5022 (N_5022,N_4137,N_4865);
and U5023 (N_5023,N_4644,N_3670);
nor U5024 (N_5024,N_4603,N_4838);
xor U5025 (N_5025,N_4001,N_4834);
and U5026 (N_5026,N_4774,N_2823);
or U5027 (N_5027,N_4362,N_4152);
and U5028 (N_5028,N_4236,N_3247);
or U5029 (N_5029,N_4188,N_4877);
nor U5030 (N_5030,N_2596,N_4692);
nand U5031 (N_5031,N_3109,N_4035);
nand U5032 (N_5032,N_3830,N_3129);
nand U5033 (N_5033,N_3497,N_3607);
xor U5034 (N_5034,N_4114,N_3553);
xor U5035 (N_5035,N_3523,N_4915);
and U5036 (N_5036,N_4457,N_4239);
nand U5037 (N_5037,N_4786,N_2548);
or U5038 (N_5038,N_3041,N_2894);
nand U5039 (N_5039,N_3000,N_4343);
and U5040 (N_5040,N_4396,N_4672);
nor U5041 (N_5041,N_3593,N_4076);
nor U5042 (N_5042,N_4088,N_2668);
nand U5043 (N_5043,N_3775,N_2501);
nand U5044 (N_5044,N_2614,N_3103);
and U5045 (N_5045,N_2976,N_4017);
and U5046 (N_5046,N_2930,N_4111);
nand U5047 (N_5047,N_4156,N_4046);
xor U5048 (N_5048,N_2860,N_3626);
or U5049 (N_5049,N_3199,N_3810);
nor U5050 (N_5050,N_4686,N_3112);
or U5051 (N_5051,N_3716,N_4119);
and U5052 (N_5052,N_4683,N_4292);
xor U5053 (N_5053,N_3703,N_3495);
nor U5054 (N_5054,N_3496,N_4730);
and U5055 (N_5055,N_4179,N_4828);
xor U5056 (N_5056,N_2628,N_3086);
and U5057 (N_5057,N_4162,N_4320);
or U5058 (N_5058,N_3250,N_3011);
nor U5059 (N_5059,N_2568,N_3032);
nand U5060 (N_5060,N_4344,N_2907);
xnor U5061 (N_5061,N_3663,N_4328);
and U5062 (N_5062,N_4702,N_2964);
xnor U5063 (N_5063,N_4671,N_3913);
nand U5064 (N_5064,N_4492,N_3408);
nand U5065 (N_5065,N_3976,N_4388);
nand U5066 (N_5066,N_4888,N_2863);
nor U5067 (N_5067,N_2772,N_4742);
nor U5068 (N_5068,N_4975,N_2936);
nand U5069 (N_5069,N_3870,N_2928);
nand U5070 (N_5070,N_4129,N_3474);
or U5071 (N_5071,N_2890,N_2839);
nand U5072 (N_5072,N_2705,N_4178);
or U5073 (N_5073,N_3794,N_4715);
nor U5074 (N_5074,N_2747,N_4850);
or U5075 (N_5075,N_4727,N_4766);
xnor U5076 (N_5076,N_4613,N_4094);
and U5077 (N_5077,N_3277,N_2933);
nor U5078 (N_5078,N_4777,N_4995);
nor U5079 (N_5079,N_2808,N_4375);
nor U5080 (N_5080,N_2695,N_2723);
xor U5081 (N_5081,N_4147,N_3182);
or U5082 (N_5082,N_4946,N_2656);
nor U5083 (N_5083,N_2749,N_4658);
and U5084 (N_5084,N_4005,N_4670);
nor U5085 (N_5085,N_4050,N_3157);
nor U5086 (N_5086,N_4918,N_3194);
xor U5087 (N_5087,N_4845,N_4409);
nand U5088 (N_5088,N_3627,N_4606);
or U5089 (N_5089,N_4532,N_3565);
nand U5090 (N_5090,N_4793,N_4879);
and U5091 (N_5091,N_4754,N_4745);
and U5092 (N_5092,N_3248,N_3908);
nor U5093 (N_5093,N_4294,N_4181);
or U5094 (N_5094,N_3123,N_4627);
or U5095 (N_5095,N_2554,N_4841);
nand U5096 (N_5096,N_2720,N_3325);
nor U5097 (N_5097,N_3685,N_3615);
nand U5098 (N_5098,N_2531,N_3279);
or U5099 (N_5099,N_4779,N_4552);
nand U5100 (N_5100,N_4165,N_4169);
and U5101 (N_5101,N_3842,N_4269);
nor U5102 (N_5102,N_2550,N_3773);
or U5103 (N_5103,N_3216,N_4894);
nor U5104 (N_5104,N_2711,N_4191);
and U5105 (N_5105,N_3057,N_4473);
and U5106 (N_5106,N_3768,N_4010);
nand U5107 (N_5107,N_2630,N_4529);
nor U5108 (N_5108,N_3375,N_3879);
nor U5109 (N_5109,N_4430,N_3145);
xor U5110 (N_5110,N_4947,N_3146);
nor U5111 (N_5111,N_4788,N_4726);
and U5112 (N_5112,N_2732,N_4661);
xor U5113 (N_5113,N_4531,N_3718);
nor U5114 (N_5114,N_3107,N_3394);
xor U5115 (N_5115,N_2972,N_3273);
nand U5116 (N_5116,N_3823,N_2675);
nor U5117 (N_5117,N_3075,N_4940);
xor U5118 (N_5118,N_2731,N_4124);
xor U5119 (N_5119,N_3820,N_3736);
xnor U5120 (N_5120,N_3336,N_4610);
xor U5121 (N_5121,N_2619,N_4330);
and U5122 (N_5122,N_2858,N_3033);
xnor U5123 (N_5123,N_3480,N_3727);
and U5124 (N_5124,N_2811,N_3809);
or U5125 (N_5125,N_2694,N_4674);
nand U5126 (N_5126,N_4681,N_3306);
or U5127 (N_5127,N_2995,N_3875);
nand U5128 (N_5128,N_2582,N_2951);
nand U5129 (N_5129,N_4589,N_2799);
or U5130 (N_5130,N_3027,N_4075);
nand U5131 (N_5131,N_3108,N_4371);
nor U5132 (N_5132,N_3907,N_3330);
and U5133 (N_5133,N_4536,N_4134);
xnor U5134 (N_5134,N_4632,N_3237);
xor U5135 (N_5135,N_2909,N_3758);
nand U5136 (N_5136,N_4876,N_2757);
xor U5137 (N_5137,N_4569,N_4813);
or U5138 (N_5138,N_4520,N_3945);
and U5139 (N_5139,N_2920,N_4666);
xnor U5140 (N_5140,N_4827,N_4423);
and U5141 (N_5141,N_2817,N_3585);
nand U5142 (N_5142,N_4283,N_3993);
xnor U5143 (N_5143,N_4937,N_4460);
nor U5144 (N_5144,N_4471,N_2954);
nor U5145 (N_5145,N_2804,N_2622);
and U5146 (N_5146,N_2555,N_3686);
and U5147 (N_5147,N_3743,N_4612);
or U5148 (N_5148,N_4298,N_3035);
or U5149 (N_5149,N_3457,N_2781);
nor U5150 (N_5150,N_4802,N_3084);
or U5151 (N_5151,N_3421,N_4693);
and U5152 (N_5152,N_4192,N_3555);
and U5153 (N_5153,N_3964,N_3452);
nand U5154 (N_5154,N_3456,N_2900);
nor U5155 (N_5155,N_4986,N_3921);
nand U5156 (N_5156,N_4537,N_2540);
xnor U5157 (N_5157,N_4893,N_4357);
nor U5158 (N_5158,N_4541,N_4695);
nor U5159 (N_5159,N_3988,N_4780);
and U5160 (N_5160,N_3056,N_3475);
or U5161 (N_5161,N_3811,N_4826);
and U5162 (N_5162,N_4381,N_4122);
nor U5163 (N_5163,N_4920,N_2827);
xnor U5164 (N_5164,N_2657,N_3046);
xnor U5165 (N_5165,N_4347,N_4271);
xnor U5166 (N_5166,N_4200,N_3415);
and U5167 (N_5167,N_3183,N_3601);
or U5168 (N_5168,N_2880,N_3938);
nor U5169 (N_5169,N_3096,N_4107);
nor U5170 (N_5170,N_3333,N_4450);
and U5171 (N_5171,N_4452,N_3625);
nand U5172 (N_5172,N_3239,N_3857);
nand U5173 (N_5173,N_4118,N_3040);
nand U5174 (N_5174,N_3085,N_4891);
nand U5175 (N_5175,N_2681,N_4437);
nor U5176 (N_5176,N_2785,N_2896);
nor U5177 (N_5177,N_4572,N_4416);
xor U5178 (N_5178,N_4775,N_3749);
and U5179 (N_5179,N_4483,N_3803);
xor U5180 (N_5180,N_4135,N_4096);
xnor U5181 (N_5181,N_3577,N_2690);
or U5182 (N_5182,N_4168,N_3587);
nand U5183 (N_5183,N_4277,N_4494);
or U5184 (N_5184,N_2979,N_3659);
nor U5185 (N_5185,N_3047,N_4718);
and U5186 (N_5186,N_4036,N_4484);
nand U5187 (N_5187,N_3087,N_4313);
nor U5188 (N_5188,N_3490,N_4262);
or U5189 (N_5189,N_3562,N_3789);
nand U5190 (N_5190,N_4739,N_4407);
and U5191 (N_5191,N_4800,N_4394);
and U5192 (N_5192,N_4020,N_2924);
xor U5193 (N_5193,N_3828,N_3090);
or U5194 (N_5194,N_3242,N_2561);
nand U5195 (N_5195,N_4664,N_4822);
nor U5196 (N_5196,N_3631,N_4317);
nand U5197 (N_5197,N_4098,N_4849);
nor U5198 (N_5198,N_4756,N_4854);
xnor U5199 (N_5199,N_4436,N_4032);
nor U5200 (N_5200,N_3481,N_3037);
xor U5201 (N_5201,N_3853,N_4190);
xor U5202 (N_5202,N_3644,N_3192);
nand U5203 (N_5203,N_3765,N_2788);
nand U5204 (N_5204,N_3016,N_4753);
or U5205 (N_5205,N_4382,N_2868);
nor U5206 (N_5206,N_3002,N_3966);
nor U5207 (N_5207,N_3606,N_2780);
or U5208 (N_5208,N_3787,N_3967);
or U5209 (N_5209,N_4089,N_2906);
xor U5210 (N_5210,N_3638,N_4044);
xnor U5211 (N_5211,N_2769,N_2629);
nand U5212 (N_5212,N_3939,N_3518);
and U5213 (N_5213,N_3095,N_2641);
xor U5214 (N_5214,N_4984,N_3837);
xnor U5215 (N_5215,N_3845,N_2997);
xnor U5216 (N_5216,N_2574,N_3259);
and U5217 (N_5217,N_2946,N_4377);
xnor U5218 (N_5218,N_4475,N_3671);
nand U5219 (N_5219,N_4791,N_3222);
nand U5220 (N_5220,N_3714,N_2605);
nor U5221 (N_5221,N_2973,N_4335);
and U5222 (N_5222,N_3717,N_3063);
or U5223 (N_5223,N_2506,N_4863);
or U5224 (N_5224,N_4732,N_3263);
nand U5225 (N_5225,N_3550,N_2787);
nor U5226 (N_5226,N_4799,N_3719);
nor U5227 (N_5227,N_4112,N_2524);
nor U5228 (N_5228,N_2625,N_3398);
and U5229 (N_5229,N_3253,N_3927);
nor U5230 (N_5230,N_2702,N_4604);
nand U5231 (N_5231,N_4812,N_3317);
or U5232 (N_5232,N_3458,N_3079);
nand U5233 (N_5233,N_4364,N_2576);
or U5234 (N_5234,N_2722,N_4213);
and U5235 (N_5235,N_4640,N_4723);
and U5236 (N_5236,N_3185,N_2833);
nor U5237 (N_5237,N_3159,N_4787);
nor U5238 (N_5238,N_3704,N_3249);
nor U5239 (N_5239,N_3175,N_3489);
or U5240 (N_5240,N_4143,N_3750);
nand U5241 (N_5241,N_3233,N_4591);
or U5242 (N_5242,N_4719,N_4261);
nor U5243 (N_5243,N_3600,N_4105);
nand U5244 (N_5244,N_2762,N_4016);
nand U5245 (N_5245,N_4852,N_4289);
nor U5246 (N_5246,N_2761,N_4383);
nand U5247 (N_5247,N_3397,N_3683);
and U5248 (N_5248,N_3323,N_4758);
nand U5249 (N_5249,N_3150,N_3653);
nand U5250 (N_5250,N_3563,N_3180);
nand U5251 (N_5251,N_3635,N_4138);
nor U5252 (N_5252,N_3948,N_3039);
or U5253 (N_5253,N_3729,N_3203);
nor U5254 (N_5254,N_4620,N_4291);
nor U5255 (N_5255,N_3384,N_2878);
xor U5256 (N_5256,N_4059,N_2969);
or U5257 (N_5257,N_4060,N_3302);
or U5258 (N_5258,N_3440,N_4468);
nand U5259 (N_5259,N_4744,N_4028);
nor U5260 (N_5260,N_4015,N_3486);
nand U5261 (N_5261,N_3891,N_3118);
nor U5262 (N_5262,N_2618,N_2527);
nor U5263 (N_5263,N_2663,N_4021);
and U5264 (N_5264,N_3545,N_4687);
nand U5265 (N_5265,N_4594,N_3774);
and U5266 (N_5266,N_3982,N_4548);
or U5267 (N_5267,N_2856,N_4585);
or U5268 (N_5268,N_4817,N_3825);
xor U5269 (N_5269,N_3660,N_2834);
or U5270 (N_5270,N_3706,N_3382);
and U5271 (N_5271,N_2935,N_4270);
and U5272 (N_5272,N_4284,N_3965);
xor U5273 (N_5273,N_4696,N_4159);
or U5274 (N_5274,N_4194,N_3065);
and U5275 (N_5275,N_3633,N_4631);
and U5276 (N_5276,N_2740,N_2961);
nor U5277 (N_5277,N_2719,N_3077);
xor U5278 (N_5278,N_4938,N_2899);
xnor U5279 (N_5279,N_2836,N_4480);
or U5280 (N_5280,N_4533,N_4209);
nor U5281 (N_5281,N_4338,N_3070);
xnor U5282 (N_5282,N_4916,N_3331);
nand U5283 (N_5283,N_3556,N_3334);
or U5284 (N_5284,N_3448,N_2543);
or U5285 (N_5285,N_2566,N_4587);
nand U5286 (N_5286,N_4078,N_4008);
nand U5287 (N_5287,N_4039,N_3636);
nand U5288 (N_5288,N_4225,N_3464);
nand U5289 (N_5289,N_3312,N_3113);
nand U5290 (N_5290,N_3925,N_3023);
nand U5291 (N_5291,N_4575,N_2507);
xnor U5292 (N_5292,N_4106,N_3733);
nand U5293 (N_5293,N_4265,N_4414);
xor U5294 (N_5294,N_4033,N_2931);
nor U5295 (N_5295,N_2638,N_3444);
nor U5296 (N_5296,N_2883,N_2825);
and U5297 (N_5297,N_4303,N_3932);
xor U5298 (N_5298,N_3735,N_3260);
nand U5299 (N_5299,N_4951,N_3238);
xnor U5300 (N_5300,N_3790,N_3501);
and U5301 (N_5301,N_2877,N_4231);
xnor U5302 (N_5302,N_2591,N_3015);
nand U5303 (N_5303,N_2750,N_2955);
and U5304 (N_5304,N_3591,N_3427);
nor U5305 (N_5305,N_4797,N_3903);
xnor U5306 (N_5306,N_2818,N_4496);
or U5307 (N_5307,N_4971,N_3447);
nor U5308 (N_5308,N_4934,N_2903);
nand U5309 (N_5309,N_3882,N_3169);
nor U5310 (N_5310,N_4691,N_3788);
and U5311 (N_5311,N_4148,N_3224);
and U5312 (N_5312,N_4058,N_2978);
and U5313 (N_5313,N_2876,N_4222);
nand U5314 (N_5314,N_3575,N_3962);
or U5315 (N_5315,N_4856,N_3554);
xor U5316 (N_5316,N_3251,N_2801);
and U5317 (N_5317,N_4830,N_4901);
nor U5318 (N_5318,N_4281,N_4969);
xor U5319 (N_5319,N_3099,N_4196);
nor U5320 (N_5320,N_2957,N_3286);
and U5321 (N_5321,N_2721,N_2819);
nand U5322 (N_5322,N_3763,N_4630);
nand U5323 (N_5323,N_2956,N_3779);
or U5324 (N_5324,N_3466,N_4871);
or U5325 (N_5325,N_4511,N_4646);
xor U5326 (N_5326,N_3564,N_3505);
nand U5327 (N_5327,N_2841,N_2926);
xnor U5328 (N_5328,N_3656,N_3576);
xor U5329 (N_5329,N_3485,N_3119);
and U5330 (N_5330,N_4996,N_2797);
and U5331 (N_5331,N_3167,N_3209);
or U5332 (N_5332,N_3934,N_4930);
or U5333 (N_5333,N_3269,N_3975);
nand U5334 (N_5334,N_2689,N_3815);
xor U5335 (N_5335,N_3073,N_3141);
xnor U5336 (N_5336,N_4085,N_3731);
or U5337 (N_5337,N_3400,N_4710);
and U5338 (N_5338,N_2885,N_4175);
or U5339 (N_5339,N_3477,N_4030);
and U5340 (N_5340,N_4706,N_3886);
nand U5341 (N_5341,N_2828,N_4223);
and U5342 (N_5342,N_4052,N_3111);
xor U5343 (N_5343,N_2942,N_4326);
and U5344 (N_5344,N_3206,N_4921);
nand U5345 (N_5345,N_4559,N_3091);
xor U5346 (N_5346,N_3702,N_4546);
or U5347 (N_5347,N_4355,N_4578);
and U5348 (N_5348,N_4245,N_4704);
xor U5349 (N_5349,N_4100,N_4656);
nor U5350 (N_5350,N_4022,N_3877);
or U5351 (N_5351,N_3949,N_4673);
and U5352 (N_5352,N_4491,N_3493);
and U5353 (N_5353,N_2547,N_2952);
nand U5354 (N_5354,N_4919,N_3609);
nand U5355 (N_5355,N_3017,N_3429);
or U5356 (N_5356,N_2790,N_3313);
nor U5357 (N_5357,N_4093,N_2700);
nand U5358 (N_5358,N_3275,N_3435);
xnor U5359 (N_5359,N_4931,N_4514);
nand U5360 (N_5360,N_3019,N_2832);
or U5361 (N_5361,N_2653,N_3177);
nor U5362 (N_5362,N_4498,N_3786);
and U5363 (N_5363,N_2744,N_3281);
and U5364 (N_5364,N_3613,N_4340);
nand U5365 (N_5365,N_3060,N_3363);
nand U5366 (N_5366,N_3816,N_2789);
or U5367 (N_5367,N_4914,N_2533);
or U5368 (N_5368,N_4110,N_3403);
xnor U5369 (N_5369,N_4810,N_4214);
nor U5370 (N_5370,N_4750,N_3896);
nor U5371 (N_5371,N_3933,N_2518);
xor U5372 (N_5372,N_4346,N_2599);
or U5373 (N_5373,N_2684,N_2831);
nor U5374 (N_5374,N_3149,N_3619);
or U5375 (N_5375,N_4998,N_4728);
or U5376 (N_5376,N_3143,N_3827);
nand U5377 (N_5377,N_2805,N_4067);
and U5378 (N_5378,N_3236,N_3798);
nand U5379 (N_5379,N_3272,N_3904);
xnor U5380 (N_5380,N_4385,N_4682);
and U5381 (N_5381,N_3287,N_2937);
nand U5382 (N_5382,N_2893,N_3531);
xor U5383 (N_5383,N_3324,N_3179);
or U5384 (N_5384,N_4054,N_4349);
nand U5385 (N_5385,N_3001,N_4642);
nand U5386 (N_5386,N_4463,N_4935);
xor U5387 (N_5387,N_3130,N_4391);
or U5388 (N_5388,N_3424,N_4905);
or U5389 (N_5389,N_3516,N_4250);
nor U5390 (N_5390,N_3158,N_4623);
and U5391 (N_5391,N_3561,N_3290);
nand U5392 (N_5392,N_2774,N_2796);
xnor U5393 (N_5393,N_2777,N_2746);
and U5394 (N_5394,N_4829,N_4499);
nand U5395 (N_5395,N_4136,N_4814);
and U5396 (N_5396,N_3165,N_4146);
nand U5397 (N_5397,N_3854,N_4676);
xnor U5398 (N_5398,N_3871,N_4583);
xor U5399 (N_5399,N_4123,N_4086);
and U5400 (N_5400,N_2636,N_4257);
nor U5401 (N_5401,N_4244,N_3559);
nor U5402 (N_5402,N_4833,N_2680);
xor U5403 (N_5403,N_4065,N_3229);
nor U5404 (N_5404,N_4882,N_3045);
nor U5405 (N_5405,N_3658,N_4772);
nor U5406 (N_5406,N_3105,N_4639);
or U5407 (N_5407,N_4331,N_3335);
nand U5408 (N_5408,N_4868,N_3161);
and U5409 (N_5409,N_3164,N_4577);
xnor U5410 (N_5410,N_2609,N_3321);
xnor U5411 (N_5411,N_4104,N_4677);
nor U5412 (N_5412,N_3527,N_4449);
xnor U5413 (N_5413,N_4778,N_3127);
and U5414 (N_5414,N_4519,N_2598);
nor U5415 (N_5415,N_3732,N_4847);
and U5416 (N_5416,N_4345,N_2644);
or U5417 (N_5417,N_4297,N_4012);
nor U5418 (N_5418,N_2813,N_3978);
xnor U5419 (N_5419,N_4819,N_4525);
xor U5420 (N_5420,N_3571,N_4967);
nand U5421 (N_5421,N_3232,N_4694);
or U5422 (N_5422,N_3172,N_4816);
or U5423 (N_5423,N_3944,N_4070);
or U5424 (N_5424,N_4304,N_3973);
xnor U5425 (N_5425,N_2532,N_3217);
xor U5426 (N_5426,N_2600,N_4109);
and U5427 (N_5427,N_3818,N_3241);
and U5428 (N_5428,N_3012,N_4007);
or U5429 (N_5429,N_2579,N_3928);
xor U5430 (N_5430,N_4942,N_2522);
xnor U5431 (N_5431,N_4528,N_2503);
or U5432 (N_5432,N_3740,N_3692);
nor U5433 (N_5433,N_4506,N_2914);
or U5434 (N_5434,N_4764,N_4835);
xor U5435 (N_5435,N_4132,N_3142);
nand U5436 (N_5436,N_4429,N_4063);
nand U5437 (N_5437,N_2853,N_3826);
xnor U5438 (N_5438,N_4066,N_3430);
or U5439 (N_5439,N_2575,N_4264);
or U5440 (N_5440,N_2939,N_3899);
nand U5441 (N_5441,N_3337,N_3885);
xor U5442 (N_5442,N_4853,N_3739);
or U5443 (N_5443,N_3914,N_3067);
nand U5444 (N_5444,N_4679,N_4376);
nand U5445 (N_5445,N_3560,N_3592);
nor U5446 (N_5446,N_3301,N_3152);
nor U5447 (N_5447,N_3409,N_3952);
xor U5448 (N_5448,N_2908,N_3646);
or U5449 (N_5449,N_3053,N_3100);
and U5450 (N_5450,N_3256,N_3544);
xor U5451 (N_5451,N_4806,N_3418);
or U5452 (N_5452,N_3097,N_3009);
xor U5453 (N_5453,N_2620,N_3339);
or U5454 (N_5454,N_4462,N_4549);
or U5455 (N_5455,N_2814,N_3372);
or U5456 (N_5456,N_3522,N_2505);
nand U5457 (N_5457,N_2658,N_3906);
or U5458 (N_5458,N_3329,N_3543);
or U5459 (N_5459,N_3864,N_2651);
and U5460 (N_5460,N_3166,N_2755);
and U5461 (N_5461,N_3911,N_4943);
nor U5462 (N_5462,N_3190,N_4576);
nand U5463 (N_5463,N_3467,N_4968);
nor U5464 (N_5464,N_3681,N_4051);
nor U5465 (N_5465,N_4773,N_3630);
or U5466 (N_5466,N_3147,N_4267);
nor U5467 (N_5467,N_4153,N_4205);
nand U5468 (N_5468,N_3364,N_4570);
nand U5469 (N_5469,N_4461,N_2923);
nand U5470 (N_5470,N_4072,N_2770);
xnor U5471 (N_5471,N_2730,N_2637);
nor U5472 (N_5472,N_4489,N_4402);
nor U5473 (N_5473,N_4950,N_3246);
or U5474 (N_5474,N_2557,N_4482);
and U5475 (N_5475,N_4831,N_2685);
xnor U5476 (N_5476,N_4464,N_3723);
xor U5477 (N_5477,N_3122,N_3767);
or U5478 (N_5478,N_4097,N_3266);
and U5479 (N_5479,N_4226,N_2634);
nor U5480 (N_5480,N_3868,N_2516);
and U5481 (N_5481,N_3862,N_2551);
and U5482 (N_5482,N_2915,N_4509);
nand U5483 (N_5483,N_4796,N_3425);
nor U5484 (N_5484,N_2882,N_3170);
xor U5485 (N_5485,N_3349,N_3299);
nand U5486 (N_5486,N_2845,N_4011);
nand U5487 (N_5487,N_3201,N_2822);
or U5488 (N_5488,N_2643,N_3220);
xnor U5489 (N_5489,N_3833,N_4069);
xnor U5490 (N_5490,N_3205,N_4434);
nor U5491 (N_5491,N_4280,N_4081);
nor U5492 (N_5492,N_3006,N_3184);
or U5493 (N_5493,N_2968,N_4405);
xnor U5494 (N_5494,N_2712,N_2703);
and U5495 (N_5495,N_4717,N_3772);
or U5496 (N_5496,N_4889,N_4367);
xor U5497 (N_5497,N_2606,N_2699);
nand U5498 (N_5498,N_4422,N_3262);
nor U5499 (N_5499,N_4203,N_3937);
nand U5500 (N_5500,N_3744,N_2670);
and U5501 (N_5501,N_3007,N_3089);
nor U5502 (N_5502,N_2611,N_4649);
and U5503 (N_5503,N_3389,N_4352);
or U5504 (N_5504,N_4844,N_4880);
xnor U5505 (N_5505,N_2602,N_4374);
nor U5506 (N_5506,N_3987,N_4903);
or U5507 (N_5507,N_4419,N_4332);
nor U5508 (N_5508,N_4055,N_3700);
nand U5509 (N_5509,N_3243,N_2558);
nand U5510 (N_5510,N_3315,N_2862);
xnor U5511 (N_5511,N_4972,N_3589);
nand U5512 (N_5512,N_3647,N_3542);
or U5513 (N_5513,N_3698,N_4392);
and U5514 (N_5514,N_4418,N_4933);
or U5515 (N_5515,N_4939,N_2713);
nand U5516 (N_5516,N_3665,N_3140);
and U5517 (N_5517,N_4420,N_2521);
nand U5518 (N_5518,N_4554,N_4133);
nand U5519 (N_5519,N_2578,N_4397);
and U5520 (N_5520,N_4435,N_3655);
xor U5521 (N_5521,N_3133,N_2612);
xnor U5522 (N_5522,N_3411,N_3283);
or U5523 (N_5523,N_4440,N_4295);
nor U5524 (N_5524,N_2879,N_3274);
nor U5525 (N_5525,N_3764,N_3661);
nand U5526 (N_5526,N_3196,N_4144);
xnor U5527 (N_5527,N_2552,N_3472);
and U5528 (N_5528,N_3135,N_4729);
or U5529 (N_5529,N_4892,N_4019);
nor U5530 (N_5530,N_4873,N_4233);
nand U5531 (N_5531,N_4314,N_4206);
nor U5532 (N_5532,N_4928,N_3792);
nand U5533 (N_5533,N_3422,N_2671);
xnor U5534 (N_5534,N_4142,N_3368);
nand U5535 (N_5535,N_4163,N_4792);
nand U5536 (N_5536,N_4099,N_2660);
xor U5537 (N_5537,N_3838,N_2645);
nor U5538 (N_5538,N_3612,N_4259);
nand U5539 (N_5539,N_3395,N_2970);
xor U5540 (N_5540,N_2659,N_3226);
nor U5541 (N_5541,N_3618,N_4960);
and U5542 (N_5542,N_4542,N_2706);
nor U5543 (N_5543,N_3876,N_4763);
xnor U5544 (N_5544,N_3342,N_3104);
xnor U5545 (N_5545,N_4130,N_4411);
nand U5546 (N_5546,N_3841,N_3114);
xor U5547 (N_5547,N_2872,N_2704);
or U5548 (N_5548,N_3955,N_4755);
xnor U5549 (N_5549,N_2631,N_2534);
or U5550 (N_5550,N_4645,N_3541);
nor U5551 (N_5551,N_4700,N_2812);
and U5552 (N_5552,N_4446,N_3080);
nor U5553 (N_5553,N_3320,N_2595);
xor U5554 (N_5554,N_2556,N_3509);
nand U5555 (N_5555,N_2873,N_2691);
or U5556 (N_5556,N_3822,N_3920);
nand U5557 (N_5557,N_4186,N_2642);
or U5558 (N_5558,N_2993,N_3651);
and U5559 (N_5559,N_4386,N_4539);
or U5560 (N_5560,N_4954,N_3981);
xnor U5561 (N_5561,N_3672,N_3432);
or U5562 (N_5562,N_4860,N_3461);
nand U5563 (N_5563,N_4629,N_3054);
xor U5564 (N_5564,N_4917,N_4116);
or U5565 (N_5565,N_2840,N_4053);
and U5566 (N_5566,N_3980,N_4848);
and U5567 (N_5567,N_4472,N_2918);
nand U5568 (N_5568,N_3622,N_4474);
xor U5569 (N_5569,N_3709,N_2911);
or U5570 (N_5570,N_3861,N_3293);
and U5571 (N_5571,N_3352,N_4278);
nand U5572 (N_5572,N_3092,N_3345);
nor U5573 (N_5573,N_2994,N_3800);
nand U5574 (N_5574,N_4329,N_2948);
nor U5575 (N_5575,N_3401,N_3793);
and U5576 (N_5576,N_3898,N_4958);
nand U5577 (N_5577,N_2925,N_3599);
xnor U5578 (N_5578,N_3610,N_2701);
nor U5579 (N_5579,N_3947,N_2708);
nand U5580 (N_5580,N_4713,N_4584);
or U5581 (N_5581,N_3381,N_3062);
nor U5582 (N_5582,N_4333,N_2775);
and U5583 (N_5583,N_2621,N_4650);
nor U5584 (N_5584,N_4373,N_2960);
and U5585 (N_5585,N_3346,N_3549);
nor U5586 (N_5586,N_2849,N_4803);
nand U5587 (N_5587,N_3420,N_4992);
and U5588 (N_5588,N_3308,N_4454);
and U5589 (N_5589,N_2892,N_2661);
nor U5590 (N_5590,N_3197,N_3757);
and U5591 (N_5591,N_3712,N_2953);
or U5592 (N_5592,N_3617,N_3551);
xnor U5593 (N_5593,N_3225,N_3428);
nand U5594 (N_5594,N_2766,N_4279);
nand U5595 (N_5595,N_4361,N_3124);
nand U5596 (N_5596,N_3374,N_4228);
nor U5597 (N_5597,N_3369,N_4601);
nor U5598 (N_5598,N_3696,N_2586);
and U5599 (N_5599,N_3371,N_4299);
nand U5600 (N_5600,N_4746,N_2517);
nand U5601 (N_5601,N_2679,N_3362);
nor U5602 (N_5602,N_3835,N_3572);
or U5603 (N_5603,N_2523,N_4018);
nor U5604 (N_5604,N_4736,N_4247);
and U5605 (N_5605,N_2767,N_3866);
nand U5606 (N_5606,N_2977,N_3901);
and U5607 (N_5607,N_4157,N_3968);
and U5608 (N_5608,N_4956,N_3780);
nor U5609 (N_5609,N_2682,N_2692);
and U5610 (N_5610,N_3603,N_2698);
and U5611 (N_5611,N_3511,N_4199);
nand U5612 (N_5612,N_3332,N_3088);
xnor U5613 (N_5613,N_4651,N_3471);
nor U5614 (N_5614,N_3050,N_3126);
nand U5615 (N_5615,N_3873,N_3652);
xor U5616 (N_5616,N_2824,N_4353);
xnor U5617 (N_5617,N_3227,N_4404);
and U5618 (N_5618,N_4155,N_4515);
xnor U5619 (N_5619,N_4310,N_3155);
nand U5620 (N_5620,N_4837,N_2583);
and U5621 (N_5621,N_4592,N_4895);
nand U5622 (N_5622,N_2635,N_4851);
nor U5623 (N_5623,N_2962,N_3528);
or U5624 (N_5624,N_4354,N_2927);
or U5625 (N_5625,N_4964,N_3446);
or U5626 (N_5626,N_2916,N_4246);
and U5627 (N_5627,N_4957,N_3162);
xor U5628 (N_5628,N_4013,N_3951);
nor U5629 (N_5629,N_3358,N_3726);
nand U5630 (N_5630,N_3918,N_3081);
nand U5631 (N_5631,N_4769,N_4535);
nor U5632 (N_5632,N_4721,N_3021);
or U5633 (N_5633,N_3300,N_4274);
or U5634 (N_5634,N_4216,N_4530);
xnor U5635 (N_5635,N_4202,N_3693);
xnor U5636 (N_5636,N_2854,N_3529);
nor U5637 (N_5637,N_3284,N_3799);
xor U5638 (N_5638,N_3878,N_4125);
or U5639 (N_5639,N_3341,N_2861);
and U5640 (N_5640,N_3643,N_3116);
or U5641 (N_5641,N_3602,N_3344);
nor U5642 (N_5642,N_4709,N_4581);
xnor U5643 (N_5643,N_3996,N_4365);
and U5644 (N_5644,N_4510,N_4823);
xor U5645 (N_5645,N_4653,N_4734);
or U5646 (N_5646,N_3986,N_3688);
or U5647 (N_5647,N_2569,N_3074);
nor U5648 (N_5648,N_4487,N_3642);
or U5649 (N_5649,N_3526,N_2565);
nor U5650 (N_5650,N_3365,N_4395);
nor U5651 (N_5651,N_4907,N_4316);
nand U5652 (N_5652,N_3191,N_4809);
nor U5653 (N_5653,N_2971,N_4512);
nor U5654 (N_5654,N_4023,N_4605);
nor U5655 (N_5655,N_4558,N_4522);
xor U5656 (N_5656,N_3624,N_3831);
xnor U5657 (N_5657,N_3905,N_4061);
nand U5658 (N_5658,N_3066,N_3052);
or U5659 (N_5659,N_3055,N_4049);
nand U5660 (N_5660,N_4170,N_3436);
or U5661 (N_5661,N_3473,N_3832);
or U5662 (N_5662,N_4818,N_4242);
or U5663 (N_5663,N_3093,N_3900);
or U5664 (N_5664,N_3514,N_2654);
nand U5665 (N_5665,N_3347,N_4309);
and U5666 (N_5666,N_4985,N_2815);
or U5667 (N_5667,N_3722,N_4300);
or U5668 (N_5668,N_4469,N_2929);
nand U5669 (N_5669,N_3061,N_2647);
nand U5670 (N_5670,N_2603,N_3476);
xnor U5671 (N_5671,N_3210,N_4253);
nand U5672 (N_5672,N_2745,N_3212);
or U5673 (N_5673,N_3043,N_4562);
nor U5674 (N_5674,N_2593,N_4628);
and U5675 (N_5675,N_4808,N_3759);
nand U5676 (N_5676,N_2662,N_4249);
nor U5677 (N_5677,N_2829,N_4290);
xor U5678 (N_5678,N_2984,N_4641);
and U5679 (N_5679,N_4161,N_2587);
nor U5680 (N_5680,N_2958,N_4488);
nor U5681 (N_5681,N_3355,N_4749);
nand U5682 (N_5682,N_2715,N_4003);
xnor U5683 (N_5683,N_4881,N_3847);
and U5684 (N_5684,N_4824,N_4618);
and U5685 (N_5685,N_2633,N_2592);
nand U5686 (N_5686,N_4204,N_4767);
or U5687 (N_5687,N_2806,N_4478);
nand U5688 (N_5688,N_3390,N_4636);
nand U5689 (N_5689,N_3863,N_4741);
xnor U5690 (N_5690,N_4553,N_2664);
and U5691 (N_5691,N_4322,N_4431);
xor U5692 (N_5692,N_4467,N_4801);
nor U5693 (N_5693,N_4619,N_3044);
nor U5694 (N_5694,N_3462,N_3517);
nor U5695 (N_5695,N_3296,N_3228);
nand U5696 (N_5696,N_3431,N_3747);
and U5697 (N_5697,N_3778,N_4428);
nand U5698 (N_5698,N_2535,N_3682);
and U5699 (N_5699,N_4617,N_3265);
nand U5700 (N_5700,N_3851,N_4567);
nor U5701 (N_5701,N_3770,N_3223);
or U5702 (N_5702,N_3846,N_3508);
nand U5703 (N_5703,N_3405,N_3957);
nor U5704 (N_5704,N_2783,N_4164);
nor U5705 (N_5705,N_3632,N_2826);
or U5706 (N_5706,N_2843,N_4311);
xnor U5707 (N_5707,N_3557,N_2975);
nor U5708 (N_5708,N_4215,N_2545);
nor U5709 (N_5709,N_3525,N_4243);
nand U5710 (N_5710,N_3282,N_4308);
xor U5711 (N_5711,N_3797,N_4870);
xnor U5712 (N_5712,N_4323,N_4557);
xor U5713 (N_5713,N_4504,N_2864);
nor U5714 (N_5714,N_3134,N_3171);
nand U5715 (N_5715,N_2509,N_2784);
and U5716 (N_5716,N_2904,N_4846);
and U5717 (N_5717,N_2607,N_2999);
nor U5718 (N_5718,N_4427,N_3805);
and U5719 (N_5719,N_4248,N_3416);
nand U5720 (N_5720,N_3558,N_4887);
nand U5721 (N_5721,N_2865,N_3098);
nor U5722 (N_5722,N_3038,N_4568);
nand U5723 (N_5723,N_4534,N_3388);
xor U5724 (N_5724,N_4565,N_3762);
or U5725 (N_5725,N_3322,N_4057);
nor U5726 (N_5726,N_2897,N_3897);
or U5727 (N_5727,N_4115,N_3608);
nand U5728 (N_5728,N_3639,N_4716);
nand U5729 (N_5729,N_2624,N_3984);
nor U5730 (N_5730,N_4432,N_4976);
nor U5731 (N_5731,N_4258,N_2738);
nand U5732 (N_5732,N_4439,N_2669);
nand U5733 (N_5733,N_3844,N_3453);
nand U5734 (N_5734,N_3504,N_4667);
and U5735 (N_5735,N_2648,N_4731);
nor U5736 (N_5736,N_3953,N_4227);
nand U5737 (N_5737,N_4183,N_2943);
or U5738 (N_5738,N_4254,N_3929);
or U5739 (N_5739,N_4221,N_3465);
nor U5740 (N_5740,N_3994,N_3568);
xor U5741 (N_5741,N_3434,N_2563);
or U5742 (N_5742,N_3340,N_4009);
or U5743 (N_5743,N_2763,N_4370);
nand U5744 (N_5744,N_4595,N_2895);
and U5745 (N_5745,N_2794,N_3580);
nor U5746 (N_5746,N_4875,N_4771);
or U5747 (N_5747,N_4301,N_3552);
xnor U5748 (N_5748,N_4707,N_2526);
and U5749 (N_5749,N_3451,N_4701);
nor U5750 (N_5750,N_2760,N_3922);
nand U5751 (N_5751,N_3574,N_3760);
or U5752 (N_5752,N_4680,N_4735);
and U5753 (N_5753,N_4408,N_2696);
xnor U5754 (N_5754,N_4500,N_4043);
nand U5755 (N_5755,N_3880,N_4720);
and U5756 (N_5756,N_3721,N_2728);
or U5757 (N_5757,N_3178,N_4955);
and U5758 (N_5758,N_3271,N_3578);
nand U5759 (N_5759,N_4497,N_4091);
or U5760 (N_5760,N_3950,N_3917);
and U5761 (N_5761,N_4648,N_4952);
nor U5762 (N_5762,N_4897,N_3515);
and U5763 (N_5763,N_4229,N_3536);
or U5764 (N_5764,N_3959,N_3013);
xor U5765 (N_5765,N_3971,N_4635);
and U5766 (N_5766,N_3289,N_4869);
xnor U5767 (N_5767,N_2887,N_3594);
and U5768 (N_5768,N_3524,N_3817);
nand U5769 (N_5769,N_2905,N_2617);
nand U5770 (N_5770,N_3298,N_4647);
nor U5771 (N_5771,N_4366,N_4318);
xnor U5772 (N_5772,N_3343,N_4493);
xor U5773 (N_5773,N_3776,N_4521);
or U5774 (N_5774,N_4878,N_2921);
nand U5775 (N_5775,N_3998,N_3742);
and U5776 (N_5776,N_4027,N_4445);
nor U5777 (N_5777,N_4150,N_4783);
nor U5778 (N_5778,N_2809,N_3361);
or U5779 (N_5779,N_3648,N_4784);
and U5780 (N_5780,N_3292,N_4126);
xor U5781 (N_5781,N_4582,N_2980);
nand U5782 (N_5782,N_3005,N_4321);
and U5783 (N_5783,N_4965,N_4073);
nand U5784 (N_5784,N_2934,N_4184);
and U5785 (N_5785,N_3958,N_2779);
nand U5786 (N_5786,N_4286,N_4140);
or U5787 (N_5787,N_3521,N_4149);
nor U5788 (N_5788,N_4997,N_4158);
xor U5789 (N_5789,N_2716,N_4193);
or U5790 (N_5790,N_4688,N_2726);
and U5791 (N_5791,N_3437,N_3026);
and U5792 (N_5792,N_3316,N_4447);
and U5793 (N_5793,N_3753,N_3028);
xor U5794 (N_5794,N_2559,N_4762);
xnor U5795 (N_5795,N_4425,N_4890);
and U5796 (N_5796,N_4390,N_2564);
nand U5797 (N_5797,N_4363,N_3720);
nand U5798 (N_5798,N_3507,N_4798);
xnor U5799 (N_5799,N_4293,N_4961);
nand U5800 (N_5800,N_3255,N_4987);
nand U5801 (N_5801,N_2758,N_3478);
and U5802 (N_5802,N_4516,N_2632);
or U5803 (N_5803,N_2571,N_3829);
nand U5804 (N_5804,N_3537,N_3189);
nor U5805 (N_5805,N_3668,N_3806);
nand U5806 (N_5806,N_2537,N_4765);
and U5807 (N_5807,N_3221,N_3479);
xnor U5808 (N_5808,N_4944,N_4490);
nor U5809 (N_5809,N_2525,N_4160);
nor U5810 (N_5810,N_3010,N_4224);
nand U5811 (N_5811,N_4302,N_3510);
nor U5812 (N_5812,N_3782,N_2683);
or U5813 (N_5813,N_4443,N_4624);
or U5814 (N_5814,N_4426,N_3443);
or U5815 (N_5815,N_3106,N_2990);
and U5816 (N_5816,N_3120,N_4859);
and U5817 (N_5817,N_3889,N_2714);
nor U5818 (N_5818,N_4782,N_2674);
and U5819 (N_5819,N_2922,N_3231);
and U5820 (N_5820,N_3311,N_2649);
and U5821 (N_5821,N_3699,N_3059);
xnor U5822 (N_5822,N_4285,N_4182);
xor U5823 (N_5823,N_3943,N_4752);
nor U5824 (N_5824,N_4609,N_4953);
nand U5825 (N_5825,N_3588,N_3498);
xor U5826 (N_5826,N_3819,N_3969);
and U5827 (N_5827,N_2989,N_2742);
nor U5828 (N_5828,N_4638,N_4560);
or U5829 (N_5829,N_3491,N_3125);
nor U5830 (N_5830,N_3751,N_4858);
nor U5831 (N_5831,N_4235,N_3741);
nand U5832 (N_5832,N_4747,N_4232);
or U5833 (N_5833,N_3278,N_4387);
or U5834 (N_5834,N_4077,N_4962);
and U5835 (N_5835,N_3596,N_3049);
nor U5836 (N_5836,N_3173,N_3884);
nor U5837 (N_5837,N_3519,N_2870);
nand U5838 (N_5838,N_2963,N_2678);
nand U5839 (N_5839,N_4857,N_3995);
nand U5840 (N_5840,N_3586,N_3314);
nor U5841 (N_5841,N_4372,N_2538);
or U5842 (N_5842,N_4324,N_3769);
nand U5843 (N_5843,N_3200,N_3148);
nor U5844 (N_5844,N_4973,N_2816);
nor U5845 (N_5845,N_4872,N_4433);
and U5846 (N_5846,N_2998,N_4805);
nand U5847 (N_5847,N_4759,N_4038);
or U5848 (N_5848,N_4171,N_2567);
nand U5849 (N_5849,N_4477,N_4689);
nor U5850 (N_5850,N_4966,N_4655);
or U5851 (N_5851,N_4633,N_3083);
or U5852 (N_5852,N_3883,N_4866);
or U5853 (N_5853,N_3530,N_4665);
nand U5854 (N_5854,N_4255,N_3366);
nor U5855 (N_5855,N_2687,N_3611);
xnor U5856 (N_5856,N_4839,N_4599);
and U5857 (N_5857,N_4090,N_4359);
or U5858 (N_5858,N_4615,N_4999);
or U5859 (N_5859,N_4794,N_2898);
or U5860 (N_5860,N_3667,N_2776);
nor U5861 (N_5861,N_4384,N_3319);
xor U5862 (N_5862,N_4748,N_4369);
nand U5863 (N_5863,N_2729,N_3198);
and U5864 (N_5864,N_3303,N_4368);
xnor U5865 (N_5865,N_3791,N_3208);
nor U5866 (N_5866,N_4982,N_3020);
nand U5867 (N_5867,N_3396,N_3677);
and U5868 (N_5868,N_4843,N_3318);
nor U5869 (N_5869,N_3890,N_2519);
or U5870 (N_5870,N_3684,N_3752);
xor U5871 (N_5871,N_4117,N_4312);
nor U5872 (N_5872,N_2752,N_3724);
and U5873 (N_5873,N_3348,N_2737);
xor U5874 (N_5874,N_3992,N_3777);
or U5875 (N_5875,N_3399,N_4652);
xnor U5876 (N_5876,N_3781,N_4527);
and U5877 (N_5877,N_4698,N_3350);
and U5878 (N_5878,N_4177,N_4507);
nand U5879 (N_5879,N_3455,N_4561);
and U5880 (N_5880,N_3121,N_2590);
xor U5881 (N_5881,N_3912,N_3705);
nor U5882 (N_5882,N_2912,N_2983);
or U5883 (N_5883,N_3494,N_3439);
and U5884 (N_5884,N_2718,N_3930);
and U5885 (N_5885,N_4690,N_3076);
nor U5886 (N_5886,N_2857,N_4062);
nor U5887 (N_5887,N_3484,N_3025);
nand U5888 (N_5888,N_4564,N_3977);
or U5889 (N_5889,N_4508,N_4451);
or U5890 (N_5890,N_3482,N_3983);
nand U5891 (N_5891,N_3583,N_4978);
or U5892 (N_5892,N_4448,N_3621);
nand U5893 (N_5893,N_2585,N_2773);
xor U5894 (N_5894,N_4219,N_4356);
or U5895 (N_5895,N_2615,N_4563);
xnor U5896 (N_5896,N_3354,N_2666);
xnor U5897 (N_5897,N_2597,N_3414);
or U5898 (N_5898,N_2562,N_3872);
nand U5899 (N_5899,N_4167,N_2810);
or U5900 (N_5900,N_3860,N_3295);
xor U5901 (N_5901,N_3297,N_3662);
and U5902 (N_5902,N_4025,N_2778);
xor U5903 (N_5903,N_3756,N_4087);
xnor U5904 (N_5904,N_4867,N_3926);
nor U5905 (N_5905,N_2988,N_2967);
or U5906 (N_5906,N_4131,N_4757);
nor U5907 (N_5907,N_3402,N_3391);
nand U5908 (N_5908,N_3701,N_4526);
and U5909 (N_5909,N_4327,N_4785);
or U5910 (N_5910,N_3310,N_3469);
or U5911 (N_5911,N_4948,N_4174);
or U5912 (N_5912,N_4337,N_3064);
nand U5913 (N_5913,N_3470,N_2504);
or U5914 (N_5914,N_3024,N_4415);
nor U5915 (N_5915,N_2549,N_4502);
nand U5916 (N_5916,N_4825,N_3734);
xor U5917 (N_5917,N_3500,N_3940);
and U5918 (N_5918,N_4724,N_3036);
xnor U5919 (N_5919,N_2610,N_3417);
and U5920 (N_5920,N_4523,N_3441);
or U5921 (N_5921,N_3252,N_4151);
xnor U5922 (N_5922,N_3022,N_4064);
nand U5923 (N_5923,N_3582,N_3326);
or U5924 (N_5924,N_4524,N_4517);
and U5925 (N_5925,N_3030,N_3202);
nand U5926 (N_5926,N_3357,N_4002);
and U5927 (N_5927,N_3069,N_3393);
and U5928 (N_5928,N_3280,N_3570);
nor U5929 (N_5929,N_4237,N_2855);
nor U5930 (N_5930,N_4212,N_3307);
or U5931 (N_5931,N_3285,N_4453);
nand U5932 (N_5932,N_2717,N_2795);
nand U5933 (N_5933,N_2981,N_3168);
nand U5934 (N_5934,N_3710,N_3187);
xnor U5935 (N_5935,N_4811,N_4417);
xnor U5936 (N_5936,N_4217,N_3499);
or U5937 (N_5937,N_4685,N_4513);
nand U5938 (N_5938,N_2623,N_3188);
and U5939 (N_5939,N_2693,N_3997);
xor U5940 (N_5940,N_3546,N_3532);
xnor U5941 (N_5941,N_4543,N_3139);
and U5942 (N_5942,N_3204,N_4864);
nand U5943 (N_5943,N_3909,N_3616);
and U5944 (N_5944,N_4885,N_4006);
nor U5945 (N_5945,N_3468,N_4172);
nor U5946 (N_5946,N_3261,N_3654);
xnor U5947 (N_5947,N_4602,N_4139);
or U5948 (N_5948,N_3153,N_2686);
nand U5949 (N_5949,N_3244,N_2875);
nor U5950 (N_5950,N_4675,N_4621);
nand U5951 (N_5951,N_4014,N_3808);
nand U5952 (N_5952,N_4378,N_3814);
or U5953 (N_5953,N_4909,N_3902);
nor U5954 (N_5954,N_3338,N_2743);
nand U5955 (N_5955,N_2553,N_2764);
or U5956 (N_5956,N_3730,N_2665);
and U5957 (N_5957,N_2835,N_3264);
xor U5958 (N_5958,N_3946,N_3356);
xnor U5959 (N_5959,N_4899,N_3839);
or U5960 (N_5960,N_3567,N_4820);
nand U5961 (N_5961,N_2581,N_2842);
and U5962 (N_5962,N_3645,N_4908);
nor U5963 (N_5963,N_4056,N_2901);
xor U5964 (N_5964,N_3795,N_4358);
nand U5965 (N_5965,N_4252,N_4127);
or U5966 (N_5966,N_3919,N_2751);
xnor U5967 (N_5967,N_3008,N_3761);
and U5968 (N_5968,N_3605,N_4579);
xor U5969 (N_5969,N_4141,N_4551);
or U5970 (N_5970,N_3160,N_3132);
or U5971 (N_5971,N_2688,N_4041);
xnor U5972 (N_5972,N_2677,N_4616);
nand U5973 (N_5973,N_4485,N_4977);
nor U5974 (N_5974,N_4990,N_3410);
or U5975 (N_5975,N_3327,N_3385);
and U5976 (N_5976,N_4268,N_3512);
nor U5977 (N_5977,N_4886,N_2511);
nor U5978 (N_5978,N_4260,N_4173);
or U5979 (N_5979,N_4034,N_3915);
and U5980 (N_5980,N_2919,N_3131);
and U5981 (N_5981,N_2673,N_3614);
and U5982 (N_5982,N_3392,N_2965);
and U5983 (N_5983,N_2851,N_4501);
and U5984 (N_5984,N_3117,N_3438);
and U5985 (N_5985,N_4821,N_4912);
nor U5986 (N_5986,N_4711,N_4970);
xor U5987 (N_5987,N_4024,N_3386);
nand U5988 (N_5988,N_2910,N_3931);
nand U5989 (N_5989,N_4084,N_4983);
and U5990 (N_5990,N_4470,N_4101);
nor U5991 (N_5991,N_2982,N_4234);
nor U5992 (N_5992,N_4923,N_2850);
or U5993 (N_5993,N_3691,N_4862);
xnor U5994 (N_5994,N_2513,N_4697);
and U5995 (N_5995,N_4703,N_4959);
and U5996 (N_5996,N_4668,N_3031);
and U5997 (N_5997,N_3708,N_2544);
nand U5998 (N_5998,N_3972,N_4608);
or U5999 (N_5999,N_3042,N_4319);
and U6000 (N_6000,N_2771,N_2830);
or U6001 (N_6001,N_3460,N_4571);
and U6002 (N_6002,N_4074,N_4936);
nand U6003 (N_6003,N_4220,N_4684);
xor U6004 (N_6004,N_3328,N_4714);
nor U6005 (N_6005,N_4288,N_3669);
and U6006 (N_6006,N_4336,N_4276);
nand U6007 (N_6007,N_3304,N_3211);
nor U6008 (N_6008,N_4305,N_3029);
xor U6009 (N_6009,N_3449,N_4708);
or U6010 (N_6010,N_3640,N_2886);
nor U6011 (N_6011,N_4465,N_2725);
or U6012 (N_6012,N_2640,N_2510);
nand U6013 (N_6013,N_2577,N_2866);
nor U6014 (N_6014,N_4994,N_4398);
xor U6015 (N_6015,N_3634,N_4348);
and U6016 (N_6016,N_4238,N_2724);
xnor U6017 (N_6017,N_4896,N_4768);
nand U6018 (N_6018,N_4790,N_3137);
xor U6019 (N_6019,N_2938,N_3413);
xor U6020 (N_6020,N_4596,N_4037);
xor U6021 (N_6021,N_4740,N_2756);
xor U6022 (N_6022,N_3535,N_3305);
or U6023 (N_6023,N_2512,N_3849);
xnor U6024 (N_6024,N_3533,N_2733);
and U6025 (N_6025,N_2626,N_3459);
nor U6026 (N_6026,N_3679,N_4989);
and U6027 (N_6027,N_3004,N_3445);
and U6028 (N_6028,N_3869,N_3359);
and U6029 (N_6029,N_4108,N_2869);
xor U6030 (N_6030,N_2874,N_4306);
nor U6031 (N_6031,N_4092,N_3270);
or U6032 (N_6032,N_4412,N_4883);
and U6033 (N_6033,N_2739,N_3181);
nand U6034 (N_6034,N_4538,N_3641);
xor U6035 (N_6035,N_3373,N_3895);
nand U6036 (N_6036,N_3240,N_4287);
nand U6037 (N_6037,N_2754,N_3843);
or U6038 (N_6038,N_4555,N_3887);
or U6039 (N_6039,N_4207,N_4910);
nor U6040 (N_6040,N_3859,N_4832);
or U6041 (N_6041,N_4458,N_3276);
nor U6042 (N_6042,N_2542,N_3807);
nor U6043 (N_6043,N_3623,N_4240);
and U6044 (N_6044,N_3487,N_4456);
nor U6045 (N_6045,N_3664,N_3234);
xnor U6046 (N_6046,N_3378,N_4379);
xnor U6047 (N_6047,N_4904,N_2539);
or U6048 (N_6048,N_2902,N_3213);
or U6049 (N_6049,N_2741,N_4545);
nand U6050 (N_6050,N_4981,N_2846);
nor U6051 (N_6051,N_2800,N_3695);
or U6052 (N_6052,N_3268,N_3383);
nor U6053 (N_6053,N_2639,N_3783);
nor U6054 (N_6054,N_3072,N_3407);
xnor U6055 (N_6055,N_3068,N_3892);
and U6056 (N_6056,N_4874,N_3291);
nor U6057 (N_6057,N_4654,N_3954);
xor U6058 (N_6058,N_3979,N_4401);
or U6059 (N_6059,N_2974,N_3492);
and U6060 (N_6060,N_3094,N_4725);
nor U6061 (N_6061,N_4607,N_4743);
nor U6062 (N_6062,N_3620,N_3581);
xor U6063 (N_6063,N_2848,N_3974);
or U6064 (N_6064,N_4884,N_3824);
and U6065 (N_6065,N_3483,N_4518);
nor U6066 (N_6066,N_3058,N_2821);
and U6067 (N_6067,N_4988,N_3856);
nor U6068 (N_6068,N_4421,N_3697);
and U6069 (N_6069,N_4325,N_3694);
or U6070 (N_6070,N_4993,N_2572);
and U6071 (N_6071,N_2881,N_4503);
nand U6072 (N_6072,N_3888,N_3387);
nand U6073 (N_6073,N_2798,N_4660);
nor U6074 (N_6074,N_3579,N_3218);
nor U6075 (N_6075,N_4926,N_4444);
or U6076 (N_6076,N_3048,N_4556);
or U6077 (N_6077,N_4505,N_2859);
xor U6078 (N_6078,N_4083,N_3785);
and U6079 (N_6079,N_3858,N_4922);
nand U6080 (N_6080,N_3230,N_2985);
xnor U6081 (N_6081,N_2949,N_4082);
xnor U6082 (N_6082,N_4927,N_2768);
and U6083 (N_6083,N_2992,N_4459);
or U6084 (N_6084,N_2710,N_4307);
xnor U6085 (N_6085,N_4218,N_3258);
and U6086 (N_6086,N_3649,N_2786);
xor U6087 (N_6087,N_3989,N_2588);
xnor U6088 (N_6088,N_3991,N_3923);
and U6089 (N_6089,N_4399,N_3353);
and U6090 (N_6090,N_2529,N_3834);
nand U6091 (N_6091,N_4597,N_2676);
nor U6092 (N_6092,N_4282,N_3351);
xor U6093 (N_6093,N_4042,N_3503);
nand U6094 (N_6094,N_3894,N_3215);
nor U6095 (N_6095,N_2734,N_4198);
and U6096 (N_6096,N_4980,N_3942);
or U6097 (N_6097,N_4113,N_3569);
xnor U6098 (N_6098,N_4855,N_2594);
or U6099 (N_6099,N_4079,N_4176);
nor U6100 (N_6100,N_2959,N_3380);
nor U6101 (N_6101,N_4342,N_4634);
and U6102 (N_6102,N_4166,N_3539);
or U6103 (N_6103,N_2837,N_4836);
and U6104 (N_6104,N_4574,N_4341);
xnor U6105 (N_6105,N_4230,N_3804);
nand U6106 (N_6106,N_4963,N_3071);
and U6107 (N_6107,N_2530,N_4103);
and U6108 (N_6108,N_3101,N_4442);
or U6109 (N_6109,N_2560,N_3433);
or U6110 (N_6110,N_4815,N_3836);
or U6111 (N_6111,N_3725,N_3003);
nand U6112 (N_6112,N_4380,N_3637);
nor U6113 (N_6113,N_3566,N_3186);
xnor U6114 (N_6114,N_4751,N_4272);
nor U6115 (N_6115,N_4211,N_3573);
or U6116 (N_6116,N_4712,N_4080);
and U6117 (N_6117,N_3746,N_3848);
nor U6118 (N_6118,N_2966,N_3963);
and U6119 (N_6119,N_3078,N_2932);
xor U6120 (N_6120,N_2652,N_3214);
nand U6121 (N_6121,N_4842,N_4145);
or U6122 (N_6122,N_3257,N_2589);
or U6123 (N_6123,N_4737,N_4334);
xor U6124 (N_6124,N_4406,N_3855);
nor U6125 (N_6125,N_3680,N_4360);
nand U6126 (N_6126,N_2820,N_4251);
nor U6127 (N_6127,N_3910,N_4657);
nor U6128 (N_6128,N_3690,N_4949);
or U6129 (N_6129,N_3676,N_2891);
xnor U6130 (N_6130,N_2888,N_2844);
xnor U6131 (N_6131,N_4486,N_3488);
or U6132 (N_6132,N_3018,N_3110);
xor U6133 (N_6133,N_4781,N_4550);
and U6134 (N_6134,N_4776,N_3597);
xor U6135 (N_6135,N_4479,N_3138);
xor U6136 (N_6136,N_2709,N_3082);
xor U6137 (N_6137,N_4128,N_2502);
or U6138 (N_6138,N_2996,N_4924);
nand U6139 (N_6139,N_3534,N_3235);
and U6140 (N_6140,N_2940,N_2627);
and U6141 (N_6141,N_2867,N_3595);
nand U6142 (N_6142,N_3219,N_3737);
nor U6143 (N_6143,N_2608,N_4068);
nor U6144 (N_6144,N_3675,N_4566);
nor U6145 (N_6145,N_2514,N_3156);
xnor U6146 (N_6146,N_2736,N_3689);
or U6147 (N_6147,N_3309,N_3852);
or U6148 (N_6148,N_2520,N_3144);
nand U6149 (N_6149,N_3590,N_4048);
nand U6150 (N_6150,N_4945,N_4789);
and U6151 (N_6151,N_3874,N_4622);
and U6152 (N_6152,N_2735,N_3370);
nand U6153 (N_6153,N_2950,N_3840);
or U6154 (N_6154,N_4898,N_2707);
nor U6155 (N_6155,N_3195,N_3051);
xor U6156 (N_6156,N_3245,N_3379);
xnor U6157 (N_6157,N_2697,N_4410);
nand U6158 (N_6158,N_2508,N_3673);
or U6159 (N_6159,N_4004,N_3812);
xnor U6160 (N_6160,N_4733,N_4189);
and U6161 (N_6161,N_3713,N_3985);
nand U6162 (N_6162,N_3463,N_2847);
and U6163 (N_6163,N_3547,N_2667);
nand U6164 (N_6164,N_3628,N_4466);
or U6165 (N_6165,N_3711,N_2753);
nand U6166 (N_6166,N_3754,N_4991);
and U6167 (N_6167,N_3941,N_2672);
xnor U6168 (N_6168,N_4102,N_4659);
xor U6169 (N_6169,N_4540,N_2987);
nand U6170 (N_6170,N_3163,N_3771);
xnor U6171 (N_6171,N_3404,N_3102);
and U6172 (N_6172,N_3423,N_3821);
or U6173 (N_6173,N_3294,N_3598);
and U6174 (N_6174,N_4941,N_2986);
and U6175 (N_6175,N_4403,N_2573);
or U6176 (N_6176,N_3865,N_4187);
xnor U6177 (N_6177,N_3936,N_2646);
nor U6178 (N_6178,N_2616,N_4722);
or U6179 (N_6179,N_4804,N_4760);
nand U6180 (N_6180,N_4154,N_3584);
xor U6181 (N_6181,N_4273,N_3999);
and U6182 (N_6182,N_4544,N_3960);
nand U6183 (N_6183,N_2917,N_4045);
and U6184 (N_6184,N_4201,N_2792);
and U6185 (N_6185,N_2515,N_3893);
nand U6186 (N_6186,N_2500,N_2570);
xor U6187 (N_6187,N_4662,N_3502);
xor U6188 (N_6188,N_4637,N_3115);
xor U6189 (N_6189,N_2650,N_3801);
xor U6190 (N_6190,N_2852,N_4614);
nor U6191 (N_6191,N_3538,N_4208);
nor U6192 (N_6192,N_3254,N_2991);
nor U6193 (N_6193,N_4339,N_4275);
and U6194 (N_6194,N_3412,N_3034);
xor U6195 (N_6195,N_4663,N_4593);
nand U6196 (N_6196,N_4861,N_2884);
and U6197 (N_6197,N_4180,N_4807);
or U6198 (N_6198,N_4241,N_4840);
or U6199 (N_6199,N_3935,N_3796);
nand U6200 (N_6200,N_2913,N_4413);
xor U6201 (N_6201,N_3360,N_4699);
nand U6202 (N_6202,N_3924,N_4900);
nor U6203 (N_6203,N_3207,N_2782);
nand U6204 (N_6204,N_3267,N_4600);
and U6205 (N_6205,N_4974,N_3766);
nor U6206 (N_6206,N_3881,N_4761);
nor U6207 (N_6207,N_3367,N_4588);
or U6208 (N_6208,N_3426,N_2793);
or U6209 (N_6209,N_3151,N_2945);
nor U6210 (N_6210,N_2727,N_3014);
and U6211 (N_6211,N_4643,N_2803);
or U6212 (N_6212,N_3176,N_4031);
and U6213 (N_6213,N_4455,N_4580);
or U6214 (N_6214,N_4121,N_3174);
nand U6215 (N_6215,N_4350,N_4573);
and U6216 (N_6216,N_2528,N_3916);
and U6217 (N_6217,N_3513,N_4586);
nor U6218 (N_6218,N_4210,N_4476);
xnor U6219 (N_6219,N_3450,N_4590);
or U6220 (N_6220,N_3128,N_3154);
xor U6221 (N_6221,N_3650,N_2941);
nand U6222 (N_6222,N_4626,N_2580);
nand U6223 (N_6223,N_2655,N_2802);
nand U6224 (N_6224,N_4263,N_4351);
and U6225 (N_6225,N_2947,N_4424);
or U6226 (N_6226,N_4795,N_3970);
xnor U6227 (N_6227,N_2765,N_4611);
nand U6228 (N_6228,N_3666,N_3850);
nand U6229 (N_6229,N_3288,N_4266);
xnor U6230 (N_6230,N_3506,N_4902);
nand U6231 (N_6231,N_2601,N_3755);
nand U6232 (N_6232,N_3728,N_2871);
nor U6233 (N_6233,N_3745,N_3961);
nor U6234 (N_6234,N_2748,N_3604);
nand U6235 (N_6235,N_4911,N_4481);
nor U6236 (N_6236,N_4495,N_3678);
nor U6237 (N_6237,N_3956,N_4047);
nor U6238 (N_6238,N_3738,N_4913);
xor U6239 (N_6239,N_2541,N_3377);
nor U6240 (N_6240,N_4185,N_4979);
nand U6241 (N_6241,N_3657,N_4738);
xnor U6242 (N_6242,N_4932,N_4393);
xnor U6243 (N_6243,N_4000,N_3136);
nor U6244 (N_6244,N_4669,N_2838);
nor U6245 (N_6245,N_3629,N_3748);
or U6246 (N_6246,N_2584,N_4625);
nand U6247 (N_6247,N_4400,N_2536);
xnor U6248 (N_6248,N_3548,N_4120);
nand U6249 (N_6249,N_3454,N_4906);
nand U6250 (N_6250,N_3416,N_3571);
or U6251 (N_6251,N_4384,N_4298);
nor U6252 (N_6252,N_3584,N_4775);
or U6253 (N_6253,N_3504,N_3883);
xor U6254 (N_6254,N_4070,N_3722);
xnor U6255 (N_6255,N_2639,N_3690);
or U6256 (N_6256,N_4218,N_4724);
or U6257 (N_6257,N_4763,N_3785);
and U6258 (N_6258,N_3839,N_2519);
nand U6259 (N_6259,N_4540,N_3585);
nor U6260 (N_6260,N_4895,N_2576);
nor U6261 (N_6261,N_2672,N_4845);
xor U6262 (N_6262,N_3054,N_4127);
nor U6263 (N_6263,N_4389,N_2581);
nand U6264 (N_6264,N_3543,N_4564);
nor U6265 (N_6265,N_2747,N_3544);
nand U6266 (N_6266,N_2984,N_4016);
nand U6267 (N_6267,N_4701,N_3657);
xnor U6268 (N_6268,N_2815,N_2880);
nor U6269 (N_6269,N_4163,N_2618);
or U6270 (N_6270,N_3953,N_3660);
xnor U6271 (N_6271,N_3373,N_4557);
and U6272 (N_6272,N_3269,N_4307);
nor U6273 (N_6273,N_2820,N_2952);
xor U6274 (N_6274,N_3528,N_4173);
nand U6275 (N_6275,N_4008,N_4747);
xor U6276 (N_6276,N_3267,N_4035);
or U6277 (N_6277,N_3592,N_4757);
nand U6278 (N_6278,N_3082,N_4280);
or U6279 (N_6279,N_2895,N_3957);
or U6280 (N_6280,N_3834,N_4309);
xnor U6281 (N_6281,N_4227,N_3151);
xor U6282 (N_6282,N_4910,N_3669);
xnor U6283 (N_6283,N_3511,N_4187);
xor U6284 (N_6284,N_4645,N_3376);
nand U6285 (N_6285,N_2736,N_2697);
xnor U6286 (N_6286,N_4304,N_3602);
or U6287 (N_6287,N_4379,N_3986);
nand U6288 (N_6288,N_3930,N_4086);
and U6289 (N_6289,N_3175,N_4707);
xnor U6290 (N_6290,N_2657,N_4935);
xor U6291 (N_6291,N_3322,N_4451);
or U6292 (N_6292,N_2620,N_4292);
and U6293 (N_6293,N_4543,N_3016);
nand U6294 (N_6294,N_4148,N_4604);
xnor U6295 (N_6295,N_4326,N_2684);
and U6296 (N_6296,N_3340,N_2781);
nor U6297 (N_6297,N_4415,N_2838);
nand U6298 (N_6298,N_3829,N_4478);
nand U6299 (N_6299,N_2577,N_4780);
nand U6300 (N_6300,N_3082,N_3486);
nor U6301 (N_6301,N_4684,N_2819);
nor U6302 (N_6302,N_3913,N_3441);
nand U6303 (N_6303,N_4996,N_3960);
xnor U6304 (N_6304,N_4542,N_4733);
nand U6305 (N_6305,N_4934,N_3251);
and U6306 (N_6306,N_3619,N_3889);
nand U6307 (N_6307,N_4149,N_3049);
nand U6308 (N_6308,N_2783,N_4120);
and U6309 (N_6309,N_3056,N_4820);
nand U6310 (N_6310,N_3668,N_4288);
xor U6311 (N_6311,N_4680,N_3818);
nand U6312 (N_6312,N_3864,N_3017);
nor U6313 (N_6313,N_3337,N_4797);
and U6314 (N_6314,N_4782,N_3622);
nor U6315 (N_6315,N_4820,N_3490);
nor U6316 (N_6316,N_2831,N_3629);
nand U6317 (N_6317,N_3389,N_3541);
or U6318 (N_6318,N_4236,N_3747);
nor U6319 (N_6319,N_3568,N_3627);
nor U6320 (N_6320,N_3411,N_4260);
xnor U6321 (N_6321,N_4535,N_4595);
nand U6322 (N_6322,N_4738,N_4169);
or U6323 (N_6323,N_4867,N_4753);
or U6324 (N_6324,N_2502,N_2833);
nand U6325 (N_6325,N_4755,N_3649);
xor U6326 (N_6326,N_4088,N_4807);
nor U6327 (N_6327,N_4183,N_3052);
xnor U6328 (N_6328,N_2593,N_4298);
nand U6329 (N_6329,N_3980,N_4622);
nand U6330 (N_6330,N_2689,N_3795);
xor U6331 (N_6331,N_4386,N_4702);
xnor U6332 (N_6332,N_4476,N_3364);
and U6333 (N_6333,N_4509,N_4878);
xnor U6334 (N_6334,N_3773,N_3920);
nor U6335 (N_6335,N_3942,N_4189);
nand U6336 (N_6336,N_3594,N_3344);
nor U6337 (N_6337,N_2670,N_4355);
nand U6338 (N_6338,N_4030,N_4816);
and U6339 (N_6339,N_3979,N_3069);
nor U6340 (N_6340,N_3101,N_4134);
or U6341 (N_6341,N_3334,N_3733);
and U6342 (N_6342,N_4479,N_3038);
nor U6343 (N_6343,N_2524,N_3330);
and U6344 (N_6344,N_3844,N_3234);
and U6345 (N_6345,N_4690,N_4441);
xor U6346 (N_6346,N_3644,N_3229);
or U6347 (N_6347,N_4615,N_3285);
nor U6348 (N_6348,N_4363,N_4162);
nor U6349 (N_6349,N_4914,N_2778);
xor U6350 (N_6350,N_3992,N_4418);
or U6351 (N_6351,N_4840,N_4658);
xnor U6352 (N_6352,N_4103,N_4474);
or U6353 (N_6353,N_4416,N_3548);
xnor U6354 (N_6354,N_4864,N_3492);
nand U6355 (N_6355,N_3383,N_4884);
nand U6356 (N_6356,N_3312,N_4925);
or U6357 (N_6357,N_3421,N_4744);
nand U6358 (N_6358,N_3997,N_4347);
and U6359 (N_6359,N_4002,N_4963);
nand U6360 (N_6360,N_4378,N_3286);
xnor U6361 (N_6361,N_3280,N_4056);
xnor U6362 (N_6362,N_3215,N_4497);
nor U6363 (N_6363,N_4894,N_3639);
and U6364 (N_6364,N_3699,N_2681);
and U6365 (N_6365,N_3494,N_3108);
nor U6366 (N_6366,N_3243,N_3572);
or U6367 (N_6367,N_3109,N_3599);
nand U6368 (N_6368,N_2983,N_2571);
nand U6369 (N_6369,N_2986,N_3624);
or U6370 (N_6370,N_3674,N_3033);
nor U6371 (N_6371,N_3556,N_4625);
nand U6372 (N_6372,N_4153,N_4925);
nand U6373 (N_6373,N_3438,N_4509);
xnor U6374 (N_6374,N_3360,N_3910);
xor U6375 (N_6375,N_4002,N_3974);
nand U6376 (N_6376,N_4831,N_3905);
or U6377 (N_6377,N_2912,N_4798);
nor U6378 (N_6378,N_3902,N_2875);
nor U6379 (N_6379,N_2960,N_2715);
or U6380 (N_6380,N_4099,N_2751);
and U6381 (N_6381,N_3889,N_4839);
nand U6382 (N_6382,N_4357,N_4581);
nand U6383 (N_6383,N_2520,N_4181);
and U6384 (N_6384,N_3792,N_3966);
or U6385 (N_6385,N_4027,N_2991);
or U6386 (N_6386,N_3372,N_2699);
xor U6387 (N_6387,N_2574,N_3260);
xnor U6388 (N_6388,N_4230,N_3331);
xnor U6389 (N_6389,N_4035,N_3703);
nor U6390 (N_6390,N_4805,N_4059);
nor U6391 (N_6391,N_2715,N_2639);
or U6392 (N_6392,N_3132,N_2727);
and U6393 (N_6393,N_3337,N_3184);
xnor U6394 (N_6394,N_2879,N_4552);
nand U6395 (N_6395,N_3939,N_2856);
xor U6396 (N_6396,N_4387,N_4218);
nor U6397 (N_6397,N_3625,N_2802);
and U6398 (N_6398,N_3469,N_3614);
or U6399 (N_6399,N_3730,N_4527);
nor U6400 (N_6400,N_4318,N_3322);
or U6401 (N_6401,N_4219,N_2699);
xnor U6402 (N_6402,N_3309,N_2997);
xnor U6403 (N_6403,N_4713,N_2689);
xor U6404 (N_6404,N_2710,N_4361);
and U6405 (N_6405,N_4036,N_4562);
and U6406 (N_6406,N_2553,N_2662);
and U6407 (N_6407,N_4006,N_4730);
xnor U6408 (N_6408,N_4241,N_2628);
nor U6409 (N_6409,N_4376,N_2565);
nor U6410 (N_6410,N_3512,N_3543);
nand U6411 (N_6411,N_3045,N_2890);
xnor U6412 (N_6412,N_4700,N_2955);
and U6413 (N_6413,N_2877,N_2669);
nor U6414 (N_6414,N_4239,N_4073);
nand U6415 (N_6415,N_4769,N_4272);
and U6416 (N_6416,N_2882,N_3698);
nand U6417 (N_6417,N_3866,N_4368);
nand U6418 (N_6418,N_3458,N_2839);
nand U6419 (N_6419,N_4295,N_2756);
xnor U6420 (N_6420,N_4425,N_3652);
and U6421 (N_6421,N_2538,N_2622);
nor U6422 (N_6422,N_3806,N_4247);
xor U6423 (N_6423,N_2787,N_3528);
nor U6424 (N_6424,N_2975,N_4317);
nor U6425 (N_6425,N_3965,N_4046);
nor U6426 (N_6426,N_3754,N_4926);
and U6427 (N_6427,N_3570,N_3414);
nand U6428 (N_6428,N_3339,N_3919);
xor U6429 (N_6429,N_3973,N_4025);
xor U6430 (N_6430,N_2639,N_3488);
or U6431 (N_6431,N_2923,N_3401);
xor U6432 (N_6432,N_4581,N_3130);
nor U6433 (N_6433,N_4764,N_4852);
and U6434 (N_6434,N_3615,N_3416);
nand U6435 (N_6435,N_3760,N_3904);
or U6436 (N_6436,N_3387,N_2509);
or U6437 (N_6437,N_4968,N_3568);
nor U6438 (N_6438,N_3285,N_2908);
nor U6439 (N_6439,N_4432,N_4051);
or U6440 (N_6440,N_3818,N_4156);
or U6441 (N_6441,N_3580,N_4598);
and U6442 (N_6442,N_4308,N_3357);
and U6443 (N_6443,N_3135,N_4052);
and U6444 (N_6444,N_4398,N_2829);
nand U6445 (N_6445,N_3200,N_2822);
nor U6446 (N_6446,N_4379,N_4415);
or U6447 (N_6447,N_3690,N_3142);
and U6448 (N_6448,N_3268,N_3371);
nor U6449 (N_6449,N_3326,N_4468);
or U6450 (N_6450,N_2693,N_4485);
or U6451 (N_6451,N_4851,N_3488);
xor U6452 (N_6452,N_3272,N_2621);
xor U6453 (N_6453,N_2612,N_2639);
nor U6454 (N_6454,N_3309,N_3064);
xor U6455 (N_6455,N_3371,N_4296);
xor U6456 (N_6456,N_3983,N_4840);
xor U6457 (N_6457,N_4069,N_2682);
or U6458 (N_6458,N_2919,N_4499);
and U6459 (N_6459,N_4368,N_2507);
nand U6460 (N_6460,N_3456,N_4218);
nand U6461 (N_6461,N_3483,N_4267);
nor U6462 (N_6462,N_2910,N_4314);
nand U6463 (N_6463,N_4324,N_4561);
xnor U6464 (N_6464,N_2688,N_2844);
xnor U6465 (N_6465,N_3799,N_2751);
xor U6466 (N_6466,N_4890,N_3362);
or U6467 (N_6467,N_4832,N_2604);
nor U6468 (N_6468,N_3510,N_4526);
and U6469 (N_6469,N_3732,N_4463);
and U6470 (N_6470,N_3959,N_3174);
nand U6471 (N_6471,N_3054,N_3154);
and U6472 (N_6472,N_2674,N_4263);
or U6473 (N_6473,N_3205,N_2743);
nand U6474 (N_6474,N_3761,N_3313);
nor U6475 (N_6475,N_4112,N_4350);
or U6476 (N_6476,N_4291,N_4435);
xnor U6477 (N_6477,N_3881,N_2529);
nor U6478 (N_6478,N_4716,N_4782);
xnor U6479 (N_6479,N_2507,N_3632);
nor U6480 (N_6480,N_2596,N_3753);
nand U6481 (N_6481,N_4343,N_4898);
nor U6482 (N_6482,N_3725,N_3917);
xnor U6483 (N_6483,N_3993,N_2777);
nand U6484 (N_6484,N_3979,N_4639);
and U6485 (N_6485,N_4028,N_3664);
and U6486 (N_6486,N_3172,N_3799);
xnor U6487 (N_6487,N_4944,N_4695);
or U6488 (N_6488,N_3217,N_4288);
nand U6489 (N_6489,N_3374,N_4318);
and U6490 (N_6490,N_3943,N_4392);
nor U6491 (N_6491,N_4624,N_3985);
and U6492 (N_6492,N_4802,N_2525);
and U6493 (N_6493,N_2903,N_3139);
nor U6494 (N_6494,N_3087,N_2988);
and U6495 (N_6495,N_2728,N_2791);
nor U6496 (N_6496,N_4950,N_3761);
or U6497 (N_6497,N_3593,N_4473);
or U6498 (N_6498,N_4466,N_2619);
or U6499 (N_6499,N_4037,N_3022);
or U6500 (N_6500,N_4975,N_3251);
xnor U6501 (N_6501,N_3121,N_3494);
xnor U6502 (N_6502,N_3890,N_3551);
or U6503 (N_6503,N_4641,N_2537);
nand U6504 (N_6504,N_4156,N_4894);
and U6505 (N_6505,N_4637,N_3664);
nand U6506 (N_6506,N_2592,N_3052);
or U6507 (N_6507,N_2962,N_4736);
xor U6508 (N_6508,N_3176,N_3116);
and U6509 (N_6509,N_2689,N_4478);
and U6510 (N_6510,N_4853,N_3527);
nor U6511 (N_6511,N_4539,N_4208);
and U6512 (N_6512,N_4745,N_2831);
nor U6513 (N_6513,N_3677,N_2969);
nand U6514 (N_6514,N_3621,N_4833);
xor U6515 (N_6515,N_2830,N_3104);
nor U6516 (N_6516,N_3509,N_3359);
and U6517 (N_6517,N_4909,N_2596);
xor U6518 (N_6518,N_2777,N_3480);
and U6519 (N_6519,N_4214,N_4970);
xor U6520 (N_6520,N_3726,N_4027);
nor U6521 (N_6521,N_3034,N_3463);
nor U6522 (N_6522,N_3289,N_3662);
nor U6523 (N_6523,N_2893,N_2890);
xor U6524 (N_6524,N_4584,N_4893);
nor U6525 (N_6525,N_3282,N_2501);
nand U6526 (N_6526,N_4389,N_2916);
nand U6527 (N_6527,N_3453,N_3858);
nor U6528 (N_6528,N_4961,N_3224);
nor U6529 (N_6529,N_4998,N_4344);
or U6530 (N_6530,N_4783,N_3689);
and U6531 (N_6531,N_2523,N_4229);
or U6532 (N_6532,N_4305,N_2811);
and U6533 (N_6533,N_4357,N_3149);
or U6534 (N_6534,N_4421,N_2762);
xnor U6535 (N_6535,N_2939,N_3898);
or U6536 (N_6536,N_4370,N_4301);
nor U6537 (N_6537,N_3271,N_2627);
nand U6538 (N_6538,N_4117,N_4681);
xor U6539 (N_6539,N_3573,N_3171);
and U6540 (N_6540,N_2589,N_3525);
nor U6541 (N_6541,N_3318,N_4994);
xor U6542 (N_6542,N_2715,N_4878);
nor U6543 (N_6543,N_4832,N_3046);
or U6544 (N_6544,N_2588,N_3464);
nor U6545 (N_6545,N_3770,N_3228);
and U6546 (N_6546,N_4295,N_3501);
nand U6547 (N_6547,N_2820,N_3724);
and U6548 (N_6548,N_3790,N_3972);
nand U6549 (N_6549,N_4192,N_3240);
or U6550 (N_6550,N_3410,N_4839);
and U6551 (N_6551,N_2819,N_4318);
nand U6552 (N_6552,N_3554,N_2798);
and U6553 (N_6553,N_4882,N_4042);
or U6554 (N_6554,N_4621,N_3131);
xnor U6555 (N_6555,N_3732,N_3344);
or U6556 (N_6556,N_4618,N_2763);
nor U6557 (N_6557,N_4272,N_4444);
and U6558 (N_6558,N_4951,N_3101);
or U6559 (N_6559,N_3631,N_4900);
or U6560 (N_6560,N_3032,N_2665);
nor U6561 (N_6561,N_3118,N_2712);
nand U6562 (N_6562,N_2777,N_2662);
nand U6563 (N_6563,N_3490,N_3449);
nor U6564 (N_6564,N_4796,N_4062);
and U6565 (N_6565,N_3699,N_4166);
nor U6566 (N_6566,N_4113,N_4674);
nand U6567 (N_6567,N_2710,N_3082);
nand U6568 (N_6568,N_3309,N_4618);
xnor U6569 (N_6569,N_3624,N_3778);
and U6570 (N_6570,N_4096,N_3565);
nand U6571 (N_6571,N_3499,N_4563);
nand U6572 (N_6572,N_3985,N_3685);
or U6573 (N_6573,N_3085,N_4434);
nand U6574 (N_6574,N_3424,N_3408);
xnor U6575 (N_6575,N_3546,N_3615);
and U6576 (N_6576,N_3917,N_4255);
nand U6577 (N_6577,N_2519,N_3788);
nor U6578 (N_6578,N_3173,N_2901);
or U6579 (N_6579,N_4665,N_4398);
and U6580 (N_6580,N_3887,N_3601);
and U6581 (N_6581,N_4017,N_3609);
and U6582 (N_6582,N_3023,N_4396);
and U6583 (N_6583,N_4111,N_3859);
and U6584 (N_6584,N_3035,N_3422);
or U6585 (N_6585,N_3253,N_2544);
xor U6586 (N_6586,N_2579,N_3424);
nand U6587 (N_6587,N_4193,N_3742);
and U6588 (N_6588,N_4599,N_2718);
nor U6589 (N_6589,N_3039,N_4076);
or U6590 (N_6590,N_3154,N_3830);
or U6591 (N_6591,N_4533,N_4620);
nor U6592 (N_6592,N_3222,N_4914);
or U6593 (N_6593,N_3573,N_4252);
and U6594 (N_6594,N_4175,N_3064);
xor U6595 (N_6595,N_4299,N_4991);
nand U6596 (N_6596,N_4384,N_3233);
and U6597 (N_6597,N_3072,N_3138);
xor U6598 (N_6598,N_3006,N_2981);
xnor U6599 (N_6599,N_4884,N_4845);
and U6600 (N_6600,N_4304,N_4846);
or U6601 (N_6601,N_4803,N_3433);
or U6602 (N_6602,N_3853,N_3174);
and U6603 (N_6603,N_3679,N_4842);
and U6604 (N_6604,N_2697,N_4201);
or U6605 (N_6605,N_2783,N_3950);
nor U6606 (N_6606,N_2591,N_3460);
or U6607 (N_6607,N_3501,N_4677);
or U6608 (N_6608,N_4872,N_4828);
nor U6609 (N_6609,N_3828,N_3050);
and U6610 (N_6610,N_3596,N_4509);
nor U6611 (N_6611,N_3801,N_4535);
nand U6612 (N_6612,N_4844,N_4238);
nor U6613 (N_6613,N_4246,N_3576);
and U6614 (N_6614,N_4043,N_3637);
xor U6615 (N_6615,N_4587,N_3493);
nand U6616 (N_6616,N_4189,N_4646);
nor U6617 (N_6617,N_3577,N_3822);
and U6618 (N_6618,N_2562,N_3496);
and U6619 (N_6619,N_4780,N_4972);
nor U6620 (N_6620,N_3241,N_3228);
xnor U6621 (N_6621,N_3058,N_4567);
and U6622 (N_6622,N_3013,N_2906);
and U6623 (N_6623,N_3060,N_4667);
nor U6624 (N_6624,N_3950,N_3425);
nor U6625 (N_6625,N_4662,N_4164);
and U6626 (N_6626,N_3755,N_4670);
nand U6627 (N_6627,N_4374,N_4290);
or U6628 (N_6628,N_3696,N_4474);
nor U6629 (N_6629,N_2849,N_4812);
nand U6630 (N_6630,N_2536,N_2585);
nand U6631 (N_6631,N_3525,N_2532);
and U6632 (N_6632,N_3874,N_4929);
nor U6633 (N_6633,N_2913,N_2690);
nor U6634 (N_6634,N_4937,N_2738);
nand U6635 (N_6635,N_3937,N_2628);
nor U6636 (N_6636,N_3680,N_2986);
nor U6637 (N_6637,N_3929,N_4597);
nand U6638 (N_6638,N_4064,N_2848);
xor U6639 (N_6639,N_4334,N_4522);
nor U6640 (N_6640,N_4953,N_4856);
and U6641 (N_6641,N_4698,N_3040);
or U6642 (N_6642,N_2536,N_4646);
or U6643 (N_6643,N_3363,N_4655);
nor U6644 (N_6644,N_3117,N_4044);
or U6645 (N_6645,N_3437,N_3465);
nor U6646 (N_6646,N_4462,N_3639);
and U6647 (N_6647,N_2926,N_2980);
nand U6648 (N_6648,N_3590,N_3597);
nor U6649 (N_6649,N_4231,N_4886);
nor U6650 (N_6650,N_4291,N_4811);
and U6651 (N_6651,N_4561,N_4158);
xnor U6652 (N_6652,N_4849,N_4898);
or U6653 (N_6653,N_4906,N_3172);
nor U6654 (N_6654,N_2546,N_4212);
and U6655 (N_6655,N_3845,N_4296);
nand U6656 (N_6656,N_4963,N_3865);
and U6657 (N_6657,N_2907,N_2617);
or U6658 (N_6658,N_4307,N_3987);
and U6659 (N_6659,N_4139,N_2805);
or U6660 (N_6660,N_3674,N_2692);
and U6661 (N_6661,N_4751,N_3461);
xnor U6662 (N_6662,N_2676,N_2945);
nand U6663 (N_6663,N_3813,N_4728);
nand U6664 (N_6664,N_2734,N_4295);
xnor U6665 (N_6665,N_3949,N_3121);
nand U6666 (N_6666,N_2936,N_4024);
and U6667 (N_6667,N_2984,N_4845);
nand U6668 (N_6668,N_3901,N_4452);
or U6669 (N_6669,N_3009,N_4673);
and U6670 (N_6670,N_2541,N_4797);
nor U6671 (N_6671,N_4094,N_4365);
xnor U6672 (N_6672,N_4794,N_4435);
nor U6673 (N_6673,N_4246,N_2938);
nor U6674 (N_6674,N_3295,N_4475);
or U6675 (N_6675,N_2834,N_3922);
nand U6676 (N_6676,N_4739,N_3648);
or U6677 (N_6677,N_2581,N_3255);
nand U6678 (N_6678,N_3563,N_4915);
nor U6679 (N_6679,N_3621,N_2835);
xor U6680 (N_6680,N_4863,N_4980);
xor U6681 (N_6681,N_3689,N_3160);
nor U6682 (N_6682,N_2813,N_2739);
and U6683 (N_6683,N_3106,N_4554);
nor U6684 (N_6684,N_3089,N_3918);
nor U6685 (N_6685,N_4164,N_3724);
and U6686 (N_6686,N_4992,N_3183);
xnor U6687 (N_6687,N_2702,N_4359);
and U6688 (N_6688,N_3081,N_2527);
and U6689 (N_6689,N_4270,N_2682);
and U6690 (N_6690,N_3251,N_4992);
nand U6691 (N_6691,N_2721,N_2799);
or U6692 (N_6692,N_2922,N_4708);
nand U6693 (N_6693,N_3327,N_2546);
and U6694 (N_6694,N_2691,N_4545);
and U6695 (N_6695,N_4278,N_2813);
xor U6696 (N_6696,N_3736,N_3793);
or U6697 (N_6697,N_4939,N_3620);
or U6698 (N_6698,N_3359,N_3111);
and U6699 (N_6699,N_2878,N_4107);
or U6700 (N_6700,N_4632,N_3846);
nor U6701 (N_6701,N_4635,N_3019);
xor U6702 (N_6702,N_2830,N_3388);
or U6703 (N_6703,N_3556,N_4782);
xor U6704 (N_6704,N_4538,N_4015);
or U6705 (N_6705,N_3867,N_4704);
and U6706 (N_6706,N_3977,N_3263);
xor U6707 (N_6707,N_2652,N_4991);
and U6708 (N_6708,N_3983,N_4018);
and U6709 (N_6709,N_4459,N_4959);
xor U6710 (N_6710,N_2991,N_4248);
or U6711 (N_6711,N_4732,N_3792);
and U6712 (N_6712,N_4785,N_4169);
and U6713 (N_6713,N_4265,N_3469);
and U6714 (N_6714,N_3842,N_4658);
nor U6715 (N_6715,N_4854,N_4660);
nor U6716 (N_6716,N_3834,N_4051);
xor U6717 (N_6717,N_4236,N_2929);
nor U6718 (N_6718,N_4380,N_3158);
nor U6719 (N_6719,N_4664,N_3868);
xnor U6720 (N_6720,N_2564,N_3026);
and U6721 (N_6721,N_2566,N_4735);
nor U6722 (N_6722,N_3201,N_4777);
and U6723 (N_6723,N_3820,N_3827);
and U6724 (N_6724,N_3161,N_3281);
xor U6725 (N_6725,N_3035,N_2874);
or U6726 (N_6726,N_3534,N_3719);
or U6727 (N_6727,N_4459,N_4641);
nand U6728 (N_6728,N_4622,N_4664);
or U6729 (N_6729,N_2525,N_4882);
or U6730 (N_6730,N_3358,N_4303);
xor U6731 (N_6731,N_4807,N_2806);
or U6732 (N_6732,N_2787,N_4083);
nand U6733 (N_6733,N_4529,N_3942);
and U6734 (N_6734,N_2853,N_2743);
xor U6735 (N_6735,N_3442,N_4346);
and U6736 (N_6736,N_4823,N_3247);
or U6737 (N_6737,N_3138,N_4523);
xnor U6738 (N_6738,N_3035,N_4433);
xnor U6739 (N_6739,N_3937,N_3843);
or U6740 (N_6740,N_3836,N_2579);
or U6741 (N_6741,N_3078,N_3721);
nand U6742 (N_6742,N_3665,N_3970);
nand U6743 (N_6743,N_3832,N_3393);
or U6744 (N_6744,N_3887,N_4395);
nor U6745 (N_6745,N_3265,N_2663);
xnor U6746 (N_6746,N_2578,N_4146);
xnor U6747 (N_6747,N_4362,N_3207);
nor U6748 (N_6748,N_4631,N_3121);
xor U6749 (N_6749,N_3599,N_4528);
nand U6750 (N_6750,N_3680,N_2922);
or U6751 (N_6751,N_2731,N_2799);
and U6752 (N_6752,N_4367,N_4359);
nor U6753 (N_6753,N_4436,N_3743);
nor U6754 (N_6754,N_3114,N_4701);
nor U6755 (N_6755,N_3114,N_4285);
or U6756 (N_6756,N_3404,N_4782);
and U6757 (N_6757,N_3702,N_4762);
and U6758 (N_6758,N_4239,N_2553);
or U6759 (N_6759,N_2691,N_3868);
xnor U6760 (N_6760,N_2777,N_4324);
or U6761 (N_6761,N_4872,N_2831);
nand U6762 (N_6762,N_3612,N_3651);
xnor U6763 (N_6763,N_4321,N_4614);
nor U6764 (N_6764,N_4154,N_3257);
nor U6765 (N_6765,N_4262,N_3336);
nand U6766 (N_6766,N_3571,N_2588);
and U6767 (N_6767,N_3439,N_3150);
xnor U6768 (N_6768,N_2519,N_4083);
and U6769 (N_6769,N_2624,N_3856);
nor U6770 (N_6770,N_2575,N_4104);
or U6771 (N_6771,N_3330,N_3911);
and U6772 (N_6772,N_2857,N_4876);
and U6773 (N_6773,N_4449,N_2611);
and U6774 (N_6774,N_3125,N_3906);
and U6775 (N_6775,N_3166,N_3818);
nand U6776 (N_6776,N_4731,N_3065);
or U6777 (N_6777,N_2900,N_4120);
nand U6778 (N_6778,N_3739,N_3368);
or U6779 (N_6779,N_4340,N_4031);
or U6780 (N_6780,N_4148,N_4167);
or U6781 (N_6781,N_2685,N_3815);
nor U6782 (N_6782,N_2847,N_4422);
nand U6783 (N_6783,N_2863,N_4240);
or U6784 (N_6784,N_4835,N_2517);
or U6785 (N_6785,N_4762,N_3009);
nor U6786 (N_6786,N_3385,N_4996);
or U6787 (N_6787,N_2521,N_2675);
nor U6788 (N_6788,N_3298,N_4134);
or U6789 (N_6789,N_3298,N_4745);
and U6790 (N_6790,N_4411,N_2587);
nor U6791 (N_6791,N_3484,N_4846);
and U6792 (N_6792,N_4418,N_3060);
xor U6793 (N_6793,N_3308,N_3002);
and U6794 (N_6794,N_2531,N_4308);
nand U6795 (N_6795,N_2951,N_4401);
nor U6796 (N_6796,N_2861,N_4295);
and U6797 (N_6797,N_4785,N_3329);
or U6798 (N_6798,N_3693,N_4431);
xnor U6799 (N_6799,N_4409,N_2843);
nor U6800 (N_6800,N_3259,N_4877);
nand U6801 (N_6801,N_2926,N_4269);
nand U6802 (N_6802,N_3637,N_2823);
or U6803 (N_6803,N_2712,N_3578);
and U6804 (N_6804,N_4897,N_4267);
and U6805 (N_6805,N_4416,N_3713);
xor U6806 (N_6806,N_3880,N_4056);
nor U6807 (N_6807,N_3172,N_4178);
or U6808 (N_6808,N_4551,N_4863);
and U6809 (N_6809,N_4597,N_2794);
or U6810 (N_6810,N_2729,N_3471);
and U6811 (N_6811,N_4148,N_3053);
nor U6812 (N_6812,N_4587,N_2776);
nand U6813 (N_6813,N_4069,N_2581);
xnor U6814 (N_6814,N_3537,N_4359);
and U6815 (N_6815,N_4760,N_3525);
xor U6816 (N_6816,N_3795,N_3752);
nor U6817 (N_6817,N_4182,N_4217);
or U6818 (N_6818,N_2697,N_4680);
xor U6819 (N_6819,N_2647,N_4220);
xnor U6820 (N_6820,N_4844,N_3085);
and U6821 (N_6821,N_3938,N_3561);
nor U6822 (N_6822,N_2535,N_2595);
nand U6823 (N_6823,N_4646,N_4196);
or U6824 (N_6824,N_3504,N_3337);
or U6825 (N_6825,N_4792,N_3119);
nor U6826 (N_6826,N_3722,N_4251);
xor U6827 (N_6827,N_3179,N_3074);
nand U6828 (N_6828,N_4903,N_3574);
or U6829 (N_6829,N_4420,N_4547);
xor U6830 (N_6830,N_3896,N_4951);
xor U6831 (N_6831,N_2803,N_3448);
or U6832 (N_6832,N_3803,N_4103);
nor U6833 (N_6833,N_2624,N_3263);
nand U6834 (N_6834,N_4192,N_2794);
or U6835 (N_6835,N_3021,N_3610);
or U6836 (N_6836,N_3399,N_3807);
xor U6837 (N_6837,N_4198,N_3098);
xnor U6838 (N_6838,N_2847,N_4247);
nor U6839 (N_6839,N_3734,N_3649);
and U6840 (N_6840,N_3689,N_4341);
or U6841 (N_6841,N_4868,N_2885);
nand U6842 (N_6842,N_3638,N_4731);
nor U6843 (N_6843,N_4083,N_3593);
nand U6844 (N_6844,N_3659,N_3343);
and U6845 (N_6845,N_3021,N_4398);
nand U6846 (N_6846,N_4163,N_3200);
and U6847 (N_6847,N_3010,N_3969);
nor U6848 (N_6848,N_3580,N_3961);
nand U6849 (N_6849,N_2583,N_3176);
and U6850 (N_6850,N_3504,N_3880);
nand U6851 (N_6851,N_4410,N_4127);
or U6852 (N_6852,N_4041,N_3935);
or U6853 (N_6853,N_3229,N_3033);
or U6854 (N_6854,N_4384,N_2588);
nand U6855 (N_6855,N_3276,N_4372);
and U6856 (N_6856,N_3702,N_4949);
nor U6857 (N_6857,N_3688,N_3893);
xor U6858 (N_6858,N_3800,N_4498);
nor U6859 (N_6859,N_4362,N_3673);
or U6860 (N_6860,N_2518,N_3520);
nand U6861 (N_6861,N_3882,N_2510);
nand U6862 (N_6862,N_3819,N_4126);
nand U6863 (N_6863,N_3840,N_4693);
and U6864 (N_6864,N_2523,N_3681);
and U6865 (N_6865,N_4130,N_3083);
nand U6866 (N_6866,N_4202,N_4151);
nor U6867 (N_6867,N_4640,N_3565);
nand U6868 (N_6868,N_3710,N_4578);
and U6869 (N_6869,N_3081,N_2936);
nor U6870 (N_6870,N_3515,N_4073);
nand U6871 (N_6871,N_4500,N_3254);
nor U6872 (N_6872,N_2912,N_4405);
nand U6873 (N_6873,N_3776,N_4277);
or U6874 (N_6874,N_2589,N_4734);
xnor U6875 (N_6875,N_4645,N_4895);
and U6876 (N_6876,N_3799,N_2787);
and U6877 (N_6877,N_2722,N_4930);
or U6878 (N_6878,N_4535,N_2538);
xnor U6879 (N_6879,N_4779,N_3610);
nand U6880 (N_6880,N_4349,N_4789);
xor U6881 (N_6881,N_2862,N_2743);
nand U6882 (N_6882,N_4890,N_4348);
xnor U6883 (N_6883,N_2579,N_3008);
nor U6884 (N_6884,N_3894,N_3451);
and U6885 (N_6885,N_4553,N_4368);
nand U6886 (N_6886,N_2618,N_2606);
or U6887 (N_6887,N_3028,N_3927);
nand U6888 (N_6888,N_4799,N_4446);
xnor U6889 (N_6889,N_3180,N_3673);
nand U6890 (N_6890,N_4376,N_4395);
xnor U6891 (N_6891,N_4481,N_3089);
or U6892 (N_6892,N_4120,N_4962);
nor U6893 (N_6893,N_3736,N_2562);
nor U6894 (N_6894,N_4193,N_2899);
nand U6895 (N_6895,N_4550,N_3099);
or U6896 (N_6896,N_4443,N_2703);
xnor U6897 (N_6897,N_2594,N_3936);
nand U6898 (N_6898,N_3711,N_4698);
or U6899 (N_6899,N_2819,N_2534);
and U6900 (N_6900,N_4843,N_4215);
and U6901 (N_6901,N_2534,N_4611);
nand U6902 (N_6902,N_2634,N_4231);
nor U6903 (N_6903,N_3251,N_4712);
and U6904 (N_6904,N_4127,N_3828);
nand U6905 (N_6905,N_3927,N_4641);
nand U6906 (N_6906,N_3152,N_2941);
and U6907 (N_6907,N_3265,N_3775);
and U6908 (N_6908,N_2738,N_4198);
xor U6909 (N_6909,N_3123,N_3760);
xnor U6910 (N_6910,N_2663,N_3425);
or U6911 (N_6911,N_4696,N_3378);
nor U6912 (N_6912,N_3178,N_2750);
and U6913 (N_6913,N_3865,N_4196);
xnor U6914 (N_6914,N_4012,N_4791);
and U6915 (N_6915,N_3743,N_2513);
or U6916 (N_6916,N_4534,N_4846);
and U6917 (N_6917,N_3827,N_3491);
and U6918 (N_6918,N_3656,N_4493);
or U6919 (N_6919,N_2939,N_4339);
or U6920 (N_6920,N_4773,N_4408);
xor U6921 (N_6921,N_4928,N_4030);
and U6922 (N_6922,N_4229,N_2969);
nand U6923 (N_6923,N_3451,N_4579);
or U6924 (N_6924,N_4300,N_3698);
nor U6925 (N_6925,N_3268,N_3732);
and U6926 (N_6926,N_3705,N_2968);
nand U6927 (N_6927,N_2507,N_3366);
and U6928 (N_6928,N_2837,N_4841);
or U6929 (N_6929,N_3786,N_3002);
xnor U6930 (N_6930,N_2650,N_2581);
nand U6931 (N_6931,N_3967,N_3757);
and U6932 (N_6932,N_3116,N_3237);
or U6933 (N_6933,N_4864,N_2617);
xor U6934 (N_6934,N_3849,N_4763);
nor U6935 (N_6935,N_4303,N_3437);
nor U6936 (N_6936,N_4200,N_3504);
or U6937 (N_6937,N_4127,N_4609);
xor U6938 (N_6938,N_3133,N_4927);
xor U6939 (N_6939,N_4096,N_4345);
nor U6940 (N_6940,N_3938,N_4250);
or U6941 (N_6941,N_4573,N_3124);
nor U6942 (N_6942,N_4848,N_4652);
xnor U6943 (N_6943,N_2845,N_2570);
xor U6944 (N_6944,N_2871,N_3319);
and U6945 (N_6945,N_2532,N_2982);
xor U6946 (N_6946,N_4004,N_3886);
and U6947 (N_6947,N_4381,N_4349);
xor U6948 (N_6948,N_3968,N_2969);
nand U6949 (N_6949,N_2921,N_4281);
xor U6950 (N_6950,N_2908,N_4492);
xor U6951 (N_6951,N_3611,N_4250);
nand U6952 (N_6952,N_3800,N_4563);
and U6953 (N_6953,N_3154,N_3363);
nand U6954 (N_6954,N_3980,N_4708);
and U6955 (N_6955,N_3329,N_4942);
nand U6956 (N_6956,N_3074,N_4643);
nand U6957 (N_6957,N_4363,N_3478);
and U6958 (N_6958,N_4055,N_4588);
xnor U6959 (N_6959,N_3217,N_3604);
nor U6960 (N_6960,N_3770,N_4877);
xnor U6961 (N_6961,N_2880,N_2802);
nor U6962 (N_6962,N_2840,N_4049);
and U6963 (N_6963,N_3122,N_4077);
xor U6964 (N_6964,N_4465,N_3510);
xnor U6965 (N_6965,N_2644,N_3482);
nand U6966 (N_6966,N_3283,N_3502);
xor U6967 (N_6967,N_3523,N_4379);
xnor U6968 (N_6968,N_2668,N_2657);
xnor U6969 (N_6969,N_3806,N_3978);
nor U6970 (N_6970,N_4027,N_3886);
xnor U6971 (N_6971,N_3134,N_4202);
nor U6972 (N_6972,N_4544,N_4592);
nor U6973 (N_6973,N_4830,N_3676);
nor U6974 (N_6974,N_2782,N_4185);
or U6975 (N_6975,N_3024,N_2939);
nor U6976 (N_6976,N_4803,N_4698);
or U6977 (N_6977,N_4933,N_3795);
or U6978 (N_6978,N_3738,N_3113);
xnor U6979 (N_6979,N_2673,N_4805);
xnor U6980 (N_6980,N_4490,N_2601);
nand U6981 (N_6981,N_2658,N_4409);
nand U6982 (N_6982,N_4555,N_2921);
and U6983 (N_6983,N_4866,N_2595);
nand U6984 (N_6984,N_4281,N_2961);
nand U6985 (N_6985,N_2616,N_2951);
nor U6986 (N_6986,N_4454,N_4594);
xor U6987 (N_6987,N_4518,N_2790);
xnor U6988 (N_6988,N_4179,N_3665);
or U6989 (N_6989,N_3079,N_3619);
or U6990 (N_6990,N_4497,N_2816);
nor U6991 (N_6991,N_3473,N_2602);
and U6992 (N_6992,N_4760,N_3727);
nand U6993 (N_6993,N_3717,N_3291);
xor U6994 (N_6994,N_3891,N_4800);
nor U6995 (N_6995,N_3815,N_2737);
nand U6996 (N_6996,N_2606,N_2782);
or U6997 (N_6997,N_4817,N_4176);
and U6998 (N_6998,N_2888,N_4047);
nand U6999 (N_6999,N_4493,N_4453);
and U7000 (N_7000,N_4044,N_3351);
xor U7001 (N_7001,N_4589,N_4981);
nand U7002 (N_7002,N_3355,N_3273);
and U7003 (N_7003,N_2870,N_3122);
or U7004 (N_7004,N_4233,N_4294);
or U7005 (N_7005,N_4162,N_3886);
or U7006 (N_7006,N_4560,N_2680);
xnor U7007 (N_7007,N_3619,N_3890);
nor U7008 (N_7008,N_4171,N_4512);
or U7009 (N_7009,N_3593,N_3027);
and U7010 (N_7010,N_2917,N_4179);
or U7011 (N_7011,N_3739,N_3809);
nor U7012 (N_7012,N_4021,N_4943);
or U7013 (N_7013,N_3085,N_3224);
and U7014 (N_7014,N_2944,N_4941);
and U7015 (N_7015,N_4828,N_3213);
nor U7016 (N_7016,N_4972,N_4700);
nor U7017 (N_7017,N_3567,N_4229);
or U7018 (N_7018,N_2607,N_3280);
nand U7019 (N_7019,N_4720,N_3889);
xor U7020 (N_7020,N_4676,N_3803);
nand U7021 (N_7021,N_3738,N_2905);
xor U7022 (N_7022,N_3948,N_4520);
nor U7023 (N_7023,N_2901,N_4136);
xnor U7024 (N_7024,N_3296,N_4629);
or U7025 (N_7025,N_4247,N_3332);
nor U7026 (N_7026,N_2764,N_3807);
xnor U7027 (N_7027,N_4952,N_3108);
nand U7028 (N_7028,N_4010,N_2850);
nand U7029 (N_7029,N_3284,N_2800);
and U7030 (N_7030,N_3266,N_2820);
and U7031 (N_7031,N_3680,N_4502);
or U7032 (N_7032,N_2742,N_4125);
nand U7033 (N_7033,N_3913,N_3643);
and U7034 (N_7034,N_3081,N_2614);
or U7035 (N_7035,N_4975,N_2998);
nand U7036 (N_7036,N_4154,N_3926);
and U7037 (N_7037,N_4781,N_2642);
or U7038 (N_7038,N_3671,N_4699);
and U7039 (N_7039,N_2968,N_3824);
and U7040 (N_7040,N_3569,N_2755);
and U7041 (N_7041,N_4948,N_4472);
and U7042 (N_7042,N_4162,N_4424);
and U7043 (N_7043,N_3607,N_4905);
or U7044 (N_7044,N_4978,N_3502);
nand U7045 (N_7045,N_3462,N_4729);
nor U7046 (N_7046,N_4702,N_4030);
and U7047 (N_7047,N_2826,N_3624);
nor U7048 (N_7048,N_4164,N_3246);
and U7049 (N_7049,N_3306,N_2831);
nor U7050 (N_7050,N_3333,N_2798);
or U7051 (N_7051,N_4973,N_3478);
nand U7052 (N_7052,N_4755,N_2679);
or U7053 (N_7053,N_4357,N_4617);
and U7054 (N_7054,N_4801,N_3234);
xor U7055 (N_7055,N_3630,N_4397);
nand U7056 (N_7056,N_4367,N_2664);
xnor U7057 (N_7057,N_2961,N_4866);
or U7058 (N_7058,N_3309,N_3550);
or U7059 (N_7059,N_4057,N_2759);
nand U7060 (N_7060,N_2632,N_2854);
and U7061 (N_7061,N_4718,N_4542);
or U7062 (N_7062,N_3378,N_3401);
nor U7063 (N_7063,N_4768,N_4614);
xor U7064 (N_7064,N_3306,N_2714);
nor U7065 (N_7065,N_4771,N_4654);
xnor U7066 (N_7066,N_2938,N_3384);
xnor U7067 (N_7067,N_4761,N_2521);
or U7068 (N_7068,N_3738,N_4170);
nor U7069 (N_7069,N_2577,N_2826);
or U7070 (N_7070,N_4926,N_3902);
nor U7071 (N_7071,N_3440,N_4133);
nor U7072 (N_7072,N_3616,N_3040);
or U7073 (N_7073,N_2646,N_3107);
nand U7074 (N_7074,N_4515,N_2887);
and U7075 (N_7075,N_4118,N_4163);
xor U7076 (N_7076,N_3795,N_3823);
and U7077 (N_7077,N_2510,N_3437);
nand U7078 (N_7078,N_3789,N_4466);
and U7079 (N_7079,N_4708,N_3839);
and U7080 (N_7080,N_3277,N_3058);
xnor U7081 (N_7081,N_4022,N_4412);
and U7082 (N_7082,N_4926,N_3568);
nand U7083 (N_7083,N_4707,N_4172);
nor U7084 (N_7084,N_3157,N_4779);
nor U7085 (N_7085,N_4476,N_3271);
nand U7086 (N_7086,N_4901,N_4469);
or U7087 (N_7087,N_3281,N_4099);
nand U7088 (N_7088,N_2824,N_4510);
or U7089 (N_7089,N_4534,N_3289);
xor U7090 (N_7090,N_3984,N_4548);
xor U7091 (N_7091,N_4986,N_4543);
nor U7092 (N_7092,N_4451,N_3717);
xnor U7093 (N_7093,N_4689,N_4942);
and U7094 (N_7094,N_3646,N_3990);
or U7095 (N_7095,N_4813,N_4435);
xor U7096 (N_7096,N_3095,N_4393);
nand U7097 (N_7097,N_3274,N_2698);
nor U7098 (N_7098,N_4257,N_4950);
nand U7099 (N_7099,N_4683,N_2901);
and U7100 (N_7100,N_4522,N_3036);
or U7101 (N_7101,N_4574,N_3122);
nor U7102 (N_7102,N_3914,N_4018);
or U7103 (N_7103,N_2702,N_3738);
xor U7104 (N_7104,N_2779,N_3177);
and U7105 (N_7105,N_3168,N_3838);
nor U7106 (N_7106,N_2740,N_2879);
xnor U7107 (N_7107,N_3267,N_4008);
nand U7108 (N_7108,N_4729,N_3586);
nor U7109 (N_7109,N_4887,N_3626);
nand U7110 (N_7110,N_3311,N_2912);
or U7111 (N_7111,N_4035,N_3514);
nand U7112 (N_7112,N_2500,N_2675);
or U7113 (N_7113,N_2966,N_4968);
or U7114 (N_7114,N_4258,N_3888);
and U7115 (N_7115,N_2869,N_2729);
and U7116 (N_7116,N_4482,N_3640);
or U7117 (N_7117,N_3248,N_4193);
and U7118 (N_7118,N_4847,N_3760);
or U7119 (N_7119,N_4586,N_3795);
and U7120 (N_7120,N_4078,N_3982);
and U7121 (N_7121,N_4768,N_2678);
or U7122 (N_7122,N_4502,N_4582);
nand U7123 (N_7123,N_4076,N_4992);
and U7124 (N_7124,N_4252,N_3385);
xnor U7125 (N_7125,N_2517,N_3151);
or U7126 (N_7126,N_3554,N_2652);
and U7127 (N_7127,N_3641,N_3653);
nor U7128 (N_7128,N_3794,N_3848);
and U7129 (N_7129,N_4203,N_2561);
xor U7130 (N_7130,N_4057,N_3112);
xnor U7131 (N_7131,N_2535,N_4741);
nand U7132 (N_7132,N_2721,N_2696);
or U7133 (N_7133,N_3982,N_3247);
and U7134 (N_7134,N_2776,N_2688);
and U7135 (N_7135,N_4356,N_2671);
nand U7136 (N_7136,N_4494,N_3998);
and U7137 (N_7137,N_4173,N_4620);
nor U7138 (N_7138,N_3123,N_3818);
or U7139 (N_7139,N_4319,N_4621);
and U7140 (N_7140,N_3666,N_2712);
or U7141 (N_7141,N_4544,N_3207);
nor U7142 (N_7142,N_3788,N_2604);
nand U7143 (N_7143,N_4999,N_3506);
or U7144 (N_7144,N_2973,N_4016);
nand U7145 (N_7145,N_2802,N_3287);
or U7146 (N_7146,N_3175,N_3383);
nor U7147 (N_7147,N_3079,N_4010);
and U7148 (N_7148,N_3619,N_2788);
and U7149 (N_7149,N_3105,N_3412);
xor U7150 (N_7150,N_2728,N_3761);
nand U7151 (N_7151,N_3339,N_3778);
or U7152 (N_7152,N_4725,N_2888);
xor U7153 (N_7153,N_4745,N_3681);
nor U7154 (N_7154,N_4009,N_4283);
xor U7155 (N_7155,N_3462,N_3431);
or U7156 (N_7156,N_3479,N_4011);
xor U7157 (N_7157,N_3527,N_4577);
and U7158 (N_7158,N_4986,N_3868);
nand U7159 (N_7159,N_3549,N_2974);
nand U7160 (N_7160,N_4016,N_4255);
and U7161 (N_7161,N_4142,N_3026);
nand U7162 (N_7162,N_3815,N_4663);
nand U7163 (N_7163,N_3220,N_3145);
nand U7164 (N_7164,N_4002,N_4918);
nand U7165 (N_7165,N_4718,N_4972);
nand U7166 (N_7166,N_3195,N_4891);
nor U7167 (N_7167,N_4854,N_4570);
xor U7168 (N_7168,N_3675,N_3181);
or U7169 (N_7169,N_4405,N_3955);
nand U7170 (N_7170,N_4156,N_4882);
or U7171 (N_7171,N_3224,N_4264);
or U7172 (N_7172,N_2683,N_2812);
or U7173 (N_7173,N_4002,N_4287);
xor U7174 (N_7174,N_3244,N_3087);
xnor U7175 (N_7175,N_3938,N_3194);
xnor U7176 (N_7176,N_4189,N_3047);
and U7177 (N_7177,N_3643,N_3763);
xnor U7178 (N_7178,N_2782,N_4574);
xnor U7179 (N_7179,N_3588,N_2975);
xnor U7180 (N_7180,N_3629,N_4737);
nor U7181 (N_7181,N_3813,N_4274);
or U7182 (N_7182,N_2620,N_4187);
nand U7183 (N_7183,N_4154,N_2994);
nand U7184 (N_7184,N_4496,N_3378);
or U7185 (N_7185,N_4691,N_3776);
xnor U7186 (N_7186,N_3490,N_3036);
and U7187 (N_7187,N_3468,N_3077);
or U7188 (N_7188,N_4682,N_3427);
nand U7189 (N_7189,N_2853,N_3034);
nor U7190 (N_7190,N_3856,N_3759);
nor U7191 (N_7191,N_3194,N_3689);
xnor U7192 (N_7192,N_3957,N_3925);
and U7193 (N_7193,N_3981,N_3205);
nand U7194 (N_7194,N_2847,N_4291);
and U7195 (N_7195,N_4042,N_3675);
and U7196 (N_7196,N_4857,N_4687);
xor U7197 (N_7197,N_2626,N_3406);
or U7198 (N_7198,N_2813,N_2651);
xor U7199 (N_7199,N_3861,N_4063);
and U7200 (N_7200,N_3423,N_3297);
and U7201 (N_7201,N_2524,N_3005);
or U7202 (N_7202,N_2716,N_3174);
nor U7203 (N_7203,N_4018,N_4838);
nand U7204 (N_7204,N_3318,N_3387);
or U7205 (N_7205,N_4873,N_3246);
nor U7206 (N_7206,N_4946,N_3139);
nor U7207 (N_7207,N_4944,N_3676);
xor U7208 (N_7208,N_4951,N_3366);
or U7209 (N_7209,N_3387,N_3422);
and U7210 (N_7210,N_4838,N_4503);
and U7211 (N_7211,N_4720,N_4957);
nand U7212 (N_7212,N_3209,N_3682);
or U7213 (N_7213,N_4303,N_2568);
and U7214 (N_7214,N_3091,N_2995);
nand U7215 (N_7215,N_3507,N_3806);
xor U7216 (N_7216,N_4028,N_4734);
and U7217 (N_7217,N_4570,N_2797);
and U7218 (N_7218,N_4294,N_4931);
or U7219 (N_7219,N_3580,N_3145);
xor U7220 (N_7220,N_2965,N_4673);
nor U7221 (N_7221,N_4563,N_3827);
or U7222 (N_7222,N_4015,N_4363);
and U7223 (N_7223,N_2781,N_4401);
or U7224 (N_7224,N_4117,N_4766);
nand U7225 (N_7225,N_2611,N_2795);
nor U7226 (N_7226,N_4458,N_3318);
and U7227 (N_7227,N_4961,N_4298);
nor U7228 (N_7228,N_3813,N_2567);
nor U7229 (N_7229,N_2719,N_3303);
nor U7230 (N_7230,N_4963,N_4532);
xor U7231 (N_7231,N_3784,N_4739);
nor U7232 (N_7232,N_2829,N_4389);
and U7233 (N_7233,N_4275,N_3450);
nand U7234 (N_7234,N_4582,N_3980);
or U7235 (N_7235,N_4038,N_3053);
nand U7236 (N_7236,N_3482,N_3270);
xor U7237 (N_7237,N_4689,N_2630);
or U7238 (N_7238,N_4594,N_2911);
nor U7239 (N_7239,N_4844,N_4040);
nand U7240 (N_7240,N_4300,N_3123);
or U7241 (N_7241,N_3114,N_3515);
nand U7242 (N_7242,N_3983,N_4278);
and U7243 (N_7243,N_2813,N_3200);
nor U7244 (N_7244,N_3695,N_2871);
and U7245 (N_7245,N_2927,N_4041);
xnor U7246 (N_7246,N_2584,N_4667);
or U7247 (N_7247,N_3504,N_4606);
nand U7248 (N_7248,N_4508,N_3056);
xnor U7249 (N_7249,N_4391,N_4047);
or U7250 (N_7250,N_3212,N_4289);
or U7251 (N_7251,N_3671,N_3740);
nor U7252 (N_7252,N_4728,N_2665);
and U7253 (N_7253,N_4474,N_3307);
and U7254 (N_7254,N_4250,N_3006);
or U7255 (N_7255,N_3512,N_3846);
nor U7256 (N_7256,N_3005,N_3144);
nor U7257 (N_7257,N_2559,N_3408);
nand U7258 (N_7258,N_3080,N_2716);
xnor U7259 (N_7259,N_2863,N_3286);
xnor U7260 (N_7260,N_3137,N_4194);
and U7261 (N_7261,N_3393,N_4478);
nor U7262 (N_7262,N_3594,N_4293);
nand U7263 (N_7263,N_3298,N_3393);
nand U7264 (N_7264,N_2605,N_2769);
or U7265 (N_7265,N_3972,N_4533);
nand U7266 (N_7266,N_4451,N_4640);
nor U7267 (N_7267,N_3794,N_4091);
xnor U7268 (N_7268,N_3056,N_3341);
xor U7269 (N_7269,N_2658,N_3865);
nand U7270 (N_7270,N_4414,N_4564);
nor U7271 (N_7271,N_4742,N_2786);
xnor U7272 (N_7272,N_2569,N_2843);
nor U7273 (N_7273,N_2899,N_2621);
nand U7274 (N_7274,N_4340,N_4633);
xor U7275 (N_7275,N_3022,N_4083);
xnor U7276 (N_7276,N_4149,N_3583);
and U7277 (N_7277,N_4415,N_4541);
and U7278 (N_7278,N_3371,N_4962);
and U7279 (N_7279,N_4942,N_4590);
and U7280 (N_7280,N_4923,N_3340);
and U7281 (N_7281,N_3737,N_4959);
nand U7282 (N_7282,N_2913,N_3216);
and U7283 (N_7283,N_2515,N_3806);
nor U7284 (N_7284,N_3018,N_4523);
or U7285 (N_7285,N_4349,N_4061);
and U7286 (N_7286,N_4427,N_4291);
nor U7287 (N_7287,N_3788,N_4580);
and U7288 (N_7288,N_2815,N_3616);
and U7289 (N_7289,N_3277,N_2634);
and U7290 (N_7290,N_2611,N_3389);
nand U7291 (N_7291,N_2589,N_3345);
and U7292 (N_7292,N_2796,N_4589);
and U7293 (N_7293,N_4370,N_4077);
nand U7294 (N_7294,N_3266,N_4070);
nor U7295 (N_7295,N_2886,N_2965);
nor U7296 (N_7296,N_3926,N_4015);
nor U7297 (N_7297,N_4148,N_4375);
nand U7298 (N_7298,N_2511,N_3634);
and U7299 (N_7299,N_3243,N_4760);
xor U7300 (N_7300,N_4671,N_4630);
or U7301 (N_7301,N_4441,N_3348);
xor U7302 (N_7302,N_3920,N_4041);
nand U7303 (N_7303,N_4823,N_2645);
or U7304 (N_7304,N_4144,N_4759);
xnor U7305 (N_7305,N_2513,N_4232);
xnor U7306 (N_7306,N_2500,N_3654);
and U7307 (N_7307,N_4728,N_2642);
or U7308 (N_7308,N_4250,N_3435);
or U7309 (N_7309,N_2879,N_3902);
or U7310 (N_7310,N_3943,N_4438);
xor U7311 (N_7311,N_4156,N_2888);
and U7312 (N_7312,N_4325,N_3906);
and U7313 (N_7313,N_2798,N_3314);
xnor U7314 (N_7314,N_3914,N_3735);
nor U7315 (N_7315,N_4082,N_3478);
xnor U7316 (N_7316,N_3212,N_4460);
and U7317 (N_7317,N_4168,N_2953);
nand U7318 (N_7318,N_4208,N_2685);
nor U7319 (N_7319,N_4442,N_2831);
xnor U7320 (N_7320,N_3941,N_2847);
nor U7321 (N_7321,N_4519,N_4709);
nand U7322 (N_7322,N_3716,N_4646);
nor U7323 (N_7323,N_4586,N_4169);
xor U7324 (N_7324,N_2895,N_3924);
nor U7325 (N_7325,N_2683,N_4100);
nor U7326 (N_7326,N_3375,N_4647);
xor U7327 (N_7327,N_3920,N_3282);
and U7328 (N_7328,N_3448,N_4167);
xnor U7329 (N_7329,N_4776,N_4409);
nand U7330 (N_7330,N_2562,N_4781);
and U7331 (N_7331,N_3983,N_4652);
nand U7332 (N_7332,N_3636,N_4762);
nor U7333 (N_7333,N_3955,N_4929);
xor U7334 (N_7334,N_2539,N_4775);
and U7335 (N_7335,N_2627,N_3807);
and U7336 (N_7336,N_3096,N_3416);
xnor U7337 (N_7337,N_3159,N_3914);
nand U7338 (N_7338,N_4994,N_2697);
xnor U7339 (N_7339,N_3162,N_4461);
and U7340 (N_7340,N_4912,N_2793);
xnor U7341 (N_7341,N_4397,N_4208);
or U7342 (N_7342,N_2919,N_4914);
or U7343 (N_7343,N_3914,N_3046);
nor U7344 (N_7344,N_3067,N_2896);
nand U7345 (N_7345,N_4009,N_3946);
xnor U7346 (N_7346,N_4825,N_3454);
nand U7347 (N_7347,N_4347,N_4546);
nor U7348 (N_7348,N_4756,N_2670);
xor U7349 (N_7349,N_3522,N_3504);
or U7350 (N_7350,N_3303,N_4521);
or U7351 (N_7351,N_4836,N_3495);
nor U7352 (N_7352,N_3691,N_4437);
nand U7353 (N_7353,N_2543,N_2861);
xor U7354 (N_7354,N_2964,N_4932);
and U7355 (N_7355,N_4231,N_4166);
and U7356 (N_7356,N_4492,N_2735);
nor U7357 (N_7357,N_3868,N_3540);
or U7358 (N_7358,N_3651,N_3111);
xnor U7359 (N_7359,N_3875,N_4375);
or U7360 (N_7360,N_4960,N_3526);
nand U7361 (N_7361,N_3364,N_4067);
and U7362 (N_7362,N_4798,N_3612);
nor U7363 (N_7363,N_4935,N_3626);
xor U7364 (N_7364,N_4819,N_4708);
and U7365 (N_7365,N_2864,N_2659);
nor U7366 (N_7366,N_3826,N_4291);
and U7367 (N_7367,N_4018,N_2584);
xnor U7368 (N_7368,N_4689,N_4234);
or U7369 (N_7369,N_2523,N_4862);
and U7370 (N_7370,N_3139,N_4506);
nor U7371 (N_7371,N_2769,N_2844);
xor U7372 (N_7372,N_4663,N_2640);
xnor U7373 (N_7373,N_3775,N_4664);
or U7374 (N_7374,N_3166,N_2784);
nor U7375 (N_7375,N_4534,N_4125);
nand U7376 (N_7376,N_3321,N_3897);
or U7377 (N_7377,N_2694,N_3868);
nor U7378 (N_7378,N_3748,N_4032);
xnor U7379 (N_7379,N_3690,N_4248);
or U7380 (N_7380,N_4601,N_3043);
and U7381 (N_7381,N_4171,N_4394);
xor U7382 (N_7382,N_4214,N_3995);
nor U7383 (N_7383,N_3840,N_3514);
or U7384 (N_7384,N_3989,N_4906);
xor U7385 (N_7385,N_2889,N_3383);
nor U7386 (N_7386,N_4866,N_3058);
or U7387 (N_7387,N_4827,N_3960);
nor U7388 (N_7388,N_2753,N_2620);
nor U7389 (N_7389,N_2947,N_3859);
or U7390 (N_7390,N_3075,N_4935);
xnor U7391 (N_7391,N_3990,N_3238);
or U7392 (N_7392,N_4196,N_3131);
and U7393 (N_7393,N_2861,N_3231);
or U7394 (N_7394,N_3744,N_3166);
or U7395 (N_7395,N_2885,N_4998);
and U7396 (N_7396,N_2859,N_3695);
and U7397 (N_7397,N_2658,N_4048);
and U7398 (N_7398,N_4096,N_3554);
xnor U7399 (N_7399,N_3374,N_3710);
xor U7400 (N_7400,N_3595,N_4782);
nand U7401 (N_7401,N_4104,N_2839);
and U7402 (N_7402,N_3736,N_2681);
or U7403 (N_7403,N_4784,N_4966);
nor U7404 (N_7404,N_2947,N_4047);
nor U7405 (N_7405,N_4426,N_3422);
and U7406 (N_7406,N_4546,N_3773);
or U7407 (N_7407,N_3639,N_4637);
or U7408 (N_7408,N_3152,N_4795);
nand U7409 (N_7409,N_4541,N_2785);
nand U7410 (N_7410,N_2889,N_4940);
or U7411 (N_7411,N_3195,N_3920);
and U7412 (N_7412,N_3812,N_3771);
or U7413 (N_7413,N_3533,N_3147);
nand U7414 (N_7414,N_3231,N_2794);
or U7415 (N_7415,N_2977,N_3381);
nand U7416 (N_7416,N_4482,N_3656);
or U7417 (N_7417,N_2756,N_3425);
and U7418 (N_7418,N_4345,N_3471);
nor U7419 (N_7419,N_4296,N_4021);
and U7420 (N_7420,N_4074,N_4830);
nor U7421 (N_7421,N_4094,N_4620);
xnor U7422 (N_7422,N_2764,N_2630);
nor U7423 (N_7423,N_3887,N_3412);
and U7424 (N_7424,N_2757,N_3725);
nand U7425 (N_7425,N_4166,N_2588);
and U7426 (N_7426,N_4888,N_3830);
nand U7427 (N_7427,N_2511,N_4000);
nor U7428 (N_7428,N_3747,N_2775);
xnor U7429 (N_7429,N_3836,N_4578);
nand U7430 (N_7430,N_4963,N_2982);
and U7431 (N_7431,N_4991,N_3294);
and U7432 (N_7432,N_2638,N_3517);
xnor U7433 (N_7433,N_4057,N_4177);
nand U7434 (N_7434,N_3402,N_2883);
and U7435 (N_7435,N_3735,N_2704);
or U7436 (N_7436,N_3553,N_4670);
and U7437 (N_7437,N_3276,N_4793);
nor U7438 (N_7438,N_3611,N_3836);
xor U7439 (N_7439,N_3308,N_4530);
nand U7440 (N_7440,N_4864,N_3234);
nor U7441 (N_7441,N_2783,N_3434);
and U7442 (N_7442,N_4342,N_4969);
or U7443 (N_7443,N_3182,N_2848);
or U7444 (N_7444,N_4275,N_4592);
or U7445 (N_7445,N_3595,N_3828);
nor U7446 (N_7446,N_2589,N_3153);
and U7447 (N_7447,N_3004,N_2646);
xnor U7448 (N_7448,N_4075,N_3385);
xnor U7449 (N_7449,N_3078,N_4340);
nor U7450 (N_7450,N_4865,N_3126);
nand U7451 (N_7451,N_3735,N_4423);
nor U7452 (N_7452,N_3784,N_3469);
xor U7453 (N_7453,N_4113,N_4873);
nor U7454 (N_7454,N_4007,N_3149);
or U7455 (N_7455,N_3719,N_4927);
xnor U7456 (N_7456,N_3046,N_3891);
nor U7457 (N_7457,N_3385,N_4529);
or U7458 (N_7458,N_2636,N_2655);
xor U7459 (N_7459,N_4322,N_3796);
and U7460 (N_7460,N_3591,N_4701);
nor U7461 (N_7461,N_3367,N_3595);
nand U7462 (N_7462,N_2811,N_4291);
nor U7463 (N_7463,N_4809,N_4472);
and U7464 (N_7464,N_3145,N_3646);
or U7465 (N_7465,N_3301,N_2968);
nor U7466 (N_7466,N_3998,N_3680);
and U7467 (N_7467,N_3953,N_4004);
nor U7468 (N_7468,N_4938,N_3921);
xor U7469 (N_7469,N_3153,N_4892);
xor U7470 (N_7470,N_3300,N_3631);
nand U7471 (N_7471,N_2612,N_2819);
and U7472 (N_7472,N_4061,N_4272);
xnor U7473 (N_7473,N_4036,N_4714);
nor U7474 (N_7474,N_4251,N_2765);
nand U7475 (N_7475,N_3655,N_3277);
nor U7476 (N_7476,N_3584,N_4296);
or U7477 (N_7477,N_4366,N_4248);
nor U7478 (N_7478,N_4914,N_3093);
nand U7479 (N_7479,N_4029,N_3707);
and U7480 (N_7480,N_3339,N_4288);
or U7481 (N_7481,N_3571,N_4271);
or U7482 (N_7482,N_3720,N_4867);
nor U7483 (N_7483,N_4867,N_2573);
nor U7484 (N_7484,N_4334,N_3137);
or U7485 (N_7485,N_3929,N_3750);
nor U7486 (N_7486,N_3592,N_3178);
nand U7487 (N_7487,N_2781,N_4201);
xor U7488 (N_7488,N_4092,N_4119);
xnor U7489 (N_7489,N_3994,N_3449);
nand U7490 (N_7490,N_3235,N_3063);
and U7491 (N_7491,N_4378,N_3394);
nor U7492 (N_7492,N_4922,N_3730);
xnor U7493 (N_7493,N_4890,N_4693);
nor U7494 (N_7494,N_3185,N_2877);
and U7495 (N_7495,N_3162,N_3868);
or U7496 (N_7496,N_3597,N_3734);
and U7497 (N_7497,N_4894,N_4461);
xnor U7498 (N_7498,N_3297,N_3188);
and U7499 (N_7499,N_4641,N_4454);
xnor U7500 (N_7500,N_6998,N_5409);
nand U7501 (N_7501,N_7418,N_5797);
and U7502 (N_7502,N_6172,N_5402);
xnor U7503 (N_7503,N_6057,N_7033);
nand U7504 (N_7504,N_6807,N_5931);
xor U7505 (N_7505,N_6498,N_5668);
nor U7506 (N_7506,N_7448,N_7120);
nand U7507 (N_7507,N_7248,N_5353);
and U7508 (N_7508,N_7353,N_5433);
xor U7509 (N_7509,N_6175,N_5026);
nor U7510 (N_7510,N_5669,N_7491);
or U7511 (N_7511,N_5348,N_6647);
and U7512 (N_7512,N_5974,N_7151);
or U7513 (N_7513,N_5335,N_7222);
xor U7514 (N_7514,N_6126,N_6889);
xor U7515 (N_7515,N_6244,N_5986);
or U7516 (N_7516,N_7417,N_6742);
xnor U7517 (N_7517,N_7457,N_6664);
and U7518 (N_7518,N_5435,N_6623);
or U7519 (N_7519,N_7066,N_5852);
xnor U7520 (N_7520,N_5819,N_6718);
or U7521 (N_7521,N_6363,N_5473);
xor U7522 (N_7522,N_5236,N_5599);
or U7523 (N_7523,N_6227,N_5573);
nor U7524 (N_7524,N_7153,N_6088);
nor U7525 (N_7525,N_5648,N_6365);
or U7526 (N_7526,N_6787,N_6333);
nand U7527 (N_7527,N_5781,N_5924);
and U7528 (N_7528,N_5664,N_5954);
xor U7529 (N_7529,N_6453,N_6967);
and U7530 (N_7530,N_6912,N_6938);
nand U7531 (N_7531,N_5037,N_5138);
xor U7532 (N_7532,N_6235,N_6286);
or U7533 (N_7533,N_5084,N_5719);
or U7534 (N_7534,N_7069,N_5831);
nor U7535 (N_7535,N_7133,N_6338);
and U7536 (N_7536,N_7005,N_5491);
nand U7537 (N_7537,N_7013,N_5330);
xnor U7538 (N_7538,N_5126,N_7402);
xor U7539 (N_7539,N_6595,N_5210);
or U7540 (N_7540,N_5653,N_6193);
nand U7541 (N_7541,N_5841,N_5769);
xnor U7542 (N_7542,N_7320,N_5096);
and U7543 (N_7543,N_7115,N_7302);
and U7544 (N_7544,N_6852,N_6467);
or U7545 (N_7545,N_5703,N_6234);
nor U7546 (N_7546,N_7392,N_5893);
xnor U7547 (N_7547,N_6368,N_7297);
nand U7548 (N_7548,N_5298,N_7056);
nand U7549 (N_7549,N_5321,N_6408);
nand U7550 (N_7550,N_5522,N_5608);
xnor U7551 (N_7551,N_5293,N_5625);
nor U7552 (N_7552,N_5890,N_7160);
and U7553 (N_7553,N_7057,N_7458);
nor U7554 (N_7554,N_5067,N_5045);
nand U7555 (N_7555,N_7312,N_5981);
and U7556 (N_7556,N_7241,N_5100);
and U7557 (N_7557,N_5665,N_5802);
and U7558 (N_7558,N_6135,N_6853);
nor U7559 (N_7559,N_5169,N_6715);
and U7560 (N_7560,N_7233,N_6307);
or U7561 (N_7561,N_5405,N_7028);
and U7562 (N_7562,N_6671,N_6560);
nor U7563 (N_7563,N_6434,N_6061);
or U7564 (N_7564,N_6021,N_5289);
nor U7565 (N_7565,N_5271,N_5998);
xnor U7566 (N_7566,N_5763,N_6496);
and U7567 (N_7567,N_5922,N_7373);
xor U7568 (N_7568,N_5206,N_5844);
nand U7569 (N_7569,N_5675,N_5952);
xor U7570 (N_7570,N_7391,N_6031);
and U7571 (N_7571,N_5810,N_6051);
and U7572 (N_7572,N_7067,N_5276);
or U7573 (N_7573,N_5883,N_5116);
or U7574 (N_7574,N_7189,N_6890);
nand U7575 (N_7575,N_6200,N_6656);
xnor U7576 (N_7576,N_5311,N_6452);
or U7577 (N_7577,N_6440,N_6747);
xor U7578 (N_7578,N_7346,N_6955);
xor U7579 (N_7579,N_5315,N_6778);
or U7580 (N_7580,N_6101,N_6373);
xor U7581 (N_7581,N_6987,N_7243);
nor U7582 (N_7582,N_5550,N_5476);
or U7583 (N_7583,N_6585,N_6424);
or U7584 (N_7584,N_5219,N_5520);
xnor U7585 (N_7585,N_6500,N_6661);
xor U7586 (N_7586,N_5278,N_5261);
nand U7587 (N_7587,N_5707,N_6737);
nor U7588 (N_7588,N_6525,N_7215);
or U7589 (N_7589,N_6002,N_7226);
xor U7590 (N_7590,N_7105,N_5006);
and U7591 (N_7591,N_6753,N_7106);
and U7592 (N_7592,N_7228,N_7411);
nand U7593 (N_7593,N_6176,N_6809);
nand U7594 (N_7594,N_6136,N_5149);
or U7595 (N_7595,N_5495,N_6226);
xor U7596 (N_7596,N_6161,N_6866);
nor U7597 (N_7597,N_5065,N_7250);
nor U7598 (N_7598,N_5372,N_7253);
xor U7599 (N_7599,N_7044,N_7092);
nor U7600 (N_7600,N_6102,N_6845);
nor U7601 (N_7601,N_5848,N_6120);
and U7602 (N_7602,N_6055,N_7301);
nand U7603 (N_7603,N_5381,N_6382);
or U7604 (N_7604,N_7239,N_5422);
nor U7605 (N_7605,N_6924,N_5766);
and U7606 (N_7606,N_6377,N_6682);
xor U7607 (N_7607,N_6963,N_5316);
and U7608 (N_7608,N_6904,N_6013);
nand U7609 (N_7609,N_5756,N_6222);
nor U7610 (N_7610,N_5263,N_6763);
and U7611 (N_7611,N_7264,N_5558);
nor U7612 (N_7612,N_5077,N_6238);
xnor U7613 (N_7613,N_6838,N_5370);
and U7614 (N_7614,N_7355,N_5387);
nor U7615 (N_7615,N_6374,N_5367);
nand U7616 (N_7616,N_6961,N_6230);
or U7617 (N_7617,N_5907,N_5089);
and U7618 (N_7618,N_5184,N_6393);
nor U7619 (N_7619,N_6037,N_7280);
xor U7620 (N_7620,N_7366,N_7370);
and U7621 (N_7621,N_6203,N_6545);
nor U7622 (N_7622,N_7313,N_5812);
nor U7623 (N_7623,N_6684,N_7277);
or U7624 (N_7624,N_5297,N_6881);
nand U7625 (N_7625,N_5286,N_6009);
and U7626 (N_7626,N_7481,N_5328);
nor U7627 (N_7627,N_5865,N_7337);
xor U7628 (N_7628,N_6877,N_6299);
nand U7629 (N_7629,N_5317,N_6976);
nor U7630 (N_7630,N_5878,N_5139);
xor U7631 (N_7631,N_5171,N_7388);
nand U7632 (N_7632,N_5785,N_7210);
nand U7633 (N_7633,N_7142,N_5343);
nand U7634 (N_7634,N_5765,N_5566);
or U7635 (N_7635,N_6953,N_6336);
nor U7636 (N_7636,N_7180,N_6237);
or U7637 (N_7637,N_6131,N_6911);
or U7638 (N_7638,N_5512,N_6156);
or U7639 (N_7639,N_5109,N_7156);
and U7640 (N_7640,N_6649,N_5754);
nand U7641 (N_7641,N_5136,N_7444);
or U7642 (N_7642,N_5121,N_6644);
or U7643 (N_7643,N_5203,N_5780);
or U7644 (N_7644,N_6068,N_5811);
nand U7645 (N_7645,N_7109,N_6287);
or U7646 (N_7646,N_6533,N_5418);
nor U7647 (N_7647,N_5031,N_6815);
or U7648 (N_7648,N_5061,N_6657);
and U7649 (N_7649,N_7000,N_5966);
nor U7650 (N_7650,N_6069,N_7242);
nor U7651 (N_7651,N_5043,N_6213);
nand U7652 (N_7652,N_6125,N_5284);
xor U7653 (N_7653,N_6750,N_7255);
xnor U7654 (N_7654,N_5245,N_5038);
or U7655 (N_7655,N_7147,N_6015);
nor U7656 (N_7656,N_5420,N_5634);
xnor U7657 (N_7657,N_5611,N_6704);
xor U7658 (N_7658,N_5997,N_5521);
or U7659 (N_7659,N_6764,N_5985);
nor U7660 (N_7660,N_6908,N_6048);
and U7661 (N_7661,N_5709,N_6501);
and U7662 (N_7662,N_5972,N_5723);
xor U7663 (N_7663,N_6642,N_6695);
nor U7664 (N_7664,N_6876,N_6354);
nand U7665 (N_7665,N_6872,N_5630);
and U7666 (N_7666,N_6306,N_5487);
and U7667 (N_7667,N_5104,N_7185);
and U7668 (N_7668,N_5478,N_5228);
and U7669 (N_7669,N_6942,N_5440);
or U7670 (N_7670,N_6401,N_5517);
nor U7671 (N_7671,N_7045,N_7084);
nand U7672 (N_7672,N_6367,N_7178);
or U7673 (N_7673,N_5807,N_7341);
and U7674 (N_7674,N_7298,N_6384);
or U7675 (N_7675,N_7083,N_7177);
nand U7676 (N_7676,N_6993,N_6793);
xnor U7677 (N_7677,N_5281,N_5073);
nand U7678 (N_7678,N_6552,N_6786);
or U7679 (N_7679,N_6956,N_6670);
or U7680 (N_7680,N_6794,N_5718);
nand U7681 (N_7681,N_5386,N_6597);
nand U7682 (N_7682,N_5357,N_5578);
nor U7683 (N_7683,N_5783,N_7303);
and U7684 (N_7684,N_6263,N_7082);
nand U7685 (N_7685,N_6350,N_5205);
xnor U7686 (N_7686,N_5078,N_5469);
nor U7687 (N_7687,N_6006,N_6951);
xor U7688 (N_7688,N_6814,N_7051);
and U7689 (N_7689,N_5744,N_6492);
or U7690 (N_7690,N_6047,N_6907);
or U7691 (N_7691,N_6471,N_7111);
nor U7692 (N_7692,N_5933,N_6933);
nor U7693 (N_7693,N_6514,N_6518);
and U7694 (N_7694,N_6790,N_6611);
or U7695 (N_7695,N_7382,N_5294);
nand U7696 (N_7696,N_6673,N_5074);
nor U7697 (N_7697,N_7441,N_5150);
and U7698 (N_7698,N_6861,N_5361);
nand U7699 (N_7699,N_5932,N_7251);
nor U7700 (N_7700,N_6157,N_6271);
nand U7701 (N_7701,N_5870,N_5364);
and U7702 (N_7702,N_5671,N_6108);
or U7703 (N_7703,N_6683,N_7396);
xnor U7704 (N_7704,N_5235,N_7181);
xnor U7705 (N_7705,N_6667,N_5696);
xnor U7706 (N_7706,N_5523,N_5855);
xor U7707 (N_7707,N_6112,N_5773);
and U7708 (N_7708,N_5876,N_6968);
xnor U7709 (N_7709,N_7062,N_7318);
xor U7710 (N_7710,N_6537,N_5181);
or U7711 (N_7711,N_6544,N_6085);
and U7712 (N_7712,N_6023,N_6969);
nand U7713 (N_7713,N_6940,N_6189);
xor U7714 (N_7714,N_7347,N_5208);
nand U7715 (N_7715,N_7237,N_5246);
nor U7716 (N_7716,N_5410,N_5708);
nor U7717 (N_7717,N_5334,N_6334);
nand U7718 (N_7718,N_7221,N_6732);
and U7719 (N_7719,N_5768,N_6302);
nor U7720 (N_7720,N_7383,N_5660);
nor U7721 (N_7721,N_6736,N_5000);
nand U7722 (N_7722,N_6739,N_5864);
nand U7723 (N_7723,N_6729,N_6168);
or U7724 (N_7724,N_5651,N_6705);
nor U7725 (N_7725,N_6685,N_6045);
xor U7726 (N_7726,N_6455,N_5467);
xnor U7727 (N_7727,N_5501,N_5151);
nand U7728 (N_7728,N_6358,N_6818);
and U7729 (N_7729,N_7266,N_5331);
and U7730 (N_7730,N_6550,N_6971);
nor U7731 (N_7731,N_5157,N_5107);
nor U7732 (N_7732,N_5302,N_6724);
xnor U7733 (N_7733,N_5720,N_7128);
nor U7734 (N_7734,N_5982,N_5818);
and U7735 (N_7735,N_6843,N_5993);
or U7736 (N_7736,N_5882,N_5048);
nor U7737 (N_7737,N_5590,N_6910);
or U7738 (N_7738,N_6355,N_7398);
and U7739 (N_7739,N_5698,N_5141);
and U7740 (N_7740,N_5195,N_6551);
nand U7741 (N_7741,N_6081,N_5592);
nand U7742 (N_7742,N_6746,N_6318);
or U7743 (N_7743,N_6655,N_7283);
and U7744 (N_7744,N_6127,N_5706);
nor U7745 (N_7745,N_5062,N_6796);
and U7746 (N_7746,N_6722,N_5233);
xnor U7747 (N_7747,N_5212,N_5484);
or U7748 (N_7748,N_6592,N_7342);
and U7749 (N_7749,N_6208,N_6110);
nor U7750 (N_7750,N_7421,N_5240);
and U7751 (N_7751,N_5808,N_5329);
nor U7752 (N_7752,N_5761,N_6160);
and U7753 (N_7753,N_6308,N_6205);
and U7754 (N_7754,N_5684,N_5693);
and U7755 (N_7755,N_5979,N_5034);
xnor U7756 (N_7756,N_6282,N_5951);
nand U7757 (N_7757,N_5401,N_5490);
or U7758 (N_7758,N_5688,N_5099);
nor U7759 (N_7759,N_6152,N_7073);
nand U7760 (N_7760,N_7438,N_6485);
xnor U7761 (N_7761,N_5486,N_5724);
or U7762 (N_7762,N_6144,N_5631);
or U7763 (N_7763,N_7480,N_5231);
nor U7764 (N_7764,N_5640,N_6844);
and U7765 (N_7765,N_6840,N_6820);
nor U7766 (N_7766,N_7261,N_6666);
nand U7767 (N_7767,N_6425,N_5414);
and U7768 (N_7768,N_7247,N_6507);
and U7769 (N_7769,N_5362,N_7324);
and U7770 (N_7770,N_7208,N_7344);
nor U7771 (N_7771,N_5510,N_5462);
and U7772 (N_7772,N_5341,N_5003);
or U7773 (N_7773,N_6948,N_5249);
xor U7774 (N_7774,N_6626,N_5570);
and U7775 (N_7775,N_5359,N_7489);
nand U7776 (N_7776,N_6030,N_5344);
or U7777 (N_7777,N_7350,N_5845);
or U7778 (N_7778,N_7220,N_6313);
nand U7779 (N_7779,N_7371,N_5589);
nand U7780 (N_7780,N_6000,N_5862);
nor U7781 (N_7781,N_6719,N_5498);
and U7782 (N_7782,N_7424,N_5040);
and U7783 (N_7783,N_5185,N_7401);
or U7784 (N_7784,N_5962,N_6224);
nand U7785 (N_7785,N_7459,N_5324);
and U7786 (N_7786,N_7130,N_7478);
or U7787 (N_7787,N_6254,N_6099);
or U7788 (N_7788,N_7087,N_7245);
and U7789 (N_7789,N_5733,N_5291);
and U7790 (N_7790,N_6072,N_6687);
xnor U7791 (N_7791,N_6219,N_7258);
and U7792 (N_7792,N_6008,N_6730);
and U7793 (N_7793,N_7482,N_6782);
or U7794 (N_7794,N_6417,N_6605);
nand U7795 (N_7795,N_5775,N_6476);
xor U7796 (N_7796,N_6097,N_6926);
or U7797 (N_7797,N_5180,N_6232);
and U7798 (N_7798,N_6138,N_5853);
nor U7799 (N_7799,N_5957,N_5729);
nand U7800 (N_7800,N_7123,N_7148);
nand U7801 (N_7801,N_7016,N_7462);
xnor U7802 (N_7802,N_5969,N_5252);
or U7803 (N_7803,N_6770,N_5135);
nand U7804 (N_7804,N_5223,N_6331);
and U7805 (N_7805,N_6209,N_7206);
or U7806 (N_7806,N_7168,N_6115);
and U7807 (N_7807,N_7121,N_5944);
xor U7808 (N_7808,N_6608,N_6241);
nor U7809 (N_7809,N_5854,N_5105);
nand U7810 (N_7810,N_7385,N_5977);
xnor U7811 (N_7811,N_6752,N_6721);
or U7812 (N_7812,N_7081,N_6280);
nor U7813 (N_7813,N_5187,N_6154);
nor U7814 (N_7814,N_6491,N_5567);
xnor U7815 (N_7815,N_5055,N_7452);
and U7816 (N_7816,N_5145,N_7024);
nor U7817 (N_7817,N_5505,N_5943);
or U7818 (N_7818,N_6053,N_6916);
xor U7819 (N_7819,N_7175,N_5909);
nor U7820 (N_7820,N_5429,N_5008);
nor U7821 (N_7821,N_6821,N_5477);
nand U7822 (N_7822,N_7381,N_6974);
nand U7823 (N_7823,N_5304,N_6837);
nor U7824 (N_7824,N_5452,N_6615);
and U7825 (N_7825,N_6091,N_6040);
and U7826 (N_7826,N_6356,N_6530);
nor U7827 (N_7827,N_7187,N_5027);
and U7828 (N_7828,N_6247,N_5166);
nand U7829 (N_7829,N_6293,N_5148);
nand U7830 (N_7830,N_6634,N_7360);
and U7831 (N_7831,N_5011,N_6986);
nor U7832 (N_7832,N_6033,N_6012);
nor U7833 (N_7833,N_7377,N_5287);
or U7834 (N_7834,N_5224,N_6631);
nand U7835 (N_7835,N_6599,N_7466);
or U7836 (N_7836,N_6195,N_7488);
nor U7837 (N_7837,N_5313,N_5253);
nand U7838 (N_7838,N_5118,N_5991);
nand U7839 (N_7839,N_7223,N_5595);
or U7840 (N_7840,N_5774,N_5356);
or U7841 (N_7841,N_5103,N_5295);
or U7842 (N_7842,N_6950,N_6410);
or U7843 (N_7843,N_5757,N_5413);
nor U7844 (N_7844,N_6409,N_5533);
and U7845 (N_7845,N_7289,N_7116);
xor U7846 (N_7846,N_5175,N_6320);
or U7847 (N_7847,N_5963,N_7330);
and U7848 (N_7848,N_5973,N_6726);
and U7849 (N_7849,N_5778,N_6576);
nor U7850 (N_7850,N_5619,N_7329);
nor U7851 (N_7851,N_6166,N_5274);
and U7852 (N_7852,N_6577,N_5308);
nor U7853 (N_7853,N_6475,N_5004);
nand U7854 (N_7854,N_5441,N_7477);
or U7855 (N_7855,N_6979,N_7412);
xor U7856 (N_7856,N_6429,N_6830);
or U7857 (N_7857,N_5872,N_5090);
xor U7858 (N_7858,N_5913,N_5389);
nand U7859 (N_7859,N_5444,N_7122);
nor U7860 (N_7860,N_6495,N_5900);
nand U7861 (N_7861,N_6992,N_6964);
and U7862 (N_7862,N_5456,N_7030);
xor U7863 (N_7863,N_6645,N_5525);
nor U7864 (N_7864,N_6810,N_6621);
nand U7865 (N_7865,N_5758,N_6194);
or U7866 (N_7866,N_6484,N_6878);
xor U7867 (N_7867,N_7173,N_6079);
nor U7868 (N_7868,N_6106,N_5489);
xnor U7869 (N_7869,N_6819,N_6936);
and U7870 (N_7870,N_5543,N_6357);
nand U7871 (N_7871,N_5574,N_6801);
or U7872 (N_7872,N_6388,N_6415);
or U7873 (N_7873,N_6329,N_6442);
and U7874 (N_7874,N_7157,N_5835);
and U7875 (N_7875,N_6935,N_5735);
or U7876 (N_7876,N_6311,N_5687);
xnor U7877 (N_7877,N_5244,N_6283);
or U7878 (N_7878,N_5504,N_6927);
and U7879 (N_7879,N_6113,N_5102);
nor U7880 (N_7880,N_7027,N_5094);
nor U7881 (N_7881,N_5562,N_5580);
or U7882 (N_7882,N_6489,N_5010);
nor U7883 (N_7883,N_5283,N_5247);
nor U7884 (N_7884,N_5686,N_7420);
nand U7885 (N_7885,N_6740,N_6481);
or U7886 (N_7886,N_6019,N_6301);
nor U7887 (N_7887,N_5929,N_7335);
or U7888 (N_7888,N_5397,N_6180);
or U7889 (N_7889,N_6902,N_5650);
xor U7890 (N_7890,N_6882,N_6930);
nand U7891 (N_7891,N_6188,N_5358);
or U7892 (N_7892,N_7091,N_5955);
nor U7893 (N_7893,N_6458,N_7055);
nor U7894 (N_7894,N_6231,N_6352);
nor U7895 (N_7895,N_5447,N_7049);
or U7896 (N_7896,N_7046,N_5170);
nand U7897 (N_7897,N_5602,N_7202);
nor U7898 (N_7898,N_6825,N_7099);
and U7899 (N_7899,N_5494,N_6353);
or U7900 (N_7900,N_6210,N_5548);
nand U7901 (N_7901,N_5920,N_6223);
or U7902 (N_7902,N_6708,N_6400);
nor U7903 (N_7903,N_6733,N_6182);
and U7904 (N_7904,N_5927,N_5838);
or U7905 (N_7905,N_5647,N_6038);
xor U7906 (N_7906,N_6562,N_5956);
or U7907 (N_7907,N_5753,N_6829);
and U7908 (N_7908,N_6349,N_7378);
or U7909 (N_7909,N_6319,N_7025);
and U7910 (N_7910,N_5174,N_6462);
and U7911 (N_7911,N_5577,N_6398);
nand U7912 (N_7912,N_7204,N_6433);
nor U7913 (N_7913,N_7135,N_7119);
nand U7914 (N_7914,N_5468,N_7172);
nand U7915 (N_7915,N_7262,N_6994);
nor U7916 (N_7916,N_6637,N_6867);
nand U7917 (N_7917,N_7265,N_6427);
nor U7918 (N_7918,N_5147,N_6606);
xor U7919 (N_7919,N_6917,N_5060);
nor U7920 (N_7920,N_6119,N_7451);
or U7921 (N_7921,N_7137,N_7031);
nor U7922 (N_7922,N_6269,N_5019);
nand U7923 (N_7923,N_7166,N_5782);
nor U7924 (N_7924,N_5158,N_5680);
nor U7925 (N_7925,N_6668,N_7072);
nand U7926 (N_7926,N_6849,N_7158);
nor U7927 (N_7927,N_6909,N_7494);
nor U7928 (N_7928,N_5275,N_5216);
and U7929 (N_7929,N_7340,N_6075);
xor U7930 (N_7930,N_5503,N_6698);
xnor U7931 (N_7931,N_6050,N_5137);
nor U7932 (N_7932,N_5789,N_6122);
xor U7933 (N_7933,N_5482,N_5336);
and U7934 (N_7934,N_6406,N_7354);
and U7935 (N_7935,N_5842,N_6369);
nand U7936 (N_7936,N_6294,N_7319);
and U7937 (N_7937,N_5571,N_6859);
and U7938 (N_7938,N_5598,N_5895);
or U7939 (N_7939,N_7176,N_7107);
or U7940 (N_7940,N_7012,N_6768);
xnor U7941 (N_7941,N_5588,N_5770);
xnor U7942 (N_7942,N_5417,N_6170);
or U7943 (N_7943,N_6860,N_5155);
xnor U7944 (N_7944,N_6713,N_5113);
or U7945 (N_7945,N_5117,N_7205);
and U7946 (N_7946,N_5070,N_6111);
and U7947 (N_7947,N_7167,N_6364);
xor U7948 (N_7948,N_7427,N_7282);
or U7949 (N_7949,N_6520,N_5163);
nor U7950 (N_7950,N_6688,N_7188);
xnor U7951 (N_7951,N_6337,N_5211);
or U7952 (N_7952,N_6042,N_6117);
nand U7953 (N_7953,N_7352,N_7363);
nor U7954 (N_7954,N_6022,N_5946);
nor U7955 (N_7955,N_6268,N_5989);
xor U7956 (N_7956,N_6982,N_7375);
and U7957 (N_7957,N_7096,N_6542);
nand U7958 (N_7958,N_6761,N_5799);
nor U7959 (N_7959,N_6177,N_6946);
xnor U7960 (N_7960,N_6524,N_5677);
or U7961 (N_7961,N_5860,N_5967);
or U7962 (N_7962,N_7379,N_6016);
nor U7963 (N_7963,N_6158,N_5165);
nand U7964 (N_7964,N_6291,N_6939);
or U7965 (N_7965,N_7114,N_5824);
nand U7966 (N_7966,N_6565,N_7328);
nand U7967 (N_7967,N_6905,N_6610);
or U7968 (N_7968,N_6679,N_6614);
or U7969 (N_7969,N_5251,N_6202);
or U7970 (N_7970,N_5083,N_6755);
xor U7971 (N_7971,N_5197,N_6447);
xor U7972 (N_7972,N_7098,N_5930);
nand U7973 (N_7973,N_5914,N_5600);
and U7974 (N_7974,N_7089,N_7244);
xor U7975 (N_7975,N_5106,N_6295);
nand U7976 (N_7976,N_6303,N_6497);
xnor U7977 (N_7977,N_6243,N_6164);
or U7978 (N_7978,N_5264,N_6529);
xor U7979 (N_7979,N_6375,N_6141);
and U7980 (N_7980,N_5636,N_5351);
nor U7981 (N_7981,N_6339,N_6714);
and U7982 (N_7982,N_5921,N_6710);
and U7983 (N_7983,N_5800,N_7292);
or U7984 (N_7984,N_7490,N_6052);
and U7985 (N_7985,N_6880,N_5267);
nor U7986 (N_7986,N_5097,N_5268);
nand U7987 (N_7987,N_5213,N_5587);
xor U7988 (N_7988,N_6104,N_6548);
or U7989 (N_7989,N_5806,N_7063);
nand U7990 (N_7990,N_7061,N_5805);
xor U7991 (N_7991,N_6781,N_6522);
xor U7992 (N_7992,N_5325,N_6779);
and U7993 (N_7993,N_5237,N_6932);
xnor U7994 (N_7994,N_5915,N_6680);
nand U7995 (N_7995,N_7086,N_7331);
and U7996 (N_7996,N_5064,N_7487);
nor U7997 (N_7997,N_5152,N_7409);
and U7998 (N_7998,N_5001,N_5199);
and U7999 (N_7999,N_7395,N_5232);
nand U8000 (N_8000,N_6376,N_7278);
or U8001 (N_8001,N_6245,N_7094);
xor U8002 (N_8002,N_6490,N_5939);
nor U8003 (N_8003,N_5851,N_6056);
or U8004 (N_8004,N_5556,N_6273);
and U8005 (N_8005,N_6506,N_7279);
nor U8006 (N_8006,N_6450,N_5649);
xnor U8007 (N_8007,N_7413,N_6887);
or U8008 (N_8008,N_6572,N_7240);
or U8009 (N_8009,N_5887,N_6646);
and U8010 (N_8010,N_6635,N_5258);
or U8011 (N_8011,N_5350,N_6588);
nor U8012 (N_8012,N_5305,N_6470);
nand U8013 (N_8013,N_5710,N_6020);
or U8014 (N_8014,N_6931,N_6390);
nand U8015 (N_8015,N_6625,N_7134);
nor U8016 (N_8016,N_5443,N_7334);
nor U8017 (N_8017,N_5345,N_7394);
nor U8018 (N_8018,N_6727,N_6561);
and U8019 (N_8019,N_6891,N_6527);
and U8020 (N_8020,N_6385,N_7495);
nor U8021 (N_8021,N_6504,N_7422);
xnor U8022 (N_8022,N_5029,N_5129);
or U8023 (N_8023,N_5050,N_7085);
nand U8024 (N_8024,N_7017,N_6811);
xnor U8025 (N_8025,N_5762,N_7486);
nor U8026 (N_8026,N_6486,N_5419);
nand U8027 (N_8027,N_6477,N_7110);
and U8028 (N_8028,N_6575,N_5866);
or U8029 (N_8029,N_6791,N_5926);
nand U8030 (N_8030,N_5460,N_5925);
or U8031 (N_8031,N_7071,N_6792);
nand U8032 (N_8032,N_6569,N_6773);
xor U8033 (N_8033,N_6011,N_6672);
nand U8034 (N_8034,N_7150,N_5398);
nor U8035 (N_8035,N_5987,N_5792);
nor U8036 (N_8036,N_5391,N_6423);
or U8037 (N_8037,N_7213,N_5705);
xnor U8038 (N_8038,N_5749,N_7454);
nor U8039 (N_8039,N_5218,N_6555);
nor U8040 (N_8040,N_6328,N_6316);
nor U8041 (N_8041,N_7273,N_7093);
or U8042 (N_8042,N_6065,N_6827);
nor U8043 (N_8043,N_6469,N_5044);
nor U8044 (N_8044,N_5087,N_5430);
xor U8045 (N_8045,N_6510,N_7372);
nor U8046 (N_8046,N_5057,N_5285);
and U8047 (N_8047,N_5942,N_6503);
nand U8048 (N_8048,N_6092,N_6381);
and U8049 (N_8049,N_7311,N_5821);
xor U8050 (N_8050,N_7006,N_5912);
nand U8051 (N_8051,N_6321,N_6925);
nand U8052 (N_8052,N_5751,N_7060);
xor U8053 (N_8053,N_5292,N_5380);
nor U8054 (N_8054,N_5624,N_6066);
xnor U8055 (N_8055,N_6788,N_5479);
or U8056 (N_8056,N_5934,N_6071);
xnor U8057 (N_8057,N_5672,N_6564);
nand U8058 (N_8058,N_5500,N_7274);
and U8059 (N_8059,N_7275,N_5881);
or U8060 (N_8060,N_6310,N_6007);
nor U8061 (N_8061,N_6207,N_5375);
or U8062 (N_8062,N_5968,N_5066);
nor U8063 (N_8063,N_6312,N_6633);
and U8064 (N_8064,N_7325,N_6431);
or U8065 (N_8065,N_5254,N_6010);
and U8066 (N_8066,N_6978,N_7052);
xor U8067 (N_8067,N_6184,N_5047);
or U8068 (N_8068,N_6686,N_7426);
nor U8069 (N_8069,N_6183,N_6145);
nor U8070 (N_8070,N_6093,N_5453);
and U8071 (N_8071,N_7095,N_6578);
and U8072 (N_8072,N_6248,N_6412);
or U8073 (N_8073,N_6554,N_5470);
nand U8074 (N_8074,N_7432,N_6426);
xnor U8075 (N_8075,N_5327,N_6619);
or U8076 (N_8076,N_5960,N_5615);
or U8077 (N_8077,N_6894,N_5421);
nand U8078 (N_8078,N_6511,N_7469);
nor U8079 (N_8079,N_6919,N_5700);
nor U8080 (N_8080,N_6414,N_7231);
nand U8081 (N_8081,N_5178,N_5017);
or U8082 (N_8082,N_5269,N_6900);
or U8083 (N_8083,N_5691,N_7132);
xnor U8084 (N_8084,N_5767,N_5201);
or U8085 (N_8085,N_7269,N_6004);
nor U8086 (N_8086,N_6532,N_6918);
or U8087 (N_8087,N_5013,N_6459);
nand U8088 (N_8088,N_7456,N_6817);
and U8089 (N_8089,N_5436,N_5499);
or U8090 (N_8090,N_7183,N_6465);
or U8091 (N_8091,N_5407,N_7357);
or U8092 (N_8092,N_5695,N_6808);
xnor U8093 (N_8093,N_7410,N_6921);
nand U8094 (N_8094,N_6669,N_6806);
xor U8095 (N_8095,N_5459,N_5488);
nand U8096 (N_8096,N_5875,N_7284);
nor U8097 (N_8097,N_7036,N_6613);
xnor U8098 (N_8098,N_7256,N_6903);
nor U8099 (N_8099,N_6134,N_7358);
or U8100 (N_8100,N_6132,N_7165);
nand U8101 (N_8101,N_6720,N_5053);
nor U8102 (N_8102,N_5918,N_6662);
and U8103 (N_8103,N_5604,N_5829);
or U8104 (N_8104,N_5547,N_5221);
nor U8105 (N_8105,N_7201,N_5347);
xor U8106 (N_8106,N_5874,N_6451);
nor U8107 (N_8107,N_7356,N_7333);
nand U8108 (N_8108,N_5072,N_6432);
xnor U8109 (N_8109,N_5183,N_5728);
xnor U8110 (N_8110,N_5256,N_6945);
xor U8111 (N_8111,N_7435,N_6923);
and U8112 (N_8112,N_5813,N_7041);
nor U8113 (N_8113,N_6151,N_6762);
xor U8114 (N_8114,N_6983,N_6094);
and U8115 (N_8115,N_7414,N_5411);
xnor U8116 (N_8116,N_6641,N_5022);
nand U8117 (N_8117,N_6841,N_5400);
or U8118 (N_8118,N_7040,N_5492);
and U8119 (N_8119,N_7475,N_5623);
nand U8120 (N_8120,N_5739,N_6118);
nand U8121 (N_8121,N_7026,N_6246);
nand U8122 (N_8122,N_5310,N_7445);
and U8123 (N_8123,N_6396,N_5239);
xor U8124 (N_8124,N_6262,N_7368);
xnor U8125 (N_8125,N_6947,N_6989);
or U8126 (N_8126,N_5899,N_6553);
and U8127 (N_8127,N_7100,N_5740);
nand U8128 (N_8128,N_6332,N_5360);
nor U8129 (N_8129,N_6833,N_7113);
or U8130 (N_8130,N_7326,N_6812);
nor U8131 (N_8131,N_6711,N_6580);
nor U8132 (N_8132,N_5796,N_6896);
nor U8133 (N_8133,N_7323,N_7097);
xnor U8134 (N_8134,N_5509,N_6402);
and U8135 (N_8135,N_7008,N_6257);
nor U8136 (N_8136,N_6289,N_5667);
nand U8137 (N_8137,N_5309,N_6323);
nor U8138 (N_8138,N_7076,N_6058);
xor U8139 (N_8139,N_7455,N_6759);
nor U8140 (N_8140,N_7304,N_5888);
and U8141 (N_8141,N_6153,N_6109);
xor U8142 (N_8142,N_7212,N_6281);
xor U8143 (N_8143,N_7203,N_7485);
nand U8144 (N_8144,N_6985,N_6479);
nand U8145 (N_8145,N_5474,N_5823);
xor U8146 (N_8146,N_6913,N_7327);
xor U8147 (N_8147,N_7020,N_6028);
nand U8148 (N_8148,N_6883,N_5259);
nor U8149 (N_8149,N_5828,N_5427);
nand U8150 (N_8150,N_5204,N_7286);
nor U8151 (N_8151,N_6928,N_5033);
and U8152 (N_8152,N_6225,N_5338);
or U8153 (N_8153,N_7364,N_7035);
nand U8154 (N_8154,N_5849,N_5455);
or U8155 (N_8155,N_6826,N_5681);
nand U8156 (N_8156,N_5685,N_5601);
and U8157 (N_8157,N_5978,N_6345);
xor U8158 (N_8158,N_5377,N_7470);
and U8159 (N_8159,N_5349,N_7281);
nor U8160 (N_8160,N_6379,N_6421);
and U8161 (N_8161,N_6601,N_5658);
xnor U8162 (N_8162,N_6566,N_6018);
or U8163 (N_8163,N_5186,N_6439);
or U8164 (N_8164,N_5859,N_5657);
and U8165 (N_8165,N_5861,N_6064);
and U8166 (N_8166,N_5643,N_6960);
nor U8167 (N_8167,N_7305,N_7074);
nand U8168 (N_8168,N_5633,N_6253);
nor U8169 (N_8169,N_6835,N_5847);
nor U8170 (N_8170,N_5994,N_6080);
nand U8171 (N_8171,N_6103,N_7144);
xnor U8172 (N_8172,N_6589,N_6915);
or U8173 (N_8173,N_6839,N_7217);
xnor U8174 (N_8174,N_5156,N_6265);
and U8175 (N_8175,N_6003,N_6139);
or U8176 (N_8176,N_5759,N_7064);
and U8177 (N_8177,N_6137,N_7195);
xor U8178 (N_8178,N_7461,N_6214);
or U8179 (N_8179,N_5908,N_6513);
nor U8180 (N_8180,N_7349,N_7054);
nand U8181 (N_8181,N_5917,N_6725);
nor U8182 (N_8182,N_6803,N_5376);
nor U8183 (N_8183,N_5115,N_5858);
xor U8184 (N_8184,N_5629,N_6990);
and U8185 (N_8185,N_5904,N_7433);
xor U8186 (N_8186,N_6831,N_6996);
nor U8187 (N_8187,N_6954,N_6699);
or U8188 (N_8188,N_5738,N_5101);
nand U8189 (N_8189,N_5748,N_5322);
nor U8190 (N_8190,N_7453,N_5790);
and U8191 (N_8191,N_5659,N_5025);
and U8192 (N_8192,N_6777,N_7070);
or U8193 (N_8193,N_5193,N_5300);
nor U8194 (N_8194,N_7294,N_6677);
nor U8195 (N_8195,N_6025,N_6389);
and U8196 (N_8196,N_6549,N_5564);
and U8197 (N_8197,N_6178,N_6186);
and U8198 (N_8198,N_5527,N_5192);
nor U8199 (N_8199,N_5059,N_6628);
or U8200 (N_8200,N_6460,N_6975);
xnor U8201 (N_8201,N_5086,N_5215);
or U8202 (N_8202,N_5379,N_5603);
and U8203 (N_8203,N_5128,N_6654);
xor U8204 (N_8204,N_6300,N_6351);
xnor U8205 (N_8205,N_5750,N_5983);
or U8206 (N_8206,N_5280,N_7161);
nor U8207 (N_8207,N_6029,N_6114);
nand U8208 (N_8208,N_5938,N_5046);
or U8209 (N_8209,N_6944,N_7218);
or U8210 (N_8210,N_6970,N_6749);
and U8211 (N_8211,N_5575,N_6797);
nand U8212 (N_8212,N_6744,N_6590);
or U8213 (N_8213,N_7224,N_6892);
xnor U8214 (N_8214,N_6574,N_7317);
nor U8215 (N_8215,N_7446,N_5058);
nor U8216 (N_8216,N_6348,N_5697);
or U8217 (N_8217,N_6516,N_7345);
or U8218 (N_8218,N_6692,N_6446);
and U8219 (N_8219,N_5817,N_5016);
and U8220 (N_8220,N_6073,N_6546);
or U8221 (N_8221,N_5873,N_5711);
nand U8222 (N_8222,N_7009,N_7002);
xnor U8223 (N_8223,N_6236,N_6422);
and U8224 (N_8224,N_7050,N_7384);
and U8225 (N_8225,N_6828,N_7170);
or U8226 (N_8226,N_5257,N_5822);
nand U8227 (N_8227,N_6870,N_7287);
xor U8228 (N_8228,N_6392,N_5606);
xor U8229 (N_8229,N_6239,N_5736);
xnor U8230 (N_8230,N_6571,N_6305);
nand U8231 (N_8231,N_7343,N_6731);
nand U8232 (N_8232,N_5996,N_5337);
xor U8233 (N_8233,N_5130,N_6612);
xnor U8234 (N_8234,N_7117,N_5154);
and U8235 (N_8235,N_6330,N_5076);
and U8236 (N_8236,N_5530,N_5980);
xnor U8237 (N_8237,N_5771,N_6032);
nor U8238 (N_8238,N_6842,N_6528);
or U8239 (N_8239,N_5255,N_6784);
xnor U8240 (N_8240,N_6728,N_6256);
or U8241 (N_8241,N_6034,N_7047);
xnor U8242 (N_8242,N_5801,N_5704);
nand U8243 (N_8243,N_5052,N_6314);
xnor U8244 (N_8244,N_7252,N_7004);
nor U8245 (N_8245,N_7484,N_6060);
or U8246 (N_8246,N_5553,N_5516);
nor U8247 (N_8247,N_6420,N_5439);
and U8248 (N_8248,N_6167,N_7029);
nand U8249 (N_8249,N_7152,N_7316);
xor U8250 (N_8250,N_7214,N_6893);
and U8251 (N_8251,N_6143,N_6579);
and U8252 (N_8252,N_5423,N_6163);
and U8253 (N_8253,N_6934,N_5365);
nand U8254 (N_8254,N_6622,N_7429);
nand U8255 (N_8255,N_5472,N_7285);
and U8256 (N_8256,N_7042,N_5133);
and U8257 (N_8257,N_5905,N_6594);
nand U8258 (N_8258,N_7225,N_7472);
nor U8259 (N_8259,N_7300,N_6276);
nand U8260 (N_8260,N_5557,N_5140);
or U8261 (N_8261,N_5226,N_6361);
nand U8262 (N_8262,N_5826,N_7496);
xnor U8263 (N_8263,N_7007,N_6716);
nor U8264 (N_8264,N_7186,N_5177);
and U8265 (N_8265,N_6875,N_7443);
or U8266 (N_8266,N_6620,N_5314);
nand U8267 (N_8267,N_5448,N_7037);
nand U8268 (N_8268,N_5428,N_6046);
nand U8269 (N_8269,N_5333,N_7423);
nand U8270 (N_8270,N_6150,N_6823);
nand U8271 (N_8271,N_5613,N_5307);
xnor U8272 (N_8272,N_6380,N_5082);
and U8273 (N_8273,N_6584,N_6798);
nand U8274 (N_8274,N_7361,N_6534);
nor U8275 (N_8275,N_6804,N_6116);
nand U8276 (N_8276,N_6886,N_6738);
nand U8277 (N_8277,N_7367,N_7390);
xor U8278 (N_8278,N_7023,N_7314);
xnor U8279 (N_8279,N_5815,N_6952);
nand U8280 (N_8280,N_6067,N_7291);
xor U8281 (N_8281,N_6326,N_5020);
or U8282 (N_8282,N_6922,N_5528);
xnor U8283 (N_8283,N_5551,N_5437);
nor U8284 (N_8284,N_5777,N_6660);
xor U8285 (N_8285,N_7032,N_5496);
nand U8286 (N_8286,N_5132,N_5787);
xnor U8287 (N_8287,N_5674,N_5355);
xnor U8288 (N_8288,N_5877,N_6767);
xnor U8289 (N_8289,N_6407,N_7088);
or U8290 (N_8290,N_6617,N_5742);
nor U8291 (N_8291,N_5673,N_5632);
xnor U8292 (N_8292,N_5318,N_5340);
xnor U8293 (N_8293,N_5586,N_5424);
nor U8294 (N_8294,N_7190,N_6920);
nor U8295 (N_8295,N_5088,N_5886);
xor U8296 (N_8296,N_6769,N_5014);
and U8297 (N_8297,N_6972,N_5610);
nand U8298 (N_8298,N_6665,N_6017);
nor U8299 (N_8299,N_6371,N_5538);
and U8300 (N_8300,N_5884,N_7149);
nand U8301 (N_8301,N_6394,N_6404);
and U8302 (N_8302,N_6199,N_5737);
or U8303 (N_8303,N_5628,N_6813);
or U8304 (N_8304,N_5273,N_5572);
xor U8305 (N_8305,N_5953,N_5816);
or U8306 (N_8306,N_5730,N_5301);
or U8307 (N_8307,N_6847,N_6822);
nor U8308 (N_8308,N_6502,N_5692);
nor U8309 (N_8309,N_6539,N_5248);
or U8310 (N_8310,N_6604,N_5012);
nand U8311 (N_8311,N_5230,N_5579);
nor U8312 (N_8312,N_7257,N_5889);
xnor U8313 (N_8313,N_5162,N_5198);
nand U8314 (N_8314,N_7108,N_5095);
or U8315 (N_8315,N_5069,N_7310);
and U8316 (N_8316,N_5833,N_5524);
xnor U8317 (N_8317,N_6512,N_5493);
nor U8318 (N_8318,N_6327,N_7232);
nand U8319 (N_8319,N_6965,N_5732);
xnor U8320 (N_8320,N_6395,N_6284);
and U8321 (N_8321,N_7118,N_5299);
nor U8322 (N_8322,N_5032,N_7043);
nand U8323 (N_8323,N_5279,N_5637);
nor U8324 (N_8324,N_6278,N_6463);
nand U8325 (N_8325,N_5005,N_6609);
xnor U8326 (N_8326,N_6342,N_7386);
or U8327 (N_8327,N_5332,N_5901);
nand U8328 (N_8328,N_6179,N_7474);
and U8329 (N_8329,N_5127,N_6499);
or U8330 (N_8330,N_5194,N_6760);
and U8331 (N_8331,N_5390,N_5593);
and U8332 (N_8332,N_5712,N_7124);
nand U8333 (N_8333,N_5641,N_5042);
and U8334 (N_8334,N_6914,N_6443);
and U8335 (N_8335,N_6586,N_5063);
or U8336 (N_8336,N_6086,N_7174);
nor U8337 (N_8337,N_5857,N_6074);
nor U8338 (N_8338,N_6632,N_6220);
nor U8339 (N_8339,N_5036,N_7162);
and U8340 (N_8340,N_6658,N_5971);
and U8341 (N_8341,N_6386,N_5947);
and U8342 (N_8342,N_6461,N_5189);
xnor U8343 (N_8343,N_6472,N_7348);
xor U8344 (N_8344,N_5683,N_6766);
and U8345 (N_8345,N_5385,N_5085);
or U8346 (N_8346,N_7339,N_7351);
xor U8347 (N_8347,N_6059,N_7018);
nor U8348 (N_8348,N_6581,N_5124);
nand U8349 (N_8349,N_5715,N_6517);
xnor U8350 (N_8350,N_5465,N_7336);
nor U8351 (N_8351,N_5200,N_7125);
nand U8352 (N_8352,N_6221,N_5597);
or U8353 (N_8353,N_6702,N_6515);
or U8354 (N_8354,N_5892,N_5621);
nor U8355 (N_8355,N_7196,N_5445);
or U8356 (N_8356,N_7163,N_5949);
and U8357 (N_8357,N_6888,N_5879);
or U8358 (N_8358,N_6098,N_6343);
xor U8359 (N_8359,N_5481,N_5975);
nand U8360 (N_8360,N_5988,N_6648);
nand U8361 (N_8361,N_6538,N_5612);
and U8362 (N_8362,N_5970,N_6036);
nand U8363 (N_8363,N_6089,N_6795);
nor U8364 (N_8364,N_5395,N_6899);
xnor U8365 (N_8365,N_6559,N_5442);
nand U8366 (N_8366,N_6140,N_6027);
xor U8367 (N_8367,N_5717,N_5897);
nor U8368 (N_8368,N_6958,N_7464);
nand U8369 (N_8369,N_5383,N_5791);
xor U8370 (N_8370,N_5755,N_6258);
xnor U8371 (N_8371,N_5202,N_5111);
and U8372 (N_8372,N_5123,N_5160);
or U8373 (N_8373,N_6233,N_7011);
nand U8374 (N_8374,N_6765,N_7428);
and U8375 (N_8375,N_6674,N_6570);
or U8376 (N_8376,N_6723,N_5368);
nor U8377 (N_8377,N_5655,N_7171);
and U8378 (N_8378,N_7080,N_7437);
xor U8379 (N_8379,N_6482,N_5190);
nor U8380 (N_8380,N_5176,N_6603);
or U8381 (N_8381,N_5911,N_6508);
xnor U8382 (N_8382,N_6531,N_6317);
nand U8383 (N_8383,N_6799,N_6526);
or U8384 (N_8384,N_6898,N_5354);
nor U8385 (N_8385,N_6416,N_7308);
nand U8386 (N_8386,N_5995,N_6242);
and U8387 (N_8387,N_5303,N_5565);
xor U8388 (N_8388,N_6618,N_6128);
nor U8389 (N_8389,N_5396,N_5609);
and U8390 (N_8390,N_6264,N_6748);
xnor U8391 (N_8391,N_5793,N_5541);
and U8392 (N_8392,N_5803,N_5161);
xnor U8393 (N_8393,N_6943,N_5209);
or U8394 (N_8394,N_5108,N_6428);
xor U8395 (N_8395,N_7169,N_7102);
or U8396 (N_8396,N_5945,N_7268);
and U8397 (N_8397,N_5662,N_6309);
and U8398 (N_8398,N_6780,N_6855);
xnor U8399 (N_8399,N_6879,N_5568);
nand U8400 (N_8400,N_6745,N_5173);
xnor U8401 (N_8401,N_5374,N_7408);
nand U8402 (N_8402,N_6062,N_5843);
nor U8403 (N_8403,N_5403,N_5776);
nor U8404 (N_8404,N_6703,N_5569);
nor U8405 (N_8405,N_7219,N_5188);
nor U8406 (N_8406,N_5747,N_5282);
nand U8407 (N_8407,N_5701,N_6981);
or U8408 (N_8408,N_6436,N_6629);
nand U8409 (N_8409,N_5222,N_5238);
xor U8410 (N_8410,N_6962,N_6616);
xnor U8411 (N_8411,N_5546,N_7288);
and U8412 (N_8412,N_5555,N_5471);
nand U8413 (N_8413,N_6602,N_7001);
or U8414 (N_8414,N_5234,N_6587);
and U8415 (N_8415,N_5265,N_7059);
nor U8416 (N_8416,N_5039,N_7362);
and U8417 (N_8417,N_5663,N_7199);
and U8418 (N_8418,N_6474,N_6959);
nand U8419 (N_8419,N_5272,N_5772);
or U8420 (N_8420,N_6370,N_6541);
nand U8421 (N_8421,N_6678,N_6607);
and U8422 (N_8422,N_5961,N_5814);
nand U8423 (N_8423,N_5049,N_6488);
or U8424 (N_8424,N_5451,N_7103);
nand U8425 (N_8425,N_5894,N_7315);
and U8426 (N_8426,N_6627,N_6556);
or U8427 (N_8427,N_7234,N_6251);
nor U8428 (N_8428,N_6785,N_7184);
or U8429 (N_8429,N_6418,N_6204);
or U8430 (N_8430,N_6988,N_7293);
nand U8431 (N_8431,N_7471,N_5856);
or U8432 (N_8432,N_5784,N_6717);
and U8433 (N_8433,N_7374,N_6691);
or U8434 (N_8434,N_6681,N_6285);
nand U8435 (N_8435,N_5519,N_6095);
nand U8436 (N_8436,N_5678,N_5134);
or U8437 (N_8437,N_7216,N_6709);
nand U8438 (N_8438,N_5415,N_6165);
and U8439 (N_8439,N_5098,N_6854);
and U8440 (N_8440,N_6024,N_5559);
nand U8441 (N_8441,N_5119,N_7207);
nand U8442 (N_8442,N_6142,N_5051);
and U8443 (N_8443,N_6378,N_6783);
nor U8444 (N_8444,N_6147,N_6190);
nor U8445 (N_8445,N_5714,N_6324);
xor U8446 (N_8446,N_5399,N_7492);
xor U8447 (N_8447,N_6457,N_6984);
and U8448 (N_8448,N_6659,N_6279);
xnor U8449 (N_8449,N_5028,N_5694);
or U8450 (N_8450,N_7154,N_6274);
and U8451 (N_8451,N_6694,N_5018);
nor U8452 (N_8452,N_5964,N_7380);
nor U8453 (N_8453,N_7463,N_5532);
nor U8454 (N_8454,N_6430,N_6756);
and U8455 (N_8455,N_7143,N_7129);
or U8456 (N_8456,N_7192,N_5958);
nand U8457 (N_8457,N_6383,N_5935);
or U8458 (N_8458,N_6372,N_7296);
and U8459 (N_8459,N_6690,N_6043);
xnor U8460 (N_8460,N_6832,N_6836);
and U8461 (N_8461,N_5607,N_7473);
nand U8462 (N_8462,N_6929,N_7299);
xor U8463 (N_8463,N_5581,N_6201);
nor U8464 (N_8464,N_7246,N_7365);
xor U8465 (N_8465,N_5936,N_6991);
or U8466 (N_8466,N_5242,N_5466);
or U8467 (N_8467,N_6901,N_6206);
or U8468 (N_8468,N_5288,N_5537);
and U8469 (N_8469,N_5871,N_7321);
xor U8470 (N_8470,N_7200,N_6624);
nor U8471 (N_8471,N_6366,N_5850);
and U8472 (N_8472,N_7359,N_5446);
nor U8473 (N_8473,N_6857,N_5661);
and U8474 (N_8474,N_6105,N_6846);
and U8475 (N_8475,N_6162,N_7164);
and U8476 (N_8476,N_7397,N_6260);
nor U8477 (N_8477,N_5645,N_5722);
xor U8478 (N_8478,N_6448,N_5903);
nor U8479 (N_8479,N_5999,N_6456);
and U8480 (N_8480,N_7465,N_6212);
and U8481 (N_8481,N_7450,N_5371);
nor U8482 (N_8482,N_5179,N_5120);
nor U8483 (N_8483,N_5622,N_6676);
or U8484 (N_8484,N_7127,N_6229);
or U8485 (N_8485,N_6884,N_5809);
xnor U8486 (N_8486,N_6873,N_5458);
xnor U8487 (N_8487,N_6776,N_5545);
and U8488 (N_8488,N_6159,N_5081);
and U8489 (N_8489,N_6653,N_6129);
nand U8490 (N_8490,N_7022,N_6583);
nand U8491 (N_8491,N_7449,N_6639);
xor U8492 (N_8492,N_6121,N_6980);
and U8493 (N_8493,N_7419,N_5552);
xor U8494 (N_8494,N_7039,N_7079);
nand U8495 (N_8495,N_6315,N_5798);
xnor U8496 (N_8496,N_5727,N_5461);
xor U8497 (N_8497,N_6413,N_6487);
nand U8498 (N_8498,N_5079,N_6596);
nand U8499 (N_8499,N_6155,N_6249);
xnor U8500 (N_8500,N_5670,N_6636);
and U8501 (N_8501,N_7155,N_7235);
nand U8502 (N_8502,N_5425,N_6148);
nand U8503 (N_8503,N_5312,N_6078);
xor U8504 (N_8504,N_6494,N_6735);
nor U8505 (N_8505,N_6483,N_6906);
nor U8506 (N_8506,N_5725,N_6706);
nand U8507 (N_8507,N_6949,N_5122);
and U8508 (N_8508,N_7405,N_7254);
or U8509 (N_8509,N_6344,N_6054);
xnor U8510 (N_8510,N_6341,N_5627);
and U8511 (N_8511,N_6340,N_7058);
and U8512 (N_8512,N_5863,N_6437);
nand U8513 (N_8513,N_5626,N_5306);
and U8514 (N_8514,N_5068,N_6399);
and U8515 (N_8515,N_5576,N_6824);
and U8516 (N_8516,N_6039,N_5406);
nand U8517 (N_8517,N_5438,N_6593);
xor U8518 (N_8518,N_6444,N_6995);
or U8519 (N_8519,N_6266,N_7400);
nand U8520 (N_8520,N_7077,N_7197);
xor U8521 (N_8521,N_7179,N_5617);
nor U8522 (N_8522,N_6192,N_5041);
nor U8523 (N_8523,N_5716,N_7260);
and U8524 (N_8524,N_6734,N_5092);
nor U8525 (N_8525,N_6519,N_6049);
nor U8526 (N_8526,N_7227,N_6107);
and U8527 (N_8527,N_5511,N_5689);
nand U8528 (N_8528,N_5745,N_5825);
nor U8529 (N_8529,N_6885,N_5656);
nand U8530 (N_8530,N_5638,N_5035);
nor U8531 (N_8531,N_6663,N_5614);
and U8532 (N_8532,N_7434,N_5164);
xor U8533 (N_8533,N_5277,N_6438);
nand U8534 (N_8534,N_7425,N_6638);
or U8535 (N_8535,N_7476,N_5959);
nor U8536 (N_8536,N_7249,N_5373);
nand U8537 (N_8537,N_5091,N_6897);
or U8538 (N_8538,N_7276,N_5896);
nor U8539 (N_8539,N_6360,N_6651);
nand U8540 (N_8540,N_6044,N_5250);
or U8541 (N_8541,N_6435,N_5840);
or U8542 (N_8542,N_6751,N_6215);
nand U8543 (N_8543,N_6848,N_5270);
nor U8544 (N_8544,N_7198,N_5384);
nand U8545 (N_8545,N_7439,N_6999);
nor U8546 (N_8546,N_5990,N_6169);
nand U8547 (N_8547,N_5549,N_5323);
nor U8548 (N_8548,N_5319,N_6288);
and U8549 (N_8549,N_5940,N_5560);
or U8550 (N_8550,N_6743,N_7447);
or U8551 (N_8551,N_5544,N_6403);
nand U8552 (N_8552,N_7440,N_6650);
or U8553 (N_8553,N_5654,N_5168);
and U8554 (N_8554,N_5056,N_5928);
and U8555 (N_8555,N_6480,N_7393);
nor U8556 (N_8556,N_5867,N_7415);
or U8557 (N_8557,N_6087,N_6405);
and U8558 (N_8558,N_6563,N_7322);
xnor U8559 (N_8559,N_5652,N_6096);
and U8560 (N_8560,N_5114,N_7131);
or U8561 (N_8561,N_5923,N_5225);
nor U8562 (N_8562,N_5431,N_6547);
or U8563 (N_8563,N_6133,N_6973);
xor U8564 (N_8564,N_6521,N_6449);
nor U8565 (N_8565,N_5363,N_7159);
nand U8566 (N_8566,N_6441,N_7078);
nand U8567 (N_8567,N_6464,N_5112);
and U8568 (N_8568,N_5635,N_6123);
and U8569 (N_8569,N_6858,N_7259);
xor U8570 (N_8570,N_6277,N_6146);
and U8571 (N_8571,N_6582,N_5902);
and U8572 (N_8572,N_5666,N_6077);
nand U8573 (N_8573,N_5214,N_5021);
nor U8574 (N_8574,N_5326,N_6869);
nor U8575 (N_8575,N_6774,N_5346);
nor U8576 (N_8576,N_7389,N_5015);
or U8577 (N_8577,N_7271,N_7306);
nand U8578 (N_8578,N_5885,N_5497);
nand U8579 (N_8579,N_5002,N_5804);
xnor U8580 (N_8580,N_7053,N_5260);
xor U8581 (N_8581,N_7404,N_5146);
nand U8582 (N_8582,N_7416,N_7104);
xnor U8583 (N_8583,N_6240,N_5620);
nand U8584 (N_8584,N_6250,N_7460);
nor U8585 (N_8585,N_6346,N_7270);
nand U8586 (N_8586,N_5820,N_5992);
xnor U8587 (N_8587,N_6997,N_5690);
or U8588 (N_8588,N_7090,N_5846);
nor U8589 (N_8589,N_5536,N_5404);
nor U8590 (N_8590,N_6567,N_5699);
nand U8591 (N_8591,N_6261,N_6640);
and U8592 (N_8592,N_6568,N_6966);
and U8593 (N_8593,N_7272,N_7307);
xor U8594 (N_8594,N_6874,N_6325);
or U8595 (N_8595,N_6275,N_7338);
nand U8596 (N_8596,N_6800,N_5526);
nor U8597 (N_8597,N_5948,N_6445);
or U8598 (N_8598,N_5554,N_5167);
xnor U8599 (N_8599,N_6076,N_7048);
xor U8600 (N_8600,N_6149,N_6493);
nand U8601 (N_8601,N_5320,N_5795);
xor U8602 (N_8602,N_5752,N_5898);
or U8603 (N_8603,N_7145,N_5220);
and U8604 (N_8604,N_6362,N_7230);
and U8605 (N_8605,N_6834,N_5030);
nor U8606 (N_8606,N_6218,N_5207);
nand U8607 (N_8607,N_5734,N_7290);
xor U8608 (N_8608,N_6290,N_6758);
nand U8609 (N_8609,N_6757,N_6523);
or U8610 (N_8610,N_7038,N_5594);
and U8611 (N_8611,N_5071,N_5642);
xnor U8612 (N_8612,N_5788,N_6124);
nor U8613 (N_8613,N_5394,N_5432);
and U8614 (N_8614,N_7209,N_7467);
nor U8615 (N_8615,N_6689,N_6185);
xor U8616 (N_8616,N_5682,N_6387);
nand U8617 (N_8617,N_6191,N_6505);
xor U8618 (N_8618,N_7014,N_5024);
nor U8619 (N_8619,N_6335,N_7498);
or U8620 (N_8620,N_6292,N_6198);
nand U8621 (N_8621,N_7479,N_5646);
and U8622 (N_8622,N_5513,N_7499);
and U8623 (N_8623,N_5794,N_7267);
nand U8624 (N_8624,N_5965,N_5153);
nor U8625 (N_8625,N_6865,N_7387);
xnor U8626 (N_8626,N_5464,N_6540);
nand U8627 (N_8627,N_6937,N_5352);
nor U8628 (N_8628,N_5540,N_6197);
nor U8629 (N_8629,N_5463,N_5426);
nand U8630 (N_8630,N_6543,N_5506);
xor U8631 (N_8631,N_6856,N_6187);
nand U8632 (N_8632,N_5342,N_5382);
nand U8633 (N_8633,N_5243,N_5412);
xor U8634 (N_8634,N_5731,N_5764);
nor U8635 (N_8635,N_5743,N_6868);
or U8636 (N_8636,N_5339,N_5392);
nor U8637 (N_8637,N_7211,N_6805);
and U8638 (N_8638,N_6466,N_6558);
nand U8639 (N_8639,N_7126,N_5480);
or U8640 (N_8640,N_5502,N_5450);
nor U8641 (N_8641,N_5839,N_6630);
nor U8642 (N_8642,N_6001,N_5891);
and U8643 (N_8643,N_6941,N_5779);
or U8644 (N_8644,N_6598,N_5618);
nand U8645 (N_8645,N_5836,N_7003);
nand U8646 (N_8646,N_5054,N_5229);
nand U8647 (N_8647,N_7193,N_6675);
nand U8648 (N_8648,N_5644,N_6084);
or U8649 (N_8649,N_5093,N_6391);
nand U8650 (N_8650,N_5534,N_6509);
and U8651 (N_8651,N_5976,N_5296);
xor U8652 (N_8652,N_5475,N_5542);
nand U8653 (N_8653,N_6297,N_7399);
nor U8654 (N_8654,N_5434,N_5485);
nor U8655 (N_8655,N_6772,N_5950);
xor U8656 (N_8656,N_6536,N_6397);
nor U8657 (N_8657,N_7136,N_7141);
and U8658 (N_8658,N_5454,N_5726);
and U8659 (N_8659,N_7431,N_5369);
or U8660 (N_8660,N_7010,N_7263);
or U8661 (N_8661,N_5880,N_6419);
or U8662 (N_8662,N_6700,N_6228);
or U8663 (N_8663,N_5535,N_7332);
xor U8664 (N_8664,N_5561,N_5131);
and U8665 (N_8665,N_7236,N_5582);
and U8666 (N_8666,N_6014,N_5596);
xor U8667 (N_8667,N_6304,N_6557);
nor U8668 (N_8668,N_6272,N_5266);
nor U8669 (N_8669,N_5366,N_6771);
or U8670 (N_8670,N_7497,N_6741);
nand U8671 (N_8671,N_6712,N_7139);
or U8672 (N_8672,N_6259,N_5182);
nand U8673 (N_8673,N_7068,N_6454);
or U8674 (N_8674,N_5702,N_6063);
nand U8675 (N_8675,N_6600,N_5241);
or U8676 (N_8676,N_5388,N_5531);
nand U8677 (N_8677,N_5009,N_7436);
nand U8678 (N_8678,N_7112,N_5159);
nor U8679 (N_8679,N_5143,N_6895);
or U8680 (N_8680,N_6754,N_5906);
or U8681 (N_8681,N_6041,N_6216);
or U8682 (N_8682,N_5416,N_6252);
and U8683 (N_8683,N_7065,N_5679);
nand U8684 (N_8684,N_5142,N_5515);
xor U8685 (N_8685,N_6863,N_6478);
and U8686 (N_8686,N_6701,N_5916);
and U8687 (N_8687,N_5746,N_5508);
xnor U8688 (N_8688,N_6070,N_7406);
xor U8689 (N_8689,N_6035,N_7369);
nor U8690 (N_8690,N_7238,N_5539);
and U8691 (N_8691,N_5290,N_5080);
or U8692 (N_8692,N_7407,N_7138);
nor U8693 (N_8693,N_6643,N_5941);
nor U8694 (N_8694,N_5110,N_6322);
or U8695 (N_8695,N_5830,N_6696);
and U8696 (N_8696,N_6652,N_6862);
xor U8697 (N_8697,N_7295,N_6850);
nand U8698 (N_8698,N_6707,N_5023);
nor U8699 (N_8699,N_5827,N_6267);
nor U8700 (N_8700,N_6005,N_6359);
and U8701 (N_8701,N_5868,N_7376);
nor U8702 (N_8702,N_7403,N_6083);
xor U8703 (N_8703,N_6270,N_6255);
nand U8704 (N_8704,N_6090,N_7194);
and U8705 (N_8705,N_5191,N_5007);
and U8706 (N_8706,N_6957,N_6082);
nand U8707 (N_8707,N_6697,N_5457);
nor U8708 (N_8708,N_6977,N_6298);
or U8709 (N_8709,N_7191,N_5910);
or U8710 (N_8710,N_7021,N_5217);
xor U8711 (N_8711,N_5378,N_5919);
nand U8712 (N_8712,N_6816,N_6347);
nand U8713 (N_8713,N_5075,N_7101);
nor U8714 (N_8714,N_6693,N_5449);
xnor U8715 (N_8715,N_5483,N_7140);
and U8716 (N_8716,N_5832,N_6473);
nor U8717 (N_8717,N_5227,N_5721);
xnor U8718 (N_8718,N_6851,N_5125);
nand U8719 (N_8719,N_6573,N_6026);
nand U8720 (N_8720,N_6775,N_5196);
nand U8721 (N_8721,N_5584,N_6802);
nor U8722 (N_8722,N_5262,N_6864);
nand U8723 (N_8723,N_6468,N_5984);
and U8724 (N_8724,N_5786,N_6411);
or U8725 (N_8725,N_6174,N_5713);
xnor U8726 (N_8726,N_5514,N_6173);
nor U8727 (N_8727,N_5393,N_5937);
or U8728 (N_8728,N_6211,N_6591);
nor U8729 (N_8729,N_6100,N_5616);
xor U8730 (N_8730,N_5605,N_5741);
or U8731 (N_8731,N_7019,N_7075);
nand U8732 (N_8732,N_5760,N_7034);
or U8733 (N_8733,N_5507,N_5529);
or U8734 (N_8734,N_5837,N_7468);
nor U8735 (N_8735,N_7483,N_5172);
xnor U8736 (N_8736,N_6871,N_7430);
and U8737 (N_8737,N_7229,N_7146);
and U8738 (N_8738,N_6130,N_6171);
nor U8739 (N_8739,N_5585,N_6789);
or U8740 (N_8740,N_7442,N_5676);
and U8741 (N_8741,N_5639,N_6196);
or U8742 (N_8742,N_5591,N_6296);
xnor U8743 (N_8743,N_7493,N_5869);
and U8744 (N_8744,N_5834,N_7015);
and U8745 (N_8745,N_7182,N_6181);
xor U8746 (N_8746,N_6535,N_6217);
or U8747 (N_8747,N_5583,N_5408);
and U8748 (N_8748,N_5144,N_5518);
xnor U8749 (N_8749,N_5563,N_7309);
or U8750 (N_8750,N_6862,N_5662);
and U8751 (N_8751,N_6147,N_7149);
nand U8752 (N_8752,N_5099,N_5119);
or U8753 (N_8753,N_7045,N_7402);
nor U8754 (N_8754,N_6538,N_7307);
nor U8755 (N_8755,N_5232,N_6723);
or U8756 (N_8756,N_6602,N_5187);
nor U8757 (N_8757,N_5373,N_6535);
xor U8758 (N_8758,N_7310,N_5365);
or U8759 (N_8759,N_5826,N_7070);
nand U8760 (N_8760,N_5775,N_6526);
nor U8761 (N_8761,N_7051,N_5675);
xor U8762 (N_8762,N_6034,N_6164);
nand U8763 (N_8763,N_5851,N_5573);
nand U8764 (N_8764,N_5658,N_6086);
xor U8765 (N_8765,N_7211,N_6600);
or U8766 (N_8766,N_6392,N_6171);
xor U8767 (N_8767,N_5334,N_5691);
nand U8768 (N_8768,N_6918,N_5890);
or U8769 (N_8769,N_7187,N_5439);
xnor U8770 (N_8770,N_6756,N_6772);
nand U8771 (N_8771,N_7025,N_5410);
xor U8772 (N_8772,N_5463,N_7421);
nor U8773 (N_8773,N_6699,N_6406);
nand U8774 (N_8774,N_7149,N_5891);
or U8775 (N_8775,N_7395,N_5598);
xor U8776 (N_8776,N_5791,N_6690);
xor U8777 (N_8777,N_5820,N_6355);
nor U8778 (N_8778,N_6521,N_7076);
and U8779 (N_8779,N_5387,N_6264);
and U8780 (N_8780,N_5418,N_7434);
or U8781 (N_8781,N_6717,N_5277);
nor U8782 (N_8782,N_6276,N_5443);
nand U8783 (N_8783,N_7162,N_5735);
xor U8784 (N_8784,N_5283,N_5538);
nor U8785 (N_8785,N_6331,N_6205);
xnor U8786 (N_8786,N_6200,N_6592);
nor U8787 (N_8787,N_7413,N_5508);
xnor U8788 (N_8788,N_5790,N_5176);
or U8789 (N_8789,N_6100,N_6931);
and U8790 (N_8790,N_6176,N_5260);
and U8791 (N_8791,N_7213,N_6803);
and U8792 (N_8792,N_6982,N_7277);
or U8793 (N_8793,N_5911,N_5121);
nand U8794 (N_8794,N_6391,N_6506);
nor U8795 (N_8795,N_5920,N_5122);
and U8796 (N_8796,N_6390,N_7236);
nor U8797 (N_8797,N_6751,N_6789);
or U8798 (N_8798,N_6513,N_6461);
nor U8799 (N_8799,N_5264,N_6652);
or U8800 (N_8800,N_6457,N_7281);
nand U8801 (N_8801,N_5853,N_6350);
and U8802 (N_8802,N_5691,N_6927);
nor U8803 (N_8803,N_6196,N_6432);
nand U8804 (N_8804,N_6261,N_6881);
nand U8805 (N_8805,N_7120,N_7311);
nand U8806 (N_8806,N_7375,N_6917);
nor U8807 (N_8807,N_7305,N_5636);
nand U8808 (N_8808,N_5443,N_5986);
nor U8809 (N_8809,N_6656,N_6132);
and U8810 (N_8810,N_6895,N_7461);
and U8811 (N_8811,N_6321,N_6105);
nor U8812 (N_8812,N_5392,N_5013);
nand U8813 (N_8813,N_6798,N_6481);
or U8814 (N_8814,N_5655,N_6520);
and U8815 (N_8815,N_6016,N_7417);
xnor U8816 (N_8816,N_5347,N_6842);
and U8817 (N_8817,N_5680,N_5156);
nand U8818 (N_8818,N_5866,N_7157);
and U8819 (N_8819,N_5565,N_6713);
nand U8820 (N_8820,N_5329,N_5041);
or U8821 (N_8821,N_7064,N_6643);
or U8822 (N_8822,N_7408,N_6927);
xor U8823 (N_8823,N_6706,N_7011);
nor U8824 (N_8824,N_5168,N_5576);
nand U8825 (N_8825,N_6036,N_6295);
xor U8826 (N_8826,N_7434,N_5594);
xor U8827 (N_8827,N_6410,N_6206);
xnor U8828 (N_8828,N_6072,N_6830);
nor U8829 (N_8829,N_7402,N_7029);
nand U8830 (N_8830,N_5722,N_5630);
nor U8831 (N_8831,N_6315,N_6404);
and U8832 (N_8832,N_5979,N_5791);
xor U8833 (N_8833,N_5301,N_5363);
nor U8834 (N_8834,N_5950,N_6551);
and U8835 (N_8835,N_5315,N_6313);
or U8836 (N_8836,N_5135,N_5232);
nand U8837 (N_8837,N_5285,N_6165);
nand U8838 (N_8838,N_6575,N_6084);
nand U8839 (N_8839,N_5702,N_5616);
and U8840 (N_8840,N_6355,N_7417);
nor U8841 (N_8841,N_7091,N_6392);
nor U8842 (N_8842,N_5366,N_6254);
xnor U8843 (N_8843,N_5220,N_6570);
xnor U8844 (N_8844,N_6127,N_5229);
or U8845 (N_8845,N_5874,N_6382);
or U8846 (N_8846,N_6602,N_5944);
nand U8847 (N_8847,N_5485,N_6718);
or U8848 (N_8848,N_6716,N_6002);
and U8849 (N_8849,N_5186,N_7073);
nand U8850 (N_8850,N_6928,N_5626);
xor U8851 (N_8851,N_7282,N_5174);
nor U8852 (N_8852,N_7406,N_5443);
and U8853 (N_8853,N_5606,N_6251);
xor U8854 (N_8854,N_6084,N_6304);
and U8855 (N_8855,N_6952,N_6777);
nand U8856 (N_8856,N_5239,N_7208);
nor U8857 (N_8857,N_5765,N_6946);
nor U8858 (N_8858,N_6946,N_6048);
or U8859 (N_8859,N_7131,N_5889);
or U8860 (N_8860,N_7282,N_5106);
nand U8861 (N_8861,N_7143,N_6885);
nand U8862 (N_8862,N_6920,N_7064);
nand U8863 (N_8863,N_6042,N_5086);
nand U8864 (N_8864,N_6053,N_7147);
nand U8865 (N_8865,N_6339,N_7226);
nor U8866 (N_8866,N_6431,N_7239);
nand U8867 (N_8867,N_6386,N_6354);
or U8868 (N_8868,N_5142,N_5905);
and U8869 (N_8869,N_5053,N_5174);
and U8870 (N_8870,N_5874,N_5292);
nor U8871 (N_8871,N_5359,N_5241);
nor U8872 (N_8872,N_5594,N_5962);
xor U8873 (N_8873,N_6425,N_6811);
nor U8874 (N_8874,N_5569,N_7370);
xnor U8875 (N_8875,N_6926,N_7413);
and U8876 (N_8876,N_7298,N_5975);
xor U8877 (N_8877,N_7016,N_6634);
xnor U8878 (N_8878,N_7108,N_5656);
xnor U8879 (N_8879,N_6217,N_6775);
xnor U8880 (N_8880,N_5829,N_6672);
and U8881 (N_8881,N_5553,N_5949);
nor U8882 (N_8882,N_5545,N_5308);
and U8883 (N_8883,N_6573,N_7004);
nor U8884 (N_8884,N_6197,N_7472);
and U8885 (N_8885,N_6133,N_5001);
and U8886 (N_8886,N_5318,N_6819);
xor U8887 (N_8887,N_7017,N_5333);
and U8888 (N_8888,N_5758,N_5342);
xor U8889 (N_8889,N_6817,N_5974);
or U8890 (N_8890,N_5613,N_7201);
nor U8891 (N_8891,N_5234,N_5967);
nor U8892 (N_8892,N_6007,N_6891);
or U8893 (N_8893,N_6824,N_5433);
and U8894 (N_8894,N_6435,N_7069);
nand U8895 (N_8895,N_7029,N_6540);
or U8896 (N_8896,N_7487,N_5125);
xor U8897 (N_8897,N_7026,N_6614);
nor U8898 (N_8898,N_6099,N_5947);
and U8899 (N_8899,N_7390,N_6642);
xor U8900 (N_8900,N_5246,N_5824);
and U8901 (N_8901,N_6034,N_7350);
and U8902 (N_8902,N_6554,N_7408);
nor U8903 (N_8903,N_5133,N_5722);
nor U8904 (N_8904,N_5422,N_6598);
xor U8905 (N_8905,N_5559,N_6476);
nor U8906 (N_8906,N_6936,N_6365);
xnor U8907 (N_8907,N_6249,N_6760);
nor U8908 (N_8908,N_5261,N_5295);
or U8909 (N_8909,N_6221,N_5068);
and U8910 (N_8910,N_6678,N_6114);
nand U8911 (N_8911,N_6805,N_5783);
or U8912 (N_8912,N_7071,N_5971);
nand U8913 (N_8913,N_7074,N_7472);
nand U8914 (N_8914,N_7436,N_6257);
xor U8915 (N_8915,N_5983,N_7199);
or U8916 (N_8916,N_5281,N_5936);
and U8917 (N_8917,N_6472,N_6969);
and U8918 (N_8918,N_7089,N_5531);
nor U8919 (N_8919,N_5207,N_5123);
nand U8920 (N_8920,N_7355,N_5323);
nand U8921 (N_8921,N_6923,N_5537);
xnor U8922 (N_8922,N_6007,N_7086);
nand U8923 (N_8923,N_5096,N_6199);
and U8924 (N_8924,N_5048,N_6167);
xnor U8925 (N_8925,N_5647,N_6593);
nor U8926 (N_8926,N_6637,N_6726);
and U8927 (N_8927,N_7333,N_6770);
nor U8928 (N_8928,N_7043,N_6692);
and U8929 (N_8929,N_5990,N_6047);
or U8930 (N_8930,N_6566,N_5089);
or U8931 (N_8931,N_7282,N_6333);
or U8932 (N_8932,N_5183,N_7432);
and U8933 (N_8933,N_5136,N_5927);
nor U8934 (N_8934,N_7143,N_7089);
xnor U8935 (N_8935,N_5750,N_5131);
nor U8936 (N_8936,N_5362,N_7301);
xor U8937 (N_8937,N_5671,N_6607);
and U8938 (N_8938,N_6210,N_6465);
nor U8939 (N_8939,N_7460,N_6997);
and U8940 (N_8940,N_6927,N_5579);
xnor U8941 (N_8941,N_7039,N_5066);
xor U8942 (N_8942,N_5518,N_7377);
or U8943 (N_8943,N_5842,N_6859);
or U8944 (N_8944,N_6265,N_7380);
nor U8945 (N_8945,N_6858,N_6387);
nand U8946 (N_8946,N_7389,N_5106);
or U8947 (N_8947,N_6434,N_6877);
nand U8948 (N_8948,N_7372,N_6247);
or U8949 (N_8949,N_5976,N_6248);
xnor U8950 (N_8950,N_5339,N_6198);
or U8951 (N_8951,N_7387,N_7065);
nand U8952 (N_8952,N_7475,N_6446);
nor U8953 (N_8953,N_6900,N_6767);
or U8954 (N_8954,N_5909,N_5316);
or U8955 (N_8955,N_7055,N_5056);
nand U8956 (N_8956,N_5465,N_7379);
nor U8957 (N_8957,N_5415,N_6860);
or U8958 (N_8958,N_5345,N_6106);
xnor U8959 (N_8959,N_5033,N_7425);
and U8960 (N_8960,N_5518,N_6402);
and U8961 (N_8961,N_5655,N_7069);
nor U8962 (N_8962,N_7352,N_6749);
nor U8963 (N_8963,N_6223,N_5853);
or U8964 (N_8964,N_6738,N_5776);
and U8965 (N_8965,N_6455,N_5119);
xor U8966 (N_8966,N_5037,N_6022);
xnor U8967 (N_8967,N_5554,N_5706);
nor U8968 (N_8968,N_5782,N_5826);
xnor U8969 (N_8969,N_6478,N_5054);
nand U8970 (N_8970,N_7160,N_5539);
nand U8971 (N_8971,N_5570,N_6871);
nand U8972 (N_8972,N_7340,N_6134);
nor U8973 (N_8973,N_6001,N_6917);
nand U8974 (N_8974,N_5065,N_7311);
or U8975 (N_8975,N_5276,N_7010);
and U8976 (N_8976,N_5592,N_7305);
or U8977 (N_8977,N_6067,N_6422);
nor U8978 (N_8978,N_6403,N_5135);
nand U8979 (N_8979,N_6185,N_6960);
xor U8980 (N_8980,N_5690,N_5328);
and U8981 (N_8981,N_7236,N_5330);
xnor U8982 (N_8982,N_6028,N_6990);
xor U8983 (N_8983,N_6766,N_5803);
or U8984 (N_8984,N_6774,N_7148);
xor U8985 (N_8985,N_7141,N_6441);
nand U8986 (N_8986,N_6315,N_6464);
and U8987 (N_8987,N_5612,N_7422);
or U8988 (N_8988,N_5577,N_6647);
nand U8989 (N_8989,N_5432,N_5102);
xnor U8990 (N_8990,N_6483,N_7384);
nor U8991 (N_8991,N_5116,N_7360);
and U8992 (N_8992,N_7341,N_6495);
or U8993 (N_8993,N_5826,N_6537);
and U8994 (N_8994,N_7333,N_6668);
nor U8995 (N_8995,N_6595,N_5454);
or U8996 (N_8996,N_6885,N_5033);
xor U8997 (N_8997,N_5713,N_5957);
nand U8998 (N_8998,N_6028,N_6350);
nand U8999 (N_8999,N_6402,N_5708);
xor U9000 (N_9000,N_6864,N_5503);
and U9001 (N_9001,N_6518,N_7022);
or U9002 (N_9002,N_5456,N_6980);
and U9003 (N_9003,N_7247,N_6148);
or U9004 (N_9004,N_6717,N_7005);
and U9005 (N_9005,N_7385,N_7494);
and U9006 (N_9006,N_6297,N_7398);
or U9007 (N_9007,N_6847,N_5782);
and U9008 (N_9008,N_5073,N_6586);
and U9009 (N_9009,N_7433,N_5065);
and U9010 (N_9010,N_5775,N_6405);
nand U9011 (N_9011,N_7073,N_6390);
or U9012 (N_9012,N_6586,N_5128);
nand U9013 (N_9013,N_5075,N_7446);
xnor U9014 (N_9014,N_7143,N_5058);
and U9015 (N_9015,N_7132,N_5201);
and U9016 (N_9016,N_7399,N_6029);
nand U9017 (N_9017,N_5097,N_6810);
nor U9018 (N_9018,N_6236,N_5466);
or U9019 (N_9019,N_5294,N_5730);
nor U9020 (N_9020,N_6267,N_7010);
xor U9021 (N_9021,N_5017,N_6947);
xor U9022 (N_9022,N_6832,N_5395);
or U9023 (N_9023,N_6659,N_5336);
nor U9024 (N_9024,N_7428,N_7219);
and U9025 (N_9025,N_6788,N_5127);
nand U9026 (N_9026,N_5134,N_5271);
or U9027 (N_9027,N_5080,N_5308);
or U9028 (N_9028,N_5705,N_5396);
nand U9029 (N_9029,N_6180,N_7210);
nand U9030 (N_9030,N_6460,N_5380);
nor U9031 (N_9031,N_5184,N_5781);
nor U9032 (N_9032,N_6591,N_5456);
or U9033 (N_9033,N_5058,N_5321);
nor U9034 (N_9034,N_6514,N_5632);
xor U9035 (N_9035,N_5568,N_6232);
nand U9036 (N_9036,N_6866,N_5217);
nor U9037 (N_9037,N_6519,N_6934);
nor U9038 (N_9038,N_5861,N_5485);
or U9039 (N_9039,N_5673,N_5924);
xnor U9040 (N_9040,N_5598,N_6011);
nor U9041 (N_9041,N_7383,N_5830);
xor U9042 (N_9042,N_5605,N_6263);
and U9043 (N_9043,N_7230,N_6814);
nor U9044 (N_9044,N_6622,N_7270);
and U9045 (N_9045,N_6317,N_6482);
or U9046 (N_9046,N_7405,N_7450);
or U9047 (N_9047,N_5876,N_5622);
xor U9048 (N_9048,N_6873,N_5078);
xnor U9049 (N_9049,N_5508,N_7107);
and U9050 (N_9050,N_6822,N_6877);
nor U9051 (N_9051,N_7108,N_7063);
nand U9052 (N_9052,N_6857,N_5262);
nor U9053 (N_9053,N_5015,N_6821);
and U9054 (N_9054,N_6044,N_7326);
and U9055 (N_9055,N_6092,N_7453);
nand U9056 (N_9056,N_6949,N_5938);
xnor U9057 (N_9057,N_6152,N_6281);
nor U9058 (N_9058,N_6506,N_6081);
xnor U9059 (N_9059,N_5752,N_6571);
and U9060 (N_9060,N_6378,N_6264);
or U9061 (N_9061,N_5508,N_6264);
and U9062 (N_9062,N_6562,N_7155);
nand U9063 (N_9063,N_7353,N_7106);
nor U9064 (N_9064,N_5153,N_6242);
nand U9065 (N_9065,N_5346,N_6170);
nand U9066 (N_9066,N_5988,N_5937);
or U9067 (N_9067,N_7115,N_6405);
nor U9068 (N_9068,N_5601,N_5800);
nor U9069 (N_9069,N_7377,N_7239);
nand U9070 (N_9070,N_7009,N_5842);
nand U9071 (N_9071,N_6724,N_5293);
or U9072 (N_9072,N_5822,N_7187);
nor U9073 (N_9073,N_5197,N_5841);
or U9074 (N_9074,N_5166,N_6462);
nor U9075 (N_9075,N_6583,N_7306);
or U9076 (N_9076,N_7269,N_7131);
and U9077 (N_9077,N_5970,N_5400);
nor U9078 (N_9078,N_6827,N_7328);
nand U9079 (N_9079,N_6267,N_5498);
nor U9080 (N_9080,N_6571,N_6696);
nor U9081 (N_9081,N_7420,N_7267);
or U9082 (N_9082,N_7382,N_5859);
and U9083 (N_9083,N_5090,N_6630);
or U9084 (N_9084,N_5618,N_5085);
nor U9085 (N_9085,N_6463,N_5647);
xnor U9086 (N_9086,N_7058,N_5845);
xor U9087 (N_9087,N_7011,N_5178);
nand U9088 (N_9088,N_6556,N_5142);
or U9089 (N_9089,N_5584,N_6475);
xnor U9090 (N_9090,N_6003,N_5938);
nor U9091 (N_9091,N_5281,N_5824);
nand U9092 (N_9092,N_6077,N_5144);
xnor U9093 (N_9093,N_6984,N_6943);
xor U9094 (N_9094,N_7028,N_5159);
xor U9095 (N_9095,N_7158,N_6612);
and U9096 (N_9096,N_5781,N_6705);
nand U9097 (N_9097,N_5422,N_6018);
nor U9098 (N_9098,N_6742,N_5141);
and U9099 (N_9099,N_5393,N_5333);
nand U9100 (N_9100,N_6925,N_7187);
nor U9101 (N_9101,N_6286,N_7294);
or U9102 (N_9102,N_5226,N_5120);
or U9103 (N_9103,N_6102,N_7412);
or U9104 (N_9104,N_5319,N_5690);
xnor U9105 (N_9105,N_6837,N_5442);
nand U9106 (N_9106,N_6365,N_5137);
and U9107 (N_9107,N_5684,N_5928);
nand U9108 (N_9108,N_6495,N_6096);
nor U9109 (N_9109,N_6982,N_5572);
or U9110 (N_9110,N_6865,N_6304);
nor U9111 (N_9111,N_6040,N_5061);
and U9112 (N_9112,N_6690,N_6559);
nor U9113 (N_9113,N_5676,N_6393);
nor U9114 (N_9114,N_5250,N_6841);
xor U9115 (N_9115,N_6126,N_7011);
nand U9116 (N_9116,N_6202,N_5704);
or U9117 (N_9117,N_6254,N_6263);
xor U9118 (N_9118,N_5803,N_5566);
and U9119 (N_9119,N_5571,N_6735);
and U9120 (N_9120,N_7027,N_6041);
nor U9121 (N_9121,N_7271,N_6575);
and U9122 (N_9122,N_5405,N_5011);
nor U9123 (N_9123,N_6921,N_5415);
or U9124 (N_9124,N_5771,N_6878);
or U9125 (N_9125,N_6488,N_5313);
nand U9126 (N_9126,N_5402,N_5517);
or U9127 (N_9127,N_5147,N_5365);
nand U9128 (N_9128,N_5904,N_5121);
xor U9129 (N_9129,N_6774,N_5129);
nand U9130 (N_9130,N_6408,N_5573);
nor U9131 (N_9131,N_6882,N_7186);
xnor U9132 (N_9132,N_5986,N_5425);
or U9133 (N_9133,N_7384,N_5309);
nor U9134 (N_9134,N_5679,N_5000);
and U9135 (N_9135,N_6426,N_5012);
or U9136 (N_9136,N_6830,N_6999);
nand U9137 (N_9137,N_6646,N_5088);
nor U9138 (N_9138,N_5900,N_7221);
and U9139 (N_9139,N_5653,N_6184);
nor U9140 (N_9140,N_6748,N_7035);
xor U9141 (N_9141,N_6579,N_5661);
and U9142 (N_9142,N_5088,N_5916);
nand U9143 (N_9143,N_7210,N_5774);
nor U9144 (N_9144,N_5645,N_6755);
nand U9145 (N_9145,N_6696,N_7320);
nor U9146 (N_9146,N_7312,N_5973);
or U9147 (N_9147,N_7342,N_7169);
or U9148 (N_9148,N_6576,N_6235);
and U9149 (N_9149,N_5118,N_7255);
or U9150 (N_9150,N_7204,N_6689);
and U9151 (N_9151,N_6933,N_6287);
and U9152 (N_9152,N_5303,N_5265);
and U9153 (N_9153,N_6901,N_6674);
nor U9154 (N_9154,N_6657,N_6009);
nand U9155 (N_9155,N_5036,N_5657);
xnor U9156 (N_9156,N_6586,N_5854);
nand U9157 (N_9157,N_5699,N_5298);
nand U9158 (N_9158,N_6667,N_5313);
and U9159 (N_9159,N_5448,N_5115);
and U9160 (N_9160,N_6810,N_5106);
and U9161 (N_9161,N_6598,N_6990);
nand U9162 (N_9162,N_5304,N_6171);
xnor U9163 (N_9163,N_6183,N_7163);
nor U9164 (N_9164,N_5480,N_7014);
nand U9165 (N_9165,N_6314,N_5183);
or U9166 (N_9166,N_6604,N_6267);
nand U9167 (N_9167,N_5167,N_6165);
xor U9168 (N_9168,N_7184,N_5111);
nand U9169 (N_9169,N_7158,N_7245);
nor U9170 (N_9170,N_7183,N_7082);
nor U9171 (N_9171,N_6514,N_6917);
or U9172 (N_9172,N_5719,N_5770);
and U9173 (N_9173,N_7473,N_5278);
nor U9174 (N_9174,N_5765,N_6992);
or U9175 (N_9175,N_5722,N_6676);
nand U9176 (N_9176,N_6670,N_5776);
or U9177 (N_9177,N_5001,N_5873);
xor U9178 (N_9178,N_7206,N_6851);
or U9179 (N_9179,N_6221,N_6184);
nand U9180 (N_9180,N_7336,N_7194);
and U9181 (N_9181,N_6396,N_5932);
xor U9182 (N_9182,N_5535,N_6755);
and U9183 (N_9183,N_7281,N_5698);
nor U9184 (N_9184,N_5603,N_5309);
nor U9185 (N_9185,N_7001,N_7194);
nor U9186 (N_9186,N_7363,N_5731);
nand U9187 (N_9187,N_5365,N_5006);
or U9188 (N_9188,N_5553,N_6442);
and U9189 (N_9189,N_6089,N_6698);
nor U9190 (N_9190,N_6750,N_6570);
or U9191 (N_9191,N_5757,N_5042);
nand U9192 (N_9192,N_5267,N_5715);
nand U9193 (N_9193,N_5890,N_6321);
and U9194 (N_9194,N_6728,N_7064);
xnor U9195 (N_9195,N_6234,N_7165);
and U9196 (N_9196,N_7096,N_7260);
or U9197 (N_9197,N_5329,N_5509);
nor U9198 (N_9198,N_5277,N_6118);
nor U9199 (N_9199,N_6362,N_6915);
or U9200 (N_9200,N_6408,N_5600);
and U9201 (N_9201,N_5591,N_5936);
nor U9202 (N_9202,N_6189,N_5367);
nand U9203 (N_9203,N_6949,N_5151);
or U9204 (N_9204,N_5630,N_7100);
nand U9205 (N_9205,N_7488,N_6748);
xnor U9206 (N_9206,N_5523,N_5143);
nor U9207 (N_9207,N_7380,N_5575);
nor U9208 (N_9208,N_5354,N_6542);
xor U9209 (N_9209,N_6596,N_6628);
or U9210 (N_9210,N_7093,N_6245);
and U9211 (N_9211,N_5337,N_6428);
nand U9212 (N_9212,N_6549,N_5037);
nand U9213 (N_9213,N_6829,N_5150);
or U9214 (N_9214,N_5989,N_5506);
nor U9215 (N_9215,N_7171,N_6526);
or U9216 (N_9216,N_5465,N_6918);
nor U9217 (N_9217,N_5864,N_5472);
nor U9218 (N_9218,N_5227,N_5988);
xor U9219 (N_9219,N_6214,N_5104);
or U9220 (N_9220,N_5342,N_7215);
or U9221 (N_9221,N_5471,N_5473);
xnor U9222 (N_9222,N_5795,N_7105);
and U9223 (N_9223,N_6263,N_6182);
nand U9224 (N_9224,N_7471,N_7491);
nand U9225 (N_9225,N_5560,N_6747);
nor U9226 (N_9226,N_5569,N_7324);
nor U9227 (N_9227,N_6259,N_6211);
nand U9228 (N_9228,N_6788,N_5405);
nor U9229 (N_9229,N_6608,N_7358);
xnor U9230 (N_9230,N_5651,N_6061);
nor U9231 (N_9231,N_6024,N_5202);
and U9232 (N_9232,N_5167,N_5026);
xor U9233 (N_9233,N_7443,N_7115);
or U9234 (N_9234,N_5016,N_5039);
or U9235 (N_9235,N_6072,N_5561);
and U9236 (N_9236,N_6973,N_6779);
or U9237 (N_9237,N_6098,N_5408);
nor U9238 (N_9238,N_6122,N_6495);
nand U9239 (N_9239,N_5921,N_5899);
or U9240 (N_9240,N_6725,N_6973);
and U9241 (N_9241,N_6416,N_6461);
xnor U9242 (N_9242,N_6946,N_5196);
and U9243 (N_9243,N_6986,N_7133);
and U9244 (N_9244,N_5183,N_6971);
nand U9245 (N_9245,N_7319,N_6630);
and U9246 (N_9246,N_6624,N_6723);
or U9247 (N_9247,N_6649,N_6070);
nand U9248 (N_9248,N_6948,N_6706);
and U9249 (N_9249,N_7471,N_6094);
and U9250 (N_9250,N_6107,N_7147);
and U9251 (N_9251,N_6813,N_7261);
nand U9252 (N_9252,N_7388,N_5924);
xnor U9253 (N_9253,N_6002,N_5193);
nor U9254 (N_9254,N_5713,N_7134);
xnor U9255 (N_9255,N_7468,N_7145);
and U9256 (N_9256,N_5652,N_5077);
xor U9257 (N_9257,N_6607,N_6735);
xnor U9258 (N_9258,N_5533,N_5180);
xor U9259 (N_9259,N_5335,N_6282);
and U9260 (N_9260,N_6693,N_6468);
xnor U9261 (N_9261,N_6294,N_6478);
xor U9262 (N_9262,N_7017,N_7117);
or U9263 (N_9263,N_5144,N_6482);
nand U9264 (N_9264,N_5679,N_5524);
nor U9265 (N_9265,N_5065,N_6678);
and U9266 (N_9266,N_7282,N_5871);
or U9267 (N_9267,N_7005,N_5531);
nand U9268 (N_9268,N_7136,N_6423);
and U9269 (N_9269,N_7385,N_5077);
nand U9270 (N_9270,N_7095,N_5562);
and U9271 (N_9271,N_7154,N_6567);
and U9272 (N_9272,N_6122,N_6878);
nor U9273 (N_9273,N_5809,N_7146);
and U9274 (N_9274,N_6987,N_5509);
xnor U9275 (N_9275,N_7446,N_5225);
xnor U9276 (N_9276,N_5602,N_5797);
or U9277 (N_9277,N_6712,N_5001);
nor U9278 (N_9278,N_7431,N_6138);
or U9279 (N_9279,N_6896,N_5795);
or U9280 (N_9280,N_5567,N_5556);
or U9281 (N_9281,N_6864,N_5857);
nand U9282 (N_9282,N_6303,N_5181);
xor U9283 (N_9283,N_5134,N_6350);
nor U9284 (N_9284,N_7361,N_5454);
xnor U9285 (N_9285,N_6158,N_5811);
or U9286 (N_9286,N_5309,N_6691);
nand U9287 (N_9287,N_6458,N_6680);
and U9288 (N_9288,N_6739,N_5280);
nor U9289 (N_9289,N_6993,N_6309);
or U9290 (N_9290,N_6111,N_6165);
nor U9291 (N_9291,N_5309,N_6820);
nand U9292 (N_9292,N_7332,N_5751);
nor U9293 (N_9293,N_7216,N_5227);
or U9294 (N_9294,N_7260,N_5673);
and U9295 (N_9295,N_5804,N_5601);
or U9296 (N_9296,N_6547,N_5436);
xnor U9297 (N_9297,N_6014,N_5098);
nor U9298 (N_9298,N_6194,N_5415);
nor U9299 (N_9299,N_5645,N_5823);
xnor U9300 (N_9300,N_6138,N_5632);
and U9301 (N_9301,N_5156,N_6890);
xnor U9302 (N_9302,N_5541,N_5168);
or U9303 (N_9303,N_5863,N_6114);
xnor U9304 (N_9304,N_7479,N_6289);
nor U9305 (N_9305,N_5673,N_6066);
or U9306 (N_9306,N_6285,N_6329);
nand U9307 (N_9307,N_6512,N_5517);
or U9308 (N_9308,N_7114,N_7428);
or U9309 (N_9309,N_5193,N_5098);
and U9310 (N_9310,N_6516,N_6412);
xor U9311 (N_9311,N_6438,N_5237);
nor U9312 (N_9312,N_5589,N_7177);
nand U9313 (N_9313,N_5118,N_6471);
and U9314 (N_9314,N_7470,N_6034);
and U9315 (N_9315,N_5966,N_6690);
and U9316 (N_9316,N_6770,N_5496);
and U9317 (N_9317,N_6817,N_5930);
nor U9318 (N_9318,N_7225,N_6106);
xor U9319 (N_9319,N_7278,N_5709);
or U9320 (N_9320,N_7404,N_6809);
and U9321 (N_9321,N_5806,N_7464);
nand U9322 (N_9322,N_6276,N_6378);
and U9323 (N_9323,N_7315,N_6706);
or U9324 (N_9324,N_6722,N_5160);
nand U9325 (N_9325,N_6261,N_7476);
xor U9326 (N_9326,N_6254,N_6918);
and U9327 (N_9327,N_7015,N_7428);
xnor U9328 (N_9328,N_5232,N_5498);
xor U9329 (N_9329,N_7312,N_6013);
nor U9330 (N_9330,N_6094,N_7069);
xor U9331 (N_9331,N_6542,N_5735);
nor U9332 (N_9332,N_6354,N_5290);
or U9333 (N_9333,N_5323,N_6302);
xnor U9334 (N_9334,N_5153,N_7236);
xnor U9335 (N_9335,N_6908,N_6255);
or U9336 (N_9336,N_5624,N_6172);
xnor U9337 (N_9337,N_5119,N_6655);
or U9338 (N_9338,N_5351,N_5822);
or U9339 (N_9339,N_5277,N_5443);
and U9340 (N_9340,N_5387,N_5076);
xor U9341 (N_9341,N_5213,N_5917);
xnor U9342 (N_9342,N_5905,N_7499);
nand U9343 (N_9343,N_5462,N_6099);
or U9344 (N_9344,N_5191,N_5587);
or U9345 (N_9345,N_5985,N_5612);
xnor U9346 (N_9346,N_5321,N_5005);
nor U9347 (N_9347,N_6747,N_5756);
nor U9348 (N_9348,N_6140,N_5797);
xor U9349 (N_9349,N_6858,N_6378);
nand U9350 (N_9350,N_5302,N_6156);
and U9351 (N_9351,N_6535,N_6106);
nand U9352 (N_9352,N_6722,N_6509);
xor U9353 (N_9353,N_6985,N_5953);
xnor U9354 (N_9354,N_5481,N_7139);
nor U9355 (N_9355,N_6555,N_5991);
xor U9356 (N_9356,N_7287,N_5260);
or U9357 (N_9357,N_7170,N_6406);
and U9358 (N_9358,N_5234,N_6543);
nor U9359 (N_9359,N_6698,N_7039);
and U9360 (N_9360,N_6663,N_5227);
nor U9361 (N_9361,N_7389,N_5877);
nand U9362 (N_9362,N_7204,N_6805);
nand U9363 (N_9363,N_6493,N_6025);
or U9364 (N_9364,N_7009,N_5600);
and U9365 (N_9365,N_6825,N_6983);
nand U9366 (N_9366,N_7192,N_6239);
nor U9367 (N_9367,N_5044,N_5540);
xor U9368 (N_9368,N_6694,N_5745);
nor U9369 (N_9369,N_7217,N_6604);
xor U9370 (N_9370,N_5889,N_6324);
xor U9371 (N_9371,N_7492,N_5513);
and U9372 (N_9372,N_5543,N_5616);
nor U9373 (N_9373,N_5170,N_6806);
xnor U9374 (N_9374,N_6168,N_6296);
nand U9375 (N_9375,N_7073,N_5434);
or U9376 (N_9376,N_5738,N_7160);
and U9377 (N_9377,N_7099,N_5055);
nand U9378 (N_9378,N_5287,N_5925);
and U9379 (N_9379,N_6624,N_5268);
xnor U9380 (N_9380,N_7192,N_5120);
or U9381 (N_9381,N_5190,N_5778);
nand U9382 (N_9382,N_7388,N_6808);
nor U9383 (N_9383,N_5206,N_7387);
and U9384 (N_9384,N_5060,N_6152);
or U9385 (N_9385,N_7358,N_6495);
and U9386 (N_9386,N_6173,N_6910);
nand U9387 (N_9387,N_5654,N_5834);
nand U9388 (N_9388,N_6054,N_7464);
and U9389 (N_9389,N_6770,N_7393);
and U9390 (N_9390,N_5101,N_5581);
nand U9391 (N_9391,N_7423,N_7110);
xnor U9392 (N_9392,N_6810,N_7296);
or U9393 (N_9393,N_6695,N_7325);
xnor U9394 (N_9394,N_6687,N_7340);
and U9395 (N_9395,N_6226,N_6932);
xor U9396 (N_9396,N_5205,N_6373);
nor U9397 (N_9397,N_6671,N_5053);
nand U9398 (N_9398,N_6553,N_5304);
nand U9399 (N_9399,N_5029,N_6136);
and U9400 (N_9400,N_6295,N_7315);
or U9401 (N_9401,N_6331,N_5874);
xor U9402 (N_9402,N_5107,N_5423);
or U9403 (N_9403,N_6605,N_5253);
and U9404 (N_9404,N_7216,N_6982);
and U9405 (N_9405,N_5222,N_5503);
or U9406 (N_9406,N_6420,N_6508);
nand U9407 (N_9407,N_6566,N_5570);
xnor U9408 (N_9408,N_6563,N_5140);
and U9409 (N_9409,N_6035,N_5737);
nand U9410 (N_9410,N_7187,N_7428);
or U9411 (N_9411,N_5985,N_6991);
or U9412 (N_9412,N_6441,N_5595);
nor U9413 (N_9413,N_5962,N_5784);
and U9414 (N_9414,N_5635,N_5765);
and U9415 (N_9415,N_7429,N_6947);
nor U9416 (N_9416,N_6848,N_5380);
or U9417 (N_9417,N_5992,N_5619);
nor U9418 (N_9418,N_7390,N_7140);
nor U9419 (N_9419,N_5808,N_5068);
nand U9420 (N_9420,N_5851,N_5506);
and U9421 (N_9421,N_5274,N_6310);
xnor U9422 (N_9422,N_5492,N_5312);
nand U9423 (N_9423,N_5569,N_6784);
xor U9424 (N_9424,N_7024,N_7014);
nor U9425 (N_9425,N_6796,N_5193);
and U9426 (N_9426,N_6461,N_6298);
or U9427 (N_9427,N_7354,N_5295);
nand U9428 (N_9428,N_6513,N_7039);
or U9429 (N_9429,N_6047,N_6128);
nand U9430 (N_9430,N_6908,N_6330);
and U9431 (N_9431,N_6022,N_5124);
xnor U9432 (N_9432,N_6512,N_5511);
or U9433 (N_9433,N_5566,N_7413);
and U9434 (N_9434,N_5208,N_6079);
xnor U9435 (N_9435,N_5512,N_5283);
xnor U9436 (N_9436,N_6473,N_6751);
or U9437 (N_9437,N_7155,N_6240);
and U9438 (N_9438,N_7409,N_6392);
or U9439 (N_9439,N_6729,N_7107);
xnor U9440 (N_9440,N_7209,N_6321);
or U9441 (N_9441,N_5913,N_5632);
and U9442 (N_9442,N_5517,N_5343);
and U9443 (N_9443,N_6387,N_6970);
xor U9444 (N_9444,N_7299,N_6373);
xnor U9445 (N_9445,N_5966,N_6871);
xor U9446 (N_9446,N_6645,N_5524);
nand U9447 (N_9447,N_6337,N_7147);
and U9448 (N_9448,N_6634,N_5398);
or U9449 (N_9449,N_7058,N_5432);
xnor U9450 (N_9450,N_5328,N_6112);
nand U9451 (N_9451,N_5344,N_5971);
nor U9452 (N_9452,N_5739,N_6895);
or U9453 (N_9453,N_7244,N_5788);
nor U9454 (N_9454,N_5611,N_5954);
and U9455 (N_9455,N_7235,N_7497);
or U9456 (N_9456,N_6366,N_5899);
or U9457 (N_9457,N_5915,N_5868);
and U9458 (N_9458,N_5726,N_5604);
nand U9459 (N_9459,N_6198,N_5900);
nor U9460 (N_9460,N_6641,N_6020);
and U9461 (N_9461,N_5254,N_6109);
nor U9462 (N_9462,N_6234,N_7315);
or U9463 (N_9463,N_6062,N_7258);
or U9464 (N_9464,N_5171,N_7206);
nor U9465 (N_9465,N_6583,N_6154);
nor U9466 (N_9466,N_5912,N_5369);
or U9467 (N_9467,N_6008,N_6039);
nand U9468 (N_9468,N_5998,N_6625);
and U9469 (N_9469,N_5603,N_7067);
or U9470 (N_9470,N_7097,N_5184);
nand U9471 (N_9471,N_6856,N_6315);
or U9472 (N_9472,N_5306,N_5562);
nor U9473 (N_9473,N_5138,N_7201);
and U9474 (N_9474,N_6669,N_5160);
or U9475 (N_9475,N_5563,N_6718);
or U9476 (N_9476,N_6550,N_6051);
nor U9477 (N_9477,N_5505,N_7263);
nand U9478 (N_9478,N_7470,N_6254);
nand U9479 (N_9479,N_5447,N_5763);
nand U9480 (N_9480,N_6797,N_7110);
xor U9481 (N_9481,N_5268,N_7270);
nand U9482 (N_9482,N_5299,N_7456);
nor U9483 (N_9483,N_7287,N_5825);
nand U9484 (N_9484,N_5595,N_6608);
nand U9485 (N_9485,N_7438,N_6600);
nand U9486 (N_9486,N_6293,N_7267);
nand U9487 (N_9487,N_6386,N_6548);
or U9488 (N_9488,N_5449,N_6020);
xor U9489 (N_9489,N_6994,N_7274);
and U9490 (N_9490,N_5316,N_7345);
and U9491 (N_9491,N_5485,N_5611);
nor U9492 (N_9492,N_5041,N_6116);
nor U9493 (N_9493,N_5825,N_6001);
xnor U9494 (N_9494,N_7219,N_5042);
nand U9495 (N_9495,N_7061,N_7290);
nor U9496 (N_9496,N_7217,N_6000);
nor U9497 (N_9497,N_6609,N_5909);
xor U9498 (N_9498,N_6676,N_6046);
nand U9499 (N_9499,N_6281,N_5862);
and U9500 (N_9500,N_5721,N_5037);
or U9501 (N_9501,N_5775,N_5403);
or U9502 (N_9502,N_5639,N_6717);
xnor U9503 (N_9503,N_5390,N_7283);
nor U9504 (N_9504,N_5251,N_6812);
nor U9505 (N_9505,N_6354,N_6408);
nand U9506 (N_9506,N_7378,N_5203);
xor U9507 (N_9507,N_6466,N_5186);
or U9508 (N_9508,N_5781,N_6488);
nor U9509 (N_9509,N_6442,N_5601);
and U9510 (N_9510,N_6244,N_7295);
nand U9511 (N_9511,N_6556,N_5880);
nand U9512 (N_9512,N_7046,N_6862);
and U9513 (N_9513,N_6262,N_7057);
nor U9514 (N_9514,N_7375,N_5655);
nor U9515 (N_9515,N_7232,N_5399);
or U9516 (N_9516,N_6036,N_6731);
nand U9517 (N_9517,N_6907,N_6791);
nand U9518 (N_9518,N_5523,N_6299);
nand U9519 (N_9519,N_7160,N_6827);
and U9520 (N_9520,N_6123,N_6488);
nand U9521 (N_9521,N_5440,N_7266);
and U9522 (N_9522,N_6126,N_6320);
and U9523 (N_9523,N_5992,N_6718);
or U9524 (N_9524,N_6524,N_7467);
nor U9525 (N_9525,N_5980,N_5320);
nand U9526 (N_9526,N_7397,N_5317);
nand U9527 (N_9527,N_5640,N_6026);
nor U9528 (N_9528,N_5453,N_6047);
nand U9529 (N_9529,N_6962,N_5536);
nor U9530 (N_9530,N_5498,N_5301);
nor U9531 (N_9531,N_7426,N_5314);
nand U9532 (N_9532,N_6493,N_6305);
and U9533 (N_9533,N_6112,N_6565);
or U9534 (N_9534,N_5453,N_6278);
nor U9535 (N_9535,N_5407,N_6735);
and U9536 (N_9536,N_6255,N_6052);
nand U9537 (N_9537,N_6961,N_6369);
nand U9538 (N_9538,N_5204,N_6338);
nand U9539 (N_9539,N_7245,N_6905);
and U9540 (N_9540,N_6771,N_6998);
or U9541 (N_9541,N_5596,N_7491);
and U9542 (N_9542,N_6179,N_5362);
or U9543 (N_9543,N_5406,N_5261);
nand U9544 (N_9544,N_5874,N_5142);
nor U9545 (N_9545,N_7372,N_6328);
xnor U9546 (N_9546,N_7446,N_5368);
nor U9547 (N_9547,N_6918,N_5926);
nand U9548 (N_9548,N_6767,N_7402);
or U9549 (N_9549,N_5463,N_5301);
nor U9550 (N_9550,N_5402,N_5143);
or U9551 (N_9551,N_6138,N_7111);
xnor U9552 (N_9552,N_5828,N_7154);
and U9553 (N_9553,N_6711,N_7298);
xor U9554 (N_9554,N_6118,N_6172);
nand U9555 (N_9555,N_7390,N_5558);
or U9556 (N_9556,N_5163,N_6297);
nand U9557 (N_9557,N_6140,N_7451);
nor U9558 (N_9558,N_5386,N_7207);
nand U9559 (N_9559,N_6729,N_5237);
or U9560 (N_9560,N_5766,N_6430);
or U9561 (N_9561,N_5622,N_6327);
nand U9562 (N_9562,N_6999,N_7316);
xnor U9563 (N_9563,N_5423,N_7061);
xor U9564 (N_9564,N_7148,N_6818);
or U9565 (N_9565,N_6680,N_6465);
xnor U9566 (N_9566,N_7343,N_5620);
and U9567 (N_9567,N_5915,N_6546);
nor U9568 (N_9568,N_6025,N_6265);
or U9569 (N_9569,N_6462,N_5498);
nor U9570 (N_9570,N_6052,N_5456);
nand U9571 (N_9571,N_5104,N_6626);
and U9572 (N_9572,N_5105,N_5845);
or U9573 (N_9573,N_6799,N_5762);
xor U9574 (N_9574,N_5049,N_5505);
and U9575 (N_9575,N_5484,N_6320);
nand U9576 (N_9576,N_6614,N_6781);
and U9577 (N_9577,N_6105,N_5022);
or U9578 (N_9578,N_6177,N_5110);
nor U9579 (N_9579,N_6641,N_6240);
nand U9580 (N_9580,N_5097,N_5464);
and U9581 (N_9581,N_5920,N_5424);
xnor U9582 (N_9582,N_6704,N_6451);
nand U9583 (N_9583,N_5520,N_5630);
and U9584 (N_9584,N_5403,N_7488);
nand U9585 (N_9585,N_5399,N_7407);
nand U9586 (N_9586,N_5959,N_7331);
nand U9587 (N_9587,N_7193,N_5311);
or U9588 (N_9588,N_5896,N_5980);
nor U9589 (N_9589,N_6857,N_6370);
nand U9590 (N_9590,N_6509,N_5141);
and U9591 (N_9591,N_7200,N_6732);
and U9592 (N_9592,N_6482,N_7195);
or U9593 (N_9593,N_6630,N_6168);
nand U9594 (N_9594,N_5006,N_5585);
nand U9595 (N_9595,N_7399,N_7248);
xor U9596 (N_9596,N_7290,N_6587);
nand U9597 (N_9597,N_5363,N_6350);
nand U9598 (N_9598,N_6743,N_5166);
nand U9599 (N_9599,N_5957,N_7303);
xnor U9600 (N_9600,N_6803,N_6014);
and U9601 (N_9601,N_6618,N_7160);
or U9602 (N_9602,N_6078,N_6599);
or U9603 (N_9603,N_6949,N_5073);
and U9604 (N_9604,N_5160,N_6979);
and U9605 (N_9605,N_5061,N_5149);
xor U9606 (N_9606,N_6219,N_5215);
nor U9607 (N_9607,N_7025,N_6365);
nand U9608 (N_9608,N_5573,N_6394);
xnor U9609 (N_9609,N_5710,N_7086);
or U9610 (N_9610,N_5877,N_5012);
xnor U9611 (N_9611,N_5449,N_7371);
xnor U9612 (N_9612,N_6357,N_6316);
or U9613 (N_9613,N_5376,N_6764);
and U9614 (N_9614,N_6901,N_7496);
nand U9615 (N_9615,N_7203,N_7075);
nand U9616 (N_9616,N_5721,N_5921);
or U9617 (N_9617,N_5140,N_5740);
nand U9618 (N_9618,N_6075,N_6063);
xor U9619 (N_9619,N_5603,N_6521);
or U9620 (N_9620,N_6789,N_5469);
and U9621 (N_9621,N_5663,N_7334);
nand U9622 (N_9622,N_6836,N_6928);
or U9623 (N_9623,N_5154,N_6195);
nor U9624 (N_9624,N_5766,N_5734);
nand U9625 (N_9625,N_7221,N_7404);
or U9626 (N_9626,N_7226,N_6029);
nand U9627 (N_9627,N_5754,N_6714);
or U9628 (N_9628,N_5949,N_6650);
xnor U9629 (N_9629,N_5541,N_6354);
nand U9630 (N_9630,N_5247,N_6706);
nand U9631 (N_9631,N_6704,N_7024);
xor U9632 (N_9632,N_6261,N_5522);
xnor U9633 (N_9633,N_6240,N_5038);
nor U9634 (N_9634,N_7423,N_7106);
nor U9635 (N_9635,N_6120,N_5198);
and U9636 (N_9636,N_7405,N_6205);
or U9637 (N_9637,N_5268,N_7395);
nor U9638 (N_9638,N_5775,N_5228);
and U9639 (N_9639,N_5892,N_5156);
and U9640 (N_9640,N_6532,N_6935);
xnor U9641 (N_9641,N_6114,N_5648);
xor U9642 (N_9642,N_6779,N_5318);
xor U9643 (N_9643,N_5693,N_6412);
and U9644 (N_9644,N_7081,N_7134);
nand U9645 (N_9645,N_5699,N_5774);
nor U9646 (N_9646,N_7356,N_6531);
xor U9647 (N_9647,N_6452,N_6990);
nand U9648 (N_9648,N_6746,N_5755);
nand U9649 (N_9649,N_6065,N_7487);
and U9650 (N_9650,N_6024,N_5556);
or U9651 (N_9651,N_6072,N_7065);
or U9652 (N_9652,N_5815,N_5552);
or U9653 (N_9653,N_6052,N_7233);
xnor U9654 (N_9654,N_7256,N_6479);
xor U9655 (N_9655,N_7073,N_5717);
xnor U9656 (N_9656,N_6603,N_6900);
nand U9657 (N_9657,N_6050,N_6271);
or U9658 (N_9658,N_6701,N_6621);
and U9659 (N_9659,N_5580,N_7189);
nor U9660 (N_9660,N_5537,N_5327);
xnor U9661 (N_9661,N_6484,N_6436);
and U9662 (N_9662,N_6073,N_6016);
xnor U9663 (N_9663,N_5006,N_5544);
xnor U9664 (N_9664,N_6721,N_5077);
and U9665 (N_9665,N_5394,N_6404);
nand U9666 (N_9666,N_6730,N_5554);
nand U9667 (N_9667,N_5192,N_5318);
or U9668 (N_9668,N_5990,N_6508);
nand U9669 (N_9669,N_6678,N_5322);
or U9670 (N_9670,N_7249,N_6756);
or U9671 (N_9671,N_5068,N_6986);
nor U9672 (N_9672,N_7086,N_5246);
and U9673 (N_9673,N_5265,N_6966);
or U9674 (N_9674,N_7219,N_6427);
and U9675 (N_9675,N_6448,N_5367);
and U9676 (N_9676,N_6469,N_7063);
xor U9677 (N_9677,N_6233,N_5166);
nand U9678 (N_9678,N_7495,N_5378);
xor U9679 (N_9679,N_5143,N_7212);
nor U9680 (N_9680,N_7328,N_6625);
and U9681 (N_9681,N_6093,N_6092);
nand U9682 (N_9682,N_6150,N_6140);
nand U9683 (N_9683,N_5430,N_5214);
nand U9684 (N_9684,N_5606,N_6984);
nand U9685 (N_9685,N_6814,N_5014);
nand U9686 (N_9686,N_7426,N_6868);
nor U9687 (N_9687,N_5731,N_5192);
xnor U9688 (N_9688,N_6844,N_6526);
xor U9689 (N_9689,N_5473,N_5822);
and U9690 (N_9690,N_7205,N_5252);
or U9691 (N_9691,N_5703,N_6431);
and U9692 (N_9692,N_5843,N_5439);
or U9693 (N_9693,N_5290,N_7430);
or U9694 (N_9694,N_6541,N_5361);
nor U9695 (N_9695,N_5934,N_7102);
or U9696 (N_9696,N_7474,N_6582);
nand U9697 (N_9697,N_7176,N_5149);
or U9698 (N_9698,N_5912,N_7453);
and U9699 (N_9699,N_7394,N_5027);
nand U9700 (N_9700,N_6421,N_5127);
or U9701 (N_9701,N_5512,N_5023);
and U9702 (N_9702,N_6096,N_5125);
nor U9703 (N_9703,N_7464,N_5936);
xnor U9704 (N_9704,N_6347,N_7264);
or U9705 (N_9705,N_6630,N_5810);
or U9706 (N_9706,N_7387,N_6617);
and U9707 (N_9707,N_6399,N_6411);
xnor U9708 (N_9708,N_6348,N_7065);
xnor U9709 (N_9709,N_7382,N_7147);
xor U9710 (N_9710,N_6278,N_6898);
nand U9711 (N_9711,N_7019,N_6842);
and U9712 (N_9712,N_6774,N_6561);
or U9713 (N_9713,N_5069,N_6010);
xnor U9714 (N_9714,N_6470,N_6133);
xnor U9715 (N_9715,N_5199,N_5672);
and U9716 (N_9716,N_6647,N_5508);
and U9717 (N_9717,N_5597,N_6509);
nor U9718 (N_9718,N_7084,N_5333);
and U9719 (N_9719,N_6836,N_7374);
xor U9720 (N_9720,N_6244,N_5999);
and U9721 (N_9721,N_6595,N_7124);
xnor U9722 (N_9722,N_5819,N_5664);
or U9723 (N_9723,N_5565,N_5753);
nand U9724 (N_9724,N_5664,N_7371);
nand U9725 (N_9725,N_6205,N_7071);
nand U9726 (N_9726,N_6315,N_7418);
xor U9727 (N_9727,N_6224,N_6283);
or U9728 (N_9728,N_7295,N_7426);
xor U9729 (N_9729,N_5352,N_5906);
nor U9730 (N_9730,N_7487,N_6958);
nand U9731 (N_9731,N_7186,N_5433);
nand U9732 (N_9732,N_5684,N_5216);
nor U9733 (N_9733,N_7480,N_5523);
or U9734 (N_9734,N_6825,N_5102);
nand U9735 (N_9735,N_7250,N_6511);
or U9736 (N_9736,N_5563,N_7246);
nand U9737 (N_9737,N_6802,N_6913);
or U9738 (N_9738,N_5772,N_5608);
or U9739 (N_9739,N_7052,N_5089);
nand U9740 (N_9740,N_6288,N_5882);
nor U9741 (N_9741,N_5417,N_7353);
nand U9742 (N_9742,N_5361,N_6611);
nor U9743 (N_9743,N_6899,N_6260);
nand U9744 (N_9744,N_5741,N_6699);
nor U9745 (N_9745,N_7129,N_5882);
nor U9746 (N_9746,N_7327,N_6174);
nor U9747 (N_9747,N_6185,N_6754);
xor U9748 (N_9748,N_6321,N_5580);
and U9749 (N_9749,N_6542,N_7114);
nand U9750 (N_9750,N_5587,N_5278);
and U9751 (N_9751,N_6650,N_6088);
or U9752 (N_9752,N_6681,N_6271);
and U9753 (N_9753,N_6806,N_5614);
and U9754 (N_9754,N_5705,N_6365);
nand U9755 (N_9755,N_5452,N_6502);
nand U9756 (N_9756,N_5008,N_6091);
nand U9757 (N_9757,N_6078,N_5696);
xor U9758 (N_9758,N_5822,N_6904);
nand U9759 (N_9759,N_6215,N_6834);
or U9760 (N_9760,N_6770,N_5345);
xnor U9761 (N_9761,N_6765,N_6299);
and U9762 (N_9762,N_6135,N_6842);
and U9763 (N_9763,N_6223,N_6834);
or U9764 (N_9764,N_7132,N_7487);
or U9765 (N_9765,N_5916,N_5089);
xor U9766 (N_9766,N_6101,N_5717);
or U9767 (N_9767,N_6563,N_5906);
nand U9768 (N_9768,N_6097,N_6750);
xnor U9769 (N_9769,N_5996,N_7136);
or U9770 (N_9770,N_5216,N_5968);
nand U9771 (N_9771,N_6353,N_6062);
or U9772 (N_9772,N_6184,N_5242);
nor U9773 (N_9773,N_5035,N_6632);
nand U9774 (N_9774,N_6819,N_7136);
or U9775 (N_9775,N_5644,N_5864);
nor U9776 (N_9776,N_5897,N_5844);
or U9777 (N_9777,N_5633,N_5295);
xnor U9778 (N_9778,N_5686,N_5243);
xor U9779 (N_9779,N_6390,N_6585);
xnor U9780 (N_9780,N_6921,N_6470);
nor U9781 (N_9781,N_5433,N_5776);
and U9782 (N_9782,N_5599,N_7360);
nand U9783 (N_9783,N_7148,N_5920);
nand U9784 (N_9784,N_6422,N_6458);
and U9785 (N_9785,N_5728,N_5358);
or U9786 (N_9786,N_7300,N_6498);
xor U9787 (N_9787,N_6132,N_6813);
nor U9788 (N_9788,N_6378,N_6554);
nand U9789 (N_9789,N_6426,N_5250);
nand U9790 (N_9790,N_6111,N_6062);
nand U9791 (N_9791,N_7014,N_5750);
or U9792 (N_9792,N_5366,N_5123);
and U9793 (N_9793,N_6482,N_5369);
xor U9794 (N_9794,N_6020,N_6970);
or U9795 (N_9795,N_5112,N_7479);
nor U9796 (N_9796,N_7008,N_6603);
nor U9797 (N_9797,N_5802,N_5955);
xor U9798 (N_9798,N_7265,N_7003);
xnor U9799 (N_9799,N_7029,N_6189);
or U9800 (N_9800,N_5449,N_6148);
and U9801 (N_9801,N_7185,N_5376);
xnor U9802 (N_9802,N_5812,N_5071);
nand U9803 (N_9803,N_7196,N_5598);
xor U9804 (N_9804,N_6398,N_7425);
xnor U9805 (N_9805,N_5289,N_5340);
xnor U9806 (N_9806,N_7304,N_6531);
xor U9807 (N_9807,N_7128,N_5387);
xnor U9808 (N_9808,N_5374,N_5603);
or U9809 (N_9809,N_6308,N_5449);
nor U9810 (N_9810,N_5495,N_6425);
xnor U9811 (N_9811,N_5939,N_5807);
or U9812 (N_9812,N_7493,N_5066);
and U9813 (N_9813,N_5620,N_5395);
or U9814 (N_9814,N_5380,N_5468);
or U9815 (N_9815,N_5916,N_7011);
and U9816 (N_9816,N_5414,N_6857);
nor U9817 (N_9817,N_6055,N_6053);
nor U9818 (N_9818,N_5558,N_6558);
nor U9819 (N_9819,N_5262,N_6158);
xnor U9820 (N_9820,N_6729,N_5457);
xnor U9821 (N_9821,N_6535,N_5855);
xnor U9822 (N_9822,N_5690,N_6116);
nor U9823 (N_9823,N_6588,N_7219);
or U9824 (N_9824,N_6209,N_5585);
nor U9825 (N_9825,N_5523,N_5577);
nand U9826 (N_9826,N_5296,N_6982);
nor U9827 (N_9827,N_5683,N_5412);
and U9828 (N_9828,N_5764,N_6754);
xor U9829 (N_9829,N_6562,N_5074);
nor U9830 (N_9830,N_5811,N_6011);
or U9831 (N_9831,N_5587,N_6088);
or U9832 (N_9832,N_7321,N_5436);
and U9833 (N_9833,N_5940,N_5290);
xor U9834 (N_9834,N_6088,N_7244);
and U9835 (N_9835,N_5972,N_6199);
nand U9836 (N_9836,N_5977,N_6751);
nor U9837 (N_9837,N_7478,N_5527);
nand U9838 (N_9838,N_7400,N_6372);
nor U9839 (N_9839,N_7108,N_6744);
xor U9840 (N_9840,N_7420,N_5528);
and U9841 (N_9841,N_6293,N_5448);
nand U9842 (N_9842,N_5775,N_7236);
or U9843 (N_9843,N_7416,N_7056);
or U9844 (N_9844,N_6986,N_5706);
nand U9845 (N_9845,N_5855,N_6224);
nand U9846 (N_9846,N_7038,N_6486);
and U9847 (N_9847,N_5928,N_6547);
nand U9848 (N_9848,N_7331,N_5578);
xor U9849 (N_9849,N_5700,N_5628);
nor U9850 (N_9850,N_6070,N_6479);
and U9851 (N_9851,N_6954,N_7249);
nor U9852 (N_9852,N_6470,N_5731);
xor U9853 (N_9853,N_6820,N_7202);
or U9854 (N_9854,N_5502,N_6679);
xnor U9855 (N_9855,N_5238,N_6126);
or U9856 (N_9856,N_5548,N_5683);
nand U9857 (N_9857,N_5645,N_6128);
nor U9858 (N_9858,N_6166,N_7354);
and U9859 (N_9859,N_7335,N_5172);
nand U9860 (N_9860,N_6119,N_5461);
xor U9861 (N_9861,N_6026,N_5070);
nor U9862 (N_9862,N_5432,N_6422);
nor U9863 (N_9863,N_5742,N_5105);
or U9864 (N_9864,N_5971,N_7274);
and U9865 (N_9865,N_6106,N_5380);
xnor U9866 (N_9866,N_6764,N_7283);
xnor U9867 (N_9867,N_7170,N_5494);
nor U9868 (N_9868,N_7180,N_5402);
xnor U9869 (N_9869,N_5468,N_5751);
nand U9870 (N_9870,N_5705,N_6303);
or U9871 (N_9871,N_5017,N_6871);
nand U9872 (N_9872,N_7381,N_6503);
and U9873 (N_9873,N_6444,N_6355);
and U9874 (N_9874,N_5014,N_5279);
and U9875 (N_9875,N_7434,N_5545);
or U9876 (N_9876,N_6328,N_7383);
and U9877 (N_9877,N_5308,N_7322);
or U9878 (N_9878,N_5439,N_6337);
or U9879 (N_9879,N_5054,N_7357);
nor U9880 (N_9880,N_6227,N_5295);
xor U9881 (N_9881,N_6463,N_7017);
xor U9882 (N_9882,N_5790,N_5216);
xnor U9883 (N_9883,N_6967,N_6491);
nor U9884 (N_9884,N_6170,N_6062);
nand U9885 (N_9885,N_6438,N_6563);
and U9886 (N_9886,N_6327,N_6411);
nor U9887 (N_9887,N_5878,N_5212);
nor U9888 (N_9888,N_5397,N_5618);
nand U9889 (N_9889,N_5966,N_6092);
nor U9890 (N_9890,N_6494,N_5489);
or U9891 (N_9891,N_6951,N_5132);
nand U9892 (N_9892,N_5127,N_5432);
nand U9893 (N_9893,N_7086,N_5037);
and U9894 (N_9894,N_5293,N_5154);
nor U9895 (N_9895,N_6093,N_7259);
and U9896 (N_9896,N_7296,N_5131);
xor U9897 (N_9897,N_6928,N_6483);
xnor U9898 (N_9898,N_6063,N_7324);
nor U9899 (N_9899,N_6943,N_6865);
and U9900 (N_9900,N_5146,N_5710);
and U9901 (N_9901,N_6951,N_5373);
nor U9902 (N_9902,N_5650,N_5357);
or U9903 (N_9903,N_6027,N_5886);
nor U9904 (N_9904,N_6866,N_6252);
xnor U9905 (N_9905,N_5587,N_5774);
xnor U9906 (N_9906,N_6770,N_6179);
or U9907 (N_9907,N_5948,N_7092);
and U9908 (N_9908,N_7231,N_5061);
nor U9909 (N_9909,N_6409,N_6701);
or U9910 (N_9910,N_7253,N_6623);
and U9911 (N_9911,N_7251,N_6034);
nor U9912 (N_9912,N_7108,N_7145);
or U9913 (N_9913,N_7467,N_5641);
and U9914 (N_9914,N_5241,N_7062);
nand U9915 (N_9915,N_6151,N_5815);
or U9916 (N_9916,N_5975,N_6787);
nand U9917 (N_9917,N_7117,N_6881);
and U9918 (N_9918,N_5948,N_6157);
xor U9919 (N_9919,N_6860,N_5912);
nor U9920 (N_9920,N_5955,N_6010);
nand U9921 (N_9921,N_5991,N_7169);
nor U9922 (N_9922,N_6703,N_5492);
or U9923 (N_9923,N_7478,N_6690);
xnor U9924 (N_9924,N_6069,N_6566);
nand U9925 (N_9925,N_5191,N_7251);
and U9926 (N_9926,N_6939,N_5757);
and U9927 (N_9927,N_6866,N_6538);
nor U9928 (N_9928,N_6145,N_6139);
and U9929 (N_9929,N_6922,N_6121);
or U9930 (N_9930,N_5554,N_6828);
nand U9931 (N_9931,N_5746,N_5790);
xnor U9932 (N_9932,N_6921,N_5986);
or U9933 (N_9933,N_5235,N_5226);
nor U9934 (N_9934,N_7118,N_6955);
nand U9935 (N_9935,N_6523,N_7165);
nor U9936 (N_9936,N_5266,N_5130);
nand U9937 (N_9937,N_5239,N_6722);
xnor U9938 (N_9938,N_7334,N_5297);
or U9939 (N_9939,N_5064,N_7234);
nor U9940 (N_9940,N_5191,N_6300);
and U9941 (N_9941,N_7298,N_6613);
xor U9942 (N_9942,N_6310,N_7210);
xnor U9943 (N_9943,N_5336,N_5174);
or U9944 (N_9944,N_5705,N_5147);
nor U9945 (N_9945,N_6239,N_7407);
nand U9946 (N_9946,N_5221,N_6048);
or U9947 (N_9947,N_5180,N_7003);
nor U9948 (N_9948,N_5474,N_6863);
xor U9949 (N_9949,N_5914,N_5142);
or U9950 (N_9950,N_5532,N_5286);
nor U9951 (N_9951,N_6629,N_6211);
nor U9952 (N_9952,N_6685,N_7290);
xnor U9953 (N_9953,N_6889,N_5400);
and U9954 (N_9954,N_5521,N_5537);
or U9955 (N_9955,N_5085,N_7338);
nor U9956 (N_9956,N_6404,N_6400);
xor U9957 (N_9957,N_6688,N_5181);
xor U9958 (N_9958,N_6543,N_6240);
nand U9959 (N_9959,N_7408,N_7222);
and U9960 (N_9960,N_5158,N_5930);
or U9961 (N_9961,N_5392,N_5813);
xnor U9962 (N_9962,N_5024,N_5716);
nor U9963 (N_9963,N_7233,N_7485);
xnor U9964 (N_9964,N_7117,N_5458);
nand U9965 (N_9965,N_5425,N_7213);
nor U9966 (N_9966,N_6660,N_5016);
or U9967 (N_9967,N_7231,N_5619);
and U9968 (N_9968,N_5997,N_6166);
xnor U9969 (N_9969,N_6824,N_6518);
xnor U9970 (N_9970,N_6305,N_6023);
and U9971 (N_9971,N_7282,N_6123);
xnor U9972 (N_9972,N_7499,N_6210);
and U9973 (N_9973,N_5795,N_6736);
nand U9974 (N_9974,N_6375,N_5116);
nand U9975 (N_9975,N_5384,N_6216);
nand U9976 (N_9976,N_5994,N_5862);
nor U9977 (N_9977,N_6346,N_5933);
xnor U9978 (N_9978,N_6313,N_6683);
nand U9979 (N_9979,N_7456,N_6875);
nand U9980 (N_9980,N_7401,N_6986);
and U9981 (N_9981,N_7157,N_5843);
or U9982 (N_9982,N_5712,N_5605);
nor U9983 (N_9983,N_5250,N_5969);
nand U9984 (N_9984,N_6562,N_6601);
or U9985 (N_9985,N_5735,N_7067);
and U9986 (N_9986,N_6629,N_7463);
nor U9987 (N_9987,N_6472,N_6747);
xor U9988 (N_9988,N_6373,N_5968);
nand U9989 (N_9989,N_6101,N_5385);
nand U9990 (N_9990,N_5193,N_6606);
nand U9991 (N_9991,N_6301,N_5144);
and U9992 (N_9992,N_5319,N_7191);
nor U9993 (N_9993,N_7372,N_6958);
nor U9994 (N_9994,N_7341,N_6830);
or U9995 (N_9995,N_7066,N_7107);
xnor U9996 (N_9996,N_7361,N_7461);
and U9997 (N_9997,N_6566,N_6863);
xnor U9998 (N_9998,N_6307,N_6009);
nand U9999 (N_9999,N_6687,N_6163);
nor UO_0 (O_0,N_8815,N_8414);
and UO_1 (O_1,N_7852,N_9064);
nor UO_2 (O_2,N_9210,N_7579);
or UO_3 (O_3,N_8500,N_9509);
xor UO_4 (O_4,N_9183,N_8595);
nor UO_5 (O_5,N_8631,N_9944);
xor UO_6 (O_6,N_9535,N_9129);
xnor UO_7 (O_7,N_8741,N_9729);
nand UO_8 (O_8,N_9585,N_8635);
xnor UO_9 (O_9,N_7509,N_8093);
xor UO_10 (O_10,N_8400,N_8603);
nor UO_11 (O_11,N_9415,N_9085);
and UO_12 (O_12,N_9516,N_9340);
nand UO_13 (O_13,N_9855,N_7636);
nand UO_14 (O_14,N_8764,N_7573);
nor UO_15 (O_15,N_8811,N_9756);
xnor UO_16 (O_16,N_7850,N_8489);
or UO_17 (O_17,N_8460,N_8597);
nand UO_18 (O_18,N_8553,N_8096);
nand UO_19 (O_19,N_9547,N_9333);
nand UO_20 (O_20,N_8024,N_9815);
or UO_21 (O_21,N_9053,N_9996);
or UO_22 (O_22,N_9031,N_9993);
or UO_23 (O_23,N_9706,N_9599);
or UO_24 (O_24,N_7841,N_9147);
nand UO_25 (O_25,N_9660,N_9778);
nor UO_26 (O_26,N_8275,N_9066);
or UO_27 (O_27,N_8733,N_7688);
xor UO_28 (O_28,N_7857,N_7723);
nor UO_29 (O_29,N_8454,N_8744);
nor UO_30 (O_30,N_9707,N_9310);
and UO_31 (O_31,N_7574,N_9046);
or UO_32 (O_32,N_7724,N_8940);
nor UO_33 (O_33,N_9838,N_7618);
or UO_34 (O_34,N_8245,N_8911);
nand UO_35 (O_35,N_8194,N_8680);
nand UO_36 (O_36,N_9363,N_8347);
and UO_37 (O_37,N_9238,N_9135);
or UO_38 (O_38,N_9105,N_8295);
or UO_39 (O_39,N_7631,N_8143);
xnor UO_40 (O_40,N_8497,N_8386);
nand UO_41 (O_41,N_9079,N_7848);
and UO_42 (O_42,N_9819,N_8466);
nand UO_43 (O_43,N_7878,N_7621);
nand UO_44 (O_44,N_8541,N_9564);
nor UO_45 (O_45,N_9545,N_9762);
and UO_46 (O_46,N_8622,N_8159);
and UO_47 (O_47,N_8828,N_8762);
nor UO_48 (O_48,N_8936,N_8486);
or UO_49 (O_49,N_8151,N_8901);
nand UO_50 (O_50,N_9661,N_8258);
nand UO_51 (O_51,N_8506,N_7785);
nor UO_52 (O_52,N_9335,N_8441);
or UO_53 (O_53,N_7668,N_8459);
and UO_54 (O_54,N_9752,N_8915);
nand UO_55 (O_55,N_7641,N_8077);
and UO_56 (O_56,N_9686,N_7746);
or UO_57 (O_57,N_9475,N_8920);
and UO_58 (O_58,N_9833,N_8327);
xor UO_59 (O_59,N_9791,N_7715);
xnor UO_60 (O_60,N_7976,N_8246);
xnor UO_61 (O_61,N_9241,N_7823);
xnor UO_62 (O_62,N_7686,N_9020);
xnor UO_63 (O_63,N_9169,N_9469);
nor UO_64 (O_64,N_9750,N_7750);
or UO_65 (O_65,N_7781,N_8705);
nand UO_66 (O_66,N_9731,N_9471);
and UO_67 (O_67,N_8044,N_8191);
nand UO_68 (O_68,N_9655,N_8370);
nand UO_69 (O_69,N_9744,N_7953);
nand UO_70 (O_70,N_8239,N_8367);
or UO_71 (O_71,N_8904,N_9269);
and UO_72 (O_72,N_9417,N_9149);
xnor UO_73 (O_73,N_9159,N_9100);
xnor UO_74 (O_74,N_9161,N_9919);
xnor UO_75 (O_75,N_7828,N_9579);
or UO_76 (O_76,N_7513,N_8638);
nand UO_77 (O_77,N_8129,N_8543);
and UO_78 (O_78,N_8814,N_8594);
xor UO_79 (O_79,N_9111,N_9747);
nand UO_80 (O_80,N_9146,N_8994);
nor UO_81 (O_81,N_7890,N_9621);
xnor UO_82 (O_82,N_8606,N_7766);
xnor UO_83 (O_83,N_8127,N_9866);
or UO_84 (O_84,N_7662,N_9235);
or UO_85 (O_85,N_7928,N_9894);
xor UO_86 (O_86,N_7695,N_9005);
xor UO_87 (O_87,N_9843,N_9376);
nor UO_88 (O_88,N_8887,N_7967);
xor UO_89 (O_89,N_7542,N_9027);
and UO_90 (O_90,N_9945,N_9581);
and UO_91 (O_91,N_9905,N_9828);
and UO_92 (O_92,N_8062,N_9913);
or UO_93 (O_93,N_9711,N_7786);
nand UO_94 (O_94,N_9739,N_8822);
or UO_95 (O_95,N_9302,N_9280);
and UO_96 (O_96,N_8910,N_8254);
xor UO_97 (O_97,N_9757,N_8425);
and UO_98 (O_98,N_9764,N_9180);
and UO_99 (O_99,N_7560,N_8927);
or UO_100 (O_100,N_9804,N_7589);
xnor UO_101 (O_101,N_9718,N_9935);
and UO_102 (O_102,N_7888,N_7827);
or UO_103 (O_103,N_8291,N_8107);
nand UO_104 (O_104,N_9278,N_7569);
xor UO_105 (O_105,N_8823,N_9613);
and UO_106 (O_106,N_8690,N_8616);
xnor UO_107 (O_107,N_8673,N_9330);
nor UO_108 (O_108,N_8854,N_9240);
nor UO_109 (O_109,N_7563,N_8114);
nand UO_110 (O_110,N_8008,N_9970);
and UO_111 (O_111,N_9219,N_7821);
nor UO_112 (O_112,N_7664,N_9862);
and UO_113 (O_113,N_9308,N_8753);
nor UO_114 (O_114,N_9504,N_9200);
nor UO_115 (O_115,N_8394,N_8119);
xnor UO_116 (O_116,N_9156,N_9732);
xor UO_117 (O_117,N_7859,N_7792);
and UO_118 (O_118,N_9533,N_8001);
and UO_119 (O_119,N_9758,N_8505);
and UO_120 (O_120,N_9976,N_8440);
nand UO_121 (O_121,N_7815,N_8260);
nor UO_122 (O_122,N_8080,N_7773);
or UO_123 (O_123,N_8780,N_9868);
and UO_124 (O_124,N_7814,N_9923);
and UO_125 (O_125,N_8329,N_8659);
xor UO_126 (O_126,N_8368,N_9624);
nor UO_127 (O_127,N_8446,N_9709);
nor UO_128 (O_128,N_8951,N_9125);
or UO_129 (O_129,N_8178,N_8433);
or UO_130 (O_130,N_9746,N_8689);
and UO_131 (O_131,N_8643,N_9749);
and UO_132 (O_132,N_8054,N_9687);
nand UO_133 (O_133,N_8304,N_7844);
xnor UO_134 (O_134,N_8161,N_9072);
nand UO_135 (O_135,N_7936,N_8049);
nor UO_136 (O_136,N_9481,N_9258);
xor UO_137 (O_137,N_9262,N_8771);
xor UO_138 (O_138,N_8075,N_8973);
nand UO_139 (O_139,N_8878,N_9304);
and UO_140 (O_140,N_8538,N_7514);
xor UO_141 (O_141,N_7570,N_9421);
nor UO_142 (O_142,N_9846,N_9849);
and UO_143 (O_143,N_9629,N_7860);
and UO_144 (O_144,N_9979,N_8526);
nand UO_145 (O_145,N_9666,N_8092);
and UO_146 (O_146,N_9370,N_8132);
and UO_147 (O_147,N_8840,N_7948);
and UO_148 (O_148,N_8421,N_7501);
and UO_149 (O_149,N_7701,N_8410);
or UO_150 (O_150,N_9225,N_9755);
xnor UO_151 (O_151,N_8311,N_9852);
xor UO_152 (O_152,N_8736,N_9999);
and UO_153 (O_153,N_7637,N_7632);
nand UO_154 (O_154,N_7939,N_7580);
nand UO_155 (O_155,N_7903,N_9783);
xor UO_156 (O_156,N_9268,N_7721);
or UO_157 (O_157,N_7753,N_8221);
or UO_158 (O_158,N_8135,N_8913);
or UO_159 (O_159,N_8584,N_9179);
xnor UO_160 (O_160,N_7764,N_8747);
xnor UO_161 (O_161,N_8626,N_9879);
xnor UO_162 (O_162,N_7806,N_9039);
nand UO_163 (O_163,N_8919,N_7608);
xor UO_164 (O_164,N_9283,N_9000);
nor UO_165 (O_165,N_9356,N_9048);
or UO_166 (O_166,N_7969,N_8533);
nand UO_167 (O_167,N_8222,N_8248);
and UO_168 (O_168,N_9910,N_9338);
nor UO_169 (O_169,N_9980,N_9860);
or UO_170 (O_170,N_9355,N_9953);
nor UO_171 (O_171,N_8396,N_9554);
xnor UO_172 (O_172,N_9679,N_9320);
or UO_173 (O_173,N_9371,N_8265);
nand UO_174 (O_174,N_9394,N_9780);
nor UO_175 (O_175,N_8312,N_9524);
and UO_176 (O_176,N_9300,N_8059);
nand UO_177 (O_177,N_9658,N_9657);
xnor UO_178 (O_178,N_8856,N_8413);
xnor UO_179 (O_179,N_8398,N_9315);
nand UO_180 (O_180,N_8802,N_8409);
xnor UO_181 (O_181,N_8227,N_8319);
or UO_182 (O_182,N_8022,N_8478);
or UO_183 (O_183,N_8542,N_8165);
nor UO_184 (O_184,N_7812,N_8580);
or UO_185 (O_185,N_8534,N_9276);
xnor UO_186 (O_186,N_7898,N_8152);
and UO_187 (O_187,N_8464,N_9196);
or UO_188 (O_188,N_8945,N_7527);
or UO_189 (O_189,N_8145,N_9576);
nor UO_190 (O_190,N_9137,N_8401);
or UO_191 (O_191,N_7795,N_9632);
nor UO_192 (O_192,N_9802,N_9830);
xnor UO_193 (O_193,N_9119,N_7867);
nand UO_194 (O_194,N_8448,N_8859);
or UO_195 (O_195,N_8423,N_9068);
and UO_196 (O_196,N_9503,N_7972);
xnor UO_197 (O_197,N_9045,N_9487);
xor UO_198 (O_198,N_8081,N_9432);
xnor UO_199 (O_199,N_8742,N_9735);
and UO_200 (O_200,N_8346,N_9202);
xnor UO_201 (O_201,N_7762,N_7713);
nor UO_202 (O_202,N_7789,N_8349);
and UO_203 (O_203,N_7627,N_8789);
nor UO_204 (O_204,N_8213,N_9412);
and UO_205 (O_205,N_9143,N_9033);
nand UO_206 (O_206,N_8471,N_8038);
and UO_207 (O_207,N_8184,N_9737);
or UO_208 (O_208,N_7562,N_9633);
or UO_209 (O_209,N_8284,N_7597);
or UO_210 (O_210,N_8966,N_9592);
or UO_211 (O_211,N_7524,N_9152);
nor UO_212 (O_212,N_7633,N_9406);
and UO_213 (O_213,N_7986,N_9987);
nor UO_214 (O_214,N_9456,N_7919);
nor UO_215 (O_215,N_7659,N_8271);
or UO_216 (O_216,N_9274,N_8773);
nand UO_217 (O_217,N_7653,N_8750);
nor UO_218 (O_218,N_9150,N_9069);
nor UO_219 (O_219,N_9028,N_9299);
xnor UO_220 (O_220,N_7772,N_9844);
or UO_221 (O_221,N_9257,N_8849);
and UO_222 (O_222,N_9230,N_8261);
and UO_223 (O_223,N_8361,N_8405);
nor UO_224 (O_224,N_9035,N_9604);
nand UO_225 (O_225,N_7949,N_8267);
xor UO_226 (O_226,N_8693,N_8691);
xor UO_227 (O_227,N_8279,N_8617);
nand UO_228 (O_228,N_9422,N_9001);
nand UO_229 (O_229,N_9559,N_8600);
nor UO_230 (O_230,N_8906,N_9622);
xor UO_231 (O_231,N_8810,N_8094);
nor UO_232 (O_232,N_8028,N_9431);
or UO_233 (O_233,N_9378,N_7736);
nand UO_234 (O_234,N_9223,N_9337);
or UO_235 (O_235,N_7630,N_9386);
or UO_236 (O_236,N_9113,N_7797);
and UO_237 (O_237,N_8109,N_8696);
and UO_238 (O_238,N_7571,N_8030);
or UO_239 (O_239,N_8984,N_8676);
nand UO_240 (O_240,N_8937,N_8422);
xnor UO_241 (O_241,N_9895,N_8982);
nor UO_242 (O_242,N_9864,N_9556);
and UO_243 (O_243,N_8513,N_9982);
nor UO_244 (O_244,N_8457,N_9584);
and UO_245 (O_245,N_8527,N_8941);
and UO_246 (O_246,N_9008,N_8384);
xor UO_247 (O_247,N_9091,N_9204);
xor UO_248 (O_248,N_8628,N_9022);
and UO_249 (O_249,N_9742,N_8939);
or UO_250 (O_250,N_9051,N_8494);
and UO_251 (O_251,N_9591,N_7914);
and UO_252 (O_252,N_9336,N_9936);
nor UO_253 (O_253,N_9126,N_8954);
and UO_254 (O_254,N_9322,N_9187);
nand UO_255 (O_255,N_8025,N_8155);
nand UO_256 (O_256,N_7520,N_9733);
nor UO_257 (O_257,N_9414,N_7535);
nor UO_258 (O_258,N_8399,N_9975);
or UO_259 (O_259,N_7930,N_9662);
nand UO_260 (O_260,N_7744,N_9642);
or UO_261 (O_261,N_9647,N_7853);
and UO_262 (O_262,N_8266,N_8359);
nor UO_263 (O_263,N_9796,N_8962);
nor UO_264 (O_264,N_9586,N_7554);
nand UO_265 (O_265,N_8636,N_8540);
or UO_266 (O_266,N_9527,N_8447);
or UO_267 (O_267,N_9854,N_9245);
nand UO_268 (O_268,N_9728,N_8051);
or UO_269 (O_269,N_8066,N_7741);
nor UO_270 (O_270,N_9295,N_9443);
or UO_271 (O_271,N_8324,N_9608);
nand UO_272 (O_272,N_7768,N_9676);
or UO_273 (O_273,N_8979,N_8259);
and UO_274 (O_274,N_7564,N_7959);
and UO_275 (O_275,N_9789,N_9198);
xnor UO_276 (O_276,N_8047,N_8065);
or UO_277 (O_277,N_8196,N_8436);
and UO_278 (O_278,N_9148,N_9779);
nand UO_279 (O_279,N_9437,N_8826);
xor UO_280 (O_280,N_7583,N_9943);
or UO_281 (O_281,N_9270,N_7816);
nor UO_282 (O_282,N_7505,N_8894);
and UO_283 (O_283,N_9346,N_9157);
nor UO_284 (O_284,N_9771,N_8099);
or UO_285 (O_285,N_9721,N_8640);
and UO_286 (O_286,N_9428,N_9674);
nand UO_287 (O_287,N_8662,N_8943);
and UO_288 (O_288,N_9244,N_9929);
xor UO_289 (O_289,N_8511,N_7916);
nand UO_290 (O_290,N_9070,N_8088);
xor UO_291 (O_291,N_7738,N_8432);
nand UO_292 (O_292,N_9402,N_7984);
or UO_293 (O_293,N_9181,N_9812);
nand UO_294 (O_294,N_8768,N_8864);
nor UO_295 (O_295,N_8176,N_7887);
nor UO_296 (O_296,N_9102,N_7722);
xor UO_297 (O_297,N_7669,N_7690);
nor UO_298 (O_298,N_8276,N_9857);
and UO_299 (O_299,N_9347,N_9582);
nand UO_300 (O_300,N_7800,N_8665);
or UO_301 (O_301,N_9413,N_8668);
nor UO_302 (O_302,N_9447,N_9824);
xor UO_303 (O_303,N_7547,N_7731);
nand UO_304 (O_304,N_9882,N_8530);
nand UO_305 (O_305,N_8407,N_7693);
xor UO_306 (O_306,N_8234,N_8344);
nand UO_307 (O_307,N_9185,N_9600);
or UO_308 (O_308,N_7550,N_8375);
and UO_309 (O_309,N_8743,N_9160);
xnor UO_310 (O_310,N_7622,N_8362);
nand UO_311 (O_311,N_8732,N_8599);
nand UO_312 (O_312,N_9172,N_7747);
or UO_313 (O_313,N_9388,N_8095);
and UO_314 (O_314,N_7896,N_7709);
nand UO_315 (O_315,N_8063,N_9967);
xnor UO_316 (O_316,N_8701,N_9365);
nand UO_317 (O_317,N_8649,N_8969);
or UO_318 (O_318,N_8769,N_7791);
and UO_319 (O_319,N_7796,N_8148);
and UO_320 (O_320,N_8577,N_9792);
nand UO_321 (O_321,N_8201,N_9389);
nand UO_322 (O_322,N_9252,N_7658);
nor UO_323 (O_323,N_7805,N_9653);
nand UO_324 (O_324,N_9457,N_8663);
or UO_325 (O_325,N_9671,N_7742);
and UO_326 (O_326,N_7774,N_8443);
xnor UO_327 (O_327,N_7672,N_9877);
xor UO_328 (O_328,N_7963,N_7757);
nand UO_329 (O_329,N_8847,N_8342);
and UO_330 (O_330,N_9738,N_9464);
xnor UO_331 (O_331,N_8761,N_9578);
nor UO_332 (O_332,N_8935,N_7975);
and UO_333 (O_333,N_7956,N_9442);
nor UO_334 (O_334,N_9800,N_7523);
or UO_335 (O_335,N_8113,N_8593);
xor UO_336 (O_336,N_9941,N_9536);
and UO_337 (O_337,N_7683,N_8090);
nor UO_338 (O_338,N_8153,N_9817);
xor UO_339 (O_339,N_9221,N_9859);
xnor UO_340 (O_340,N_9641,N_7754);
nand UO_341 (O_341,N_9587,N_9191);
or UO_342 (O_342,N_9141,N_8130);
nand UO_343 (O_343,N_7990,N_8158);
nor UO_344 (O_344,N_8235,N_8108);
or UO_345 (O_345,N_8351,N_8071);
nor UO_346 (O_346,N_9133,N_8830);
nor UO_347 (O_347,N_8551,N_7537);
or UO_348 (O_348,N_8816,N_7617);
xnor UO_349 (O_349,N_7946,N_9360);
or UO_350 (O_350,N_8253,N_8115);
nand UO_351 (O_351,N_8598,N_9358);
nand UO_352 (O_352,N_7784,N_7932);
nor UO_353 (O_353,N_8147,N_9960);
nor UO_354 (O_354,N_8412,N_8805);
xor UO_355 (O_355,N_7638,N_9942);
or UO_356 (O_356,N_8179,N_7615);
or UO_357 (O_357,N_8681,N_8523);
or UO_358 (O_358,N_8417,N_8765);
and UO_359 (O_359,N_8559,N_9924);
xnor UO_360 (O_360,N_8790,N_9741);
xor UO_361 (O_361,N_9690,N_9215);
and UO_362 (O_362,N_9520,N_9659);
or UO_363 (O_363,N_8870,N_9768);
or UO_364 (O_364,N_9399,N_8204);
xnor UO_365 (O_365,N_9806,N_8924);
nor UO_366 (O_366,N_9004,N_9572);
and UO_367 (O_367,N_8007,N_8150);
nand UO_368 (O_368,N_9153,N_8565);
nand UO_369 (O_369,N_9018,N_8990);
nand UO_370 (O_370,N_7977,N_8575);
xor UO_371 (O_371,N_9213,N_8453);
xor UO_372 (O_372,N_8382,N_9781);
nand UO_373 (O_373,N_9809,N_9023);
or UO_374 (O_374,N_9610,N_7954);
nor UO_375 (O_375,N_7904,N_9243);
xnor UO_376 (O_376,N_7943,N_8579);
and UO_377 (O_377,N_8468,N_8069);
nand UO_378 (O_378,N_9491,N_8480);
or UO_379 (O_379,N_9981,N_8999);
nand UO_380 (O_380,N_9209,N_8252);
xor UO_381 (O_381,N_9871,N_9829);
or UO_382 (O_382,N_8653,N_9896);
and UO_383 (O_383,N_8907,N_7807);
nor UO_384 (O_384,N_8385,N_8091);
nand UO_385 (O_385,N_9727,N_7679);
and UO_386 (O_386,N_8331,N_8012);
or UO_387 (O_387,N_9101,N_7720);
nand UO_388 (O_388,N_8499,N_9284);
and UO_389 (O_389,N_7831,N_9229);
nor UO_390 (O_390,N_9205,N_8820);
nand UO_391 (O_391,N_8376,N_8861);
xor UO_392 (O_392,N_9593,N_9379);
xnor UO_393 (O_393,N_9061,N_9760);
nor UO_394 (O_394,N_9753,N_9555);
or UO_395 (O_395,N_9530,N_9436);
nand UO_396 (O_396,N_8685,N_9248);
nand UO_397 (O_397,N_7871,N_8144);
nand UO_398 (O_398,N_8726,N_7941);
nand UO_399 (O_399,N_8525,N_8948);
xnor UO_400 (O_400,N_8782,N_8137);
xnor UO_401 (O_401,N_7538,N_8492);
xnor UO_402 (O_402,N_8290,N_8989);
nor UO_403 (O_403,N_9962,N_7988);
nand UO_404 (O_404,N_7906,N_9416);
and UO_405 (O_405,N_9407,N_8219);
or UO_406 (O_406,N_8909,N_9260);
xor UO_407 (O_407,N_7870,N_9523);
xnor UO_408 (O_408,N_9502,N_9907);
and UO_409 (O_409,N_9251,N_9228);
or UO_410 (O_410,N_9314,N_9607);
or UO_411 (O_411,N_8032,N_9540);
nand UO_412 (O_412,N_9271,N_7801);
nor UO_413 (O_413,N_9439,N_9013);
xnor UO_414 (O_414,N_9345,N_8629);
nor UO_415 (O_415,N_9513,N_7897);
and UO_416 (O_416,N_9548,N_9664);
xnor UO_417 (O_417,N_7869,N_8833);
xnor UO_418 (O_418,N_9900,N_8437);
nor UO_419 (O_419,N_9353,N_9420);
and UO_420 (O_420,N_9788,N_9254);
nor UO_421 (O_421,N_8763,N_8287);
nor UO_422 (O_422,N_7872,N_7868);
xor UO_423 (O_423,N_9165,N_8532);
nand UO_424 (O_424,N_8023,N_7955);
or UO_425 (O_425,N_8884,N_8719);
and UO_426 (O_426,N_8652,N_9626);
nand UO_427 (O_427,N_7861,N_8714);
nor UO_428 (O_428,N_7541,N_9850);
and UO_429 (O_429,N_8498,N_7737);
nand UO_430 (O_430,N_8841,N_8985);
xor UO_431 (O_431,N_8043,N_8852);
xnor UO_432 (O_432,N_9144,N_7830);
nand UO_433 (O_433,N_7656,N_8517);
nand UO_434 (O_434,N_7855,N_9192);
nand UO_435 (O_435,N_9708,N_8465);
and UO_436 (O_436,N_9208,N_9403);
xnor UO_437 (O_437,N_8000,N_9317);
and UO_438 (O_438,N_7603,N_8713);
and UO_439 (O_439,N_7749,N_7759);
nor UO_440 (O_440,N_8503,N_9845);
nand UO_441 (O_441,N_9019,N_8122);
xor UO_442 (O_442,N_8341,N_8953);
xor UO_443 (O_443,N_8117,N_9343);
nor UO_444 (O_444,N_9901,N_8717);
nand UO_445 (O_445,N_8903,N_8784);
nor UO_446 (O_446,N_9207,N_7655);
and UO_447 (O_447,N_7593,N_9627);
nor UO_448 (O_448,N_7838,N_8146);
nand UO_449 (O_449,N_8957,N_7769);
or UO_450 (O_450,N_8605,N_9327);
xnor UO_451 (O_451,N_9878,N_7775);
nand UO_452 (O_452,N_8749,N_7676);
nor UO_453 (O_453,N_7767,N_9751);
or UO_454 (O_454,N_7725,N_9383);
nand UO_455 (O_455,N_9296,N_7694);
and UO_456 (O_456,N_8273,N_8257);
or UO_457 (O_457,N_9594,N_8801);
nor UO_458 (O_458,N_9015,N_8174);
and UO_459 (O_459,N_8018,N_9688);
xor UO_460 (O_460,N_7743,N_9853);
and UO_461 (O_461,N_9303,N_8632);
and UO_462 (O_462,N_8930,N_8426);
and UO_463 (O_463,N_8079,N_8991);
nor UO_464 (O_464,N_8374,N_8862);
xnor UO_465 (O_465,N_9381,N_8225);
or UO_466 (O_466,N_7654,N_8186);
and UO_467 (O_467,N_8029,N_8495);
xnor UO_468 (O_468,N_8658,N_8111);
xnor UO_469 (O_469,N_8098,N_8212);
nand UO_470 (O_470,N_8420,N_8809);
and UO_471 (O_471,N_9617,N_9890);
xnor UO_472 (O_472,N_8157,N_7665);
or UO_473 (O_473,N_8670,N_9140);
nor UO_474 (O_474,N_9098,N_9142);
or UO_475 (O_475,N_9211,N_8781);
or UO_476 (O_476,N_7596,N_8633);
or UO_477 (O_477,N_8912,N_9644);
nor UO_478 (O_478,N_9212,N_8574);
xnor UO_479 (O_479,N_8845,N_9518);
or UO_480 (O_480,N_8269,N_9324);
or UO_481 (O_481,N_8928,N_9500);
or UO_482 (O_482,N_8596,N_8562);
or UO_483 (O_483,N_9357,N_8315);
nor UO_484 (O_484,N_8730,N_8348);
and UO_485 (O_485,N_8485,N_8140);
or UO_486 (O_486,N_9026,N_7817);
and UO_487 (O_487,N_9495,N_8639);
nand UO_488 (O_488,N_9589,N_7696);
and UO_489 (O_489,N_8268,N_9774);
and UO_490 (O_490,N_8377,N_8255);
and UO_491 (O_491,N_8981,N_8877);
xnor UO_492 (O_492,N_9206,N_9190);
nor UO_493 (O_493,N_8381,N_7539);
or UO_494 (O_494,N_8893,N_8683);
nor UO_495 (O_495,N_9261,N_9329);
nand UO_496 (O_496,N_8476,N_9730);
xnor UO_497 (O_497,N_8104,N_7921);
or UO_498 (O_498,N_8672,N_8720);
xnor UO_499 (O_499,N_8272,N_9164);
nor UO_500 (O_500,N_8578,N_8898);
xor UO_501 (O_501,N_8218,N_8961);
or UO_502 (O_502,N_9998,N_9775);
xor UO_503 (O_503,N_8918,N_9695);
nand UO_504 (O_504,N_8293,N_7782);
or UO_505 (O_505,N_8777,N_8739);
and UO_506 (O_506,N_9832,N_7549);
nand UO_507 (O_507,N_8914,N_9231);
nand UO_508 (O_508,N_7697,N_7646);
nor UO_509 (O_509,N_7612,N_7504);
and UO_510 (O_510,N_9972,N_8886);
or UO_511 (O_511,N_9726,N_8800);
nor UO_512 (O_512,N_9798,N_8334);
or UO_513 (O_513,N_9888,N_8380);
or UO_514 (O_514,N_9770,N_8702);
nor UO_515 (O_515,N_9927,N_9865);
and UO_516 (O_516,N_9567,N_9095);
nor UO_517 (O_517,N_8923,N_8164);
nand UO_518 (O_518,N_7556,N_9650);
and UO_519 (O_519,N_9049,N_8408);
xor UO_520 (O_520,N_8428,N_9339);
or UO_521 (O_521,N_9784,N_9876);
xor UO_522 (O_522,N_8281,N_7595);
and UO_523 (O_523,N_9193,N_9598);
and UO_524 (O_524,N_9037,N_8475);
nor UO_525 (O_525,N_9349,N_8189);
nor UO_526 (O_526,N_9233,N_9813);
xnor UO_527 (O_527,N_9321,N_7856);
nand UO_528 (O_528,N_8306,N_8057);
nand UO_529 (O_529,N_7847,N_8558);
and UO_530 (O_530,N_7752,N_7891);
xor UO_531 (O_531,N_9423,N_9628);
nand UO_532 (O_532,N_7704,N_9404);
xor UO_533 (O_533,N_9831,N_8325);
xnor UO_534 (O_534,N_9342,N_8872);
and UO_535 (O_535,N_9766,N_9656);
and UO_536 (O_536,N_8775,N_8838);
or UO_537 (O_537,N_7783,N_8804);
nor UO_538 (O_538,N_8048,N_7918);
or UO_539 (O_539,N_8889,N_9427);
nor UO_540 (O_540,N_9908,N_9638);
and UO_541 (O_541,N_8902,N_9021);
nand UO_542 (O_542,N_8456,N_9918);
or UO_543 (O_543,N_7522,N_7577);
nand UO_544 (O_544,N_9915,N_7698);
and UO_545 (O_545,N_9724,N_8895);
nor UO_546 (O_546,N_8364,N_8006);
and UO_547 (O_547,N_7794,N_9801);
nand UO_548 (O_548,N_8230,N_7707);
nor UO_549 (O_549,N_8602,N_8586);
nor UO_550 (O_550,N_9625,N_8017);
xnor UO_551 (O_551,N_9562,N_7517);
nand UO_552 (O_552,N_9712,N_8014);
and UO_553 (O_553,N_9006,N_9186);
or UO_554 (O_554,N_8835,N_9848);
or UO_555 (O_555,N_8869,N_8524);
and UO_556 (O_556,N_7712,N_8993);
nand UO_557 (O_557,N_7982,N_8074);
nand UO_558 (O_558,N_8045,N_8850);
nor UO_559 (O_559,N_9958,N_8671);
xor UO_560 (O_560,N_9362,N_8788);
nor UO_561 (O_561,N_9418,N_9574);
and UO_562 (O_562,N_9065,N_9350);
xor UO_563 (O_563,N_8876,N_8926);
nor UO_564 (O_564,N_8350,N_8149);
nand UO_565 (O_565,N_8118,N_7915);
xor UO_566 (O_566,N_9790,N_8326);
nand UO_567 (O_567,N_8323,N_8883);
xor UO_568 (O_568,N_9086,N_7661);
nor UO_569 (O_569,N_8974,N_8875);
nand UO_570 (O_570,N_8288,N_8687);
or UO_571 (O_571,N_8226,N_7981);
and UO_572 (O_572,N_9002,N_9694);
xnor UO_573 (O_573,N_8031,N_9869);
xor UO_574 (O_574,N_8187,N_8064);
or UO_575 (O_575,N_8619,N_7687);
nor UO_576 (O_576,N_8621,N_9974);
nor UO_577 (O_577,N_7635,N_9038);
xnor UO_578 (O_578,N_9501,N_7881);
or UO_579 (O_579,N_7719,N_7950);
nand UO_580 (O_580,N_9114,N_8708);
nand UO_581 (O_581,N_7854,N_9275);
or UO_582 (O_582,N_8755,N_9636);
nand UO_583 (O_583,N_7863,N_9009);
or UO_584 (O_584,N_8335,N_9397);
nor UO_585 (O_585,N_9703,N_9445);
nor UO_586 (O_586,N_9400,N_8393);
nor UO_587 (O_587,N_8821,N_9596);
or UO_588 (O_588,N_9606,N_9189);
nor UO_589 (O_589,N_9118,N_8808);
or UO_590 (O_590,N_9203,N_9036);
or UO_591 (O_591,N_9692,N_7989);
or UO_592 (O_592,N_8899,N_8424);
nor UO_593 (O_593,N_9089,N_7515);
nor UO_594 (O_594,N_8866,N_7908);
nor UO_595 (O_595,N_8576,N_8917);
and UO_596 (O_596,N_7645,N_9103);
xor UO_597 (O_597,N_9930,N_9060);
and UO_598 (O_598,N_8116,N_8208);
nand UO_599 (O_599,N_7651,N_8977);
nor UO_600 (O_600,N_9909,N_9474);
xnor UO_601 (O_601,N_8379,N_7923);
nand UO_602 (O_602,N_9216,N_9887);
or UO_603 (O_603,N_9145,N_9047);
xor UO_604 (O_604,N_7952,N_8112);
or UO_605 (O_605,N_9971,N_8390);
xnor UO_606 (O_606,N_8729,N_8836);
and UO_607 (O_607,N_7578,N_8795);
nor UO_608 (O_608,N_7760,N_7947);
nor UO_609 (O_609,N_8103,N_9134);
and UO_610 (O_610,N_9588,N_7985);
and UO_611 (O_611,N_9977,N_8699);
or UO_612 (O_612,N_9226,N_7528);
and UO_613 (O_613,N_9512,N_8863);
or UO_614 (O_614,N_7974,N_7729);
and UO_615 (O_615,N_9099,N_8880);
nand UO_616 (O_616,N_7642,N_8087);
nor UO_617 (O_617,N_7810,N_9289);
xor UO_618 (O_618,N_9517,N_9816);
xor UO_619 (O_619,N_9580,N_9870);
xor UO_620 (O_620,N_8655,N_9597);
nand UO_621 (O_621,N_8190,N_9259);
nor UO_622 (O_622,N_8608,N_8660);
or UO_623 (O_623,N_7788,N_8046);
nand UO_624 (O_624,N_8358,N_8625);
and UO_625 (O_625,N_8537,N_9369);
and UO_626 (O_626,N_7840,N_9384);
nor UO_627 (O_627,N_9348,N_8614);
nor UO_628 (O_628,N_9242,N_7545);
xor UO_629 (O_629,N_8703,N_8039);
nand UO_630 (O_630,N_9990,N_9479);
and UO_631 (O_631,N_8160,N_9106);
and UO_632 (O_632,N_8604,N_9640);
nand UO_633 (O_633,N_9522,N_8223);
xor UO_634 (O_634,N_9305,N_9032);
and UO_635 (O_635,N_7702,N_9331);
nor UO_636 (O_636,N_9799,N_7973);
nor UO_637 (O_637,N_9067,N_8387);
nor UO_638 (O_638,N_9956,N_9620);
and UO_639 (O_639,N_8797,N_8013);
and UO_640 (O_640,N_9218,N_9785);
or UO_641 (O_641,N_7809,N_7811);
nand UO_642 (O_642,N_7971,N_8637);
nand UO_643 (O_643,N_8516,N_8216);
nand UO_644 (O_644,N_9030,N_7978);
nor UO_645 (O_645,N_8561,N_9438);
nor UO_646 (O_646,N_9398,N_7600);
nand UO_647 (O_647,N_9040,N_8648);
and UO_648 (O_648,N_8921,N_9863);
nor UO_649 (O_649,N_9978,N_9392);
and UO_650 (O_650,N_8716,N_9544);
nand UO_651 (O_651,N_9117,N_9459);
nand UO_652 (O_652,N_9450,N_9435);
or UO_653 (O_653,N_8274,N_7901);
or UO_654 (O_654,N_8126,N_7818);
or UO_655 (O_655,N_7516,N_7937);
or UO_656 (O_656,N_8607,N_8916);
nor UO_657 (O_657,N_8570,N_7909);
and UO_658 (O_658,N_9634,N_8944);
xor UO_659 (O_659,N_9480,N_9612);
or UO_660 (O_660,N_8321,N_8698);
xor UO_661 (O_661,N_8536,N_9188);
nor UO_662 (O_662,N_8055,N_8353);
or UO_663 (O_663,N_7951,N_9078);
nand UO_664 (O_664,N_9094,N_7931);
nor UO_665 (O_665,N_9532,N_8547);
nand UO_666 (O_666,N_7590,N_8490);
or UO_667 (O_667,N_9493,N_9946);
nand UO_668 (O_668,N_8645,N_9434);
nor UO_669 (O_669,N_8978,N_8972);
or UO_670 (O_670,N_8727,N_7670);
or UO_671 (O_671,N_8089,N_8539);
and UO_672 (O_672,N_8169,N_7691);
or UO_673 (O_673,N_8664,N_8173);
and UO_674 (O_674,N_9367,N_9470);
nor UO_675 (O_675,N_8479,N_7700);
xor UO_676 (O_676,N_9563,N_9841);
xnor UO_677 (O_677,N_9639,N_8209);
xnor UO_678 (O_678,N_8215,N_8888);
nand UO_679 (O_679,N_7521,N_9197);
nor UO_680 (O_680,N_9932,N_9466);
nor UO_681 (O_681,N_8082,N_9558);
nor UO_682 (O_682,N_9096,N_7771);
nor UO_683 (O_683,N_9409,N_9814);
xor UO_684 (O_684,N_9534,N_9673);
and UO_685 (O_685,N_7576,N_8167);
nor UO_686 (O_686,N_7519,N_8449);
nor UO_687 (O_687,N_7561,N_7534);
nor UO_688 (O_688,N_7877,N_8706);
nand UO_689 (O_689,N_8731,N_9669);
or UO_690 (O_690,N_9482,N_8488);
xnor UO_691 (O_691,N_9452,N_8515);
or UO_692 (O_692,N_7648,N_9717);
xor UO_693 (O_693,N_8592,N_9154);
xor UO_694 (O_694,N_8582,N_8998);
nand UO_695 (O_695,N_8163,N_7910);
and UO_696 (O_696,N_8086,N_9121);
and UO_697 (O_697,N_8996,N_7613);
nand UO_698 (O_698,N_9460,N_8980);
and UO_699 (O_699,N_9682,N_8020);
nor UO_700 (O_700,N_7606,N_8960);
xor UO_701 (O_701,N_9247,N_8270);
nand UO_702 (O_702,N_8556,N_8738);
or UO_703 (O_703,N_7591,N_8783);
nand UO_704 (O_704,N_8493,N_9107);
xor UO_705 (O_705,N_7965,N_8299);
nand UO_706 (O_706,N_9822,N_7674);
nand UO_707 (O_707,N_9429,N_9618);
nor UO_708 (O_708,N_7607,N_7531);
nand UO_709 (O_709,N_7506,N_7629);
xor UO_710 (O_710,N_8812,N_7907);
xnor UO_711 (O_711,N_9914,N_9736);
nor UO_712 (O_712,N_7902,N_8166);
nand UO_713 (O_713,N_8477,N_7685);
xnor UO_714 (O_714,N_8793,N_9041);
nor UO_715 (O_715,N_9898,N_8787);
and UO_716 (O_716,N_7944,N_9341);
and UO_717 (O_717,N_8955,N_7566);
nor UO_718 (O_718,N_8737,N_8613);
and UO_719 (O_719,N_7678,N_8037);
nand UO_720 (O_720,N_7751,N_8858);
xnor UO_721 (O_721,N_9926,N_8857);
nand UO_722 (O_722,N_8162,N_8369);
nand UO_723 (O_723,N_9285,N_9237);
xor UO_724 (O_724,N_9772,N_7778);
xnor UO_725 (O_725,N_8568,N_7970);
nand UO_726 (O_726,N_9525,N_8004);
xnor UO_727 (O_727,N_9922,N_9467);
and UO_728 (O_728,N_7508,N_9902);
and UO_729 (O_729,N_8651,N_8963);
nor UO_730 (O_730,N_9484,N_9334);
nand UO_731 (O_731,N_9010,N_9665);
nand UO_732 (O_732,N_9668,N_9820);
nor UO_733 (O_733,N_9537,N_7755);
nor UO_734 (O_734,N_9700,N_9997);
and UO_735 (O_735,N_9382,N_8496);
xnor UO_736 (O_736,N_8068,N_8302);
nor UO_737 (O_737,N_9851,N_9131);
xor UO_738 (O_738,N_9797,N_8976);
nor UO_739 (O_739,N_8583,N_8388);
or UO_740 (O_740,N_7604,N_8199);
and UO_741 (O_741,N_9082,N_7846);
nand UO_742 (O_742,N_8931,N_9623);
nand UO_743 (O_743,N_8711,N_8332);
nand UO_744 (O_744,N_8778,N_9301);
or UO_745 (O_745,N_8892,N_7997);
nand UO_746 (O_746,N_8874,N_7733);
xor UO_747 (O_747,N_9920,N_8752);
xnor UO_748 (O_748,N_8491,N_9652);
xor UO_749 (O_749,N_8233,N_9316);
nor UO_750 (O_750,N_8470,N_7945);
nor UO_751 (O_751,N_9227,N_9492);
or UO_752 (O_752,N_9825,N_8220);
and UO_753 (O_753,N_9601,N_8310);
and UO_754 (O_754,N_7819,N_8686);
xor UO_755 (O_755,N_8366,N_9093);
xor UO_756 (O_756,N_9426,N_9498);
nor UO_757 (O_757,N_8294,N_8827);
and UO_758 (O_758,N_9433,N_9539);
nand UO_759 (O_759,N_9875,N_8995);
and UO_760 (O_760,N_7663,N_8785);
and UO_761 (O_761,N_8198,N_8180);
and UO_762 (O_762,N_8759,N_8725);
or UO_763 (O_763,N_9818,N_9366);
nor UO_764 (O_764,N_8644,N_8307);
nor UO_765 (O_765,N_9505,N_9328);
nand UO_766 (O_766,N_9521,N_9326);
xor UO_767 (O_767,N_9163,N_8700);
and UO_768 (O_768,N_9077,N_8992);
or UO_769 (O_769,N_8452,N_9722);
xnor UO_770 (O_770,N_8581,N_7835);
nand UO_771 (O_771,N_9352,N_9080);
xor UO_772 (O_772,N_8217,N_8510);
or UO_773 (O_773,N_9266,N_7652);
nand UO_774 (O_774,N_7598,N_7917);
nor UO_775 (O_775,N_8925,N_9483);
xnor UO_776 (O_776,N_9776,N_9224);
xnor UO_777 (O_777,N_9454,N_8019);
or UO_778 (O_778,N_7862,N_9025);
nor UO_779 (O_779,N_9570,N_9344);
xor UO_780 (O_780,N_7588,N_7532);
and UO_781 (O_781,N_8550,N_8956);
nand UO_782 (O_782,N_9494,N_7839);
nand UO_783 (O_783,N_9307,N_9011);
nor UO_784 (O_784,N_9834,N_8360);
or UO_785 (O_785,N_9490,N_7924);
or UO_786 (O_786,N_7703,N_9294);
xor UO_787 (O_787,N_7649,N_7540);
or UO_788 (O_788,N_8560,N_8712);
nor UO_789 (O_789,N_8365,N_9827);
nor UO_790 (O_790,N_8303,N_8754);
and UO_791 (O_791,N_9973,N_9777);
and UO_792 (O_792,N_8070,N_8439);
or UO_793 (O_793,N_9583,N_8469);
or UO_794 (O_794,N_9387,N_7730);
or UO_795 (O_795,N_9112,N_9496);
nor UO_796 (O_796,N_9615,N_9549);
and UO_797 (O_797,N_8084,N_7502);
nor UO_798 (O_798,N_9891,N_8682);
and UO_799 (O_799,N_7581,N_8389);
or UO_800 (O_800,N_9934,N_8590);
or UO_801 (O_801,N_8964,N_8242);
nand UO_802 (O_802,N_9497,N_7609);
and UO_803 (O_803,N_8610,N_9507);
and UO_804 (O_804,N_9680,N_8842);
and UO_805 (O_805,N_8734,N_8723);
or UO_806 (O_806,N_9292,N_7585);
or UO_807 (O_807,N_9763,N_7824);
nand UO_808 (O_808,N_8848,N_7822);
nand UO_809 (O_809,N_7610,N_7647);
nor UO_810 (O_810,N_7876,N_9063);
nand UO_811 (O_811,N_7594,N_8519);
and UO_812 (O_812,N_8724,N_7883);
and UO_813 (O_813,N_9995,N_9162);
and UO_814 (O_814,N_8286,N_7734);
xnor UO_815 (O_815,N_9773,N_7675);
nand UO_816 (O_816,N_9391,N_9984);
and UO_817 (O_817,N_8101,N_8684);
or UO_818 (O_818,N_8474,N_8879);
xor UO_819 (O_819,N_7551,N_7993);
xor UO_820 (O_820,N_9611,N_8908);
and UO_821 (O_821,N_9232,N_9050);
xor UO_822 (O_822,N_9839,N_9478);
xnor UO_823 (O_823,N_8796,N_9903);
nor UO_824 (O_824,N_8052,N_7826);
nand UO_825 (O_825,N_9290,N_7927);
nor UO_826 (O_826,N_8256,N_9265);
and UO_827 (O_827,N_9239,N_8654);
or UO_828 (O_828,N_7920,N_9477);
nand UO_829 (O_829,N_9351,N_9071);
nor UO_830 (O_830,N_8283,N_9528);
nand UO_831 (O_831,N_9155,N_9743);
or UO_832 (O_832,N_8710,N_8988);
xor UO_833 (O_833,N_9255,N_8548);
or UO_834 (O_834,N_9602,N_9952);
nor UO_835 (O_835,N_7568,N_8322);
xor UO_836 (O_836,N_9949,N_7748);
nor UO_837 (O_837,N_9410,N_9782);
nand UO_838 (O_838,N_8967,N_8544);
nor UO_839 (O_839,N_9560,N_8514);
xor UO_840 (O_840,N_9759,N_9115);
and UO_841 (O_841,N_7799,N_8378);
nor UO_842 (O_842,N_9715,N_8061);
or UO_843 (O_843,N_8481,N_8056);
or UO_844 (O_844,N_8746,N_9899);
nor UO_845 (O_845,N_9681,N_9424);
and UO_846 (O_846,N_9823,N_8243);
nand UO_847 (O_847,N_9983,N_8704);
nor UO_848 (O_848,N_7567,N_9840);
and UO_849 (O_849,N_8249,N_7836);
or UO_850 (O_850,N_8328,N_9765);
nor UO_851 (O_851,N_7845,N_8589);
xnor UO_852 (O_852,N_9693,N_8355);
or UO_853 (O_853,N_8067,N_7892);
nand UO_854 (O_854,N_9506,N_9373);
nand UO_855 (O_855,N_7726,N_9201);
and UO_856 (O_856,N_9948,N_9176);
xnor UO_857 (O_857,N_9955,N_8938);
and UO_858 (O_858,N_8050,N_9177);
nor UO_859 (O_859,N_9076,N_9007);
and UO_860 (O_860,N_8588,N_8552);
nor UO_861 (O_861,N_9017,N_8110);
xnor UO_862 (O_862,N_9055,N_8211);
or UO_863 (O_863,N_7964,N_9769);
xnor UO_864 (O_864,N_9014,N_9550);
xor UO_865 (O_865,N_8015,N_8555);
or UO_866 (O_866,N_9256,N_9648);
nand UO_867 (O_867,N_7565,N_9485);
nor UO_868 (O_868,N_8563,N_7572);
nor UO_869 (O_869,N_8278,N_8142);
xnor UO_870 (O_870,N_7739,N_8175);
xor UO_871 (O_871,N_9911,N_8250);
and UO_872 (O_872,N_7875,N_9058);
xnor UO_873 (O_873,N_9168,N_9951);
or UO_874 (O_874,N_7804,N_9396);
nor UO_875 (O_875,N_8983,N_8609);
or UO_876 (O_876,N_9710,N_8666);
xnor UO_877 (O_877,N_9917,N_8003);
nor UO_878 (O_878,N_9453,N_7756);
xnor UO_879 (O_879,N_9748,N_8669);
or UO_880 (O_880,N_9921,N_9723);
nor UO_881 (O_881,N_8642,N_8832);
or UO_882 (O_882,N_9856,N_8692);
xnor UO_883 (O_883,N_9184,N_7548);
nand UO_884 (O_884,N_8508,N_8825);
nor UO_885 (O_885,N_7832,N_8231);
nand UO_886 (O_886,N_8766,N_9097);
xnor UO_887 (O_887,N_9510,N_8416);
nor UO_888 (O_888,N_8868,N_9938);
nand UO_889 (O_889,N_8210,N_9122);
nor UO_890 (O_890,N_7718,N_9553);
xor UO_891 (O_891,N_9873,N_9933);
nand UO_892 (O_892,N_7834,N_8415);
and UO_893 (O_893,N_7958,N_9222);
nor UO_894 (O_894,N_7599,N_8799);
and UO_895 (O_895,N_9637,N_9670);
and UO_896 (O_896,N_9214,N_8748);
or UO_897 (O_897,N_7843,N_7999);
nor UO_898 (O_898,N_7820,N_9440);
or UO_899 (O_899,N_9236,N_8141);
xor UO_900 (O_900,N_9286,N_8431);
nor UO_901 (O_901,N_8442,N_8333);
nand UO_902 (O_902,N_9034,N_8502);
nor UO_903 (O_903,N_9968,N_7833);
nor UO_904 (O_904,N_9702,N_7770);
nand UO_905 (O_905,N_8027,N_7968);
nand UO_906 (O_906,N_8383,N_8522);
nor UO_907 (O_907,N_8839,N_9701);
and UO_908 (O_908,N_9994,N_8813);
nor UO_909 (O_909,N_9906,N_7732);
nand UO_910 (O_910,N_8297,N_9306);
and UO_911 (O_911,N_9127,N_8202);
and UO_912 (O_912,N_7546,N_8803);
nand UO_913 (O_913,N_7681,N_9472);
or UO_914 (O_914,N_8473,N_9697);
xnor UO_915 (O_915,N_8922,N_9311);
and UO_916 (O_916,N_9551,N_8392);
and UO_917 (O_917,N_9318,N_9199);
nor UO_918 (O_918,N_9959,N_8891);
or UO_919 (O_919,N_8564,N_8314);
xnor UO_920 (O_920,N_8520,N_7640);
nand UO_921 (O_921,N_8183,N_9965);
xor UO_922 (O_922,N_9138,N_8317);
or UO_923 (O_923,N_9511,N_9264);
or UO_924 (O_924,N_7728,N_9847);
nor UO_925 (O_925,N_7644,N_8501);
and UO_926 (O_926,N_8033,N_9139);
or UO_927 (O_927,N_9635,N_7525);
and UO_928 (O_928,N_7825,N_9795);
or UO_929 (O_929,N_8285,N_9298);
xnor UO_930 (O_930,N_7922,N_8549);
or UO_931 (O_931,N_8853,N_8450);
and UO_932 (O_932,N_9786,N_9805);
nor UO_933 (O_933,N_7758,N_8300);
xor UO_934 (O_934,N_9109,N_9964);
and UO_935 (O_935,N_7714,N_8756);
and UO_936 (O_936,N_8444,N_9281);
nand UO_937 (O_937,N_7692,N_9288);
or UO_938 (O_938,N_8040,N_9803);
and UO_939 (O_939,N_9872,N_8240);
or UO_940 (O_940,N_9519,N_9678);
xnor UO_941 (O_941,N_8512,N_9566);
or UO_942 (O_942,N_9425,N_8072);
nor UO_943 (O_943,N_9514,N_7942);
or UO_944 (O_944,N_9761,N_9486);
and UO_945 (O_945,N_7994,N_9489);
and UO_946 (O_946,N_8078,N_8207);
or UO_947 (O_947,N_7864,N_7934);
nand UO_948 (O_948,N_8679,N_7708);
nand UO_949 (O_949,N_9542,N_9925);
xor UO_950 (O_950,N_7682,N_9074);
nor UO_951 (O_951,N_9401,N_8138);
or UO_952 (O_952,N_9577,N_8567);
or UO_953 (O_953,N_9631,N_7790);
nor UO_954 (O_954,N_7667,N_7616);
or UO_955 (O_955,N_8445,N_8280);
xor UO_956 (O_956,N_9568,N_8105);
xnor UO_957 (O_957,N_9408,N_7884);
nand UO_958 (O_958,N_7889,N_9719);
nor UO_959 (O_959,N_9880,N_8612);
nor UO_960 (O_960,N_8336,N_9893);
or UO_961 (O_961,N_7625,N_7780);
xor UO_962 (O_962,N_8707,N_8034);
and UO_963 (O_963,N_9734,N_8195);
nand UO_964 (O_964,N_9448,N_8694);
xor UO_965 (O_965,N_8675,N_7587);
nor UO_966 (O_966,N_8837,N_9473);
and UO_967 (O_967,N_8337,N_9090);
nand UO_968 (O_968,N_9961,N_7643);
nor UO_969 (O_969,N_7512,N_8002);
or UO_970 (O_970,N_9088,N_9947);
nor UO_971 (O_971,N_8403,N_9573);
nor UO_972 (O_972,N_9740,N_8236);
nor UO_973 (O_973,N_8289,N_8168);
nand UO_974 (O_974,N_9745,N_8397);
and UO_975 (O_975,N_8363,N_9136);
nor UO_976 (O_976,N_8238,N_8968);
nor UO_977 (O_977,N_9884,N_7912);
nor UO_978 (O_978,N_8076,N_7620);
or UO_979 (O_979,N_8975,N_7503);
or UO_980 (O_980,N_8965,N_8933);
nand UO_981 (O_981,N_8035,N_9220);
and UO_982 (O_982,N_9546,N_8618);
or UO_983 (O_983,N_8085,N_7961);
nand UO_984 (O_984,N_7611,N_9364);
xnor UO_985 (O_985,N_9116,N_9449);
and UO_986 (O_986,N_8831,N_8554);
nor UO_987 (O_987,N_8083,N_7507);
nand UO_988 (O_988,N_9515,N_9954);
or UO_989 (O_989,N_8834,N_8264);
and UO_990 (O_990,N_7657,N_8060);
and UO_991 (O_991,N_9787,N_8036);
nand UO_992 (O_992,N_8794,N_7874);
xnor UO_993 (O_993,N_7966,N_8343);
xor UO_994 (O_994,N_8531,N_8646);
nand UO_995 (O_995,N_8518,N_9835);
and UO_996 (O_996,N_8718,N_8402);
nor UO_997 (O_997,N_9886,N_8601);
and UO_998 (O_998,N_8709,N_9928);
xnor UO_999 (O_999,N_7837,N_8952);
and UO_1000 (O_1000,N_7813,N_8472);
nor UO_1001 (O_1001,N_9279,N_8009);
nand UO_1002 (O_1002,N_9012,N_8170);
or UO_1003 (O_1003,N_7582,N_8192);
or UO_1004 (O_1004,N_8467,N_7776);
or UO_1005 (O_1005,N_8172,N_8345);
nand UO_1006 (O_1006,N_8106,N_8740);
nand UO_1007 (O_1007,N_8356,N_7929);
nand UO_1008 (O_1008,N_9043,N_9720);
nand UO_1009 (O_1009,N_8193,N_8905);
nor UO_1010 (O_1010,N_9253,N_9123);
xor UO_1011 (O_1011,N_8282,N_9217);
nor UO_1012 (O_1012,N_7911,N_8934);
nand UO_1013 (O_1013,N_9458,N_8011);
nand UO_1014 (O_1014,N_9654,N_8427);
or UO_1015 (O_1015,N_7575,N_9590);
and UO_1016 (O_1016,N_8010,N_8571);
or UO_1017 (O_1017,N_8843,N_8484);
nand UO_1018 (O_1018,N_9616,N_8241);
nor UO_1019 (O_1019,N_8958,N_8156);
nand UO_1020 (O_1020,N_9696,N_9182);
xnor UO_1021 (O_1021,N_7991,N_8757);
nor UO_1022 (O_1022,N_7558,N_8177);
or UO_1023 (O_1023,N_9499,N_9042);
nand UO_1024 (O_1024,N_9081,N_8772);
nor UO_1025 (O_1025,N_7885,N_7933);
xor UO_1026 (O_1026,N_9649,N_9684);
xnor UO_1027 (O_1027,N_9092,N_8569);
xor UO_1028 (O_1028,N_8487,N_8545);
and UO_1029 (O_1029,N_8650,N_7699);
nand UO_1030 (O_1030,N_8097,N_9992);
and UO_1031 (O_1031,N_7980,N_8124);
nand UO_1032 (O_1032,N_8715,N_7926);
nor UO_1033 (O_1033,N_9529,N_9713);
xnor UO_1034 (O_1034,N_8728,N_9249);
xor UO_1035 (O_1035,N_8391,N_9075);
and UO_1036 (O_1036,N_7740,N_9151);
or UO_1037 (O_1037,N_8404,N_9754);
and UO_1038 (O_1038,N_8296,N_8897);
xnor UO_1039 (O_1039,N_9293,N_9837);
nor UO_1040 (O_1040,N_8946,N_8251);
xor UO_1041 (O_1041,N_8305,N_8674);
xor UO_1042 (O_1042,N_9561,N_9931);
and UO_1043 (O_1043,N_9174,N_7605);
xnor UO_1044 (O_1044,N_7987,N_7842);
and UO_1045 (O_1045,N_9988,N_7586);
or UO_1046 (O_1046,N_9444,N_8461);
nand UO_1047 (O_1047,N_8131,N_9468);
or UO_1048 (O_1048,N_8776,N_8354);
nand UO_1049 (O_1049,N_9937,N_7880);
xnor UO_1050 (O_1050,N_9704,N_7602);
xnor UO_1051 (O_1051,N_8237,N_8851);
or UO_1052 (O_1052,N_9234,N_7866);
nor UO_1053 (O_1053,N_8352,N_8846);
nand UO_1054 (O_1054,N_7882,N_9939);
and UO_1055 (O_1055,N_9393,N_9377);
or UO_1056 (O_1056,N_7650,N_8121);
nand UO_1057 (O_1057,N_8102,N_8572);
or UO_1058 (O_1058,N_7763,N_7660);
nand UO_1059 (O_1059,N_9385,N_9565);
and UO_1060 (O_1060,N_8406,N_8987);
or UO_1061 (O_1061,N_8482,N_8214);
nor UO_1062 (O_1062,N_9361,N_9087);
nand UO_1063 (O_1063,N_9643,N_8182);
or UO_1064 (O_1064,N_8123,N_7905);
nand UO_1065 (O_1065,N_8434,N_8760);
or UO_1066 (O_1066,N_8134,N_8185);
or UO_1067 (O_1067,N_7900,N_9374);
or UO_1068 (O_1068,N_9889,N_8949);
or UO_1069 (O_1069,N_8896,N_8136);
nor UO_1070 (O_1070,N_9821,N_8509);
and UO_1071 (O_1071,N_7526,N_8959);
nand UO_1072 (O_1072,N_8244,N_8751);
or UO_1073 (O_1073,N_8890,N_8818);
xor UO_1074 (O_1074,N_9104,N_9912);
and UO_1075 (O_1075,N_9619,N_8100);
xor UO_1076 (O_1076,N_9195,N_7858);
and UO_1077 (O_1077,N_8873,N_9167);
nor UO_1078 (O_1078,N_8807,N_9645);
xnor UO_1079 (O_1079,N_9683,N_9685);
or UO_1080 (O_1080,N_8819,N_7689);
xor UO_1081 (O_1081,N_9287,N_8900);
and UO_1082 (O_1082,N_8483,N_8247);
nand UO_1083 (O_1083,N_9390,N_8462);
and UO_1084 (O_1084,N_7717,N_9323);
xor UO_1085 (O_1085,N_8611,N_9950);
xor UO_1086 (O_1086,N_7634,N_7706);
nor UO_1087 (O_1087,N_7530,N_9698);
nand UO_1088 (O_1088,N_7995,N_7899);
and UO_1089 (O_1089,N_8678,N_9465);
or UO_1090 (O_1090,N_9488,N_7684);
nor UO_1091 (O_1091,N_8139,N_9016);
and UO_1092 (O_1092,N_8463,N_8774);
or UO_1093 (O_1093,N_9858,N_8932);
xor UO_1094 (O_1094,N_7873,N_8429);
xor UO_1095 (O_1095,N_8824,N_8200);
or UO_1096 (O_1096,N_9170,N_8677);
and UO_1097 (O_1097,N_8855,N_9571);
nor UO_1098 (O_1098,N_8507,N_8779);
nand UO_1099 (O_1099,N_8330,N_8338);
xnor UO_1100 (O_1100,N_9171,N_9541);
nand UO_1101 (O_1101,N_7518,N_7960);
nand UO_1102 (O_1102,N_8817,N_8947);
nor UO_1103 (O_1103,N_8641,N_9108);
nand UO_1104 (O_1104,N_8197,N_7895);
or UO_1105 (O_1105,N_7894,N_7761);
nor UO_1106 (O_1106,N_8357,N_8929);
xor UO_1107 (O_1107,N_8206,N_9867);
nor UO_1108 (O_1108,N_8430,N_9595);
and UO_1109 (O_1109,N_9881,N_8372);
nor UO_1110 (O_1110,N_9508,N_8042);
or UO_1111 (O_1111,N_8181,N_9166);
xnor UO_1112 (O_1112,N_9084,N_9044);
nand UO_1113 (O_1113,N_8735,N_8997);
nand UO_1114 (O_1114,N_8128,N_8301);
nor UO_1115 (O_1115,N_9989,N_9405);
nor UO_1116 (O_1116,N_7979,N_9663);
or UO_1117 (O_1117,N_7671,N_8224);
and UO_1118 (O_1118,N_8667,N_9552);
and UO_1119 (O_1119,N_9029,N_8656);
nand UO_1120 (O_1120,N_9651,N_9716);
and UO_1121 (O_1121,N_7727,N_9725);
or UO_1122 (O_1122,N_8745,N_8721);
and UO_1123 (O_1123,N_9024,N_7536);
or UO_1124 (O_1124,N_8418,N_7957);
xnor UO_1125 (O_1125,N_9614,N_9411);
or UO_1126 (O_1126,N_8971,N_9380);
and UO_1127 (O_1127,N_7787,N_9158);
xnor UO_1128 (O_1128,N_9057,N_9430);
xor UO_1129 (O_1129,N_9985,N_9826);
and UO_1130 (O_1130,N_8791,N_8860);
nor UO_1131 (O_1131,N_8205,N_9957);
and UO_1132 (O_1132,N_7851,N_8395);
nand UO_1133 (O_1133,N_8697,N_9699);
xnor UO_1134 (O_1134,N_8504,N_8277);
xor UO_1135 (O_1135,N_9130,N_8844);
and UO_1136 (O_1136,N_8058,N_8120);
and UO_1137 (O_1137,N_9557,N_8133);
xor UO_1138 (O_1138,N_9675,N_9667);
nand UO_1139 (O_1139,N_8829,N_8566);
or UO_1140 (O_1140,N_9609,N_8419);
nor UO_1141 (O_1141,N_9603,N_9526);
xor UO_1142 (O_1142,N_7983,N_7500);
or UO_1143 (O_1143,N_7893,N_8630);
nand UO_1144 (O_1144,N_8881,N_7745);
or UO_1145 (O_1145,N_7793,N_8316);
and UO_1146 (O_1146,N_9277,N_9309);
or UO_1147 (O_1147,N_7735,N_9810);
xor UO_1148 (O_1148,N_9441,N_8627);
nand UO_1149 (O_1149,N_7533,N_8308);
and UO_1150 (O_1150,N_8318,N_8770);
xnor UO_1151 (O_1151,N_8647,N_9714);
nor UO_1152 (O_1152,N_8722,N_9883);
xnor UO_1153 (O_1153,N_8053,N_7543);
or UO_1154 (O_1154,N_9966,N_8154);
nand UO_1155 (O_1155,N_8435,N_8528);
nor UO_1156 (O_1156,N_7849,N_9173);
xor UO_1157 (O_1157,N_8882,N_8546);
or UO_1158 (O_1158,N_8657,N_9003);
xnor UO_1159 (O_1159,N_7639,N_8798);
or UO_1160 (O_1160,N_7666,N_8455);
or UO_1161 (O_1161,N_9359,N_8340);
and UO_1162 (O_1162,N_7802,N_7716);
and UO_1163 (O_1163,N_8371,N_7680);
nand UO_1164 (O_1164,N_8623,N_9461);
nor UO_1165 (O_1165,N_8320,N_9083);
xor UO_1166 (O_1166,N_8950,N_9885);
and UO_1167 (O_1167,N_8228,N_7559);
xnor UO_1168 (O_1168,N_9319,N_7529);
nand UO_1169 (O_1169,N_8758,N_9297);
xnor UO_1170 (O_1170,N_9605,N_7601);
and UO_1171 (O_1171,N_9575,N_8529);
xnor UO_1172 (O_1172,N_8557,N_8313);
nand UO_1173 (O_1173,N_7677,N_8688);
nand UO_1174 (O_1174,N_9178,N_9916);
and UO_1175 (O_1175,N_7711,N_8188);
nor UO_1176 (O_1176,N_9120,N_9892);
nand UO_1177 (O_1177,N_9543,N_7552);
nor UO_1178 (O_1178,N_8942,N_8339);
or UO_1179 (O_1179,N_9132,N_9073);
xnor UO_1180 (O_1180,N_8970,N_7803);
or UO_1181 (O_1181,N_8292,N_7938);
and UO_1182 (O_1182,N_8041,N_9273);
xnor UO_1183 (O_1183,N_9263,N_7614);
nand UO_1184 (O_1184,N_7555,N_9808);
xnor UO_1185 (O_1185,N_7628,N_9372);
xor UO_1186 (O_1186,N_8867,N_9267);
nor UO_1187 (O_1187,N_8203,N_7624);
nand UO_1188 (O_1188,N_7886,N_8986);
nand UO_1189 (O_1189,N_9451,N_9969);
and UO_1190 (O_1190,N_8695,N_7623);
or UO_1191 (O_1191,N_9354,N_8005);
nand UO_1192 (O_1192,N_9807,N_8309);
nand UO_1193 (O_1193,N_9062,N_8411);
xor UO_1194 (O_1194,N_9476,N_7705);
and UO_1195 (O_1195,N_7808,N_9368);
xnor UO_1196 (O_1196,N_7619,N_9811);
nor UO_1197 (O_1197,N_8620,N_9291);
or UO_1198 (O_1198,N_9110,N_9646);
xnor UO_1199 (O_1199,N_8298,N_8229);
or UO_1200 (O_1200,N_7765,N_7996);
or UO_1201 (O_1201,N_9446,N_7925);
nor UO_1202 (O_1202,N_9874,N_7935);
xnor UO_1203 (O_1203,N_9691,N_8792);
xnor UO_1204 (O_1204,N_9246,N_7557);
nand UO_1205 (O_1205,N_9861,N_8521);
or UO_1206 (O_1206,N_9689,N_9940);
xor UO_1207 (O_1207,N_9419,N_7710);
nand UO_1208 (O_1208,N_9325,N_8458);
xor UO_1209 (O_1209,N_9128,N_9282);
nand UO_1210 (O_1210,N_9250,N_7879);
nor UO_1211 (O_1211,N_7626,N_9677);
nor UO_1212 (O_1212,N_8871,N_8021);
xor UO_1213 (O_1213,N_8016,N_8661);
nor UO_1214 (O_1214,N_9272,N_9395);
and UO_1215 (O_1215,N_8615,N_9794);
and UO_1216 (O_1216,N_8171,N_9569);
or UO_1217 (O_1217,N_9194,N_8438);
and UO_1218 (O_1218,N_9332,N_7829);
or UO_1219 (O_1219,N_9904,N_9991);
nand UO_1220 (O_1220,N_9793,N_7998);
and UO_1221 (O_1221,N_9705,N_9375);
or UO_1222 (O_1222,N_8263,N_7777);
xnor UO_1223 (O_1223,N_8232,N_9531);
or UO_1224 (O_1224,N_7544,N_9842);
xor UO_1225 (O_1225,N_7510,N_9054);
or UO_1226 (O_1226,N_8451,N_8767);
or UO_1227 (O_1227,N_8885,N_9672);
or UO_1228 (O_1228,N_8373,N_8624);
xor UO_1229 (O_1229,N_8806,N_8591);
xnor UO_1230 (O_1230,N_8125,N_9059);
nand UO_1231 (O_1231,N_9463,N_7865);
and UO_1232 (O_1232,N_8634,N_9836);
nor UO_1233 (O_1233,N_9630,N_9538);
nor UO_1234 (O_1234,N_7673,N_8786);
xnor UO_1235 (O_1235,N_9462,N_8535);
nor UO_1236 (O_1236,N_8587,N_9963);
and UO_1237 (O_1237,N_7940,N_8573);
nor UO_1238 (O_1238,N_7798,N_9052);
xor UO_1239 (O_1239,N_7962,N_9455);
nor UO_1240 (O_1240,N_8073,N_9312);
xor UO_1241 (O_1241,N_8262,N_8865);
nand UO_1242 (O_1242,N_9175,N_7779);
xor UO_1243 (O_1243,N_7992,N_8585);
nor UO_1244 (O_1244,N_9056,N_7592);
and UO_1245 (O_1245,N_9897,N_7511);
xor UO_1246 (O_1246,N_9767,N_8026);
nor UO_1247 (O_1247,N_7913,N_9124);
xnor UO_1248 (O_1248,N_9313,N_7553);
nor UO_1249 (O_1249,N_9986,N_7584);
xor UO_1250 (O_1250,N_8206,N_9977);
xnor UO_1251 (O_1251,N_9441,N_9289);
nand UO_1252 (O_1252,N_8572,N_9071);
nor UO_1253 (O_1253,N_8016,N_8647);
nor UO_1254 (O_1254,N_9499,N_7970);
and UO_1255 (O_1255,N_7552,N_9469);
or UO_1256 (O_1256,N_7960,N_7687);
xor UO_1257 (O_1257,N_9934,N_7912);
nor UO_1258 (O_1258,N_7687,N_9483);
or UO_1259 (O_1259,N_7679,N_8181);
and UO_1260 (O_1260,N_9328,N_7711);
xor UO_1261 (O_1261,N_7945,N_9704);
nand UO_1262 (O_1262,N_9994,N_9022);
nor UO_1263 (O_1263,N_9391,N_7568);
or UO_1264 (O_1264,N_8456,N_7887);
and UO_1265 (O_1265,N_9948,N_8239);
nor UO_1266 (O_1266,N_9140,N_7570);
nand UO_1267 (O_1267,N_9107,N_9569);
xnor UO_1268 (O_1268,N_9680,N_9390);
or UO_1269 (O_1269,N_8739,N_7862);
nand UO_1270 (O_1270,N_9502,N_9158);
nor UO_1271 (O_1271,N_9071,N_8485);
xor UO_1272 (O_1272,N_9561,N_7625);
or UO_1273 (O_1273,N_9213,N_8160);
nor UO_1274 (O_1274,N_7920,N_9857);
nor UO_1275 (O_1275,N_8335,N_7767);
nand UO_1276 (O_1276,N_8265,N_8745);
xor UO_1277 (O_1277,N_8630,N_9709);
nand UO_1278 (O_1278,N_9150,N_7949);
and UO_1279 (O_1279,N_8526,N_9527);
and UO_1280 (O_1280,N_8470,N_9811);
and UO_1281 (O_1281,N_7958,N_9066);
and UO_1282 (O_1282,N_8152,N_9194);
nor UO_1283 (O_1283,N_8022,N_7535);
nor UO_1284 (O_1284,N_8263,N_8957);
and UO_1285 (O_1285,N_9752,N_8484);
nor UO_1286 (O_1286,N_8611,N_8494);
nor UO_1287 (O_1287,N_8886,N_8695);
and UO_1288 (O_1288,N_8996,N_9959);
nand UO_1289 (O_1289,N_7623,N_8029);
nand UO_1290 (O_1290,N_9972,N_9291);
xor UO_1291 (O_1291,N_9369,N_8361);
xor UO_1292 (O_1292,N_9076,N_9466);
xnor UO_1293 (O_1293,N_8835,N_9734);
or UO_1294 (O_1294,N_7663,N_9127);
nand UO_1295 (O_1295,N_9172,N_9290);
xor UO_1296 (O_1296,N_9660,N_9673);
and UO_1297 (O_1297,N_9564,N_8755);
and UO_1298 (O_1298,N_8767,N_8554);
or UO_1299 (O_1299,N_8292,N_9595);
or UO_1300 (O_1300,N_8389,N_9899);
nand UO_1301 (O_1301,N_8415,N_9642);
nand UO_1302 (O_1302,N_8274,N_9186);
nand UO_1303 (O_1303,N_8844,N_8880);
xor UO_1304 (O_1304,N_8035,N_7750);
or UO_1305 (O_1305,N_9920,N_9684);
nand UO_1306 (O_1306,N_9783,N_9174);
nand UO_1307 (O_1307,N_9093,N_8942);
and UO_1308 (O_1308,N_7593,N_8792);
nand UO_1309 (O_1309,N_8209,N_8389);
nand UO_1310 (O_1310,N_9906,N_8155);
and UO_1311 (O_1311,N_9730,N_9588);
or UO_1312 (O_1312,N_9027,N_8189);
nor UO_1313 (O_1313,N_8928,N_9063);
and UO_1314 (O_1314,N_9350,N_8889);
nor UO_1315 (O_1315,N_8712,N_8873);
nand UO_1316 (O_1316,N_7729,N_8150);
and UO_1317 (O_1317,N_8357,N_8069);
or UO_1318 (O_1318,N_7994,N_9771);
xor UO_1319 (O_1319,N_9527,N_9490);
nor UO_1320 (O_1320,N_9528,N_9857);
and UO_1321 (O_1321,N_9720,N_8227);
xnor UO_1322 (O_1322,N_9848,N_9171);
nand UO_1323 (O_1323,N_9853,N_8533);
or UO_1324 (O_1324,N_7939,N_9991);
nor UO_1325 (O_1325,N_8110,N_9267);
or UO_1326 (O_1326,N_7730,N_7525);
nand UO_1327 (O_1327,N_8330,N_9939);
xor UO_1328 (O_1328,N_9575,N_8145);
or UO_1329 (O_1329,N_7561,N_8936);
and UO_1330 (O_1330,N_8466,N_9827);
nand UO_1331 (O_1331,N_8054,N_8255);
nand UO_1332 (O_1332,N_8218,N_8786);
and UO_1333 (O_1333,N_9042,N_9375);
xor UO_1334 (O_1334,N_8342,N_7686);
xor UO_1335 (O_1335,N_8132,N_9616);
or UO_1336 (O_1336,N_9164,N_8966);
nand UO_1337 (O_1337,N_8215,N_8536);
xnor UO_1338 (O_1338,N_8506,N_7851);
nand UO_1339 (O_1339,N_7936,N_9278);
or UO_1340 (O_1340,N_9183,N_8818);
nor UO_1341 (O_1341,N_9055,N_8389);
nor UO_1342 (O_1342,N_9706,N_8675);
or UO_1343 (O_1343,N_8527,N_8608);
or UO_1344 (O_1344,N_8181,N_9448);
or UO_1345 (O_1345,N_8612,N_8471);
and UO_1346 (O_1346,N_8157,N_7788);
nand UO_1347 (O_1347,N_7592,N_7917);
and UO_1348 (O_1348,N_9038,N_8759);
nor UO_1349 (O_1349,N_9691,N_8950);
or UO_1350 (O_1350,N_8980,N_7808);
nand UO_1351 (O_1351,N_9110,N_7946);
and UO_1352 (O_1352,N_9805,N_8244);
and UO_1353 (O_1353,N_9703,N_8964);
or UO_1354 (O_1354,N_7796,N_8292);
or UO_1355 (O_1355,N_9776,N_7887);
or UO_1356 (O_1356,N_8090,N_8648);
and UO_1357 (O_1357,N_8750,N_8318);
or UO_1358 (O_1358,N_8076,N_7621);
xor UO_1359 (O_1359,N_8013,N_8450);
and UO_1360 (O_1360,N_9751,N_9293);
xor UO_1361 (O_1361,N_8375,N_7754);
xnor UO_1362 (O_1362,N_9068,N_9926);
nand UO_1363 (O_1363,N_9567,N_8319);
nand UO_1364 (O_1364,N_7665,N_8781);
nand UO_1365 (O_1365,N_9999,N_9846);
or UO_1366 (O_1366,N_9361,N_7737);
and UO_1367 (O_1367,N_9540,N_7834);
or UO_1368 (O_1368,N_9697,N_8481);
xnor UO_1369 (O_1369,N_8685,N_8051);
nor UO_1370 (O_1370,N_9569,N_8018);
and UO_1371 (O_1371,N_8677,N_9213);
nand UO_1372 (O_1372,N_8768,N_7748);
nor UO_1373 (O_1373,N_9775,N_9393);
nand UO_1374 (O_1374,N_9263,N_9304);
xnor UO_1375 (O_1375,N_8812,N_7611);
nor UO_1376 (O_1376,N_7537,N_9137);
or UO_1377 (O_1377,N_8551,N_8597);
and UO_1378 (O_1378,N_8717,N_9748);
nor UO_1379 (O_1379,N_9272,N_8575);
xor UO_1380 (O_1380,N_8479,N_9663);
nor UO_1381 (O_1381,N_9566,N_9425);
and UO_1382 (O_1382,N_9311,N_9765);
and UO_1383 (O_1383,N_9569,N_9796);
or UO_1384 (O_1384,N_9857,N_8853);
nor UO_1385 (O_1385,N_8923,N_9650);
nor UO_1386 (O_1386,N_8411,N_7629);
xor UO_1387 (O_1387,N_9202,N_7954);
nand UO_1388 (O_1388,N_7925,N_8509);
and UO_1389 (O_1389,N_8644,N_7573);
or UO_1390 (O_1390,N_8941,N_8728);
and UO_1391 (O_1391,N_8931,N_9732);
xor UO_1392 (O_1392,N_8861,N_9250);
or UO_1393 (O_1393,N_8325,N_8067);
nor UO_1394 (O_1394,N_9772,N_8941);
and UO_1395 (O_1395,N_7501,N_8970);
nor UO_1396 (O_1396,N_9378,N_9333);
or UO_1397 (O_1397,N_8007,N_9028);
and UO_1398 (O_1398,N_9866,N_8170);
xor UO_1399 (O_1399,N_8186,N_9005);
or UO_1400 (O_1400,N_9585,N_8909);
and UO_1401 (O_1401,N_7730,N_7858);
nand UO_1402 (O_1402,N_8466,N_9229);
xnor UO_1403 (O_1403,N_8119,N_7966);
nand UO_1404 (O_1404,N_9374,N_8995);
nor UO_1405 (O_1405,N_8276,N_8596);
nand UO_1406 (O_1406,N_9083,N_9012);
xor UO_1407 (O_1407,N_8376,N_7759);
nand UO_1408 (O_1408,N_9597,N_8187);
nand UO_1409 (O_1409,N_7669,N_8014);
xor UO_1410 (O_1410,N_9027,N_8975);
nor UO_1411 (O_1411,N_7518,N_7966);
and UO_1412 (O_1412,N_8040,N_8288);
nand UO_1413 (O_1413,N_8927,N_9637);
or UO_1414 (O_1414,N_9936,N_7772);
and UO_1415 (O_1415,N_9681,N_8540);
xor UO_1416 (O_1416,N_9590,N_9588);
xor UO_1417 (O_1417,N_9323,N_9155);
or UO_1418 (O_1418,N_8736,N_9517);
nand UO_1419 (O_1419,N_9238,N_9333);
or UO_1420 (O_1420,N_9764,N_8309);
nor UO_1421 (O_1421,N_8889,N_8346);
and UO_1422 (O_1422,N_8760,N_7760);
xnor UO_1423 (O_1423,N_8251,N_9712);
nand UO_1424 (O_1424,N_8014,N_9493);
nor UO_1425 (O_1425,N_9104,N_9769);
and UO_1426 (O_1426,N_8382,N_7891);
and UO_1427 (O_1427,N_8017,N_8388);
nor UO_1428 (O_1428,N_8041,N_8006);
xor UO_1429 (O_1429,N_8329,N_7913);
nand UO_1430 (O_1430,N_9139,N_9966);
xnor UO_1431 (O_1431,N_8493,N_7569);
or UO_1432 (O_1432,N_8283,N_8937);
or UO_1433 (O_1433,N_9057,N_9506);
nand UO_1434 (O_1434,N_7655,N_8348);
and UO_1435 (O_1435,N_8519,N_8400);
nor UO_1436 (O_1436,N_8202,N_8069);
and UO_1437 (O_1437,N_8621,N_8576);
and UO_1438 (O_1438,N_9385,N_8857);
xnor UO_1439 (O_1439,N_7921,N_9711);
nand UO_1440 (O_1440,N_8710,N_8322);
or UO_1441 (O_1441,N_8774,N_8477);
nor UO_1442 (O_1442,N_8447,N_7660);
and UO_1443 (O_1443,N_8960,N_9944);
nand UO_1444 (O_1444,N_9427,N_9950);
nand UO_1445 (O_1445,N_8182,N_7954);
nor UO_1446 (O_1446,N_9511,N_8787);
or UO_1447 (O_1447,N_9707,N_9141);
xnor UO_1448 (O_1448,N_9000,N_8615);
nor UO_1449 (O_1449,N_7762,N_7612);
nand UO_1450 (O_1450,N_9331,N_8188);
or UO_1451 (O_1451,N_9687,N_9784);
nor UO_1452 (O_1452,N_8562,N_9518);
and UO_1453 (O_1453,N_7779,N_9532);
or UO_1454 (O_1454,N_8718,N_7902);
and UO_1455 (O_1455,N_9782,N_9363);
xor UO_1456 (O_1456,N_8359,N_9571);
and UO_1457 (O_1457,N_8726,N_9564);
and UO_1458 (O_1458,N_9489,N_8723);
or UO_1459 (O_1459,N_8020,N_8066);
nor UO_1460 (O_1460,N_7838,N_7528);
or UO_1461 (O_1461,N_9072,N_9080);
xnor UO_1462 (O_1462,N_7943,N_8772);
or UO_1463 (O_1463,N_9902,N_8130);
and UO_1464 (O_1464,N_8647,N_8418);
nor UO_1465 (O_1465,N_9736,N_8392);
xnor UO_1466 (O_1466,N_9640,N_9542);
or UO_1467 (O_1467,N_9186,N_8585);
and UO_1468 (O_1468,N_9982,N_9969);
or UO_1469 (O_1469,N_9353,N_8140);
nor UO_1470 (O_1470,N_7864,N_7553);
nor UO_1471 (O_1471,N_8359,N_8977);
or UO_1472 (O_1472,N_8158,N_9015);
xor UO_1473 (O_1473,N_7659,N_8399);
or UO_1474 (O_1474,N_9260,N_8322);
or UO_1475 (O_1475,N_7686,N_9198);
and UO_1476 (O_1476,N_9314,N_8328);
nor UO_1477 (O_1477,N_9705,N_9837);
nand UO_1478 (O_1478,N_9538,N_9984);
nand UO_1479 (O_1479,N_8093,N_9082);
nand UO_1480 (O_1480,N_9839,N_8973);
and UO_1481 (O_1481,N_8377,N_8193);
xnor UO_1482 (O_1482,N_7938,N_8885);
nor UO_1483 (O_1483,N_8757,N_9035);
or UO_1484 (O_1484,N_8898,N_8303);
xnor UO_1485 (O_1485,N_8682,N_9598);
and UO_1486 (O_1486,N_8377,N_9067);
and UO_1487 (O_1487,N_9038,N_8136);
or UO_1488 (O_1488,N_8940,N_9403);
nor UO_1489 (O_1489,N_9945,N_8685);
and UO_1490 (O_1490,N_8100,N_7787);
nor UO_1491 (O_1491,N_9827,N_8903);
xor UO_1492 (O_1492,N_9387,N_8280);
and UO_1493 (O_1493,N_8921,N_7954);
or UO_1494 (O_1494,N_9925,N_7549);
and UO_1495 (O_1495,N_8264,N_8650);
nor UO_1496 (O_1496,N_8828,N_8142);
nand UO_1497 (O_1497,N_9361,N_9449);
nor UO_1498 (O_1498,N_9821,N_9901);
nand UO_1499 (O_1499,N_8683,N_8649);
endmodule