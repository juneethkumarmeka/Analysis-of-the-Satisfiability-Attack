module basic_500_3000_500_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_100,In_316);
or U1 (N_1,In_81,In_193);
or U2 (N_2,In_480,In_459);
nand U3 (N_3,In_268,In_447);
and U4 (N_4,In_61,In_138);
and U5 (N_5,In_259,In_214);
xnor U6 (N_6,In_420,In_494);
xor U7 (N_7,In_261,In_102);
or U8 (N_8,In_51,In_380);
nor U9 (N_9,In_19,In_91);
nand U10 (N_10,In_310,In_256);
and U11 (N_11,In_129,In_250);
nor U12 (N_12,In_74,In_416);
or U13 (N_13,In_403,In_121);
and U14 (N_14,In_495,In_169);
or U15 (N_15,In_227,In_435);
and U16 (N_16,In_251,In_392);
or U17 (N_17,In_276,In_49);
or U18 (N_18,In_341,In_181);
or U19 (N_19,In_84,In_455);
or U20 (N_20,In_357,In_212);
or U21 (N_21,In_104,In_389);
or U22 (N_22,In_469,In_474);
and U23 (N_23,In_188,In_233);
nand U24 (N_24,In_490,In_153);
nand U25 (N_25,In_488,In_364);
and U26 (N_26,In_171,In_359);
xnor U27 (N_27,In_228,In_203);
or U28 (N_28,In_56,In_464);
and U29 (N_29,In_471,In_194);
and U30 (N_30,In_337,In_429);
nand U31 (N_31,In_77,In_344);
xor U32 (N_32,In_30,In_462);
or U33 (N_33,In_98,In_85);
and U34 (N_34,In_107,In_334);
xnor U35 (N_35,In_140,In_443);
or U36 (N_36,In_299,In_406);
nor U37 (N_37,In_90,In_279);
and U38 (N_38,In_387,In_286);
xor U39 (N_39,In_108,In_208);
nand U40 (N_40,In_277,In_249);
or U41 (N_41,In_12,In_80);
xnor U42 (N_42,In_426,In_313);
xnor U43 (N_43,In_444,In_258);
nand U44 (N_44,In_161,In_178);
xnor U45 (N_45,In_65,In_103);
xnor U46 (N_46,In_473,In_69);
xnor U47 (N_47,In_42,In_385);
nand U48 (N_48,In_144,In_418);
or U49 (N_49,In_309,In_283);
nand U50 (N_50,In_175,In_423);
or U51 (N_51,In_67,In_115);
nand U52 (N_52,In_37,In_430);
nor U53 (N_53,In_127,In_457);
xnor U54 (N_54,In_415,In_89);
and U55 (N_55,In_7,In_45);
nand U56 (N_56,In_340,In_266);
xor U57 (N_57,In_305,In_414);
xor U58 (N_58,In_463,In_489);
and U59 (N_59,In_396,In_157);
or U60 (N_60,In_167,In_219);
and U61 (N_61,In_246,In_395);
nand U62 (N_62,In_59,In_441);
or U63 (N_63,In_232,In_26);
or U64 (N_64,In_238,In_29);
nand U65 (N_65,In_215,In_173);
nor U66 (N_66,In_141,In_314);
and U67 (N_67,In_295,In_269);
nand U68 (N_68,In_252,In_497);
or U69 (N_69,In_271,In_163);
and U70 (N_70,In_476,In_202);
nor U71 (N_71,In_148,In_165);
xor U72 (N_72,In_413,In_105);
or U73 (N_73,In_343,In_240);
or U74 (N_74,In_123,In_466);
and U75 (N_75,In_382,In_460);
xor U76 (N_76,In_330,In_290);
nor U77 (N_77,In_3,In_86);
nor U78 (N_78,In_366,In_159);
and U79 (N_79,In_229,In_437);
or U80 (N_80,In_231,In_199);
nor U81 (N_81,In_483,In_36);
or U82 (N_82,In_301,In_472);
nand U83 (N_83,In_216,In_94);
nand U84 (N_84,In_164,In_244);
xnor U85 (N_85,In_180,In_13);
or U86 (N_86,In_222,In_260);
or U87 (N_87,In_38,In_124);
or U88 (N_88,In_303,In_424);
xnor U89 (N_89,In_191,In_35);
and U90 (N_90,In_493,In_436);
or U91 (N_91,In_323,In_431);
nand U92 (N_92,In_207,In_183);
nor U93 (N_93,In_428,In_449);
xnor U94 (N_94,In_446,In_353);
or U95 (N_95,In_147,In_306);
or U96 (N_96,In_421,In_210);
xnor U97 (N_97,In_106,In_190);
and U98 (N_98,In_274,In_198);
nor U99 (N_99,In_312,In_130);
or U100 (N_100,In_377,In_39);
or U101 (N_101,In_454,In_451);
and U102 (N_102,In_376,In_41);
nand U103 (N_103,In_226,In_257);
nand U104 (N_104,In_481,In_367);
nor U105 (N_105,In_111,In_53);
and U106 (N_106,In_267,In_358);
nand U107 (N_107,In_204,In_384);
xor U108 (N_108,In_43,In_339);
nor U109 (N_109,In_14,In_79);
nor U110 (N_110,In_118,In_52);
nand U111 (N_111,In_55,In_96);
and U112 (N_112,In_186,In_221);
or U113 (N_113,In_408,In_73);
nand U114 (N_114,In_346,In_125);
and U115 (N_115,In_245,In_336);
nand U116 (N_116,In_189,In_78);
xnor U117 (N_117,In_327,In_253);
nand U118 (N_118,In_15,In_425);
or U119 (N_119,In_170,In_97);
xnor U120 (N_120,In_66,In_275);
nor U121 (N_121,In_402,In_287);
and U122 (N_122,In_46,In_348);
nand U123 (N_123,In_272,In_338);
and U124 (N_124,In_302,In_417);
and U125 (N_125,In_247,In_294);
xnor U126 (N_126,In_197,In_399);
xor U127 (N_127,In_355,In_179);
xor U128 (N_128,In_347,In_223);
or U129 (N_129,In_142,In_70);
nand U130 (N_130,In_95,In_475);
xor U131 (N_131,In_442,In_8);
nand U132 (N_132,In_291,In_18);
and U133 (N_133,In_195,In_72);
or U134 (N_134,In_200,In_304);
nor U135 (N_135,In_182,In_22);
and U136 (N_136,In_342,In_325);
xnor U137 (N_137,In_438,In_150);
and U138 (N_138,In_71,In_322);
xnor U139 (N_139,In_211,In_434);
nand U140 (N_140,In_388,In_439);
and U141 (N_141,In_82,In_492);
nand U142 (N_142,In_284,In_363);
or U143 (N_143,In_468,In_136);
nor U144 (N_144,In_405,In_93);
or U145 (N_145,In_6,In_401);
xor U146 (N_146,In_120,In_465);
xor U147 (N_147,In_135,In_166);
and U148 (N_148,In_154,In_375);
xnor U149 (N_149,In_461,In_288);
xnor U150 (N_150,In_285,In_452);
or U151 (N_151,In_298,In_25);
nand U152 (N_152,In_34,In_235);
xor U153 (N_153,In_119,In_192);
nand U154 (N_154,In_484,In_264);
and U155 (N_155,In_224,In_368);
nor U156 (N_156,In_27,In_308);
xor U157 (N_157,In_467,In_112);
nand U158 (N_158,In_206,In_371);
or U159 (N_159,In_177,In_297);
nor U160 (N_160,In_390,In_254);
nand U161 (N_161,In_33,In_209);
and U162 (N_162,In_239,In_263);
xnor U163 (N_163,In_372,In_132);
and U164 (N_164,In_311,In_185);
xor U165 (N_165,In_354,In_440);
nor U166 (N_166,In_498,In_137);
nand U167 (N_167,In_57,In_374);
nand U168 (N_168,In_48,In_44);
or U169 (N_169,In_499,In_76);
and U170 (N_170,In_496,In_158);
nor U171 (N_171,In_92,In_187);
or U172 (N_172,In_128,In_356);
xor U173 (N_173,In_237,In_242);
nor U174 (N_174,In_448,In_241);
nand U175 (N_175,In_21,In_58);
and U176 (N_176,In_381,In_398);
or U177 (N_177,In_139,In_361);
nor U178 (N_178,In_379,In_151);
nand U179 (N_179,In_40,In_63);
nand U180 (N_180,In_332,In_391);
or U181 (N_181,In_149,In_273);
nor U182 (N_182,In_335,In_419);
xnor U183 (N_183,In_174,In_378);
nor U184 (N_184,In_168,In_422);
xor U185 (N_185,In_282,In_220);
nand U186 (N_186,In_11,In_450);
and U187 (N_187,In_133,In_24);
nor U188 (N_188,In_410,In_296);
nor U189 (N_189,In_281,In_433);
or U190 (N_190,In_23,In_386);
and U191 (N_191,In_248,In_265);
nor U192 (N_192,In_318,In_360);
nor U193 (N_193,In_155,In_101);
and U194 (N_194,In_2,In_362);
xor U195 (N_195,In_478,In_196);
and U196 (N_196,In_225,In_68);
nand U197 (N_197,In_470,In_324);
nand U198 (N_198,In_152,In_393);
nand U199 (N_199,In_1,In_345);
or U200 (N_200,In_117,In_255);
nor U201 (N_201,In_126,In_482);
or U202 (N_202,In_369,In_270);
xnor U203 (N_203,In_184,In_331);
xnor U204 (N_204,In_230,In_62);
and U205 (N_205,In_243,In_427);
xnor U206 (N_206,In_50,In_292);
nand U207 (N_207,In_394,In_397);
xnor U208 (N_208,In_116,In_485);
nand U209 (N_209,In_9,In_319);
nor U210 (N_210,In_321,In_300);
xnor U211 (N_211,In_278,In_10);
nand U212 (N_212,In_64,In_5);
xor U213 (N_213,In_293,In_326);
or U214 (N_214,In_307,In_404);
nor U215 (N_215,In_60,In_47);
nand U216 (N_216,In_217,In_350);
or U217 (N_217,In_432,In_315);
xnor U218 (N_218,In_99,In_134);
nor U219 (N_219,In_17,In_87);
or U220 (N_220,In_143,In_411);
xor U221 (N_221,In_328,In_262);
nor U222 (N_222,In_365,In_412);
nor U223 (N_223,In_456,In_351);
xnor U224 (N_224,In_201,In_486);
nand U225 (N_225,In_453,In_16);
or U226 (N_226,In_122,In_75);
and U227 (N_227,In_146,In_289);
xnor U228 (N_228,In_113,In_88);
and U229 (N_229,In_28,In_383);
xnor U230 (N_230,In_352,In_329);
and U231 (N_231,In_32,In_477);
nand U232 (N_232,In_83,In_407);
and U233 (N_233,In_4,In_370);
nor U234 (N_234,In_54,In_409);
or U235 (N_235,In_162,In_487);
and U236 (N_236,In_234,In_172);
nand U237 (N_237,In_160,In_109);
xnor U238 (N_238,In_491,In_280);
and U239 (N_239,In_213,In_400);
nand U240 (N_240,In_445,In_145);
and U241 (N_241,In_131,In_320);
nor U242 (N_242,In_114,In_349);
or U243 (N_243,In_20,In_458);
nand U244 (N_244,In_176,In_317);
nand U245 (N_245,In_236,In_156);
nand U246 (N_246,In_0,In_333);
or U247 (N_247,In_110,In_205);
and U248 (N_248,In_479,In_218);
and U249 (N_249,In_31,In_373);
or U250 (N_250,In_325,In_321);
and U251 (N_251,In_365,In_162);
xor U252 (N_252,In_25,In_452);
nand U253 (N_253,In_6,In_362);
xnor U254 (N_254,In_370,In_151);
nor U255 (N_255,In_425,In_135);
and U256 (N_256,In_389,In_258);
xor U257 (N_257,In_397,In_203);
nand U258 (N_258,In_419,In_115);
nor U259 (N_259,In_54,In_79);
xnor U260 (N_260,In_464,In_457);
and U261 (N_261,In_122,In_225);
or U262 (N_262,In_488,In_437);
and U263 (N_263,In_186,In_246);
or U264 (N_264,In_490,In_186);
nor U265 (N_265,In_215,In_442);
or U266 (N_266,In_88,In_248);
nand U267 (N_267,In_191,In_204);
nand U268 (N_268,In_464,In_83);
and U269 (N_269,In_438,In_274);
xnor U270 (N_270,In_29,In_333);
or U271 (N_271,In_213,In_269);
nand U272 (N_272,In_7,In_304);
nand U273 (N_273,In_16,In_66);
nor U274 (N_274,In_322,In_257);
nand U275 (N_275,In_300,In_462);
or U276 (N_276,In_204,In_219);
xnor U277 (N_277,In_97,In_370);
nor U278 (N_278,In_322,In_178);
or U279 (N_279,In_46,In_499);
or U280 (N_280,In_417,In_130);
or U281 (N_281,In_348,In_160);
xnor U282 (N_282,In_441,In_74);
xor U283 (N_283,In_498,In_182);
nand U284 (N_284,In_294,In_96);
xnor U285 (N_285,In_437,In_206);
nand U286 (N_286,In_129,In_106);
or U287 (N_287,In_188,In_304);
or U288 (N_288,In_413,In_267);
and U289 (N_289,In_431,In_383);
and U290 (N_290,In_478,In_378);
or U291 (N_291,In_320,In_27);
or U292 (N_292,In_214,In_161);
nand U293 (N_293,In_484,In_327);
nand U294 (N_294,In_453,In_60);
and U295 (N_295,In_118,In_338);
and U296 (N_296,In_82,In_103);
xnor U297 (N_297,In_416,In_12);
or U298 (N_298,In_13,In_126);
nor U299 (N_299,In_120,In_108);
nor U300 (N_300,In_50,In_219);
xor U301 (N_301,In_441,In_254);
nor U302 (N_302,In_167,In_7);
or U303 (N_303,In_12,In_408);
and U304 (N_304,In_4,In_257);
or U305 (N_305,In_18,In_338);
nand U306 (N_306,In_167,In_479);
xnor U307 (N_307,In_335,In_7);
nor U308 (N_308,In_385,In_388);
xnor U309 (N_309,In_404,In_430);
xnor U310 (N_310,In_196,In_171);
nand U311 (N_311,In_245,In_362);
nor U312 (N_312,In_28,In_65);
xnor U313 (N_313,In_369,In_94);
nor U314 (N_314,In_215,In_469);
nor U315 (N_315,In_376,In_440);
or U316 (N_316,In_262,In_173);
or U317 (N_317,In_358,In_343);
nor U318 (N_318,In_340,In_85);
nor U319 (N_319,In_41,In_266);
and U320 (N_320,In_356,In_383);
xnor U321 (N_321,In_56,In_385);
and U322 (N_322,In_221,In_276);
or U323 (N_323,In_248,In_240);
nor U324 (N_324,In_363,In_84);
or U325 (N_325,In_342,In_278);
or U326 (N_326,In_52,In_299);
or U327 (N_327,In_339,In_158);
xor U328 (N_328,In_444,In_99);
or U329 (N_329,In_185,In_47);
and U330 (N_330,In_215,In_294);
nor U331 (N_331,In_8,In_295);
nand U332 (N_332,In_409,In_401);
and U333 (N_333,In_249,In_27);
xor U334 (N_334,In_377,In_92);
xor U335 (N_335,In_213,In_188);
or U336 (N_336,In_487,In_240);
nor U337 (N_337,In_456,In_427);
and U338 (N_338,In_117,In_238);
nand U339 (N_339,In_412,In_149);
or U340 (N_340,In_418,In_486);
nor U341 (N_341,In_252,In_288);
and U342 (N_342,In_64,In_0);
nor U343 (N_343,In_351,In_222);
xnor U344 (N_344,In_319,In_58);
nand U345 (N_345,In_229,In_283);
and U346 (N_346,In_294,In_375);
nor U347 (N_347,In_389,In_290);
and U348 (N_348,In_151,In_29);
and U349 (N_349,In_468,In_350);
nand U350 (N_350,In_283,In_12);
nand U351 (N_351,In_381,In_100);
or U352 (N_352,In_278,In_468);
xor U353 (N_353,In_486,In_346);
xnor U354 (N_354,In_173,In_107);
nand U355 (N_355,In_304,In_86);
or U356 (N_356,In_145,In_376);
xor U357 (N_357,In_243,In_78);
and U358 (N_358,In_400,In_59);
nor U359 (N_359,In_315,In_334);
and U360 (N_360,In_369,In_30);
nor U361 (N_361,In_412,In_357);
and U362 (N_362,In_29,In_110);
and U363 (N_363,In_365,In_311);
or U364 (N_364,In_12,In_245);
or U365 (N_365,In_146,In_203);
and U366 (N_366,In_464,In_9);
nand U367 (N_367,In_6,In_398);
nor U368 (N_368,In_91,In_472);
and U369 (N_369,In_36,In_464);
nor U370 (N_370,In_42,In_350);
nor U371 (N_371,In_28,In_314);
nand U372 (N_372,In_221,In_499);
or U373 (N_373,In_184,In_123);
nor U374 (N_374,In_405,In_445);
or U375 (N_375,In_218,In_463);
and U376 (N_376,In_89,In_159);
nand U377 (N_377,In_231,In_387);
xor U378 (N_378,In_220,In_252);
or U379 (N_379,In_395,In_193);
xnor U380 (N_380,In_390,In_468);
nand U381 (N_381,In_479,In_493);
or U382 (N_382,In_107,In_335);
nand U383 (N_383,In_9,In_372);
nor U384 (N_384,In_323,In_499);
or U385 (N_385,In_385,In_322);
or U386 (N_386,In_278,In_133);
xnor U387 (N_387,In_153,In_131);
xor U388 (N_388,In_321,In_269);
or U389 (N_389,In_180,In_285);
or U390 (N_390,In_23,In_65);
or U391 (N_391,In_188,In_11);
nor U392 (N_392,In_31,In_365);
or U393 (N_393,In_395,In_239);
nand U394 (N_394,In_274,In_384);
and U395 (N_395,In_355,In_478);
nor U396 (N_396,In_335,In_79);
xnor U397 (N_397,In_27,In_6);
or U398 (N_398,In_343,In_320);
xor U399 (N_399,In_491,In_399);
nor U400 (N_400,In_163,In_149);
and U401 (N_401,In_255,In_308);
and U402 (N_402,In_161,In_370);
nor U403 (N_403,In_150,In_221);
xnor U404 (N_404,In_101,In_486);
nor U405 (N_405,In_390,In_421);
or U406 (N_406,In_471,In_349);
xnor U407 (N_407,In_386,In_170);
xnor U408 (N_408,In_96,In_236);
nand U409 (N_409,In_400,In_311);
and U410 (N_410,In_229,In_108);
xor U411 (N_411,In_261,In_276);
nor U412 (N_412,In_446,In_61);
nor U413 (N_413,In_345,In_353);
nand U414 (N_414,In_319,In_482);
nor U415 (N_415,In_306,In_180);
nor U416 (N_416,In_303,In_91);
nor U417 (N_417,In_364,In_268);
or U418 (N_418,In_342,In_35);
or U419 (N_419,In_311,In_377);
nor U420 (N_420,In_290,In_315);
xor U421 (N_421,In_115,In_72);
xnor U422 (N_422,In_80,In_114);
or U423 (N_423,In_235,In_28);
or U424 (N_424,In_323,In_24);
nor U425 (N_425,In_412,In_21);
and U426 (N_426,In_44,In_496);
or U427 (N_427,In_414,In_222);
xnor U428 (N_428,In_387,In_94);
nand U429 (N_429,In_431,In_185);
xnor U430 (N_430,In_27,In_86);
and U431 (N_431,In_131,In_56);
nand U432 (N_432,In_290,In_464);
nand U433 (N_433,In_385,In_345);
nor U434 (N_434,In_162,In_363);
xnor U435 (N_435,In_405,In_321);
or U436 (N_436,In_105,In_385);
nor U437 (N_437,In_73,In_289);
or U438 (N_438,In_77,In_22);
xor U439 (N_439,In_183,In_25);
or U440 (N_440,In_83,In_33);
or U441 (N_441,In_321,In_100);
nor U442 (N_442,In_254,In_375);
nor U443 (N_443,In_204,In_88);
nor U444 (N_444,In_226,In_459);
nand U445 (N_445,In_185,In_352);
nand U446 (N_446,In_385,In_257);
or U447 (N_447,In_139,In_331);
nand U448 (N_448,In_142,In_211);
nand U449 (N_449,In_248,In_66);
nand U450 (N_450,In_218,In_106);
or U451 (N_451,In_382,In_428);
nor U452 (N_452,In_447,In_205);
and U453 (N_453,In_273,In_181);
xnor U454 (N_454,In_422,In_62);
nand U455 (N_455,In_374,In_265);
or U456 (N_456,In_341,In_277);
nor U457 (N_457,In_286,In_81);
or U458 (N_458,In_246,In_340);
or U459 (N_459,In_253,In_122);
xor U460 (N_460,In_142,In_499);
nand U461 (N_461,In_130,In_346);
nor U462 (N_462,In_220,In_204);
nor U463 (N_463,In_472,In_467);
and U464 (N_464,In_64,In_59);
or U465 (N_465,In_185,In_221);
nor U466 (N_466,In_164,In_127);
nor U467 (N_467,In_361,In_352);
and U468 (N_468,In_240,In_375);
nor U469 (N_469,In_34,In_264);
nor U470 (N_470,In_363,In_64);
nor U471 (N_471,In_234,In_223);
and U472 (N_472,In_490,In_389);
or U473 (N_473,In_58,In_472);
or U474 (N_474,In_143,In_409);
or U475 (N_475,In_271,In_343);
nand U476 (N_476,In_316,In_28);
nor U477 (N_477,In_29,In_215);
and U478 (N_478,In_103,In_260);
xnor U479 (N_479,In_272,In_427);
nand U480 (N_480,In_93,In_415);
nand U481 (N_481,In_356,In_418);
and U482 (N_482,In_36,In_277);
nor U483 (N_483,In_270,In_469);
xor U484 (N_484,In_60,In_50);
and U485 (N_485,In_419,In_62);
nand U486 (N_486,In_423,In_222);
xnor U487 (N_487,In_409,In_309);
and U488 (N_488,In_270,In_454);
and U489 (N_489,In_479,In_499);
xor U490 (N_490,In_329,In_222);
nor U491 (N_491,In_343,In_110);
and U492 (N_492,In_251,In_128);
and U493 (N_493,In_183,In_140);
xnor U494 (N_494,In_55,In_12);
or U495 (N_495,In_440,In_339);
or U496 (N_496,In_387,In_279);
or U497 (N_497,In_301,In_258);
and U498 (N_498,In_287,In_313);
xnor U499 (N_499,In_238,In_69);
or U500 (N_500,In_435,In_231);
nand U501 (N_501,In_405,In_439);
xor U502 (N_502,In_207,In_458);
nor U503 (N_503,In_10,In_232);
or U504 (N_504,In_328,In_51);
nor U505 (N_505,In_334,In_269);
xor U506 (N_506,In_29,In_452);
nand U507 (N_507,In_136,In_146);
xor U508 (N_508,In_410,In_231);
xnor U509 (N_509,In_14,In_289);
xor U510 (N_510,In_58,In_369);
nand U511 (N_511,In_269,In_70);
xnor U512 (N_512,In_312,In_374);
xor U513 (N_513,In_36,In_418);
nand U514 (N_514,In_373,In_375);
xnor U515 (N_515,In_315,In_141);
or U516 (N_516,In_344,In_320);
nor U517 (N_517,In_7,In_254);
or U518 (N_518,In_119,In_36);
or U519 (N_519,In_416,In_3);
nor U520 (N_520,In_23,In_396);
xnor U521 (N_521,In_81,In_453);
xnor U522 (N_522,In_375,In_419);
nand U523 (N_523,In_271,In_232);
nand U524 (N_524,In_198,In_440);
nand U525 (N_525,In_187,In_250);
or U526 (N_526,In_260,In_214);
xnor U527 (N_527,In_112,In_174);
xnor U528 (N_528,In_393,In_173);
or U529 (N_529,In_416,In_152);
nand U530 (N_530,In_417,In_40);
and U531 (N_531,In_51,In_401);
and U532 (N_532,In_432,In_240);
xnor U533 (N_533,In_377,In_492);
nand U534 (N_534,In_113,In_59);
nor U535 (N_535,In_227,In_36);
and U536 (N_536,In_116,In_498);
nand U537 (N_537,In_304,In_112);
and U538 (N_538,In_416,In_460);
or U539 (N_539,In_357,In_338);
and U540 (N_540,In_63,In_473);
nor U541 (N_541,In_266,In_212);
or U542 (N_542,In_247,In_357);
nand U543 (N_543,In_216,In_7);
and U544 (N_544,In_367,In_51);
nand U545 (N_545,In_426,In_17);
and U546 (N_546,In_179,In_307);
or U547 (N_547,In_158,In_340);
xnor U548 (N_548,In_8,In_269);
xnor U549 (N_549,In_477,In_175);
and U550 (N_550,In_93,In_286);
nand U551 (N_551,In_263,In_324);
and U552 (N_552,In_49,In_254);
nor U553 (N_553,In_146,In_470);
xnor U554 (N_554,In_435,In_278);
xnor U555 (N_555,In_476,In_347);
and U556 (N_556,In_315,In_442);
nand U557 (N_557,In_3,In_205);
and U558 (N_558,In_429,In_323);
nor U559 (N_559,In_383,In_433);
nor U560 (N_560,In_359,In_297);
nor U561 (N_561,In_294,In_372);
nand U562 (N_562,In_18,In_98);
or U563 (N_563,In_238,In_138);
nand U564 (N_564,In_236,In_356);
and U565 (N_565,In_490,In_354);
xnor U566 (N_566,In_18,In_41);
and U567 (N_567,In_195,In_170);
nor U568 (N_568,In_256,In_65);
or U569 (N_569,In_129,In_339);
xnor U570 (N_570,In_499,In_136);
xor U571 (N_571,In_143,In_158);
nor U572 (N_572,In_158,In_200);
and U573 (N_573,In_55,In_459);
xnor U574 (N_574,In_443,In_377);
or U575 (N_575,In_157,In_134);
and U576 (N_576,In_458,In_253);
or U577 (N_577,In_329,In_494);
xnor U578 (N_578,In_276,In_206);
nand U579 (N_579,In_387,In_436);
xor U580 (N_580,In_176,In_415);
or U581 (N_581,In_139,In_11);
xor U582 (N_582,In_498,In_456);
nor U583 (N_583,In_456,In_258);
and U584 (N_584,In_137,In_82);
nand U585 (N_585,In_174,In_114);
nand U586 (N_586,In_327,In_264);
and U587 (N_587,In_232,In_293);
nor U588 (N_588,In_226,In_162);
xor U589 (N_589,In_87,In_165);
or U590 (N_590,In_86,In_281);
or U591 (N_591,In_290,In_60);
or U592 (N_592,In_142,In_350);
and U593 (N_593,In_30,In_378);
nor U594 (N_594,In_436,In_466);
or U595 (N_595,In_172,In_283);
xor U596 (N_596,In_456,In_288);
xnor U597 (N_597,In_77,In_280);
or U598 (N_598,In_415,In_139);
nor U599 (N_599,In_496,In_294);
nor U600 (N_600,N_424,N_209);
and U601 (N_601,N_237,N_488);
or U602 (N_602,N_293,N_289);
or U603 (N_603,N_321,N_21);
or U604 (N_604,N_287,N_368);
xnor U605 (N_605,N_579,N_25);
nand U606 (N_606,N_60,N_67);
or U607 (N_607,N_81,N_345);
nand U608 (N_608,N_296,N_212);
nor U609 (N_609,N_537,N_340);
nor U610 (N_610,N_421,N_17);
nand U611 (N_611,N_46,N_255);
or U612 (N_612,N_335,N_78);
nor U613 (N_613,N_360,N_250);
or U614 (N_614,N_74,N_247);
or U615 (N_615,N_544,N_466);
or U616 (N_616,N_549,N_158);
xor U617 (N_617,N_526,N_408);
nand U618 (N_618,N_556,N_199);
or U619 (N_619,N_571,N_348);
nand U620 (N_620,N_410,N_225);
nor U621 (N_621,N_532,N_282);
xnor U622 (N_622,N_319,N_135);
or U623 (N_623,N_505,N_290);
xor U624 (N_624,N_73,N_206);
nor U625 (N_625,N_361,N_437);
xnor U626 (N_626,N_351,N_198);
or U627 (N_627,N_477,N_307);
nand U628 (N_628,N_99,N_308);
nor U629 (N_629,N_381,N_175);
nor U630 (N_630,N_582,N_66);
nand U631 (N_631,N_275,N_405);
xor U632 (N_632,N_43,N_414);
and U633 (N_633,N_333,N_353);
or U634 (N_634,N_301,N_504);
nand U635 (N_635,N_40,N_513);
nand U636 (N_636,N_173,N_597);
or U637 (N_637,N_11,N_427);
xor U638 (N_638,N_285,N_502);
or U639 (N_639,N_178,N_129);
xor U640 (N_640,N_476,N_33);
or U641 (N_641,N_469,N_363);
xnor U642 (N_642,N_27,N_591);
or U643 (N_643,N_403,N_387);
nor U644 (N_644,N_177,N_569);
xnor U645 (N_645,N_208,N_318);
xnor U646 (N_646,N_281,N_525);
xor U647 (N_647,N_13,N_251);
nor U648 (N_648,N_134,N_415);
nor U649 (N_649,N_231,N_136);
or U650 (N_650,N_113,N_510);
and U651 (N_651,N_214,N_184);
and U652 (N_652,N_352,N_283);
and U653 (N_653,N_234,N_367);
nor U654 (N_654,N_35,N_356);
nand U655 (N_655,N_261,N_48);
nor U656 (N_656,N_191,N_259);
and U657 (N_657,N_546,N_151);
nor U658 (N_658,N_131,N_270);
xor U659 (N_659,N_436,N_118);
and U660 (N_660,N_244,N_14);
xor U661 (N_661,N_75,N_535);
or U662 (N_662,N_79,N_145);
and U663 (N_663,N_369,N_143);
or U664 (N_664,N_64,N_599);
nor U665 (N_665,N_419,N_82);
xnor U666 (N_666,N_432,N_305);
xor U667 (N_667,N_164,N_18);
nor U668 (N_668,N_383,N_106);
nor U669 (N_669,N_380,N_71);
nor U670 (N_670,N_552,N_426);
xnor U671 (N_671,N_550,N_501);
nand U672 (N_672,N_105,N_323);
nand U673 (N_673,N_30,N_422);
or U674 (N_674,N_562,N_389);
nand U675 (N_675,N_377,N_76);
or U676 (N_676,N_534,N_574);
nand U677 (N_677,N_386,N_51);
or U678 (N_678,N_317,N_563);
nand U679 (N_679,N_311,N_447);
nor U680 (N_680,N_218,N_215);
and U681 (N_681,N_420,N_481);
xnor U682 (N_682,N_5,N_109);
xor U683 (N_683,N_338,N_37);
and U684 (N_684,N_529,N_220);
nand U685 (N_685,N_428,N_245);
nand U686 (N_686,N_34,N_107);
nand U687 (N_687,N_96,N_418);
or U688 (N_688,N_385,N_0);
xor U689 (N_689,N_401,N_486);
nor U690 (N_690,N_61,N_464);
nand U691 (N_691,N_475,N_190);
xnor U692 (N_692,N_503,N_174);
or U693 (N_693,N_104,N_97);
nor U694 (N_694,N_50,N_112);
xnor U695 (N_695,N_86,N_366);
and U696 (N_696,N_578,N_47);
xor U697 (N_697,N_445,N_595);
and U698 (N_698,N_266,N_23);
or U699 (N_699,N_110,N_400);
nand U700 (N_700,N_442,N_413);
nand U701 (N_701,N_519,N_489);
xnor U702 (N_702,N_253,N_547);
or U703 (N_703,N_520,N_384);
or U704 (N_704,N_458,N_396);
or U705 (N_705,N_327,N_358);
nor U706 (N_706,N_233,N_269);
xnor U707 (N_707,N_416,N_391);
xor U708 (N_708,N_194,N_376);
and U709 (N_709,N_496,N_350);
nor U710 (N_710,N_453,N_431);
nand U711 (N_711,N_395,N_298);
and U712 (N_712,N_465,N_197);
or U713 (N_713,N_31,N_334);
xnor U714 (N_714,N_555,N_241);
and U715 (N_715,N_449,N_373);
nand U716 (N_716,N_506,N_146);
nor U717 (N_717,N_8,N_258);
or U718 (N_718,N_111,N_68);
or U719 (N_719,N_375,N_156);
nand U720 (N_720,N_201,N_583);
and U721 (N_721,N_125,N_238);
and U722 (N_722,N_339,N_117);
or U723 (N_723,N_541,N_203);
nor U724 (N_724,N_515,N_273);
nand U725 (N_725,N_101,N_313);
and U726 (N_726,N_183,N_320);
nand U727 (N_727,N_277,N_62);
xnor U728 (N_728,N_159,N_172);
xor U729 (N_729,N_256,N_130);
and U730 (N_730,N_217,N_39);
and U731 (N_731,N_236,N_148);
nand U732 (N_732,N_157,N_192);
or U733 (N_733,N_397,N_56);
nand U734 (N_734,N_355,N_402);
or U735 (N_735,N_326,N_240);
and U736 (N_736,N_474,N_349);
and U737 (N_737,N_324,N_160);
nand U738 (N_738,N_412,N_58);
nor U739 (N_739,N_278,N_28);
nand U740 (N_740,N_411,N_171);
xnor U741 (N_741,N_216,N_128);
and U742 (N_742,N_357,N_429);
or U743 (N_743,N_235,N_140);
or U744 (N_744,N_10,N_227);
xnor U745 (N_745,N_226,N_155);
and U746 (N_746,N_388,N_138);
or U747 (N_747,N_57,N_124);
or U748 (N_748,N_181,N_16);
or U749 (N_749,N_557,N_119);
and U750 (N_750,N_297,N_254);
or U751 (N_751,N_438,N_538);
and U752 (N_752,N_570,N_589);
nand U753 (N_753,N_492,N_470);
nor U754 (N_754,N_480,N_167);
nor U755 (N_755,N_100,N_598);
xnor U756 (N_756,N_263,N_268);
and U757 (N_757,N_430,N_116);
and U758 (N_758,N_139,N_439);
and U759 (N_759,N_149,N_249);
and U760 (N_760,N_499,N_560);
nand U761 (N_761,N_186,N_205);
nand U762 (N_762,N_500,N_302);
and U763 (N_763,N_77,N_221);
and U764 (N_764,N_200,N_122);
xnor U765 (N_765,N_179,N_398);
nand U766 (N_766,N_463,N_284);
nor U767 (N_767,N_312,N_487);
nor U768 (N_768,N_374,N_596);
and U769 (N_769,N_90,N_126);
xnor U770 (N_770,N_123,N_455);
and U771 (N_771,N_141,N_581);
or U772 (N_772,N_72,N_288);
or U773 (N_773,N_94,N_276);
nand U774 (N_774,N_166,N_342);
and U775 (N_775,N_267,N_102);
nand U776 (N_776,N_440,N_142);
nand U777 (N_777,N_92,N_461);
nand U778 (N_778,N_390,N_185);
xnor U779 (N_779,N_91,N_147);
or U780 (N_780,N_451,N_204);
or U781 (N_781,N_45,N_272);
xor U782 (N_782,N_232,N_70);
and U783 (N_783,N_531,N_63);
xor U784 (N_784,N_450,N_44);
or U785 (N_785,N_262,N_89);
nor U786 (N_786,N_354,N_587);
and U787 (N_787,N_572,N_425);
nor U788 (N_788,N_26,N_95);
nor U789 (N_789,N_310,N_180);
and U790 (N_790,N_478,N_32);
nand U791 (N_791,N_84,N_392);
or U792 (N_792,N_163,N_378);
and U793 (N_793,N_576,N_545);
nor U794 (N_794,N_210,N_260);
nand U795 (N_795,N_444,N_341);
nor U796 (N_796,N_566,N_80);
nor U797 (N_797,N_271,N_170);
nand U798 (N_798,N_264,N_512);
and U799 (N_799,N_379,N_228);
nor U800 (N_800,N_36,N_115);
nor U801 (N_801,N_359,N_536);
or U802 (N_802,N_29,N_554);
nand U803 (N_803,N_55,N_304);
or U804 (N_804,N_362,N_239);
nand U805 (N_805,N_484,N_20);
and U806 (N_806,N_332,N_306);
nand U807 (N_807,N_471,N_495);
and U808 (N_808,N_417,N_559);
nor U809 (N_809,N_548,N_452);
and U810 (N_810,N_460,N_328);
xnor U811 (N_811,N_230,N_514);
and U812 (N_812,N_539,N_528);
and U813 (N_813,N_229,N_573);
or U814 (N_814,N_182,N_144);
and U815 (N_815,N_482,N_193);
and U816 (N_816,N_586,N_219);
nand U817 (N_817,N_24,N_564);
or U818 (N_818,N_542,N_543);
nor U819 (N_819,N_409,N_567);
nor U820 (N_820,N_364,N_473);
and U821 (N_821,N_522,N_114);
nand U822 (N_822,N_511,N_83);
or U823 (N_823,N_490,N_279);
and U824 (N_824,N_207,N_551);
nor U825 (N_825,N_524,N_292);
or U826 (N_826,N_423,N_568);
nand U827 (N_827,N_472,N_406);
nor U828 (N_828,N_133,N_347);
or U829 (N_829,N_88,N_223);
nand U830 (N_830,N_314,N_331);
nand U831 (N_831,N_343,N_9);
nand U832 (N_832,N_483,N_590);
and U833 (N_833,N_517,N_322);
and U834 (N_834,N_592,N_516);
and U835 (N_835,N_467,N_493);
nor U836 (N_836,N_103,N_3);
xor U837 (N_837,N_300,N_577);
or U838 (N_838,N_42,N_161);
nor U839 (N_839,N_213,N_195);
and U840 (N_840,N_188,N_315);
xor U841 (N_841,N_365,N_252);
nand U842 (N_842,N_165,N_457);
or U843 (N_843,N_22,N_433);
and U844 (N_844,N_523,N_176);
nand U845 (N_845,N_152,N_530);
xor U846 (N_846,N_580,N_265);
nand U847 (N_847,N_98,N_533);
or U848 (N_848,N_54,N_382);
nor U849 (N_849,N_187,N_150);
nand U850 (N_850,N_69,N_393);
and U851 (N_851,N_127,N_132);
or U852 (N_852,N_407,N_462);
and U853 (N_853,N_448,N_459);
and U854 (N_854,N_337,N_4);
nand U855 (N_855,N_370,N_85);
or U856 (N_856,N_49,N_19);
xor U857 (N_857,N_575,N_168);
nand U858 (N_858,N_120,N_291);
nand U859 (N_859,N_479,N_154);
nand U860 (N_860,N_169,N_53);
nand U861 (N_861,N_41,N_257);
nor U862 (N_862,N_468,N_242);
and U863 (N_863,N_196,N_372);
xnor U864 (N_864,N_446,N_336);
and U865 (N_865,N_246,N_434);
nor U866 (N_866,N_508,N_594);
xor U867 (N_867,N_121,N_498);
and U868 (N_868,N_299,N_137);
or U869 (N_869,N_303,N_202);
nor U870 (N_870,N_509,N_189);
or U871 (N_871,N_280,N_224);
nand U872 (N_872,N_65,N_243);
nor U873 (N_873,N_584,N_399);
nand U874 (N_874,N_325,N_561);
nor U875 (N_875,N_248,N_52);
nor U876 (N_876,N_456,N_565);
and U877 (N_877,N_316,N_346);
nand U878 (N_878,N_404,N_309);
and U879 (N_879,N_435,N_344);
or U880 (N_880,N_211,N_162);
and U881 (N_881,N_286,N_443);
and U882 (N_882,N_108,N_87);
nor U883 (N_883,N_518,N_494);
nor U884 (N_884,N_294,N_497);
or U885 (N_885,N_222,N_15);
or U886 (N_886,N_274,N_330);
and U887 (N_887,N_593,N_521);
nand U888 (N_888,N_153,N_59);
and U889 (N_889,N_507,N_585);
nand U890 (N_890,N_7,N_329);
nand U891 (N_891,N_553,N_12);
xor U892 (N_892,N_2,N_93);
and U893 (N_893,N_38,N_491);
nand U894 (N_894,N_295,N_540);
and U895 (N_895,N_394,N_441);
and U896 (N_896,N_6,N_588);
nor U897 (N_897,N_371,N_454);
xnor U898 (N_898,N_1,N_558);
xnor U899 (N_899,N_485,N_527);
and U900 (N_900,N_139,N_59);
and U901 (N_901,N_405,N_98);
and U902 (N_902,N_202,N_264);
or U903 (N_903,N_47,N_151);
nor U904 (N_904,N_121,N_39);
nor U905 (N_905,N_49,N_582);
xor U906 (N_906,N_34,N_215);
nor U907 (N_907,N_450,N_552);
nor U908 (N_908,N_136,N_79);
nand U909 (N_909,N_20,N_100);
nor U910 (N_910,N_437,N_405);
nand U911 (N_911,N_356,N_539);
nand U912 (N_912,N_245,N_442);
nor U913 (N_913,N_247,N_262);
nand U914 (N_914,N_278,N_261);
or U915 (N_915,N_269,N_76);
and U916 (N_916,N_33,N_507);
nor U917 (N_917,N_532,N_285);
nor U918 (N_918,N_75,N_239);
or U919 (N_919,N_358,N_411);
or U920 (N_920,N_333,N_433);
nand U921 (N_921,N_389,N_319);
or U922 (N_922,N_471,N_127);
nand U923 (N_923,N_587,N_385);
or U924 (N_924,N_257,N_84);
nor U925 (N_925,N_226,N_70);
nand U926 (N_926,N_321,N_83);
nor U927 (N_927,N_389,N_175);
nand U928 (N_928,N_513,N_441);
nor U929 (N_929,N_204,N_96);
xnor U930 (N_930,N_184,N_580);
and U931 (N_931,N_75,N_340);
and U932 (N_932,N_437,N_445);
or U933 (N_933,N_236,N_200);
nand U934 (N_934,N_344,N_347);
and U935 (N_935,N_138,N_73);
nor U936 (N_936,N_353,N_514);
nor U937 (N_937,N_297,N_463);
xnor U938 (N_938,N_227,N_257);
xor U939 (N_939,N_155,N_65);
xor U940 (N_940,N_560,N_485);
nand U941 (N_941,N_561,N_48);
nor U942 (N_942,N_172,N_36);
nor U943 (N_943,N_503,N_562);
nand U944 (N_944,N_127,N_325);
or U945 (N_945,N_353,N_289);
nor U946 (N_946,N_396,N_275);
and U947 (N_947,N_311,N_172);
xnor U948 (N_948,N_267,N_293);
nor U949 (N_949,N_327,N_234);
nor U950 (N_950,N_340,N_213);
and U951 (N_951,N_269,N_573);
or U952 (N_952,N_292,N_548);
nor U953 (N_953,N_147,N_278);
nor U954 (N_954,N_571,N_507);
and U955 (N_955,N_336,N_202);
xnor U956 (N_956,N_431,N_162);
and U957 (N_957,N_79,N_478);
nor U958 (N_958,N_530,N_506);
or U959 (N_959,N_312,N_209);
and U960 (N_960,N_499,N_242);
and U961 (N_961,N_404,N_439);
and U962 (N_962,N_487,N_185);
or U963 (N_963,N_464,N_356);
xnor U964 (N_964,N_568,N_41);
and U965 (N_965,N_404,N_455);
nand U966 (N_966,N_199,N_414);
and U967 (N_967,N_562,N_462);
xnor U968 (N_968,N_122,N_249);
or U969 (N_969,N_139,N_588);
nor U970 (N_970,N_577,N_271);
xnor U971 (N_971,N_494,N_493);
nand U972 (N_972,N_544,N_47);
and U973 (N_973,N_510,N_508);
or U974 (N_974,N_132,N_551);
nand U975 (N_975,N_548,N_88);
nand U976 (N_976,N_160,N_290);
nand U977 (N_977,N_510,N_213);
nand U978 (N_978,N_345,N_34);
nor U979 (N_979,N_174,N_540);
nand U980 (N_980,N_234,N_575);
nand U981 (N_981,N_393,N_129);
nor U982 (N_982,N_598,N_433);
xnor U983 (N_983,N_410,N_194);
xor U984 (N_984,N_580,N_130);
and U985 (N_985,N_271,N_86);
nor U986 (N_986,N_239,N_126);
or U987 (N_987,N_377,N_300);
nor U988 (N_988,N_306,N_120);
nor U989 (N_989,N_308,N_517);
nor U990 (N_990,N_403,N_473);
nand U991 (N_991,N_234,N_7);
and U992 (N_992,N_319,N_56);
nor U993 (N_993,N_481,N_304);
and U994 (N_994,N_292,N_212);
nand U995 (N_995,N_439,N_328);
or U996 (N_996,N_192,N_435);
nor U997 (N_997,N_449,N_224);
nor U998 (N_998,N_555,N_443);
nor U999 (N_999,N_192,N_387);
nor U1000 (N_1000,N_236,N_312);
xnor U1001 (N_1001,N_66,N_31);
or U1002 (N_1002,N_380,N_0);
and U1003 (N_1003,N_262,N_370);
nand U1004 (N_1004,N_164,N_369);
and U1005 (N_1005,N_328,N_501);
nand U1006 (N_1006,N_322,N_186);
or U1007 (N_1007,N_176,N_490);
or U1008 (N_1008,N_39,N_114);
and U1009 (N_1009,N_183,N_421);
nor U1010 (N_1010,N_146,N_315);
nand U1011 (N_1011,N_503,N_205);
nand U1012 (N_1012,N_241,N_592);
or U1013 (N_1013,N_297,N_32);
nor U1014 (N_1014,N_567,N_213);
and U1015 (N_1015,N_88,N_396);
or U1016 (N_1016,N_390,N_531);
and U1017 (N_1017,N_567,N_476);
nor U1018 (N_1018,N_179,N_81);
nor U1019 (N_1019,N_545,N_0);
nor U1020 (N_1020,N_228,N_444);
nor U1021 (N_1021,N_535,N_70);
nor U1022 (N_1022,N_277,N_368);
xnor U1023 (N_1023,N_563,N_467);
and U1024 (N_1024,N_477,N_550);
nand U1025 (N_1025,N_181,N_74);
and U1026 (N_1026,N_474,N_141);
and U1027 (N_1027,N_339,N_366);
nor U1028 (N_1028,N_272,N_490);
or U1029 (N_1029,N_47,N_166);
and U1030 (N_1030,N_38,N_533);
or U1031 (N_1031,N_319,N_274);
xnor U1032 (N_1032,N_561,N_544);
nor U1033 (N_1033,N_373,N_52);
or U1034 (N_1034,N_426,N_440);
xnor U1035 (N_1035,N_238,N_279);
xnor U1036 (N_1036,N_40,N_506);
xor U1037 (N_1037,N_548,N_445);
or U1038 (N_1038,N_499,N_320);
nor U1039 (N_1039,N_386,N_82);
nor U1040 (N_1040,N_47,N_263);
nor U1041 (N_1041,N_158,N_424);
xor U1042 (N_1042,N_207,N_424);
and U1043 (N_1043,N_230,N_196);
nand U1044 (N_1044,N_120,N_222);
nand U1045 (N_1045,N_74,N_142);
xor U1046 (N_1046,N_176,N_21);
and U1047 (N_1047,N_54,N_215);
or U1048 (N_1048,N_379,N_443);
nand U1049 (N_1049,N_391,N_406);
nor U1050 (N_1050,N_394,N_208);
xor U1051 (N_1051,N_212,N_295);
nand U1052 (N_1052,N_142,N_73);
nor U1053 (N_1053,N_275,N_348);
nand U1054 (N_1054,N_296,N_298);
or U1055 (N_1055,N_16,N_226);
nor U1056 (N_1056,N_542,N_283);
and U1057 (N_1057,N_393,N_450);
nand U1058 (N_1058,N_424,N_211);
nand U1059 (N_1059,N_297,N_17);
xor U1060 (N_1060,N_401,N_150);
xnor U1061 (N_1061,N_160,N_491);
or U1062 (N_1062,N_326,N_536);
or U1063 (N_1063,N_49,N_24);
xor U1064 (N_1064,N_526,N_302);
or U1065 (N_1065,N_421,N_141);
nand U1066 (N_1066,N_513,N_161);
or U1067 (N_1067,N_393,N_324);
or U1068 (N_1068,N_101,N_370);
xor U1069 (N_1069,N_288,N_146);
and U1070 (N_1070,N_378,N_176);
nand U1071 (N_1071,N_372,N_38);
nor U1072 (N_1072,N_485,N_595);
or U1073 (N_1073,N_214,N_220);
nand U1074 (N_1074,N_190,N_508);
nor U1075 (N_1075,N_220,N_204);
or U1076 (N_1076,N_558,N_215);
or U1077 (N_1077,N_253,N_239);
xor U1078 (N_1078,N_517,N_154);
and U1079 (N_1079,N_41,N_180);
nand U1080 (N_1080,N_234,N_473);
xor U1081 (N_1081,N_268,N_577);
or U1082 (N_1082,N_114,N_52);
xor U1083 (N_1083,N_518,N_125);
nor U1084 (N_1084,N_425,N_406);
nand U1085 (N_1085,N_0,N_156);
nor U1086 (N_1086,N_457,N_598);
xnor U1087 (N_1087,N_98,N_473);
nor U1088 (N_1088,N_359,N_24);
or U1089 (N_1089,N_319,N_377);
nor U1090 (N_1090,N_23,N_539);
and U1091 (N_1091,N_195,N_164);
nor U1092 (N_1092,N_405,N_203);
xor U1093 (N_1093,N_73,N_63);
and U1094 (N_1094,N_430,N_362);
xnor U1095 (N_1095,N_517,N_597);
and U1096 (N_1096,N_304,N_296);
nand U1097 (N_1097,N_276,N_223);
nor U1098 (N_1098,N_549,N_13);
or U1099 (N_1099,N_447,N_322);
nor U1100 (N_1100,N_53,N_8);
nand U1101 (N_1101,N_537,N_567);
xor U1102 (N_1102,N_423,N_25);
nor U1103 (N_1103,N_253,N_446);
xor U1104 (N_1104,N_487,N_222);
xor U1105 (N_1105,N_511,N_473);
and U1106 (N_1106,N_325,N_489);
nor U1107 (N_1107,N_474,N_566);
nand U1108 (N_1108,N_148,N_566);
nor U1109 (N_1109,N_436,N_202);
xor U1110 (N_1110,N_508,N_188);
and U1111 (N_1111,N_13,N_41);
and U1112 (N_1112,N_219,N_92);
or U1113 (N_1113,N_583,N_460);
or U1114 (N_1114,N_219,N_400);
and U1115 (N_1115,N_228,N_504);
nor U1116 (N_1116,N_439,N_590);
and U1117 (N_1117,N_92,N_196);
or U1118 (N_1118,N_5,N_49);
nand U1119 (N_1119,N_18,N_244);
nor U1120 (N_1120,N_268,N_369);
nand U1121 (N_1121,N_230,N_537);
and U1122 (N_1122,N_134,N_264);
nand U1123 (N_1123,N_159,N_590);
or U1124 (N_1124,N_371,N_222);
and U1125 (N_1125,N_549,N_246);
and U1126 (N_1126,N_323,N_559);
nand U1127 (N_1127,N_435,N_333);
nor U1128 (N_1128,N_120,N_207);
nor U1129 (N_1129,N_102,N_402);
or U1130 (N_1130,N_361,N_307);
or U1131 (N_1131,N_166,N_505);
or U1132 (N_1132,N_45,N_110);
or U1133 (N_1133,N_116,N_242);
and U1134 (N_1134,N_352,N_113);
and U1135 (N_1135,N_391,N_190);
or U1136 (N_1136,N_571,N_238);
xnor U1137 (N_1137,N_385,N_458);
or U1138 (N_1138,N_492,N_519);
nand U1139 (N_1139,N_131,N_383);
and U1140 (N_1140,N_205,N_258);
nand U1141 (N_1141,N_55,N_562);
nand U1142 (N_1142,N_446,N_425);
nor U1143 (N_1143,N_211,N_58);
and U1144 (N_1144,N_169,N_286);
xor U1145 (N_1145,N_511,N_328);
and U1146 (N_1146,N_469,N_548);
and U1147 (N_1147,N_238,N_84);
nand U1148 (N_1148,N_472,N_273);
nor U1149 (N_1149,N_339,N_107);
nand U1150 (N_1150,N_259,N_79);
and U1151 (N_1151,N_247,N_449);
xnor U1152 (N_1152,N_167,N_171);
xnor U1153 (N_1153,N_222,N_175);
xor U1154 (N_1154,N_537,N_108);
nor U1155 (N_1155,N_366,N_408);
nor U1156 (N_1156,N_235,N_276);
nand U1157 (N_1157,N_485,N_186);
nor U1158 (N_1158,N_189,N_476);
nor U1159 (N_1159,N_420,N_586);
and U1160 (N_1160,N_176,N_263);
and U1161 (N_1161,N_584,N_234);
or U1162 (N_1162,N_104,N_99);
and U1163 (N_1163,N_565,N_102);
or U1164 (N_1164,N_58,N_481);
nand U1165 (N_1165,N_37,N_376);
nand U1166 (N_1166,N_590,N_230);
nand U1167 (N_1167,N_47,N_528);
xnor U1168 (N_1168,N_485,N_559);
and U1169 (N_1169,N_332,N_447);
or U1170 (N_1170,N_567,N_19);
xnor U1171 (N_1171,N_221,N_223);
or U1172 (N_1172,N_165,N_131);
and U1173 (N_1173,N_394,N_312);
nor U1174 (N_1174,N_379,N_130);
xor U1175 (N_1175,N_229,N_594);
or U1176 (N_1176,N_117,N_367);
xor U1177 (N_1177,N_598,N_547);
and U1178 (N_1178,N_572,N_239);
nand U1179 (N_1179,N_420,N_131);
xnor U1180 (N_1180,N_444,N_521);
nor U1181 (N_1181,N_83,N_415);
nand U1182 (N_1182,N_367,N_278);
nor U1183 (N_1183,N_372,N_127);
or U1184 (N_1184,N_199,N_1);
xor U1185 (N_1185,N_120,N_188);
nand U1186 (N_1186,N_208,N_441);
and U1187 (N_1187,N_549,N_466);
or U1188 (N_1188,N_593,N_155);
xnor U1189 (N_1189,N_563,N_550);
or U1190 (N_1190,N_565,N_197);
or U1191 (N_1191,N_409,N_586);
xor U1192 (N_1192,N_152,N_29);
or U1193 (N_1193,N_124,N_4);
nor U1194 (N_1194,N_385,N_379);
and U1195 (N_1195,N_309,N_72);
and U1196 (N_1196,N_542,N_438);
nor U1197 (N_1197,N_382,N_231);
or U1198 (N_1198,N_404,N_58);
and U1199 (N_1199,N_454,N_339);
nand U1200 (N_1200,N_1172,N_1092);
xnor U1201 (N_1201,N_644,N_1184);
or U1202 (N_1202,N_1190,N_723);
xnor U1203 (N_1203,N_671,N_818);
and U1204 (N_1204,N_995,N_978);
xor U1205 (N_1205,N_785,N_884);
nor U1206 (N_1206,N_1125,N_801);
nand U1207 (N_1207,N_639,N_805);
xor U1208 (N_1208,N_1164,N_969);
nor U1209 (N_1209,N_889,N_989);
nor U1210 (N_1210,N_1036,N_614);
or U1211 (N_1211,N_701,N_1144);
and U1212 (N_1212,N_632,N_925);
nand U1213 (N_1213,N_651,N_630);
xnor U1214 (N_1214,N_781,N_893);
nand U1215 (N_1215,N_1014,N_1102);
or U1216 (N_1216,N_1162,N_763);
xnor U1217 (N_1217,N_638,N_856);
or U1218 (N_1218,N_771,N_849);
xor U1219 (N_1219,N_985,N_615);
and U1220 (N_1220,N_1173,N_980);
xor U1221 (N_1221,N_600,N_1143);
nor U1222 (N_1222,N_887,N_888);
nand U1223 (N_1223,N_761,N_735);
or U1224 (N_1224,N_1131,N_959);
and U1225 (N_1225,N_619,N_691);
or U1226 (N_1226,N_729,N_720);
nand U1227 (N_1227,N_1191,N_939);
and U1228 (N_1228,N_1115,N_1098);
or U1229 (N_1229,N_862,N_1060);
or U1230 (N_1230,N_690,N_853);
nor U1231 (N_1231,N_695,N_997);
xnor U1232 (N_1232,N_869,N_882);
nor U1233 (N_1233,N_738,N_610);
nand U1234 (N_1234,N_859,N_611);
or U1235 (N_1235,N_1076,N_830);
nor U1236 (N_1236,N_758,N_660);
nand U1237 (N_1237,N_672,N_979);
nor U1238 (N_1238,N_784,N_1166);
nand U1239 (N_1239,N_1029,N_663);
xnor U1240 (N_1240,N_1185,N_1159);
xnor U1241 (N_1241,N_1196,N_800);
xnor U1242 (N_1242,N_659,N_773);
or U1243 (N_1243,N_1012,N_649);
nand U1244 (N_1244,N_1199,N_1118);
and U1245 (N_1245,N_652,N_824);
nor U1246 (N_1246,N_850,N_1157);
nor U1247 (N_1247,N_861,N_1152);
xor U1248 (N_1248,N_1129,N_1073);
nor U1249 (N_1249,N_950,N_832);
and U1250 (N_1250,N_1160,N_1198);
nand U1251 (N_1251,N_694,N_993);
xnor U1252 (N_1252,N_1178,N_1021);
and U1253 (N_1253,N_909,N_836);
nand U1254 (N_1254,N_971,N_1111);
or U1255 (N_1255,N_1141,N_713);
nand U1256 (N_1256,N_725,N_1007);
or U1257 (N_1257,N_747,N_1083);
xnor U1258 (N_1258,N_1019,N_1182);
or U1259 (N_1259,N_791,N_780);
nand U1260 (N_1260,N_878,N_1193);
or U1261 (N_1261,N_870,N_838);
nand U1262 (N_1262,N_911,N_1024);
or U1263 (N_1263,N_1179,N_696);
xnor U1264 (N_1264,N_1097,N_745);
xnor U1265 (N_1265,N_966,N_1120);
nor U1266 (N_1266,N_762,N_1080);
or U1267 (N_1267,N_721,N_679);
xor U1268 (N_1268,N_846,N_1009);
nor U1269 (N_1269,N_1049,N_743);
xor U1270 (N_1270,N_1069,N_1169);
or U1271 (N_1271,N_627,N_1081);
and U1272 (N_1272,N_689,N_1057);
nor U1273 (N_1273,N_1026,N_932);
nor U1274 (N_1274,N_683,N_1041);
xor U1275 (N_1275,N_907,N_931);
and U1276 (N_1276,N_1124,N_1093);
nand U1277 (N_1277,N_914,N_858);
or U1278 (N_1278,N_955,N_899);
or U1279 (N_1279,N_718,N_1094);
xnor U1280 (N_1280,N_618,N_647);
nor U1281 (N_1281,N_839,N_686);
nand U1282 (N_1282,N_1065,N_999);
and U1283 (N_1283,N_712,N_1064);
xor U1284 (N_1284,N_965,N_1058);
and U1285 (N_1285,N_1110,N_827);
or U1286 (N_1286,N_952,N_736);
nand U1287 (N_1287,N_885,N_898);
nand U1288 (N_1288,N_1035,N_669);
and U1289 (N_1289,N_769,N_936);
nand U1290 (N_1290,N_1071,N_788);
or U1291 (N_1291,N_626,N_837);
or U1292 (N_1292,N_646,N_891);
xnor U1293 (N_1293,N_1194,N_1126);
nor U1294 (N_1294,N_670,N_1084);
or U1295 (N_1295,N_992,N_1167);
and U1296 (N_1296,N_752,N_730);
nand U1297 (N_1297,N_977,N_746);
xor U1298 (N_1298,N_1105,N_928);
and U1299 (N_1299,N_819,N_1062);
nor U1300 (N_1300,N_879,N_783);
nand U1301 (N_1301,N_1030,N_903);
and U1302 (N_1302,N_1015,N_806);
nand U1303 (N_1303,N_1032,N_1011);
nor U1304 (N_1304,N_883,N_854);
nand U1305 (N_1305,N_820,N_1176);
and U1306 (N_1306,N_643,N_620);
and U1307 (N_1307,N_1042,N_1135);
nor U1308 (N_1308,N_943,N_1170);
nand U1309 (N_1309,N_601,N_662);
xor U1310 (N_1310,N_1163,N_896);
nor U1311 (N_1311,N_1089,N_812);
nand U1312 (N_1312,N_717,N_641);
or U1313 (N_1313,N_1122,N_1139);
or U1314 (N_1314,N_1038,N_1028);
nor U1315 (N_1315,N_948,N_1180);
nand U1316 (N_1316,N_933,N_940);
nand U1317 (N_1317,N_692,N_1077);
xnor U1318 (N_1318,N_779,N_634);
nand U1319 (N_1319,N_960,N_942);
xor U1320 (N_1320,N_1040,N_727);
or U1321 (N_1321,N_1006,N_704);
or U1322 (N_1322,N_816,N_1186);
nor U1323 (N_1323,N_1103,N_857);
or U1324 (N_1324,N_1043,N_777);
and U1325 (N_1325,N_617,N_922);
and U1326 (N_1326,N_635,N_828);
and U1327 (N_1327,N_1059,N_871);
nand U1328 (N_1328,N_860,N_708);
or U1329 (N_1329,N_1020,N_1161);
and U1330 (N_1330,N_908,N_865);
nand U1331 (N_1331,N_719,N_1044);
nand U1332 (N_1332,N_1133,N_797);
xor U1333 (N_1333,N_1134,N_938);
nand U1334 (N_1334,N_776,N_890);
nor U1335 (N_1335,N_757,N_741);
nand U1336 (N_1336,N_749,N_902);
and U1337 (N_1337,N_616,N_687);
nor U1338 (N_1338,N_786,N_789);
nor U1339 (N_1339,N_673,N_920);
or U1340 (N_1340,N_733,N_1121);
xnor U1341 (N_1341,N_608,N_768);
nand U1342 (N_1342,N_603,N_1087);
and U1343 (N_1343,N_655,N_904);
or U1344 (N_1344,N_653,N_1000);
nor U1345 (N_1345,N_956,N_748);
and U1346 (N_1346,N_935,N_1096);
or U1347 (N_1347,N_1188,N_919);
and U1348 (N_1348,N_764,N_724);
or U1349 (N_1349,N_778,N_905);
nor U1350 (N_1350,N_740,N_1066);
nand U1351 (N_1351,N_848,N_1106);
xor U1352 (N_1352,N_961,N_983);
and U1353 (N_1353,N_732,N_866);
nand U1354 (N_1354,N_991,N_715);
and U1355 (N_1355,N_1068,N_1095);
xor U1356 (N_1356,N_1154,N_640);
nor U1357 (N_1357,N_803,N_633);
or U1358 (N_1358,N_607,N_731);
or U1359 (N_1359,N_1136,N_613);
xor U1360 (N_1360,N_996,N_1148);
and U1361 (N_1361,N_901,N_1055);
nand U1362 (N_1362,N_1100,N_954);
and U1363 (N_1363,N_1048,N_872);
or U1364 (N_1364,N_1189,N_946);
nor U1365 (N_1365,N_825,N_1197);
nor U1366 (N_1366,N_1079,N_648);
or U1367 (N_1367,N_1017,N_897);
or U1368 (N_1368,N_787,N_875);
or U1369 (N_1369,N_759,N_976);
nor U1370 (N_1370,N_900,N_1023);
nor U1371 (N_1371,N_750,N_705);
and U1372 (N_1372,N_967,N_760);
or U1373 (N_1373,N_1054,N_913);
and U1374 (N_1374,N_1132,N_821);
nand U1375 (N_1375,N_700,N_947);
nand U1376 (N_1376,N_681,N_794);
or U1377 (N_1377,N_612,N_918);
nand U1378 (N_1378,N_877,N_1099);
or U1379 (N_1379,N_957,N_605);
xor U1380 (N_1380,N_1177,N_988);
and U1381 (N_1381,N_1010,N_1153);
nor U1382 (N_1382,N_894,N_804);
nor U1383 (N_1383,N_751,N_1123);
and U1384 (N_1384,N_728,N_929);
and U1385 (N_1385,N_1072,N_667);
and U1386 (N_1386,N_814,N_685);
xor U1387 (N_1387,N_1142,N_1151);
nor U1388 (N_1388,N_772,N_765);
and U1389 (N_1389,N_906,N_756);
or U1390 (N_1390,N_1074,N_964);
nand U1391 (N_1391,N_972,N_628);
nor U1392 (N_1392,N_684,N_709);
nor U1393 (N_1393,N_974,N_1149);
or U1394 (N_1394,N_1114,N_1047);
nor U1395 (N_1395,N_1104,N_1085);
and U1396 (N_1396,N_910,N_767);
or U1397 (N_1397,N_1016,N_1187);
nand U1398 (N_1398,N_968,N_1061);
or U1399 (N_1399,N_833,N_984);
and U1400 (N_1400,N_822,N_637);
nor U1401 (N_1401,N_624,N_987);
or U1402 (N_1402,N_1165,N_1018);
nor U1403 (N_1403,N_739,N_829);
and U1404 (N_1404,N_1116,N_1001);
nor U1405 (N_1405,N_766,N_676);
and U1406 (N_1406,N_699,N_1051);
xor U1407 (N_1407,N_881,N_1128);
or U1408 (N_1408,N_606,N_1145);
and U1409 (N_1409,N_847,N_722);
nand U1410 (N_1410,N_675,N_798);
and U1411 (N_1411,N_1181,N_698);
and U1412 (N_1412,N_1091,N_1146);
nor U1413 (N_1413,N_625,N_1127);
and U1414 (N_1414,N_1025,N_710);
or U1415 (N_1415,N_1070,N_795);
and U1416 (N_1416,N_944,N_842);
nor U1417 (N_1417,N_963,N_873);
xor U1418 (N_1418,N_915,N_1031);
xor U1419 (N_1419,N_753,N_1003);
xor U1420 (N_1420,N_657,N_799);
nand U1421 (N_1421,N_937,N_845);
or U1422 (N_1422,N_868,N_927);
xnor U1423 (N_1423,N_986,N_1174);
and U1424 (N_1424,N_975,N_1067);
and U1425 (N_1425,N_934,N_941);
and U1426 (N_1426,N_755,N_1138);
nand U1427 (N_1427,N_1192,N_754);
and U1428 (N_1428,N_949,N_835);
xor U1429 (N_1429,N_770,N_1022);
and U1430 (N_1430,N_1130,N_665);
and U1431 (N_1431,N_664,N_930);
or U1432 (N_1432,N_1195,N_834);
or U1433 (N_1433,N_734,N_623);
xnor U1434 (N_1434,N_823,N_1156);
nor U1435 (N_1435,N_1052,N_994);
nand U1436 (N_1436,N_656,N_1109);
nand U1437 (N_1437,N_1056,N_923);
or U1438 (N_1438,N_668,N_714);
xor U1439 (N_1439,N_711,N_742);
xor U1440 (N_1440,N_1013,N_962);
and U1441 (N_1441,N_645,N_1168);
xor U1442 (N_1442,N_843,N_1039);
nor U1443 (N_1443,N_1086,N_1112);
and U1444 (N_1444,N_707,N_796);
nor U1445 (N_1445,N_1002,N_982);
and U1446 (N_1446,N_677,N_726);
and U1447 (N_1447,N_990,N_790);
nor U1448 (N_1448,N_867,N_809);
nand U1449 (N_1449,N_831,N_921);
xor U1450 (N_1450,N_678,N_1078);
nor U1451 (N_1451,N_1137,N_737);
and U1452 (N_1452,N_1027,N_1101);
nor U1453 (N_1453,N_693,N_863);
nand U1454 (N_1454,N_1158,N_661);
or U1455 (N_1455,N_774,N_706);
or U1456 (N_1456,N_841,N_631);
or U1457 (N_1457,N_916,N_792);
xor U1458 (N_1458,N_658,N_945);
nor U1459 (N_1459,N_973,N_951);
or U1460 (N_1460,N_636,N_926);
or U1461 (N_1461,N_650,N_1117);
and U1462 (N_1462,N_688,N_1045);
or U1463 (N_1463,N_981,N_642);
or U1464 (N_1464,N_1037,N_1005);
or U1465 (N_1465,N_622,N_1171);
nor U1466 (N_1466,N_1063,N_1113);
nand U1467 (N_1467,N_1147,N_844);
or U1468 (N_1468,N_998,N_1034);
nand U1469 (N_1469,N_654,N_1183);
nand U1470 (N_1470,N_782,N_602);
and U1471 (N_1471,N_851,N_958);
xor U1472 (N_1472,N_840,N_917);
or U1473 (N_1473,N_1108,N_924);
xor U1474 (N_1474,N_1155,N_702);
or U1475 (N_1475,N_793,N_666);
nor U1476 (N_1476,N_953,N_1175);
nor U1477 (N_1477,N_1004,N_680);
xnor U1478 (N_1478,N_1088,N_802);
or U1479 (N_1479,N_629,N_1140);
nor U1480 (N_1480,N_864,N_1090);
or U1481 (N_1481,N_775,N_1046);
xor U1482 (N_1482,N_621,N_1119);
nor U1483 (N_1483,N_892,N_604);
nor U1484 (N_1484,N_1033,N_674);
nor U1485 (N_1485,N_682,N_876);
and U1486 (N_1486,N_895,N_813);
or U1487 (N_1487,N_970,N_807);
nand U1488 (N_1488,N_1075,N_697);
nor U1489 (N_1489,N_874,N_912);
and U1490 (N_1490,N_703,N_815);
xor U1491 (N_1491,N_810,N_1150);
nand U1492 (N_1492,N_811,N_1082);
and U1493 (N_1493,N_716,N_1107);
nor U1494 (N_1494,N_817,N_1050);
xor U1495 (N_1495,N_826,N_852);
and U1496 (N_1496,N_1053,N_609);
or U1497 (N_1497,N_855,N_744);
nor U1498 (N_1498,N_808,N_1008);
xnor U1499 (N_1499,N_886,N_880);
xor U1500 (N_1500,N_872,N_897);
nor U1501 (N_1501,N_888,N_750);
and U1502 (N_1502,N_1080,N_1191);
and U1503 (N_1503,N_685,N_1154);
or U1504 (N_1504,N_749,N_623);
or U1505 (N_1505,N_1184,N_679);
or U1506 (N_1506,N_669,N_683);
and U1507 (N_1507,N_954,N_842);
nor U1508 (N_1508,N_1010,N_627);
nand U1509 (N_1509,N_968,N_868);
and U1510 (N_1510,N_1047,N_785);
xnor U1511 (N_1511,N_1016,N_1087);
and U1512 (N_1512,N_673,N_927);
xor U1513 (N_1513,N_895,N_906);
and U1514 (N_1514,N_734,N_920);
xnor U1515 (N_1515,N_624,N_670);
and U1516 (N_1516,N_1093,N_958);
nand U1517 (N_1517,N_835,N_1020);
xnor U1518 (N_1518,N_756,N_707);
or U1519 (N_1519,N_1088,N_833);
xor U1520 (N_1520,N_838,N_731);
and U1521 (N_1521,N_701,N_1105);
or U1522 (N_1522,N_776,N_875);
and U1523 (N_1523,N_606,N_842);
nor U1524 (N_1524,N_1091,N_902);
xnor U1525 (N_1525,N_908,N_1170);
and U1526 (N_1526,N_1152,N_600);
nand U1527 (N_1527,N_1113,N_966);
nor U1528 (N_1528,N_1126,N_610);
and U1529 (N_1529,N_742,N_1087);
and U1530 (N_1530,N_1021,N_1001);
nor U1531 (N_1531,N_675,N_620);
nand U1532 (N_1532,N_911,N_1131);
nand U1533 (N_1533,N_1019,N_979);
nor U1534 (N_1534,N_852,N_749);
nor U1535 (N_1535,N_627,N_738);
xnor U1536 (N_1536,N_892,N_717);
xnor U1537 (N_1537,N_1010,N_616);
xnor U1538 (N_1538,N_1027,N_1137);
nor U1539 (N_1539,N_802,N_1106);
or U1540 (N_1540,N_643,N_960);
nand U1541 (N_1541,N_879,N_1174);
nor U1542 (N_1542,N_667,N_681);
or U1543 (N_1543,N_812,N_790);
nor U1544 (N_1544,N_1168,N_803);
nor U1545 (N_1545,N_921,N_1136);
xor U1546 (N_1546,N_1050,N_647);
or U1547 (N_1547,N_633,N_955);
xor U1548 (N_1548,N_1081,N_1053);
and U1549 (N_1549,N_1095,N_670);
xnor U1550 (N_1550,N_1051,N_1036);
or U1551 (N_1551,N_783,N_960);
nand U1552 (N_1552,N_660,N_669);
and U1553 (N_1553,N_723,N_971);
or U1554 (N_1554,N_1195,N_780);
nand U1555 (N_1555,N_706,N_737);
nor U1556 (N_1556,N_1033,N_844);
or U1557 (N_1557,N_960,N_861);
or U1558 (N_1558,N_1136,N_775);
and U1559 (N_1559,N_921,N_973);
and U1560 (N_1560,N_1163,N_1036);
nor U1561 (N_1561,N_882,N_1119);
nand U1562 (N_1562,N_1055,N_1093);
or U1563 (N_1563,N_987,N_1125);
nand U1564 (N_1564,N_1067,N_782);
or U1565 (N_1565,N_854,N_1125);
xnor U1566 (N_1566,N_682,N_668);
xnor U1567 (N_1567,N_739,N_907);
nor U1568 (N_1568,N_724,N_994);
and U1569 (N_1569,N_604,N_753);
or U1570 (N_1570,N_1058,N_975);
or U1571 (N_1571,N_717,N_837);
nor U1572 (N_1572,N_1143,N_863);
and U1573 (N_1573,N_927,N_777);
and U1574 (N_1574,N_1091,N_1156);
or U1575 (N_1575,N_696,N_1029);
and U1576 (N_1576,N_833,N_970);
xnor U1577 (N_1577,N_841,N_899);
nor U1578 (N_1578,N_786,N_936);
nor U1579 (N_1579,N_678,N_1018);
nand U1580 (N_1580,N_1175,N_805);
xnor U1581 (N_1581,N_651,N_828);
and U1582 (N_1582,N_760,N_711);
and U1583 (N_1583,N_750,N_1107);
or U1584 (N_1584,N_709,N_650);
or U1585 (N_1585,N_1093,N_1008);
xnor U1586 (N_1586,N_815,N_1050);
nand U1587 (N_1587,N_788,N_951);
and U1588 (N_1588,N_1030,N_1178);
or U1589 (N_1589,N_702,N_893);
xnor U1590 (N_1590,N_822,N_1054);
and U1591 (N_1591,N_1007,N_679);
nand U1592 (N_1592,N_1158,N_637);
xor U1593 (N_1593,N_937,N_995);
nand U1594 (N_1594,N_695,N_755);
nor U1595 (N_1595,N_994,N_836);
xor U1596 (N_1596,N_607,N_895);
or U1597 (N_1597,N_1019,N_656);
nand U1598 (N_1598,N_1175,N_995);
or U1599 (N_1599,N_632,N_1042);
nand U1600 (N_1600,N_897,N_968);
nor U1601 (N_1601,N_604,N_870);
nor U1602 (N_1602,N_771,N_605);
nand U1603 (N_1603,N_1098,N_718);
nor U1604 (N_1604,N_1061,N_844);
or U1605 (N_1605,N_962,N_808);
or U1606 (N_1606,N_1068,N_1133);
nor U1607 (N_1607,N_861,N_1093);
and U1608 (N_1608,N_1082,N_932);
nand U1609 (N_1609,N_619,N_1010);
and U1610 (N_1610,N_1155,N_1067);
nand U1611 (N_1611,N_935,N_841);
nand U1612 (N_1612,N_996,N_1037);
and U1613 (N_1613,N_1013,N_788);
xnor U1614 (N_1614,N_1176,N_834);
xnor U1615 (N_1615,N_1157,N_664);
or U1616 (N_1616,N_798,N_925);
and U1617 (N_1617,N_689,N_1035);
and U1618 (N_1618,N_1000,N_857);
or U1619 (N_1619,N_819,N_631);
nor U1620 (N_1620,N_1172,N_974);
xnor U1621 (N_1621,N_1055,N_907);
nand U1622 (N_1622,N_794,N_601);
nor U1623 (N_1623,N_713,N_1180);
nand U1624 (N_1624,N_899,N_1057);
or U1625 (N_1625,N_641,N_1035);
nor U1626 (N_1626,N_698,N_999);
or U1627 (N_1627,N_1108,N_624);
and U1628 (N_1628,N_973,N_1055);
nand U1629 (N_1629,N_854,N_1028);
xor U1630 (N_1630,N_604,N_839);
xnor U1631 (N_1631,N_684,N_1068);
or U1632 (N_1632,N_1069,N_621);
and U1633 (N_1633,N_714,N_690);
xnor U1634 (N_1634,N_1040,N_691);
and U1635 (N_1635,N_768,N_733);
or U1636 (N_1636,N_1070,N_816);
nor U1637 (N_1637,N_622,N_619);
nor U1638 (N_1638,N_960,N_980);
nor U1639 (N_1639,N_838,N_667);
or U1640 (N_1640,N_999,N_765);
and U1641 (N_1641,N_643,N_690);
nand U1642 (N_1642,N_1173,N_748);
xnor U1643 (N_1643,N_777,N_806);
xnor U1644 (N_1644,N_923,N_991);
xnor U1645 (N_1645,N_938,N_692);
nor U1646 (N_1646,N_782,N_856);
xnor U1647 (N_1647,N_1025,N_1044);
nor U1648 (N_1648,N_1068,N_655);
and U1649 (N_1649,N_1146,N_945);
xnor U1650 (N_1650,N_1130,N_657);
and U1651 (N_1651,N_616,N_1111);
or U1652 (N_1652,N_1189,N_1049);
nand U1653 (N_1653,N_706,N_613);
nor U1654 (N_1654,N_1039,N_919);
xor U1655 (N_1655,N_907,N_888);
and U1656 (N_1656,N_963,N_689);
and U1657 (N_1657,N_1106,N_609);
nor U1658 (N_1658,N_743,N_887);
xor U1659 (N_1659,N_1129,N_658);
or U1660 (N_1660,N_982,N_718);
nand U1661 (N_1661,N_933,N_1117);
xnor U1662 (N_1662,N_773,N_922);
nor U1663 (N_1663,N_737,N_623);
and U1664 (N_1664,N_1007,N_969);
nand U1665 (N_1665,N_1116,N_1047);
xor U1666 (N_1666,N_1144,N_610);
xor U1667 (N_1667,N_653,N_855);
or U1668 (N_1668,N_822,N_606);
and U1669 (N_1669,N_724,N_1019);
xor U1670 (N_1670,N_763,N_1112);
xnor U1671 (N_1671,N_912,N_694);
nand U1672 (N_1672,N_869,N_935);
nor U1673 (N_1673,N_688,N_978);
and U1674 (N_1674,N_747,N_820);
or U1675 (N_1675,N_661,N_741);
and U1676 (N_1676,N_784,N_864);
nand U1677 (N_1677,N_696,N_1144);
nor U1678 (N_1678,N_627,N_749);
and U1679 (N_1679,N_742,N_1029);
nand U1680 (N_1680,N_906,N_1035);
nand U1681 (N_1681,N_628,N_936);
xor U1682 (N_1682,N_1123,N_838);
xor U1683 (N_1683,N_766,N_1169);
nor U1684 (N_1684,N_873,N_879);
or U1685 (N_1685,N_876,N_811);
or U1686 (N_1686,N_614,N_1070);
nor U1687 (N_1687,N_1027,N_838);
or U1688 (N_1688,N_846,N_854);
xnor U1689 (N_1689,N_813,N_841);
nor U1690 (N_1690,N_1071,N_1173);
xor U1691 (N_1691,N_1042,N_954);
nor U1692 (N_1692,N_1089,N_855);
or U1693 (N_1693,N_908,N_1185);
xor U1694 (N_1694,N_837,N_1107);
and U1695 (N_1695,N_919,N_887);
xnor U1696 (N_1696,N_1131,N_1049);
nand U1697 (N_1697,N_1014,N_830);
xnor U1698 (N_1698,N_764,N_601);
and U1699 (N_1699,N_983,N_1151);
nor U1700 (N_1700,N_1134,N_904);
nor U1701 (N_1701,N_715,N_1168);
xor U1702 (N_1702,N_969,N_973);
xnor U1703 (N_1703,N_1186,N_1068);
and U1704 (N_1704,N_797,N_667);
or U1705 (N_1705,N_768,N_1027);
or U1706 (N_1706,N_929,N_780);
nor U1707 (N_1707,N_1089,N_720);
or U1708 (N_1708,N_986,N_892);
and U1709 (N_1709,N_786,N_1181);
and U1710 (N_1710,N_798,N_690);
or U1711 (N_1711,N_635,N_1194);
xor U1712 (N_1712,N_1169,N_685);
nor U1713 (N_1713,N_608,N_861);
and U1714 (N_1714,N_1112,N_899);
nor U1715 (N_1715,N_779,N_839);
or U1716 (N_1716,N_631,N_806);
nor U1717 (N_1717,N_717,N_662);
and U1718 (N_1718,N_601,N_1108);
xnor U1719 (N_1719,N_842,N_1128);
or U1720 (N_1720,N_821,N_620);
xor U1721 (N_1721,N_876,N_867);
nand U1722 (N_1722,N_912,N_881);
and U1723 (N_1723,N_1160,N_707);
nand U1724 (N_1724,N_763,N_939);
nand U1725 (N_1725,N_715,N_860);
nor U1726 (N_1726,N_825,N_706);
xor U1727 (N_1727,N_871,N_833);
or U1728 (N_1728,N_1110,N_763);
nor U1729 (N_1729,N_950,N_640);
and U1730 (N_1730,N_786,N_1003);
xnor U1731 (N_1731,N_608,N_870);
and U1732 (N_1732,N_803,N_984);
xnor U1733 (N_1733,N_931,N_773);
and U1734 (N_1734,N_814,N_821);
xnor U1735 (N_1735,N_643,N_1014);
nand U1736 (N_1736,N_734,N_706);
xnor U1737 (N_1737,N_709,N_1100);
xor U1738 (N_1738,N_822,N_1121);
nor U1739 (N_1739,N_744,N_655);
and U1740 (N_1740,N_764,N_826);
nor U1741 (N_1741,N_711,N_720);
and U1742 (N_1742,N_752,N_994);
nand U1743 (N_1743,N_992,N_904);
or U1744 (N_1744,N_744,N_1015);
xor U1745 (N_1745,N_1035,N_1102);
and U1746 (N_1746,N_1132,N_860);
nand U1747 (N_1747,N_665,N_1095);
or U1748 (N_1748,N_766,N_1095);
nand U1749 (N_1749,N_948,N_956);
xor U1750 (N_1750,N_1129,N_838);
or U1751 (N_1751,N_1122,N_958);
nand U1752 (N_1752,N_1148,N_1085);
and U1753 (N_1753,N_1125,N_935);
xor U1754 (N_1754,N_737,N_1183);
or U1755 (N_1755,N_838,N_620);
and U1756 (N_1756,N_648,N_618);
xnor U1757 (N_1757,N_1094,N_856);
nor U1758 (N_1758,N_1178,N_726);
nor U1759 (N_1759,N_649,N_690);
and U1760 (N_1760,N_823,N_875);
nor U1761 (N_1761,N_751,N_969);
and U1762 (N_1762,N_1017,N_1093);
or U1763 (N_1763,N_600,N_1096);
and U1764 (N_1764,N_935,N_1073);
nand U1765 (N_1765,N_895,N_799);
or U1766 (N_1766,N_1102,N_1052);
xor U1767 (N_1767,N_627,N_774);
or U1768 (N_1768,N_731,N_1195);
xor U1769 (N_1769,N_727,N_628);
xor U1770 (N_1770,N_703,N_647);
or U1771 (N_1771,N_668,N_989);
nand U1772 (N_1772,N_848,N_754);
and U1773 (N_1773,N_1154,N_916);
and U1774 (N_1774,N_992,N_1110);
or U1775 (N_1775,N_843,N_958);
and U1776 (N_1776,N_835,N_976);
and U1777 (N_1777,N_1178,N_1162);
xor U1778 (N_1778,N_771,N_979);
or U1779 (N_1779,N_859,N_626);
xor U1780 (N_1780,N_928,N_744);
xor U1781 (N_1781,N_1040,N_815);
xor U1782 (N_1782,N_930,N_953);
or U1783 (N_1783,N_682,N_1001);
or U1784 (N_1784,N_693,N_813);
or U1785 (N_1785,N_629,N_1099);
nor U1786 (N_1786,N_730,N_832);
nand U1787 (N_1787,N_830,N_765);
nand U1788 (N_1788,N_654,N_823);
nand U1789 (N_1789,N_768,N_839);
or U1790 (N_1790,N_609,N_895);
and U1791 (N_1791,N_927,N_700);
and U1792 (N_1792,N_601,N_929);
nor U1793 (N_1793,N_929,N_765);
nor U1794 (N_1794,N_918,N_939);
xnor U1795 (N_1795,N_655,N_883);
nor U1796 (N_1796,N_868,N_1055);
nor U1797 (N_1797,N_1198,N_896);
and U1798 (N_1798,N_870,N_845);
xnor U1799 (N_1799,N_857,N_932);
and U1800 (N_1800,N_1427,N_1319);
or U1801 (N_1801,N_1221,N_1532);
and U1802 (N_1802,N_1323,N_1224);
nand U1803 (N_1803,N_1615,N_1249);
nor U1804 (N_1804,N_1527,N_1585);
xnor U1805 (N_1805,N_1459,N_1611);
nand U1806 (N_1806,N_1663,N_1783);
xor U1807 (N_1807,N_1481,N_1302);
xor U1808 (N_1808,N_1708,N_1778);
or U1809 (N_1809,N_1274,N_1538);
xor U1810 (N_1810,N_1376,N_1790);
xor U1811 (N_1811,N_1333,N_1410);
and U1812 (N_1812,N_1666,N_1702);
and U1813 (N_1813,N_1613,N_1502);
nand U1814 (N_1814,N_1200,N_1524);
and U1815 (N_1815,N_1353,N_1286);
xor U1816 (N_1816,N_1514,N_1581);
or U1817 (N_1817,N_1354,N_1639);
nand U1818 (N_1818,N_1272,N_1248);
xnor U1819 (N_1819,N_1363,N_1775);
nor U1820 (N_1820,N_1657,N_1403);
nor U1821 (N_1821,N_1564,N_1776);
xor U1822 (N_1822,N_1288,N_1505);
and U1823 (N_1823,N_1710,N_1223);
and U1824 (N_1824,N_1406,N_1332);
or U1825 (N_1825,N_1392,N_1417);
and U1826 (N_1826,N_1537,N_1294);
or U1827 (N_1827,N_1308,N_1281);
nand U1828 (N_1828,N_1706,N_1741);
nand U1829 (N_1829,N_1371,N_1599);
xor U1830 (N_1830,N_1602,N_1364);
and U1831 (N_1831,N_1667,N_1669);
or U1832 (N_1832,N_1253,N_1445);
nand U1833 (N_1833,N_1316,N_1604);
nand U1834 (N_1834,N_1550,N_1289);
xnor U1835 (N_1835,N_1408,N_1765);
or U1836 (N_1836,N_1265,N_1263);
nand U1837 (N_1837,N_1299,N_1689);
nand U1838 (N_1838,N_1356,N_1518);
and U1839 (N_1839,N_1589,N_1405);
or U1840 (N_1840,N_1691,N_1269);
nor U1841 (N_1841,N_1566,N_1322);
and U1842 (N_1842,N_1767,N_1206);
and U1843 (N_1843,N_1284,N_1535);
and U1844 (N_1844,N_1653,N_1305);
or U1845 (N_1845,N_1303,N_1693);
or U1846 (N_1846,N_1509,N_1492);
and U1847 (N_1847,N_1777,N_1222);
xnor U1848 (N_1848,N_1215,N_1692);
nand U1849 (N_1849,N_1632,N_1714);
or U1850 (N_1850,N_1598,N_1655);
nand U1851 (N_1851,N_1385,N_1780);
xor U1852 (N_1852,N_1601,N_1362);
nor U1853 (N_1853,N_1750,N_1234);
or U1854 (N_1854,N_1623,N_1497);
xor U1855 (N_1855,N_1225,N_1799);
and U1856 (N_1856,N_1243,N_1203);
or U1857 (N_1857,N_1582,N_1791);
nor U1858 (N_1858,N_1747,N_1619);
or U1859 (N_1859,N_1675,N_1761);
nand U1860 (N_1860,N_1477,N_1300);
or U1861 (N_1861,N_1740,N_1246);
xnor U1862 (N_1862,N_1454,N_1226);
or U1863 (N_1863,N_1268,N_1577);
nand U1864 (N_1864,N_1312,N_1484);
nor U1865 (N_1865,N_1526,N_1314);
xor U1866 (N_1866,N_1561,N_1315);
and U1867 (N_1867,N_1375,N_1628);
or U1868 (N_1868,N_1608,N_1549);
xor U1869 (N_1869,N_1307,N_1404);
xor U1870 (N_1870,N_1531,N_1437);
nand U1871 (N_1871,N_1503,N_1291);
nand U1872 (N_1872,N_1510,N_1489);
xnor U1873 (N_1873,N_1430,N_1600);
nand U1874 (N_1874,N_1681,N_1436);
and U1875 (N_1875,N_1652,N_1335);
nand U1876 (N_1876,N_1712,N_1355);
nor U1877 (N_1877,N_1208,N_1723);
nor U1878 (N_1878,N_1321,N_1352);
nand U1879 (N_1879,N_1540,N_1447);
nor U1880 (N_1880,N_1565,N_1758);
nand U1881 (N_1881,N_1482,N_1380);
nor U1882 (N_1882,N_1487,N_1627);
nand U1883 (N_1883,N_1432,N_1400);
and U1884 (N_1884,N_1409,N_1209);
nor U1885 (N_1885,N_1673,N_1256);
nor U1886 (N_1886,N_1368,N_1416);
xor U1887 (N_1887,N_1597,N_1635);
nand U1888 (N_1888,N_1202,N_1466);
xnor U1889 (N_1889,N_1782,N_1377);
xor U1890 (N_1890,N_1606,N_1562);
or U1891 (N_1891,N_1343,N_1516);
or U1892 (N_1892,N_1748,N_1647);
nand U1893 (N_1893,N_1444,N_1528);
and U1894 (N_1894,N_1396,N_1625);
nand U1895 (N_1895,N_1727,N_1230);
nor U1896 (N_1896,N_1580,N_1773);
xor U1897 (N_1897,N_1533,N_1501);
nor U1898 (N_1898,N_1751,N_1402);
xor U1899 (N_1899,N_1297,N_1434);
or U1900 (N_1900,N_1211,N_1794);
xor U1901 (N_1901,N_1388,N_1545);
and U1902 (N_1902,N_1257,N_1755);
nand U1903 (N_1903,N_1373,N_1245);
nor U1904 (N_1904,N_1424,N_1270);
and U1905 (N_1905,N_1534,N_1548);
nand U1906 (N_1906,N_1688,N_1590);
or U1907 (N_1907,N_1645,N_1218);
nor U1908 (N_1908,N_1413,N_1738);
xnor U1909 (N_1909,N_1563,N_1769);
or U1910 (N_1910,N_1576,N_1423);
nand U1911 (N_1911,N_1654,N_1390);
and U1912 (N_1912,N_1469,N_1442);
and U1913 (N_1913,N_1523,N_1642);
nand U1914 (N_1914,N_1609,N_1781);
nand U1915 (N_1915,N_1440,N_1631);
nand U1916 (N_1916,N_1347,N_1293);
nor U1917 (N_1917,N_1275,N_1217);
and U1918 (N_1918,N_1351,N_1212);
nor U1919 (N_1919,N_1586,N_1728);
and U1920 (N_1920,N_1746,N_1330);
xnor U1921 (N_1921,N_1683,N_1792);
nand U1922 (N_1922,N_1638,N_1743);
and U1923 (N_1923,N_1557,N_1651);
xnor U1924 (N_1924,N_1350,N_1662);
nor U1925 (N_1925,N_1273,N_1520);
xor U1926 (N_1926,N_1734,N_1278);
nor U1927 (N_1927,N_1344,N_1493);
nand U1928 (N_1928,N_1317,N_1467);
nand U1929 (N_1929,N_1452,N_1766);
xnor U1930 (N_1930,N_1480,N_1729);
or U1931 (N_1931,N_1719,N_1551);
or U1932 (N_1932,N_1742,N_1515);
and U1933 (N_1933,N_1641,N_1367);
nor U1934 (N_1934,N_1461,N_1471);
nand U1935 (N_1935,N_1235,N_1379);
nand U1936 (N_1936,N_1560,N_1438);
and U1937 (N_1937,N_1517,N_1340);
nor U1938 (N_1938,N_1709,N_1448);
or U1939 (N_1939,N_1703,N_1698);
xnor U1940 (N_1940,N_1610,N_1694);
or U1941 (N_1941,N_1787,N_1711);
nand U1942 (N_1942,N_1690,N_1659);
and U1943 (N_1943,N_1525,N_1282);
nand U1944 (N_1944,N_1313,N_1365);
and U1945 (N_1945,N_1578,N_1626);
or U1946 (N_1946,N_1464,N_1213);
nand U1947 (N_1947,N_1456,N_1513);
nand U1948 (N_1948,N_1399,N_1425);
and U1949 (N_1949,N_1473,N_1287);
nor U1950 (N_1950,N_1401,N_1369);
nor U1951 (N_1951,N_1228,N_1559);
nand U1952 (N_1952,N_1721,N_1779);
xnor U1953 (N_1953,N_1393,N_1682);
or U1954 (N_1954,N_1359,N_1391);
xor U1955 (N_1955,N_1762,N_1499);
xor U1956 (N_1956,N_1737,N_1646);
nor U1957 (N_1957,N_1558,N_1543);
nand U1958 (N_1958,N_1680,N_1726);
nand U1959 (N_1959,N_1552,N_1267);
xnor U1960 (N_1960,N_1650,N_1668);
nand U1961 (N_1961,N_1414,N_1784);
nand U1962 (N_1962,N_1759,N_1412);
nand U1963 (N_1963,N_1595,N_1259);
nor U1964 (N_1964,N_1725,N_1536);
or U1965 (N_1965,N_1756,N_1700);
nor U1966 (N_1966,N_1227,N_1512);
and U1967 (N_1967,N_1588,N_1389);
xnor U1968 (N_1968,N_1507,N_1342);
xnor U1969 (N_1969,N_1327,N_1339);
and U1970 (N_1970,N_1629,N_1519);
and U1971 (N_1971,N_1617,N_1271);
and U1972 (N_1972,N_1656,N_1772);
nor U1973 (N_1973,N_1384,N_1205);
nor U1974 (N_1974,N_1449,N_1546);
or U1975 (N_1975,N_1699,N_1311);
xnor U1976 (N_1976,N_1242,N_1357);
nor U1977 (N_1977,N_1630,N_1522);
or U1978 (N_1978,N_1696,N_1572);
nor U1979 (N_1979,N_1660,N_1705);
and U1980 (N_1980,N_1504,N_1511);
nor U1981 (N_1981,N_1435,N_1574);
xor U1982 (N_1982,N_1240,N_1397);
nor U1983 (N_1983,N_1496,N_1798);
xor U1984 (N_1984,N_1443,N_1500);
and U1985 (N_1985,N_1260,N_1796);
nand U1986 (N_1986,N_1764,N_1422);
nor U1987 (N_1987,N_1621,N_1789);
or U1988 (N_1988,N_1648,N_1745);
nand U1989 (N_1989,N_1661,N_1664);
xnor U1990 (N_1990,N_1567,N_1716);
nor U1991 (N_1991,N_1382,N_1407);
or U1992 (N_1992,N_1338,N_1450);
xnor U1993 (N_1993,N_1633,N_1429);
and U1994 (N_1994,N_1383,N_1475);
or U1995 (N_1995,N_1236,N_1325);
xor U1996 (N_1996,N_1361,N_1460);
nand U1997 (N_1997,N_1279,N_1250);
nand U1998 (N_1998,N_1793,N_1658);
xor U1999 (N_1999,N_1326,N_1398);
xnor U2000 (N_2000,N_1569,N_1718);
xnor U2001 (N_2001,N_1283,N_1207);
nor U2002 (N_2002,N_1622,N_1266);
nor U2003 (N_2003,N_1770,N_1607);
nand U2004 (N_2004,N_1555,N_1547);
nor U2005 (N_2005,N_1553,N_1395);
xor U2006 (N_2006,N_1570,N_1468);
nor U2007 (N_2007,N_1679,N_1331);
or U2008 (N_2008,N_1470,N_1672);
and U2009 (N_2009,N_1421,N_1214);
and U2010 (N_2010,N_1634,N_1320);
nor U2011 (N_2011,N_1735,N_1612);
xnor U2012 (N_2012,N_1584,N_1695);
nand U2013 (N_2013,N_1329,N_1378);
nand U2014 (N_2014,N_1684,N_1483);
nand U2015 (N_2015,N_1579,N_1730);
nand U2016 (N_2016,N_1453,N_1381);
nand U2017 (N_2017,N_1788,N_1757);
or U2018 (N_2018,N_1310,N_1446);
nor U2019 (N_2019,N_1462,N_1508);
xnor U2020 (N_2020,N_1754,N_1760);
and U2021 (N_2021,N_1605,N_1345);
nand U2022 (N_2022,N_1678,N_1201);
nand U2023 (N_2023,N_1304,N_1276);
nand U2024 (N_2024,N_1797,N_1341);
and U2025 (N_2025,N_1334,N_1328);
nor U2026 (N_2026,N_1583,N_1318);
or U2027 (N_2027,N_1458,N_1624);
nand U2028 (N_2028,N_1665,N_1258);
nand U2029 (N_2029,N_1697,N_1620);
and U2030 (N_2030,N_1337,N_1204);
or U2031 (N_2031,N_1336,N_1370);
nor U2032 (N_2032,N_1616,N_1433);
nor U2033 (N_2033,N_1372,N_1387);
or U2034 (N_2034,N_1231,N_1255);
or U2035 (N_2035,N_1591,N_1731);
and U2036 (N_2036,N_1704,N_1426);
or U2037 (N_2037,N_1592,N_1237);
nor U2038 (N_2038,N_1457,N_1476);
nor U2039 (N_2039,N_1455,N_1571);
nand U2040 (N_2040,N_1394,N_1229);
nand U2041 (N_2041,N_1254,N_1292);
xnor U2042 (N_2042,N_1431,N_1262);
nor U2043 (N_2043,N_1349,N_1506);
and U2044 (N_2044,N_1324,N_1238);
or U2045 (N_2045,N_1771,N_1774);
or U2046 (N_2046,N_1795,N_1587);
nand U2047 (N_2047,N_1753,N_1306);
nor U2048 (N_2048,N_1707,N_1358);
nand U2049 (N_2049,N_1749,N_1247);
xor U2050 (N_2050,N_1251,N_1239);
and U2051 (N_2051,N_1309,N_1277);
nor U2052 (N_2052,N_1539,N_1744);
or U2053 (N_2053,N_1596,N_1441);
nand U2054 (N_2054,N_1219,N_1722);
or U2055 (N_2055,N_1530,N_1261);
nor U2056 (N_2056,N_1244,N_1301);
and U2057 (N_2057,N_1415,N_1374);
and U2058 (N_2058,N_1210,N_1541);
nand U2059 (N_2059,N_1736,N_1713);
nor U2060 (N_2060,N_1348,N_1439);
nand U2061 (N_2061,N_1686,N_1474);
nand U2062 (N_2062,N_1640,N_1644);
xor U2063 (N_2063,N_1490,N_1544);
or U2064 (N_2064,N_1485,N_1732);
nor U2065 (N_2065,N_1542,N_1280);
nor U2066 (N_2066,N_1419,N_1252);
or U2067 (N_2067,N_1360,N_1676);
nand U2068 (N_2068,N_1685,N_1594);
nand U2069 (N_2069,N_1701,N_1498);
nand U2070 (N_2070,N_1285,N_1495);
nand U2071 (N_2071,N_1529,N_1593);
or U2072 (N_2072,N_1479,N_1346);
nor U2073 (N_2073,N_1298,N_1216);
nor U2074 (N_2074,N_1290,N_1494);
or U2075 (N_2075,N_1603,N_1739);
and U2076 (N_2076,N_1573,N_1637);
or U2077 (N_2077,N_1687,N_1521);
nor U2078 (N_2078,N_1478,N_1556);
or U2079 (N_2079,N_1752,N_1232);
nor U2080 (N_2080,N_1671,N_1428);
or U2081 (N_2081,N_1670,N_1386);
nor U2082 (N_2082,N_1554,N_1488);
xnor U2083 (N_2083,N_1674,N_1241);
xor U2084 (N_2084,N_1575,N_1472);
nand U2085 (N_2085,N_1643,N_1618);
and U2086 (N_2086,N_1724,N_1233);
nor U2087 (N_2087,N_1636,N_1465);
and U2088 (N_2088,N_1295,N_1720);
and U2089 (N_2089,N_1785,N_1568);
or U2090 (N_2090,N_1677,N_1411);
or U2091 (N_2091,N_1614,N_1296);
xnor U2092 (N_2092,N_1463,N_1264);
nand U2093 (N_2093,N_1649,N_1763);
nor U2094 (N_2094,N_1366,N_1491);
nor U2095 (N_2095,N_1220,N_1717);
or U2096 (N_2096,N_1786,N_1733);
xnor U2097 (N_2097,N_1486,N_1418);
or U2098 (N_2098,N_1420,N_1768);
or U2099 (N_2099,N_1451,N_1715);
nor U2100 (N_2100,N_1250,N_1738);
and U2101 (N_2101,N_1716,N_1770);
nand U2102 (N_2102,N_1578,N_1285);
nor U2103 (N_2103,N_1302,N_1665);
nand U2104 (N_2104,N_1294,N_1712);
xor U2105 (N_2105,N_1557,N_1736);
nand U2106 (N_2106,N_1284,N_1365);
nand U2107 (N_2107,N_1340,N_1745);
nor U2108 (N_2108,N_1345,N_1283);
and U2109 (N_2109,N_1621,N_1521);
and U2110 (N_2110,N_1762,N_1476);
and U2111 (N_2111,N_1713,N_1461);
nor U2112 (N_2112,N_1396,N_1456);
nand U2113 (N_2113,N_1225,N_1388);
and U2114 (N_2114,N_1553,N_1372);
nor U2115 (N_2115,N_1609,N_1700);
nand U2116 (N_2116,N_1659,N_1724);
and U2117 (N_2117,N_1573,N_1361);
nand U2118 (N_2118,N_1667,N_1273);
or U2119 (N_2119,N_1608,N_1246);
and U2120 (N_2120,N_1286,N_1536);
xnor U2121 (N_2121,N_1667,N_1514);
and U2122 (N_2122,N_1301,N_1586);
xnor U2123 (N_2123,N_1596,N_1467);
nor U2124 (N_2124,N_1450,N_1755);
nor U2125 (N_2125,N_1554,N_1782);
xnor U2126 (N_2126,N_1680,N_1207);
and U2127 (N_2127,N_1355,N_1332);
or U2128 (N_2128,N_1470,N_1696);
nand U2129 (N_2129,N_1622,N_1624);
nor U2130 (N_2130,N_1331,N_1270);
nand U2131 (N_2131,N_1787,N_1738);
and U2132 (N_2132,N_1287,N_1224);
xnor U2133 (N_2133,N_1325,N_1511);
xor U2134 (N_2134,N_1743,N_1626);
nor U2135 (N_2135,N_1363,N_1367);
and U2136 (N_2136,N_1562,N_1274);
and U2137 (N_2137,N_1526,N_1796);
nor U2138 (N_2138,N_1610,N_1746);
or U2139 (N_2139,N_1508,N_1513);
or U2140 (N_2140,N_1232,N_1254);
and U2141 (N_2141,N_1247,N_1668);
or U2142 (N_2142,N_1472,N_1482);
xnor U2143 (N_2143,N_1221,N_1376);
and U2144 (N_2144,N_1262,N_1496);
and U2145 (N_2145,N_1669,N_1701);
nand U2146 (N_2146,N_1716,N_1446);
or U2147 (N_2147,N_1368,N_1259);
nand U2148 (N_2148,N_1582,N_1538);
or U2149 (N_2149,N_1203,N_1218);
and U2150 (N_2150,N_1748,N_1746);
nor U2151 (N_2151,N_1217,N_1269);
xnor U2152 (N_2152,N_1627,N_1441);
or U2153 (N_2153,N_1216,N_1713);
and U2154 (N_2154,N_1584,N_1780);
nor U2155 (N_2155,N_1395,N_1543);
xnor U2156 (N_2156,N_1634,N_1351);
xor U2157 (N_2157,N_1259,N_1353);
and U2158 (N_2158,N_1466,N_1490);
or U2159 (N_2159,N_1678,N_1294);
and U2160 (N_2160,N_1498,N_1601);
nand U2161 (N_2161,N_1345,N_1744);
nor U2162 (N_2162,N_1233,N_1406);
xor U2163 (N_2163,N_1649,N_1539);
nor U2164 (N_2164,N_1439,N_1458);
xor U2165 (N_2165,N_1451,N_1468);
or U2166 (N_2166,N_1723,N_1588);
nor U2167 (N_2167,N_1275,N_1779);
xnor U2168 (N_2168,N_1343,N_1738);
xnor U2169 (N_2169,N_1301,N_1222);
xor U2170 (N_2170,N_1638,N_1293);
or U2171 (N_2171,N_1236,N_1481);
nor U2172 (N_2172,N_1716,N_1625);
or U2173 (N_2173,N_1223,N_1402);
or U2174 (N_2174,N_1617,N_1543);
xnor U2175 (N_2175,N_1642,N_1619);
xnor U2176 (N_2176,N_1354,N_1725);
xor U2177 (N_2177,N_1287,N_1659);
and U2178 (N_2178,N_1678,N_1448);
nand U2179 (N_2179,N_1656,N_1661);
and U2180 (N_2180,N_1605,N_1549);
and U2181 (N_2181,N_1383,N_1225);
nor U2182 (N_2182,N_1488,N_1443);
or U2183 (N_2183,N_1610,N_1390);
or U2184 (N_2184,N_1564,N_1758);
nand U2185 (N_2185,N_1307,N_1568);
or U2186 (N_2186,N_1732,N_1424);
or U2187 (N_2187,N_1582,N_1384);
or U2188 (N_2188,N_1630,N_1443);
and U2189 (N_2189,N_1513,N_1543);
and U2190 (N_2190,N_1275,N_1553);
xnor U2191 (N_2191,N_1461,N_1741);
and U2192 (N_2192,N_1682,N_1319);
or U2193 (N_2193,N_1544,N_1214);
nor U2194 (N_2194,N_1278,N_1454);
nor U2195 (N_2195,N_1736,N_1637);
and U2196 (N_2196,N_1449,N_1337);
or U2197 (N_2197,N_1468,N_1283);
and U2198 (N_2198,N_1301,N_1787);
nor U2199 (N_2199,N_1386,N_1253);
and U2200 (N_2200,N_1690,N_1302);
nand U2201 (N_2201,N_1435,N_1226);
or U2202 (N_2202,N_1484,N_1784);
xnor U2203 (N_2203,N_1711,N_1700);
and U2204 (N_2204,N_1589,N_1323);
xor U2205 (N_2205,N_1542,N_1519);
xor U2206 (N_2206,N_1411,N_1247);
nand U2207 (N_2207,N_1470,N_1747);
and U2208 (N_2208,N_1468,N_1694);
xor U2209 (N_2209,N_1768,N_1244);
xor U2210 (N_2210,N_1257,N_1789);
or U2211 (N_2211,N_1328,N_1336);
nand U2212 (N_2212,N_1205,N_1316);
nand U2213 (N_2213,N_1639,N_1352);
xor U2214 (N_2214,N_1581,N_1597);
xor U2215 (N_2215,N_1381,N_1542);
nor U2216 (N_2216,N_1247,N_1473);
and U2217 (N_2217,N_1242,N_1776);
and U2218 (N_2218,N_1445,N_1329);
and U2219 (N_2219,N_1268,N_1636);
or U2220 (N_2220,N_1410,N_1389);
or U2221 (N_2221,N_1251,N_1721);
nand U2222 (N_2222,N_1234,N_1458);
and U2223 (N_2223,N_1736,N_1440);
or U2224 (N_2224,N_1507,N_1362);
and U2225 (N_2225,N_1252,N_1246);
and U2226 (N_2226,N_1369,N_1218);
or U2227 (N_2227,N_1217,N_1434);
nor U2228 (N_2228,N_1425,N_1317);
xor U2229 (N_2229,N_1253,N_1565);
nor U2230 (N_2230,N_1375,N_1289);
nor U2231 (N_2231,N_1434,N_1432);
and U2232 (N_2232,N_1221,N_1605);
nand U2233 (N_2233,N_1398,N_1588);
and U2234 (N_2234,N_1545,N_1684);
xnor U2235 (N_2235,N_1408,N_1731);
nor U2236 (N_2236,N_1460,N_1348);
nand U2237 (N_2237,N_1434,N_1693);
or U2238 (N_2238,N_1316,N_1566);
and U2239 (N_2239,N_1302,N_1691);
and U2240 (N_2240,N_1343,N_1261);
nand U2241 (N_2241,N_1202,N_1640);
nand U2242 (N_2242,N_1782,N_1573);
and U2243 (N_2243,N_1610,N_1310);
or U2244 (N_2244,N_1762,N_1647);
xor U2245 (N_2245,N_1268,N_1495);
xnor U2246 (N_2246,N_1406,N_1555);
nor U2247 (N_2247,N_1602,N_1581);
nand U2248 (N_2248,N_1703,N_1709);
nor U2249 (N_2249,N_1217,N_1681);
or U2250 (N_2250,N_1201,N_1422);
nand U2251 (N_2251,N_1480,N_1473);
xnor U2252 (N_2252,N_1680,N_1560);
or U2253 (N_2253,N_1341,N_1548);
or U2254 (N_2254,N_1666,N_1715);
nor U2255 (N_2255,N_1459,N_1461);
nor U2256 (N_2256,N_1533,N_1598);
and U2257 (N_2257,N_1672,N_1507);
nor U2258 (N_2258,N_1540,N_1567);
and U2259 (N_2259,N_1688,N_1612);
nor U2260 (N_2260,N_1360,N_1348);
nand U2261 (N_2261,N_1245,N_1597);
xnor U2262 (N_2262,N_1518,N_1612);
xnor U2263 (N_2263,N_1645,N_1740);
or U2264 (N_2264,N_1349,N_1553);
xor U2265 (N_2265,N_1639,N_1578);
xor U2266 (N_2266,N_1444,N_1631);
nor U2267 (N_2267,N_1438,N_1229);
nor U2268 (N_2268,N_1625,N_1510);
nand U2269 (N_2269,N_1411,N_1432);
xor U2270 (N_2270,N_1272,N_1387);
nor U2271 (N_2271,N_1743,N_1565);
or U2272 (N_2272,N_1231,N_1628);
xnor U2273 (N_2273,N_1760,N_1428);
xor U2274 (N_2274,N_1653,N_1204);
nand U2275 (N_2275,N_1364,N_1233);
xor U2276 (N_2276,N_1360,N_1329);
nand U2277 (N_2277,N_1511,N_1737);
and U2278 (N_2278,N_1624,N_1393);
or U2279 (N_2279,N_1389,N_1717);
xor U2280 (N_2280,N_1668,N_1474);
nor U2281 (N_2281,N_1693,N_1785);
nand U2282 (N_2282,N_1441,N_1261);
nor U2283 (N_2283,N_1738,N_1634);
nand U2284 (N_2284,N_1751,N_1367);
and U2285 (N_2285,N_1684,N_1410);
xnor U2286 (N_2286,N_1287,N_1631);
nand U2287 (N_2287,N_1467,N_1767);
xor U2288 (N_2288,N_1446,N_1220);
nand U2289 (N_2289,N_1286,N_1453);
or U2290 (N_2290,N_1340,N_1266);
nand U2291 (N_2291,N_1564,N_1244);
xor U2292 (N_2292,N_1330,N_1558);
or U2293 (N_2293,N_1786,N_1234);
or U2294 (N_2294,N_1467,N_1379);
xnor U2295 (N_2295,N_1324,N_1252);
nor U2296 (N_2296,N_1757,N_1541);
xnor U2297 (N_2297,N_1631,N_1699);
and U2298 (N_2298,N_1626,N_1270);
and U2299 (N_2299,N_1472,N_1718);
nand U2300 (N_2300,N_1466,N_1651);
nand U2301 (N_2301,N_1522,N_1349);
nor U2302 (N_2302,N_1690,N_1585);
nand U2303 (N_2303,N_1596,N_1745);
nand U2304 (N_2304,N_1258,N_1320);
and U2305 (N_2305,N_1771,N_1718);
or U2306 (N_2306,N_1293,N_1543);
nand U2307 (N_2307,N_1467,N_1699);
and U2308 (N_2308,N_1545,N_1422);
and U2309 (N_2309,N_1555,N_1721);
nor U2310 (N_2310,N_1671,N_1783);
or U2311 (N_2311,N_1707,N_1706);
xnor U2312 (N_2312,N_1619,N_1663);
and U2313 (N_2313,N_1506,N_1611);
nor U2314 (N_2314,N_1569,N_1273);
nor U2315 (N_2315,N_1262,N_1794);
nand U2316 (N_2316,N_1639,N_1571);
nor U2317 (N_2317,N_1562,N_1666);
and U2318 (N_2318,N_1785,N_1707);
xor U2319 (N_2319,N_1746,N_1245);
xnor U2320 (N_2320,N_1238,N_1437);
and U2321 (N_2321,N_1772,N_1549);
or U2322 (N_2322,N_1302,N_1539);
and U2323 (N_2323,N_1449,N_1535);
nor U2324 (N_2324,N_1727,N_1710);
nand U2325 (N_2325,N_1605,N_1798);
nor U2326 (N_2326,N_1792,N_1507);
nand U2327 (N_2327,N_1300,N_1710);
and U2328 (N_2328,N_1286,N_1527);
or U2329 (N_2329,N_1417,N_1633);
xor U2330 (N_2330,N_1647,N_1597);
nor U2331 (N_2331,N_1741,N_1229);
xor U2332 (N_2332,N_1632,N_1672);
or U2333 (N_2333,N_1602,N_1492);
or U2334 (N_2334,N_1748,N_1544);
nor U2335 (N_2335,N_1623,N_1352);
or U2336 (N_2336,N_1445,N_1509);
and U2337 (N_2337,N_1284,N_1780);
nand U2338 (N_2338,N_1788,N_1338);
xnor U2339 (N_2339,N_1525,N_1513);
nor U2340 (N_2340,N_1252,N_1332);
or U2341 (N_2341,N_1227,N_1638);
or U2342 (N_2342,N_1428,N_1465);
xnor U2343 (N_2343,N_1604,N_1288);
or U2344 (N_2344,N_1365,N_1305);
and U2345 (N_2345,N_1299,N_1705);
nor U2346 (N_2346,N_1687,N_1373);
nand U2347 (N_2347,N_1248,N_1686);
or U2348 (N_2348,N_1282,N_1751);
nand U2349 (N_2349,N_1684,N_1626);
and U2350 (N_2350,N_1539,N_1505);
nor U2351 (N_2351,N_1622,N_1550);
nor U2352 (N_2352,N_1414,N_1552);
xor U2353 (N_2353,N_1532,N_1356);
nand U2354 (N_2354,N_1352,N_1643);
nand U2355 (N_2355,N_1621,N_1722);
nand U2356 (N_2356,N_1358,N_1298);
nand U2357 (N_2357,N_1763,N_1259);
or U2358 (N_2358,N_1656,N_1465);
xnor U2359 (N_2359,N_1357,N_1769);
xor U2360 (N_2360,N_1206,N_1363);
nand U2361 (N_2361,N_1275,N_1205);
nor U2362 (N_2362,N_1269,N_1466);
or U2363 (N_2363,N_1606,N_1501);
and U2364 (N_2364,N_1780,N_1575);
xor U2365 (N_2365,N_1489,N_1520);
nand U2366 (N_2366,N_1585,N_1625);
or U2367 (N_2367,N_1289,N_1607);
nor U2368 (N_2368,N_1424,N_1205);
and U2369 (N_2369,N_1724,N_1441);
and U2370 (N_2370,N_1269,N_1442);
xnor U2371 (N_2371,N_1568,N_1646);
xnor U2372 (N_2372,N_1474,N_1579);
or U2373 (N_2373,N_1670,N_1328);
or U2374 (N_2374,N_1263,N_1412);
nor U2375 (N_2375,N_1203,N_1566);
nand U2376 (N_2376,N_1544,N_1503);
nor U2377 (N_2377,N_1506,N_1742);
and U2378 (N_2378,N_1778,N_1319);
and U2379 (N_2379,N_1525,N_1226);
or U2380 (N_2380,N_1737,N_1770);
nor U2381 (N_2381,N_1625,N_1717);
or U2382 (N_2382,N_1543,N_1498);
or U2383 (N_2383,N_1317,N_1269);
or U2384 (N_2384,N_1753,N_1315);
nand U2385 (N_2385,N_1463,N_1649);
nand U2386 (N_2386,N_1498,N_1680);
nor U2387 (N_2387,N_1258,N_1750);
or U2388 (N_2388,N_1323,N_1594);
nor U2389 (N_2389,N_1593,N_1227);
xor U2390 (N_2390,N_1608,N_1654);
or U2391 (N_2391,N_1771,N_1282);
nand U2392 (N_2392,N_1716,N_1276);
xor U2393 (N_2393,N_1222,N_1288);
nor U2394 (N_2394,N_1496,N_1507);
or U2395 (N_2395,N_1583,N_1579);
nand U2396 (N_2396,N_1311,N_1475);
nor U2397 (N_2397,N_1691,N_1399);
nor U2398 (N_2398,N_1366,N_1574);
and U2399 (N_2399,N_1475,N_1686);
xor U2400 (N_2400,N_1977,N_2087);
or U2401 (N_2401,N_1917,N_2130);
nor U2402 (N_2402,N_1848,N_1942);
or U2403 (N_2403,N_2330,N_2394);
xor U2404 (N_2404,N_2154,N_2344);
nand U2405 (N_2405,N_1924,N_2237);
nor U2406 (N_2406,N_1934,N_2262);
xor U2407 (N_2407,N_2263,N_2086);
nand U2408 (N_2408,N_2239,N_2260);
xor U2409 (N_2409,N_1935,N_2001);
and U2410 (N_2410,N_2010,N_2080);
nand U2411 (N_2411,N_1945,N_1998);
nand U2412 (N_2412,N_2204,N_1810);
nor U2413 (N_2413,N_2186,N_2279);
xor U2414 (N_2414,N_2129,N_2090);
nor U2415 (N_2415,N_2385,N_2377);
nand U2416 (N_2416,N_1939,N_2210);
or U2417 (N_2417,N_1954,N_2399);
or U2418 (N_2418,N_2326,N_2290);
nor U2419 (N_2419,N_2347,N_1873);
and U2420 (N_2420,N_2067,N_2276);
nand U2421 (N_2421,N_2142,N_2048);
xnor U2422 (N_2422,N_1824,N_2144);
xnor U2423 (N_2423,N_2302,N_1883);
or U2424 (N_2424,N_1807,N_2157);
or U2425 (N_2425,N_2216,N_2065);
or U2426 (N_2426,N_2228,N_1811);
nand U2427 (N_2427,N_2307,N_1949);
xor U2428 (N_2428,N_2343,N_1843);
nor U2429 (N_2429,N_2119,N_2208);
and U2430 (N_2430,N_2238,N_1878);
or U2431 (N_2431,N_2245,N_1813);
xnor U2432 (N_2432,N_1832,N_2059);
nor U2433 (N_2433,N_2299,N_2350);
or U2434 (N_2434,N_2259,N_2166);
xor U2435 (N_2435,N_2085,N_1845);
nand U2436 (N_2436,N_2063,N_2207);
xnor U2437 (N_2437,N_2200,N_2380);
or U2438 (N_2438,N_1879,N_2281);
and U2439 (N_2439,N_2220,N_2012);
or U2440 (N_2440,N_2098,N_1896);
and U2441 (N_2441,N_1973,N_2134);
xnor U2442 (N_2442,N_1978,N_2387);
xor U2443 (N_2443,N_2293,N_2179);
and U2444 (N_2444,N_2064,N_1950);
xor U2445 (N_2445,N_2390,N_2247);
nor U2446 (N_2446,N_2317,N_2004);
xnor U2447 (N_2447,N_2122,N_2389);
or U2448 (N_2448,N_2248,N_1804);
nor U2449 (N_2449,N_2155,N_2329);
xnor U2450 (N_2450,N_2391,N_2163);
or U2451 (N_2451,N_2335,N_2043);
or U2452 (N_2452,N_2363,N_2088);
nor U2453 (N_2453,N_2214,N_1927);
nand U2454 (N_2454,N_2374,N_2131);
xnor U2455 (N_2455,N_2147,N_2211);
nor U2456 (N_2456,N_1850,N_2309);
and U2457 (N_2457,N_1818,N_1836);
or U2458 (N_2458,N_2274,N_2023);
or U2459 (N_2459,N_2174,N_2139);
or U2460 (N_2460,N_2325,N_2320);
nand U2461 (N_2461,N_2075,N_2256);
nor U2462 (N_2462,N_1864,N_2049);
nor U2463 (N_2463,N_1961,N_2189);
and U2464 (N_2464,N_1969,N_1964);
or U2465 (N_2465,N_2272,N_1853);
xor U2466 (N_2466,N_2355,N_2244);
or U2467 (N_2467,N_2145,N_2013);
or U2468 (N_2468,N_2046,N_2252);
xor U2469 (N_2469,N_2255,N_2103);
nor U2470 (N_2470,N_1892,N_2162);
nor U2471 (N_2471,N_2017,N_2352);
xor U2472 (N_2472,N_1870,N_2342);
nor U2473 (N_2473,N_2068,N_2025);
and U2474 (N_2474,N_2108,N_2002);
nand U2475 (N_2475,N_2183,N_2106);
nand U2476 (N_2476,N_2036,N_1971);
and U2477 (N_2477,N_2303,N_1840);
or U2478 (N_2478,N_2124,N_2097);
nand U2479 (N_2479,N_1923,N_2288);
nor U2480 (N_2480,N_2202,N_2104);
nand U2481 (N_2481,N_2327,N_2198);
nor U2482 (N_2482,N_2366,N_2304);
and U2483 (N_2483,N_1842,N_2125);
nor U2484 (N_2484,N_2242,N_2332);
xnor U2485 (N_2485,N_2024,N_1898);
xnor U2486 (N_2486,N_2072,N_2322);
and U2487 (N_2487,N_2146,N_2267);
nand U2488 (N_2488,N_2345,N_2209);
xnor U2489 (N_2489,N_1865,N_1869);
or U2490 (N_2490,N_1839,N_2339);
xnor U2491 (N_2491,N_1893,N_1930);
nand U2492 (N_2492,N_2213,N_2081);
nand U2493 (N_2493,N_1966,N_2037);
or U2494 (N_2494,N_1970,N_2235);
xnor U2495 (N_2495,N_1905,N_2061);
nor U2496 (N_2496,N_2315,N_1863);
xnor U2497 (N_2497,N_2176,N_1963);
or U2498 (N_2498,N_1929,N_2082);
nand U2499 (N_2499,N_1981,N_1991);
xnor U2500 (N_2500,N_2027,N_2045);
xor U2501 (N_2501,N_1861,N_2378);
or U2502 (N_2502,N_2319,N_2221);
and U2503 (N_2503,N_2365,N_2234);
or U2504 (N_2504,N_2253,N_1936);
nand U2505 (N_2505,N_2133,N_2201);
xnor U2506 (N_2506,N_2241,N_1874);
xnor U2507 (N_2507,N_2052,N_2051);
xnor U2508 (N_2508,N_2160,N_2386);
or U2509 (N_2509,N_2019,N_2392);
nor U2510 (N_2510,N_2184,N_2101);
xor U2511 (N_2511,N_1938,N_2148);
nand U2512 (N_2512,N_1837,N_2055);
nand U2513 (N_2513,N_2218,N_2217);
nor U2514 (N_2514,N_1829,N_1925);
nor U2515 (N_2515,N_2398,N_2128);
and U2516 (N_2516,N_2312,N_1996);
nor U2517 (N_2517,N_2257,N_2269);
and U2518 (N_2518,N_1812,N_2136);
or U2519 (N_2519,N_1986,N_1826);
nor U2520 (N_2520,N_2215,N_2300);
nor U2521 (N_2521,N_2289,N_2324);
or U2522 (N_2522,N_1851,N_1994);
nand U2523 (N_2523,N_1830,N_1984);
nand U2524 (N_2524,N_2323,N_1989);
or U2525 (N_2525,N_2178,N_1946);
and U2526 (N_2526,N_1867,N_2219);
or U2527 (N_2527,N_1844,N_2268);
and U2528 (N_2528,N_2192,N_2029);
nand U2529 (N_2529,N_1899,N_1907);
and U2530 (N_2530,N_2314,N_2137);
nor U2531 (N_2531,N_2156,N_2000);
nand U2532 (N_2532,N_2318,N_2250);
nand U2533 (N_2533,N_2271,N_1968);
nor U2534 (N_2534,N_2116,N_2368);
or U2535 (N_2535,N_2190,N_1992);
nand U2536 (N_2536,N_2076,N_2354);
nand U2537 (N_2537,N_1814,N_2038);
nor U2538 (N_2538,N_2197,N_2328);
and U2539 (N_2539,N_2351,N_2285);
nand U2540 (N_2540,N_2138,N_1862);
xor U2541 (N_2541,N_2275,N_2341);
xnor U2542 (N_2542,N_1831,N_2287);
nand U2543 (N_2543,N_2100,N_2305);
nor U2544 (N_2544,N_2346,N_2032);
xnor U2545 (N_2545,N_2383,N_1955);
nor U2546 (N_2546,N_1957,N_2353);
or U2547 (N_2547,N_1941,N_2236);
nor U2548 (N_2548,N_1904,N_1900);
or U2549 (N_2549,N_1960,N_2294);
nand U2550 (N_2550,N_2270,N_1965);
nor U2551 (N_2551,N_2077,N_2246);
and U2552 (N_2552,N_2396,N_1920);
xor U2553 (N_2553,N_2232,N_2360);
nor U2554 (N_2554,N_1889,N_1884);
or U2555 (N_2555,N_1952,N_1858);
nand U2556 (N_2556,N_2071,N_2127);
nand U2557 (N_2557,N_2170,N_1913);
nor U2558 (N_2558,N_2140,N_2376);
and U2559 (N_2559,N_2056,N_1909);
and U2560 (N_2560,N_1866,N_1816);
nor U2561 (N_2561,N_2397,N_2364);
or U2562 (N_2562,N_2298,N_2371);
xnor U2563 (N_2563,N_2313,N_1922);
nor U2564 (N_2564,N_2028,N_2308);
xnor U2565 (N_2565,N_2135,N_1958);
xor U2566 (N_2566,N_2044,N_2333);
and U2567 (N_2567,N_2132,N_2181);
nand U2568 (N_2568,N_1979,N_2243);
nand U2569 (N_2569,N_1895,N_2338);
and U2570 (N_2570,N_2062,N_2282);
and U2571 (N_2571,N_1849,N_1983);
nor U2572 (N_2572,N_1805,N_2011);
or U2573 (N_2573,N_2393,N_2277);
nand U2574 (N_2574,N_1821,N_2151);
or U2575 (N_2575,N_2054,N_2283);
nand U2576 (N_2576,N_2362,N_1817);
xor U2577 (N_2577,N_1856,N_2379);
or U2578 (N_2578,N_2005,N_2167);
and U2579 (N_2579,N_2331,N_2286);
or U2580 (N_2580,N_2105,N_2370);
nand U2581 (N_2581,N_2018,N_2030);
nor U2582 (N_2582,N_2382,N_1921);
or U2583 (N_2583,N_2336,N_2016);
xnor U2584 (N_2584,N_2278,N_2251);
xor U2585 (N_2585,N_2224,N_2079);
and U2586 (N_2586,N_2060,N_1823);
nand U2587 (N_2587,N_2117,N_2008);
nand U2588 (N_2588,N_2310,N_1902);
nand U2589 (N_2589,N_1891,N_2053);
nand U2590 (N_2590,N_2265,N_2089);
or U2591 (N_2591,N_1872,N_2057);
xnor U2592 (N_2592,N_1852,N_2058);
and U2593 (N_2593,N_1887,N_2375);
nand U2594 (N_2594,N_2042,N_1997);
nor U2595 (N_2595,N_2115,N_2091);
or U2596 (N_2596,N_2111,N_2113);
nand U2597 (N_2597,N_2047,N_2143);
and U2598 (N_2598,N_2205,N_2357);
nand U2599 (N_2599,N_2112,N_2007);
or U2600 (N_2600,N_1901,N_2195);
and U2601 (N_2601,N_2123,N_2171);
and U2602 (N_2602,N_2280,N_1999);
nand U2603 (N_2603,N_2039,N_1841);
xnor U2604 (N_2604,N_2034,N_2295);
xor U2605 (N_2605,N_1916,N_2165);
xor U2606 (N_2606,N_1912,N_1886);
nand U2607 (N_2607,N_2191,N_2040);
nor U2608 (N_2608,N_1882,N_2321);
and U2609 (N_2609,N_1855,N_1988);
nand U2610 (N_2610,N_1894,N_1985);
nor U2611 (N_2611,N_2297,N_1933);
nand U2612 (N_2612,N_2388,N_2153);
nand U2613 (N_2613,N_1990,N_1888);
or U2614 (N_2614,N_1833,N_2381);
nand U2615 (N_2615,N_2227,N_1803);
or U2616 (N_2616,N_1835,N_2070);
nor U2617 (N_2617,N_2340,N_2296);
nand U2618 (N_2618,N_1914,N_2222);
xnor U2619 (N_2619,N_1806,N_1975);
or U2620 (N_2620,N_2206,N_2121);
nand U2621 (N_2621,N_2229,N_2150);
nor U2622 (N_2622,N_2021,N_2110);
nor U2623 (N_2623,N_1908,N_2126);
and U2624 (N_2624,N_2020,N_2284);
xor U2625 (N_2625,N_2050,N_2177);
or U2626 (N_2626,N_2369,N_2026);
nor U2627 (N_2627,N_2006,N_1932);
nor U2628 (N_2628,N_2022,N_2182);
and U2629 (N_2629,N_1911,N_2266);
nand U2630 (N_2630,N_2014,N_2033);
nand U2631 (N_2631,N_2273,N_2009);
nor U2632 (N_2632,N_2003,N_1974);
nand U2633 (N_2633,N_1982,N_2095);
and U2634 (N_2634,N_2372,N_2031);
and U2635 (N_2635,N_2169,N_2083);
or U2636 (N_2636,N_1819,N_2301);
xnor U2637 (N_2637,N_2141,N_2258);
and U2638 (N_2638,N_2194,N_2196);
or U2639 (N_2639,N_1903,N_2212);
or U2640 (N_2640,N_2102,N_2384);
nand U2641 (N_2641,N_2074,N_1822);
nand U2642 (N_2642,N_2172,N_2373);
nand U2643 (N_2643,N_2069,N_2306);
nand U2644 (N_2644,N_2118,N_1834);
nand U2645 (N_2645,N_1838,N_2225);
and U2646 (N_2646,N_1802,N_2264);
nor U2647 (N_2647,N_1995,N_1815);
nor U2648 (N_2648,N_2161,N_1915);
xnor U2649 (N_2649,N_1890,N_2231);
or U2650 (N_2650,N_1947,N_1940);
and U2651 (N_2651,N_1881,N_2249);
nor U2652 (N_2652,N_1828,N_1868);
nor U2653 (N_2653,N_2254,N_1987);
nand U2654 (N_2654,N_2316,N_2120);
xor U2655 (N_2655,N_1919,N_2092);
and U2656 (N_2656,N_1897,N_1962);
or U2657 (N_2657,N_2168,N_1993);
xnor U2658 (N_2658,N_1820,N_2187);
xnor U2659 (N_2659,N_2164,N_2015);
nand U2660 (N_2660,N_2078,N_2152);
nor U2661 (N_2661,N_1808,N_2096);
or U2662 (N_2662,N_2223,N_1800);
xor U2663 (N_2663,N_1967,N_2073);
xnor U2664 (N_2664,N_1825,N_1847);
nor U2665 (N_2665,N_1931,N_2159);
nand U2666 (N_2666,N_2180,N_1976);
nor U2667 (N_2667,N_2292,N_2084);
or U2668 (N_2668,N_2114,N_2185);
and U2669 (N_2669,N_2173,N_2041);
nor U2670 (N_2670,N_2107,N_1943);
and U2671 (N_2671,N_2367,N_1801);
xnor U2672 (N_2672,N_1880,N_2226);
or U2673 (N_2673,N_1959,N_2158);
and U2674 (N_2674,N_1875,N_1885);
and U2675 (N_2675,N_1871,N_2199);
and U2676 (N_2676,N_1910,N_1846);
nand U2677 (N_2677,N_2035,N_1980);
nand U2678 (N_2678,N_2356,N_1809);
and U2679 (N_2679,N_2334,N_1953);
nor U2680 (N_2680,N_1876,N_1951);
and U2681 (N_2681,N_2149,N_1877);
nand U2682 (N_2682,N_2337,N_2230);
xnor U2683 (N_2683,N_1906,N_2348);
and U2684 (N_2684,N_1854,N_1859);
nand U2685 (N_2685,N_2094,N_1937);
nor U2686 (N_2686,N_1956,N_1944);
or U2687 (N_2687,N_1928,N_1972);
nor U2688 (N_2688,N_1948,N_2240);
xnor U2689 (N_2689,N_2066,N_2311);
nor U2690 (N_2690,N_2233,N_2261);
and U2691 (N_2691,N_2099,N_1827);
and U2692 (N_2692,N_2358,N_2359);
xnor U2693 (N_2693,N_2395,N_1860);
and U2694 (N_2694,N_2175,N_2291);
or U2695 (N_2695,N_2188,N_2349);
and U2696 (N_2696,N_2109,N_1926);
and U2697 (N_2697,N_2193,N_1918);
nor U2698 (N_2698,N_2361,N_1857);
xor U2699 (N_2699,N_2093,N_2203);
xor U2700 (N_2700,N_2345,N_1878);
xnor U2701 (N_2701,N_2248,N_2216);
and U2702 (N_2702,N_2065,N_1815);
xnor U2703 (N_2703,N_1839,N_2353);
or U2704 (N_2704,N_2051,N_2275);
or U2705 (N_2705,N_1882,N_2098);
nor U2706 (N_2706,N_1934,N_2169);
or U2707 (N_2707,N_2016,N_2383);
and U2708 (N_2708,N_2028,N_1874);
nor U2709 (N_2709,N_1875,N_2349);
xor U2710 (N_2710,N_2175,N_1944);
nor U2711 (N_2711,N_1952,N_2311);
xnor U2712 (N_2712,N_1883,N_2116);
or U2713 (N_2713,N_2112,N_2236);
nand U2714 (N_2714,N_2055,N_2111);
and U2715 (N_2715,N_2033,N_2000);
and U2716 (N_2716,N_2268,N_2170);
nand U2717 (N_2717,N_2302,N_2029);
nand U2718 (N_2718,N_2296,N_2355);
nor U2719 (N_2719,N_2264,N_1883);
nand U2720 (N_2720,N_2272,N_1884);
or U2721 (N_2721,N_1809,N_2120);
or U2722 (N_2722,N_1836,N_1844);
and U2723 (N_2723,N_2392,N_1914);
nand U2724 (N_2724,N_2181,N_1946);
xnor U2725 (N_2725,N_1860,N_1835);
nand U2726 (N_2726,N_1992,N_1962);
nor U2727 (N_2727,N_2066,N_2218);
nand U2728 (N_2728,N_1823,N_2082);
or U2729 (N_2729,N_2222,N_2362);
nor U2730 (N_2730,N_1982,N_1895);
or U2731 (N_2731,N_1951,N_2129);
nand U2732 (N_2732,N_1972,N_2265);
xnor U2733 (N_2733,N_2318,N_1887);
or U2734 (N_2734,N_1886,N_2159);
and U2735 (N_2735,N_1999,N_2348);
nor U2736 (N_2736,N_2227,N_2009);
xnor U2737 (N_2737,N_2215,N_2152);
nand U2738 (N_2738,N_1827,N_2081);
nand U2739 (N_2739,N_2398,N_2177);
nor U2740 (N_2740,N_2104,N_1912);
xnor U2741 (N_2741,N_2365,N_2141);
or U2742 (N_2742,N_2197,N_1972);
or U2743 (N_2743,N_1803,N_2142);
nor U2744 (N_2744,N_2284,N_2062);
or U2745 (N_2745,N_2276,N_1943);
nor U2746 (N_2746,N_2376,N_2182);
and U2747 (N_2747,N_2203,N_1806);
or U2748 (N_2748,N_2288,N_1849);
xor U2749 (N_2749,N_2160,N_2038);
and U2750 (N_2750,N_2197,N_1942);
or U2751 (N_2751,N_2318,N_2133);
nor U2752 (N_2752,N_1863,N_2307);
nand U2753 (N_2753,N_1929,N_2354);
nor U2754 (N_2754,N_1817,N_2181);
nor U2755 (N_2755,N_2115,N_1961);
nand U2756 (N_2756,N_2211,N_1867);
nor U2757 (N_2757,N_1807,N_2130);
nand U2758 (N_2758,N_2040,N_2184);
nor U2759 (N_2759,N_2272,N_1934);
nor U2760 (N_2760,N_2395,N_1847);
xnor U2761 (N_2761,N_2122,N_2322);
nor U2762 (N_2762,N_2218,N_2255);
nor U2763 (N_2763,N_1842,N_2024);
nor U2764 (N_2764,N_1869,N_2308);
and U2765 (N_2765,N_2276,N_1953);
and U2766 (N_2766,N_2383,N_1896);
or U2767 (N_2767,N_2169,N_1863);
and U2768 (N_2768,N_2190,N_2183);
nand U2769 (N_2769,N_1930,N_1857);
nor U2770 (N_2770,N_1998,N_1983);
nand U2771 (N_2771,N_2374,N_2301);
nand U2772 (N_2772,N_2246,N_1823);
nor U2773 (N_2773,N_2194,N_2389);
or U2774 (N_2774,N_1866,N_1915);
or U2775 (N_2775,N_2213,N_1858);
nand U2776 (N_2776,N_1940,N_2312);
nand U2777 (N_2777,N_2157,N_2214);
xor U2778 (N_2778,N_2254,N_2386);
nor U2779 (N_2779,N_2393,N_2170);
xnor U2780 (N_2780,N_1984,N_2186);
nand U2781 (N_2781,N_2342,N_2227);
nand U2782 (N_2782,N_2181,N_1825);
nand U2783 (N_2783,N_2093,N_2198);
nor U2784 (N_2784,N_2273,N_2293);
nor U2785 (N_2785,N_2254,N_1951);
nor U2786 (N_2786,N_2165,N_2071);
xor U2787 (N_2787,N_1818,N_2050);
nand U2788 (N_2788,N_2012,N_2047);
nand U2789 (N_2789,N_2131,N_2014);
xnor U2790 (N_2790,N_1880,N_2256);
xnor U2791 (N_2791,N_2379,N_1836);
nor U2792 (N_2792,N_2127,N_2162);
nand U2793 (N_2793,N_1981,N_2147);
nand U2794 (N_2794,N_1852,N_2026);
or U2795 (N_2795,N_1984,N_1824);
xnor U2796 (N_2796,N_2072,N_1866);
xnor U2797 (N_2797,N_1886,N_1849);
and U2798 (N_2798,N_2033,N_1927);
or U2799 (N_2799,N_2176,N_2220);
nor U2800 (N_2800,N_1963,N_2261);
and U2801 (N_2801,N_1951,N_2212);
or U2802 (N_2802,N_1819,N_2117);
or U2803 (N_2803,N_1976,N_2124);
or U2804 (N_2804,N_2300,N_1944);
nor U2805 (N_2805,N_1852,N_1925);
xor U2806 (N_2806,N_2039,N_1891);
or U2807 (N_2807,N_2218,N_2271);
nand U2808 (N_2808,N_2353,N_2357);
xor U2809 (N_2809,N_1977,N_1800);
nor U2810 (N_2810,N_2020,N_2361);
and U2811 (N_2811,N_1998,N_2359);
and U2812 (N_2812,N_2050,N_2290);
nand U2813 (N_2813,N_1920,N_2386);
or U2814 (N_2814,N_2171,N_2178);
nor U2815 (N_2815,N_2086,N_2262);
or U2816 (N_2816,N_1998,N_2283);
nor U2817 (N_2817,N_2191,N_1960);
or U2818 (N_2818,N_1989,N_1970);
nor U2819 (N_2819,N_2226,N_1955);
or U2820 (N_2820,N_1871,N_1894);
and U2821 (N_2821,N_1878,N_1949);
nand U2822 (N_2822,N_2116,N_2279);
or U2823 (N_2823,N_1924,N_2317);
xnor U2824 (N_2824,N_2316,N_2038);
xnor U2825 (N_2825,N_2006,N_2097);
xnor U2826 (N_2826,N_2190,N_1988);
or U2827 (N_2827,N_1849,N_2026);
nor U2828 (N_2828,N_2318,N_2043);
and U2829 (N_2829,N_1969,N_2148);
and U2830 (N_2830,N_2314,N_2074);
or U2831 (N_2831,N_2042,N_2027);
and U2832 (N_2832,N_1978,N_2236);
nand U2833 (N_2833,N_1897,N_2060);
xnor U2834 (N_2834,N_2335,N_1926);
and U2835 (N_2835,N_1866,N_1833);
and U2836 (N_2836,N_2173,N_2009);
xnor U2837 (N_2837,N_2141,N_2394);
or U2838 (N_2838,N_1887,N_2177);
nor U2839 (N_2839,N_1859,N_1947);
nand U2840 (N_2840,N_2368,N_2259);
or U2841 (N_2841,N_2267,N_2334);
xnor U2842 (N_2842,N_2273,N_2343);
and U2843 (N_2843,N_2121,N_1848);
xor U2844 (N_2844,N_1849,N_2215);
nand U2845 (N_2845,N_2259,N_2360);
nand U2846 (N_2846,N_2084,N_1839);
and U2847 (N_2847,N_2227,N_2184);
nand U2848 (N_2848,N_1905,N_2057);
nor U2849 (N_2849,N_1829,N_1992);
xnor U2850 (N_2850,N_2060,N_1988);
xnor U2851 (N_2851,N_1991,N_1998);
nor U2852 (N_2852,N_2091,N_2049);
xor U2853 (N_2853,N_2203,N_1942);
or U2854 (N_2854,N_2258,N_2243);
or U2855 (N_2855,N_2192,N_2398);
nand U2856 (N_2856,N_2274,N_1998);
and U2857 (N_2857,N_2352,N_2201);
nand U2858 (N_2858,N_2390,N_2316);
nand U2859 (N_2859,N_2301,N_2054);
nand U2860 (N_2860,N_2170,N_2018);
xnor U2861 (N_2861,N_1903,N_2007);
or U2862 (N_2862,N_2290,N_1880);
nand U2863 (N_2863,N_2313,N_1859);
xnor U2864 (N_2864,N_2012,N_2163);
and U2865 (N_2865,N_2215,N_2263);
or U2866 (N_2866,N_2275,N_2371);
xnor U2867 (N_2867,N_2374,N_1817);
xor U2868 (N_2868,N_2154,N_2386);
or U2869 (N_2869,N_1851,N_2021);
and U2870 (N_2870,N_2249,N_2196);
or U2871 (N_2871,N_2326,N_2209);
xor U2872 (N_2872,N_1920,N_1912);
or U2873 (N_2873,N_2262,N_1819);
xnor U2874 (N_2874,N_1848,N_1832);
nor U2875 (N_2875,N_2345,N_2001);
xnor U2876 (N_2876,N_1947,N_2380);
xnor U2877 (N_2877,N_1972,N_2208);
nand U2878 (N_2878,N_1814,N_2332);
nor U2879 (N_2879,N_2152,N_1981);
or U2880 (N_2880,N_2329,N_2292);
xor U2881 (N_2881,N_2353,N_1928);
nor U2882 (N_2882,N_1960,N_2281);
nor U2883 (N_2883,N_2185,N_1841);
nand U2884 (N_2884,N_2124,N_1896);
xnor U2885 (N_2885,N_1946,N_2306);
or U2886 (N_2886,N_1922,N_2080);
or U2887 (N_2887,N_2136,N_1949);
xnor U2888 (N_2888,N_2270,N_2297);
nand U2889 (N_2889,N_2096,N_2224);
nand U2890 (N_2890,N_1840,N_1838);
or U2891 (N_2891,N_2169,N_2204);
nor U2892 (N_2892,N_1952,N_2300);
xnor U2893 (N_2893,N_1864,N_1868);
or U2894 (N_2894,N_2001,N_1809);
nand U2895 (N_2895,N_2235,N_2219);
or U2896 (N_2896,N_1845,N_1816);
nand U2897 (N_2897,N_2094,N_1830);
or U2898 (N_2898,N_2153,N_2267);
xnor U2899 (N_2899,N_2005,N_2279);
nand U2900 (N_2900,N_2339,N_2059);
nor U2901 (N_2901,N_1828,N_2128);
or U2902 (N_2902,N_2218,N_2227);
nand U2903 (N_2903,N_2247,N_2350);
or U2904 (N_2904,N_2360,N_2159);
and U2905 (N_2905,N_2335,N_2103);
nand U2906 (N_2906,N_2020,N_2129);
and U2907 (N_2907,N_2109,N_2225);
nor U2908 (N_2908,N_1855,N_1906);
or U2909 (N_2909,N_2232,N_1916);
xnor U2910 (N_2910,N_2036,N_1829);
xnor U2911 (N_2911,N_2167,N_1850);
nand U2912 (N_2912,N_2067,N_2394);
nand U2913 (N_2913,N_2045,N_1961);
nand U2914 (N_2914,N_2171,N_2311);
nor U2915 (N_2915,N_1837,N_2203);
or U2916 (N_2916,N_1924,N_1855);
and U2917 (N_2917,N_1816,N_2166);
nor U2918 (N_2918,N_2135,N_2149);
nand U2919 (N_2919,N_1838,N_2153);
nor U2920 (N_2920,N_1844,N_2315);
nor U2921 (N_2921,N_2031,N_2390);
nor U2922 (N_2922,N_2209,N_1806);
nand U2923 (N_2923,N_2007,N_1866);
or U2924 (N_2924,N_2272,N_2028);
and U2925 (N_2925,N_1857,N_2082);
xor U2926 (N_2926,N_2286,N_2239);
nand U2927 (N_2927,N_2153,N_2082);
or U2928 (N_2928,N_2040,N_2000);
or U2929 (N_2929,N_1841,N_1990);
xnor U2930 (N_2930,N_1927,N_2074);
and U2931 (N_2931,N_1888,N_2264);
or U2932 (N_2932,N_2358,N_2344);
and U2933 (N_2933,N_2349,N_2273);
or U2934 (N_2934,N_2278,N_1835);
nand U2935 (N_2935,N_2341,N_2129);
nor U2936 (N_2936,N_2070,N_1845);
nor U2937 (N_2937,N_1893,N_2326);
and U2938 (N_2938,N_1807,N_2079);
nor U2939 (N_2939,N_2100,N_2163);
and U2940 (N_2940,N_1862,N_1837);
nand U2941 (N_2941,N_2365,N_2216);
nor U2942 (N_2942,N_2093,N_2015);
xor U2943 (N_2943,N_2216,N_1985);
nor U2944 (N_2944,N_2123,N_2366);
nand U2945 (N_2945,N_2397,N_2037);
or U2946 (N_2946,N_2159,N_2085);
xnor U2947 (N_2947,N_2116,N_1954);
nand U2948 (N_2948,N_1965,N_2031);
and U2949 (N_2949,N_1884,N_1979);
xnor U2950 (N_2950,N_1800,N_2353);
and U2951 (N_2951,N_1919,N_2388);
and U2952 (N_2952,N_2092,N_1998);
or U2953 (N_2953,N_1941,N_2007);
and U2954 (N_2954,N_2356,N_2178);
xnor U2955 (N_2955,N_2070,N_2245);
nor U2956 (N_2956,N_1866,N_1854);
nor U2957 (N_2957,N_2267,N_2326);
nor U2958 (N_2958,N_2008,N_1867);
or U2959 (N_2959,N_1802,N_2232);
and U2960 (N_2960,N_1957,N_2209);
nor U2961 (N_2961,N_2124,N_2362);
nor U2962 (N_2962,N_1873,N_1935);
xor U2963 (N_2963,N_2138,N_1810);
and U2964 (N_2964,N_1939,N_2039);
xor U2965 (N_2965,N_2291,N_1926);
nand U2966 (N_2966,N_1952,N_1888);
xnor U2967 (N_2967,N_1964,N_1810);
nor U2968 (N_2968,N_2062,N_2127);
or U2969 (N_2969,N_1997,N_2189);
xnor U2970 (N_2970,N_1936,N_1970);
nand U2971 (N_2971,N_2294,N_1979);
and U2972 (N_2972,N_1889,N_2202);
xnor U2973 (N_2973,N_2219,N_2114);
nor U2974 (N_2974,N_1870,N_2214);
and U2975 (N_2975,N_2392,N_1801);
or U2976 (N_2976,N_2112,N_2055);
nand U2977 (N_2977,N_1803,N_2310);
xnor U2978 (N_2978,N_2301,N_2121);
and U2979 (N_2979,N_2148,N_2114);
and U2980 (N_2980,N_2127,N_2395);
nor U2981 (N_2981,N_1810,N_1972);
or U2982 (N_2982,N_2273,N_2267);
nand U2983 (N_2983,N_2034,N_2156);
or U2984 (N_2984,N_1935,N_2198);
nor U2985 (N_2985,N_1929,N_2337);
xnor U2986 (N_2986,N_2057,N_2237);
nor U2987 (N_2987,N_2037,N_2149);
or U2988 (N_2988,N_2150,N_1989);
xor U2989 (N_2989,N_1957,N_2039);
and U2990 (N_2990,N_1971,N_1866);
nand U2991 (N_2991,N_2243,N_2269);
xnor U2992 (N_2992,N_1919,N_2030);
and U2993 (N_2993,N_2021,N_2345);
or U2994 (N_2994,N_2116,N_2113);
or U2995 (N_2995,N_1835,N_1958);
or U2996 (N_2996,N_2193,N_2081);
xor U2997 (N_2997,N_2223,N_2361);
nand U2998 (N_2998,N_2136,N_2063);
or U2999 (N_2999,N_2132,N_1800);
or UO_0 (O_0,N_2817,N_2868);
nand UO_1 (O_1,N_2540,N_2653);
or UO_2 (O_2,N_2624,N_2793);
nor UO_3 (O_3,N_2758,N_2963);
nor UO_4 (O_4,N_2880,N_2443);
and UO_5 (O_5,N_2630,N_2730);
nand UO_6 (O_6,N_2469,N_2587);
or UO_7 (O_7,N_2706,N_2826);
and UO_8 (O_8,N_2908,N_2850);
xor UO_9 (O_9,N_2935,N_2507);
and UO_10 (O_10,N_2831,N_2494);
nor UO_11 (O_11,N_2522,N_2895);
nor UO_12 (O_12,N_2805,N_2909);
nand UO_13 (O_13,N_2661,N_2537);
xor UO_14 (O_14,N_2486,N_2433);
or UO_15 (O_15,N_2421,N_2997);
and UO_16 (O_16,N_2533,N_2775);
or UO_17 (O_17,N_2778,N_2479);
nand UO_18 (O_18,N_2442,N_2874);
and UO_19 (O_19,N_2626,N_2768);
nand UO_20 (O_20,N_2663,N_2838);
or UO_21 (O_21,N_2921,N_2840);
xnor UO_22 (O_22,N_2965,N_2957);
xor UO_23 (O_23,N_2687,N_2500);
nor UO_24 (O_24,N_2643,N_2407);
and UO_25 (O_25,N_2847,N_2893);
xor UO_26 (O_26,N_2857,N_2526);
or UO_27 (O_27,N_2815,N_2670);
nor UO_28 (O_28,N_2401,N_2604);
or UO_29 (O_29,N_2445,N_2923);
xor UO_30 (O_30,N_2767,N_2532);
xnor UO_31 (O_31,N_2959,N_2889);
and UO_32 (O_32,N_2419,N_2867);
nor UO_33 (O_33,N_2927,N_2415);
or UO_34 (O_34,N_2460,N_2422);
nor UO_35 (O_35,N_2844,N_2948);
xnor UO_36 (O_36,N_2735,N_2766);
and UO_37 (O_37,N_2552,N_2404);
nand UO_38 (O_38,N_2698,N_2635);
and UO_39 (O_39,N_2848,N_2430);
nor UO_40 (O_40,N_2697,N_2859);
nand UO_41 (O_41,N_2747,N_2456);
nand UO_42 (O_42,N_2651,N_2993);
xnor UO_43 (O_43,N_2922,N_2406);
or UO_44 (O_44,N_2524,N_2646);
nand UO_45 (O_45,N_2905,N_2994);
or UO_46 (O_46,N_2400,N_2739);
nand UO_47 (O_47,N_2614,N_2517);
and UO_48 (O_48,N_2928,N_2438);
nand UO_49 (O_49,N_2956,N_2878);
nor UO_50 (O_50,N_2610,N_2551);
nand UO_51 (O_51,N_2518,N_2571);
nor UO_52 (O_52,N_2839,N_2416);
nand UO_53 (O_53,N_2477,N_2535);
and UO_54 (O_54,N_2936,N_2951);
or UO_55 (O_55,N_2509,N_2764);
and UO_56 (O_56,N_2884,N_2435);
or UO_57 (O_57,N_2876,N_2666);
nand UO_58 (O_58,N_2668,N_2870);
and UO_59 (O_59,N_2591,N_2757);
and UO_60 (O_60,N_2882,N_2966);
nor UO_61 (O_61,N_2784,N_2737);
xor UO_62 (O_62,N_2420,N_2836);
nor UO_63 (O_63,N_2937,N_2811);
xnor UO_64 (O_64,N_2631,N_2871);
xor UO_65 (O_65,N_2919,N_2934);
or UO_66 (O_66,N_2545,N_2402);
and UO_67 (O_67,N_2744,N_2515);
or UO_68 (O_68,N_2695,N_2762);
and UO_69 (O_69,N_2642,N_2930);
nor UO_70 (O_70,N_2891,N_2875);
and UO_71 (O_71,N_2453,N_2502);
and UO_72 (O_72,N_2572,N_2405);
nand UO_73 (O_73,N_2558,N_2904);
nand UO_74 (O_74,N_2869,N_2851);
xor UO_75 (O_75,N_2669,N_2593);
or UO_76 (O_76,N_2557,N_2929);
nand UO_77 (O_77,N_2563,N_2579);
nor UO_78 (O_78,N_2411,N_2506);
or UO_79 (O_79,N_2588,N_2647);
or UO_80 (O_80,N_2656,N_2898);
nand UO_81 (O_81,N_2603,N_2931);
nor UO_82 (O_82,N_2724,N_2525);
nor UO_83 (O_83,N_2822,N_2933);
xnor UO_84 (O_84,N_2426,N_2632);
or UO_85 (O_85,N_2861,N_2717);
and UO_86 (O_86,N_2681,N_2789);
or UO_87 (O_87,N_2577,N_2621);
nor UO_88 (O_88,N_2711,N_2719);
and UO_89 (O_89,N_2746,N_2846);
nor UO_90 (O_90,N_2423,N_2903);
nor UO_91 (O_91,N_2629,N_2710);
xnor UO_92 (O_92,N_2704,N_2489);
or UO_93 (O_93,N_2733,N_2449);
or UO_94 (O_94,N_2684,N_2498);
nor UO_95 (O_95,N_2776,N_2829);
or UO_96 (O_96,N_2598,N_2541);
nand UO_97 (O_97,N_2821,N_2873);
nand UO_98 (O_98,N_2660,N_2452);
xor UO_99 (O_99,N_2978,N_2677);
xor UO_100 (O_100,N_2641,N_2977);
nor UO_101 (O_101,N_2655,N_2550);
xnor UO_102 (O_102,N_2788,N_2812);
or UO_103 (O_103,N_2576,N_2800);
xor UO_104 (O_104,N_2440,N_2796);
nor UO_105 (O_105,N_2731,N_2490);
nand UO_106 (O_106,N_2939,N_2454);
nor UO_107 (O_107,N_2819,N_2879);
nor UO_108 (O_108,N_2544,N_2781);
and UO_109 (O_109,N_2485,N_2947);
xnor UO_110 (O_110,N_2856,N_2925);
xnor UO_111 (O_111,N_2801,N_2476);
nand UO_112 (O_112,N_2536,N_2917);
xor UO_113 (O_113,N_2592,N_2464);
xnor UO_114 (O_114,N_2804,N_2451);
and UO_115 (O_115,N_2990,N_2495);
nand UO_116 (O_116,N_2664,N_2832);
and UO_117 (O_117,N_2803,N_2619);
or UO_118 (O_118,N_2914,N_2508);
and UO_119 (O_119,N_2749,N_2470);
or UO_120 (O_120,N_2809,N_2699);
or UO_121 (O_121,N_2648,N_2566);
or UO_122 (O_122,N_2862,N_2763);
or UO_123 (O_123,N_2940,N_2946);
nor UO_124 (O_124,N_2599,N_2465);
xor UO_125 (O_125,N_2662,N_2645);
xnor UO_126 (O_126,N_2410,N_2570);
nor UO_127 (O_127,N_2618,N_2751);
nor UO_128 (O_128,N_2478,N_2975);
and UO_129 (O_129,N_2998,N_2896);
or UO_130 (O_130,N_2752,N_2813);
nand UO_131 (O_131,N_2807,N_2802);
and UO_132 (O_132,N_2753,N_2561);
xor UO_133 (O_133,N_2491,N_2770);
xor UO_134 (O_134,N_2617,N_2949);
nand UO_135 (O_135,N_2968,N_2623);
xor UO_136 (O_136,N_2596,N_2825);
xor UO_137 (O_137,N_2657,N_2759);
and UO_138 (O_138,N_2855,N_2823);
nor UO_139 (O_139,N_2732,N_2611);
xor UO_140 (O_140,N_2530,N_2534);
or UO_141 (O_141,N_2582,N_2787);
and UO_142 (O_142,N_2511,N_2713);
nor UO_143 (O_143,N_2890,N_2496);
or UO_144 (O_144,N_2864,N_2429);
nor UO_145 (O_145,N_2595,N_2488);
or UO_146 (O_146,N_2771,N_2484);
nor UO_147 (O_147,N_2542,N_2709);
nand UO_148 (O_148,N_2455,N_2471);
nand UO_149 (O_149,N_2911,N_2436);
nor UO_150 (O_150,N_2858,N_2521);
nand UO_151 (O_151,N_2792,N_2602);
nand UO_152 (O_152,N_2584,N_2637);
nor UO_153 (O_153,N_2459,N_2625);
nor UO_154 (O_154,N_2980,N_2761);
nor UO_155 (O_155,N_2519,N_2721);
xnor UO_156 (O_156,N_2413,N_2633);
nor UO_157 (O_157,N_2955,N_2818);
and UO_158 (O_158,N_2988,N_2981);
and UO_159 (O_159,N_2466,N_2497);
or UO_160 (O_160,N_2707,N_2575);
nor UO_161 (O_161,N_2481,N_2608);
nor UO_162 (O_162,N_2690,N_2634);
and UO_163 (O_163,N_2720,N_2573);
nor UO_164 (O_164,N_2529,N_2915);
and UO_165 (O_165,N_2835,N_2510);
nor UO_166 (O_166,N_2984,N_2808);
nand UO_167 (O_167,N_2750,N_2703);
and UO_168 (O_168,N_2692,N_2913);
or UO_169 (O_169,N_2590,N_2565);
xnor UO_170 (O_170,N_2547,N_2597);
nand UO_171 (O_171,N_2600,N_2854);
nand UO_172 (O_172,N_2897,N_2887);
xor UO_173 (O_173,N_2673,N_2727);
and UO_174 (O_174,N_2417,N_2463);
nand UO_175 (O_175,N_2457,N_2468);
xnor UO_176 (O_176,N_2999,N_2798);
nand UO_177 (O_177,N_2493,N_2782);
and UO_178 (O_178,N_2601,N_2568);
or UO_179 (O_179,N_2652,N_2425);
nor UO_180 (O_180,N_2740,N_2567);
or UO_181 (O_181,N_2546,N_2691);
nor UO_182 (O_182,N_2672,N_2837);
nand UO_183 (O_183,N_2888,N_2627);
xor UO_184 (O_184,N_2961,N_2986);
nor UO_185 (O_185,N_2820,N_2441);
nor UO_186 (O_186,N_2701,N_2754);
nor UO_187 (O_187,N_2501,N_2786);
and UO_188 (O_188,N_2556,N_2841);
nor UO_189 (O_189,N_2555,N_2444);
nand UO_190 (O_190,N_2885,N_2971);
or UO_191 (O_191,N_2434,N_2683);
xnor UO_192 (O_192,N_2799,N_2943);
or UO_193 (O_193,N_2830,N_2659);
nor UO_194 (O_194,N_2866,N_2976);
or UO_195 (O_195,N_2685,N_2979);
xnor UO_196 (O_196,N_2605,N_2554);
and UO_197 (O_197,N_2680,N_2738);
xor UO_198 (O_198,N_2810,N_2458);
nor UO_199 (O_199,N_2883,N_2446);
xnor UO_200 (O_200,N_2970,N_2613);
nand UO_201 (O_201,N_2972,N_2718);
and UO_202 (O_202,N_2578,N_2755);
and UO_203 (O_203,N_2628,N_2480);
and UO_204 (O_204,N_2562,N_2772);
xor UO_205 (O_205,N_2676,N_2606);
nand UO_206 (O_206,N_2688,N_2726);
and UO_207 (O_207,N_2926,N_2992);
and UO_208 (O_208,N_2828,N_2513);
nand UO_209 (O_209,N_2872,N_2954);
or UO_210 (O_210,N_2722,N_2475);
xnor UO_211 (O_211,N_2408,N_2686);
or UO_212 (O_212,N_2589,N_2708);
xnor UO_213 (O_213,N_2523,N_2725);
and UO_214 (O_214,N_2900,N_2845);
nor UO_215 (O_215,N_2682,N_2962);
nand UO_216 (O_216,N_2785,N_2765);
nand UO_217 (O_217,N_2678,N_2548);
nor UO_218 (O_218,N_2414,N_2969);
or UO_219 (O_219,N_2615,N_2638);
and UO_220 (O_220,N_2539,N_2428);
or UO_221 (O_221,N_2418,N_2991);
nor UO_222 (O_222,N_2806,N_2472);
xnor UO_223 (O_223,N_2607,N_2942);
xnor UO_224 (O_224,N_2985,N_2640);
nor UO_225 (O_225,N_2989,N_2403);
nor UO_226 (O_226,N_2512,N_2729);
xor UO_227 (O_227,N_2748,N_2996);
or UO_228 (O_228,N_2920,N_2894);
or UO_229 (O_229,N_2877,N_2487);
nor UO_230 (O_230,N_2499,N_2409);
nand UO_231 (O_231,N_2667,N_2938);
and UO_232 (O_232,N_2474,N_2745);
or UO_233 (O_233,N_2842,N_2531);
nand UO_234 (O_234,N_2983,N_2492);
and UO_235 (O_235,N_2960,N_2723);
and UO_236 (O_236,N_2482,N_2843);
nand UO_237 (O_237,N_2527,N_2712);
nand UO_238 (O_238,N_2743,N_2549);
and UO_239 (O_239,N_2675,N_2714);
and UO_240 (O_240,N_2514,N_2461);
or UO_241 (O_241,N_2953,N_2932);
nor UO_242 (O_242,N_2794,N_2580);
nand UO_243 (O_243,N_2447,N_2901);
and UO_244 (O_244,N_2504,N_2916);
and UO_245 (O_245,N_2437,N_2860);
xor UO_246 (O_246,N_2791,N_2696);
xor UO_247 (O_247,N_2483,N_2431);
nand UO_248 (O_248,N_2756,N_2674);
or UO_249 (O_249,N_2814,N_2964);
or UO_250 (O_250,N_2622,N_2503);
or UO_251 (O_251,N_2967,N_2612);
and UO_252 (O_252,N_2987,N_2543);
and UO_253 (O_253,N_2944,N_2728);
nand UO_254 (O_254,N_2973,N_2952);
xor UO_255 (O_255,N_2780,N_2777);
xnor UO_256 (O_256,N_2769,N_2790);
nand UO_257 (O_257,N_2693,N_2941);
nor UO_258 (O_258,N_2824,N_2918);
xnor UO_259 (O_259,N_2553,N_2650);
xnor UO_260 (O_260,N_2564,N_2899);
or UO_261 (O_261,N_2594,N_2609);
or UO_262 (O_262,N_2865,N_2907);
nand UO_263 (O_263,N_2715,N_2424);
or UO_264 (O_264,N_2795,N_2639);
nor UO_265 (O_265,N_2924,N_2982);
nand UO_266 (O_266,N_2702,N_2671);
nand UO_267 (O_267,N_2902,N_2679);
and UO_268 (O_268,N_2774,N_2620);
xor UO_269 (O_269,N_2516,N_2520);
xnor UO_270 (O_270,N_2574,N_2797);
nor UO_271 (O_271,N_2760,N_2559);
nor UO_272 (O_272,N_2560,N_2462);
xor UO_273 (O_273,N_2432,N_2742);
nand UO_274 (O_274,N_2773,N_2412);
or UO_275 (O_275,N_2649,N_2505);
nand UO_276 (O_276,N_2528,N_2834);
or UO_277 (O_277,N_2616,N_2849);
nand UO_278 (O_278,N_2636,N_2950);
nor UO_279 (O_279,N_2910,N_2586);
or UO_280 (O_280,N_2833,N_2827);
xnor UO_281 (O_281,N_2427,N_2658);
or UO_282 (O_282,N_2450,N_2912);
or UO_283 (O_283,N_2448,N_2853);
xor UO_284 (O_284,N_2886,N_2705);
nor UO_285 (O_285,N_2700,N_2467);
nand UO_286 (O_286,N_2892,N_2665);
or UO_287 (O_287,N_2783,N_2569);
and UO_288 (O_288,N_2654,N_2439);
nand UO_289 (O_289,N_2995,N_2816);
xnor UO_290 (O_290,N_2585,N_2538);
xnor UO_291 (O_291,N_2734,N_2945);
and UO_292 (O_292,N_2779,N_2881);
xor UO_293 (O_293,N_2694,N_2581);
or UO_294 (O_294,N_2741,N_2958);
and UO_295 (O_295,N_2863,N_2716);
nor UO_296 (O_296,N_2583,N_2689);
nor UO_297 (O_297,N_2644,N_2852);
nand UO_298 (O_298,N_2974,N_2473);
nand UO_299 (O_299,N_2906,N_2736);
and UO_300 (O_300,N_2635,N_2823);
and UO_301 (O_301,N_2403,N_2425);
xnor UO_302 (O_302,N_2889,N_2720);
or UO_303 (O_303,N_2904,N_2813);
xnor UO_304 (O_304,N_2901,N_2943);
xor UO_305 (O_305,N_2718,N_2925);
xor UO_306 (O_306,N_2741,N_2480);
xor UO_307 (O_307,N_2527,N_2930);
or UO_308 (O_308,N_2896,N_2553);
nand UO_309 (O_309,N_2676,N_2483);
nand UO_310 (O_310,N_2417,N_2565);
xnor UO_311 (O_311,N_2663,N_2719);
xor UO_312 (O_312,N_2705,N_2931);
and UO_313 (O_313,N_2536,N_2807);
nor UO_314 (O_314,N_2409,N_2674);
xor UO_315 (O_315,N_2881,N_2809);
nand UO_316 (O_316,N_2537,N_2816);
xor UO_317 (O_317,N_2579,N_2647);
or UO_318 (O_318,N_2477,N_2835);
or UO_319 (O_319,N_2467,N_2547);
nand UO_320 (O_320,N_2410,N_2660);
or UO_321 (O_321,N_2936,N_2592);
or UO_322 (O_322,N_2629,N_2891);
or UO_323 (O_323,N_2875,N_2826);
and UO_324 (O_324,N_2986,N_2937);
nand UO_325 (O_325,N_2858,N_2940);
and UO_326 (O_326,N_2838,N_2672);
xor UO_327 (O_327,N_2799,N_2928);
nand UO_328 (O_328,N_2538,N_2579);
nand UO_329 (O_329,N_2814,N_2590);
nor UO_330 (O_330,N_2886,N_2550);
or UO_331 (O_331,N_2510,N_2545);
nor UO_332 (O_332,N_2718,N_2947);
xor UO_333 (O_333,N_2846,N_2554);
nand UO_334 (O_334,N_2848,N_2516);
xor UO_335 (O_335,N_2779,N_2735);
nor UO_336 (O_336,N_2936,N_2412);
or UO_337 (O_337,N_2667,N_2699);
nand UO_338 (O_338,N_2491,N_2409);
or UO_339 (O_339,N_2441,N_2725);
xor UO_340 (O_340,N_2465,N_2986);
and UO_341 (O_341,N_2941,N_2701);
xor UO_342 (O_342,N_2905,N_2631);
nor UO_343 (O_343,N_2543,N_2671);
or UO_344 (O_344,N_2658,N_2459);
or UO_345 (O_345,N_2935,N_2527);
or UO_346 (O_346,N_2943,N_2618);
nor UO_347 (O_347,N_2673,N_2774);
xor UO_348 (O_348,N_2700,N_2531);
nand UO_349 (O_349,N_2968,N_2589);
and UO_350 (O_350,N_2710,N_2549);
nand UO_351 (O_351,N_2537,N_2439);
and UO_352 (O_352,N_2795,N_2752);
or UO_353 (O_353,N_2713,N_2418);
xor UO_354 (O_354,N_2740,N_2858);
xnor UO_355 (O_355,N_2416,N_2410);
nand UO_356 (O_356,N_2722,N_2844);
or UO_357 (O_357,N_2738,N_2496);
and UO_358 (O_358,N_2536,N_2707);
and UO_359 (O_359,N_2794,N_2564);
nand UO_360 (O_360,N_2580,N_2593);
and UO_361 (O_361,N_2595,N_2965);
and UO_362 (O_362,N_2712,N_2759);
and UO_363 (O_363,N_2623,N_2574);
nand UO_364 (O_364,N_2701,N_2699);
nand UO_365 (O_365,N_2461,N_2830);
and UO_366 (O_366,N_2846,N_2655);
xor UO_367 (O_367,N_2499,N_2415);
nand UO_368 (O_368,N_2867,N_2982);
or UO_369 (O_369,N_2670,N_2434);
or UO_370 (O_370,N_2991,N_2921);
nand UO_371 (O_371,N_2801,N_2605);
xor UO_372 (O_372,N_2589,N_2421);
and UO_373 (O_373,N_2856,N_2824);
xnor UO_374 (O_374,N_2554,N_2581);
or UO_375 (O_375,N_2510,N_2929);
and UO_376 (O_376,N_2655,N_2456);
or UO_377 (O_377,N_2896,N_2621);
xnor UO_378 (O_378,N_2774,N_2709);
or UO_379 (O_379,N_2794,N_2834);
nor UO_380 (O_380,N_2676,N_2708);
or UO_381 (O_381,N_2957,N_2644);
xnor UO_382 (O_382,N_2602,N_2606);
xnor UO_383 (O_383,N_2709,N_2579);
nor UO_384 (O_384,N_2864,N_2936);
and UO_385 (O_385,N_2765,N_2710);
or UO_386 (O_386,N_2789,N_2942);
nand UO_387 (O_387,N_2790,N_2747);
nor UO_388 (O_388,N_2749,N_2452);
nor UO_389 (O_389,N_2948,N_2686);
nor UO_390 (O_390,N_2763,N_2592);
nor UO_391 (O_391,N_2630,N_2512);
nor UO_392 (O_392,N_2851,N_2866);
or UO_393 (O_393,N_2855,N_2726);
and UO_394 (O_394,N_2553,N_2957);
xor UO_395 (O_395,N_2805,N_2801);
and UO_396 (O_396,N_2847,N_2873);
nor UO_397 (O_397,N_2999,N_2695);
and UO_398 (O_398,N_2844,N_2976);
nor UO_399 (O_399,N_2577,N_2861);
or UO_400 (O_400,N_2902,N_2453);
and UO_401 (O_401,N_2482,N_2651);
nor UO_402 (O_402,N_2624,N_2432);
nor UO_403 (O_403,N_2584,N_2804);
xor UO_404 (O_404,N_2874,N_2949);
or UO_405 (O_405,N_2691,N_2485);
nor UO_406 (O_406,N_2799,N_2481);
nand UO_407 (O_407,N_2428,N_2660);
or UO_408 (O_408,N_2853,N_2543);
nor UO_409 (O_409,N_2562,N_2971);
or UO_410 (O_410,N_2422,N_2929);
xnor UO_411 (O_411,N_2540,N_2645);
nor UO_412 (O_412,N_2440,N_2687);
xnor UO_413 (O_413,N_2407,N_2848);
nor UO_414 (O_414,N_2484,N_2952);
and UO_415 (O_415,N_2422,N_2853);
and UO_416 (O_416,N_2969,N_2916);
nor UO_417 (O_417,N_2505,N_2450);
nor UO_418 (O_418,N_2913,N_2503);
xor UO_419 (O_419,N_2915,N_2842);
and UO_420 (O_420,N_2682,N_2627);
xnor UO_421 (O_421,N_2781,N_2512);
xor UO_422 (O_422,N_2945,N_2465);
nand UO_423 (O_423,N_2968,N_2657);
or UO_424 (O_424,N_2793,N_2417);
and UO_425 (O_425,N_2572,N_2573);
or UO_426 (O_426,N_2512,N_2904);
nor UO_427 (O_427,N_2883,N_2602);
nand UO_428 (O_428,N_2853,N_2937);
and UO_429 (O_429,N_2669,N_2615);
xor UO_430 (O_430,N_2511,N_2711);
nand UO_431 (O_431,N_2574,N_2695);
nor UO_432 (O_432,N_2720,N_2437);
nor UO_433 (O_433,N_2705,N_2436);
or UO_434 (O_434,N_2538,N_2464);
nand UO_435 (O_435,N_2749,N_2809);
and UO_436 (O_436,N_2545,N_2601);
nor UO_437 (O_437,N_2717,N_2912);
nand UO_438 (O_438,N_2544,N_2799);
or UO_439 (O_439,N_2998,N_2885);
and UO_440 (O_440,N_2425,N_2969);
or UO_441 (O_441,N_2783,N_2950);
and UO_442 (O_442,N_2563,N_2779);
nor UO_443 (O_443,N_2950,N_2588);
and UO_444 (O_444,N_2643,N_2472);
and UO_445 (O_445,N_2403,N_2984);
nor UO_446 (O_446,N_2732,N_2527);
nor UO_447 (O_447,N_2949,N_2868);
xnor UO_448 (O_448,N_2721,N_2404);
or UO_449 (O_449,N_2403,N_2630);
or UO_450 (O_450,N_2915,N_2764);
or UO_451 (O_451,N_2576,N_2403);
nand UO_452 (O_452,N_2912,N_2485);
or UO_453 (O_453,N_2869,N_2401);
nand UO_454 (O_454,N_2927,N_2631);
nand UO_455 (O_455,N_2711,N_2505);
nand UO_456 (O_456,N_2797,N_2607);
nand UO_457 (O_457,N_2823,N_2707);
xnor UO_458 (O_458,N_2702,N_2909);
and UO_459 (O_459,N_2605,N_2494);
nand UO_460 (O_460,N_2921,N_2963);
or UO_461 (O_461,N_2867,N_2927);
or UO_462 (O_462,N_2667,N_2533);
and UO_463 (O_463,N_2626,N_2707);
xnor UO_464 (O_464,N_2860,N_2481);
xor UO_465 (O_465,N_2999,N_2641);
nor UO_466 (O_466,N_2697,N_2443);
nor UO_467 (O_467,N_2902,N_2408);
and UO_468 (O_468,N_2657,N_2734);
xor UO_469 (O_469,N_2886,N_2612);
xnor UO_470 (O_470,N_2871,N_2734);
nand UO_471 (O_471,N_2874,N_2483);
or UO_472 (O_472,N_2947,N_2899);
nor UO_473 (O_473,N_2636,N_2628);
xor UO_474 (O_474,N_2870,N_2688);
and UO_475 (O_475,N_2470,N_2815);
or UO_476 (O_476,N_2714,N_2557);
or UO_477 (O_477,N_2542,N_2907);
nand UO_478 (O_478,N_2755,N_2787);
and UO_479 (O_479,N_2907,N_2956);
nor UO_480 (O_480,N_2993,N_2839);
nor UO_481 (O_481,N_2626,N_2655);
nand UO_482 (O_482,N_2992,N_2704);
and UO_483 (O_483,N_2723,N_2979);
or UO_484 (O_484,N_2415,N_2642);
nand UO_485 (O_485,N_2406,N_2636);
and UO_486 (O_486,N_2861,N_2875);
nand UO_487 (O_487,N_2957,N_2855);
xor UO_488 (O_488,N_2556,N_2699);
and UO_489 (O_489,N_2601,N_2889);
nor UO_490 (O_490,N_2753,N_2507);
or UO_491 (O_491,N_2561,N_2794);
and UO_492 (O_492,N_2813,N_2564);
or UO_493 (O_493,N_2469,N_2892);
or UO_494 (O_494,N_2606,N_2917);
nor UO_495 (O_495,N_2972,N_2856);
nor UO_496 (O_496,N_2886,N_2478);
or UO_497 (O_497,N_2522,N_2996);
and UO_498 (O_498,N_2742,N_2773);
nor UO_499 (O_499,N_2494,N_2953);
endmodule