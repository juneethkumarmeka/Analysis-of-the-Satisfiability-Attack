module basic_1000_10000_1500_4_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_174,In_977);
nand U1 (N_1,In_380,In_95);
or U2 (N_2,In_610,In_713);
nor U3 (N_3,In_776,In_406);
and U4 (N_4,In_354,In_491);
nand U5 (N_5,In_457,In_134);
nand U6 (N_6,In_205,In_54);
nand U7 (N_7,In_312,In_161);
or U8 (N_8,In_908,In_316);
or U9 (N_9,In_510,In_912);
nor U10 (N_10,In_709,In_347);
xor U11 (N_11,In_999,In_627);
nor U12 (N_12,In_72,In_771);
and U13 (N_13,In_2,In_973);
and U14 (N_14,In_869,In_433);
or U15 (N_15,In_261,In_129);
or U16 (N_16,In_145,In_343);
nand U17 (N_17,In_669,In_690);
and U18 (N_18,In_310,In_583);
or U19 (N_19,In_43,In_360);
nand U20 (N_20,In_692,In_516);
or U21 (N_21,In_863,In_611);
nor U22 (N_22,In_110,In_270);
or U23 (N_23,In_202,In_720);
or U24 (N_24,In_582,In_472);
and U25 (N_25,In_846,In_671);
nor U26 (N_26,In_1,In_336);
and U27 (N_27,In_702,In_634);
nor U28 (N_28,In_127,In_988);
nand U29 (N_29,In_641,In_169);
nor U30 (N_30,In_166,In_984);
nor U31 (N_31,In_682,In_961);
nand U32 (N_32,In_666,In_707);
and U33 (N_33,In_477,In_640);
nand U34 (N_34,In_564,In_440);
nor U35 (N_35,In_920,In_880);
and U36 (N_36,In_629,In_475);
or U37 (N_37,In_294,In_957);
and U38 (N_38,In_88,In_409);
xnor U39 (N_39,In_591,In_455);
nand U40 (N_40,In_703,In_235);
xnor U41 (N_41,In_27,In_58);
or U42 (N_42,In_162,In_264);
nor U43 (N_43,In_228,In_509);
nand U44 (N_44,In_974,In_394);
and U45 (N_45,In_520,In_885);
and U46 (N_46,In_293,In_534);
nor U47 (N_47,In_266,In_584);
or U48 (N_48,In_302,In_291);
nand U49 (N_49,In_375,In_946);
nand U50 (N_50,In_956,In_327);
or U51 (N_51,In_792,In_78);
and U52 (N_52,In_827,In_315);
xor U53 (N_53,In_92,In_6);
nand U54 (N_54,In_898,In_934);
or U55 (N_55,In_185,In_960);
nor U56 (N_56,In_943,In_239);
nor U57 (N_57,In_987,In_19);
or U58 (N_58,In_779,In_60);
or U59 (N_59,In_431,In_546);
nor U60 (N_60,In_416,In_49);
or U61 (N_61,In_501,In_816);
or U62 (N_62,In_408,In_888);
or U63 (N_63,In_979,In_989);
or U64 (N_64,In_899,In_916);
and U65 (N_65,In_405,In_972);
or U66 (N_66,In_372,In_502);
nand U67 (N_67,In_278,In_780);
or U68 (N_68,In_111,In_545);
nand U69 (N_69,In_11,In_396);
or U70 (N_70,In_348,In_981);
or U71 (N_71,In_335,In_337);
nor U72 (N_72,In_824,In_998);
nor U73 (N_73,In_919,In_819);
nor U74 (N_74,In_480,In_855);
nor U75 (N_75,In_462,In_643);
nor U76 (N_76,In_361,In_924);
and U77 (N_77,In_171,In_823);
nor U78 (N_78,In_388,In_263);
nor U79 (N_79,In_925,In_808);
nand U80 (N_80,In_829,In_874);
or U81 (N_81,In_445,In_559);
or U82 (N_82,In_598,In_642);
or U83 (N_83,In_673,In_203);
xor U84 (N_84,In_993,In_283);
nand U85 (N_85,In_208,In_186);
nand U86 (N_86,In_333,In_482);
or U87 (N_87,In_190,In_281);
and U88 (N_88,In_801,In_646);
nand U89 (N_89,In_104,In_747);
nor U90 (N_90,In_179,In_437);
nand U91 (N_91,In_505,In_524);
or U92 (N_92,In_726,In_872);
nand U93 (N_93,In_153,In_45);
or U94 (N_94,In_744,In_966);
xnor U95 (N_95,In_746,In_840);
nand U96 (N_96,In_672,In_907);
xnor U97 (N_97,In_470,In_909);
or U98 (N_98,In_149,In_124);
nand U99 (N_99,In_198,In_3);
and U100 (N_100,In_130,In_137);
and U101 (N_101,In_484,In_68);
nand U102 (N_102,In_851,In_459);
nor U103 (N_103,In_217,In_825);
and U104 (N_104,In_541,In_918);
nor U105 (N_105,In_249,In_188);
or U106 (N_106,In_288,In_342);
or U107 (N_107,In_414,In_248);
nor U108 (N_108,In_773,In_962);
nor U109 (N_109,In_30,In_154);
or U110 (N_110,In_511,In_426);
xor U111 (N_111,In_97,In_652);
or U112 (N_112,In_942,In_842);
nand U113 (N_113,In_800,In_573);
and U114 (N_114,In_101,In_12);
or U115 (N_115,In_826,In_533);
nand U116 (N_116,In_531,In_292);
and U117 (N_117,In_128,In_280);
nor U118 (N_118,In_114,In_600);
and U119 (N_119,In_471,In_811);
or U120 (N_120,In_170,In_9);
or U121 (N_121,In_948,In_536);
and U122 (N_122,In_799,In_172);
nor U123 (N_123,In_305,In_653);
or U124 (N_124,In_767,In_844);
nand U125 (N_125,In_499,In_522);
nand U126 (N_126,In_893,In_492);
nand U127 (N_127,In_309,In_861);
nor U128 (N_128,In_135,In_745);
or U129 (N_129,In_63,In_637);
nor U130 (N_130,In_847,In_70);
or U131 (N_131,In_102,In_173);
nor U132 (N_132,In_15,In_216);
nor U133 (N_133,In_308,In_233);
or U134 (N_134,In_705,In_715);
xor U135 (N_135,In_62,In_421);
nand U136 (N_136,In_879,In_26);
nand U137 (N_137,In_64,In_731);
nor U138 (N_138,In_512,In_857);
nor U139 (N_139,In_719,In_763);
or U140 (N_140,In_706,In_814);
nor U141 (N_141,In_123,In_366);
nand U142 (N_142,In_741,In_782);
or U143 (N_143,In_759,In_377);
nor U144 (N_144,In_300,In_914);
and U145 (N_145,In_915,In_976);
or U146 (N_146,In_526,In_341);
nor U147 (N_147,In_439,In_834);
nand U148 (N_148,In_680,In_122);
nand U149 (N_149,In_887,In_606);
and U150 (N_150,In_685,In_31);
nand U151 (N_151,In_397,In_77);
nand U152 (N_152,In_772,In_220);
xnor U153 (N_153,In_136,In_143);
or U154 (N_154,In_454,In_14);
or U155 (N_155,In_498,In_200);
or U156 (N_156,In_662,In_109);
nand U157 (N_157,In_786,In_635);
nand U158 (N_158,In_797,In_699);
and U159 (N_159,In_521,In_906);
nand U160 (N_160,In_750,In_483);
nand U161 (N_161,In_619,In_46);
nand U162 (N_162,In_419,In_314);
nor U163 (N_163,In_151,In_453);
nor U164 (N_164,In_65,In_578);
and U165 (N_165,In_441,In_785);
xnor U166 (N_166,In_631,In_784);
xor U167 (N_167,In_716,In_287);
or U168 (N_168,In_89,In_44);
and U169 (N_169,In_955,In_362);
and U170 (N_170,In_905,In_739);
and U171 (N_171,In_859,In_896);
xor U172 (N_172,In_251,In_935);
and U173 (N_173,In_399,In_450);
nand U174 (N_174,In_940,In_883);
nand U175 (N_175,In_146,In_359);
nand U176 (N_176,In_428,In_903);
nand U177 (N_177,In_489,In_992);
or U178 (N_178,In_996,In_275);
and U179 (N_179,In_886,In_13);
or U180 (N_180,In_478,In_544);
nor U181 (N_181,In_736,In_687);
and U182 (N_182,In_810,In_479);
nand U183 (N_183,In_383,In_994);
nand U184 (N_184,In_738,In_451);
or U185 (N_185,In_116,In_488);
and U186 (N_186,In_182,In_626);
nor U187 (N_187,In_193,In_950);
and U188 (N_188,In_237,In_749);
and U189 (N_189,In_322,In_507);
nor U190 (N_190,In_538,In_625);
xor U191 (N_191,In_345,In_107);
or U192 (N_192,In_225,In_947);
and U193 (N_193,In_167,In_301);
nor U194 (N_194,In_50,In_730);
and U195 (N_195,In_659,In_403);
nand U196 (N_196,In_997,In_32);
nor U197 (N_197,In_820,In_307);
and U198 (N_198,In_422,In_815);
nand U199 (N_199,In_17,In_214);
nor U200 (N_200,In_762,In_681);
nand U201 (N_201,In_504,In_781);
nand U202 (N_202,In_932,In_94);
and U203 (N_203,In_938,In_630);
xnor U204 (N_204,In_242,In_332);
and U205 (N_205,In_390,In_794);
nor U206 (N_206,In_740,In_51);
nand U207 (N_207,In_882,In_490);
nand U208 (N_208,In_215,In_722);
nand U209 (N_209,In_931,In_609);
and U210 (N_210,In_742,In_565);
or U211 (N_211,In_513,In_679);
or U212 (N_212,In_602,In_930);
nor U213 (N_213,In_425,In_777);
xnor U214 (N_214,In_61,In_100);
nand U215 (N_215,In_518,In_766);
nand U216 (N_216,In_614,In_959);
nor U217 (N_217,In_339,In_636);
or U218 (N_218,In_751,In_620);
or U219 (N_219,In_543,In_676);
or U220 (N_220,In_423,In_265);
nand U221 (N_221,In_245,In_900);
nor U222 (N_222,In_210,In_276);
nor U223 (N_223,In_554,In_805);
nand U224 (N_224,In_866,In_382);
and U225 (N_225,In_96,In_648);
nand U226 (N_226,In_668,In_570);
nand U227 (N_227,In_607,In_85);
and U228 (N_228,In_392,In_481);
or U229 (N_229,In_941,In_349);
or U230 (N_230,In_219,In_369);
or U231 (N_231,In_356,In_579);
nand U232 (N_232,In_737,In_184);
or U233 (N_233,In_73,In_537);
and U234 (N_234,In_895,In_473);
or U235 (N_235,In_204,In_628);
nand U236 (N_236,In_298,In_822);
and U237 (N_237,In_69,In_158);
nand U238 (N_238,In_809,In_655);
nand U239 (N_239,In_753,In_683);
nand U240 (N_240,In_663,In_791);
nor U241 (N_241,In_858,In_467);
nor U242 (N_242,In_556,In_862);
nand U243 (N_243,In_191,In_351);
and U244 (N_244,In_563,In_571);
nor U245 (N_245,In_304,In_120);
nor U246 (N_246,In_980,In_187);
or U247 (N_247,In_461,In_211);
or U248 (N_248,In_227,In_807);
and U249 (N_249,In_639,In_557);
or U250 (N_250,In_456,In_255);
and U251 (N_251,In_160,In_649);
or U252 (N_252,In_698,In_175);
nor U253 (N_253,In_689,In_150);
and U254 (N_254,In_868,In_141);
and U255 (N_255,In_37,In_789);
nor U256 (N_256,In_694,In_113);
nand U257 (N_257,In_10,In_657);
or U258 (N_258,In_4,In_82);
nor U259 (N_259,In_644,In_376);
nor U260 (N_260,In_894,In_953);
nand U261 (N_261,In_774,In_661);
nor U262 (N_262,In_241,In_904);
or U263 (N_263,In_432,In_121);
nand U264 (N_264,In_420,In_199);
and U265 (N_265,In_108,In_494);
or U266 (N_266,In_231,In_415);
nor U267 (N_267,In_593,In_528);
nor U268 (N_268,In_207,In_272);
xnor U269 (N_269,In_358,In_581);
and U270 (N_270,In_448,In_764);
nor U271 (N_271,In_317,In_945);
nor U272 (N_272,In_778,In_74);
or U273 (N_273,In_849,In_575);
and U274 (N_274,In_212,In_732);
nand U275 (N_275,In_465,In_770);
nor U276 (N_276,In_497,In_284);
nand U277 (N_277,In_438,In_697);
and U278 (N_278,In_970,In_458);
nand U279 (N_279,In_371,In_991);
and U280 (N_280,In_56,In_176);
nand U281 (N_281,In_20,In_608);
nand U282 (N_282,In_367,In_447);
nand U283 (N_283,In_760,In_658);
or U284 (N_284,In_22,In_90);
nor U285 (N_285,In_67,In_395);
or U286 (N_286,In_389,In_381);
and U287 (N_287,In_936,In_87);
nor U288 (N_288,In_838,In_86);
nand U289 (N_289,In_177,In_542);
or U290 (N_290,In_986,In_232);
or U291 (N_291,In_667,In_257);
nand U292 (N_292,In_147,In_319);
nor U293 (N_293,In_155,In_765);
nand U294 (N_294,In_708,In_892);
or U295 (N_295,In_240,In_891);
or U296 (N_296,In_837,In_647);
nor U297 (N_297,In_508,In_968);
and U298 (N_298,In_500,In_547);
and U299 (N_299,In_47,In_601);
or U300 (N_300,In_540,In_285);
nand U301 (N_301,In_180,In_693);
nor U302 (N_302,In_684,In_365);
or U303 (N_303,In_645,In_517);
or U304 (N_304,In_975,In_831);
xor U305 (N_305,In_875,In_24);
nand U306 (N_306,In_410,In_260);
nand U307 (N_307,In_350,In_318);
nor U308 (N_308,In_328,In_413);
nand U309 (N_309,In_818,In_181);
or U310 (N_310,In_443,In_446);
or U311 (N_311,In_969,In_576);
and U312 (N_312,In_572,In_7);
nand U313 (N_313,In_552,In_864);
nand U314 (N_314,In_402,In_412);
nor U315 (N_315,In_76,In_468);
and U316 (N_316,In_677,In_400);
nor U317 (N_317,In_612,In_853);
nor U318 (N_318,In_118,In_718);
and U319 (N_319,In_615,In_353);
and U320 (N_320,In_452,In_954);
nor U321 (N_321,In_133,In_725);
or U322 (N_322,In_340,In_560);
nor U323 (N_323,In_525,In_321);
and U324 (N_324,In_258,In_860);
nand U325 (N_325,In_664,In_18);
and U326 (N_326,In_618,In_870);
and U327 (N_327,In_995,In_144);
or U328 (N_328,In_99,In_368);
and U329 (N_329,In_599,In_93);
or U330 (N_330,In_971,In_464);
nor U331 (N_331,In_357,In_138);
and U332 (N_332,In_355,In_469);
nor U333 (N_333,In_674,In_733);
and U334 (N_334,In_616,In_878);
xor U335 (N_335,In_33,In_804);
nand U336 (N_336,In_551,In_250);
and U337 (N_337,In_192,In_913);
and U338 (N_338,In_66,In_585);
or U339 (N_339,In_460,In_890);
and U340 (N_340,In_295,In_435);
or U341 (N_341,In_474,In_271);
or U342 (N_342,In_743,In_877);
and U343 (N_343,In_821,In_463);
nor U344 (N_344,In_704,In_194);
or U345 (N_345,In_373,In_411);
nor U346 (N_346,In_603,In_434);
nand U347 (N_347,In_230,In_487);
nor U348 (N_348,In_613,In_29);
and U349 (N_349,In_35,In_41);
nor U350 (N_350,In_580,In_597);
nand U351 (N_351,In_712,In_503);
or U352 (N_352,In_568,In_183);
nand U353 (N_353,In_401,In_700);
and U354 (N_354,In_795,In_982);
nand U355 (N_355,In_754,In_277);
nor U356 (N_356,In_835,In_269);
nand U357 (N_357,In_8,In_75);
nor U358 (N_358,In_79,In_427);
nor U359 (N_359,In_555,In_752);
nand U360 (N_360,In_243,In_798);
nor U361 (N_361,In_757,In_48);
and U362 (N_362,In_370,In_28);
or U363 (N_363,In_654,In_928);
nor U364 (N_364,In_178,In_132);
and U365 (N_365,In_466,In_485);
or U366 (N_366,In_939,In_836);
nand U367 (N_367,In_313,In_802);
and U368 (N_368,In_140,In_735);
and U369 (N_369,In_921,In_444);
xnor U370 (N_370,In_247,In_106);
and U371 (N_371,In_268,In_334);
nor U372 (N_372,In_553,In_796);
xor U373 (N_373,In_841,In_91);
xnor U374 (N_374,In_539,In_244);
and U375 (N_375,In_933,In_695);
nor U376 (N_376,In_52,In_696);
nand U377 (N_377,In_624,In_429);
and U378 (N_378,In_103,In_519);
nand U379 (N_379,In_964,In_515);
and U380 (N_380,In_320,In_55);
nor U381 (N_381,In_25,In_16);
nand U382 (N_382,In_476,In_152);
nand U383 (N_383,In_978,In_574);
nand U384 (N_384,In_352,In_952);
nor U385 (N_385,In_717,In_621);
and U386 (N_386,In_633,In_398);
nor U387 (N_387,In_832,In_527);
nand U388 (N_388,In_833,In_605);
and U389 (N_389,In_549,In_843);
nand U390 (N_390,In_0,In_81);
nor U391 (N_391,In_867,In_157);
nor U392 (N_392,In_569,In_282);
nand U393 (N_393,In_206,In_329);
and U394 (N_394,In_638,In_246);
and U395 (N_395,In_670,In_691);
or U396 (N_396,In_828,In_38);
and U397 (N_397,In_363,In_562);
nand U398 (N_398,In_949,In_164);
nor U399 (N_399,In_131,In_963);
nor U400 (N_400,In_852,In_21);
or U401 (N_401,In_660,In_163);
nand U402 (N_402,In_148,In_678);
nand U403 (N_403,In_23,In_675);
xor U404 (N_404,In_378,In_876);
and U405 (N_405,In_229,In_793);
nor U406 (N_406,In_723,In_812);
xnor U407 (N_407,In_926,In_253);
nor U408 (N_408,In_755,In_632);
and U409 (N_409,In_985,In_262);
or U410 (N_410,In_297,In_53);
or U411 (N_411,In_506,In_561);
nand U412 (N_412,In_604,In_259);
nand U413 (N_413,In_937,In_839);
nor U414 (N_414,In_156,In_529);
nand U415 (N_415,In_927,In_404);
or U416 (N_416,In_126,In_850);
and U417 (N_417,In_387,In_865);
or U418 (N_418,In_418,In_566);
and U419 (N_419,In_768,In_594);
and U420 (N_420,In_486,In_727);
nand U421 (N_421,In_787,In_817);
nor U422 (N_422,In_535,In_922);
nor U423 (N_423,In_424,In_990);
nand U424 (N_424,In_495,In_386);
nor U425 (N_425,In_59,In_845);
or U426 (N_426,In_338,In_587);
nor U427 (N_427,In_273,In_236);
nand U428 (N_428,In_57,In_967);
and U429 (N_429,In_238,In_213);
nand U430 (N_430,In_721,In_222);
nor U431 (N_431,In_944,In_83);
and U432 (N_432,In_769,In_761);
nor U433 (N_433,In_165,In_112);
xor U434 (N_434,In_391,In_929);
or U435 (N_435,In_923,In_951);
nor U436 (N_436,In_196,In_848);
nor U437 (N_437,In_550,In_530);
nand U438 (N_438,In_758,In_39);
and U439 (N_439,In_756,In_622);
nand U440 (N_440,In_286,In_119);
nand U441 (N_441,In_856,In_430);
nand U442 (N_442,In_902,In_854);
and U443 (N_443,In_701,In_274);
nand U444 (N_444,In_656,In_40);
xnor U445 (N_445,In_897,In_965);
xnor U446 (N_446,In_384,In_588);
or U447 (N_447,In_299,In_650);
nand U448 (N_448,In_330,In_592);
and U449 (N_449,In_256,In_189);
and U450 (N_450,In_234,In_830);
or U451 (N_451,In_252,In_324);
nand U452 (N_452,In_224,In_617);
nor U453 (N_453,In_803,In_496);
or U454 (N_454,In_665,In_686);
or U455 (N_455,In_385,In_724);
and U456 (N_456,In_323,In_449);
and U457 (N_457,In_442,In_195);
nand U458 (N_458,In_871,In_201);
nor U459 (N_459,In_586,In_84);
nor U460 (N_460,In_748,In_296);
nand U461 (N_461,In_958,In_374);
and U462 (N_462,In_532,In_558);
nor U463 (N_463,In_596,In_36);
nor U464 (N_464,In_325,In_117);
nand U465 (N_465,In_590,In_125);
nand U466 (N_466,In_209,In_267);
or U467 (N_467,In_577,In_159);
nor U468 (N_468,In_623,In_98);
xnor U469 (N_469,In_142,In_514);
nand U470 (N_470,In_910,In_729);
and U471 (N_471,In_775,In_710);
nor U472 (N_472,In_889,In_42);
nand U473 (N_473,In_567,In_279);
nor U474 (N_474,In_589,In_417);
and U475 (N_475,In_436,In_254);
nand U476 (N_476,In_311,In_734);
nand U477 (N_477,In_688,In_5);
and U478 (N_478,In_728,In_344);
or U479 (N_479,In_218,In_651);
nand U480 (N_480,In_901,In_34);
nand U481 (N_481,In_290,In_379);
and U482 (N_482,In_917,In_393);
or U483 (N_483,In_221,In_346);
and U484 (N_484,In_788,In_80);
or U485 (N_485,In_493,In_197);
and U486 (N_486,In_331,In_873);
or U487 (N_487,In_168,In_881);
xor U488 (N_488,In_105,In_289);
nand U489 (N_489,In_884,In_226);
nor U490 (N_490,In_595,In_364);
or U491 (N_491,In_911,In_813);
or U492 (N_492,In_983,In_326);
xor U493 (N_493,In_306,In_223);
or U494 (N_494,In_139,In_711);
nand U495 (N_495,In_115,In_783);
and U496 (N_496,In_714,In_407);
and U497 (N_497,In_548,In_71);
nand U498 (N_498,In_303,In_806);
and U499 (N_499,In_790,In_523);
or U500 (N_500,In_3,In_881);
nand U501 (N_501,In_272,In_639);
nand U502 (N_502,In_261,In_977);
or U503 (N_503,In_293,In_286);
and U504 (N_504,In_670,In_186);
nand U505 (N_505,In_799,In_696);
nand U506 (N_506,In_234,In_340);
nand U507 (N_507,In_203,In_772);
or U508 (N_508,In_91,In_148);
or U509 (N_509,In_182,In_263);
and U510 (N_510,In_260,In_716);
nor U511 (N_511,In_150,In_134);
nand U512 (N_512,In_958,In_539);
and U513 (N_513,In_275,In_622);
or U514 (N_514,In_803,In_584);
and U515 (N_515,In_309,In_539);
nor U516 (N_516,In_895,In_388);
nor U517 (N_517,In_524,In_378);
nor U518 (N_518,In_997,In_237);
nor U519 (N_519,In_956,In_113);
nand U520 (N_520,In_10,In_206);
and U521 (N_521,In_897,In_75);
nand U522 (N_522,In_332,In_967);
nor U523 (N_523,In_155,In_654);
nor U524 (N_524,In_205,In_287);
nor U525 (N_525,In_364,In_654);
nand U526 (N_526,In_785,In_842);
nand U527 (N_527,In_920,In_84);
nor U528 (N_528,In_851,In_513);
or U529 (N_529,In_61,In_672);
or U530 (N_530,In_460,In_533);
nand U531 (N_531,In_146,In_408);
nand U532 (N_532,In_74,In_544);
nor U533 (N_533,In_268,In_32);
nand U534 (N_534,In_432,In_610);
nor U535 (N_535,In_144,In_13);
and U536 (N_536,In_660,In_336);
nand U537 (N_537,In_52,In_718);
nand U538 (N_538,In_58,In_659);
or U539 (N_539,In_655,In_119);
or U540 (N_540,In_291,In_848);
nand U541 (N_541,In_327,In_870);
or U542 (N_542,In_767,In_176);
nor U543 (N_543,In_675,In_462);
nand U544 (N_544,In_558,In_783);
or U545 (N_545,In_184,In_3);
nand U546 (N_546,In_977,In_251);
and U547 (N_547,In_586,In_730);
or U548 (N_548,In_155,In_374);
or U549 (N_549,In_711,In_510);
nor U550 (N_550,In_743,In_666);
nand U551 (N_551,In_17,In_475);
xor U552 (N_552,In_652,In_644);
nor U553 (N_553,In_620,In_639);
nand U554 (N_554,In_997,In_616);
and U555 (N_555,In_729,In_440);
and U556 (N_556,In_752,In_385);
nand U557 (N_557,In_330,In_566);
xor U558 (N_558,In_316,In_132);
nand U559 (N_559,In_356,In_505);
or U560 (N_560,In_18,In_773);
and U561 (N_561,In_802,In_950);
nor U562 (N_562,In_680,In_193);
nor U563 (N_563,In_97,In_131);
nand U564 (N_564,In_225,In_775);
and U565 (N_565,In_101,In_480);
nor U566 (N_566,In_645,In_680);
nor U567 (N_567,In_236,In_597);
nor U568 (N_568,In_197,In_441);
and U569 (N_569,In_373,In_876);
and U570 (N_570,In_126,In_998);
nor U571 (N_571,In_575,In_885);
or U572 (N_572,In_57,In_508);
or U573 (N_573,In_328,In_114);
nand U574 (N_574,In_289,In_490);
nand U575 (N_575,In_174,In_400);
nand U576 (N_576,In_501,In_11);
nor U577 (N_577,In_167,In_642);
and U578 (N_578,In_704,In_477);
nand U579 (N_579,In_277,In_270);
nor U580 (N_580,In_253,In_176);
nor U581 (N_581,In_362,In_212);
nand U582 (N_582,In_484,In_201);
nor U583 (N_583,In_967,In_49);
nor U584 (N_584,In_136,In_703);
nand U585 (N_585,In_921,In_434);
and U586 (N_586,In_255,In_173);
and U587 (N_587,In_411,In_58);
and U588 (N_588,In_943,In_321);
or U589 (N_589,In_767,In_797);
and U590 (N_590,In_847,In_704);
or U591 (N_591,In_274,In_797);
nor U592 (N_592,In_47,In_101);
nand U593 (N_593,In_743,In_701);
nor U594 (N_594,In_133,In_508);
nor U595 (N_595,In_497,In_274);
and U596 (N_596,In_624,In_789);
xnor U597 (N_597,In_940,In_206);
and U598 (N_598,In_291,In_474);
and U599 (N_599,In_669,In_110);
and U600 (N_600,In_186,In_594);
or U601 (N_601,In_88,In_889);
nor U602 (N_602,In_140,In_379);
nor U603 (N_603,In_182,In_115);
or U604 (N_604,In_172,In_985);
nor U605 (N_605,In_529,In_430);
or U606 (N_606,In_476,In_471);
nor U607 (N_607,In_595,In_370);
nand U608 (N_608,In_395,In_434);
nand U609 (N_609,In_67,In_838);
or U610 (N_610,In_131,In_821);
nand U611 (N_611,In_466,In_355);
or U612 (N_612,In_127,In_860);
and U613 (N_613,In_547,In_990);
nor U614 (N_614,In_256,In_523);
nand U615 (N_615,In_913,In_131);
or U616 (N_616,In_395,In_258);
nand U617 (N_617,In_619,In_183);
or U618 (N_618,In_781,In_873);
nand U619 (N_619,In_282,In_853);
nand U620 (N_620,In_279,In_716);
or U621 (N_621,In_102,In_58);
or U622 (N_622,In_371,In_50);
nor U623 (N_623,In_4,In_340);
nor U624 (N_624,In_17,In_460);
or U625 (N_625,In_858,In_195);
or U626 (N_626,In_851,In_689);
nand U627 (N_627,In_879,In_682);
and U628 (N_628,In_566,In_197);
or U629 (N_629,In_632,In_433);
nor U630 (N_630,In_14,In_307);
or U631 (N_631,In_236,In_808);
nand U632 (N_632,In_340,In_689);
or U633 (N_633,In_638,In_894);
or U634 (N_634,In_468,In_502);
or U635 (N_635,In_617,In_801);
nor U636 (N_636,In_609,In_777);
nor U637 (N_637,In_282,In_21);
xor U638 (N_638,In_676,In_77);
nand U639 (N_639,In_167,In_287);
nor U640 (N_640,In_420,In_436);
or U641 (N_641,In_977,In_86);
nand U642 (N_642,In_156,In_737);
nand U643 (N_643,In_144,In_528);
nand U644 (N_644,In_224,In_19);
or U645 (N_645,In_531,In_213);
and U646 (N_646,In_242,In_393);
nor U647 (N_647,In_310,In_605);
nor U648 (N_648,In_602,In_980);
nor U649 (N_649,In_73,In_811);
nand U650 (N_650,In_445,In_409);
nand U651 (N_651,In_604,In_14);
and U652 (N_652,In_464,In_534);
nand U653 (N_653,In_503,In_651);
nand U654 (N_654,In_398,In_760);
nand U655 (N_655,In_66,In_277);
or U656 (N_656,In_698,In_429);
or U657 (N_657,In_790,In_526);
nand U658 (N_658,In_229,In_642);
or U659 (N_659,In_777,In_384);
or U660 (N_660,In_547,In_785);
and U661 (N_661,In_983,In_912);
nor U662 (N_662,In_673,In_353);
nand U663 (N_663,In_553,In_117);
and U664 (N_664,In_862,In_525);
nor U665 (N_665,In_557,In_502);
nand U666 (N_666,In_395,In_541);
and U667 (N_667,In_694,In_823);
or U668 (N_668,In_125,In_225);
nand U669 (N_669,In_540,In_813);
or U670 (N_670,In_667,In_889);
nor U671 (N_671,In_683,In_10);
or U672 (N_672,In_844,In_566);
nor U673 (N_673,In_880,In_875);
or U674 (N_674,In_495,In_764);
nand U675 (N_675,In_127,In_70);
nand U676 (N_676,In_368,In_829);
nor U677 (N_677,In_709,In_411);
nor U678 (N_678,In_112,In_70);
or U679 (N_679,In_414,In_232);
and U680 (N_680,In_121,In_146);
nand U681 (N_681,In_127,In_597);
xnor U682 (N_682,In_856,In_834);
or U683 (N_683,In_106,In_343);
or U684 (N_684,In_83,In_951);
nor U685 (N_685,In_382,In_640);
nand U686 (N_686,In_510,In_215);
nand U687 (N_687,In_806,In_990);
nand U688 (N_688,In_104,In_667);
or U689 (N_689,In_548,In_11);
nor U690 (N_690,In_997,In_100);
or U691 (N_691,In_242,In_91);
and U692 (N_692,In_726,In_737);
or U693 (N_693,In_307,In_879);
or U694 (N_694,In_401,In_863);
and U695 (N_695,In_964,In_650);
and U696 (N_696,In_858,In_305);
and U697 (N_697,In_243,In_792);
nor U698 (N_698,In_37,In_765);
or U699 (N_699,In_242,In_404);
nand U700 (N_700,In_929,In_947);
and U701 (N_701,In_676,In_881);
or U702 (N_702,In_831,In_607);
nor U703 (N_703,In_64,In_602);
nor U704 (N_704,In_384,In_680);
nor U705 (N_705,In_422,In_472);
and U706 (N_706,In_812,In_558);
nor U707 (N_707,In_728,In_264);
nor U708 (N_708,In_791,In_254);
nand U709 (N_709,In_150,In_844);
nor U710 (N_710,In_877,In_894);
and U711 (N_711,In_361,In_561);
nor U712 (N_712,In_747,In_346);
or U713 (N_713,In_22,In_615);
nor U714 (N_714,In_727,In_179);
nand U715 (N_715,In_439,In_209);
nand U716 (N_716,In_506,In_511);
or U717 (N_717,In_149,In_172);
nor U718 (N_718,In_354,In_588);
or U719 (N_719,In_634,In_689);
and U720 (N_720,In_785,In_658);
nand U721 (N_721,In_590,In_536);
and U722 (N_722,In_107,In_620);
nand U723 (N_723,In_775,In_667);
nor U724 (N_724,In_201,In_359);
and U725 (N_725,In_695,In_409);
nor U726 (N_726,In_894,In_849);
nor U727 (N_727,In_428,In_112);
and U728 (N_728,In_291,In_632);
nor U729 (N_729,In_388,In_283);
nand U730 (N_730,In_805,In_487);
nor U731 (N_731,In_311,In_959);
nor U732 (N_732,In_93,In_463);
nand U733 (N_733,In_71,In_36);
or U734 (N_734,In_588,In_707);
and U735 (N_735,In_506,In_351);
nor U736 (N_736,In_112,In_183);
nand U737 (N_737,In_138,In_747);
or U738 (N_738,In_243,In_868);
nand U739 (N_739,In_507,In_173);
or U740 (N_740,In_462,In_361);
xor U741 (N_741,In_620,In_354);
nand U742 (N_742,In_401,In_950);
nor U743 (N_743,In_793,In_0);
nor U744 (N_744,In_53,In_795);
nor U745 (N_745,In_222,In_402);
or U746 (N_746,In_666,In_107);
and U747 (N_747,In_254,In_255);
and U748 (N_748,In_143,In_419);
and U749 (N_749,In_918,In_206);
or U750 (N_750,In_938,In_488);
and U751 (N_751,In_233,In_700);
nand U752 (N_752,In_778,In_96);
nor U753 (N_753,In_895,In_570);
nand U754 (N_754,In_782,In_647);
nor U755 (N_755,In_789,In_151);
or U756 (N_756,In_636,In_329);
or U757 (N_757,In_553,In_500);
and U758 (N_758,In_728,In_431);
nor U759 (N_759,In_918,In_621);
and U760 (N_760,In_210,In_710);
or U761 (N_761,In_438,In_516);
and U762 (N_762,In_593,In_417);
nand U763 (N_763,In_585,In_445);
or U764 (N_764,In_860,In_816);
and U765 (N_765,In_252,In_62);
nor U766 (N_766,In_627,In_123);
nor U767 (N_767,In_684,In_55);
xnor U768 (N_768,In_299,In_27);
or U769 (N_769,In_132,In_844);
nor U770 (N_770,In_494,In_486);
nand U771 (N_771,In_784,In_157);
or U772 (N_772,In_175,In_792);
xnor U773 (N_773,In_134,In_819);
or U774 (N_774,In_315,In_396);
nand U775 (N_775,In_907,In_78);
and U776 (N_776,In_8,In_852);
or U777 (N_777,In_620,In_643);
nand U778 (N_778,In_752,In_75);
nor U779 (N_779,In_229,In_226);
and U780 (N_780,In_381,In_197);
and U781 (N_781,In_434,In_537);
or U782 (N_782,In_577,In_29);
and U783 (N_783,In_930,In_53);
nand U784 (N_784,In_672,In_365);
nand U785 (N_785,In_706,In_972);
or U786 (N_786,In_276,In_391);
nand U787 (N_787,In_202,In_655);
nand U788 (N_788,In_983,In_162);
or U789 (N_789,In_431,In_349);
and U790 (N_790,In_281,In_657);
nor U791 (N_791,In_244,In_337);
nand U792 (N_792,In_270,In_922);
nand U793 (N_793,In_146,In_192);
nor U794 (N_794,In_649,In_495);
xnor U795 (N_795,In_552,In_267);
or U796 (N_796,In_392,In_459);
or U797 (N_797,In_146,In_796);
and U798 (N_798,In_925,In_964);
nor U799 (N_799,In_112,In_369);
or U800 (N_800,In_729,In_303);
nand U801 (N_801,In_20,In_482);
or U802 (N_802,In_378,In_37);
nand U803 (N_803,In_459,In_50);
xnor U804 (N_804,In_429,In_782);
and U805 (N_805,In_832,In_349);
nand U806 (N_806,In_141,In_208);
and U807 (N_807,In_678,In_961);
nor U808 (N_808,In_651,In_422);
nand U809 (N_809,In_268,In_127);
and U810 (N_810,In_879,In_246);
or U811 (N_811,In_981,In_524);
and U812 (N_812,In_900,In_43);
and U813 (N_813,In_350,In_948);
nand U814 (N_814,In_762,In_470);
nor U815 (N_815,In_394,In_391);
nand U816 (N_816,In_154,In_790);
nand U817 (N_817,In_314,In_477);
and U818 (N_818,In_226,In_553);
and U819 (N_819,In_75,In_349);
or U820 (N_820,In_332,In_881);
or U821 (N_821,In_520,In_293);
or U822 (N_822,In_358,In_344);
nor U823 (N_823,In_992,In_582);
and U824 (N_824,In_392,In_817);
nand U825 (N_825,In_484,In_364);
nand U826 (N_826,In_598,In_436);
and U827 (N_827,In_177,In_258);
nand U828 (N_828,In_619,In_204);
nand U829 (N_829,In_666,In_417);
or U830 (N_830,In_45,In_523);
and U831 (N_831,In_518,In_843);
or U832 (N_832,In_396,In_698);
nand U833 (N_833,In_12,In_256);
nor U834 (N_834,In_609,In_225);
or U835 (N_835,In_76,In_20);
and U836 (N_836,In_300,In_148);
or U837 (N_837,In_405,In_958);
nand U838 (N_838,In_550,In_479);
and U839 (N_839,In_30,In_325);
nand U840 (N_840,In_589,In_122);
nand U841 (N_841,In_790,In_267);
nand U842 (N_842,In_581,In_611);
nand U843 (N_843,In_663,In_164);
nor U844 (N_844,In_67,In_523);
and U845 (N_845,In_675,In_748);
or U846 (N_846,In_966,In_766);
or U847 (N_847,In_159,In_580);
nand U848 (N_848,In_938,In_267);
xor U849 (N_849,In_683,In_594);
nand U850 (N_850,In_205,In_511);
nand U851 (N_851,In_309,In_737);
or U852 (N_852,In_328,In_107);
nor U853 (N_853,In_618,In_366);
xor U854 (N_854,In_278,In_255);
or U855 (N_855,In_910,In_867);
and U856 (N_856,In_559,In_466);
nand U857 (N_857,In_226,In_538);
nor U858 (N_858,In_284,In_742);
and U859 (N_859,In_273,In_789);
and U860 (N_860,In_496,In_978);
or U861 (N_861,In_167,In_966);
and U862 (N_862,In_699,In_97);
nand U863 (N_863,In_894,In_594);
nand U864 (N_864,In_19,In_542);
or U865 (N_865,In_194,In_515);
nand U866 (N_866,In_854,In_86);
nor U867 (N_867,In_137,In_681);
and U868 (N_868,In_615,In_828);
nor U869 (N_869,In_2,In_198);
xnor U870 (N_870,In_183,In_970);
nand U871 (N_871,In_173,In_817);
or U872 (N_872,In_988,In_370);
and U873 (N_873,In_644,In_546);
nor U874 (N_874,In_5,In_775);
and U875 (N_875,In_322,In_212);
or U876 (N_876,In_534,In_776);
xnor U877 (N_877,In_770,In_720);
nor U878 (N_878,In_847,In_74);
nand U879 (N_879,In_956,In_682);
nand U880 (N_880,In_196,In_320);
and U881 (N_881,In_226,In_790);
nor U882 (N_882,In_37,In_968);
nand U883 (N_883,In_362,In_152);
xnor U884 (N_884,In_404,In_898);
nand U885 (N_885,In_122,In_87);
nor U886 (N_886,In_530,In_486);
and U887 (N_887,In_128,In_873);
nand U888 (N_888,In_682,In_663);
or U889 (N_889,In_534,In_456);
and U890 (N_890,In_851,In_441);
nand U891 (N_891,In_216,In_716);
nor U892 (N_892,In_50,In_11);
and U893 (N_893,In_78,In_447);
and U894 (N_894,In_628,In_556);
xor U895 (N_895,In_34,In_310);
nand U896 (N_896,In_29,In_618);
nor U897 (N_897,In_507,In_671);
and U898 (N_898,In_942,In_851);
or U899 (N_899,In_871,In_569);
and U900 (N_900,In_621,In_285);
or U901 (N_901,In_747,In_263);
and U902 (N_902,In_893,In_720);
nand U903 (N_903,In_597,In_470);
nand U904 (N_904,In_800,In_662);
or U905 (N_905,In_697,In_47);
nand U906 (N_906,In_727,In_120);
nand U907 (N_907,In_60,In_120);
or U908 (N_908,In_185,In_892);
nor U909 (N_909,In_281,In_666);
and U910 (N_910,In_52,In_392);
nand U911 (N_911,In_129,In_689);
nor U912 (N_912,In_232,In_915);
or U913 (N_913,In_911,In_670);
nand U914 (N_914,In_959,In_110);
or U915 (N_915,In_685,In_324);
and U916 (N_916,In_992,In_782);
nor U917 (N_917,In_258,In_759);
nand U918 (N_918,In_875,In_773);
xnor U919 (N_919,In_116,In_341);
nand U920 (N_920,In_443,In_494);
nand U921 (N_921,In_210,In_162);
and U922 (N_922,In_293,In_404);
or U923 (N_923,In_941,In_296);
nor U924 (N_924,In_395,In_5);
nand U925 (N_925,In_840,In_891);
nor U926 (N_926,In_998,In_343);
nor U927 (N_927,In_497,In_333);
nor U928 (N_928,In_27,In_791);
nand U929 (N_929,In_947,In_950);
or U930 (N_930,In_584,In_503);
and U931 (N_931,In_590,In_528);
nor U932 (N_932,In_818,In_487);
and U933 (N_933,In_106,In_983);
and U934 (N_934,In_379,In_61);
nand U935 (N_935,In_192,In_126);
or U936 (N_936,In_911,In_686);
or U937 (N_937,In_857,In_990);
nor U938 (N_938,In_968,In_48);
and U939 (N_939,In_15,In_515);
nand U940 (N_940,In_223,In_400);
or U941 (N_941,In_515,In_203);
and U942 (N_942,In_791,In_98);
and U943 (N_943,In_461,In_367);
or U944 (N_944,In_527,In_743);
nand U945 (N_945,In_764,In_944);
nand U946 (N_946,In_686,In_369);
or U947 (N_947,In_284,In_615);
nor U948 (N_948,In_575,In_338);
or U949 (N_949,In_995,In_719);
and U950 (N_950,In_973,In_413);
or U951 (N_951,In_354,In_656);
and U952 (N_952,In_521,In_230);
and U953 (N_953,In_193,In_184);
and U954 (N_954,In_538,In_277);
or U955 (N_955,In_808,In_585);
and U956 (N_956,In_511,In_901);
and U957 (N_957,In_917,In_354);
or U958 (N_958,In_631,In_739);
and U959 (N_959,In_570,In_989);
nor U960 (N_960,In_771,In_0);
and U961 (N_961,In_186,In_711);
nor U962 (N_962,In_193,In_281);
nand U963 (N_963,In_825,In_467);
and U964 (N_964,In_214,In_264);
and U965 (N_965,In_946,In_229);
nor U966 (N_966,In_939,In_818);
xor U967 (N_967,In_391,In_233);
and U968 (N_968,In_921,In_122);
nor U969 (N_969,In_246,In_845);
nor U970 (N_970,In_433,In_712);
nand U971 (N_971,In_93,In_780);
nand U972 (N_972,In_349,In_549);
and U973 (N_973,In_963,In_815);
nand U974 (N_974,In_78,In_304);
or U975 (N_975,In_638,In_931);
and U976 (N_976,In_668,In_512);
nor U977 (N_977,In_404,In_452);
nand U978 (N_978,In_216,In_918);
or U979 (N_979,In_948,In_450);
nand U980 (N_980,In_629,In_734);
nor U981 (N_981,In_256,In_25);
nor U982 (N_982,In_981,In_514);
nor U983 (N_983,In_195,In_77);
nand U984 (N_984,In_918,In_857);
or U985 (N_985,In_325,In_287);
and U986 (N_986,In_688,In_147);
or U987 (N_987,In_862,In_354);
or U988 (N_988,In_131,In_532);
and U989 (N_989,In_714,In_908);
or U990 (N_990,In_732,In_224);
nand U991 (N_991,In_508,In_950);
nand U992 (N_992,In_582,In_923);
or U993 (N_993,In_702,In_347);
nand U994 (N_994,In_78,In_255);
xnor U995 (N_995,In_650,In_892);
xnor U996 (N_996,In_99,In_706);
nor U997 (N_997,In_513,In_87);
nand U998 (N_998,In_13,In_31);
nor U999 (N_999,In_162,In_160);
nand U1000 (N_1000,In_863,In_527);
and U1001 (N_1001,In_90,In_565);
or U1002 (N_1002,In_646,In_248);
and U1003 (N_1003,In_759,In_425);
nand U1004 (N_1004,In_131,In_858);
and U1005 (N_1005,In_676,In_557);
nand U1006 (N_1006,In_73,In_95);
nand U1007 (N_1007,In_278,In_5);
or U1008 (N_1008,In_932,In_572);
and U1009 (N_1009,In_719,In_496);
or U1010 (N_1010,In_425,In_740);
or U1011 (N_1011,In_625,In_325);
or U1012 (N_1012,In_677,In_278);
nand U1013 (N_1013,In_241,In_525);
nand U1014 (N_1014,In_631,In_137);
and U1015 (N_1015,In_738,In_346);
nand U1016 (N_1016,In_875,In_804);
and U1017 (N_1017,In_433,In_464);
nand U1018 (N_1018,In_37,In_391);
or U1019 (N_1019,In_492,In_721);
or U1020 (N_1020,In_435,In_184);
nor U1021 (N_1021,In_230,In_916);
nor U1022 (N_1022,In_7,In_625);
nor U1023 (N_1023,In_912,In_302);
xnor U1024 (N_1024,In_876,In_254);
nand U1025 (N_1025,In_861,In_461);
or U1026 (N_1026,In_49,In_299);
or U1027 (N_1027,In_695,In_230);
and U1028 (N_1028,In_982,In_683);
or U1029 (N_1029,In_236,In_568);
nand U1030 (N_1030,In_136,In_996);
nand U1031 (N_1031,In_572,In_91);
nor U1032 (N_1032,In_372,In_227);
or U1033 (N_1033,In_47,In_924);
nor U1034 (N_1034,In_5,In_937);
nand U1035 (N_1035,In_149,In_108);
or U1036 (N_1036,In_806,In_519);
nor U1037 (N_1037,In_740,In_482);
nor U1038 (N_1038,In_688,In_766);
or U1039 (N_1039,In_254,In_364);
nand U1040 (N_1040,In_2,In_717);
nor U1041 (N_1041,In_651,In_572);
xor U1042 (N_1042,In_322,In_57);
and U1043 (N_1043,In_252,In_512);
and U1044 (N_1044,In_353,In_900);
nor U1045 (N_1045,In_484,In_79);
xnor U1046 (N_1046,In_291,In_32);
nor U1047 (N_1047,In_958,In_513);
and U1048 (N_1048,In_550,In_786);
or U1049 (N_1049,In_378,In_609);
nor U1050 (N_1050,In_409,In_725);
or U1051 (N_1051,In_251,In_682);
or U1052 (N_1052,In_260,In_635);
and U1053 (N_1053,In_554,In_933);
or U1054 (N_1054,In_886,In_441);
or U1055 (N_1055,In_93,In_327);
or U1056 (N_1056,In_842,In_456);
nor U1057 (N_1057,In_821,In_975);
nand U1058 (N_1058,In_971,In_360);
or U1059 (N_1059,In_684,In_620);
or U1060 (N_1060,In_956,In_728);
or U1061 (N_1061,In_144,In_246);
or U1062 (N_1062,In_98,In_147);
nand U1063 (N_1063,In_294,In_423);
nor U1064 (N_1064,In_966,In_489);
nor U1065 (N_1065,In_786,In_250);
and U1066 (N_1066,In_534,In_177);
nor U1067 (N_1067,In_607,In_16);
nor U1068 (N_1068,In_537,In_588);
nor U1069 (N_1069,In_56,In_9);
nor U1070 (N_1070,In_798,In_100);
or U1071 (N_1071,In_156,In_807);
and U1072 (N_1072,In_763,In_44);
nor U1073 (N_1073,In_227,In_239);
or U1074 (N_1074,In_440,In_109);
nand U1075 (N_1075,In_649,In_308);
and U1076 (N_1076,In_884,In_759);
nand U1077 (N_1077,In_272,In_981);
nor U1078 (N_1078,In_715,In_706);
nor U1079 (N_1079,In_421,In_626);
or U1080 (N_1080,In_113,In_24);
nor U1081 (N_1081,In_350,In_327);
or U1082 (N_1082,In_383,In_684);
nand U1083 (N_1083,In_494,In_88);
nor U1084 (N_1084,In_742,In_449);
xnor U1085 (N_1085,In_614,In_276);
and U1086 (N_1086,In_622,In_815);
nor U1087 (N_1087,In_126,In_782);
nand U1088 (N_1088,In_362,In_532);
or U1089 (N_1089,In_84,In_797);
or U1090 (N_1090,In_256,In_32);
or U1091 (N_1091,In_266,In_591);
nor U1092 (N_1092,In_496,In_392);
nand U1093 (N_1093,In_64,In_13);
nor U1094 (N_1094,In_527,In_459);
nand U1095 (N_1095,In_884,In_464);
or U1096 (N_1096,In_184,In_20);
or U1097 (N_1097,In_304,In_197);
or U1098 (N_1098,In_424,In_200);
xnor U1099 (N_1099,In_562,In_818);
nand U1100 (N_1100,In_397,In_492);
and U1101 (N_1101,In_515,In_709);
or U1102 (N_1102,In_163,In_300);
nor U1103 (N_1103,In_721,In_533);
or U1104 (N_1104,In_471,In_720);
or U1105 (N_1105,In_181,In_986);
nand U1106 (N_1106,In_756,In_836);
nor U1107 (N_1107,In_341,In_721);
or U1108 (N_1108,In_461,In_566);
and U1109 (N_1109,In_336,In_130);
xnor U1110 (N_1110,In_302,In_595);
nand U1111 (N_1111,In_823,In_260);
nor U1112 (N_1112,In_266,In_828);
or U1113 (N_1113,In_947,In_644);
and U1114 (N_1114,In_979,In_324);
or U1115 (N_1115,In_428,In_876);
xor U1116 (N_1116,In_204,In_158);
and U1117 (N_1117,In_460,In_517);
nor U1118 (N_1118,In_455,In_245);
or U1119 (N_1119,In_309,In_1);
and U1120 (N_1120,In_183,In_820);
and U1121 (N_1121,In_408,In_423);
or U1122 (N_1122,In_705,In_85);
and U1123 (N_1123,In_898,In_810);
nand U1124 (N_1124,In_235,In_723);
and U1125 (N_1125,In_959,In_120);
nand U1126 (N_1126,In_712,In_573);
and U1127 (N_1127,In_697,In_304);
and U1128 (N_1128,In_959,In_812);
and U1129 (N_1129,In_408,In_123);
nand U1130 (N_1130,In_894,In_332);
nor U1131 (N_1131,In_596,In_651);
or U1132 (N_1132,In_467,In_364);
nand U1133 (N_1133,In_405,In_245);
nor U1134 (N_1134,In_886,In_575);
nor U1135 (N_1135,In_794,In_717);
or U1136 (N_1136,In_995,In_283);
nand U1137 (N_1137,In_473,In_490);
nand U1138 (N_1138,In_108,In_634);
and U1139 (N_1139,In_10,In_460);
nand U1140 (N_1140,In_220,In_556);
nand U1141 (N_1141,In_456,In_990);
and U1142 (N_1142,In_148,In_4);
nor U1143 (N_1143,In_291,In_300);
or U1144 (N_1144,In_462,In_450);
nand U1145 (N_1145,In_120,In_721);
nor U1146 (N_1146,In_368,In_854);
nand U1147 (N_1147,In_944,In_608);
nand U1148 (N_1148,In_73,In_994);
and U1149 (N_1149,In_956,In_751);
and U1150 (N_1150,In_65,In_769);
xnor U1151 (N_1151,In_2,In_408);
or U1152 (N_1152,In_955,In_69);
nor U1153 (N_1153,In_672,In_458);
or U1154 (N_1154,In_215,In_541);
and U1155 (N_1155,In_889,In_502);
nor U1156 (N_1156,In_832,In_982);
and U1157 (N_1157,In_648,In_213);
and U1158 (N_1158,In_417,In_946);
or U1159 (N_1159,In_134,In_625);
nor U1160 (N_1160,In_767,In_76);
or U1161 (N_1161,In_478,In_385);
nor U1162 (N_1162,In_449,In_869);
nor U1163 (N_1163,In_351,In_145);
xnor U1164 (N_1164,In_929,In_937);
or U1165 (N_1165,In_490,In_61);
nand U1166 (N_1166,In_477,In_652);
nor U1167 (N_1167,In_717,In_220);
and U1168 (N_1168,In_665,In_129);
nor U1169 (N_1169,In_167,In_684);
xnor U1170 (N_1170,In_843,In_338);
or U1171 (N_1171,In_992,In_762);
or U1172 (N_1172,In_506,In_34);
and U1173 (N_1173,In_131,In_353);
or U1174 (N_1174,In_133,In_214);
or U1175 (N_1175,In_856,In_380);
nand U1176 (N_1176,In_629,In_253);
and U1177 (N_1177,In_626,In_323);
or U1178 (N_1178,In_274,In_284);
nand U1179 (N_1179,In_317,In_677);
or U1180 (N_1180,In_90,In_628);
nor U1181 (N_1181,In_953,In_450);
nand U1182 (N_1182,In_779,In_543);
or U1183 (N_1183,In_516,In_209);
or U1184 (N_1184,In_865,In_493);
nand U1185 (N_1185,In_256,In_693);
and U1186 (N_1186,In_173,In_935);
and U1187 (N_1187,In_668,In_767);
nor U1188 (N_1188,In_690,In_83);
or U1189 (N_1189,In_831,In_3);
and U1190 (N_1190,In_564,In_510);
and U1191 (N_1191,In_142,In_617);
nor U1192 (N_1192,In_114,In_307);
nand U1193 (N_1193,In_433,In_492);
nor U1194 (N_1194,In_403,In_29);
or U1195 (N_1195,In_664,In_561);
nor U1196 (N_1196,In_831,In_686);
nor U1197 (N_1197,In_976,In_884);
or U1198 (N_1198,In_928,In_601);
nand U1199 (N_1199,In_328,In_645);
nand U1200 (N_1200,In_9,In_681);
or U1201 (N_1201,In_873,In_778);
and U1202 (N_1202,In_122,In_131);
or U1203 (N_1203,In_680,In_137);
or U1204 (N_1204,In_841,In_743);
nor U1205 (N_1205,In_859,In_117);
and U1206 (N_1206,In_868,In_150);
nand U1207 (N_1207,In_979,In_55);
and U1208 (N_1208,In_114,In_58);
nand U1209 (N_1209,In_794,In_679);
or U1210 (N_1210,In_125,In_504);
nor U1211 (N_1211,In_584,In_553);
xor U1212 (N_1212,In_388,In_183);
or U1213 (N_1213,In_296,In_335);
nand U1214 (N_1214,In_865,In_170);
nor U1215 (N_1215,In_934,In_238);
and U1216 (N_1216,In_615,In_762);
or U1217 (N_1217,In_111,In_700);
or U1218 (N_1218,In_84,In_149);
nor U1219 (N_1219,In_59,In_280);
nand U1220 (N_1220,In_12,In_812);
nor U1221 (N_1221,In_245,In_493);
and U1222 (N_1222,In_137,In_922);
or U1223 (N_1223,In_623,In_147);
and U1224 (N_1224,In_395,In_524);
or U1225 (N_1225,In_592,In_187);
or U1226 (N_1226,In_596,In_285);
nor U1227 (N_1227,In_399,In_40);
nand U1228 (N_1228,In_346,In_971);
or U1229 (N_1229,In_629,In_376);
nor U1230 (N_1230,In_196,In_599);
nor U1231 (N_1231,In_266,In_924);
nand U1232 (N_1232,In_377,In_156);
nand U1233 (N_1233,In_224,In_767);
or U1234 (N_1234,In_982,In_983);
nor U1235 (N_1235,In_19,In_755);
or U1236 (N_1236,In_141,In_350);
nand U1237 (N_1237,In_452,In_110);
nor U1238 (N_1238,In_506,In_944);
nand U1239 (N_1239,In_594,In_757);
and U1240 (N_1240,In_691,In_106);
and U1241 (N_1241,In_614,In_147);
nand U1242 (N_1242,In_922,In_737);
or U1243 (N_1243,In_850,In_874);
nor U1244 (N_1244,In_540,In_858);
nor U1245 (N_1245,In_285,In_733);
nor U1246 (N_1246,In_202,In_777);
nor U1247 (N_1247,In_70,In_836);
and U1248 (N_1248,In_882,In_725);
or U1249 (N_1249,In_37,In_456);
nor U1250 (N_1250,In_929,In_359);
or U1251 (N_1251,In_874,In_503);
or U1252 (N_1252,In_330,In_243);
nor U1253 (N_1253,In_72,In_981);
and U1254 (N_1254,In_666,In_321);
nand U1255 (N_1255,In_806,In_134);
and U1256 (N_1256,In_625,In_971);
and U1257 (N_1257,In_541,In_22);
or U1258 (N_1258,In_511,In_816);
or U1259 (N_1259,In_873,In_717);
or U1260 (N_1260,In_730,In_503);
or U1261 (N_1261,In_335,In_636);
xor U1262 (N_1262,In_490,In_420);
nor U1263 (N_1263,In_759,In_631);
nor U1264 (N_1264,In_886,In_80);
nor U1265 (N_1265,In_658,In_533);
nand U1266 (N_1266,In_662,In_944);
nor U1267 (N_1267,In_465,In_245);
or U1268 (N_1268,In_713,In_274);
and U1269 (N_1269,In_671,In_973);
xnor U1270 (N_1270,In_471,In_402);
nand U1271 (N_1271,In_368,In_557);
and U1272 (N_1272,In_182,In_849);
nand U1273 (N_1273,In_959,In_988);
nand U1274 (N_1274,In_741,In_719);
nor U1275 (N_1275,In_478,In_400);
and U1276 (N_1276,In_415,In_910);
and U1277 (N_1277,In_843,In_863);
or U1278 (N_1278,In_850,In_455);
and U1279 (N_1279,In_40,In_98);
nand U1280 (N_1280,In_614,In_316);
nor U1281 (N_1281,In_548,In_659);
nand U1282 (N_1282,In_447,In_419);
nand U1283 (N_1283,In_731,In_412);
nor U1284 (N_1284,In_922,In_570);
and U1285 (N_1285,In_350,In_860);
nand U1286 (N_1286,In_392,In_215);
or U1287 (N_1287,In_593,In_116);
and U1288 (N_1288,In_108,In_657);
nor U1289 (N_1289,In_502,In_933);
and U1290 (N_1290,In_648,In_292);
and U1291 (N_1291,In_82,In_982);
xor U1292 (N_1292,In_182,In_773);
or U1293 (N_1293,In_856,In_979);
nand U1294 (N_1294,In_147,In_251);
or U1295 (N_1295,In_573,In_231);
or U1296 (N_1296,In_361,In_950);
and U1297 (N_1297,In_311,In_611);
nor U1298 (N_1298,In_207,In_125);
nor U1299 (N_1299,In_756,In_476);
or U1300 (N_1300,In_262,In_847);
or U1301 (N_1301,In_85,In_990);
nor U1302 (N_1302,In_773,In_894);
nor U1303 (N_1303,In_51,In_341);
xnor U1304 (N_1304,In_669,In_299);
and U1305 (N_1305,In_517,In_710);
nand U1306 (N_1306,In_740,In_361);
and U1307 (N_1307,In_808,In_827);
nand U1308 (N_1308,In_656,In_819);
and U1309 (N_1309,In_620,In_332);
and U1310 (N_1310,In_838,In_197);
or U1311 (N_1311,In_111,In_69);
and U1312 (N_1312,In_754,In_617);
nand U1313 (N_1313,In_508,In_709);
nand U1314 (N_1314,In_862,In_650);
nor U1315 (N_1315,In_969,In_859);
or U1316 (N_1316,In_164,In_511);
nand U1317 (N_1317,In_953,In_569);
nor U1318 (N_1318,In_825,In_908);
and U1319 (N_1319,In_247,In_492);
nand U1320 (N_1320,In_531,In_320);
nand U1321 (N_1321,In_24,In_363);
nor U1322 (N_1322,In_721,In_645);
and U1323 (N_1323,In_714,In_922);
or U1324 (N_1324,In_321,In_609);
and U1325 (N_1325,In_239,In_651);
and U1326 (N_1326,In_733,In_588);
or U1327 (N_1327,In_373,In_334);
or U1328 (N_1328,In_776,In_352);
nor U1329 (N_1329,In_709,In_422);
and U1330 (N_1330,In_855,In_219);
nor U1331 (N_1331,In_227,In_974);
nand U1332 (N_1332,In_584,In_642);
nand U1333 (N_1333,In_659,In_599);
nor U1334 (N_1334,In_498,In_390);
or U1335 (N_1335,In_370,In_202);
and U1336 (N_1336,In_762,In_372);
nor U1337 (N_1337,In_577,In_368);
and U1338 (N_1338,In_312,In_336);
or U1339 (N_1339,In_385,In_53);
and U1340 (N_1340,In_269,In_699);
or U1341 (N_1341,In_406,In_688);
nor U1342 (N_1342,In_530,In_55);
or U1343 (N_1343,In_87,In_58);
or U1344 (N_1344,In_579,In_411);
nand U1345 (N_1345,In_733,In_903);
or U1346 (N_1346,In_398,In_563);
nor U1347 (N_1347,In_925,In_648);
nor U1348 (N_1348,In_480,In_376);
nand U1349 (N_1349,In_472,In_561);
and U1350 (N_1350,In_725,In_177);
or U1351 (N_1351,In_707,In_200);
nand U1352 (N_1352,In_985,In_426);
nor U1353 (N_1353,In_169,In_745);
nand U1354 (N_1354,In_73,In_261);
or U1355 (N_1355,In_714,In_69);
nor U1356 (N_1356,In_952,In_267);
nand U1357 (N_1357,In_268,In_59);
and U1358 (N_1358,In_21,In_549);
or U1359 (N_1359,In_64,In_464);
nor U1360 (N_1360,In_416,In_52);
or U1361 (N_1361,In_660,In_90);
and U1362 (N_1362,In_15,In_278);
nor U1363 (N_1363,In_177,In_697);
or U1364 (N_1364,In_901,In_790);
nor U1365 (N_1365,In_305,In_774);
nor U1366 (N_1366,In_740,In_703);
nand U1367 (N_1367,In_412,In_448);
nand U1368 (N_1368,In_138,In_318);
or U1369 (N_1369,In_820,In_930);
nand U1370 (N_1370,In_710,In_778);
nand U1371 (N_1371,In_926,In_325);
nor U1372 (N_1372,In_951,In_997);
and U1373 (N_1373,In_218,In_842);
nand U1374 (N_1374,In_192,In_514);
and U1375 (N_1375,In_808,In_149);
or U1376 (N_1376,In_646,In_887);
or U1377 (N_1377,In_582,In_526);
or U1378 (N_1378,In_223,In_901);
nor U1379 (N_1379,In_41,In_137);
or U1380 (N_1380,In_432,In_255);
nand U1381 (N_1381,In_146,In_554);
and U1382 (N_1382,In_192,In_425);
or U1383 (N_1383,In_694,In_826);
or U1384 (N_1384,In_416,In_603);
or U1385 (N_1385,In_570,In_558);
nor U1386 (N_1386,In_889,In_76);
nand U1387 (N_1387,In_94,In_909);
nand U1388 (N_1388,In_639,In_656);
and U1389 (N_1389,In_706,In_865);
and U1390 (N_1390,In_33,In_855);
and U1391 (N_1391,In_78,In_867);
nor U1392 (N_1392,In_87,In_6);
nor U1393 (N_1393,In_975,In_954);
nor U1394 (N_1394,In_778,In_90);
nand U1395 (N_1395,In_282,In_760);
or U1396 (N_1396,In_415,In_496);
or U1397 (N_1397,In_555,In_392);
or U1398 (N_1398,In_587,In_525);
and U1399 (N_1399,In_890,In_845);
nor U1400 (N_1400,In_81,In_656);
and U1401 (N_1401,In_919,In_654);
or U1402 (N_1402,In_427,In_654);
nor U1403 (N_1403,In_597,In_111);
or U1404 (N_1404,In_436,In_213);
and U1405 (N_1405,In_394,In_913);
nand U1406 (N_1406,In_326,In_594);
nor U1407 (N_1407,In_588,In_750);
nor U1408 (N_1408,In_437,In_955);
nand U1409 (N_1409,In_754,In_383);
and U1410 (N_1410,In_1,In_555);
or U1411 (N_1411,In_831,In_886);
nor U1412 (N_1412,In_524,In_62);
and U1413 (N_1413,In_602,In_580);
nor U1414 (N_1414,In_491,In_901);
and U1415 (N_1415,In_349,In_997);
and U1416 (N_1416,In_861,In_186);
or U1417 (N_1417,In_140,In_119);
and U1418 (N_1418,In_704,In_815);
nor U1419 (N_1419,In_759,In_47);
nor U1420 (N_1420,In_518,In_937);
nor U1421 (N_1421,In_278,In_332);
or U1422 (N_1422,In_395,In_73);
nor U1423 (N_1423,In_96,In_39);
nor U1424 (N_1424,In_919,In_381);
nand U1425 (N_1425,In_159,In_614);
or U1426 (N_1426,In_764,In_710);
and U1427 (N_1427,In_72,In_268);
nor U1428 (N_1428,In_795,In_908);
nand U1429 (N_1429,In_274,In_558);
nand U1430 (N_1430,In_320,In_312);
and U1431 (N_1431,In_737,In_846);
or U1432 (N_1432,In_631,In_27);
and U1433 (N_1433,In_537,In_611);
nor U1434 (N_1434,In_796,In_706);
nor U1435 (N_1435,In_45,In_155);
nor U1436 (N_1436,In_645,In_460);
nor U1437 (N_1437,In_779,In_431);
nand U1438 (N_1438,In_122,In_329);
or U1439 (N_1439,In_138,In_292);
and U1440 (N_1440,In_415,In_205);
nor U1441 (N_1441,In_309,In_946);
nor U1442 (N_1442,In_65,In_689);
and U1443 (N_1443,In_914,In_147);
or U1444 (N_1444,In_417,In_954);
nand U1445 (N_1445,In_388,In_950);
nand U1446 (N_1446,In_24,In_182);
nand U1447 (N_1447,In_486,In_607);
and U1448 (N_1448,In_880,In_48);
nor U1449 (N_1449,In_943,In_631);
nor U1450 (N_1450,In_219,In_253);
and U1451 (N_1451,In_242,In_90);
or U1452 (N_1452,In_773,In_429);
nor U1453 (N_1453,In_98,In_864);
nor U1454 (N_1454,In_253,In_516);
or U1455 (N_1455,In_988,In_413);
nor U1456 (N_1456,In_989,In_978);
and U1457 (N_1457,In_245,In_775);
or U1458 (N_1458,In_680,In_834);
or U1459 (N_1459,In_954,In_143);
nand U1460 (N_1460,In_892,In_988);
nand U1461 (N_1461,In_643,In_196);
or U1462 (N_1462,In_288,In_65);
nand U1463 (N_1463,In_867,In_891);
and U1464 (N_1464,In_270,In_120);
nand U1465 (N_1465,In_123,In_721);
nor U1466 (N_1466,In_74,In_210);
or U1467 (N_1467,In_696,In_554);
nor U1468 (N_1468,In_474,In_605);
nand U1469 (N_1469,In_81,In_433);
nor U1470 (N_1470,In_390,In_433);
nand U1471 (N_1471,In_758,In_634);
or U1472 (N_1472,In_68,In_598);
and U1473 (N_1473,In_266,In_532);
nor U1474 (N_1474,In_430,In_699);
nand U1475 (N_1475,In_694,In_147);
nand U1476 (N_1476,In_332,In_870);
and U1477 (N_1477,In_276,In_56);
nand U1478 (N_1478,In_259,In_74);
and U1479 (N_1479,In_559,In_918);
nor U1480 (N_1480,In_299,In_421);
or U1481 (N_1481,In_57,In_71);
or U1482 (N_1482,In_237,In_360);
nor U1483 (N_1483,In_111,In_878);
nor U1484 (N_1484,In_110,In_618);
nand U1485 (N_1485,In_86,In_732);
or U1486 (N_1486,In_631,In_74);
nand U1487 (N_1487,In_752,In_100);
or U1488 (N_1488,In_5,In_110);
nand U1489 (N_1489,In_444,In_472);
nor U1490 (N_1490,In_514,In_769);
and U1491 (N_1491,In_825,In_20);
nand U1492 (N_1492,In_924,In_935);
nand U1493 (N_1493,In_697,In_406);
nor U1494 (N_1494,In_166,In_336);
nand U1495 (N_1495,In_379,In_644);
nand U1496 (N_1496,In_332,In_283);
or U1497 (N_1497,In_680,In_870);
nor U1498 (N_1498,In_669,In_853);
nand U1499 (N_1499,In_310,In_436);
or U1500 (N_1500,In_357,In_662);
and U1501 (N_1501,In_30,In_501);
and U1502 (N_1502,In_737,In_200);
and U1503 (N_1503,In_265,In_537);
nor U1504 (N_1504,In_40,In_224);
nor U1505 (N_1505,In_980,In_363);
xor U1506 (N_1506,In_890,In_268);
nor U1507 (N_1507,In_53,In_268);
nor U1508 (N_1508,In_200,In_33);
nor U1509 (N_1509,In_993,In_303);
or U1510 (N_1510,In_487,In_310);
nor U1511 (N_1511,In_770,In_72);
and U1512 (N_1512,In_683,In_271);
and U1513 (N_1513,In_534,In_565);
and U1514 (N_1514,In_240,In_290);
or U1515 (N_1515,In_488,In_866);
and U1516 (N_1516,In_857,In_868);
nand U1517 (N_1517,In_987,In_826);
nor U1518 (N_1518,In_196,In_84);
and U1519 (N_1519,In_318,In_720);
nor U1520 (N_1520,In_647,In_675);
nand U1521 (N_1521,In_261,In_311);
and U1522 (N_1522,In_85,In_347);
nand U1523 (N_1523,In_427,In_553);
nor U1524 (N_1524,In_869,In_740);
nor U1525 (N_1525,In_846,In_621);
or U1526 (N_1526,In_970,In_590);
or U1527 (N_1527,In_395,In_286);
and U1528 (N_1528,In_26,In_323);
nand U1529 (N_1529,In_185,In_675);
or U1530 (N_1530,In_935,In_550);
or U1531 (N_1531,In_145,In_813);
or U1532 (N_1532,In_296,In_899);
nor U1533 (N_1533,In_846,In_263);
nor U1534 (N_1534,In_667,In_288);
or U1535 (N_1535,In_646,In_561);
nand U1536 (N_1536,In_937,In_250);
nor U1537 (N_1537,In_505,In_319);
nor U1538 (N_1538,In_797,In_688);
nor U1539 (N_1539,In_944,In_159);
or U1540 (N_1540,In_45,In_173);
nand U1541 (N_1541,In_491,In_988);
or U1542 (N_1542,In_311,In_868);
nor U1543 (N_1543,In_568,In_356);
xor U1544 (N_1544,In_160,In_89);
xnor U1545 (N_1545,In_141,In_149);
nor U1546 (N_1546,In_197,In_617);
nand U1547 (N_1547,In_371,In_0);
and U1548 (N_1548,In_268,In_260);
nand U1549 (N_1549,In_603,In_787);
nor U1550 (N_1550,In_520,In_522);
or U1551 (N_1551,In_88,In_158);
and U1552 (N_1552,In_562,In_368);
nand U1553 (N_1553,In_343,In_39);
nor U1554 (N_1554,In_545,In_726);
nand U1555 (N_1555,In_938,In_607);
nand U1556 (N_1556,In_101,In_667);
or U1557 (N_1557,In_105,In_602);
nor U1558 (N_1558,In_732,In_926);
or U1559 (N_1559,In_66,In_915);
and U1560 (N_1560,In_25,In_137);
nor U1561 (N_1561,In_651,In_197);
and U1562 (N_1562,In_620,In_126);
nor U1563 (N_1563,In_926,In_505);
nand U1564 (N_1564,In_214,In_712);
or U1565 (N_1565,In_623,In_783);
nand U1566 (N_1566,In_476,In_871);
nor U1567 (N_1567,In_852,In_389);
nor U1568 (N_1568,In_226,In_169);
nand U1569 (N_1569,In_907,In_20);
nor U1570 (N_1570,In_774,In_859);
nor U1571 (N_1571,In_408,In_150);
and U1572 (N_1572,In_264,In_75);
nand U1573 (N_1573,In_644,In_543);
and U1574 (N_1574,In_488,In_718);
or U1575 (N_1575,In_683,In_817);
or U1576 (N_1576,In_610,In_247);
nand U1577 (N_1577,In_447,In_580);
and U1578 (N_1578,In_774,In_654);
nor U1579 (N_1579,In_441,In_878);
nor U1580 (N_1580,In_263,In_838);
nand U1581 (N_1581,In_589,In_918);
or U1582 (N_1582,In_222,In_299);
nor U1583 (N_1583,In_887,In_589);
nand U1584 (N_1584,In_344,In_639);
or U1585 (N_1585,In_392,In_212);
xnor U1586 (N_1586,In_505,In_258);
nor U1587 (N_1587,In_150,In_149);
and U1588 (N_1588,In_271,In_898);
nand U1589 (N_1589,In_927,In_522);
or U1590 (N_1590,In_16,In_992);
and U1591 (N_1591,In_10,In_103);
nand U1592 (N_1592,In_980,In_421);
nor U1593 (N_1593,In_23,In_549);
or U1594 (N_1594,In_318,In_66);
nand U1595 (N_1595,In_976,In_660);
and U1596 (N_1596,In_790,In_733);
nand U1597 (N_1597,In_622,In_852);
or U1598 (N_1598,In_56,In_290);
nand U1599 (N_1599,In_861,In_660);
nor U1600 (N_1600,In_390,In_664);
nand U1601 (N_1601,In_94,In_505);
xor U1602 (N_1602,In_692,In_452);
and U1603 (N_1603,In_885,In_986);
and U1604 (N_1604,In_690,In_308);
or U1605 (N_1605,In_900,In_118);
nand U1606 (N_1606,In_632,In_378);
and U1607 (N_1607,In_858,In_311);
or U1608 (N_1608,In_703,In_899);
or U1609 (N_1609,In_538,In_744);
and U1610 (N_1610,In_391,In_680);
or U1611 (N_1611,In_444,In_92);
and U1612 (N_1612,In_721,In_445);
nor U1613 (N_1613,In_331,In_854);
or U1614 (N_1614,In_353,In_884);
nor U1615 (N_1615,In_60,In_655);
or U1616 (N_1616,In_100,In_217);
and U1617 (N_1617,In_762,In_787);
or U1618 (N_1618,In_375,In_431);
nor U1619 (N_1619,In_990,In_209);
xnor U1620 (N_1620,In_38,In_519);
and U1621 (N_1621,In_554,In_203);
nor U1622 (N_1622,In_350,In_491);
and U1623 (N_1623,In_337,In_253);
or U1624 (N_1624,In_991,In_484);
nand U1625 (N_1625,In_254,In_197);
nor U1626 (N_1626,In_118,In_385);
nor U1627 (N_1627,In_394,In_13);
nor U1628 (N_1628,In_709,In_857);
xnor U1629 (N_1629,In_125,In_91);
nand U1630 (N_1630,In_645,In_704);
nand U1631 (N_1631,In_963,In_422);
nor U1632 (N_1632,In_764,In_890);
and U1633 (N_1633,In_882,In_71);
nor U1634 (N_1634,In_523,In_735);
nand U1635 (N_1635,In_684,In_204);
nor U1636 (N_1636,In_322,In_592);
nor U1637 (N_1637,In_930,In_135);
nor U1638 (N_1638,In_739,In_456);
and U1639 (N_1639,In_243,In_366);
nand U1640 (N_1640,In_425,In_525);
nor U1641 (N_1641,In_576,In_301);
xor U1642 (N_1642,In_483,In_258);
nand U1643 (N_1643,In_565,In_656);
xnor U1644 (N_1644,In_154,In_657);
or U1645 (N_1645,In_672,In_260);
and U1646 (N_1646,In_921,In_221);
and U1647 (N_1647,In_453,In_892);
and U1648 (N_1648,In_986,In_826);
or U1649 (N_1649,In_432,In_463);
and U1650 (N_1650,In_614,In_434);
nor U1651 (N_1651,In_78,In_419);
nor U1652 (N_1652,In_284,In_105);
or U1653 (N_1653,In_143,In_981);
and U1654 (N_1654,In_233,In_44);
nand U1655 (N_1655,In_527,In_446);
and U1656 (N_1656,In_940,In_102);
and U1657 (N_1657,In_213,In_350);
and U1658 (N_1658,In_400,In_356);
nor U1659 (N_1659,In_511,In_972);
or U1660 (N_1660,In_281,In_511);
and U1661 (N_1661,In_588,In_827);
nand U1662 (N_1662,In_730,In_641);
and U1663 (N_1663,In_535,In_172);
nor U1664 (N_1664,In_123,In_598);
and U1665 (N_1665,In_572,In_405);
nand U1666 (N_1666,In_867,In_883);
or U1667 (N_1667,In_120,In_399);
or U1668 (N_1668,In_579,In_164);
and U1669 (N_1669,In_745,In_718);
xnor U1670 (N_1670,In_40,In_107);
and U1671 (N_1671,In_488,In_117);
nand U1672 (N_1672,In_134,In_101);
or U1673 (N_1673,In_145,In_246);
or U1674 (N_1674,In_388,In_158);
nor U1675 (N_1675,In_974,In_31);
nand U1676 (N_1676,In_375,In_990);
nor U1677 (N_1677,In_414,In_47);
nor U1678 (N_1678,In_475,In_666);
nor U1679 (N_1679,In_525,In_973);
nor U1680 (N_1680,In_831,In_659);
or U1681 (N_1681,In_758,In_29);
nand U1682 (N_1682,In_44,In_434);
nand U1683 (N_1683,In_775,In_4);
or U1684 (N_1684,In_90,In_326);
and U1685 (N_1685,In_312,In_237);
and U1686 (N_1686,In_339,In_925);
xor U1687 (N_1687,In_609,In_714);
and U1688 (N_1688,In_569,In_84);
nand U1689 (N_1689,In_882,In_417);
nand U1690 (N_1690,In_160,In_375);
and U1691 (N_1691,In_201,In_298);
nor U1692 (N_1692,In_315,In_787);
nand U1693 (N_1693,In_816,In_683);
and U1694 (N_1694,In_303,In_228);
and U1695 (N_1695,In_499,In_858);
or U1696 (N_1696,In_195,In_693);
nor U1697 (N_1697,In_151,In_321);
or U1698 (N_1698,In_740,In_629);
and U1699 (N_1699,In_451,In_412);
or U1700 (N_1700,In_998,In_700);
nor U1701 (N_1701,In_915,In_2);
or U1702 (N_1702,In_943,In_178);
nor U1703 (N_1703,In_475,In_420);
nor U1704 (N_1704,In_113,In_969);
and U1705 (N_1705,In_994,In_629);
and U1706 (N_1706,In_372,In_271);
nand U1707 (N_1707,In_922,In_305);
nor U1708 (N_1708,In_765,In_560);
nor U1709 (N_1709,In_309,In_451);
nand U1710 (N_1710,In_300,In_498);
and U1711 (N_1711,In_368,In_387);
and U1712 (N_1712,In_549,In_860);
xnor U1713 (N_1713,In_334,In_445);
nor U1714 (N_1714,In_879,In_864);
and U1715 (N_1715,In_115,In_484);
nand U1716 (N_1716,In_719,In_725);
nor U1717 (N_1717,In_771,In_863);
nand U1718 (N_1718,In_680,In_975);
nor U1719 (N_1719,In_62,In_720);
nor U1720 (N_1720,In_486,In_688);
nand U1721 (N_1721,In_295,In_422);
or U1722 (N_1722,In_749,In_200);
and U1723 (N_1723,In_85,In_251);
and U1724 (N_1724,In_59,In_702);
nor U1725 (N_1725,In_962,In_649);
nand U1726 (N_1726,In_412,In_443);
or U1727 (N_1727,In_864,In_39);
and U1728 (N_1728,In_60,In_313);
xnor U1729 (N_1729,In_985,In_756);
nor U1730 (N_1730,In_462,In_208);
and U1731 (N_1731,In_226,In_582);
nor U1732 (N_1732,In_313,In_331);
nand U1733 (N_1733,In_923,In_555);
nor U1734 (N_1734,In_969,In_239);
or U1735 (N_1735,In_473,In_496);
and U1736 (N_1736,In_259,In_257);
or U1737 (N_1737,In_674,In_105);
and U1738 (N_1738,In_473,In_902);
and U1739 (N_1739,In_783,In_894);
nor U1740 (N_1740,In_894,In_991);
nor U1741 (N_1741,In_506,In_78);
nand U1742 (N_1742,In_243,In_630);
or U1743 (N_1743,In_820,In_99);
and U1744 (N_1744,In_718,In_785);
nand U1745 (N_1745,In_453,In_290);
nor U1746 (N_1746,In_304,In_431);
and U1747 (N_1747,In_856,In_877);
or U1748 (N_1748,In_482,In_89);
nand U1749 (N_1749,In_332,In_889);
nor U1750 (N_1750,In_133,In_838);
nor U1751 (N_1751,In_103,In_831);
and U1752 (N_1752,In_855,In_266);
and U1753 (N_1753,In_345,In_652);
and U1754 (N_1754,In_864,In_836);
or U1755 (N_1755,In_728,In_452);
or U1756 (N_1756,In_197,In_876);
or U1757 (N_1757,In_735,In_640);
nor U1758 (N_1758,In_103,In_526);
nand U1759 (N_1759,In_177,In_107);
or U1760 (N_1760,In_746,In_313);
xnor U1761 (N_1761,In_242,In_632);
nand U1762 (N_1762,In_257,In_212);
nand U1763 (N_1763,In_493,In_299);
or U1764 (N_1764,In_885,In_994);
nand U1765 (N_1765,In_267,In_472);
nand U1766 (N_1766,In_54,In_92);
nor U1767 (N_1767,In_410,In_858);
or U1768 (N_1768,In_535,In_583);
nand U1769 (N_1769,In_975,In_848);
nor U1770 (N_1770,In_4,In_640);
and U1771 (N_1771,In_11,In_810);
or U1772 (N_1772,In_116,In_297);
or U1773 (N_1773,In_843,In_320);
nand U1774 (N_1774,In_854,In_118);
nand U1775 (N_1775,In_236,In_801);
or U1776 (N_1776,In_264,In_6);
nand U1777 (N_1777,In_69,In_777);
nand U1778 (N_1778,In_992,In_543);
nand U1779 (N_1779,In_795,In_836);
xnor U1780 (N_1780,In_55,In_878);
nor U1781 (N_1781,In_70,In_363);
nor U1782 (N_1782,In_271,In_207);
nor U1783 (N_1783,In_742,In_223);
nand U1784 (N_1784,In_112,In_64);
nor U1785 (N_1785,In_198,In_683);
and U1786 (N_1786,In_143,In_701);
nor U1787 (N_1787,In_98,In_857);
and U1788 (N_1788,In_808,In_346);
xnor U1789 (N_1789,In_319,In_27);
and U1790 (N_1790,In_21,In_526);
nor U1791 (N_1791,In_367,In_49);
and U1792 (N_1792,In_583,In_245);
or U1793 (N_1793,In_593,In_564);
or U1794 (N_1794,In_615,In_383);
nand U1795 (N_1795,In_504,In_967);
or U1796 (N_1796,In_760,In_481);
nor U1797 (N_1797,In_203,In_199);
nand U1798 (N_1798,In_289,In_831);
nand U1799 (N_1799,In_882,In_650);
nand U1800 (N_1800,In_843,In_658);
and U1801 (N_1801,In_446,In_707);
nor U1802 (N_1802,In_744,In_231);
or U1803 (N_1803,In_86,In_859);
nor U1804 (N_1804,In_118,In_456);
or U1805 (N_1805,In_532,In_760);
or U1806 (N_1806,In_230,In_913);
nor U1807 (N_1807,In_645,In_936);
nor U1808 (N_1808,In_987,In_310);
nor U1809 (N_1809,In_980,In_288);
nor U1810 (N_1810,In_508,In_328);
nand U1811 (N_1811,In_752,In_524);
or U1812 (N_1812,In_84,In_867);
and U1813 (N_1813,In_249,In_163);
nand U1814 (N_1814,In_208,In_626);
nand U1815 (N_1815,In_621,In_446);
xnor U1816 (N_1816,In_717,In_162);
nor U1817 (N_1817,In_390,In_245);
or U1818 (N_1818,In_934,In_110);
and U1819 (N_1819,In_138,In_859);
nor U1820 (N_1820,In_392,In_936);
and U1821 (N_1821,In_921,In_400);
and U1822 (N_1822,In_722,In_961);
nor U1823 (N_1823,In_641,In_218);
and U1824 (N_1824,In_125,In_550);
or U1825 (N_1825,In_344,In_980);
nand U1826 (N_1826,In_961,In_480);
nor U1827 (N_1827,In_410,In_9);
nor U1828 (N_1828,In_962,In_930);
nand U1829 (N_1829,In_507,In_416);
nor U1830 (N_1830,In_910,In_363);
or U1831 (N_1831,In_217,In_971);
and U1832 (N_1832,In_802,In_262);
or U1833 (N_1833,In_242,In_125);
or U1834 (N_1834,In_822,In_76);
or U1835 (N_1835,In_395,In_45);
nand U1836 (N_1836,In_659,In_407);
nand U1837 (N_1837,In_130,In_768);
nand U1838 (N_1838,In_480,In_619);
nor U1839 (N_1839,In_152,In_668);
nand U1840 (N_1840,In_889,In_807);
or U1841 (N_1841,In_930,In_439);
nand U1842 (N_1842,In_765,In_413);
and U1843 (N_1843,In_575,In_24);
nand U1844 (N_1844,In_243,In_341);
or U1845 (N_1845,In_299,In_593);
nand U1846 (N_1846,In_966,In_670);
nand U1847 (N_1847,In_693,In_604);
nor U1848 (N_1848,In_297,In_461);
or U1849 (N_1849,In_680,In_999);
xor U1850 (N_1850,In_885,In_572);
nor U1851 (N_1851,In_863,In_737);
and U1852 (N_1852,In_0,In_250);
nor U1853 (N_1853,In_713,In_183);
or U1854 (N_1854,In_418,In_995);
or U1855 (N_1855,In_366,In_493);
nand U1856 (N_1856,In_684,In_528);
or U1857 (N_1857,In_956,In_631);
and U1858 (N_1858,In_661,In_156);
and U1859 (N_1859,In_953,In_140);
nor U1860 (N_1860,In_254,In_726);
and U1861 (N_1861,In_955,In_97);
nand U1862 (N_1862,In_49,In_17);
or U1863 (N_1863,In_858,In_612);
or U1864 (N_1864,In_115,In_513);
nand U1865 (N_1865,In_175,In_440);
xor U1866 (N_1866,In_226,In_350);
nand U1867 (N_1867,In_279,In_208);
nor U1868 (N_1868,In_302,In_738);
nor U1869 (N_1869,In_440,In_599);
or U1870 (N_1870,In_603,In_309);
and U1871 (N_1871,In_476,In_334);
or U1872 (N_1872,In_590,In_450);
nor U1873 (N_1873,In_750,In_132);
xor U1874 (N_1874,In_516,In_910);
nand U1875 (N_1875,In_97,In_681);
and U1876 (N_1876,In_4,In_707);
or U1877 (N_1877,In_342,In_542);
and U1878 (N_1878,In_757,In_881);
or U1879 (N_1879,In_874,In_815);
or U1880 (N_1880,In_171,In_782);
nor U1881 (N_1881,In_546,In_815);
or U1882 (N_1882,In_777,In_899);
nor U1883 (N_1883,In_28,In_283);
or U1884 (N_1884,In_715,In_144);
nor U1885 (N_1885,In_550,In_560);
nor U1886 (N_1886,In_345,In_836);
and U1887 (N_1887,In_444,In_139);
and U1888 (N_1888,In_439,In_4);
or U1889 (N_1889,In_3,In_778);
nor U1890 (N_1890,In_257,In_60);
or U1891 (N_1891,In_216,In_819);
nor U1892 (N_1892,In_636,In_909);
nor U1893 (N_1893,In_263,In_370);
or U1894 (N_1894,In_258,In_795);
nor U1895 (N_1895,In_765,In_896);
and U1896 (N_1896,In_690,In_391);
nor U1897 (N_1897,In_762,In_224);
nor U1898 (N_1898,In_919,In_360);
nor U1899 (N_1899,In_16,In_418);
or U1900 (N_1900,In_443,In_950);
or U1901 (N_1901,In_819,In_731);
nand U1902 (N_1902,In_217,In_107);
xnor U1903 (N_1903,In_507,In_239);
nand U1904 (N_1904,In_851,In_932);
nor U1905 (N_1905,In_772,In_265);
nand U1906 (N_1906,In_322,In_665);
or U1907 (N_1907,In_863,In_672);
nor U1908 (N_1908,In_905,In_290);
or U1909 (N_1909,In_197,In_310);
nand U1910 (N_1910,In_697,In_232);
or U1911 (N_1911,In_35,In_999);
or U1912 (N_1912,In_101,In_521);
or U1913 (N_1913,In_801,In_401);
nand U1914 (N_1914,In_637,In_876);
nor U1915 (N_1915,In_694,In_906);
nor U1916 (N_1916,In_301,In_538);
nand U1917 (N_1917,In_142,In_55);
nand U1918 (N_1918,In_666,In_539);
nor U1919 (N_1919,In_777,In_629);
or U1920 (N_1920,In_160,In_874);
nand U1921 (N_1921,In_8,In_7);
nand U1922 (N_1922,In_388,In_144);
nand U1923 (N_1923,In_519,In_276);
and U1924 (N_1924,In_526,In_105);
nand U1925 (N_1925,In_489,In_627);
nand U1926 (N_1926,In_80,In_626);
and U1927 (N_1927,In_568,In_912);
nor U1928 (N_1928,In_223,In_548);
nand U1929 (N_1929,In_34,In_858);
and U1930 (N_1930,In_333,In_728);
nor U1931 (N_1931,In_347,In_932);
and U1932 (N_1932,In_593,In_339);
nand U1933 (N_1933,In_408,In_161);
nor U1934 (N_1934,In_850,In_929);
or U1935 (N_1935,In_550,In_706);
nand U1936 (N_1936,In_845,In_821);
xor U1937 (N_1937,In_657,In_454);
and U1938 (N_1938,In_684,In_22);
nand U1939 (N_1939,In_10,In_184);
and U1940 (N_1940,In_281,In_89);
nand U1941 (N_1941,In_999,In_632);
and U1942 (N_1942,In_802,In_249);
nand U1943 (N_1943,In_500,In_540);
nor U1944 (N_1944,In_136,In_692);
nand U1945 (N_1945,In_939,In_810);
and U1946 (N_1946,In_452,In_262);
nand U1947 (N_1947,In_515,In_613);
nand U1948 (N_1948,In_879,In_333);
nor U1949 (N_1949,In_298,In_425);
nor U1950 (N_1950,In_132,In_283);
and U1951 (N_1951,In_757,In_586);
nand U1952 (N_1952,In_862,In_421);
or U1953 (N_1953,In_859,In_332);
or U1954 (N_1954,In_234,In_14);
or U1955 (N_1955,In_232,In_217);
and U1956 (N_1956,In_444,In_122);
and U1957 (N_1957,In_144,In_919);
or U1958 (N_1958,In_139,In_364);
or U1959 (N_1959,In_478,In_873);
nand U1960 (N_1960,In_495,In_530);
nand U1961 (N_1961,In_830,In_627);
and U1962 (N_1962,In_991,In_175);
and U1963 (N_1963,In_738,In_163);
and U1964 (N_1964,In_788,In_71);
and U1965 (N_1965,In_486,In_345);
nor U1966 (N_1966,In_685,In_766);
or U1967 (N_1967,In_477,In_79);
or U1968 (N_1968,In_702,In_553);
nand U1969 (N_1969,In_478,In_568);
nor U1970 (N_1970,In_994,In_635);
or U1971 (N_1971,In_324,In_86);
xor U1972 (N_1972,In_861,In_250);
nor U1973 (N_1973,In_317,In_402);
or U1974 (N_1974,In_98,In_584);
and U1975 (N_1975,In_819,In_540);
nor U1976 (N_1976,In_356,In_66);
nand U1977 (N_1977,In_351,In_704);
and U1978 (N_1978,In_455,In_82);
and U1979 (N_1979,In_516,In_787);
xnor U1980 (N_1980,In_653,In_66);
or U1981 (N_1981,In_308,In_111);
and U1982 (N_1982,In_435,In_121);
and U1983 (N_1983,In_749,In_217);
nor U1984 (N_1984,In_740,In_560);
nor U1985 (N_1985,In_885,In_560);
or U1986 (N_1986,In_427,In_221);
and U1987 (N_1987,In_232,In_312);
or U1988 (N_1988,In_554,In_973);
nor U1989 (N_1989,In_139,In_929);
xnor U1990 (N_1990,In_769,In_67);
and U1991 (N_1991,In_357,In_875);
nand U1992 (N_1992,In_105,In_496);
or U1993 (N_1993,In_771,In_597);
nand U1994 (N_1994,In_287,In_721);
and U1995 (N_1995,In_660,In_592);
nand U1996 (N_1996,In_641,In_893);
nand U1997 (N_1997,In_548,In_80);
nand U1998 (N_1998,In_589,In_980);
or U1999 (N_1999,In_446,In_516);
nor U2000 (N_2000,In_480,In_773);
and U2001 (N_2001,In_885,In_645);
nor U2002 (N_2002,In_636,In_281);
or U2003 (N_2003,In_429,In_915);
nand U2004 (N_2004,In_784,In_146);
or U2005 (N_2005,In_26,In_254);
and U2006 (N_2006,In_286,In_34);
and U2007 (N_2007,In_655,In_402);
nand U2008 (N_2008,In_663,In_557);
and U2009 (N_2009,In_407,In_724);
nor U2010 (N_2010,In_161,In_995);
and U2011 (N_2011,In_683,In_714);
and U2012 (N_2012,In_814,In_146);
and U2013 (N_2013,In_733,In_363);
and U2014 (N_2014,In_196,In_933);
and U2015 (N_2015,In_812,In_501);
nor U2016 (N_2016,In_354,In_350);
and U2017 (N_2017,In_429,In_71);
nor U2018 (N_2018,In_199,In_787);
nor U2019 (N_2019,In_530,In_904);
or U2020 (N_2020,In_742,In_706);
nand U2021 (N_2021,In_527,In_140);
and U2022 (N_2022,In_280,In_726);
nand U2023 (N_2023,In_842,In_246);
and U2024 (N_2024,In_517,In_604);
and U2025 (N_2025,In_971,In_931);
nand U2026 (N_2026,In_168,In_763);
or U2027 (N_2027,In_927,In_793);
nand U2028 (N_2028,In_198,In_920);
nor U2029 (N_2029,In_494,In_761);
nand U2030 (N_2030,In_8,In_513);
nor U2031 (N_2031,In_538,In_79);
nand U2032 (N_2032,In_139,In_56);
or U2033 (N_2033,In_867,In_340);
xnor U2034 (N_2034,In_729,In_888);
nand U2035 (N_2035,In_320,In_184);
nand U2036 (N_2036,In_735,In_472);
and U2037 (N_2037,In_322,In_297);
or U2038 (N_2038,In_178,In_645);
nand U2039 (N_2039,In_406,In_501);
nand U2040 (N_2040,In_588,In_625);
and U2041 (N_2041,In_242,In_472);
or U2042 (N_2042,In_267,In_32);
nand U2043 (N_2043,In_284,In_367);
nor U2044 (N_2044,In_212,In_277);
nor U2045 (N_2045,In_47,In_625);
nand U2046 (N_2046,In_798,In_171);
or U2047 (N_2047,In_647,In_762);
nor U2048 (N_2048,In_913,In_784);
nor U2049 (N_2049,In_337,In_227);
nor U2050 (N_2050,In_87,In_497);
and U2051 (N_2051,In_730,In_988);
nor U2052 (N_2052,In_661,In_420);
nor U2053 (N_2053,In_435,In_658);
nor U2054 (N_2054,In_921,In_630);
and U2055 (N_2055,In_128,In_67);
nand U2056 (N_2056,In_907,In_810);
nand U2057 (N_2057,In_525,In_340);
nor U2058 (N_2058,In_893,In_484);
nor U2059 (N_2059,In_738,In_335);
and U2060 (N_2060,In_784,In_41);
or U2061 (N_2061,In_829,In_778);
or U2062 (N_2062,In_716,In_248);
and U2063 (N_2063,In_199,In_52);
nor U2064 (N_2064,In_264,In_698);
and U2065 (N_2065,In_794,In_156);
and U2066 (N_2066,In_971,In_733);
and U2067 (N_2067,In_19,In_865);
or U2068 (N_2068,In_817,In_475);
or U2069 (N_2069,In_676,In_731);
and U2070 (N_2070,In_904,In_99);
nor U2071 (N_2071,In_894,In_181);
nor U2072 (N_2072,In_362,In_827);
and U2073 (N_2073,In_170,In_78);
nand U2074 (N_2074,In_113,In_172);
nor U2075 (N_2075,In_895,In_846);
nand U2076 (N_2076,In_663,In_364);
and U2077 (N_2077,In_596,In_145);
nor U2078 (N_2078,In_204,In_86);
and U2079 (N_2079,In_892,In_22);
and U2080 (N_2080,In_232,In_31);
and U2081 (N_2081,In_5,In_998);
nor U2082 (N_2082,In_500,In_33);
nor U2083 (N_2083,In_250,In_880);
and U2084 (N_2084,In_241,In_874);
or U2085 (N_2085,In_315,In_491);
nor U2086 (N_2086,In_157,In_4);
nor U2087 (N_2087,In_974,In_265);
nand U2088 (N_2088,In_813,In_921);
and U2089 (N_2089,In_491,In_827);
or U2090 (N_2090,In_5,In_108);
or U2091 (N_2091,In_540,In_564);
and U2092 (N_2092,In_170,In_429);
nor U2093 (N_2093,In_61,In_367);
nand U2094 (N_2094,In_37,In_471);
nand U2095 (N_2095,In_544,In_412);
or U2096 (N_2096,In_465,In_857);
nand U2097 (N_2097,In_942,In_39);
nand U2098 (N_2098,In_311,In_429);
and U2099 (N_2099,In_521,In_517);
xnor U2100 (N_2100,In_499,In_519);
nor U2101 (N_2101,In_289,In_995);
or U2102 (N_2102,In_481,In_90);
nor U2103 (N_2103,In_835,In_621);
and U2104 (N_2104,In_121,In_654);
nand U2105 (N_2105,In_149,In_870);
nor U2106 (N_2106,In_999,In_691);
nor U2107 (N_2107,In_936,In_663);
and U2108 (N_2108,In_626,In_301);
or U2109 (N_2109,In_946,In_759);
or U2110 (N_2110,In_181,In_358);
and U2111 (N_2111,In_883,In_180);
or U2112 (N_2112,In_748,In_62);
nand U2113 (N_2113,In_663,In_529);
and U2114 (N_2114,In_803,In_863);
nand U2115 (N_2115,In_622,In_193);
or U2116 (N_2116,In_187,In_613);
and U2117 (N_2117,In_979,In_417);
nand U2118 (N_2118,In_992,In_227);
nand U2119 (N_2119,In_870,In_437);
or U2120 (N_2120,In_210,In_701);
and U2121 (N_2121,In_589,In_2);
nor U2122 (N_2122,In_753,In_773);
nor U2123 (N_2123,In_367,In_790);
nand U2124 (N_2124,In_988,In_737);
and U2125 (N_2125,In_585,In_645);
and U2126 (N_2126,In_824,In_634);
nor U2127 (N_2127,In_794,In_287);
or U2128 (N_2128,In_945,In_230);
and U2129 (N_2129,In_947,In_994);
nand U2130 (N_2130,In_100,In_275);
and U2131 (N_2131,In_289,In_277);
or U2132 (N_2132,In_967,In_33);
nand U2133 (N_2133,In_453,In_580);
and U2134 (N_2134,In_461,In_599);
nor U2135 (N_2135,In_461,In_477);
or U2136 (N_2136,In_685,In_936);
nor U2137 (N_2137,In_190,In_807);
nor U2138 (N_2138,In_874,In_736);
or U2139 (N_2139,In_236,In_541);
or U2140 (N_2140,In_254,In_880);
nor U2141 (N_2141,In_110,In_656);
or U2142 (N_2142,In_361,In_962);
and U2143 (N_2143,In_243,In_652);
nand U2144 (N_2144,In_10,In_92);
and U2145 (N_2145,In_436,In_904);
nor U2146 (N_2146,In_264,In_281);
or U2147 (N_2147,In_616,In_296);
and U2148 (N_2148,In_293,In_573);
nand U2149 (N_2149,In_230,In_598);
or U2150 (N_2150,In_478,In_382);
and U2151 (N_2151,In_581,In_442);
or U2152 (N_2152,In_219,In_117);
nand U2153 (N_2153,In_701,In_806);
and U2154 (N_2154,In_662,In_439);
xnor U2155 (N_2155,In_298,In_581);
or U2156 (N_2156,In_802,In_732);
or U2157 (N_2157,In_507,In_926);
or U2158 (N_2158,In_766,In_861);
nand U2159 (N_2159,In_471,In_927);
and U2160 (N_2160,In_957,In_635);
and U2161 (N_2161,In_445,In_678);
nand U2162 (N_2162,In_735,In_299);
nor U2163 (N_2163,In_480,In_12);
nor U2164 (N_2164,In_406,In_261);
nor U2165 (N_2165,In_307,In_348);
nor U2166 (N_2166,In_799,In_674);
nor U2167 (N_2167,In_763,In_675);
nand U2168 (N_2168,In_666,In_668);
and U2169 (N_2169,In_946,In_825);
nand U2170 (N_2170,In_842,In_875);
and U2171 (N_2171,In_754,In_950);
and U2172 (N_2172,In_312,In_885);
and U2173 (N_2173,In_215,In_843);
and U2174 (N_2174,In_676,In_385);
or U2175 (N_2175,In_493,In_320);
nor U2176 (N_2176,In_309,In_586);
nand U2177 (N_2177,In_380,In_532);
nand U2178 (N_2178,In_342,In_285);
nor U2179 (N_2179,In_519,In_661);
nor U2180 (N_2180,In_93,In_90);
nand U2181 (N_2181,In_935,In_805);
nor U2182 (N_2182,In_34,In_515);
nand U2183 (N_2183,In_739,In_198);
nor U2184 (N_2184,In_142,In_987);
or U2185 (N_2185,In_798,In_395);
nand U2186 (N_2186,In_247,In_475);
nand U2187 (N_2187,In_19,In_352);
xnor U2188 (N_2188,In_1,In_303);
nor U2189 (N_2189,In_122,In_538);
nand U2190 (N_2190,In_755,In_710);
nor U2191 (N_2191,In_542,In_128);
nand U2192 (N_2192,In_587,In_425);
nor U2193 (N_2193,In_974,In_283);
and U2194 (N_2194,In_512,In_200);
and U2195 (N_2195,In_459,In_487);
nor U2196 (N_2196,In_567,In_663);
or U2197 (N_2197,In_321,In_45);
nor U2198 (N_2198,In_484,In_423);
nand U2199 (N_2199,In_524,In_748);
or U2200 (N_2200,In_741,In_522);
and U2201 (N_2201,In_868,In_418);
and U2202 (N_2202,In_176,In_150);
or U2203 (N_2203,In_534,In_955);
and U2204 (N_2204,In_725,In_842);
xor U2205 (N_2205,In_620,In_664);
nor U2206 (N_2206,In_880,In_391);
nand U2207 (N_2207,In_987,In_931);
and U2208 (N_2208,In_901,In_124);
nand U2209 (N_2209,In_816,In_150);
and U2210 (N_2210,In_587,In_524);
or U2211 (N_2211,In_231,In_149);
nor U2212 (N_2212,In_648,In_350);
nand U2213 (N_2213,In_772,In_905);
or U2214 (N_2214,In_34,In_709);
nand U2215 (N_2215,In_496,In_452);
or U2216 (N_2216,In_540,In_61);
nand U2217 (N_2217,In_148,In_799);
nor U2218 (N_2218,In_411,In_70);
nand U2219 (N_2219,In_735,In_352);
nand U2220 (N_2220,In_833,In_704);
nor U2221 (N_2221,In_228,In_239);
or U2222 (N_2222,In_157,In_757);
and U2223 (N_2223,In_63,In_400);
nand U2224 (N_2224,In_83,In_63);
nand U2225 (N_2225,In_779,In_426);
or U2226 (N_2226,In_654,In_136);
and U2227 (N_2227,In_762,In_914);
and U2228 (N_2228,In_990,In_419);
and U2229 (N_2229,In_173,In_412);
or U2230 (N_2230,In_553,In_661);
and U2231 (N_2231,In_935,In_86);
nor U2232 (N_2232,In_995,In_630);
or U2233 (N_2233,In_39,In_485);
and U2234 (N_2234,In_553,In_378);
nor U2235 (N_2235,In_47,In_593);
or U2236 (N_2236,In_40,In_971);
and U2237 (N_2237,In_654,In_631);
and U2238 (N_2238,In_802,In_544);
and U2239 (N_2239,In_553,In_863);
nor U2240 (N_2240,In_972,In_783);
nor U2241 (N_2241,In_188,In_304);
nand U2242 (N_2242,In_957,In_582);
and U2243 (N_2243,In_301,In_438);
and U2244 (N_2244,In_695,In_383);
nand U2245 (N_2245,In_772,In_86);
nor U2246 (N_2246,In_318,In_965);
or U2247 (N_2247,In_429,In_58);
or U2248 (N_2248,In_868,In_343);
nor U2249 (N_2249,In_923,In_344);
nand U2250 (N_2250,In_683,In_875);
nand U2251 (N_2251,In_528,In_20);
or U2252 (N_2252,In_220,In_549);
xnor U2253 (N_2253,In_907,In_927);
nand U2254 (N_2254,In_188,In_483);
or U2255 (N_2255,In_789,In_709);
nand U2256 (N_2256,In_404,In_933);
or U2257 (N_2257,In_301,In_561);
nand U2258 (N_2258,In_876,In_874);
or U2259 (N_2259,In_597,In_278);
nor U2260 (N_2260,In_191,In_30);
nand U2261 (N_2261,In_418,In_976);
nand U2262 (N_2262,In_432,In_37);
nand U2263 (N_2263,In_167,In_296);
nand U2264 (N_2264,In_104,In_592);
nor U2265 (N_2265,In_272,In_518);
and U2266 (N_2266,In_784,In_527);
or U2267 (N_2267,In_856,In_820);
nor U2268 (N_2268,In_341,In_829);
nand U2269 (N_2269,In_569,In_943);
nor U2270 (N_2270,In_206,In_719);
or U2271 (N_2271,In_401,In_208);
and U2272 (N_2272,In_533,In_484);
and U2273 (N_2273,In_666,In_846);
nand U2274 (N_2274,In_323,In_344);
or U2275 (N_2275,In_166,In_25);
nor U2276 (N_2276,In_799,In_739);
and U2277 (N_2277,In_204,In_536);
and U2278 (N_2278,In_157,In_971);
nor U2279 (N_2279,In_520,In_896);
nor U2280 (N_2280,In_389,In_762);
nor U2281 (N_2281,In_65,In_527);
nor U2282 (N_2282,In_546,In_898);
nand U2283 (N_2283,In_449,In_162);
nor U2284 (N_2284,In_725,In_586);
nand U2285 (N_2285,In_965,In_565);
or U2286 (N_2286,In_871,In_869);
and U2287 (N_2287,In_982,In_222);
nand U2288 (N_2288,In_325,In_612);
or U2289 (N_2289,In_44,In_791);
nand U2290 (N_2290,In_11,In_862);
or U2291 (N_2291,In_277,In_288);
nand U2292 (N_2292,In_863,In_759);
nand U2293 (N_2293,In_255,In_385);
nor U2294 (N_2294,In_679,In_951);
nor U2295 (N_2295,In_986,In_738);
nand U2296 (N_2296,In_429,In_303);
nor U2297 (N_2297,In_742,In_445);
or U2298 (N_2298,In_144,In_507);
nand U2299 (N_2299,In_300,In_14);
and U2300 (N_2300,In_105,In_202);
or U2301 (N_2301,In_500,In_274);
nand U2302 (N_2302,In_804,In_284);
or U2303 (N_2303,In_705,In_376);
or U2304 (N_2304,In_697,In_380);
or U2305 (N_2305,In_150,In_342);
or U2306 (N_2306,In_184,In_958);
nor U2307 (N_2307,In_64,In_940);
and U2308 (N_2308,In_480,In_312);
nand U2309 (N_2309,In_365,In_116);
or U2310 (N_2310,In_677,In_125);
or U2311 (N_2311,In_182,In_999);
and U2312 (N_2312,In_553,In_42);
nor U2313 (N_2313,In_705,In_728);
and U2314 (N_2314,In_30,In_153);
nand U2315 (N_2315,In_370,In_535);
nand U2316 (N_2316,In_356,In_116);
xnor U2317 (N_2317,In_902,In_743);
nor U2318 (N_2318,In_418,In_913);
xnor U2319 (N_2319,In_208,In_514);
nor U2320 (N_2320,In_106,In_69);
and U2321 (N_2321,In_408,In_741);
and U2322 (N_2322,In_843,In_51);
and U2323 (N_2323,In_386,In_684);
nand U2324 (N_2324,In_401,In_655);
nand U2325 (N_2325,In_196,In_932);
xor U2326 (N_2326,In_743,In_700);
or U2327 (N_2327,In_821,In_99);
or U2328 (N_2328,In_73,In_627);
and U2329 (N_2329,In_356,In_395);
and U2330 (N_2330,In_319,In_158);
nand U2331 (N_2331,In_297,In_33);
nand U2332 (N_2332,In_113,In_52);
and U2333 (N_2333,In_897,In_121);
nand U2334 (N_2334,In_823,In_517);
and U2335 (N_2335,In_297,In_204);
or U2336 (N_2336,In_255,In_100);
or U2337 (N_2337,In_592,In_74);
nor U2338 (N_2338,In_335,In_330);
nor U2339 (N_2339,In_78,In_656);
nor U2340 (N_2340,In_33,In_68);
nand U2341 (N_2341,In_207,In_412);
nor U2342 (N_2342,In_203,In_338);
and U2343 (N_2343,In_315,In_530);
nor U2344 (N_2344,In_788,In_86);
nand U2345 (N_2345,In_574,In_928);
and U2346 (N_2346,In_750,In_956);
or U2347 (N_2347,In_13,In_335);
or U2348 (N_2348,In_104,In_753);
nand U2349 (N_2349,In_945,In_294);
or U2350 (N_2350,In_545,In_901);
nor U2351 (N_2351,In_84,In_564);
nor U2352 (N_2352,In_918,In_24);
and U2353 (N_2353,In_398,In_709);
or U2354 (N_2354,In_62,In_642);
or U2355 (N_2355,In_1,In_415);
xor U2356 (N_2356,In_315,In_381);
and U2357 (N_2357,In_3,In_494);
nand U2358 (N_2358,In_699,In_732);
or U2359 (N_2359,In_889,In_758);
nor U2360 (N_2360,In_57,In_126);
or U2361 (N_2361,In_256,In_480);
or U2362 (N_2362,In_636,In_140);
nor U2363 (N_2363,In_932,In_254);
nand U2364 (N_2364,In_160,In_463);
nand U2365 (N_2365,In_673,In_81);
nand U2366 (N_2366,In_471,In_10);
nor U2367 (N_2367,In_683,In_8);
and U2368 (N_2368,In_632,In_333);
and U2369 (N_2369,In_783,In_622);
nor U2370 (N_2370,In_398,In_499);
or U2371 (N_2371,In_742,In_19);
or U2372 (N_2372,In_429,In_787);
and U2373 (N_2373,In_102,In_785);
and U2374 (N_2374,In_268,In_671);
and U2375 (N_2375,In_28,In_51);
nor U2376 (N_2376,In_337,In_29);
nor U2377 (N_2377,In_923,In_717);
nand U2378 (N_2378,In_199,In_35);
and U2379 (N_2379,In_120,In_639);
nand U2380 (N_2380,In_831,In_737);
nor U2381 (N_2381,In_531,In_99);
and U2382 (N_2382,In_276,In_803);
or U2383 (N_2383,In_433,In_774);
and U2384 (N_2384,In_895,In_130);
nand U2385 (N_2385,In_521,In_202);
nor U2386 (N_2386,In_667,In_621);
or U2387 (N_2387,In_318,In_220);
nor U2388 (N_2388,In_850,In_140);
or U2389 (N_2389,In_105,In_457);
nand U2390 (N_2390,In_174,In_439);
or U2391 (N_2391,In_196,In_515);
nor U2392 (N_2392,In_280,In_718);
or U2393 (N_2393,In_623,In_921);
nand U2394 (N_2394,In_157,In_462);
or U2395 (N_2395,In_840,In_940);
nand U2396 (N_2396,In_229,In_439);
and U2397 (N_2397,In_18,In_578);
and U2398 (N_2398,In_589,In_100);
or U2399 (N_2399,In_301,In_597);
nor U2400 (N_2400,In_825,In_344);
nand U2401 (N_2401,In_870,In_298);
nand U2402 (N_2402,In_409,In_280);
nand U2403 (N_2403,In_92,In_777);
nor U2404 (N_2404,In_735,In_976);
nor U2405 (N_2405,In_333,In_515);
nor U2406 (N_2406,In_489,In_496);
and U2407 (N_2407,In_411,In_569);
and U2408 (N_2408,In_342,In_0);
nor U2409 (N_2409,In_135,In_137);
or U2410 (N_2410,In_5,In_299);
and U2411 (N_2411,In_916,In_207);
nand U2412 (N_2412,In_243,In_356);
or U2413 (N_2413,In_127,In_702);
nor U2414 (N_2414,In_215,In_220);
nor U2415 (N_2415,In_560,In_204);
nand U2416 (N_2416,In_474,In_822);
nand U2417 (N_2417,In_957,In_396);
and U2418 (N_2418,In_242,In_684);
and U2419 (N_2419,In_382,In_383);
or U2420 (N_2420,In_219,In_53);
and U2421 (N_2421,In_434,In_207);
or U2422 (N_2422,In_151,In_329);
nand U2423 (N_2423,In_410,In_148);
nor U2424 (N_2424,In_566,In_649);
and U2425 (N_2425,In_371,In_887);
nand U2426 (N_2426,In_386,In_282);
nor U2427 (N_2427,In_918,In_121);
nor U2428 (N_2428,In_666,In_665);
or U2429 (N_2429,In_765,In_642);
or U2430 (N_2430,In_844,In_359);
nand U2431 (N_2431,In_177,In_473);
or U2432 (N_2432,In_880,In_828);
nor U2433 (N_2433,In_557,In_524);
or U2434 (N_2434,In_414,In_193);
or U2435 (N_2435,In_14,In_647);
and U2436 (N_2436,In_927,In_418);
nand U2437 (N_2437,In_273,In_364);
nand U2438 (N_2438,In_739,In_211);
nand U2439 (N_2439,In_621,In_850);
nand U2440 (N_2440,In_334,In_437);
and U2441 (N_2441,In_936,In_370);
and U2442 (N_2442,In_706,In_793);
nor U2443 (N_2443,In_75,In_672);
or U2444 (N_2444,In_598,In_990);
nor U2445 (N_2445,In_803,In_151);
nand U2446 (N_2446,In_870,In_104);
nand U2447 (N_2447,In_218,In_986);
nor U2448 (N_2448,In_90,In_66);
or U2449 (N_2449,In_880,In_274);
or U2450 (N_2450,In_170,In_238);
nand U2451 (N_2451,In_34,In_196);
nor U2452 (N_2452,In_507,In_216);
or U2453 (N_2453,In_455,In_255);
or U2454 (N_2454,In_711,In_22);
or U2455 (N_2455,In_706,In_630);
or U2456 (N_2456,In_711,In_887);
nand U2457 (N_2457,In_184,In_539);
nand U2458 (N_2458,In_816,In_797);
xor U2459 (N_2459,In_222,In_376);
or U2460 (N_2460,In_424,In_620);
and U2461 (N_2461,In_403,In_36);
and U2462 (N_2462,In_100,In_763);
or U2463 (N_2463,In_452,In_141);
nor U2464 (N_2464,In_677,In_464);
or U2465 (N_2465,In_949,In_28);
or U2466 (N_2466,In_850,In_22);
and U2467 (N_2467,In_172,In_93);
or U2468 (N_2468,In_863,In_120);
or U2469 (N_2469,In_43,In_353);
nor U2470 (N_2470,In_572,In_372);
nor U2471 (N_2471,In_538,In_972);
nand U2472 (N_2472,In_178,In_213);
and U2473 (N_2473,In_633,In_877);
nor U2474 (N_2474,In_52,In_969);
or U2475 (N_2475,In_443,In_390);
nand U2476 (N_2476,In_698,In_424);
nand U2477 (N_2477,In_898,In_179);
and U2478 (N_2478,In_990,In_700);
and U2479 (N_2479,In_383,In_952);
or U2480 (N_2480,In_72,In_508);
nand U2481 (N_2481,In_55,In_341);
or U2482 (N_2482,In_716,In_288);
nand U2483 (N_2483,In_352,In_827);
nand U2484 (N_2484,In_543,In_932);
nand U2485 (N_2485,In_673,In_144);
and U2486 (N_2486,In_813,In_28);
and U2487 (N_2487,In_188,In_872);
nor U2488 (N_2488,In_588,In_924);
or U2489 (N_2489,In_764,In_470);
or U2490 (N_2490,In_953,In_456);
nor U2491 (N_2491,In_653,In_763);
nor U2492 (N_2492,In_9,In_633);
nor U2493 (N_2493,In_286,In_98);
or U2494 (N_2494,In_201,In_699);
and U2495 (N_2495,In_656,In_152);
nand U2496 (N_2496,In_165,In_503);
or U2497 (N_2497,In_386,In_616);
and U2498 (N_2498,In_952,In_303);
nor U2499 (N_2499,In_594,In_105);
or U2500 (N_2500,N_222,N_590);
and U2501 (N_2501,N_1474,N_1238);
and U2502 (N_2502,N_640,N_1586);
and U2503 (N_2503,N_1200,N_603);
nor U2504 (N_2504,N_455,N_1723);
nand U2505 (N_2505,N_1625,N_1385);
nor U2506 (N_2506,N_2317,N_1124);
or U2507 (N_2507,N_279,N_1937);
nand U2508 (N_2508,N_1577,N_1189);
or U2509 (N_2509,N_1001,N_1165);
or U2510 (N_2510,N_983,N_1966);
or U2511 (N_2511,N_732,N_2413);
nor U2512 (N_2512,N_1650,N_522);
or U2513 (N_2513,N_1348,N_1674);
and U2514 (N_2514,N_1830,N_562);
nand U2515 (N_2515,N_2145,N_2342);
nand U2516 (N_2516,N_1147,N_1459);
or U2517 (N_2517,N_234,N_1125);
and U2518 (N_2518,N_333,N_57);
or U2519 (N_2519,N_1065,N_399);
and U2520 (N_2520,N_1801,N_193);
nor U2521 (N_2521,N_2036,N_1686);
nor U2522 (N_2522,N_1356,N_2440);
and U2523 (N_2523,N_489,N_2439);
or U2524 (N_2524,N_1386,N_491);
or U2525 (N_2525,N_220,N_751);
or U2526 (N_2526,N_2048,N_1048);
and U2527 (N_2527,N_1950,N_1063);
nand U2528 (N_2528,N_864,N_366);
or U2529 (N_2529,N_1691,N_898);
nand U2530 (N_2530,N_114,N_1246);
nor U2531 (N_2531,N_1593,N_1953);
nand U2532 (N_2532,N_340,N_1399);
nand U2533 (N_2533,N_919,N_750);
or U2534 (N_2534,N_1151,N_2015);
and U2535 (N_2535,N_685,N_1914);
or U2536 (N_2536,N_192,N_1865);
or U2537 (N_2537,N_253,N_111);
and U2538 (N_2538,N_109,N_2302);
nor U2539 (N_2539,N_1143,N_2034);
and U2540 (N_2540,N_1102,N_2318);
and U2541 (N_2541,N_2049,N_200);
nand U2542 (N_2542,N_1305,N_1807);
or U2543 (N_2543,N_1741,N_1491);
nor U2544 (N_2544,N_1560,N_1714);
nand U2545 (N_2545,N_2406,N_1843);
nand U2546 (N_2546,N_1133,N_1106);
and U2547 (N_2547,N_370,N_226);
and U2548 (N_2548,N_1044,N_332);
nand U2549 (N_2549,N_1027,N_2364);
nor U2550 (N_2550,N_866,N_1997);
nand U2551 (N_2551,N_997,N_1020);
nand U2552 (N_2552,N_2299,N_1996);
and U2553 (N_2553,N_1419,N_1547);
nand U2554 (N_2554,N_257,N_807);
nor U2555 (N_2555,N_8,N_369);
and U2556 (N_2556,N_81,N_1268);
nor U2557 (N_2557,N_1538,N_1878);
nand U2558 (N_2558,N_209,N_2156);
and U2559 (N_2559,N_1852,N_238);
and U2560 (N_2560,N_2350,N_2155);
and U2561 (N_2561,N_352,N_819);
nor U2562 (N_2562,N_47,N_1248);
or U2563 (N_2563,N_1828,N_844);
or U2564 (N_2564,N_1884,N_1234);
nand U2565 (N_2565,N_2188,N_1235);
and U2566 (N_2566,N_1363,N_1528);
or U2567 (N_2567,N_2196,N_1928);
nand U2568 (N_2568,N_1506,N_523);
nor U2569 (N_2569,N_1543,N_2149);
nand U2570 (N_2570,N_2136,N_947);
or U2571 (N_2571,N_882,N_2495);
nor U2572 (N_2572,N_872,N_1082);
and U2573 (N_2573,N_1122,N_1226);
nor U2574 (N_2574,N_722,N_1427);
or U2575 (N_2575,N_258,N_555);
xnor U2576 (N_2576,N_1026,N_1249);
or U2577 (N_2577,N_1934,N_2425);
or U2578 (N_2578,N_867,N_85);
or U2579 (N_2579,N_1738,N_2434);
or U2580 (N_2580,N_402,N_275);
nand U2581 (N_2581,N_297,N_422);
and U2582 (N_2582,N_829,N_156);
nor U2583 (N_2583,N_1636,N_1777);
nand U2584 (N_2584,N_296,N_1021);
and U2585 (N_2585,N_2488,N_1033);
and U2586 (N_2586,N_1605,N_1278);
or U2587 (N_2587,N_487,N_1339);
nor U2588 (N_2588,N_2479,N_2189);
nand U2589 (N_2589,N_1508,N_2327);
nor U2590 (N_2590,N_2007,N_182);
or U2591 (N_2591,N_1324,N_535);
nor U2592 (N_2592,N_361,N_1939);
nor U2593 (N_2593,N_1377,N_641);
and U2594 (N_2594,N_34,N_716);
or U2595 (N_2595,N_1052,N_2073);
nor U2596 (N_2596,N_683,N_1397);
and U2597 (N_2597,N_2480,N_1757);
nand U2598 (N_2598,N_2276,N_1150);
or U2599 (N_2599,N_703,N_926);
or U2600 (N_2600,N_2431,N_534);
or U2601 (N_2601,N_1263,N_2260);
and U2602 (N_2602,N_1909,N_2108);
nand U2603 (N_2603,N_2450,N_1564);
or U2604 (N_2604,N_164,N_2494);
xor U2605 (N_2605,N_118,N_654);
and U2606 (N_2606,N_2037,N_2058);
or U2607 (N_2607,N_1436,N_981);
nand U2608 (N_2608,N_2198,N_1756);
or U2609 (N_2609,N_1510,N_1005);
or U2610 (N_2610,N_2152,N_319);
or U2611 (N_2611,N_1227,N_736);
xor U2612 (N_2612,N_419,N_1628);
or U2613 (N_2613,N_500,N_550);
nand U2614 (N_2614,N_1706,N_848);
nand U2615 (N_2615,N_908,N_2308);
nand U2616 (N_2616,N_2498,N_1479);
and U2617 (N_2617,N_175,N_1047);
or U2618 (N_2618,N_108,N_2201);
or U2619 (N_2619,N_2119,N_836);
or U2620 (N_2620,N_2124,N_762);
or U2621 (N_2621,N_2477,N_1844);
or U2622 (N_2622,N_1374,N_364);
or U2623 (N_2623,N_909,N_1958);
and U2624 (N_2624,N_1011,N_2447);
or U2625 (N_2625,N_2235,N_1494);
nand U2626 (N_2626,N_987,N_138);
nand U2627 (N_2627,N_1,N_350);
nor U2628 (N_2628,N_540,N_1434);
or U2629 (N_2629,N_1632,N_2286);
nand U2630 (N_2630,N_468,N_1907);
nand U2631 (N_2631,N_1422,N_430);
or U2632 (N_2632,N_502,N_771);
and U2633 (N_2633,N_1781,N_608);
nor U2634 (N_2634,N_1276,N_755);
and U2635 (N_2635,N_1432,N_2024);
and U2636 (N_2636,N_1464,N_276);
and U2637 (N_2637,N_1025,N_2292);
xnor U2638 (N_2638,N_865,N_1619);
nor U2639 (N_2639,N_835,N_407);
and U2640 (N_2640,N_244,N_1693);
or U2641 (N_2641,N_881,N_224);
nand U2642 (N_2642,N_2236,N_2252);
nand U2643 (N_2643,N_1612,N_1530);
nor U2644 (N_2644,N_1765,N_679);
nand U2645 (N_2645,N_1213,N_1664);
nand U2646 (N_2646,N_1130,N_971);
or U2647 (N_2647,N_2421,N_2291);
and U2648 (N_2648,N_2100,N_1059);
nand U2649 (N_2649,N_1146,N_273);
or U2650 (N_2650,N_2315,N_1710);
nand U2651 (N_2651,N_519,N_571);
nand U2652 (N_2652,N_1840,N_826);
and U2653 (N_2653,N_1300,N_2064);
nor U2654 (N_2654,N_39,N_1887);
or U2655 (N_2655,N_1794,N_928);
and U2656 (N_2656,N_239,N_1223);
nor U2657 (N_2657,N_1793,N_1416);
nor U2658 (N_2658,N_2401,N_996);
and U2659 (N_2659,N_301,N_870);
and U2660 (N_2660,N_1288,N_2052);
or U2661 (N_2661,N_1333,N_1180);
and U2662 (N_2662,N_681,N_1393);
nor U2663 (N_2663,N_1250,N_643);
or U2664 (N_2664,N_428,N_1796);
or U2665 (N_2665,N_2251,N_989);
or U2666 (N_2666,N_1314,N_936);
xnor U2667 (N_2667,N_2000,N_2436);
nor U2668 (N_2668,N_46,N_871);
nand U2669 (N_2669,N_1616,N_1751);
nor U2670 (N_2670,N_2372,N_1834);
nor U2671 (N_2671,N_1228,N_1407);
nor U2672 (N_2672,N_2078,N_1798);
nand U2673 (N_2673,N_1384,N_783);
and U2674 (N_2674,N_126,N_934);
nand U2675 (N_2675,N_259,N_2255);
nand U2676 (N_2676,N_1800,N_1214);
and U2677 (N_2677,N_1215,N_125);
nand U2678 (N_2678,N_1946,N_0);
xor U2679 (N_2679,N_1572,N_1003);
nand U2680 (N_2680,N_568,N_1309);
nand U2681 (N_2681,N_195,N_642);
nor U2682 (N_2682,N_1673,N_174);
or U2683 (N_2683,N_1495,N_915);
or U2684 (N_2684,N_3,N_665);
or U2685 (N_2685,N_1008,N_1343);
nand U2686 (N_2686,N_1992,N_1209);
nand U2687 (N_2687,N_1835,N_2388);
or U2688 (N_2688,N_704,N_597);
and U2689 (N_2689,N_1929,N_1651);
nor U2690 (N_2690,N_899,N_1949);
nor U2691 (N_2691,N_2120,N_1489);
nand U2692 (N_2692,N_561,N_1947);
and U2693 (N_2693,N_1859,N_2381);
nor U2694 (N_2694,N_151,N_2424);
nand U2695 (N_2695,N_1039,N_2496);
or U2696 (N_2696,N_1444,N_2127);
xnor U2697 (N_2697,N_1196,N_1264);
nor U2698 (N_2698,N_2219,N_2343);
or U2699 (N_2699,N_2375,N_1119);
nor U2700 (N_2700,N_1590,N_905);
and U2701 (N_2701,N_1131,N_2194);
and U2702 (N_2702,N_1601,N_787);
and U2703 (N_2703,N_1372,N_2077);
and U2704 (N_2704,N_1221,N_408);
or U2705 (N_2705,N_767,N_2275);
or U2706 (N_2706,N_1408,N_1321);
nor U2707 (N_2707,N_710,N_651);
nor U2708 (N_2708,N_991,N_1822);
or U2709 (N_2709,N_1779,N_932);
nor U2710 (N_2710,N_2316,N_1135);
or U2711 (N_2711,N_1607,N_820);
nand U2712 (N_2712,N_1812,N_358);
xor U2713 (N_2713,N_498,N_2337);
nor U2714 (N_2714,N_1144,N_1054);
nand U2715 (N_2715,N_717,N_2366);
xnor U2716 (N_2716,N_860,N_1977);
or U2717 (N_2717,N_1987,N_2497);
nand U2718 (N_2718,N_1160,N_1608);
and U2719 (N_2719,N_62,N_122);
and U2720 (N_2720,N_417,N_442);
nor U2721 (N_2721,N_1940,N_2322);
xor U2722 (N_2722,N_1944,N_1123);
nor U2723 (N_2723,N_60,N_621);
nand U2724 (N_2724,N_558,N_1905);
and U2725 (N_2725,N_1661,N_1916);
and U2726 (N_2726,N_1207,N_749);
and U2727 (N_2727,N_1967,N_91);
and U2728 (N_2728,N_2191,N_2033);
xor U2729 (N_2729,N_2386,N_1322);
or U2730 (N_2730,N_1079,N_270);
or U2731 (N_2731,N_413,N_344);
nand U2732 (N_2732,N_1867,N_392);
nand U2733 (N_2733,N_2223,N_1938);
and U2734 (N_2734,N_676,N_520);
nor U2735 (N_2735,N_956,N_12);
nor U2736 (N_2736,N_1960,N_566);
or U2737 (N_2737,N_400,N_1795);
and U2738 (N_2738,N_2269,N_1814);
xor U2739 (N_2739,N_2489,N_559);
nand U2740 (N_2740,N_17,N_1519);
and U2741 (N_2741,N_1137,N_287);
or U2742 (N_2742,N_1568,N_890);
or U2743 (N_2743,N_492,N_1641);
nor U2744 (N_2744,N_1627,N_1925);
and U2745 (N_2745,N_1174,N_1876);
nand U2746 (N_2746,N_201,N_2396);
nand U2747 (N_2747,N_2471,N_38);
nor U2748 (N_2748,N_499,N_2047);
or U2749 (N_2749,N_2218,N_1555);
or U2750 (N_2750,N_1291,N_1403);
or U2751 (N_2751,N_1889,N_2279);
xnor U2752 (N_2752,N_474,N_678);
nand U2753 (N_2753,N_178,N_980);
or U2754 (N_2754,N_1525,N_2206);
nand U2755 (N_2755,N_2378,N_2228);
nor U2756 (N_2756,N_1646,N_397);
and U2757 (N_2757,N_1297,N_1846);
or U2758 (N_2758,N_2423,N_1883);
or U2759 (N_2759,N_354,N_2070);
and U2760 (N_2760,N_446,N_1428);
nor U2761 (N_2761,N_1791,N_1563);
nand U2762 (N_2762,N_1580,N_2069);
nand U2763 (N_2763,N_1556,N_792);
nand U2764 (N_2764,N_2377,N_1552);
and U2765 (N_2765,N_1164,N_129);
nor U2766 (N_2766,N_806,N_803);
nor U2767 (N_2767,N_2143,N_204);
nand U2768 (N_2768,N_373,N_2487);
nand U2769 (N_2769,N_1284,N_1856);
nand U2770 (N_2770,N_2159,N_271);
nand U2771 (N_2771,N_548,N_1549);
nor U2772 (N_2772,N_1265,N_1128);
nand U2773 (N_2773,N_1837,N_1262);
or U2774 (N_2774,N_155,N_1327);
or U2775 (N_2775,N_496,N_180);
or U2776 (N_2776,N_218,N_2084);
or U2777 (N_2777,N_472,N_1923);
and U2778 (N_2778,N_158,N_35);
nand U2779 (N_2779,N_1936,N_99);
nor U2780 (N_2780,N_1985,N_2131);
nor U2781 (N_2781,N_1685,N_2474);
nand U2782 (N_2782,N_1726,N_395);
or U2783 (N_2783,N_1388,N_900);
nor U2784 (N_2784,N_1755,N_1753);
nor U2785 (N_2785,N_1918,N_849);
nor U2786 (N_2786,N_1329,N_733);
or U2787 (N_2787,N_1711,N_846);
and U2788 (N_2788,N_1991,N_1171);
and U2789 (N_2789,N_360,N_2349);
nor U2790 (N_2790,N_1702,N_1378);
nor U2791 (N_2791,N_2059,N_2259);
nand U2792 (N_2792,N_2150,N_1177);
and U2793 (N_2793,N_847,N_2180);
nor U2794 (N_2794,N_1340,N_2226);
xor U2795 (N_2795,N_2261,N_453);
nor U2796 (N_2796,N_2466,N_2281);
nor U2797 (N_2797,N_2250,N_675);
or U2798 (N_2798,N_1570,N_368);
or U2799 (N_2799,N_2408,N_1247);
or U2800 (N_2800,N_2167,N_2465);
nand U2801 (N_2801,N_282,N_1776);
nor U2802 (N_2802,N_521,N_2455);
nand U2803 (N_2803,N_1290,N_670);
and U2804 (N_2804,N_2220,N_691);
nor U2805 (N_2805,N_44,N_1720);
or U2806 (N_2806,N_1462,N_1891);
or U2807 (N_2807,N_1855,N_177);
or U2808 (N_2808,N_878,N_1129);
or U2809 (N_2809,N_127,N_2039);
and U2810 (N_2810,N_172,N_1470);
nand U2811 (N_2811,N_1527,N_313);
nor U2812 (N_2812,N_891,N_2384);
nand U2813 (N_2813,N_595,N_702);
nor U2814 (N_2814,N_1999,N_362);
and U2815 (N_2815,N_584,N_2444);
nand U2816 (N_2816,N_481,N_761);
nor U2817 (N_2817,N_874,N_371);
nand U2818 (N_2818,N_2456,N_144);
and U2819 (N_2819,N_1225,N_1473);
nor U2820 (N_2820,N_977,N_1698);
nand U2821 (N_2821,N_1239,N_459);
nand U2822 (N_2822,N_1456,N_1965);
nand U2823 (N_2823,N_1198,N_329);
nor U2824 (N_2824,N_470,N_563);
or U2825 (N_2825,N_1860,N_1551);
nand U2826 (N_2826,N_1353,N_930);
and U2827 (N_2827,N_1542,N_1638);
nand U2828 (N_2828,N_1733,N_2391);
and U2829 (N_2829,N_1310,N_1058);
or U2830 (N_2830,N_1886,N_758);
nor U2831 (N_2831,N_490,N_677);
nand U2832 (N_2832,N_1347,N_1790);
and U2833 (N_2833,N_213,N_944);
and U2834 (N_2834,N_901,N_2050);
nand U2835 (N_2835,N_1104,N_1271);
nor U2836 (N_2836,N_1145,N_1617);
nor U2837 (N_2837,N_1841,N_950);
nor U2838 (N_2838,N_73,N_179);
nand U2839 (N_2839,N_1451,N_2134);
nand U2840 (N_2840,N_495,N_1424);
and U2841 (N_2841,N_1369,N_1357);
and U2842 (N_2842,N_1645,N_1443);
nand U2843 (N_2843,N_1064,N_2485);
and U2844 (N_2844,N_576,N_377);
nor U2845 (N_2845,N_1758,N_634);
nand U2846 (N_2846,N_2435,N_589);
and U2847 (N_2847,N_1526,N_345);
nor U2848 (N_2848,N_1023,N_2157);
nor U2849 (N_2849,N_58,N_1240);
nor U2850 (N_2850,N_1475,N_1480);
nand U2851 (N_2851,N_715,N_1880);
and U2852 (N_2852,N_1219,N_2357);
or U2853 (N_2853,N_52,N_740);
and U2854 (N_2854,N_367,N_832);
or U2855 (N_2855,N_49,N_1854);
and U2856 (N_2856,N_2055,N_976);
nand U2857 (N_2857,N_1141,N_1739);
nor U2858 (N_2858,N_699,N_517);
or U2859 (N_2859,N_2441,N_262);
and U2860 (N_2860,N_688,N_1716);
and U2861 (N_2861,N_2148,N_538);
nand U2862 (N_2862,N_64,N_966);
or U2863 (N_2863,N_1390,N_667);
and U2864 (N_2864,N_169,N_1861);
xor U2865 (N_2865,N_277,N_1232);
xor U2866 (N_2866,N_1675,N_1810);
or U2867 (N_2867,N_2482,N_2154);
or U2868 (N_2868,N_1463,N_556);
or U2869 (N_2869,N_854,N_1986);
nand U2870 (N_2870,N_196,N_1115);
and U2871 (N_2871,N_744,N_291);
nand U2872 (N_2872,N_1010,N_1767);
nor U2873 (N_2873,N_2213,N_1236);
nand U2874 (N_2874,N_1351,N_439);
and U2875 (N_2875,N_845,N_1073);
and U2876 (N_2876,N_1975,N_1157);
or U2877 (N_2877,N_963,N_2314);
or U2878 (N_2878,N_2341,N_217);
nand U2879 (N_2879,N_1622,N_799);
nand U2880 (N_2880,N_2289,N_1098);
and U2881 (N_2881,N_2030,N_356);
or U2882 (N_2882,N_90,N_436);
nor U2883 (N_2883,N_1435,N_208);
nand U2884 (N_2884,N_69,N_1730);
nor U2885 (N_2885,N_1139,N_978);
and U2886 (N_2886,N_482,N_314);
nor U2887 (N_2887,N_1349,N_268);
or U2888 (N_2888,N_309,N_325);
nor U2889 (N_2889,N_1062,N_2017);
and U2890 (N_2890,N_84,N_117);
nor U2891 (N_2891,N_353,N_1824);
nor U2892 (N_2892,N_1640,N_1670);
and U2893 (N_2893,N_1976,N_1243);
nor U2894 (N_2894,N_1100,N_1618);
and U2895 (N_2895,N_1919,N_2319);
nor U2896 (N_2896,N_184,N_1692);
or U2897 (N_2897,N_1903,N_1574);
or U2898 (N_2898,N_1906,N_1514);
nor U2899 (N_2899,N_2493,N_75);
or U2900 (N_2900,N_54,N_1326);
and U2901 (N_2901,N_2027,N_2185);
and U2902 (N_2902,N_1414,N_2038);
nand U2903 (N_2903,N_731,N_1550);
and U2904 (N_2904,N_1500,N_1136);
nand U2905 (N_2905,N_1331,N_695);
nand U2906 (N_2906,N_2208,N_968);
nand U2907 (N_2907,N_242,N_1545);
nor U2908 (N_2908,N_541,N_2262);
or U2909 (N_2909,N_1216,N_1864);
and U2910 (N_2910,N_1731,N_1993);
nor U2911 (N_2911,N_1303,N_24);
nor U2912 (N_2912,N_1696,N_2258);
nand U2913 (N_2913,N_2405,N_1401);
and U2914 (N_2914,N_228,N_1703);
nand U2915 (N_2915,N_254,N_2014);
and U2916 (N_2916,N_389,N_2175);
or U2917 (N_2917,N_398,N_107);
and U2918 (N_2918,N_1633,N_815);
nand U2919 (N_2919,N_2162,N_2454);
nor U2920 (N_2920,N_2462,N_497);
and U2921 (N_2921,N_1541,N_1575);
nor U2922 (N_2922,N_1251,N_904);
or U2923 (N_2923,N_811,N_86);
nand U2924 (N_2924,N_2067,N_1802);
and U2925 (N_2925,N_581,N_1423);
nand U2926 (N_2926,N_2126,N_1486);
and U2927 (N_2927,N_929,N_2486);
nand U2928 (N_2928,N_1086,N_1587);
or U2929 (N_2929,N_2122,N_1358);
nor U2930 (N_2930,N_1194,N_2285);
nand U2931 (N_2931,N_910,N_2460);
and U2932 (N_2932,N_147,N_7);
nor U2933 (N_2933,N_949,N_27);
nor U2934 (N_2934,N_1567,N_914);
nand U2935 (N_2935,N_504,N_668);
nand U2936 (N_2936,N_2043,N_880);
nand U2937 (N_2937,N_1732,N_887);
nand U2938 (N_2938,N_1319,N_1121);
or U2939 (N_2939,N_2231,N_1811);
and U2940 (N_2940,N_933,N_1074);
xnor U2941 (N_2941,N_2463,N_2254);
and U2942 (N_2942,N_974,N_247);
or U2943 (N_2943,N_2344,N_788);
or U2944 (N_2944,N_2368,N_1851);
nor U2945 (N_2945,N_1736,N_1368);
nand U2946 (N_2946,N_2410,N_1666);
nor U2947 (N_2947,N_437,N_67);
nand U2948 (N_2948,N_1277,N_252);
or U2949 (N_2949,N_1566,N_269);
nor U2950 (N_2950,N_1488,N_1902);
and U2951 (N_2951,N_916,N_1138);
xor U2952 (N_2952,N_975,N_1589);
and U2953 (N_2953,N_2484,N_2382);
nor U2954 (N_2954,N_326,N_1518);
nor U2955 (N_2955,N_587,N_1292);
or U2956 (N_2956,N_2164,N_1971);
and U2957 (N_2957,N_1654,N_1789);
and U2958 (N_2958,N_1788,N_1539);
or U2959 (N_2959,N_911,N_223);
nand U2960 (N_2960,N_1261,N_267);
nor U2961 (N_2961,N_1599,N_288);
and U2962 (N_2962,N_493,N_1132);
nand U2963 (N_2963,N_1540,N_1613);
nand U2964 (N_2964,N_938,N_1689);
nor U2965 (N_2965,N_2359,N_1875);
nor U2966 (N_2966,N_1813,N_211);
nand U2967 (N_2967,N_16,N_743);
or U2968 (N_2968,N_1134,N_1648);
or U2969 (N_2969,N_42,N_505);
nand U2970 (N_2970,N_1402,N_1154);
and U2971 (N_2971,N_1620,N_387);
nor U2972 (N_2972,N_1915,N_1192);
or U2973 (N_2973,N_1325,N_578);
or U2974 (N_2974,N_2298,N_1561);
and U2975 (N_2975,N_406,N_802);
and U2976 (N_2976,N_232,N_21);
nor U2977 (N_2977,N_1012,N_656);
and U2978 (N_2978,N_645,N_89);
and U2979 (N_2979,N_2065,N_32);
nand U2980 (N_2980,N_414,N_616);
and U2981 (N_2981,N_1658,N_1956);
xor U2982 (N_2982,N_1750,N_1787);
nand U2983 (N_2983,N_1974,N_2104);
and U2984 (N_2984,N_921,N_153);
nor U2985 (N_2985,N_780,N_55);
or U2986 (N_2986,N_1890,N_1749);
or U2987 (N_2987,N_2204,N_359);
and U2988 (N_2988,N_1908,N_2002);
xor U2989 (N_2989,N_1982,N_298);
and U2990 (N_2990,N_227,N_623);
nor U2991 (N_2991,N_1360,N_1034);
nor U2992 (N_2992,N_1467,N_1306);
nor U2993 (N_2993,N_2173,N_241);
nand U2994 (N_2994,N_285,N_1274);
nor U2995 (N_2995,N_1471,N_240);
xor U2996 (N_2996,N_206,N_730);
or U2997 (N_2997,N_593,N_918);
and U2998 (N_2998,N_210,N_536);
or U2999 (N_2999,N_461,N_1148);
nor U3000 (N_3000,N_2241,N_514);
nor U3001 (N_3001,N_1220,N_225);
xnor U3002 (N_3002,N_546,N_294);
nand U3003 (N_3003,N_74,N_1799);
or U3004 (N_3004,N_610,N_1069);
or U3005 (N_3005,N_2290,N_2367);
nand U3006 (N_3006,N_588,N_1626);
nor U3007 (N_3007,N_307,N_433);
xor U3008 (N_3008,N_261,N_331);
nor U3009 (N_3009,N_1941,N_460);
nand U3010 (N_3010,N_2128,N_690);
and U3011 (N_3011,N_1819,N_859);
or U3012 (N_3012,N_2045,N_843);
or U3013 (N_3013,N_2101,N_2399);
or U3014 (N_3014,N_207,N_2054);
and U3015 (N_3015,N_1935,N_1083);
or U3016 (N_3016,N_2063,N_2020);
and U3017 (N_3017,N_1808,N_630);
nand U3018 (N_3018,N_2075,N_1804);
or U3019 (N_3019,N_619,N_1105);
nor U3020 (N_3020,N_2411,N_1771);
nor U3021 (N_3021,N_1728,N_1396);
nor U3022 (N_3022,N_374,N_2376);
nand U3023 (N_3023,N_1531,N_2112);
or U3024 (N_3024,N_973,N_411);
nand U3025 (N_3025,N_2029,N_604);
xnor U3026 (N_3026,N_1318,N_1312);
or U3027 (N_3027,N_2168,N_2227);
xnor U3028 (N_3028,N_2373,N_404);
or U3029 (N_3029,N_2211,N_29);
nor U3030 (N_3030,N_924,N_1961);
or U3031 (N_3031,N_1981,N_501);
and U3032 (N_3032,N_1643,N_1085);
and U3033 (N_3033,N_745,N_1870);
nor U3034 (N_3034,N_822,N_1273);
or U3035 (N_3035,N_1879,N_2297);
nor U3036 (N_3036,N_863,N_2453);
or U3037 (N_3037,N_547,N_2186);
nor U3038 (N_3038,N_607,N_609);
nand U3039 (N_3039,N_2040,N_2293);
nor U3040 (N_3040,N_1449,N_524);
nor U3041 (N_3041,N_575,N_265);
or U3042 (N_3042,N_2326,N_927);
and U3043 (N_3043,N_746,N_2256);
nor U3044 (N_3044,N_100,N_2325);
or U3045 (N_3045,N_1426,N_274);
and U3046 (N_3046,N_161,N_964);
and U3047 (N_3047,N_1610,N_1244);
nor U3048 (N_3048,N_1687,N_632);
and U3049 (N_3049,N_686,N_1287);
or U3050 (N_3050,N_2371,N_2392);
nor U3051 (N_3051,N_1433,N_993);
nor U3052 (N_3052,N_1370,N_1862);
and U3053 (N_3053,N_759,N_1825);
nor U3054 (N_3054,N_1683,N_78);
and U3055 (N_3055,N_2091,N_2338);
nor U3056 (N_3056,N_251,N_738);
and U3057 (N_3057,N_831,N_789);
and U3058 (N_3058,N_1095,N_1529);
xnor U3059 (N_3059,N_1181,N_510);
xor U3060 (N_3060,N_1482,N_2240);
nand U3061 (N_3061,N_37,N_378);
and U3062 (N_3062,N_1153,N_553);
and U3063 (N_3063,N_2280,N_1881);
nor U3064 (N_3064,N_868,N_765);
and U3065 (N_3065,N_321,N_264);
nor U3066 (N_3066,N_2271,N_1176);
nor U3067 (N_3067,N_1410,N_102);
nand U3068 (N_3068,N_1152,N_41);
and U3069 (N_3069,N_805,N_2200);
and U3070 (N_3070,N_2097,N_2102);
nor U3071 (N_3071,N_1653,N_1166);
or U3072 (N_3072,N_2184,N_2361);
nor U3073 (N_3073,N_2283,N_1766);
and U3074 (N_3074,N_1373,N_1904);
nand U3075 (N_3075,N_1004,N_591);
nor U3076 (N_3076,N_554,N_1679);
nand U3077 (N_3077,N_1366,N_2339);
or U3078 (N_3078,N_1553,N_824);
and U3079 (N_3079,N_2238,N_794);
nor U3080 (N_3080,N_1901,N_1258);
xor U3081 (N_3081,N_278,N_1017);
and U3082 (N_3082,N_567,N_1912);
nor U3083 (N_3083,N_1163,N_995);
xor U3084 (N_3084,N_1501,N_2088);
and U3085 (N_3085,N_445,N_1955);
nand U3086 (N_3086,N_2011,N_804);
and U3087 (N_3087,N_1898,N_2179);
nor U3088 (N_3088,N_2093,N_1655);
nand U3089 (N_3089,N_507,N_56);
nor U3090 (N_3090,N_1070,N_2430);
nand U3091 (N_3091,N_2212,N_2427);
or U3092 (N_3092,N_427,N_2183);
or U3093 (N_3093,N_1367,N_1853);
or U3094 (N_3094,N_1979,N_2451);
nor U3095 (N_3095,N_1735,N_1763);
nor U3096 (N_3096,N_1037,N_1515);
or U3097 (N_3097,N_1046,N_315);
or U3098 (N_3098,N_230,N_484);
nand U3099 (N_3099,N_1293,N_1415);
and U3100 (N_3100,N_647,N_664);
or U3101 (N_3101,N_2031,N_2130);
or U3102 (N_3102,N_249,N_311);
or U3103 (N_3103,N_1745,N_2123);
nand U3104 (N_3104,N_36,N_897);
nand U3105 (N_3105,N_1662,N_1437);
nor U3106 (N_3106,N_625,N_401);
nand U3107 (N_3107,N_653,N_2331);
and U3108 (N_3108,N_1994,N_827);
nor U3109 (N_3109,N_709,N_2478);
or U3110 (N_3110,N_992,N_1959);
and U3111 (N_3111,N_2397,N_478);
or U3112 (N_3112,N_1272,N_2442);
nor U3113 (N_3113,N_1188,N_1383);
or U3114 (N_3114,N_449,N_2202);
nor U3115 (N_3115,N_198,N_2199);
nor U3116 (N_3116,N_2415,N_2491);
nand U3117 (N_3117,N_1185,N_842);
nand U3118 (N_3118,N_2105,N_165);
nor U3119 (N_3119,N_101,N_1899);
or U3120 (N_3120,N_2012,N_873);
and U3121 (N_3121,N_2267,N_958);
nand U3122 (N_3122,N_795,N_1421);
or U3123 (N_3123,N_2174,N_30);
or U3124 (N_3124,N_2178,N_687);
and U3125 (N_3125,N_1101,N_115);
nor U3126 (N_3126,N_1933,N_1774);
or U3127 (N_3127,N_1611,N_1659);
or U3128 (N_3128,N_2244,N_644);
xor U3129 (N_3129,N_1031,N_384);
nor U3130 (N_3130,N_797,N_140);
or U3131 (N_3131,N_2324,N_292);
nand U3132 (N_3132,N_1204,N_1071);
nand U3133 (N_3133,N_9,N_166);
nand U3134 (N_3134,N_1573,N_724);
nand U3135 (N_3135,N_2295,N_1197);
and U3136 (N_3136,N_986,N_1839);
nor U3137 (N_3137,N_2265,N_1913);
or U3138 (N_3138,N_516,N_119);
or U3139 (N_3139,N_1704,N_216);
nand U3140 (N_3140,N_753,N_527);
or U3141 (N_3141,N_577,N_469);
and U3142 (N_3142,N_2044,N_1562);
or U3143 (N_3143,N_1669,N_2233);
nand U3144 (N_3144,N_339,N_63);
nand U3145 (N_3145,N_953,N_1544);
nand U3146 (N_3146,N_2432,N_2473);
and U3147 (N_3147,N_1831,N_801);
and U3148 (N_3148,N_2225,N_1663);
nor U3149 (N_3149,N_614,N_1962);
nand U3150 (N_3150,N_2166,N_2268);
and U3151 (N_3151,N_2144,N_456);
nand U3152 (N_3152,N_611,N_1595);
nor U3153 (N_3153,N_1718,N_706);
nor U3154 (N_3154,N_379,N_1087);
or U3155 (N_3155,N_88,N_1743);
and U3156 (N_3156,N_2266,N_1701);
and U3157 (N_3157,N_626,N_1007);
or U3158 (N_3158,N_1283,N_159);
nand U3159 (N_3159,N_1015,N_1301);
or U3160 (N_3160,N_1458,N_205);
nand U3161 (N_3161,N_1019,N_61);
or U3162 (N_3162,N_1270,N_766);
nor U3163 (N_3163,N_725,N_1721);
nand U3164 (N_3164,N_2278,N_2499);
or U3165 (N_3165,N_351,N_203);
or U3166 (N_3166,N_886,N_2224);
nand U3167 (N_3167,N_1637,N_2340);
nand U3168 (N_3168,N_2355,N_1768);
nor U3169 (N_3169,N_861,N_1921);
and U3170 (N_3170,N_2301,N_837);
or U3171 (N_3171,N_477,N_2282);
or U3172 (N_3172,N_2365,N_817);
nand U3173 (N_3173,N_1872,N_600);
nor U3174 (N_3174,N_1418,N_1871);
or U3175 (N_3175,N_2389,N_1920);
nor U3176 (N_3176,N_739,N_1445);
nor U3177 (N_3177,N_1623,N_1080);
nand U3178 (N_3178,N_1505,N_1490);
nand U3179 (N_3179,N_1040,N_2074);
or U3180 (N_3180,N_355,N_1448);
and U3181 (N_3181,N_96,N_1700);
nand U3182 (N_3182,N_1469,N_1404);
nand U3183 (N_3183,N_1499,N_365);
xnor U3184 (N_3184,N_300,N_1242);
xor U3185 (N_3185,N_2428,N_13);
nand U3186 (N_3186,N_2139,N_655);
and U3187 (N_3187,N_2446,N_583);
nand U3188 (N_3188,N_2061,N_2272);
or U3189 (N_3189,N_323,N_324);
nand U3190 (N_3190,N_1699,N_2412);
and U3191 (N_3191,N_530,N_1186);
nor U3192 (N_3192,N_1786,N_825);
and U3193 (N_3193,N_2449,N_342);
and U3194 (N_3194,N_1773,N_1229);
or U3195 (N_3195,N_452,N_2418);
nand U3196 (N_3196,N_508,N_1481);
or U3197 (N_3197,N_917,N_748);
nor U3198 (N_3198,N_635,N_735);
nand U3199 (N_3199,N_1089,N_458);
or U3200 (N_3200,N_776,N_711);
nor U3201 (N_3201,N_266,N_515);
and U3202 (N_3202,N_93,N_2448);
or U3203 (N_3203,N_1035,N_1684);
nor U3204 (N_3204,N_1591,N_471);
or U3205 (N_3205,N_1533,N_708);
or U3206 (N_3206,N_1964,N_2379);
nor U3207 (N_3207,N_1092,N_53);
nor U3208 (N_3208,N_602,N_479);
and U3209 (N_3209,N_1472,N_1142);
or U3210 (N_3210,N_1338,N_1558);
nand U3211 (N_3211,N_913,N_2010);
nor U3212 (N_3212,N_1895,N_1709);
or U3213 (N_3213,N_429,N_1335);
nor U3214 (N_3214,N_1968,N_1647);
nor U3215 (N_3215,N_551,N_391);
nand U3216 (N_3216,N_1042,N_2076);
nor U3217 (N_3217,N_545,N_1461);
or U3218 (N_3218,N_1569,N_2458);
nand U3219 (N_3219,N_2333,N_40);
and U3220 (N_3220,N_457,N_488);
and U3221 (N_3221,N_1320,N_962);
nand U3222 (N_3222,N_1535,N_786);
and U3223 (N_3223,N_1036,N_103);
nand U3224 (N_3224,N_1168,N_1253);
or U3225 (N_3225,N_528,N_2354);
xor U3226 (N_3226,N_2300,N_2409);
nor U3227 (N_3227,N_149,N_143);
nor U3228 (N_3228,N_2464,N_721);
nand U3229 (N_3229,N_961,N_106);
and U3230 (N_3230,N_190,N_713);
and U3231 (N_3231,N_1951,N_2437);
nor U3232 (N_3232,N_852,N_2287);
or U3233 (N_3233,N_895,N_1296);
nor U3234 (N_3234,N_1485,N_229);
and U3235 (N_3235,N_582,N_1195);
or U3236 (N_3236,N_1927,N_572);
or U3237 (N_3237,N_1998,N_1409);
or U3238 (N_3238,N_663,N_317);
and U3239 (N_3239,N_6,N_729);
nor U3240 (N_3240,N_893,N_2042);
and U3241 (N_3241,N_1536,N_2107);
nand U3242 (N_3242,N_876,N_970);
nand U3243 (N_3243,N_660,N_1405);
nand U3244 (N_3244,N_1328,N_22);
and U3245 (N_3245,N_1823,N_1604);
nor U3246 (N_3246,N_629,N_723);
xor U3247 (N_3247,N_2026,N_1817);
nand U3248 (N_3248,N_19,N_638);
and U3249 (N_3249,N_720,N_1930);
or U3250 (N_3250,N_2095,N_2402);
nor U3251 (N_3251,N_1417,N_1954);
nand U3252 (N_3252,N_246,N_1578);
and U3253 (N_3253,N_1022,N_348);
and U3254 (N_3254,N_1455,N_1747);
and U3255 (N_3255,N_1382,N_1350);
nand U3256 (N_3256,N_2417,N_2163);
or U3257 (N_3257,N_1866,N_236);
nand U3258 (N_3258,N_173,N_1516);
or U3259 (N_3259,N_1361,N_255);
nor U3260 (N_3260,N_1108,N_480);
and U3261 (N_3261,N_1056,N_666);
or U3262 (N_3262,N_969,N_295);
and U3263 (N_3263,N_286,N_336);
nand U3264 (N_3264,N_2461,N_1342);
or U3265 (N_3265,N_2263,N_128);
nor U3266 (N_3266,N_1376,N_752);
nand U3267 (N_3267,N_2374,N_237);
or U3268 (N_3268,N_171,N_1375);
or U3269 (N_3269,N_2330,N_1816);
nor U3270 (N_3270,N_1512,N_809);
or U3271 (N_3271,N_1957,N_2106);
nor U3272 (N_3272,N_1308,N_1341);
nor U3273 (N_3273,N_2414,N_513);
nor U3274 (N_3274,N_1571,N_2080);
nor U3275 (N_3275,N_965,N_1084);
and U3276 (N_3276,N_1820,N_1057);
or U3277 (N_3277,N_2475,N_2006);
and U3278 (N_3278,N_338,N_310);
nor U3279 (N_3279,N_233,N_299);
nand U3280 (N_3280,N_1922,N_1173);
nor U3281 (N_3281,N_728,N_2433);
nor U3282 (N_3282,N_1775,N_87);
nor U3283 (N_3283,N_1717,N_33);
and U3284 (N_3284,N_1690,N_902);
nor U3285 (N_3285,N_2257,N_1088);
xnor U3286 (N_3286,N_1394,N_451);
and U3287 (N_3287,N_283,N_892);
nor U3288 (N_3288,N_2304,N_2087);
nor U3289 (N_3289,N_2288,N_2099);
xor U3290 (N_3290,N_1524,N_742);
nor U3291 (N_3291,N_1468,N_2082);
nor U3292 (N_3292,N_2215,N_463);
nor U3293 (N_3293,N_772,N_1832);
or U3294 (N_3294,N_189,N_1110);
nand U3295 (N_3295,N_1983,N_839);
nand U3296 (N_3296,N_1827,N_957);
and U3297 (N_3297,N_1460,N_2008);
and U3298 (N_3298,N_2141,N_1201);
nor U3299 (N_3299,N_1869,N_1446);
nor U3300 (N_3300,N_2416,N_2062);
or U3301 (N_3301,N_1000,N_1159);
nor U3302 (N_3302,N_853,N_79);
or U3303 (N_3303,N_141,N_2360);
nor U3304 (N_3304,N_1772,N_1440);
nor U3305 (N_3305,N_1060,N_2193);
and U3306 (N_3306,N_2207,N_1797);
nor U3307 (N_3307,N_1030,N_2468);
nand U3308 (N_3308,N_1973,N_1926);
nor U3309 (N_3309,N_2140,N_1708);
nand U3310 (N_3310,N_526,N_1315);
and U3311 (N_3311,N_1208,N_70);
nand U3312 (N_3312,N_1984,N_1412);
nand U3313 (N_3313,N_2221,N_183);
or U3314 (N_3314,N_245,N_818);
nand U3315 (N_3315,N_2071,N_43);
or U3316 (N_3316,N_1624,N_903);
nor U3317 (N_3317,N_1615,N_494);
and U3318 (N_3318,N_1045,N_503);
nand U3319 (N_3319,N_2394,N_2347);
nand U3320 (N_3320,N_191,N_1096);
nor U3321 (N_3321,N_2385,N_696);
or U3322 (N_3322,N_2138,N_1093);
nand U3323 (N_3323,N_260,N_1476);
nor U3324 (N_3324,N_1199,N_1266);
or U3325 (N_3325,N_2210,N_1761);
nand U3326 (N_3326,N_2176,N_1657);
or U3327 (N_3327,N_885,N_1411);
nor U3328 (N_3328,N_66,N_322);
and U3329 (N_3329,N_2232,N_1127);
and U3330 (N_3330,N_438,N_123);
nand U3331 (N_3331,N_2090,N_130);
and U3332 (N_3332,N_2132,N_2242);
nor U3333 (N_3333,N_2203,N_760);
xnor U3334 (N_3334,N_2019,N_539);
nand U3335 (N_3335,N_757,N_884);
nor U3336 (N_3336,N_2334,N_1523);
and U3337 (N_3337,N_573,N_467);
nand U3338 (N_3338,N_98,N_2239);
nor U3339 (N_3339,N_2476,N_1502);
and U3340 (N_3340,N_1507,N_1752);
or U3341 (N_3341,N_432,N_1442);
and U3342 (N_3342,N_1169,N_1447);
or U3343 (N_3343,N_327,N_1989);
and U3344 (N_3344,N_532,N_1330);
nand U3345 (N_3345,N_2169,N_1051);
nor U3346 (N_3346,N_512,N_2323);
nor U3347 (N_3347,N_613,N_941);
nand U3348 (N_3348,N_18,N_816);
nor U3349 (N_3349,N_2028,N_2312);
or U3350 (N_3350,N_1900,N_586);
nand U3351 (N_3351,N_1492,N_1660);
nor U3352 (N_3352,N_1520,N_2151);
and U3353 (N_3353,N_869,N_1606);
and U3354 (N_3354,N_243,N_698);
nor U3355 (N_3355,N_486,N_1614);
and U3356 (N_3356,N_594,N_1695);
nor U3357 (N_3357,N_923,N_1049);
nor U3358 (N_3358,N_443,N_793);
xor U3359 (N_3359,N_674,N_1032);
nand U3360 (N_3360,N_2146,N_2321);
or U3361 (N_3361,N_1970,N_2197);
nor U3362 (N_3362,N_552,N_967);
nor U3363 (N_3363,N_2243,N_1504);
and U3364 (N_3364,N_1450,N_775);
or U3365 (N_3365,N_649,N_636);
nor U3366 (N_3366,N_1081,N_1205);
nor U3367 (N_3367,N_1754,N_662);
nand U3368 (N_3368,N_424,N_1585);
xor U3369 (N_3369,N_1061,N_110);
or U3370 (N_3370,N_1770,N_306);
and U3371 (N_3371,N_838,N_2328);
or U3372 (N_3372,N_1978,N_671);
nand U3373 (N_3373,N_560,N_2222);
nand U3374 (N_3374,N_124,N_120);
or U3375 (N_3375,N_363,N_784);
nand U3376 (N_3376,N_2103,N_1454);
or U3377 (N_3377,N_1279,N_10);
or U3378 (N_3378,N_1406,N_2422);
and U3379 (N_3379,N_284,N_2429);
or U3380 (N_3380,N_1759,N_1392);
nor U3381 (N_3381,N_682,N_2214);
nor U3382 (N_3382,N_747,N_1762);
or U3383 (N_3383,N_1697,N_2313);
nor U3384 (N_3384,N_423,N_1380);
nor U3385 (N_3385,N_1532,N_998);
nand U3386 (N_3386,N_1744,N_1212);
nor U3387 (N_3387,N_20,N_564);
xor U3388 (N_3388,N_1785,N_1942);
nor U3389 (N_3389,N_833,N_2309);
and U3390 (N_3390,N_1217,N_1782);
nand U3391 (N_3391,N_2335,N_718);
or U3392 (N_3392,N_318,N_1631);
nor U3393 (N_3393,N_113,N_1465);
and U3394 (N_3394,N_2426,N_657);
and U3395 (N_3395,N_1477,N_798);
nor U3396 (N_3396,N_231,N_2249);
nand U3397 (N_3397,N_972,N_984);
or U3398 (N_3398,N_694,N_1365);
and U3399 (N_3399,N_1224,N_2135);
nand U3400 (N_3400,N_1818,N_888);
nand U3401 (N_3401,N_858,N_1688);
or U3402 (N_3402,N_2245,N_139);
or U3403 (N_3403,N_952,N_199);
nand U3404 (N_3404,N_2016,N_303);
and U3405 (N_3405,N_410,N_790);
nand U3406 (N_3406,N_1678,N_1534);
nor U3407 (N_3407,N_1513,N_1316);
and U3408 (N_3408,N_2306,N_1231);
nor U3409 (N_3409,N_1642,N_170);
or U3410 (N_3410,N_1849,N_982);
nor U3411 (N_3411,N_1117,N_83);
or U3412 (N_3412,N_557,N_465);
and U3413 (N_3413,N_569,N_693);
and U3414 (N_3414,N_162,N_896);
xnor U3415 (N_3415,N_542,N_168);
or U3416 (N_3416,N_1639,N_1091);
or U3417 (N_3417,N_1299,N_1289);
or U3418 (N_3418,N_1630,N_1671);
nand U3419 (N_3419,N_2329,N_1943);
and U3420 (N_3420,N_426,N_289);
or U3421 (N_3421,N_1311,N_509);
and U3422 (N_3422,N_511,N_2356);
or U3423 (N_3423,N_1230,N_1203);
and U3424 (N_3424,N_1634,N_2270);
nor U3425 (N_3425,N_531,N_72);
and U3426 (N_3426,N_2060,N_768);
nor U3427 (N_3427,N_856,N_1352);
nand U3428 (N_3428,N_624,N_1842);
or U3429 (N_3429,N_48,N_937);
or U3430 (N_3430,N_939,N_862);
nor U3431 (N_3431,N_2362,N_1167);
nand U3432 (N_3432,N_1429,N_23);
nand U3433 (N_3433,N_2404,N_1803);
or U3434 (N_3434,N_1190,N_2390);
nor U3435 (N_3435,N_2009,N_1182);
or U3436 (N_3436,N_2021,N_812);
and U3437 (N_3437,N_701,N_2094);
and U3438 (N_3438,N_646,N_376);
nand U3439 (N_3439,N_1294,N_951);
or U3440 (N_3440,N_1559,N_215);
nor U3441 (N_3441,N_1267,N_741);
nand U3442 (N_3442,N_1379,N_1420);
or U3443 (N_3443,N_71,N_1055);
nand U3444 (N_3444,N_1729,N_840);
nand U3445 (N_3445,N_1910,N_383);
and U3446 (N_3446,N_2400,N_1398);
nor U3447 (N_3447,N_152,N_2443);
and U3448 (N_3448,N_650,N_637);
nand U3449 (N_3449,N_1629,N_2089);
and U3450 (N_3450,N_1438,N_412);
nor U3451 (N_3451,N_1099,N_877);
and U3452 (N_3452,N_1742,N_1740);
nor U3453 (N_3453,N_421,N_1193);
nor U3454 (N_3454,N_416,N_2086);
xnor U3455 (N_3455,N_1210,N_2395);
and U3456 (N_3456,N_305,N_754);
nand U3457 (N_3457,N_1237,N_1845);
and U3458 (N_3458,N_187,N_1737);
nor U3459 (N_3459,N_1013,N_2023);
nand U3460 (N_3460,N_1554,N_628);
nand U3461 (N_3461,N_1594,N_1521);
nor U3462 (N_3462,N_680,N_841);
or U3463 (N_3463,N_1990,N_1581);
nand U3464 (N_3464,N_1850,N_2083);
nand U3465 (N_3465,N_1222,N_1503);
nor U3466 (N_3466,N_157,N_1597);
or U3467 (N_3467,N_1713,N_1760);
or U3468 (N_3468,N_533,N_2358);
and U3469 (N_3469,N_764,N_777);
nand U3470 (N_3470,N_1498,N_212);
and U3471 (N_3471,N_1002,N_1395);
nor U3472 (N_3472,N_2005,N_2387);
xor U3473 (N_3473,N_1548,N_1780);
nor U3474 (N_3474,N_263,N_1202);
nor U3475 (N_3475,N_1635,N_1113);
or U3476 (N_3476,N_617,N_988);
nor U3477 (N_3477,N_2013,N_2237);
xnor U3478 (N_3478,N_1453,N_346);
nand U3479 (N_3479,N_121,N_506);
or U3480 (N_3480,N_954,N_1029);
nand U3481 (N_3481,N_202,N_823);
or U3482 (N_3482,N_692,N_851);
nand U3483 (N_3483,N_2403,N_1484);
nand U3484 (N_3484,N_1304,N_2311);
nand U3485 (N_3485,N_1748,N_922);
or U3486 (N_3486,N_1179,N_1323);
nor U3487 (N_3487,N_2467,N_394);
nand U3488 (N_3488,N_1911,N_393);
and U3489 (N_3489,N_97,N_347);
nand U3490 (N_3490,N_2110,N_2229);
nand U3491 (N_3491,N_1050,N_1705);
and U3492 (N_3492,N_1233,N_194);
and U3493 (N_3493,N_518,N_2153);
xor U3494 (N_3494,N_1924,N_2092);
nand U3495 (N_3495,N_1727,N_2025);
and U3496 (N_3496,N_2363,N_579);
and U3497 (N_3497,N_1211,N_1094);
and U3498 (N_3498,N_920,N_1345);
or U3499 (N_3499,N_1707,N_2181);
nand U3500 (N_3500,N_1172,N_889);
or U3501 (N_3501,N_2294,N_25);
or U3502 (N_3502,N_1972,N_684);
nand U3503 (N_3503,N_2273,N_2147);
nand U3504 (N_3504,N_1162,N_960);
nor U3505 (N_3505,N_163,N_1072);
nor U3506 (N_3506,N_707,N_2081);
or U3507 (N_3507,N_1897,N_485);
and U3508 (N_3508,N_188,N_1783);
nor U3509 (N_3509,N_585,N_1381);
and U3510 (N_3510,N_800,N_1497);
or U3511 (N_3511,N_830,N_1302);
and U3512 (N_3512,N_627,N_1874);
nand U3513 (N_3513,N_1724,N_2192);
and U3514 (N_3514,N_1511,N_2369);
nor U3515 (N_3515,N_1281,N_475);
or U3516 (N_3516,N_1116,N_1149);
and U3517 (N_3517,N_1090,N_2057);
and U3518 (N_3518,N_2115,N_2056);
and U3519 (N_3519,N_883,N_2117);
nand U3520 (N_3520,N_1592,N_791);
nand U3521 (N_3521,N_1430,N_756);
nand U3522 (N_3522,N_221,N_2353);
nor U3523 (N_3523,N_2066,N_1712);
and U3524 (N_3524,N_2111,N_1425);
nand U3525 (N_3525,N_2284,N_2346);
xnor U3526 (N_3526,N_1522,N_1126);
and U3527 (N_3527,N_714,N_782);
nand U3528 (N_3528,N_543,N_673);
and U3529 (N_3529,N_1932,N_2172);
and U3530 (N_3530,N_931,N_1952);
xor U3531 (N_3531,N_814,N_31);
and U3532 (N_3532,N_946,N_813);
or U3533 (N_3533,N_1282,N_2195);
or U3534 (N_3534,N_341,N_1206);
and U3535 (N_3535,N_1652,N_1364);
nand U3536 (N_3536,N_1603,N_1596);
nand U3537 (N_3537,N_955,N_272);
nor U3538 (N_3538,N_615,N_1576);
or U3539 (N_3539,N_134,N_473);
and U3540 (N_3540,N_1295,N_2348);
xor U3541 (N_3541,N_320,N_281);
nor U3542 (N_3542,N_935,N_652);
nand U3543 (N_3543,N_425,N_441);
and U3544 (N_3544,N_51,N_403);
nor U3545 (N_3545,N_308,N_1537);
and U3546 (N_3546,N_2161,N_335);
nand U3547 (N_3547,N_574,N_979);
nor U3548 (N_3548,N_1784,N_1517);
and U3549 (N_3549,N_1109,N_778);
and U3550 (N_3550,N_2190,N_2053);
and U3551 (N_3551,N_2303,N_1877);
nand U3552 (N_3552,N_769,N_940);
nor U3553 (N_3553,N_1280,N_1371);
or U3554 (N_3554,N_1582,N_1334);
and U3555 (N_3555,N_1565,N_1156);
nor U3556 (N_3556,N_2182,N_448);
nor U3557 (N_3557,N_612,N_396);
xnor U3558 (N_3558,N_1838,N_1722);
and U3559 (N_3559,N_2407,N_601);
nand U3560 (N_3560,N_1557,N_1255);
nor U3561 (N_3561,N_1452,N_618);
nand U3562 (N_3562,N_2001,N_1888);
and U3563 (N_3563,N_136,N_1286);
nand U3564 (N_3564,N_95,N_727);
and U3565 (N_3565,N_1075,N_1114);
or U3566 (N_3566,N_810,N_1833);
or U3567 (N_3567,N_418,N_304);
or U3568 (N_3568,N_1715,N_160);
nor U3569 (N_3569,N_2398,N_1677);
and U3570 (N_3570,N_2253,N_2380);
nor U3571 (N_3571,N_186,N_1006);
nand U3572 (N_3572,N_1389,N_2096);
and U3573 (N_3573,N_2230,N_1018);
or U3574 (N_3574,N_1896,N_2469);
and U3575 (N_3575,N_1009,N_1847);
or U3576 (N_3576,N_1931,N_2118);
nor U3577 (N_3577,N_2085,N_45);
nand U3578 (N_3578,N_737,N_1980);
xor U3579 (N_3579,N_1359,N_1332);
or U3580 (N_3580,N_781,N_167);
and U3581 (N_3581,N_2035,N_385);
nor U3582 (N_3582,N_1588,N_639);
and U3583 (N_3583,N_250,N_1313);
nand U3584 (N_3584,N_875,N_1681);
and U3585 (N_3585,N_116,N_1836);
and U3586 (N_3586,N_2133,N_2351);
nand U3587 (N_3587,N_302,N_2171);
and U3588 (N_3588,N_1041,N_1337);
nor U3589 (N_3589,N_1579,N_1868);
nand U3590 (N_3590,N_994,N_405);
nor U3591 (N_3591,N_112,N_948);
or U3592 (N_3592,N_850,N_705);
and U3593 (N_3593,N_1439,N_1487);
nor U3594 (N_3594,N_420,N_808);
nand U3595 (N_3595,N_1043,N_444);
and U3596 (N_3596,N_1118,N_1158);
and U3597 (N_3597,N_2098,N_1183);
nand U3598 (N_3598,N_312,N_1362);
or U3599 (N_3599,N_855,N_145);
nand U3600 (N_3600,N_197,N_1609);
nor U3601 (N_3601,N_1053,N_1806);
nor U3602 (N_3602,N_1694,N_712);
nor U3603 (N_3603,N_1170,N_2129);
nor U3604 (N_3604,N_1863,N_943);
or U3605 (N_3605,N_648,N_1107);
nand U3606 (N_3606,N_985,N_1259);
or U3607 (N_3607,N_1682,N_1245);
or U3608 (N_3608,N_105,N_1672);
or U3609 (N_3609,N_2125,N_2051);
nand U3610 (N_3610,N_1885,N_2352);
nand U3611 (N_3611,N_1354,N_1457);
nor U3612 (N_3612,N_857,N_580);
and U3613 (N_3613,N_131,N_785);
or U3614 (N_3614,N_565,N_440);
nand U3615 (N_3615,N_1413,N_796);
nand U3616 (N_3616,N_2320,N_135);
or U3617 (N_3617,N_483,N_380);
nor U3618 (N_3618,N_256,N_431);
nor U3619 (N_3619,N_697,N_1509);
or U3620 (N_3620,N_148,N_2116);
and U3621 (N_3621,N_658,N_669);
and U3622 (N_3622,N_328,N_912);
and U3623 (N_3623,N_906,N_1988);
nand U3624 (N_3624,N_1821,N_894);
or U3625 (N_3625,N_2022,N_999);
nor U3626 (N_3626,N_434,N_235);
nor U3627 (N_3627,N_1945,N_1256);
nand U3628 (N_3628,N_65,N_2277);
nor U3629 (N_3629,N_82,N_2177);
xnor U3630 (N_3630,N_1178,N_1848);
nand U3631 (N_3631,N_631,N_945);
and U3632 (N_3632,N_26,N_2217);
and U3633 (N_3633,N_544,N_1077);
or U3634 (N_3634,N_1400,N_2470);
or U3635 (N_3635,N_447,N_92);
nor U3636 (N_3636,N_622,N_1112);
and U3637 (N_3637,N_734,N_381);
nand U3638 (N_3638,N_2296,N_137);
and U3639 (N_3639,N_11,N_409);
and U3640 (N_3640,N_293,N_2383);
nor U3641 (N_3641,N_2393,N_2);
or U3642 (N_3642,N_388,N_1769);
nor U3643 (N_3643,N_1778,N_94);
nand U3644 (N_3644,N_435,N_290);
and U3645 (N_3645,N_1873,N_142);
or U3646 (N_3646,N_1155,N_1917);
or U3647 (N_3647,N_1111,N_1067);
nor U3648 (N_3648,N_525,N_1431);
or U3649 (N_3649,N_605,N_2345);
or U3650 (N_3650,N_661,N_2370);
nand U3651 (N_3651,N_462,N_779);
xnor U3652 (N_3652,N_50,N_529);
or U3653 (N_3653,N_2305,N_1764);
nor U3654 (N_3654,N_316,N_133);
or U3655 (N_3655,N_763,N_28);
or U3656 (N_3656,N_990,N_592);
or U3657 (N_3657,N_2248,N_570);
and U3658 (N_3658,N_959,N_1746);
or U3659 (N_3659,N_1068,N_104);
and U3660 (N_3660,N_1317,N_68);
or U3661 (N_3661,N_1191,N_633);
nand U3662 (N_3662,N_620,N_1441);
or U3663 (N_3663,N_1218,N_1466);
and U3664 (N_3664,N_1496,N_700);
and U3665 (N_3665,N_1066,N_382);
and U3666 (N_3666,N_2046,N_821);
and U3667 (N_3667,N_1355,N_2216);
nor U3668 (N_3668,N_606,N_925);
nand U3669 (N_3669,N_390,N_330);
nor U3670 (N_3670,N_2170,N_2459);
xor U3671 (N_3671,N_2137,N_1857);
xor U3672 (N_3672,N_1602,N_2004);
nand U3673 (N_3673,N_1016,N_1184);
nand U3674 (N_3674,N_1598,N_146);
nor U3675 (N_3675,N_1269,N_2209);
or U3676 (N_3676,N_2234,N_2274);
or U3677 (N_3677,N_1028,N_2068);
nand U3678 (N_3678,N_1140,N_1014);
nor U3679 (N_3679,N_1483,N_349);
and U3680 (N_3680,N_2483,N_1097);
nand U3681 (N_3681,N_907,N_1963);
and U3682 (N_3682,N_719,N_2420);
nor U3683 (N_3683,N_942,N_1120);
nand U3684 (N_3684,N_2492,N_1076);
nor U3685 (N_3685,N_1078,N_337);
nand U3686 (N_3686,N_280,N_773);
nand U3687 (N_3687,N_2472,N_1621);
nor U3688 (N_3688,N_334,N_343);
or U3689 (N_3689,N_770,N_1680);
nor U3690 (N_3690,N_1241,N_5);
nor U3691 (N_3691,N_828,N_76);
nor U3692 (N_3692,N_185,N_386);
and U3693 (N_3693,N_1298,N_1038);
nand U3694 (N_3694,N_1815,N_1346);
nand U3695 (N_3695,N_2032,N_599);
or U3696 (N_3696,N_2003,N_1024);
nand U3697 (N_3697,N_596,N_476);
or U3698 (N_3698,N_1858,N_357);
nand U3699 (N_3699,N_2438,N_1257);
nor U3700 (N_3700,N_1805,N_1995);
or U3701 (N_3701,N_2457,N_2332);
or U3702 (N_3702,N_1187,N_2079);
or U3703 (N_3703,N_1725,N_132);
and U3704 (N_3704,N_2114,N_1161);
and U3705 (N_3705,N_181,N_1948);
nand U3706 (N_3706,N_1307,N_77);
and U3707 (N_3707,N_2419,N_372);
nor U3708 (N_3708,N_1665,N_2247);
xor U3709 (N_3709,N_1252,N_1893);
or U3710 (N_3710,N_1103,N_1894);
and U3711 (N_3711,N_598,N_2187);
and U3712 (N_3712,N_1734,N_80);
and U3713 (N_3713,N_2041,N_464);
or U3714 (N_3714,N_2246,N_2113);
or U3715 (N_3715,N_1336,N_726);
nor U3716 (N_3716,N_2018,N_1829);
or U3717 (N_3717,N_1260,N_2445);
and U3718 (N_3718,N_2165,N_774);
and U3719 (N_3719,N_1644,N_2310);
or U3720 (N_3720,N_1275,N_154);
nor U3721 (N_3721,N_219,N_214);
or U3722 (N_3722,N_1649,N_2158);
nand U3723 (N_3723,N_1792,N_1656);
and U3724 (N_3724,N_537,N_248);
nand U3725 (N_3725,N_1478,N_1969);
and U3726 (N_3726,N_450,N_1254);
nand U3727 (N_3727,N_59,N_2160);
nor U3728 (N_3728,N_2490,N_1285);
nand U3729 (N_3729,N_2336,N_1676);
nand U3730 (N_3730,N_2307,N_375);
nor U3731 (N_3731,N_2072,N_1809);
and U3732 (N_3732,N_672,N_834);
nor U3733 (N_3733,N_150,N_1344);
or U3734 (N_3734,N_2109,N_466);
and U3735 (N_3735,N_14,N_4);
nor U3736 (N_3736,N_1175,N_549);
or U3737 (N_3737,N_1719,N_1493);
nand U3738 (N_3738,N_1600,N_689);
or U3739 (N_3739,N_1667,N_1882);
nor U3740 (N_3740,N_15,N_1583);
nand U3741 (N_3741,N_1387,N_1892);
nand U3742 (N_3742,N_879,N_2142);
nor U3743 (N_3743,N_2264,N_454);
nand U3744 (N_3744,N_1668,N_2452);
nand U3745 (N_3745,N_2121,N_1584);
and U3746 (N_3746,N_2481,N_2205);
and U3747 (N_3747,N_1546,N_1826);
nand U3748 (N_3748,N_176,N_415);
or U3749 (N_3749,N_659,N_1391);
and U3750 (N_3750,N_1642,N_827);
nand U3751 (N_3751,N_827,N_380);
and U3752 (N_3752,N_276,N_947);
nand U3753 (N_3753,N_1774,N_608);
and U3754 (N_3754,N_2016,N_1809);
or U3755 (N_3755,N_1569,N_1374);
nand U3756 (N_3756,N_2037,N_1204);
nand U3757 (N_3757,N_1821,N_2);
nand U3758 (N_3758,N_588,N_692);
nor U3759 (N_3759,N_885,N_1555);
nand U3760 (N_3760,N_120,N_2062);
or U3761 (N_3761,N_1614,N_1209);
xnor U3762 (N_3762,N_897,N_1161);
nor U3763 (N_3763,N_1944,N_1996);
and U3764 (N_3764,N_1377,N_482);
and U3765 (N_3765,N_1853,N_2048);
and U3766 (N_3766,N_305,N_2493);
nor U3767 (N_3767,N_2113,N_150);
xor U3768 (N_3768,N_117,N_1718);
nand U3769 (N_3769,N_1825,N_1035);
nor U3770 (N_3770,N_745,N_169);
nor U3771 (N_3771,N_809,N_187);
and U3772 (N_3772,N_411,N_377);
nand U3773 (N_3773,N_350,N_802);
and U3774 (N_3774,N_545,N_229);
nor U3775 (N_3775,N_1442,N_167);
and U3776 (N_3776,N_2365,N_33);
and U3777 (N_3777,N_1751,N_185);
and U3778 (N_3778,N_2279,N_1150);
nand U3779 (N_3779,N_784,N_548);
or U3780 (N_3780,N_550,N_961);
or U3781 (N_3781,N_571,N_2067);
or U3782 (N_3782,N_2159,N_1905);
nand U3783 (N_3783,N_855,N_279);
or U3784 (N_3784,N_1325,N_1961);
or U3785 (N_3785,N_1093,N_2447);
nor U3786 (N_3786,N_438,N_232);
or U3787 (N_3787,N_177,N_335);
and U3788 (N_3788,N_1881,N_1785);
and U3789 (N_3789,N_2462,N_2366);
or U3790 (N_3790,N_1282,N_1837);
nand U3791 (N_3791,N_890,N_1060);
or U3792 (N_3792,N_712,N_2316);
nor U3793 (N_3793,N_1790,N_1017);
nand U3794 (N_3794,N_227,N_1240);
or U3795 (N_3795,N_319,N_0);
or U3796 (N_3796,N_1399,N_1618);
nand U3797 (N_3797,N_808,N_2062);
nand U3798 (N_3798,N_936,N_537);
and U3799 (N_3799,N_1209,N_756);
nor U3800 (N_3800,N_812,N_17);
nand U3801 (N_3801,N_795,N_1003);
and U3802 (N_3802,N_1093,N_956);
and U3803 (N_3803,N_380,N_738);
or U3804 (N_3804,N_2274,N_1173);
nor U3805 (N_3805,N_1684,N_2037);
and U3806 (N_3806,N_1596,N_1292);
nor U3807 (N_3807,N_1230,N_1627);
and U3808 (N_3808,N_166,N_807);
or U3809 (N_3809,N_620,N_333);
and U3810 (N_3810,N_1693,N_11);
and U3811 (N_3811,N_2471,N_1774);
and U3812 (N_3812,N_2322,N_1956);
nor U3813 (N_3813,N_1651,N_10);
nor U3814 (N_3814,N_433,N_1785);
and U3815 (N_3815,N_392,N_1581);
and U3816 (N_3816,N_376,N_716);
and U3817 (N_3817,N_882,N_187);
nand U3818 (N_3818,N_471,N_1163);
and U3819 (N_3819,N_261,N_1972);
nand U3820 (N_3820,N_777,N_1120);
nor U3821 (N_3821,N_238,N_580);
nor U3822 (N_3822,N_1517,N_801);
xnor U3823 (N_3823,N_1084,N_2140);
and U3824 (N_3824,N_524,N_759);
or U3825 (N_3825,N_1823,N_2146);
or U3826 (N_3826,N_1242,N_895);
nor U3827 (N_3827,N_918,N_1689);
and U3828 (N_3828,N_1683,N_709);
nand U3829 (N_3829,N_1240,N_1212);
nor U3830 (N_3830,N_2462,N_847);
and U3831 (N_3831,N_129,N_91);
nand U3832 (N_3832,N_239,N_1588);
nor U3833 (N_3833,N_1960,N_1114);
nand U3834 (N_3834,N_2296,N_614);
nand U3835 (N_3835,N_1388,N_967);
or U3836 (N_3836,N_2142,N_2449);
nand U3837 (N_3837,N_1588,N_852);
or U3838 (N_3838,N_379,N_1267);
and U3839 (N_3839,N_610,N_2015);
nor U3840 (N_3840,N_232,N_2478);
nor U3841 (N_3841,N_1908,N_879);
or U3842 (N_3842,N_433,N_1552);
or U3843 (N_3843,N_1975,N_973);
nor U3844 (N_3844,N_975,N_1116);
and U3845 (N_3845,N_2171,N_1184);
or U3846 (N_3846,N_1289,N_1328);
or U3847 (N_3847,N_2046,N_1150);
or U3848 (N_3848,N_2399,N_396);
or U3849 (N_3849,N_1725,N_447);
and U3850 (N_3850,N_629,N_1853);
xnor U3851 (N_3851,N_1566,N_1798);
nor U3852 (N_3852,N_1733,N_126);
nand U3853 (N_3853,N_1875,N_256);
and U3854 (N_3854,N_448,N_1993);
xnor U3855 (N_3855,N_1763,N_2429);
and U3856 (N_3856,N_2393,N_1108);
nand U3857 (N_3857,N_2165,N_2228);
nor U3858 (N_3858,N_2339,N_378);
or U3859 (N_3859,N_1691,N_1706);
nand U3860 (N_3860,N_26,N_1810);
nor U3861 (N_3861,N_1758,N_1381);
and U3862 (N_3862,N_1410,N_130);
or U3863 (N_3863,N_1398,N_1466);
and U3864 (N_3864,N_1615,N_1701);
nand U3865 (N_3865,N_276,N_1551);
nor U3866 (N_3866,N_2085,N_1174);
nand U3867 (N_3867,N_856,N_298);
nand U3868 (N_3868,N_2271,N_2006);
and U3869 (N_3869,N_333,N_1467);
or U3870 (N_3870,N_1848,N_678);
nand U3871 (N_3871,N_1223,N_649);
and U3872 (N_3872,N_1957,N_1782);
or U3873 (N_3873,N_574,N_822);
nor U3874 (N_3874,N_1703,N_1799);
nand U3875 (N_3875,N_2020,N_1803);
nand U3876 (N_3876,N_92,N_801);
and U3877 (N_3877,N_1861,N_1296);
and U3878 (N_3878,N_2236,N_1995);
nor U3879 (N_3879,N_2078,N_1295);
and U3880 (N_3880,N_2300,N_1573);
nor U3881 (N_3881,N_1254,N_1718);
nor U3882 (N_3882,N_1394,N_40);
nand U3883 (N_3883,N_1636,N_2130);
nand U3884 (N_3884,N_1099,N_1784);
nor U3885 (N_3885,N_1478,N_1417);
nand U3886 (N_3886,N_361,N_2048);
nand U3887 (N_3887,N_1838,N_2204);
or U3888 (N_3888,N_959,N_257);
and U3889 (N_3889,N_11,N_220);
nand U3890 (N_3890,N_1864,N_69);
nor U3891 (N_3891,N_978,N_1212);
and U3892 (N_3892,N_1913,N_1302);
nand U3893 (N_3893,N_703,N_1834);
nor U3894 (N_3894,N_1164,N_660);
nor U3895 (N_3895,N_2038,N_1037);
xor U3896 (N_3896,N_486,N_230);
or U3897 (N_3897,N_23,N_1115);
nand U3898 (N_3898,N_1724,N_1232);
nand U3899 (N_3899,N_271,N_1595);
nor U3900 (N_3900,N_2110,N_137);
and U3901 (N_3901,N_2344,N_1790);
or U3902 (N_3902,N_303,N_922);
or U3903 (N_3903,N_515,N_1497);
or U3904 (N_3904,N_655,N_1400);
nand U3905 (N_3905,N_708,N_2145);
or U3906 (N_3906,N_811,N_2236);
and U3907 (N_3907,N_2422,N_949);
or U3908 (N_3908,N_1231,N_30);
or U3909 (N_3909,N_483,N_1204);
nor U3910 (N_3910,N_185,N_2283);
nor U3911 (N_3911,N_1871,N_383);
and U3912 (N_3912,N_1973,N_1909);
and U3913 (N_3913,N_2412,N_1707);
and U3914 (N_3914,N_411,N_637);
nor U3915 (N_3915,N_1629,N_1076);
or U3916 (N_3916,N_1135,N_2189);
or U3917 (N_3917,N_1285,N_2437);
xor U3918 (N_3918,N_995,N_2453);
nand U3919 (N_3919,N_548,N_2065);
nor U3920 (N_3920,N_1492,N_1321);
nand U3921 (N_3921,N_923,N_986);
and U3922 (N_3922,N_49,N_28);
or U3923 (N_3923,N_257,N_2114);
and U3924 (N_3924,N_2276,N_146);
nor U3925 (N_3925,N_1573,N_1152);
nor U3926 (N_3926,N_26,N_720);
and U3927 (N_3927,N_2349,N_1800);
and U3928 (N_3928,N_2236,N_2216);
nor U3929 (N_3929,N_836,N_2075);
or U3930 (N_3930,N_1348,N_1457);
xnor U3931 (N_3931,N_467,N_859);
nand U3932 (N_3932,N_556,N_2035);
nor U3933 (N_3933,N_828,N_2077);
or U3934 (N_3934,N_2242,N_2250);
and U3935 (N_3935,N_2369,N_2192);
and U3936 (N_3936,N_2377,N_1336);
nand U3937 (N_3937,N_506,N_1680);
nor U3938 (N_3938,N_511,N_1236);
and U3939 (N_3939,N_2057,N_1833);
nor U3940 (N_3940,N_80,N_896);
nand U3941 (N_3941,N_2132,N_2004);
or U3942 (N_3942,N_1140,N_1063);
nand U3943 (N_3943,N_1953,N_1553);
and U3944 (N_3944,N_232,N_570);
or U3945 (N_3945,N_1964,N_1678);
nand U3946 (N_3946,N_92,N_457);
or U3947 (N_3947,N_591,N_1311);
and U3948 (N_3948,N_1302,N_2187);
and U3949 (N_3949,N_57,N_1230);
and U3950 (N_3950,N_361,N_351);
and U3951 (N_3951,N_571,N_1393);
nand U3952 (N_3952,N_2467,N_1613);
or U3953 (N_3953,N_1577,N_925);
nor U3954 (N_3954,N_43,N_1018);
or U3955 (N_3955,N_1373,N_1709);
and U3956 (N_3956,N_694,N_1071);
or U3957 (N_3957,N_39,N_1568);
or U3958 (N_3958,N_2362,N_651);
and U3959 (N_3959,N_1024,N_1759);
nor U3960 (N_3960,N_613,N_935);
and U3961 (N_3961,N_1733,N_2464);
nand U3962 (N_3962,N_1833,N_712);
nor U3963 (N_3963,N_1036,N_1901);
nand U3964 (N_3964,N_1049,N_2330);
or U3965 (N_3965,N_1752,N_1253);
nand U3966 (N_3966,N_246,N_1672);
and U3967 (N_3967,N_2119,N_1228);
nand U3968 (N_3968,N_2171,N_2461);
or U3969 (N_3969,N_452,N_2282);
and U3970 (N_3970,N_395,N_1254);
and U3971 (N_3971,N_1712,N_383);
or U3972 (N_3972,N_999,N_187);
nand U3973 (N_3973,N_237,N_528);
or U3974 (N_3974,N_1939,N_2061);
nor U3975 (N_3975,N_2375,N_321);
or U3976 (N_3976,N_2236,N_1438);
and U3977 (N_3977,N_244,N_1259);
nand U3978 (N_3978,N_1601,N_83);
nor U3979 (N_3979,N_2252,N_1901);
nor U3980 (N_3980,N_1384,N_2433);
nor U3981 (N_3981,N_87,N_2169);
nor U3982 (N_3982,N_1173,N_2121);
nand U3983 (N_3983,N_1478,N_1907);
and U3984 (N_3984,N_2086,N_116);
or U3985 (N_3985,N_2282,N_202);
nor U3986 (N_3986,N_823,N_1112);
nor U3987 (N_3987,N_1480,N_1872);
and U3988 (N_3988,N_1009,N_779);
or U3989 (N_3989,N_2363,N_505);
and U3990 (N_3990,N_263,N_1665);
and U3991 (N_3991,N_702,N_1928);
and U3992 (N_3992,N_962,N_2346);
nand U3993 (N_3993,N_2407,N_334);
nand U3994 (N_3994,N_947,N_1072);
and U3995 (N_3995,N_1890,N_2274);
or U3996 (N_3996,N_781,N_2242);
or U3997 (N_3997,N_2360,N_1482);
and U3998 (N_3998,N_1251,N_1064);
nand U3999 (N_3999,N_2157,N_2054);
nor U4000 (N_4000,N_822,N_1765);
nor U4001 (N_4001,N_1135,N_1891);
and U4002 (N_4002,N_1600,N_995);
and U4003 (N_4003,N_379,N_318);
and U4004 (N_4004,N_847,N_2388);
or U4005 (N_4005,N_250,N_1152);
and U4006 (N_4006,N_1510,N_1123);
and U4007 (N_4007,N_827,N_1755);
nand U4008 (N_4008,N_37,N_1748);
xor U4009 (N_4009,N_137,N_733);
nor U4010 (N_4010,N_278,N_269);
or U4011 (N_4011,N_56,N_1658);
nand U4012 (N_4012,N_1874,N_268);
or U4013 (N_4013,N_802,N_982);
or U4014 (N_4014,N_960,N_2106);
or U4015 (N_4015,N_353,N_1843);
or U4016 (N_4016,N_1154,N_1151);
nor U4017 (N_4017,N_503,N_1662);
or U4018 (N_4018,N_519,N_1407);
nand U4019 (N_4019,N_1509,N_1781);
nor U4020 (N_4020,N_1663,N_2402);
and U4021 (N_4021,N_524,N_2459);
nor U4022 (N_4022,N_130,N_1570);
nor U4023 (N_4023,N_276,N_1599);
and U4024 (N_4024,N_786,N_979);
and U4025 (N_4025,N_415,N_2034);
nand U4026 (N_4026,N_1291,N_982);
nand U4027 (N_4027,N_667,N_2343);
or U4028 (N_4028,N_1678,N_1314);
nor U4029 (N_4029,N_584,N_1210);
or U4030 (N_4030,N_287,N_907);
and U4031 (N_4031,N_812,N_38);
or U4032 (N_4032,N_1351,N_1639);
nand U4033 (N_4033,N_584,N_567);
nand U4034 (N_4034,N_1253,N_2324);
nand U4035 (N_4035,N_1662,N_21);
or U4036 (N_4036,N_848,N_946);
nand U4037 (N_4037,N_831,N_514);
nor U4038 (N_4038,N_620,N_1598);
or U4039 (N_4039,N_753,N_1121);
nor U4040 (N_4040,N_455,N_1532);
and U4041 (N_4041,N_62,N_162);
nand U4042 (N_4042,N_2390,N_1389);
or U4043 (N_4043,N_2064,N_490);
and U4044 (N_4044,N_2023,N_1984);
or U4045 (N_4045,N_1008,N_1000);
or U4046 (N_4046,N_1275,N_1451);
nor U4047 (N_4047,N_1354,N_705);
nor U4048 (N_4048,N_1356,N_1615);
and U4049 (N_4049,N_1099,N_1396);
nor U4050 (N_4050,N_903,N_439);
and U4051 (N_4051,N_2149,N_313);
or U4052 (N_4052,N_1497,N_477);
nand U4053 (N_4053,N_2327,N_203);
nand U4054 (N_4054,N_957,N_1006);
and U4055 (N_4055,N_1032,N_165);
or U4056 (N_4056,N_2363,N_2116);
xor U4057 (N_4057,N_1435,N_253);
or U4058 (N_4058,N_2119,N_686);
nand U4059 (N_4059,N_402,N_543);
nor U4060 (N_4060,N_1431,N_1093);
nor U4061 (N_4061,N_2302,N_1752);
and U4062 (N_4062,N_500,N_421);
or U4063 (N_4063,N_154,N_172);
xor U4064 (N_4064,N_416,N_2061);
or U4065 (N_4065,N_510,N_256);
or U4066 (N_4066,N_1424,N_1836);
or U4067 (N_4067,N_1808,N_267);
or U4068 (N_4068,N_2485,N_854);
nor U4069 (N_4069,N_1786,N_174);
nor U4070 (N_4070,N_1105,N_1776);
nor U4071 (N_4071,N_2367,N_1415);
or U4072 (N_4072,N_1920,N_1710);
nand U4073 (N_4073,N_304,N_1928);
or U4074 (N_4074,N_2430,N_496);
or U4075 (N_4075,N_447,N_1496);
or U4076 (N_4076,N_1766,N_1735);
nand U4077 (N_4077,N_1418,N_1455);
nor U4078 (N_4078,N_1752,N_832);
nand U4079 (N_4079,N_1382,N_1980);
nand U4080 (N_4080,N_2026,N_504);
nor U4081 (N_4081,N_429,N_360);
and U4082 (N_4082,N_279,N_1496);
nand U4083 (N_4083,N_1395,N_1127);
and U4084 (N_4084,N_168,N_1688);
nand U4085 (N_4085,N_339,N_2441);
nor U4086 (N_4086,N_1333,N_2194);
nand U4087 (N_4087,N_383,N_471);
nor U4088 (N_4088,N_2074,N_42);
or U4089 (N_4089,N_1518,N_1434);
or U4090 (N_4090,N_552,N_597);
and U4091 (N_4091,N_1731,N_1414);
or U4092 (N_4092,N_2085,N_685);
and U4093 (N_4093,N_1367,N_514);
nand U4094 (N_4094,N_1641,N_2059);
xnor U4095 (N_4095,N_1775,N_868);
or U4096 (N_4096,N_595,N_914);
and U4097 (N_4097,N_415,N_913);
nand U4098 (N_4098,N_1275,N_1011);
or U4099 (N_4099,N_1578,N_1726);
nand U4100 (N_4100,N_1629,N_586);
and U4101 (N_4101,N_343,N_2492);
or U4102 (N_4102,N_1288,N_867);
and U4103 (N_4103,N_891,N_1651);
or U4104 (N_4104,N_1007,N_51);
and U4105 (N_4105,N_2331,N_650);
nand U4106 (N_4106,N_826,N_819);
nand U4107 (N_4107,N_1439,N_999);
or U4108 (N_4108,N_1505,N_2453);
nor U4109 (N_4109,N_88,N_2171);
or U4110 (N_4110,N_1524,N_1136);
nor U4111 (N_4111,N_2085,N_2190);
or U4112 (N_4112,N_1288,N_483);
nand U4113 (N_4113,N_2232,N_784);
or U4114 (N_4114,N_1917,N_661);
or U4115 (N_4115,N_865,N_1428);
and U4116 (N_4116,N_1782,N_1355);
xnor U4117 (N_4117,N_825,N_1859);
xor U4118 (N_4118,N_2040,N_114);
and U4119 (N_4119,N_1634,N_708);
xor U4120 (N_4120,N_2091,N_2451);
or U4121 (N_4121,N_400,N_569);
nand U4122 (N_4122,N_798,N_886);
or U4123 (N_4123,N_385,N_2124);
and U4124 (N_4124,N_336,N_1601);
or U4125 (N_4125,N_924,N_991);
nor U4126 (N_4126,N_1172,N_581);
xor U4127 (N_4127,N_466,N_1543);
nor U4128 (N_4128,N_1516,N_1994);
nand U4129 (N_4129,N_328,N_2300);
or U4130 (N_4130,N_160,N_1839);
or U4131 (N_4131,N_2361,N_2310);
nor U4132 (N_4132,N_1385,N_792);
nor U4133 (N_4133,N_1346,N_2262);
nor U4134 (N_4134,N_787,N_1143);
and U4135 (N_4135,N_133,N_1648);
or U4136 (N_4136,N_564,N_17);
and U4137 (N_4137,N_2124,N_1940);
nor U4138 (N_4138,N_189,N_264);
or U4139 (N_4139,N_843,N_725);
nand U4140 (N_4140,N_444,N_249);
and U4141 (N_4141,N_1542,N_1437);
nand U4142 (N_4142,N_571,N_583);
nand U4143 (N_4143,N_1255,N_6);
nor U4144 (N_4144,N_1819,N_1428);
nand U4145 (N_4145,N_765,N_1340);
nor U4146 (N_4146,N_1286,N_1350);
or U4147 (N_4147,N_792,N_1115);
nor U4148 (N_4148,N_804,N_1327);
nand U4149 (N_4149,N_2425,N_1291);
or U4150 (N_4150,N_1756,N_1201);
or U4151 (N_4151,N_1171,N_311);
nand U4152 (N_4152,N_1772,N_798);
nand U4153 (N_4153,N_428,N_1374);
and U4154 (N_4154,N_2293,N_134);
nand U4155 (N_4155,N_2199,N_2149);
nor U4156 (N_4156,N_2009,N_1629);
or U4157 (N_4157,N_1366,N_617);
nand U4158 (N_4158,N_2111,N_1119);
and U4159 (N_4159,N_470,N_730);
and U4160 (N_4160,N_2158,N_2427);
or U4161 (N_4161,N_1640,N_612);
xor U4162 (N_4162,N_2057,N_1188);
and U4163 (N_4163,N_1966,N_2438);
and U4164 (N_4164,N_1224,N_1105);
or U4165 (N_4165,N_1494,N_955);
and U4166 (N_4166,N_1135,N_1390);
or U4167 (N_4167,N_2347,N_22);
nand U4168 (N_4168,N_940,N_2161);
nand U4169 (N_4169,N_611,N_2344);
or U4170 (N_4170,N_1359,N_2330);
nand U4171 (N_4171,N_1985,N_2488);
nor U4172 (N_4172,N_325,N_697);
nor U4173 (N_4173,N_68,N_1558);
and U4174 (N_4174,N_476,N_6);
or U4175 (N_4175,N_2063,N_1599);
or U4176 (N_4176,N_2442,N_2096);
nor U4177 (N_4177,N_1846,N_1445);
and U4178 (N_4178,N_1317,N_1918);
and U4179 (N_4179,N_217,N_1453);
or U4180 (N_4180,N_2214,N_458);
nor U4181 (N_4181,N_124,N_1644);
and U4182 (N_4182,N_76,N_1578);
nand U4183 (N_4183,N_2419,N_1843);
nor U4184 (N_4184,N_578,N_1668);
or U4185 (N_4185,N_1532,N_385);
nor U4186 (N_4186,N_1481,N_2488);
nor U4187 (N_4187,N_1806,N_2157);
nor U4188 (N_4188,N_1289,N_2321);
or U4189 (N_4189,N_1267,N_1824);
or U4190 (N_4190,N_1996,N_413);
and U4191 (N_4191,N_1709,N_1443);
nand U4192 (N_4192,N_201,N_2028);
nand U4193 (N_4193,N_2267,N_1279);
nor U4194 (N_4194,N_1484,N_616);
nor U4195 (N_4195,N_2284,N_637);
nand U4196 (N_4196,N_1611,N_1900);
nor U4197 (N_4197,N_2249,N_1771);
and U4198 (N_4198,N_867,N_607);
or U4199 (N_4199,N_1604,N_1083);
or U4200 (N_4200,N_1778,N_1146);
nand U4201 (N_4201,N_2070,N_22);
and U4202 (N_4202,N_1564,N_1420);
or U4203 (N_4203,N_1093,N_1066);
nand U4204 (N_4204,N_1934,N_1984);
and U4205 (N_4205,N_2076,N_1878);
and U4206 (N_4206,N_670,N_477);
nand U4207 (N_4207,N_2230,N_2441);
xnor U4208 (N_4208,N_1010,N_1806);
or U4209 (N_4209,N_1179,N_1245);
nand U4210 (N_4210,N_535,N_1829);
nor U4211 (N_4211,N_784,N_628);
nand U4212 (N_4212,N_2193,N_1465);
nand U4213 (N_4213,N_1229,N_223);
or U4214 (N_4214,N_663,N_143);
nand U4215 (N_4215,N_2088,N_383);
nand U4216 (N_4216,N_2022,N_1549);
nand U4217 (N_4217,N_54,N_2387);
and U4218 (N_4218,N_2169,N_2089);
nand U4219 (N_4219,N_2375,N_50);
nand U4220 (N_4220,N_997,N_487);
and U4221 (N_4221,N_1272,N_1183);
or U4222 (N_4222,N_824,N_1017);
nand U4223 (N_4223,N_2040,N_633);
xnor U4224 (N_4224,N_1799,N_961);
and U4225 (N_4225,N_1909,N_1071);
nor U4226 (N_4226,N_1483,N_2427);
nand U4227 (N_4227,N_709,N_1006);
nand U4228 (N_4228,N_744,N_645);
and U4229 (N_4229,N_798,N_943);
and U4230 (N_4230,N_1320,N_2091);
or U4231 (N_4231,N_1678,N_1177);
nand U4232 (N_4232,N_1138,N_984);
nand U4233 (N_4233,N_1198,N_1734);
nor U4234 (N_4234,N_2315,N_476);
nand U4235 (N_4235,N_0,N_1734);
and U4236 (N_4236,N_145,N_2419);
or U4237 (N_4237,N_1362,N_592);
nand U4238 (N_4238,N_1876,N_1701);
and U4239 (N_4239,N_1410,N_1590);
and U4240 (N_4240,N_28,N_1045);
nor U4241 (N_4241,N_128,N_164);
nand U4242 (N_4242,N_945,N_1527);
or U4243 (N_4243,N_1560,N_1113);
nand U4244 (N_4244,N_927,N_567);
or U4245 (N_4245,N_858,N_1028);
nor U4246 (N_4246,N_1628,N_2442);
nor U4247 (N_4247,N_1214,N_30);
nand U4248 (N_4248,N_1456,N_1509);
nor U4249 (N_4249,N_1729,N_1162);
or U4250 (N_4250,N_764,N_217);
nand U4251 (N_4251,N_181,N_1665);
nand U4252 (N_4252,N_1921,N_1220);
or U4253 (N_4253,N_454,N_1478);
nand U4254 (N_4254,N_1542,N_1010);
nand U4255 (N_4255,N_2040,N_1642);
nor U4256 (N_4256,N_2391,N_921);
nand U4257 (N_4257,N_2020,N_2233);
nor U4258 (N_4258,N_2499,N_1981);
and U4259 (N_4259,N_325,N_477);
xor U4260 (N_4260,N_1018,N_1508);
and U4261 (N_4261,N_1159,N_864);
and U4262 (N_4262,N_2406,N_120);
nor U4263 (N_4263,N_652,N_1009);
nor U4264 (N_4264,N_1329,N_2414);
nor U4265 (N_4265,N_1410,N_402);
nor U4266 (N_4266,N_1351,N_520);
nor U4267 (N_4267,N_2251,N_1874);
nor U4268 (N_4268,N_1026,N_2004);
and U4269 (N_4269,N_322,N_1437);
nand U4270 (N_4270,N_926,N_623);
nand U4271 (N_4271,N_1311,N_2299);
nand U4272 (N_4272,N_145,N_341);
and U4273 (N_4273,N_443,N_1483);
nand U4274 (N_4274,N_1287,N_1492);
and U4275 (N_4275,N_702,N_1665);
or U4276 (N_4276,N_836,N_355);
or U4277 (N_4277,N_2153,N_2432);
nor U4278 (N_4278,N_2130,N_650);
nand U4279 (N_4279,N_875,N_2310);
and U4280 (N_4280,N_194,N_1415);
nor U4281 (N_4281,N_1798,N_287);
nor U4282 (N_4282,N_2032,N_1819);
and U4283 (N_4283,N_1747,N_283);
nor U4284 (N_4284,N_610,N_2232);
nand U4285 (N_4285,N_55,N_1849);
and U4286 (N_4286,N_1705,N_410);
nor U4287 (N_4287,N_2367,N_1743);
nor U4288 (N_4288,N_1237,N_2474);
or U4289 (N_4289,N_1329,N_1811);
and U4290 (N_4290,N_1441,N_2277);
nor U4291 (N_4291,N_2394,N_2272);
nor U4292 (N_4292,N_560,N_1107);
nand U4293 (N_4293,N_153,N_169);
or U4294 (N_4294,N_1224,N_2218);
and U4295 (N_4295,N_1999,N_1599);
and U4296 (N_4296,N_2130,N_1095);
nand U4297 (N_4297,N_1035,N_1286);
nand U4298 (N_4298,N_1255,N_414);
nor U4299 (N_4299,N_2302,N_495);
nand U4300 (N_4300,N_59,N_443);
or U4301 (N_4301,N_2069,N_1184);
nand U4302 (N_4302,N_2164,N_1807);
and U4303 (N_4303,N_739,N_1404);
nand U4304 (N_4304,N_1494,N_2453);
xor U4305 (N_4305,N_1857,N_485);
or U4306 (N_4306,N_1712,N_1485);
nor U4307 (N_4307,N_581,N_168);
or U4308 (N_4308,N_1430,N_1977);
and U4309 (N_4309,N_96,N_2254);
and U4310 (N_4310,N_1637,N_485);
nor U4311 (N_4311,N_2100,N_417);
or U4312 (N_4312,N_1793,N_2055);
nor U4313 (N_4313,N_2245,N_2463);
nor U4314 (N_4314,N_976,N_1445);
or U4315 (N_4315,N_1608,N_1190);
and U4316 (N_4316,N_1590,N_298);
and U4317 (N_4317,N_184,N_1194);
nand U4318 (N_4318,N_74,N_1268);
and U4319 (N_4319,N_408,N_757);
or U4320 (N_4320,N_779,N_154);
and U4321 (N_4321,N_537,N_1806);
nand U4322 (N_4322,N_358,N_2354);
nand U4323 (N_4323,N_2436,N_2433);
nand U4324 (N_4324,N_682,N_482);
nand U4325 (N_4325,N_1524,N_2179);
nand U4326 (N_4326,N_1992,N_1299);
nor U4327 (N_4327,N_47,N_50);
or U4328 (N_4328,N_1778,N_434);
nand U4329 (N_4329,N_74,N_1721);
or U4330 (N_4330,N_1003,N_559);
and U4331 (N_4331,N_687,N_34);
and U4332 (N_4332,N_2014,N_2398);
nand U4333 (N_4333,N_1595,N_838);
nand U4334 (N_4334,N_737,N_1855);
and U4335 (N_4335,N_528,N_1300);
nand U4336 (N_4336,N_699,N_664);
and U4337 (N_4337,N_1467,N_952);
nand U4338 (N_4338,N_471,N_392);
xor U4339 (N_4339,N_1007,N_1350);
or U4340 (N_4340,N_66,N_770);
nand U4341 (N_4341,N_184,N_1243);
nor U4342 (N_4342,N_1933,N_1615);
nor U4343 (N_4343,N_1005,N_749);
and U4344 (N_4344,N_1529,N_339);
nor U4345 (N_4345,N_1782,N_2431);
and U4346 (N_4346,N_2250,N_1375);
and U4347 (N_4347,N_2059,N_1433);
nor U4348 (N_4348,N_1793,N_2232);
and U4349 (N_4349,N_132,N_2402);
nand U4350 (N_4350,N_723,N_987);
nor U4351 (N_4351,N_1205,N_2113);
or U4352 (N_4352,N_558,N_1553);
xnor U4353 (N_4353,N_980,N_1013);
and U4354 (N_4354,N_1285,N_2413);
or U4355 (N_4355,N_1654,N_1175);
and U4356 (N_4356,N_1081,N_748);
nor U4357 (N_4357,N_111,N_2150);
nor U4358 (N_4358,N_1416,N_2213);
or U4359 (N_4359,N_323,N_527);
nand U4360 (N_4360,N_1015,N_2420);
or U4361 (N_4361,N_1588,N_1545);
nor U4362 (N_4362,N_2150,N_570);
and U4363 (N_4363,N_1612,N_11);
or U4364 (N_4364,N_371,N_500);
and U4365 (N_4365,N_1189,N_1890);
nor U4366 (N_4366,N_60,N_962);
and U4367 (N_4367,N_945,N_427);
nand U4368 (N_4368,N_565,N_983);
nand U4369 (N_4369,N_60,N_442);
nand U4370 (N_4370,N_610,N_1777);
or U4371 (N_4371,N_2465,N_1564);
or U4372 (N_4372,N_1188,N_866);
nand U4373 (N_4373,N_557,N_1163);
nand U4374 (N_4374,N_502,N_370);
and U4375 (N_4375,N_1109,N_1069);
nand U4376 (N_4376,N_634,N_2086);
or U4377 (N_4377,N_1412,N_2079);
or U4378 (N_4378,N_1967,N_1673);
xnor U4379 (N_4379,N_1504,N_495);
and U4380 (N_4380,N_902,N_519);
or U4381 (N_4381,N_2478,N_1680);
and U4382 (N_4382,N_46,N_953);
or U4383 (N_4383,N_1518,N_2330);
nor U4384 (N_4384,N_1186,N_1819);
or U4385 (N_4385,N_542,N_2322);
nor U4386 (N_4386,N_91,N_1353);
nand U4387 (N_4387,N_1396,N_22);
nand U4388 (N_4388,N_1105,N_808);
and U4389 (N_4389,N_138,N_1651);
nor U4390 (N_4390,N_1910,N_811);
nand U4391 (N_4391,N_112,N_2462);
or U4392 (N_4392,N_113,N_511);
nand U4393 (N_4393,N_342,N_1117);
or U4394 (N_4394,N_1661,N_1223);
and U4395 (N_4395,N_2088,N_319);
and U4396 (N_4396,N_2469,N_2496);
and U4397 (N_4397,N_1985,N_1734);
and U4398 (N_4398,N_1724,N_1086);
or U4399 (N_4399,N_1119,N_1278);
or U4400 (N_4400,N_364,N_1260);
nand U4401 (N_4401,N_1960,N_149);
nor U4402 (N_4402,N_715,N_1471);
nand U4403 (N_4403,N_1234,N_1635);
nand U4404 (N_4404,N_775,N_1414);
nand U4405 (N_4405,N_212,N_469);
or U4406 (N_4406,N_613,N_1752);
nor U4407 (N_4407,N_1699,N_1850);
and U4408 (N_4408,N_311,N_2217);
or U4409 (N_4409,N_1911,N_744);
xor U4410 (N_4410,N_640,N_2304);
or U4411 (N_4411,N_728,N_77);
and U4412 (N_4412,N_360,N_2293);
nand U4413 (N_4413,N_93,N_1);
nor U4414 (N_4414,N_2441,N_989);
nor U4415 (N_4415,N_1490,N_953);
nand U4416 (N_4416,N_1152,N_2042);
nand U4417 (N_4417,N_928,N_1657);
and U4418 (N_4418,N_1608,N_2386);
nand U4419 (N_4419,N_418,N_1346);
nand U4420 (N_4420,N_762,N_1267);
nor U4421 (N_4421,N_1448,N_156);
nand U4422 (N_4422,N_2120,N_890);
nand U4423 (N_4423,N_1289,N_1306);
or U4424 (N_4424,N_36,N_1183);
and U4425 (N_4425,N_488,N_2024);
or U4426 (N_4426,N_1386,N_404);
nor U4427 (N_4427,N_402,N_291);
and U4428 (N_4428,N_164,N_1660);
and U4429 (N_4429,N_1016,N_24);
nor U4430 (N_4430,N_1526,N_2423);
or U4431 (N_4431,N_588,N_2226);
nor U4432 (N_4432,N_667,N_2036);
or U4433 (N_4433,N_961,N_589);
nor U4434 (N_4434,N_2372,N_626);
and U4435 (N_4435,N_1508,N_2219);
nand U4436 (N_4436,N_1035,N_802);
nor U4437 (N_4437,N_2277,N_351);
xor U4438 (N_4438,N_2026,N_354);
nor U4439 (N_4439,N_163,N_960);
and U4440 (N_4440,N_1842,N_1773);
nor U4441 (N_4441,N_1400,N_2334);
and U4442 (N_4442,N_1359,N_92);
and U4443 (N_4443,N_1307,N_2049);
nor U4444 (N_4444,N_95,N_3);
nor U4445 (N_4445,N_917,N_2150);
xor U4446 (N_4446,N_952,N_403);
nor U4447 (N_4447,N_1979,N_1715);
or U4448 (N_4448,N_1096,N_1597);
nor U4449 (N_4449,N_621,N_1382);
nor U4450 (N_4450,N_2054,N_1220);
or U4451 (N_4451,N_929,N_589);
nand U4452 (N_4452,N_158,N_2025);
and U4453 (N_4453,N_1174,N_2078);
and U4454 (N_4454,N_318,N_2129);
or U4455 (N_4455,N_1392,N_1417);
nor U4456 (N_4456,N_242,N_2437);
and U4457 (N_4457,N_337,N_1077);
xor U4458 (N_4458,N_800,N_821);
nor U4459 (N_4459,N_2016,N_1498);
and U4460 (N_4460,N_2403,N_1844);
nor U4461 (N_4461,N_256,N_1161);
nand U4462 (N_4462,N_587,N_2056);
xnor U4463 (N_4463,N_2447,N_964);
and U4464 (N_4464,N_106,N_1044);
or U4465 (N_4465,N_106,N_1954);
and U4466 (N_4466,N_2094,N_1367);
or U4467 (N_4467,N_427,N_1428);
or U4468 (N_4468,N_457,N_704);
or U4469 (N_4469,N_1585,N_2476);
and U4470 (N_4470,N_925,N_317);
nor U4471 (N_4471,N_1105,N_1427);
or U4472 (N_4472,N_1214,N_1301);
or U4473 (N_4473,N_359,N_1399);
or U4474 (N_4474,N_1082,N_2302);
and U4475 (N_4475,N_1487,N_960);
nor U4476 (N_4476,N_1064,N_885);
xnor U4477 (N_4477,N_321,N_1579);
or U4478 (N_4478,N_2269,N_1362);
nand U4479 (N_4479,N_983,N_615);
and U4480 (N_4480,N_2440,N_652);
and U4481 (N_4481,N_1330,N_1793);
or U4482 (N_4482,N_1055,N_558);
or U4483 (N_4483,N_722,N_2379);
xnor U4484 (N_4484,N_2021,N_446);
nor U4485 (N_4485,N_2136,N_2113);
or U4486 (N_4486,N_2353,N_756);
and U4487 (N_4487,N_637,N_1440);
nand U4488 (N_4488,N_970,N_1777);
nor U4489 (N_4489,N_1068,N_136);
nor U4490 (N_4490,N_194,N_1981);
and U4491 (N_4491,N_265,N_1567);
nor U4492 (N_4492,N_2351,N_1298);
nor U4493 (N_4493,N_1840,N_1078);
or U4494 (N_4494,N_28,N_2018);
or U4495 (N_4495,N_219,N_20);
nand U4496 (N_4496,N_1844,N_966);
nand U4497 (N_4497,N_1464,N_1873);
or U4498 (N_4498,N_1951,N_1954);
and U4499 (N_4499,N_2385,N_639);
or U4500 (N_4500,N_1794,N_504);
or U4501 (N_4501,N_1934,N_1698);
or U4502 (N_4502,N_1512,N_1036);
nand U4503 (N_4503,N_2302,N_534);
nor U4504 (N_4504,N_217,N_639);
and U4505 (N_4505,N_1051,N_1573);
nor U4506 (N_4506,N_1176,N_214);
and U4507 (N_4507,N_872,N_2391);
nand U4508 (N_4508,N_605,N_2327);
nor U4509 (N_4509,N_2372,N_1476);
nand U4510 (N_4510,N_1365,N_1227);
nor U4511 (N_4511,N_2212,N_2164);
nand U4512 (N_4512,N_638,N_728);
or U4513 (N_4513,N_848,N_1329);
nor U4514 (N_4514,N_1690,N_674);
and U4515 (N_4515,N_1489,N_121);
and U4516 (N_4516,N_1100,N_437);
and U4517 (N_4517,N_1913,N_1603);
nand U4518 (N_4518,N_1921,N_685);
or U4519 (N_4519,N_2145,N_1466);
nand U4520 (N_4520,N_2328,N_121);
nor U4521 (N_4521,N_2333,N_2424);
or U4522 (N_4522,N_1815,N_1604);
or U4523 (N_4523,N_312,N_1574);
or U4524 (N_4524,N_1896,N_134);
nor U4525 (N_4525,N_1668,N_930);
nor U4526 (N_4526,N_1139,N_837);
or U4527 (N_4527,N_2299,N_1756);
nor U4528 (N_4528,N_2348,N_985);
or U4529 (N_4529,N_647,N_2331);
nand U4530 (N_4530,N_1350,N_1576);
and U4531 (N_4531,N_2371,N_841);
and U4532 (N_4532,N_2259,N_2207);
or U4533 (N_4533,N_1919,N_1477);
nand U4534 (N_4534,N_8,N_95);
nor U4535 (N_4535,N_1733,N_778);
xnor U4536 (N_4536,N_687,N_546);
nand U4537 (N_4537,N_359,N_1213);
nor U4538 (N_4538,N_2031,N_897);
nand U4539 (N_4539,N_1639,N_1179);
nor U4540 (N_4540,N_1859,N_424);
xnor U4541 (N_4541,N_1366,N_1748);
xnor U4542 (N_4542,N_2249,N_854);
nand U4543 (N_4543,N_773,N_1694);
and U4544 (N_4544,N_1010,N_1674);
and U4545 (N_4545,N_1303,N_926);
and U4546 (N_4546,N_194,N_1768);
and U4547 (N_4547,N_815,N_676);
and U4548 (N_4548,N_2038,N_506);
nor U4549 (N_4549,N_243,N_1803);
or U4550 (N_4550,N_695,N_666);
nor U4551 (N_4551,N_472,N_1941);
or U4552 (N_4552,N_829,N_1157);
nor U4553 (N_4553,N_1920,N_1972);
or U4554 (N_4554,N_1928,N_548);
and U4555 (N_4555,N_1756,N_792);
or U4556 (N_4556,N_1773,N_636);
nand U4557 (N_4557,N_1203,N_1556);
or U4558 (N_4558,N_2020,N_1241);
or U4559 (N_4559,N_1282,N_529);
or U4560 (N_4560,N_2170,N_308);
xor U4561 (N_4561,N_802,N_2072);
nor U4562 (N_4562,N_607,N_1664);
nor U4563 (N_4563,N_998,N_2053);
nor U4564 (N_4564,N_988,N_406);
nand U4565 (N_4565,N_2003,N_2175);
nor U4566 (N_4566,N_2081,N_343);
or U4567 (N_4567,N_1870,N_1181);
and U4568 (N_4568,N_194,N_563);
nor U4569 (N_4569,N_37,N_1256);
nor U4570 (N_4570,N_54,N_2133);
and U4571 (N_4571,N_352,N_1167);
nand U4572 (N_4572,N_1781,N_1092);
and U4573 (N_4573,N_1309,N_2015);
or U4574 (N_4574,N_1919,N_130);
nor U4575 (N_4575,N_187,N_1988);
and U4576 (N_4576,N_910,N_843);
nor U4577 (N_4577,N_1843,N_1747);
nand U4578 (N_4578,N_2221,N_1974);
nor U4579 (N_4579,N_541,N_1276);
or U4580 (N_4580,N_2241,N_679);
nor U4581 (N_4581,N_1948,N_944);
or U4582 (N_4582,N_354,N_2144);
nand U4583 (N_4583,N_1949,N_2280);
and U4584 (N_4584,N_612,N_816);
nor U4585 (N_4585,N_522,N_1025);
nor U4586 (N_4586,N_622,N_2450);
nor U4587 (N_4587,N_712,N_2122);
nand U4588 (N_4588,N_890,N_479);
nor U4589 (N_4589,N_1577,N_458);
nor U4590 (N_4590,N_1191,N_825);
or U4591 (N_4591,N_1016,N_158);
and U4592 (N_4592,N_1975,N_2385);
nor U4593 (N_4593,N_1435,N_2058);
nand U4594 (N_4594,N_2414,N_805);
nand U4595 (N_4595,N_803,N_705);
or U4596 (N_4596,N_1321,N_1509);
nand U4597 (N_4597,N_1662,N_133);
nor U4598 (N_4598,N_2068,N_1667);
and U4599 (N_4599,N_2213,N_2314);
or U4600 (N_4600,N_837,N_2191);
nor U4601 (N_4601,N_412,N_1094);
and U4602 (N_4602,N_1854,N_283);
nor U4603 (N_4603,N_290,N_188);
and U4604 (N_4604,N_529,N_1951);
nor U4605 (N_4605,N_915,N_375);
nand U4606 (N_4606,N_130,N_1080);
and U4607 (N_4607,N_2162,N_250);
and U4608 (N_4608,N_1602,N_2168);
or U4609 (N_4609,N_1732,N_823);
or U4610 (N_4610,N_1572,N_329);
or U4611 (N_4611,N_2184,N_1117);
nand U4612 (N_4612,N_1394,N_90);
and U4613 (N_4613,N_361,N_1223);
nand U4614 (N_4614,N_921,N_1381);
or U4615 (N_4615,N_2356,N_1098);
or U4616 (N_4616,N_1317,N_1132);
nand U4617 (N_4617,N_466,N_1598);
nand U4618 (N_4618,N_1795,N_1607);
and U4619 (N_4619,N_1660,N_2123);
and U4620 (N_4620,N_1510,N_1057);
or U4621 (N_4621,N_856,N_1512);
nand U4622 (N_4622,N_579,N_1205);
or U4623 (N_4623,N_1774,N_1058);
and U4624 (N_4624,N_257,N_1666);
and U4625 (N_4625,N_2092,N_151);
or U4626 (N_4626,N_1555,N_2450);
nor U4627 (N_4627,N_1252,N_2307);
and U4628 (N_4628,N_1348,N_1);
xor U4629 (N_4629,N_2237,N_1832);
nor U4630 (N_4630,N_869,N_732);
or U4631 (N_4631,N_1652,N_620);
nand U4632 (N_4632,N_2248,N_2471);
or U4633 (N_4633,N_260,N_2374);
nor U4634 (N_4634,N_1864,N_1461);
or U4635 (N_4635,N_1403,N_1572);
nor U4636 (N_4636,N_1276,N_1788);
or U4637 (N_4637,N_1719,N_1522);
nor U4638 (N_4638,N_644,N_853);
nand U4639 (N_4639,N_1397,N_359);
nor U4640 (N_4640,N_500,N_908);
nand U4641 (N_4641,N_2313,N_517);
xor U4642 (N_4642,N_976,N_1662);
nand U4643 (N_4643,N_413,N_748);
and U4644 (N_4644,N_106,N_1901);
or U4645 (N_4645,N_1444,N_1596);
and U4646 (N_4646,N_297,N_2295);
nand U4647 (N_4647,N_1595,N_761);
nor U4648 (N_4648,N_433,N_117);
and U4649 (N_4649,N_2134,N_989);
nand U4650 (N_4650,N_517,N_2364);
and U4651 (N_4651,N_70,N_1820);
nand U4652 (N_4652,N_507,N_1898);
nand U4653 (N_4653,N_341,N_2207);
nand U4654 (N_4654,N_1713,N_1922);
nand U4655 (N_4655,N_1083,N_1434);
nor U4656 (N_4656,N_177,N_2016);
nor U4657 (N_4657,N_2064,N_1289);
nand U4658 (N_4658,N_1043,N_1535);
and U4659 (N_4659,N_1690,N_5);
nor U4660 (N_4660,N_580,N_1539);
nor U4661 (N_4661,N_1326,N_1649);
nor U4662 (N_4662,N_1231,N_2493);
nor U4663 (N_4663,N_549,N_330);
nand U4664 (N_4664,N_2249,N_461);
nand U4665 (N_4665,N_2127,N_1007);
and U4666 (N_4666,N_804,N_2380);
nand U4667 (N_4667,N_117,N_1083);
nor U4668 (N_4668,N_193,N_2025);
or U4669 (N_4669,N_510,N_2098);
and U4670 (N_4670,N_510,N_1272);
or U4671 (N_4671,N_2071,N_114);
xor U4672 (N_4672,N_221,N_772);
and U4673 (N_4673,N_929,N_1183);
or U4674 (N_4674,N_1074,N_997);
and U4675 (N_4675,N_1344,N_238);
nor U4676 (N_4676,N_1963,N_271);
nor U4677 (N_4677,N_303,N_606);
or U4678 (N_4678,N_751,N_776);
nand U4679 (N_4679,N_246,N_2098);
nor U4680 (N_4680,N_2294,N_85);
nand U4681 (N_4681,N_767,N_1366);
or U4682 (N_4682,N_1936,N_747);
nor U4683 (N_4683,N_2084,N_1551);
nor U4684 (N_4684,N_121,N_1006);
nand U4685 (N_4685,N_1602,N_2436);
or U4686 (N_4686,N_248,N_979);
nor U4687 (N_4687,N_610,N_1647);
nor U4688 (N_4688,N_295,N_898);
or U4689 (N_4689,N_1211,N_1932);
nand U4690 (N_4690,N_2300,N_2393);
or U4691 (N_4691,N_1206,N_2048);
nand U4692 (N_4692,N_6,N_1817);
and U4693 (N_4693,N_1829,N_936);
nand U4694 (N_4694,N_1314,N_140);
nor U4695 (N_4695,N_240,N_1403);
or U4696 (N_4696,N_23,N_620);
nor U4697 (N_4697,N_2288,N_2097);
or U4698 (N_4698,N_1589,N_1468);
nor U4699 (N_4699,N_2251,N_1482);
nor U4700 (N_4700,N_1581,N_497);
nand U4701 (N_4701,N_2034,N_583);
or U4702 (N_4702,N_1097,N_640);
nand U4703 (N_4703,N_31,N_536);
or U4704 (N_4704,N_1093,N_427);
or U4705 (N_4705,N_1123,N_1602);
or U4706 (N_4706,N_1230,N_886);
nor U4707 (N_4707,N_1740,N_2251);
and U4708 (N_4708,N_361,N_1630);
nand U4709 (N_4709,N_1743,N_1206);
nand U4710 (N_4710,N_2221,N_1362);
or U4711 (N_4711,N_965,N_2459);
nand U4712 (N_4712,N_2385,N_1014);
nor U4713 (N_4713,N_663,N_1411);
nor U4714 (N_4714,N_86,N_1281);
xor U4715 (N_4715,N_923,N_1875);
and U4716 (N_4716,N_549,N_1090);
and U4717 (N_4717,N_581,N_2244);
and U4718 (N_4718,N_832,N_1568);
or U4719 (N_4719,N_2023,N_1549);
nand U4720 (N_4720,N_1129,N_430);
nand U4721 (N_4721,N_266,N_1817);
and U4722 (N_4722,N_1412,N_2462);
nor U4723 (N_4723,N_848,N_871);
or U4724 (N_4724,N_674,N_1841);
or U4725 (N_4725,N_591,N_517);
and U4726 (N_4726,N_862,N_1061);
and U4727 (N_4727,N_1692,N_2067);
nand U4728 (N_4728,N_653,N_469);
and U4729 (N_4729,N_2131,N_605);
or U4730 (N_4730,N_1511,N_1091);
or U4731 (N_4731,N_2303,N_597);
and U4732 (N_4732,N_79,N_524);
nor U4733 (N_4733,N_1343,N_1877);
and U4734 (N_4734,N_211,N_1816);
or U4735 (N_4735,N_1869,N_208);
xnor U4736 (N_4736,N_1903,N_2129);
or U4737 (N_4737,N_2371,N_1280);
nor U4738 (N_4738,N_51,N_2060);
or U4739 (N_4739,N_932,N_148);
nand U4740 (N_4740,N_558,N_229);
nand U4741 (N_4741,N_2064,N_942);
or U4742 (N_4742,N_1656,N_467);
and U4743 (N_4743,N_679,N_1145);
nand U4744 (N_4744,N_2228,N_531);
or U4745 (N_4745,N_1289,N_53);
nand U4746 (N_4746,N_355,N_1661);
nand U4747 (N_4747,N_1985,N_1375);
or U4748 (N_4748,N_1477,N_955);
or U4749 (N_4749,N_2209,N_2018);
nand U4750 (N_4750,N_2100,N_2266);
nand U4751 (N_4751,N_2356,N_187);
and U4752 (N_4752,N_2447,N_1987);
and U4753 (N_4753,N_137,N_183);
nor U4754 (N_4754,N_65,N_1785);
nor U4755 (N_4755,N_1337,N_29);
and U4756 (N_4756,N_1190,N_1724);
nor U4757 (N_4757,N_555,N_1838);
or U4758 (N_4758,N_1329,N_771);
nor U4759 (N_4759,N_956,N_183);
and U4760 (N_4760,N_2434,N_1181);
nor U4761 (N_4761,N_1185,N_568);
and U4762 (N_4762,N_1016,N_38);
or U4763 (N_4763,N_926,N_1149);
nand U4764 (N_4764,N_900,N_611);
and U4765 (N_4765,N_985,N_1337);
nand U4766 (N_4766,N_382,N_1955);
nand U4767 (N_4767,N_733,N_316);
or U4768 (N_4768,N_2130,N_207);
and U4769 (N_4769,N_1371,N_1383);
and U4770 (N_4770,N_2299,N_1245);
and U4771 (N_4771,N_90,N_1238);
nor U4772 (N_4772,N_1074,N_1073);
nor U4773 (N_4773,N_425,N_2341);
and U4774 (N_4774,N_1378,N_706);
or U4775 (N_4775,N_2116,N_859);
or U4776 (N_4776,N_2073,N_480);
or U4777 (N_4777,N_2207,N_600);
or U4778 (N_4778,N_388,N_592);
nand U4779 (N_4779,N_736,N_1178);
nor U4780 (N_4780,N_2201,N_285);
nor U4781 (N_4781,N_1366,N_572);
and U4782 (N_4782,N_241,N_1579);
nor U4783 (N_4783,N_2240,N_2276);
nand U4784 (N_4784,N_742,N_1886);
xor U4785 (N_4785,N_1406,N_2359);
nand U4786 (N_4786,N_1320,N_1145);
or U4787 (N_4787,N_1674,N_2283);
nand U4788 (N_4788,N_1655,N_1504);
nor U4789 (N_4789,N_1791,N_572);
nor U4790 (N_4790,N_1545,N_1630);
nor U4791 (N_4791,N_1480,N_2300);
nand U4792 (N_4792,N_1763,N_726);
nor U4793 (N_4793,N_222,N_1164);
or U4794 (N_4794,N_2316,N_1932);
nand U4795 (N_4795,N_844,N_1006);
and U4796 (N_4796,N_1020,N_2323);
nand U4797 (N_4797,N_2187,N_1940);
nand U4798 (N_4798,N_1733,N_1830);
nand U4799 (N_4799,N_671,N_1974);
nand U4800 (N_4800,N_264,N_2476);
nor U4801 (N_4801,N_980,N_212);
nor U4802 (N_4802,N_1753,N_2424);
or U4803 (N_4803,N_1556,N_2462);
and U4804 (N_4804,N_765,N_831);
and U4805 (N_4805,N_1118,N_2198);
nor U4806 (N_4806,N_1242,N_1340);
nand U4807 (N_4807,N_1443,N_624);
nand U4808 (N_4808,N_1659,N_1112);
and U4809 (N_4809,N_1044,N_2472);
nor U4810 (N_4810,N_1893,N_221);
or U4811 (N_4811,N_1332,N_537);
nand U4812 (N_4812,N_546,N_2228);
nor U4813 (N_4813,N_241,N_116);
nor U4814 (N_4814,N_1782,N_876);
nor U4815 (N_4815,N_632,N_1766);
nand U4816 (N_4816,N_986,N_1013);
or U4817 (N_4817,N_827,N_172);
and U4818 (N_4818,N_1974,N_2478);
nor U4819 (N_4819,N_848,N_213);
and U4820 (N_4820,N_2057,N_2357);
nor U4821 (N_4821,N_2174,N_748);
or U4822 (N_4822,N_858,N_1112);
or U4823 (N_4823,N_1306,N_2350);
or U4824 (N_4824,N_164,N_341);
and U4825 (N_4825,N_526,N_749);
and U4826 (N_4826,N_2134,N_2226);
or U4827 (N_4827,N_315,N_821);
nand U4828 (N_4828,N_1326,N_465);
or U4829 (N_4829,N_1561,N_1673);
nor U4830 (N_4830,N_1345,N_718);
nand U4831 (N_4831,N_118,N_1236);
nor U4832 (N_4832,N_1290,N_1616);
nor U4833 (N_4833,N_1977,N_1045);
nand U4834 (N_4834,N_1985,N_2394);
nand U4835 (N_4835,N_566,N_920);
or U4836 (N_4836,N_2494,N_857);
nor U4837 (N_4837,N_2322,N_679);
or U4838 (N_4838,N_1876,N_71);
or U4839 (N_4839,N_1824,N_1552);
or U4840 (N_4840,N_332,N_2357);
nand U4841 (N_4841,N_308,N_435);
or U4842 (N_4842,N_54,N_1272);
nand U4843 (N_4843,N_2435,N_757);
nand U4844 (N_4844,N_715,N_16);
nand U4845 (N_4845,N_2361,N_2394);
nor U4846 (N_4846,N_1230,N_1580);
nor U4847 (N_4847,N_2340,N_215);
nor U4848 (N_4848,N_431,N_1722);
nor U4849 (N_4849,N_1642,N_1423);
nand U4850 (N_4850,N_249,N_1466);
or U4851 (N_4851,N_2010,N_2391);
or U4852 (N_4852,N_993,N_188);
nor U4853 (N_4853,N_2090,N_1903);
nor U4854 (N_4854,N_2208,N_1703);
or U4855 (N_4855,N_1283,N_1138);
nor U4856 (N_4856,N_155,N_1126);
nand U4857 (N_4857,N_1783,N_1884);
nand U4858 (N_4858,N_2240,N_1464);
and U4859 (N_4859,N_1325,N_1809);
nand U4860 (N_4860,N_1489,N_2273);
and U4861 (N_4861,N_646,N_1720);
or U4862 (N_4862,N_199,N_436);
or U4863 (N_4863,N_1563,N_395);
and U4864 (N_4864,N_1391,N_418);
nor U4865 (N_4865,N_2153,N_482);
nor U4866 (N_4866,N_733,N_1436);
nor U4867 (N_4867,N_1951,N_1784);
and U4868 (N_4868,N_1553,N_984);
and U4869 (N_4869,N_2356,N_1326);
and U4870 (N_4870,N_432,N_1362);
nor U4871 (N_4871,N_2030,N_2481);
nor U4872 (N_4872,N_661,N_792);
nand U4873 (N_4873,N_1805,N_1320);
and U4874 (N_4874,N_1682,N_1473);
nor U4875 (N_4875,N_577,N_1032);
xnor U4876 (N_4876,N_1486,N_1738);
nand U4877 (N_4877,N_1210,N_53);
nor U4878 (N_4878,N_1916,N_38);
nand U4879 (N_4879,N_2164,N_1191);
nand U4880 (N_4880,N_1045,N_84);
nor U4881 (N_4881,N_1064,N_1484);
nand U4882 (N_4882,N_2468,N_2430);
nor U4883 (N_4883,N_2075,N_907);
nor U4884 (N_4884,N_1159,N_1692);
or U4885 (N_4885,N_186,N_146);
nand U4886 (N_4886,N_163,N_1166);
and U4887 (N_4887,N_2499,N_267);
or U4888 (N_4888,N_1919,N_700);
nor U4889 (N_4889,N_164,N_186);
or U4890 (N_4890,N_1687,N_1845);
xnor U4891 (N_4891,N_31,N_544);
and U4892 (N_4892,N_989,N_1857);
or U4893 (N_4893,N_1212,N_1767);
nand U4894 (N_4894,N_1438,N_2341);
or U4895 (N_4895,N_739,N_1735);
and U4896 (N_4896,N_1573,N_1350);
or U4897 (N_4897,N_1109,N_1304);
and U4898 (N_4898,N_2317,N_658);
and U4899 (N_4899,N_970,N_2377);
or U4900 (N_4900,N_800,N_721);
nand U4901 (N_4901,N_1153,N_1655);
or U4902 (N_4902,N_1439,N_1217);
nand U4903 (N_4903,N_861,N_2283);
nor U4904 (N_4904,N_1487,N_2250);
nand U4905 (N_4905,N_1338,N_2144);
and U4906 (N_4906,N_1310,N_1459);
nor U4907 (N_4907,N_2474,N_1948);
and U4908 (N_4908,N_1002,N_2236);
or U4909 (N_4909,N_496,N_2253);
nor U4910 (N_4910,N_2152,N_939);
nor U4911 (N_4911,N_1619,N_185);
or U4912 (N_4912,N_81,N_831);
and U4913 (N_4913,N_272,N_174);
and U4914 (N_4914,N_1085,N_1760);
nand U4915 (N_4915,N_2201,N_1409);
nor U4916 (N_4916,N_2256,N_699);
and U4917 (N_4917,N_2473,N_1842);
xnor U4918 (N_4918,N_777,N_36);
or U4919 (N_4919,N_2453,N_1884);
or U4920 (N_4920,N_1201,N_2258);
nor U4921 (N_4921,N_2356,N_1968);
and U4922 (N_4922,N_450,N_2484);
nor U4923 (N_4923,N_1898,N_1922);
nand U4924 (N_4924,N_662,N_725);
or U4925 (N_4925,N_2151,N_2371);
and U4926 (N_4926,N_404,N_1565);
nor U4927 (N_4927,N_2136,N_364);
nand U4928 (N_4928,N_294,N_2212);
and U4929 (N_4929,N_2387,N_1721);
nor U4930 (N_4930,N_1729,N_888);
or U4931 (N_4931,N_418,N_178);
or U4932 (N_4932,N_1855,N_2221);
nor U4933 (N_4933,N_504,N_2271);
nand U4934 (N_4934,N_1506,N_1179);
xor U4935 (N_4935,N_657,N_1269);
or U4936 (N_4936,N_1656,N_1207);
nand U4937 (N_4937,N_2063,N_2116);
and U4938 (N_4938,N_60,N_2470);
or U4939 (N_4939,N_974,N_1100);
nand U4940 (N_4940,N_1820,N_503);
nor U4941 (N_4941,N_466,N_1365);
nand U4942 (N_4942,N_102,N_1169);
nor U4943 (N_4943,N_635,N_819);
nor U4944 (N_4944,N_552,N_1118);
and U4945 (N_4945,N_1810,N_1955);
xnor U4946 (N_4946,N_1405,N_1659);
or U4947 (N_4947,N_1346,N_901);
and U4948 (N_4948,N_2124,N_253);
or U4949 (N_4949,N_1072,N_19);
or U4950 (N_4950,N_817,N_191);
nor U4951 (N_4951,N_589,N_1938);
nand U4952 (N_4952,N_1825,N_1753);
nand U4953 (N_4953,N_1258,N_1316);
and U4954 (N_4954,N_1542,N_1548);
and U4955 (N_4955,N_899,N_2469);
nand U4956 (N_4956,N_1522,N_2375);
and U4957 (N_4957,N_2063,N_308);
nor U4958 (N_4958,N_1673,N_321);
or U4959 (N_4959,N_630,N_746);
xor U4960 (N_4960,N_916,N_272);
nor U4961 (N_4961,N_21,N_169);
nand U4962 (N_4962,N_1520,N_1467);
and U4963 (N_4963,N_1825,N_994);
and U4964 (N_4964,N_1455,N_1282);
nand U4965 (N_4965,N_941,N_2351);
or U4966 (N_4966,N_2153,N_1173);
and U4967 (N_4967,N_1856,N_2321);
nor U4968 (N_4968,N_598,N_1300);
nor U4969 (N_4969,N_1651,N_1345);
nor U4970 (N_4970,N_618,N_1904);
nor U4971 (N_4971,N_2114,N_1034);
nand U4972 (N_4972,N_960,N_829);
and U4973 (N_4973,N_2068,N_1140);
nor U4974 (N_4974,N_884,N_461);
and U4975 (N_4975,N_804,N_2182);
and U4976 (N_4976,N_2036,N_1464);
and U4977 (N_4977,N_2027,N_208);
nor U4978 (N_4978,N_598,N_220);
and U4979 (N_4979,N_1771,N_983);
nor U4980 (N_4980,N_2190,N_1345);
nor U4981 (N_4981,N_1047,N_695);
nor U4982 (N_4982,N_855,N_1229);
or U4983 (N_4983,N_223,N_1063);
nand U4984 (N_4984,N_1865,N_2121);
or U4985 (N_4985,N_335,N_841);
nand U4986 (N_4986,N_1434,N_922);
and U4987 (N_4987,N_1443,N_158);
and U4988 (N_4988,N_1925,N_1242);
nand U4989 (N_4989,N_2008,N_644);
or U4990 (N_4990,N_906,N_1432);
nand U4991 (N_4991,N_950,N_1418);
nand U4992 (N_4992,N_648,N_1062);
or U4993 (N_4993,N_2005,N_1840);
or U4994 (N_4994,N_1052,N_2493);
or U4995 (N_4995,N_964,N_1998);
and U4996 (N_4996,N_1308,N_872);
nor U4997 (N_4997,N_1392,N_2061);
and U4998 (N_4998,N_744,N_700);
or U4999 (N_4999,N_65,N_1465);
nand U5000 (N_5000,N_2875,N_3721);
nand U5001 (N_5001,N_3934,N_4616);
nor U5002 (N_5002,N_3677,N_4752);
nand U5003 (N_5003,N_3317,N_3318);
or U5004 (N_5004,N_4679,N_3221);
and U5005 (N_5005,N_3209,N_3158);
and U5006 (N_5006,N_4685,N_3797);
nor U5007 (N_5007,N_4795,N_4542);
and U5008 (N_5008,N_4790,N_3905);
or U5009 (N_5009,N_3357,N_4171);
xnor U5010 (N_5010,N_3524,N_4260);
or U5011 (N_5011,N_3217,N_3380);
and U5012 (N_5012,N_2718,N_4675);
nand U5013 (N_5013,N_4026,N_3965);
nand U5014 (N_5014,N_2967,N_3875);
and U5015 (N_5015,N_4534,N_3798);
and U5016 (N_5016,N_3371,N_2891);
or U5017 (N_5017,N_3345,N_4486);
nand U5018 (N_5018,N_2738,N_3398);
xor U5019 (N_5019,N_4222,N_2733);
and U5020 (N_5020,N_3803,N_2779);
or U5021 (N_5021,N_3871,N_3971);
nor U5022 (N_5022,N_3021,N_2941);
nor U5023 (N_5023,N_2926,N_4794);
and U5024 (N_5024,N_4018,N_3165);
nand U5025 (N_5025,N_3402,N_3784);
or U5026 (N_5026,N_2947,N_2839);
or U5027 (N_5027,N_3177,N_4208);
or U5028 (N_5028,N_4119,N_2677);
nand U5029 (N_5029,N_4199,N_2531);
or U5030 (N_5030,N_2678,N_3469);
or U5031 (N_5031,N_3001,N_4676);
nand U5032 (N_5032,N_4370,N_3780);
nand U5033 (N_5033,N_2573,N_4813);
nand U5034 (N_5034,N_4619,N_3920);
xnor U5035 (N_5035,N_2893,N_2707);
and U5036 (N_5036,N_3585,N_3643);
or U5037 (N_5037,N_4604,N_4766);
and U5038 (N_5038,N_3758,N_3192);
nor U5039 (N_5039,N_4281,N_2562);
nor U5040 (N_5040,N_2959,N_4832);
and U5041 (N_5041,N_4721,N_3285);
or U5042 (N_5042,N_3497,N_4310);
or U5043 (N_5043,N_3054,N_4162);
nand U5044 (N_5044,N_2513,N_2866);
nor U5045 (N_5045,N_2682,N_2584);
and U5046 (N_5046,N_2772,N_3610);
and U5047 (N_5047,N_2761,N_2582);
nor U5048 (N_5048,N_3896,N_4266);
nor U5049 (N_5049,N_4016,N_3601);
nand U5050 (N_5050,N_2897,N_4241);
or U5051 (N_5051,N_3543,N_3227);
and U5052 (N_5052,N_4423,N_4157);
nand U5053 (N_5053,N_2613,N_4382);
nand U5054 (N_5054,N_2516,N_4552);
nor U5055 (N_5055,N_2590,N_4190);
and U5056 (N_5056,N_4753,N_4818);
nor U5057 (N_5057,N_3013,N_3918);
xor U5058 (N_5058,N_3478,N_4198);
nand U5059 (N_5059,N_4618,N_4891);
nor U5060 (N_5060,N_4592,N_2679);
nand U5061 (N_5061,N_3694,N_3560);
nand U5062 (N_5062,N_3249,N_4723);
nor U5063 (N_5063,N_2924,N_4535);
xor U5064 (N_5064,N_3123,N_4060);
and U5065 (N_5065,N_3439,N_4777);
nor U5066 (N_5066,N_4906,N_3026);
and U5067 (N_5067,N_4074,N_4933);
nand U5068 (N_5068,N_2537,N_4177);
and U5069 (N_5069,N_4737,N_2871);
and U5070 (N_5070,N_3471,N_2948);
nand U5071 (N_5071,N_4204,N_2931);
nor U5072 (N_5072,N_2972,N_3949);
and U5073 (N_5073,N_4901,N_4336);
or U5074 (N_5074,N_4720,N_3805);
and U5075 (N_5075,N_2828,N_4126);
and U5076 (N_5076,N_3698,N_4910);
nor U5077 (N_5077,N_4031,N_2922);
nor U5078 (N_5078,N_3518,N_3839);
nor U5079 (N_5079,N_4206,N_2715);
or U5080 (N_5080,N_3662,N_4009);
and U5081 (N_5081,N_3552,N_4203);
or U5082 (N_5082,N_4200,N_2581);
and U5083 (N_5083,N_3384,N_3600);
or U5084 (N_5084,N_4365,N_2525);
and U5085 (N_5085,N_4975,N_4750);
nand U5086 (N_5086,N_2673,N_3173);
nand U5087 (N_5087,N_4167,N_2609);
nor U5088 (N_5088,N_2669,N_4246);
nand U5089 (N_5089,N_3831,N_2712);
and U5090 (N_5090,N_4503,N_4343);
or U5091 (N_5091,N_4335,N_3790);
or U5092 (N_5092,N_4537,N_4981);
nand U5093 (N_5093,N_4660,N_3844);
nor U5094 (N_5094,N_4913,N_4209);
nand U5095 (N_5095,N_4489,N_2874);
xor U5096 (N_5096,N_3214,N_4566);
nor U5097 (N_5097,N_2505,N_3701);
nand U5098 (N_5098,N_4925,N_4288);
nor U5099 (N_5099,N_3242,N_4547);
and U5100 (N_5100,N_4352,N_2724);
or U5101 (N_5101,N_3715,N_3187);
or U5102 (N_5102,N_4648,N_4415);
nor U5103 (N_5103,N_4828,N_2971);
or U5104 (N_5104,N_4356,N_3372);
nand U5105 (N_5105,N_4248,N_2661);
nand U5106 (N_5106,N_4887,N_4130);
or U5107 (N_5107,N_2729,N_2751);
nand U5108 (N_5108,N_4582,N_3326);
nand U5109 (N_5109,N_4888,N_3311);
nand U5110 (N_5110,N_3354,N_4414);
and U5111 (N_5111,N_4277,N_4398);
and U5112 (N_5112,N_4986,N_4220);
nand U5113 (N_5113,N_2507,N_4428);
nor U5114 (N_5114,N_3286,N_4588);
and U5115 (N_5115,N_4938,N_4946);
or U5116 (N_5116,N_2620,N_4951);
or U5117 (N_5117,N_3463,N_4181);
nand U5118 (N_5118,N_3296,N_3862);
nor U5119 (N_5119,N_3594,N_3129);
nor U5120 (N_5120,N_3073,N_2687);
nand U5121 (N_5121,N_4069,N_3699);
nand U5122 (N_5122,N_4022,N_4019);
nand U5123 (N_5123,N_4175,N_2980);
nand U5124 (N_5124,N_3647,N_4254);
and U5125 (N_5125,N_4784,N_2961);
and U5126 (N_5126,N_3529,N_3951);
nand U5127 (N_5127,N_4494,N_3162);
or U5128 (N_5128,N_4061,N_3040);
or U5129 (N_5129,N_3769,N_3144);
or U5130 (N_5130,N_3281,N_4670);
and U5131 (N_5131,N_4021,N_2618);
xnor U5132 (N_5132,N_4308,N_2994);
and U5133 (N_5133,N_4464,N_4814);
and U5134 (N_5134,N_2975,N_3327);
and U5135 (N_5135,N_4185,N_2764);
nor U5136 (N_5136,N_3995,N_2704);
nor U5137 (N_5137,N_4710,N_4435);
nand U5138 (N_5138,N_4629,N_4219);
nor U5139 (N_5139,N_4112,N_3513);
and U5140 (N_5140,N_2766,N_3825);
or U5141 (N_5141,N_3508,N_3653);
nor U5142 (N_5142,N_3917,N_4425);
xor U5143 (N_5143,N_2626,N_3736);
nor U5144 (N_5144,N_4221,N_3139);
nand U5145 (N_5145,N_4524,N_2501);
nand U5146 (N_5146,N_2737,N_3800);
nand U5147 (N_5147,N_3718,N_3312);
nor U5148 (N_5148,N_3779,N_3431);
nand U5149 (N_5149,N_3974,N_3551);
nand U5150 (N_5150,N_4633,N_3952);
nor U5151 (N_5151,N_4276,N_3846);
and U5152 (N_5152,N_4194,N_4758);
nor U5153 (N_5153,N_4475,N_4066);
nor U5154 (N_5154,N_3304,N_2752);
xor U5155 (N_5155,N_3446,N_4652);
and U5156 (N_5156,N_3858,N_4327);
or U5157 (N_5157,N_4564,N_4671);
nor U5158 (N_5158,N_2774,N_3065);
xor U5159 (N_5159,N_3946,N_4205);
nor U5160 (N_5160,N_3461,N_4450);
xor U5161 (N_5161,N_3270,N_3267);
and U5162 (N_5162,N_4517,N_4232);
and U5163 (N_5163,N_4070,N_4612);
and U5164 (N_5164,N_3941,N_3120);
nor U5165 (N_5165,N_3084,N_3929);
and U5166 (N_5166,N_2728,N_3403);
nor U5167 (N_5167,N_4767,N_4081);
nor U5168 (N_5168,N_4443,N_4824);
or U5169 (N_5169,N_3093,N_3391);
nor U5170 (N_5170,N_3206,N_3130);
nand U5171 (N_5171,N_4033,N_4040);
or U5172 (N_5172,N_2625,N_4320);
nor U5173 (N_5173,N_3178,N_3131);
and U5174 (N_5174,N_4275,N_3792);
nor U5175 (N_5175,N_4339,N_3848);
or U5176 (N_5176,N_3747,N_3525);
nor U5177 (N_5177,N_3010,N_3657);
or U5178 (N_5178,N_3392,N_2749);
or U5179 (N_5179,N_2607,N_4030);
and U5180 (N_5180,N_4837,N_4877);
and U5181 (N_5181,N_3709,N_4170);
or U5182 (N_5182,N_4110,N_4318);
or U5183 (N_5183,N_3523,N_4259);
or U5184 (N_5184,N_4734,N_4809);
nand U5185 (N_5185,N_4226,N_3869);
and U5186 (N_5186,N_2653,N_3534);
xor U5187 (N_5187,N_4374,N_3443);
nor U5188 (N_5188,N_4953,N_2527);
nand U5189 (N_5189,N_4354,N_4697);
and U5190 (N_5190,N_4563,N_3099);
nor U5191 (N_5191,N_4934,N_4937);
nand U5192 (N_5192,N_4650,N_3915);
nand U5193 (N_5193,N_4118,N_4863);
nor U5194 (N_5194,N_3587,N_4396);
and U5195 (N_5195,N_4659,N_4483);
or U5196 (N_5196,N_3583,N_4367);
or U5197 (N_5197,N_2963,N_2623);
nor U5198 (N_5198,N_4967,N_4613);
or U5199 (N_5199,N_4599,N_3269);
or U5200 (N_5200,N_3331,N_4071);
nor U5201 (N_5201,N_4635,N_3190);
and U5202 (N_5202,N_4106,N_3241);
and U5203 (N_5203,N_2646,N_2663);
nor U5204 (N_5204,N_3310,N_2713);
or U5205 (N_5205,N_3686,N_3211);
nor U5206 (N_5206,N_4032,N_2950);
and U5207 (N_5207,N_2790,N_3328);
nand U5208 (N_5208,N_2912,N_4011);
and U5209 (N_5209,N_3745,N_3731);
nand U5210 (N_5210,N_4576,N_2925);
nor U5211 (N_5211,N_3549,N_4643);
or U5212 (N_5212,N_3136,N_3503);
nand U5213 (N_5213,N_2886,N_3224);
or U5214 (N_5214,N_2927,N_3894);
nand U5215 (N_5215,N_4712,N_4843);
nand U5216 (N_5216,N_3042,N_3418);
nand U5217 (N_5217,N_3383,N_4323);
nand U5218 (N_5218,N_4319,N_3091);
nand U5219 (N_5219,N_4347,N_3368);
or U5220 (N_5220,N_2548,N_4476);
and U5221 (N_5221,N_2709,N_2879);
and U5222 (N_5222,N_3171,N_2558);
and U5223 (N_5223,N_2837,N_2601);
nand U5224 (N_5224,N_4127,N_4570);
and U5225 (N_5225,N_3015,N_3734);
or U5226 (N_5226,N_2550,N_4154);
and U5227 (N_5227,N_4731,N_2763);
or U5228 (N_5228,N_3627,N_4811);
nor U5229 (N_5229,N_4492,N_4454);
nand U5230 (N_5230,N_2638,N_2668);
or U5231 (N_5231,N_3665,N_3688);
nand U5232 (N_5232,N_4600,N_3669);
or U5233 (N_5233,N_2852,N_4682);
nor U5234 (N_5234,N_4529,N_4129);
nor U5235 (N_5235,N_2571,N_3095);
nand U5236 (N_5236,N_4780,N_3504);
nand U5237 (N_5237,N_3397,N_4405);
nor U5238 (N_5238,N_2823,N_3071);
nand U5239 (N_5239,N_4176,N_2949);
nor U5240 (N_5240,N_3955,N_4816);
or U5241 (N_5241,N_2848,N_2617);
and U5242 (N_5242,N_3739,N_3239);
or U5243 (N_5243,N_4551,N_2670);
nand U5244 (N_5244,N_4587,N_4763);
or U5245 (N_5245,N_2671,N_3544);
and U5246 (N_5246,N_3847,N_3652);
or U5247 (N_5247,N_4966,N_3763);
nor U5248 (N_5248,N_3389,N_4251);
xor U5249 (N_5249,N_4855,N_2547);
and U5250 (N_5250,N_3516,N_3893);
nand U5251 (N_5251,N_4645,N_4192);
nor U5252 (N_5252,N_2642,N_3422);
nand U5253 (N_5253,N_3633,N_4840);
or U5254 (N_5254,N_4045,N_3644);
nand U5255 (N_5255,N_3890,N_3981);
nor U5256 (N_5256,N_4460,N_2987);
and U5257 (N_5257,N_4015,N_3083);
nor U5258 (N_5258,N_3256,N_3723);
nor U5259 (N_5259,N_3004,N_4124);
and U5260 (N_5260,N_4538,N_3502);
nand U5261 (N_5261,N_4362,N_4379);
nor U5262 (N_5262,N_3057,N_3976);
nor U5263 (N_5263,N_4309,N_3023);
nand U5264 (N_5264,N_4839,N_2633);
nor U5265 (N_5265,N_3744,N_3205);
xnor U5266 (N_5266,N_4802,N_2798);
nor U5267 (N_5267,N_4351,N_2845);
nand U5268 (N_5268,N_3530,N_4369);
or U5269 (N_5269,N_3999,N_3788);
nand U5270 (N_5270,N_2589,N_2857);
and U5271 (N_5271,N_3930,N_4207);
nand U5272 (N_5272,N_4485,N_4225);
nor U5273 (N_5273,N_2794,N_3755);
and U5274 (N_5274,N_3804,N_4928);
nand U5275 (N_5275,N_2878,N_4068);
and U5276 (N_5276,N_2649,N_4702);
nand U5277 (N_5277,N_4502,N_3146);
xor U5278 (N_5278,N_3152,N_3661);
xnor U5279 (N_5279,N_4897,N_4134);
nand U5280 (N_5280,N_3902,N_4451);
nand U5281 (N_5281,N_4628,N_3204);
nand U5282 (N_5282,N_4180,N_2817);
nand U5283 (N_5283,N_3801,N_4634);
or U5284 (N_5284,N_3876,N_2596);
and U5285 (N_5285,N_4001,N_2850);
nand U5286 (N_5286,N_3808,N_3456);
nor U5287 (N_5287,N_4400,N_3385);
nand U5288 (N_5288,N_3381,N_3417);
and U5289 (N_5289,N_4950,N_4010);
xnor U5290 (N_5290,N_4885,N_3339);
nor U5291 (N_5291,N_3938,N_3977);
nand U5292 (N_5292,N_4909,N_3867);
or U5293 (N_5293,N_3433,N_3877);
nor U5294 (N_5294,N_2503,N_3903);
and U5295 (N_5295,N_4695,N_3452);
or U5296 (N_5296,N_2676,N_4466);
or U5297 (N_5297,N_4678,N_4392);
nand U5298 (N_5298,N_4699,N_4630);
and U5299 (N_5299,N_4444,N_4211);
nor U5300 (N_5300,N_3609,N_3494);
and U5301 (N_5301,N_3106,N_3793);
nand U5302 (N_5302,N_3319,N_4915);
or U5303 (N_5303,N_4807,N_3589);
nand U5304 (N_5304,N_3678,N_3488);
nand U5305 (N_5305,N_4446,N_2580);
and U5306 (N_5306,N_2627,N_4305);
or U5307 (N_5307,N_3573,N_4353);
or U5308 (N_5308,N_2714,N_3997);
or U5309 (N_5309,N_2564,N_4853);
and U5310 (N_5310,N_4247,N_4783);
nand U5311 (N_5311,N_2565,N_3415);
or U5312 (N_5312,N_4526,N_2889);
or U5313 (N_5313,N_3257,N_3637);
nand U5314 (N_5314,N_2666,N_4422);
or U5315 (N_5315,N_4801,N_3343);
and U5316 (N_5316,N_4411,N_4389);
nor U5317 (N_5317,N_4713,N_3366);
nand U5318 (N_5318,N_4043,N_4883);
nand U5319 (N_5319,N_3906,N_2781);
or U5320 (N_5320,N_3958,N_3441);
and U5321 (N_5321,N_3761,N_3216);
nand U5322 (N_5322,N_3307,N_3628);
nand U5323 (N_5323,N_3298,N_3991);
and U5324 (N_5324,N_2522,N_3008);
nor U5325 (N_5325,N_4214,N_4298);
nor U5326 (N_5326,N_4083,N_2867);
nand U5327 (N_5327,N_4755,N_3515);
nand U5328 (N_5328,N_3859,N_4439);
nand U5329 (N_5329,N_2807,N_4244);
and U5330 (N_5330,N_4920,N_2880);
or U5331 (N_5331,N_4449,N_3595);
nor U5332 (N_5332,N_3466,N_3765);
nand U5333 (N_5333,N_4546,N_2693);
and U5334 (N_5334,N_3713,N_3491);
or U5335 (N_5335,N_3922,N_4929);
nand U5336 (N_5336,N_2554,N_3776);
and U5337 (N_5337,N_4578,N_3640);
nor U5338 (N_5338,N_3449,N_4666);
and U5339 (N_5339,N_4872,N_3598);
or U5340 (N_5340,N_2825,N_3170);
nor U5341 (N_5341,N_3109,N_4997);
and U5342 (N_5342,N_4869,N_3514);
and U5343 (N_5343,N_3584,N_2914);
or U5344 (N_5344,N_4873,N_3807);
nand U5345 (N_5345,N_3649,N_4841);
and U5346 (N_5346,N_3094,N_3602);
and U5347 (N_5347,N_4402,N_4456);
nor U5348 (N_5348,N_3440,N_4468);
or U5349 (N_5349,N_4845,N_3289);
nor U5350 (N_5350,N_2719,N_3295);
or U5351 (N_5351,N_4722,N_4107);
and U5352 (N_5352,N_3287,N_4879);
nor U5353 (N_5353,N_4371,N_2619);
xnor U5354 (N_5354,N_4055,N_3953);
and U5355 (N_5355,N_3648,N_4280);
nand U5356 (N_5356,N_3673,N_2716);
xnor U5357 (N_5357,N_4430,N_2635);
or U5358 (N_5358,N_4972,N_4270);
nand U5359 (N_5359,N_3615,N_2982);
nand U5360 (N_5360,N_4686,N_4589);
or U5361 (N_5361,N_2512,N_4457);
nand U5362 (N_5362,N_2890,N_4215);
and U5363 (N_5363,N_3681,N_4467);
nor U5364 (N_5364,N_4707,N_3268);
or U5365 (N_5365,N_2998,N_4625);
and U5366 (N_5366,N_3014,N_3407);
nor U5367 (N_5367,N_2883,N_4518);
and U5368 (N_5368,N_4605,N_4315);
or U5369 (N_5369,N_3244,N_3306);
or U5370 (N_5370,N_3592,N_2705);
nor U5371 (N_5371,N_2706,N_2697);
nand U5372 (N_5372,N_3199,N_4172);
nor U5373 (N_5373,N_2520,N_3393);
nor U5374 (N_5374,N_3088,N_3016);
nand U5375 (N_5375,N_4998,N_2936);
or U5376 (N_5376,N_4677,N_4036);
and U5377 (N_5377,N_4136,N_2675);
or U5378 (N_5378,N_4156,N_4963);
and U5379 (N_5379,N_4985,N_2834);
or U5380 (N_5380,N_4386,N_2758);
nand U5381 (N_5381,N_4091,N_4532);
or U5382 (N_5382,N_4622,N_3459);
and U5383 (N_5383,N_2658,N_3253);
and U5384 (N_5384,N_4004,N_3424);
xor U5385 (N_5385,N_3540,N_3670);
or U5386 (N_5386,N_2563,N_3101);
and U5387 (N_5387,N_2602,N_2616);
and U5388 (N_5388,N_4663,N_3863);
nand U5389 (N_5389,N_3833,N_3333);
and U5390 (N_5390,N_3887,N_3025);
and U5391 (N_5391,N_3056,N_3873);
and U5392 (N_5392,N_4461,N_4146);
nor U5393 (N_5393,N_4426,N_4654);
nand U5394 (N_5394,N_3237,N_3278);
or U5395 (N_5395,N_3796,N_2829);
nor U5396 (N_5396,N_2574,N_4932);
or U5397 (N_5397,N_4996,N_2502);
nor U5398 (N_5398,N_2736,N_2545);
nor U5399 (N_5399,N_4694,N_4412);
nand U5400 (N_5400,N_3264,N_2685);
nor U5401 (N_5401,N_3785,N_4905);
nor U5402 (N_5402,N_2592,N_4867);
nor U5403 (N_5403,N_4601,N_3110);
nand U5404 (N_5404,N_4427,N_3555);
nor U5405 (N_5405,N_3507,N_2734);
nand U5406 (N_5406,N_2569,N_4372);
xor U5407 (N_5407,N_4092,N_2603);
nor U5408 (N_5408,N_4544,N_3355);
nor U5409 (N_5409,N_4990,N_2664);
or U5410 (N_5410,N_4739,N_3795);
nand U5411 (N_5411,N_3842,N_3539);
and U5412 (N_5412,N_3218,N_4864);
and U5413 (N_5413,N_3334,N_3742);
nand U5414 (N_5414,N_3302,N_4961);
nand U5415 (N_5415,N_2557,N_4930);
nor U5416 (N_5416,N_3196,N_4364);
nor U5417 (N_5417,N_4408,N_4057);
or U5418 (N_5418,N_2757,N_3632);
and U5419 (N_5419,N_4886,N_3034);
xnor U5420 (N_5420,N_3185,N_4557);
and U5421 (N_5421,N_4684,N_3987);
and U5422 (N_5422,N_2686,N_2530);
and U5423 (N_5423,N_4191,N_3251);
nand U5424 (N_5424,N_4810,N_4028);
xnor U5425 (N_5425,N_2681,N_2901);
and U5426 (N_5426,N_3064,N_3105);
nor U5427 (N_5427,N_4539,N_3119);
or U5428 (N_5428,N_4269,N_4787);
nor U5429 (N_5429,N_4980,N_3752);
or U5430 (N_5430,N_3379,N_3671);
nor U5431 (N_5431,N_4142,N_3945);
and U5432 (N_5432,N_4158,N_4960);
and U5433 (N_5433,N_3291,N_2767);
nand U5434 (N_5434,N_4812,N_3651);
or U5435 (N_5435,N_2727,N_2690);
nand U5436 (N_5436,N_3853,N_3301);
or U5437 (N_5437,N_2964,N_4095);
and U5438 (N_5438,N_3926,N_3753);
nand U5439 (N_5439,N_3201,N_4756);
nand U5440 (N_5440,N_2786,N_4447);
nor U5441 (N_5441,N_2787,N_3968);
xor U5442 (N_5442,N_3003,N_4572);
and U5443 (N_5443,N_3282,N_4703);
and U5444 (N_5444,N_4056,N_4316);
and U5445 (N_5445,N_4974,N_3031);
nand U5446 (N_5446,N_4596,N_2614);
nor U5447 (N_5447,N_3143,N_3891);
or U5448 (N_5448,N_2535,N_2858);
nor U5449 (N_5449,N_4287,N_4051);
nor U5450 (N_5450,N_3750,N_2515);
nor U5451 (N_5451,N_3435,N_2954);
or U5452 (N_5452,N_3450,N_3125);
xor U5453 (N_5453,N_3591,N_4945);
nand U5454 (N_5454,N_4614,N_3787);
nor U5455 (N_5455,N_4866,N_3045);
nand U5456 (N_5456,N_4401,N_4227);
xnor U5457 (N_5457,N_3423,N_3194);
nor U5458 (N_5458,N_2610,N_2651);
nand U5459 (N_5459,N_4341,N_3828);
nor U5460 (N_5460,N_2777,N_2659);
nand U5461 (N_5461,N_2934,N_3857);
and U5462 (N_5462,N_4132,N_3618);
nand U5463 (N_5463,N_3330,N_3654);
xor U5464 (N_5464,N_4585,N_4072);
or U5465 (N_5465,N_3998,N_3794);
nor U5466 (N_5466,N_4165,N_3954);
and U5467 (N_5467,N_3980,N_2746);
and U5468 (N_5468,N_3258,N_3566);
nand U5469 (N_5469,N_3597,N_4738);
nor U5470 (N_5470,N_4597,N_4012);
nand U5471 (N_5471,N_2815,N_3581);
nand U5472 (N_5472,N_4238,N_3658);
nand U5473 (N_5473,N_2593,N_3028);
and U5474 (N_5474,N_4152,N_3262);
nand U5475 (N_5475,N_2907,N_4970);
and U5476 (N_5476,N_4123,N_4764);
or U5477 (N_5477,N_2769,N_4102);
nor U5478 (N_5478,N_3155,N_3149);
or U5479 (N_5479,N_4264,N_4317);
nand U5480 (N_5480,N_3132,N_4926);
nor U5481 (N_5481,N_3730,N_3314);
and U5482 (N_5482,N_4006,N_4978);
or U5483 (N_5483,N_3451,N_4530);
and U5484 (N_5484,N_3541,N_3252);
nor U5485 (N_5485,N_3931,N_2629);
and U5486 (N_5486,N_3145,N_2566);
nand U5487 (N_5487,N_3829,N_4272);
nor U5488 (N_5488,N_3168,N_4984);
or U5489 (N_5489,N_4302,N_2806);
or U5490 (N_5490,N_3680,N_3770);
or U5491 (N_5491,N_3517,N_2748);
nand U5492 (N_5492,N_3348,N_3834);
nor U5493 (N_5493,N_3531,N_4893);
nand U5494 (N_5494,N_4368,N_2788);
nor U5495 (N_5495,N_3836,N_4922);
nand U5496 (N_5496,N_3043,N_4882);
and U5497 (N_5497,N_4617,N_2940);
and U5498 (N_5498,N_2645,N_4063);
or U5499 (N_5499,N_3018,N_3395);
or U5500 (N_5500,N_4672,N_3569);
xnor U5501 (N_5501,N_2585,N_4312);
or U5502 (N_5502,N_3117,N_4844);
nand U5503 (N_5503,N_4892,N_4186);
or U5504 (N_5504,N_3011,N_4573);
nand U5505 (N_5505,N_4470,N_3303);
and U5506 (N_5506,N_3975,N_3340);
and U5507 (N_5507,N_4321,N_3783);
nand U5508 (N_5508,N_2521,N_2741);
and U5509 (N_5509,N_3172,N_4042);
or U5510 (N_5510,N_2918,N_3260);
and U5511 (N_5511,N_2946,N_4894);
and U5512 (N_5512,N_4301,N_3711);
nor U5513 (N_5513,N_3039,N_4442);
nor U5514 (N_5514,N_3166,N_2538);
or U5515 (N_5515,N_3716,N_2655);
nor U5516 (N_5516,N_3772,N_4299);
and U5517 (N_5517,N_2945,N_4125);
nand U5518 (N_5518,N_2683,N_4080);
nor U5519 (N_5519,N_3990,N_3728);
nor U5520 (N_5520,N_4099,N_2775);
and U5521 (N_5521,N_4409,N_4240);
nand U5522 (N_5522,N_4291,N_4778);
nand U5523 (N_5523,N_2657,N_4669);
or U5524 (N_5524,N_3719,N_4328);
nand U5525 (N_5525,N_4609,N_3468);
nand U5526 (N_5526,N_3272,N_4329);
or U5527 (N_5527,N_2939,N_2908);
or U5528 (N_5528,N_2725,N_2588);
and U5529 (N_5529,N_4880,N_2977);
or U5530 (N_5530,N_4482,N_4500);
or U5531 (N_5531,N_4416,N_2504);
nand U5532 (N_5532,N_3630,N_4595);
nor U5533 (N_5533,N_4242,N_4512);
nand U5534 (N_5534,N_4859,N_3749);
or U5535 (N_5535,N_4122,N_3409);
or U5536 (N_5536,N_3659,N_4267);
and U5537 (N_5537,N_3376,N_4520);
or U5538 (N_5538,N_4952,N_3880);
and U5539 (N_5539,N_3979,N_4338);
nor U5540 (N_5540,N_3197,N_3683);
and U5541 (N_5541,N_4821,N_4332);
nor U5542 (N_5542,N_3883,N_3126);
nand U5543 (N_5543,N_4078,N_4413);
nand U5544 (N_5544,N_4746,N_4525);
or U5545 (N_5545,N_3870,N_3292);
nand U5546 (N_5546,N_3070,N_4748);
nand U5547 (N_5547,N_3626,N_2789);
nand U5548 (N_5548,N_4113,N_3150);
nor U5549 (N_5549,N_3436,N_4047);
or U5550 (N_5550,N_3019,N_4182);
nand U5551 (N_5551,N_4084,N_4759);
and U5552 (N_5552,N_4829,N_3243);
nand U5553 (N_5553,N_3250,N_2723);
nor U5554 (N_5554,N_4135,N_4137);
and U5555 (N_5555,N_3017,N_3851);
or U5556 (N_5556,N_4120,N_3556);
nor U5557 (N_5557,N_4765,N_4819);
or U5558 (N_5558,N_3782,N_4151);
and U5559 (N_5559,N_4825,N_3548);
nand U5560 (N_5560,N_2965,N_4732);
nor U5561 (N_5561,N_3470,N_3771);
nor U5562 (N_5562,N_4098,N_4540);
nand U5563 (N_5563,N_3215,N_2770);
nand U5564 (N_5564,N_4508,N_4927);
xnor U5565 (N_5565,N_3588,N_4257);
or U5566 (N_5566,N_3473,N_3989);
nand U5567 (N_5567,N_4727,N_4065);
or U5568 (N_5568,N_2662,N_4957);
and U5569 (N_5569,N_3811,N_2692);
and U5570 (N_5570,N_2694,N_4048);
or U5571 (N_5571,N_2768,N_2543);
and U5572 (N_5572,N_4550,N_4580);
or U5573 (N_5573,N_3090,N_3737);
nor U5574 (N_5574,N_4647,N_3888);
nand U5575 (N_5575,N_4627,N_3386);
and U5576 (N_5576,N_2630,N_3823);
nor U5577 (N_5577,N_4049,N_4311);
xnor U5578 (N_5578,N_4781,N_2559);
or U5579 (N_5579,N_3757,N_4399);
nor U5580 (N_5580,N_2855,N_4776);
and U5581 (N_5581,N_4027,N_2800);
or U5582 (N_5582,N_4943,N_3489);
nor U5583 (N_5583,N_4639,N_4698);
nor U5584 (N_5584,N_3341,N_3921);
and U5585 (N_5585,N_3210,N_4568);
nand U5586 (N_5586,N_3501,N_2604);
nor U5587 (N_5587,N_3634,N_2892);
and U5588 (N_5588,N_2608,N_2597);
nor U5589 (N_5589,N_4179,N_4002);
or U5590 (N_5590,N_2567,N_3536);
nand U5591 (N_5591,N_4278,N_2993);
or U5592 (N_5592,N_4023,N_4261);
and U5593 (N_5593,N_3561,N_4631);
and U5594 (N_5594,N_3660,N_3639);
and U5595 (N_5595,N_2762,N_4688);
and U5596 (N_5596,N_2672,N_3603);
nor U5597 (N_5597,N_2698,N_3059);
and U5598 (N_5598,N_4881,N_3820);
and U5599 (N_5599,N_3029,N_4484);
and U5600 (N_5600,N_3102,N_4788);
and U5601 (N_5601,N_3055,N_4393);
nor U5602 (N_5602,N_3604,N_2587);
or U5603 (N_5603,N_4355,N_4406);
and U5604 (N_5604,N_4473,N_2991);
or U5605 (N_5605,N_3049,N_4995);
nor U5606 (N_5606,N_4846,N_3672);
or U5607 (N_5607,N_3576,N_4487);
nor U5608 (N_5608,N_3248,N_4999);
nand U5609 (N_5609,N_3148,N_2870);
nand U5610 (N_5610,N_3041,N_4141);
nor U5611 (N_5611,N_3832,N_3323);
or U5612 (N_5612,N_4808,N_4507);
nor U5613 (N_5613,N_3474,N_4224);
and U5614 (N_5614,N_2594,N_2910);
nor U5615 (N_5615,N_2730,N_3547);
nor U5616 (N_5616,N_4861,N_4554);
nand U5617 (N_5617,N_4459,N_3193);
nor U5618 (N_5618,N_4642,N_3421);
nand U5619 (N_5619,N_4977,N_3076);
and U5620 (N_5620,N_4378,N_4912);
nand U5621 (N_5621,N_4860,N_4665);
or U5622 (N_5622,N_4144,N_4159);
or U5623 (N_5623,N_3363,N_2753);
and U5624 (N_5624,N_2591,N_4025);
xnor U5625 (N_5625,N_4424,N_4350);
nand U5626 (N_5626,N_4849,N_2843);
nor U5627 (N_5627,N_4429,N_4297);
nand U5628 (N_5628,N_3759,N_2575);
nand U5629 (N_5629,N_3611,N_3476);
and U5630 (N_5630,N_3437,N_3899);
and U5631 (N_5631,N_4848,N_3572);
or U5632 (N_5632,N_4531,N_4395);
nand U5633 (N_5633,N_4289,N_4149);
nor U5634 (N_5634,N_4711,N_4878);
nand U5635 (N_5635,N_4375,N_2920);
and U5636 (N_5636,N_4097,N_2814);
nand U5637 (N_5637,N_2953,N_4700);
or U5638 (N_5638,N_3151,N_2750);
nand U5639 (N_5639,N_2810,N_3928);
or U5640 (N_5640,N_4874,N_4662);
or U5641 (N_5641,N_2962,N_4921);
or U5642 (N_5642,N_2887,N_3308);
nor U5643 (N_5643,N_2988,N_3897);
or U5644 (N_5644,N_4363,N_2720);
or U5645 (N_5645,N_3754,N_2745);
and U5646 (N_5646,N_4761,N_3960);
or U5647 (N_5647,N_2747,N_4692);
nor U5648 (N_5648,N_4513,N_3316);
nand U5649 (N_5649,N_4094,N_3096);
or U5650 (N_5650,N_3986,N_3481);
nand U5651 (N_5651,N_4968,N_4366);
or U5652 (N_5652,N_2898,N_4575);
nand U5653 (N_5653,N_3722,N_2599);
or U5654 (N_5654,N_2583,N_2999);
and U5655 (N_5655,N_2647,N_3179);
nor U5656 (N_5656,N_4956,N_2844);
and U5657 (N_5657,N_4131,N_4150);
and U5658 (N_5658,N_4994,N_2536);
or U5659 (N_5659,N_3624,N_3147);
and U5660 (N_5660,N_2884,N_4387);
nor U5661 (N_5661,N_3137,N_3837);
nand U5662 (N_5662,N_2928,N_4850);
nor U5663 (N_5663,N_4410,N_2579);
nor U5664 (N_5664,N_4085,N_3482);
or U5665 (N_5665,N_4349,N_4252);
and U5666 (N_5666,N_3947,N_4062);
and U5667 (N_5667,N_2816,N_2882);
nor U5668 (N_5668,N_3271,N_2995);
nand U5669 (N_5669,N_3710,N_4183);
nand U5670 (N_5670,N_4046,N_4436);
nand U5671 (N_5671,N_4716,N_2578);
nand U5672 (N_5672,N_3081,N_3911);
and U5673 (N_5673,N_4751,N_4719);
and U5674 (N_5674,N_3141,N_3477);
nor U5675 (N_5675,N_4581,N_4655);
nor U5676 (N_5676,N_4948,N_3313);
nand U5677 (N_5677,N_3642,N_3985);
and U5678 (N_5678,N_2957,N_3908);
nand U5679 (N_5679,N_2944,N_2561);
or U5680 (N_5680,N_4314,N_3259);
nor U5681 (N_5681,N_3992,N_4560);
or U5682 (N_5682,N_2960,N_3212);
or U5683 (N_5683,N_3277,N_3495);
and U5684 (N_5684,N_2755,N_4117);
nor U5685 (N_5685,N_4949,N_2534);
or U5686 (N_5686,N_2933,N_3138);
xnor U5687 (N_5687,N_3612,N_4258);
xnor U5688 (N_5688,N_4733,N_3113);
or U5689 (N_5689,N_4114,N_2542);
and U5690 (N_5690,N_3100,N_4857);
and U5691 (N_5691,N_2885,N_3485);
nor U5692 (N_5692,N_3480,N_3509);
or U5693 (N_5693,N_3104,N_2811);
and U5694 (N_5694,N_3843,N_3309);
and U5695 (N_5695,N_4944,N_4555);
nand U5696 (N_5696,N_2853,N_4187);
and U5697 (N_5697,N_3963,N_4651);
nor U5698 (N_5698,N_2973,N_4743);
or U5699 (N_5699,N_4914,N_4667);
nor U5700 (N_5700,N_3786,N_2873);
nand U5701 (N_5701,N_4235,N_3593);
nand U5702 (N_5702,N_3118,N_2622);
and U5703 (N_5703,N_3505,N_4591);
nand U5704 (N_5704,N_3819,N_3726);
or U5705 (N_5705,N_4709,N_3447);
nand U5706 (N_5706,N_4624,N_2721);
nor U5707 (N_5707,N_4644,N_3086);
nand U5708 (N_5708,N_4404,N_4603);
nor U5709 (N_5709,N_3399,N_3273);
or U5710 (N_5710,N_2859,N_3464);
nor U5711 (N_5711,N_4163,N_3232);
or U5712 (N_5712,N_4865,N_4805);
or U5713 (N_5713,N_4987,N_2812);
nand U5714 (N_5714,N_3767,N_2710);
nor U5715 (N_5715,N_3520,N_4325);
or U5716 (N_5716,N_2708,N_2648);
and U5717 (N_5717,N_3571,N_2572);
and U5718 (N_5718,N_3490,N_3826);
or U5719 (N_5719,N_3982,N_3427);
nor U5720 (N_5720,N_4606,N_4223);
or U5721 (N_5721,N_3324,N_4741);
nand U5722 (N_5722,N_3886,N_3733);
nor U5723 (N_5723,N_3419,N_3578);
and U5724 (N_5724,N_3835,N_3320);
nand U5725 (N_5725,N_3635,N_4908);
and U5726 (N_5726,N_4991,N_3809);
nand U5727 (N_5727,N_2827,N_3124);
or U5728 (N_5728,N_2905,N_3280);
nand U5729 (N_5729,N_4730,N_3107);
and U5730 (N_5730,N_4931,N_4797);
and U5731 (N_5731,N_4279,N_4903);
nand U5732 (N_5732,N_4749,N_4515);
nor U5733 (N_5733,N_3284,N_2684);
and U5734 (N_5734,N_4681,N_3164);
nand U5735 (N_5735,N_4962,N_4469);
nand U5736 (N_5736,N_3866,N_4779);
nor U5737 (N_5737,N_4815,N_4621);
nand U5738 (N_5738,N_2541,N_2739);
nor U5739 (N_5739,N_3388,N_3689);
nor U5740 (N_5740,N_2689,N_3276);
or U5741 (N_5741,N_2792,N_2783);
and U5742 (N_5742,N_4044,N_4902);
nand U5743 (N_5743,N_2992,N_4488);
nand U5744 (N_5744,N_4093,N_2820);
or U5745 (N_5745,N_3619,N_3347);
or U5746 (N_5746,N_3746,N_3254);
nor U5747 (N_5747,N_3621,N_4747);
nor U5748 (N_5748,N_3493,N_3664);
nand U5749 (N_5749,N_3067,N_3983);
or U5750 (N_5750,N_4895,N_4000);
nor U5751 (N_5751,N_3050,N_3638);
and U5752 (N_5752,N_2641,N_3970);
nand U5753 (N_5753,N_2974,N_3426);
nor U5754 (N_5754,N_4969,N_3483);
nor U5755 (N_5755,N_3966,N_4197);
or U5756 (N_5756,N_4380,N_3815);
or U5757 (N_5757,N_3791,N_4109);
and U5758 (N_5758,N_2754,N_3841);
or U5759 (N_5759,N_3496,N_2702);
or U5760 (N_5760,N_3444,N_4096);
nand U5761 (N_5761,N_3768,N_4147);
nand U5762 (N_5762,N_3377,N_2722);
nor U5763 (N_5763,N_4851,N_2913);
nor U5764 (N_5764,N_2756,N_3111);
and U5765 (N_5765,N_3679,N_4029);
nand U5766 (N_5766,N_4100,N_4304);
or U5767 (N_5767,N_3641,N_3030);
or U5768 (N_5768,N_4598,N_2819);
and U5769 (N_5769,N_3226,N_3378);
nor U5770 (N_5770,N_3895,N_4620);
or U5771 (N_5771,N_4584,N_3203);
nor U5772 (N_5772,N_3373,N_3705);
nor U5773 (N_5773,N_3032,N_4611);
or U5774 (N_5774,N_4919,N_3225);
or U5775 (N_5775,N_2966,N_3623);
nor U5776 (N_5776,N_3358,N_3390);
nor U5777 (N_5777,N_3387,N_3714);
nor U5778 (N_5778,N_4827,N_3684);
and U5779 (N_5779,N_2951,N_3914);
nor U5780 (N_5780,N_4440,N_2894);
xor U5781 (N_5781,N_4303,N_2930);
xor U5782 (N_5782,N_3288,N_4104);
nor U5783 (N_5783,N_3973,N_3824);
xnor U5784 (N_5784,N_4282,N_2656);
nor U5785 (N_5785,N_4574,N_3000);
nand U5786 (N_5786,N_3527,N_3682);
nand U5787 (N_5787,N_2611,N_4623);
nor U5788 (N_5788,N_3629,N_2605);
and U5789 (N_5789,N_3020,N_2835);
and U5790 (N_5790,N_4955,N_4239);
or U5791 (N_5791,N_2628,N_3703);
or U5792 (N_5792,N_2899,N_4290);
nor U5793 (N_5793,N_4504,N_3375);
nand U5794 (N_5794,N_3036,N_3222);
nand U5795 (N_5795,N_3762,N_3830);
or U5796 (N_5796,N_4089,N_3586);
nor U5797 (N_5797,N_4657,N_4265);
and U5798 (N_5798,N_4917,N_2919);
nor U5799 (N_5799,N_4474,N_3188);
or U5800 (N_5800,N_4798,N_3557);
or U5801 (N_5801,N_3044,N_3183);
and U5802 (N_5802,N_3564,N_4330);
and U5803 (N_5803,N_4383,N_4543);
nor U5804 (N_5804,N_4431,N_3957);
nor U5805 (N_5805,N_4140,N_4195);
nor U5806 (N_5806,N_2979,N_4608);
nand U5807 (N_5807,N_3499,N_3410);
nor U5808 (N_5808,N_2860,N_4826);
nand U5809 (N_5809,N_4498,N_2586);
or U5810 (N_5810,N_2969,N_4696);
or U5811 (N_5811,N_3401,N_3511);
nand U5812 (N_5812,N_3872,N_4077);
nor U5813 (N_5813,N_4533,N_3913);
and U5814 (N_5814,N_2842,N_4506);
and U5815 (N_5815,N_4271,N_4856);
or U5816 (N_5816,N_4941,N_2923);
or U5817 (N_5817,N_4087,N_2644);
nand U5818 (N_5818,N_3936,N_2851);
and U5819 (N_5819,N_3022,N_3969);
and U5820 (N_5820,N_3616,N_4216);
nand U5821 (N_5821,N_3293,N_4740);
nor U5822 (N_5822,N_4800,N_4831);
and U5823 (N_5823,N_3806,N_4775);
nand U5824 (N_5824,N_4959,N_3338);
or U5825 (N_5825,N_3448,N_3344);
nor U5826 (N_5826,N_4823,N_3967);
and U5827 (N_5827,N_4253,N_2667);
nand U5828 (N_5828,N_3012,N_3233);
nand U5829 (N_5829,N_2808,N_2862);
nor U5830 (N_5830,N_2551,N_3599);
and U5831 (N_5831,N_3700,N_4569);
nand U5832 (N_5832,N_4237,N_2576);
nor U5833 (N_5833,N_3404,N_2981);
and U5834 (N_5834,N_4541,N_3219);
and U5835 (N_5835,N_2524,N_4876);
nor U5836 (N_5836,N_3432,N_3274);
and U5837 (N_5837,N_3724,N_3535);
nor U5838 (N_5838,N_3364,N_3087);
or U5839 (N_5839,N_4054,N_3667);
nand U5840 (N_5840,N_4556,N_4419);
nor U5841 (N_5841,N_2546,N_2632);
or U5842 (N_5842,N_2511,N_4562);
and U5843 (N_5843,N_4465,N_3396);
nor U5844 (N_5844,N_2832,N_3442);
or U5845 (N_5845,N_2881,N_3077);
nor U5846 (N_5846,N_4493,N_2553);
or U5847 (N_5847,N_4479,N_3855);
nor U5848 (N_5848,N_3693,N_4213);
and U5849 (N_5849,N_4005,N_4649);
nand U5850 (N_5850,N_3550,N_3305);
and U5851 (N_5851,N_2532,N_3741);
nand U5852 (N_5852,N_3545,N_4519);
or U5853 (N_5853,N_3840,N_3082);
nand U5854 (N_5854,N_2868,N_4417);
and U5855 (N_5855,N_4536,N_4791);
or U5856 (N_5856,N_3238,N_3625);
nor U5857 (N_5857,N_3261,N_3904);
nor U5858 (N_5858,N_3978,N_3574);
or U5859 (N_5859,N_2555,N_4637);
and U5860 (N_5860,N_3538,N_3069);
nor U5861 (N_5861,N_4148,N_3454);
nand U5862 (N_5862,N_4993,N_3717);
nor U5863 (N_5863,N_2876,N_3265);
nand U5864 (N_5864,N_4285,N_3176);
nor U5865 (N_5865,N_4835,N_3492);
xor U5866 (N_5866,N_3046,N_3901);
nand U5867 (N_5867,N_4954,N_4453);
or U5868 (N_5868,N_4717,N_3157);
or U5869 (N_5869,N_3923,N_2937);
nand U5870 (N_5870,N_3220,N_4796);
and U5871 (N_5871,N_3580,N_2833);
nor U5872 (N_5872,N_3916,N_3230);
nand U5873 (N_5873,N_4017,N_4340);
nand U5874 (N_5874,N_3361,N_2849);
xnor U5875 (N_5875,N_3245,N_4381);
nand U5876 (N_5876,N_3655,N_4153);
nor U5877 (N_5877,N_3075,N_2665);
nand U5878 (N_5878,N_4718,N_4773);
xnor U5879 (N_5879,N_4516,N_2943);
and U5880 (N_5880,N_2695,N_3153);
or U5881 (N_5881,N_4567,N_4510);
and U5882 (N_5882,N_3223,N_4725);
nand U5883 (N_5883,N_4007,N_4736);
nor U5884 (N_5884,N_4868,N_4052);
or U5885 (N_5885,N_4579,N_3738);
nor U5886 (N_5886,N_4255,N_3919);
nor U5887 (N_5887,N_3526,N_4090);
and U5888 (N_5888,N_4295,N_4348);
nor U5889 (N_5889,N_3169,N_4164);
or U5890 (N_5890,N_4742,N_4008);
nand U5891 (N_5891,N_3369,N_3329);
nor U5892 (N_5892,N_3898,N_3037);
nor U5893 (N_5893,N_3956,N_2847);
nand U5894 (N_5894,N_4230,N_2700);
or U5895 (N_5895,N_3195,N_3774);
nand U5896 (N_5896,N_4548,N_4284);
or U5897 (N_5897,N_2990,N_4769);
nand U5898 (N_5898,N_4708,N_3927);
or U5899 (N_5899,N_2539,N_3428);
nand U5900 (N_5900,N_4403,N_4434);
or U5901 (N_5901,N_4772,N_4890);
or U5902 (N_5902,N_3416,N_4690);
or U5903 (N_5903,N_4495,N_4590);
xor U5904 (N_5904,N_2711,N_4918);
and U5905 (N_5905,N_3174,N_3033);
or U5906 (N_5906,N_4073,N_3346);
and U5907 (N_5907,N_4497,N_3498);
or U5908 (N_5908,N_4210,N_3935);
and U5909 (N_5909,N_4728,N_2634);
and U5910 (N_5910,N_4345,N_3940);
or U5911 (N_5911,N_4076,N_3290);
nand U5912 (N_5912,N_3988,N_3685);
nand U5913 (N_5913,N_3676,N_4263);
and U5914 (N_5914,N_4307,N_4103);
or U5915 (N_5915,N_4610,N_2742);
nor U5916 (N_5916,N_3332,N_2514);
and U5917 (N_5917,N_3321,N_4916);
and U5918 (N_5918,N_4233,N_3706);
nor U5919 (N_5919,N_4477,N_4296);
or U5920 (N_5920,N_3563,N_4965);
and U5921 (N_5921,N_2759,N_4704);
nor U5922 (N_5922,N_3909,N_4774);
xnor U5923 (N_5923,N_4437,N_2830);
nand U5924 (N_5924,N_2916,N_4726);
and U5925 (N_5925,N_2560,N_3275);
and U5926 (N_5926,N_2598,N_4202);
xor U5927 (N_5927,N_2976,N_4294);
nor U5928 (N_5928,N_2526,N_4394);
nand U5929 (N_5929,N_2519,N_4139);
nor U5930 (N_5930,N_3707,N_4607);
nor U5931 (N_5931,N_3420,N_4691);
nor U5932 (N_5932,N_2895,N_4514);
nand U5933 (N_5933,N_2984,N_4804);
or U5934 (N_5934,N_3777,N_3300);
and U5935 (N_5935,N_3695,N_3430);
and U5936 (N_5936,N_3622,N_3114);
and U5937 (N_5937,N_4458,N_3704);
or U5938 (N_5938,N_2600,N_4421);
nand U5939 (N_5939,N_3558,N_4360);
or U5940 (N_5940,N_4664,N_2997);
nor U5941 (N_5941,N_2799,N_2533);
nor U5942 (N_5942,N_3098,N_4079);
nor U5943 (N_5943,N_3048,N_2921);
nor U5944 (N_5944,N_4357,N_4673);
or U5945 (N_5945,N_3964,N_3712);
and U5946 (N_5946,N_4138,N_2643);
or U5947 (N_5947,N_3802,N_3156);
or U5948 (N_5948,N_2688,N_4561);
or U5949 (N_5949,N_4481,N_4452);
nand U5950 (N_5950,N_3865,N_2701);
or U5951 (N_5951,N_4322,N_3532);
nand U5952 (N_5952,N_3816,N_2771);
and U5953 (N_5953,N_3325,N_4346);
nand U5954 (N_5954,N_3283,N_4822);
nor U5955 (N_5955,N_2529,N_3457);
nor U5956 (N_5956,N_2570,N_4471);
nand U5957 (N_5957,N_3479,N_4407);
nor U5958 (N_5958,N_3861,N_3115);
nor U5959 (N_5959,N_3352,N_2938);
or U5960 (N_5960,N_3053,N_3812);
nand U5961 (N_5961,N_3900,N_3608);
nand U5962 (N_5962,N_2985,N_4344);
or U5963 (N_5963,N_3646,N_4116);
and U5964 (N_5964,N_2606,N_3562);
nor U5965 (N_5965,N_3367,N_3889);
xnor U5966 (N_5966,N_3510,N_4854);
or U5967 (N_5967,N_2986,N_4646);
and U5968 (N_5968,N_2637,N_2796);
and U5969 (N_5969,N_3208,N_2773);
nor U5970 (N_5970,N_4586,N_2802);
nor U5971 (N_5971,N_2732,N_4786);
nand U5972 (N_5972,N_4377,N_3351);
xnor U5973 (N_5973,N_3154,N_4337);
nand U5974 (N_5974,N_3465,N_3687);
nor U5975 (N_5975,N_3405,N_2780);
and U5976 (N_5976,N_3134,N_2821);
or U5977 (N_5977,N_3135,N_3336);
nor U5978 (N_5978,N_3438,N_3813);
nand U5979 (N_5979,N_2776,N_3666);
or U5980 (N_5980,N_2846,N_3228);
and U5981 (N_5981,N_3060,N_2691);
and U5982 (N_5982,N_3663,N_4899);
or U5983 (N_5983,N_3720,N_3933);
and U5984 (N_5984,N_4128,N_2506);
nor U5985 (N_5985,N_4229,N_3116);
or U5986 (N_5986,N_4558,N_4274);
or U5987 (N_5987,N_4706,N_4992);
nor U5988 (N_5988,N_3537,N_4640);
or U5989 (N_5989,N_4522,N_2577);
nand U5990 (N_5990,N_3668,N_2801);
and U5991 (N_5991,N_2523,N_3849);
and U5992 (N_5992,N_4361,N_3860);
nor U5993 (N_5993,N_3236,N_2595);
and U5994 (N_5994,N_4577,N_4768);
and U5995 (N_5995,N_2989,N_3231);
nand U5996 (N_5996,N_2909,N_4923);
nor U5997 (N_5997,N_4830,N_4086);
nand U5998 (N_5998,N_3246,N_2841);
nor U5999 (N_5999,N_3937,N_2932);
nor U6000 (N_6000,N_2970,N_4896);
nand U6001 (N_6001,N_4218,N_2942);
nand U6002 (N_6002,N_3570,N_3198);
nand U6003 (N_6003,N_3590,N_2518);
or U6004 (N_6004,N_3255,N_2902);
nor U6005 (N_6005,N_4521,N_3884);
nor U6006 (N_6006,N_3943,N_4050);
or U6007 (N_6007,N_3085,N_3656);
or U6008 (N_6008,N_2784,N_2915);
or U6009 (N_6009,N_3412,N_3362);
or U6010 (N_6010,N_4034,N_3159);
nand U6011 (N_6011,N_3063,N_4661);
nor U6012 (N_6012,N_4760,N_4088);
nor U6013 (N_6013,N_3506,N_3696);
or U6014 (N_6014,N_4039,N_2822);
or U6015 (N_6015,N_4653,N_2760);
xnor U6016 (N_6016,N_2805,N_3006);
or U6017 (N_6017,N_4632,N_3727);
and U6018 (N_6018,N_4523,N_3360);
nand U6019 (N_6019,N_4256,N_4593);
nand U6020 (N_6020,N_4803,N_2838);
nor U6021 (N_6021,N_2636,N_4433);
or U6022 (N_6022,N_2650,N_3486);
nor U6023 (N_6023,N_4594,N_3462);
or U6024 (N_6024,N_3577,N_2955);
nand U6025 (N_6025,N_2652,N_3910);
nand U6026 (N_6026,N_4196,N_4490);
nand U6027 (N_6027,N_4884,N_4940);
or U6028 (N_6028,N_2958,N_3521);
and U6029 (N_6029,N_3133,N_3925);
nand U6030 (N_6030,N_2865,N_3279);
and U6031 (N_6031,N_4715,N_3778);
or U6032 (N_6032,N_2699,N_4907);
and U6033 (N_6033,N_3939,N_2797);
or U6034 (N_6034,N_3163,N_3455);
nand U6035 (N_6035,N_4833,N_4324);
nand U6036 (N_6036,N_2911,N_3263);
and U6037 (N_6037,N_2888,N_4858);
nor U6038 (N_6038,N_3868,N_2813);
and U6039 (N_6039,N_4236,N_4982);
and U6040 (N_6040,N_2615,N_3961);
nand U6041 (N_6041,N_3487,N_3702);
or U6042 (N_6042,N_4971,N_4168);
and U6043 (N_6043,N_4331,N_4989);
and U6044 (N_6044,N_4898,N_4376);
nand U6045 (N_6045,N_3200,N_4680);
nor U6046 (N_6046,N_4782,N_4771);
nor U6047 (N_6047,N_4480,N_3414);
and U6048 (N_6048,N_4059,N_3007);
and U6049 (N_6049,N_3756,N_3575);
nor U6050 (N_6050,N_2624,N_4418);
or U6051 (N_6051,N_3675,N_3697);
or U6052 (N_6052,N_3864,N_2778);
or U6053 (N_6053,N_3103,N_2791);
nand U6054 (N_6054,N_3614,N_4491);
or U6055 (N_6055,N_3691,N_3072);
and U6056 (N_6056,N_3122,N_4432);
nand U6057 (N_6057,N_2896,N_4626);
nand U6058 (N_6058,N_2740,N_3553);
and U6059 (N_6059,N_3472,N_3350);
or U6060 (N_6060,N_2840,N_3356);
nor U6061 (N_6061,N_4834,N_3892);
nor U6062 (N_6062,N_3406,N_4754);
or U6063 (N_6063,N_3740,N_2540);
nor U6064 (N_6064,N_4283,N_3005);
xor U6065 (N_6065,N_4463,N_3546);
nor U6066 (N_6066,N_4326,N_3349);
and U6067 (N_6067,N_3948,N_4744);
nor U6068 (N_6068,N_3708,N_4174);
nand U6069 (N_6069,N_4445,N_3674);
nand U6070 (N_6070,N_3429,N_4184);
nand U6071 (N_6071,N_4478,N_2568);
or U6072 (N_6072,N_4014,N_3374);
or U6073 (N_6073,N_3370,N_4583);
and U6074 (N_6074,N_3266,N_4333);
and U6075 (N_6075,N_4973,N_3743);
nand U6076 (N_6076,N_2556,N_4602);
or U6077 (N_6077,N_2864,N_4817);
nor U6078 (N_6078,N_4705,N_4115);
nor U6079 (N_6079,N_2824,N_4785);
or U6080 (N_6080,N_3690,N_3142);
or U6081 (N_6081,N_4875,N_4842);
xnor U6082 (N_6082,N_2836,N_2903);
nand U6083 (N_6083,N_3038,N_2904);
nor U6084 (N_6084,N_3213,N_2782);
and U6085 (N_6085,N_3078,N_4939);
and U6086 (N_6086,N_3554,N_2869);
nand U6087 (N_6087,N_2906,N_3567);
and U6088 (N_6088,N_3962,N_3775);
nor U6089 (N_6089,N_4108,N_4334);
or U6090 (N_6090,N_3822,N_3160);
nand U6091 (N_6091,N_4687,N_4976);
xor U6092 (N_6092,N_3191,N_3885);
and U6093 (N_6093,N_4234,N_4441);
and U6094 (N_6094,N_3062,N_2660);
or U6095 (N_6095,N_3827,N_3342);
and U6096 (N_6096,N_2517,N_3189);
nand U6097 (N_6097,N_3400,N_3460);
or U6098 (N_6098,N_3207,N_4789);
or U6099 (N_6099,N_2793,N_3852);
xor U6100 (N_6100,N_4496,N_2809);
or U6101 (N_6101,N_3315,N_3051);
nand U6102 (N_6102,N_2803,N_3732);
nor U6103 (N_6103,N_4836,N_4499);
or U6104 (N_6104,N_2500,N_3789);
nand U6105 (N_6105,N_3458,N_4820);
nand U6106 (N_6106,N_4397,N_3850);
nand U6107 (N_6107,N_3924,N_3984);
nand U6108 (N_6108,N_4035,N_3047);
or U6109 (N_6109,N_4770,N_4188);
nor U6110 (N_6110,N_4762,N_3365);
nand U6111 (N_6111,N_4075,N_4792);
nand U6112 (N_6112,N_2917,N_4193);
and U6113 (N_6113,N_3097,N_4041);
nand U6114 (N_6114,N_3127,N_3613);
nand U6115 (N_6115,N_4924,N_3579);
and U6116 (N_6116,N_2640,N_4656);
nor U6117 (N_6117,N_3821,N_4058);
or U6118 (N_6118,N_3484,N_4438);
and U6119 (N_6119,N_3878,N_4472);
nand U6120 (N_6120,N_3636,N_3180);
nand U6121 (N_6121,N_4155,N_4388);
nor U6122 (N_6122,N_3235,N_2612);
nand U6123 (N_6123,N_3559,N_4173);
or U6124 (N_6124,N_2654,N_3519);
or U6125 (N_6125,N_3607,N_3692);
and U6126 (N_6126,N_2978,N_4683);
or U6127 (N_6127,N_4020,N_4105);
or U6128 (N_6128,N_2631,N_2639);
nor U6129 (N_6129,N_4243,N_4509);
nand U6130 (N_6130,N_3182,N_3735);
or U6131 (N_6131,N_3512,N_4935);
nor U6132 (N_6132,N_4641,N_3766);
and U6133 (N_6133,N_2863,N_2983);
xor U6134 (N_6134,N_4228,N_4160);
and U6135 (N_6135,N_4714,N_3751);
and U6136 (N_6136,N_4358,N_2735);
and U6137 (N_6137,N_2968,N_4724);
and U6138 (N_6138,N_3932,N_2528);
and U6139 (N_6139,N_3434,N_3027);
nand U6140 (N_6140,N_3202,N_4390);
and U6141 (N_6141,N_4212,N_2935);
and U6142 (N_6142,N_2731,N_3838);
or U6143 (N_6143,N_2549,N_4306);
nor U6144 (N_6144,N_3337,N_3773);
or U6145 (N_6145,N_4615,N_3856);
nor U6146 (N_6146,N_4101,N_3631);
nor U6147 (N_6147,N_3817,N_4693);
and U6148 (N_6148,N_4505,N_4947);
nor U6149 (N_6149,N_2680,N_3760);
or U6150 (N_6150,N_3606,N_2744);
nand U6151 (N_6151,N_4638,N_4964);
or U6152 (N_6152,N_3061,N_3229);
or U6153 (N_6153,N_4359,N_4250);
or U6154 (N_6154,N_3413,N_3140);
nor U6155 (N_6155,N_4024,N_3079);
and U6156 (N_6156,N_3112,N_3950);
and U6157 (N_6157,N_4145,N_2956);
and U6158 (N_6158,N_4038,N_3972);
nand U6159 (N_6159,N_4286,N_4385);
and U6160 (N_6160,N_4689,N_3912);
nor U6161 (N_6161,N_4658,N_3066);
or U6162 (N_6162,N_4003,N_4313);
nor U6163 (N_6163,N_4862,N_3565);
nand U6164 (N_6164,N_3058,N_2621);
or U6165 (N_6165,N_3582,N_4300);
nor U6166 (N_6166,N_4201,N_3528);
or U6167 (N_6167,N_3240,N_3394);
nor U6168 (N_6168,N_3186,N_4942);
and U6169 (N_6169,N_3128,N_3002);
or U6170 (N_6170,N_4889,N_4082);
nand U6171 (N_6171,N_4373,N_3074);
nand U6172 (N_6172,N_4979,N_3297);
nand U6173 (N_6173,N_2900,N_2952);
and U6174 (N_6174,N_3052,N_2674);
nor U6175 (N_6175,N_4293,N_3382);
and U6176 (N_6176,N_2552,N_3814);
xnor U6177 (N_6177,N_3764,N_3645);
and U6178 (N_6178,N_2508,N_3996);
nand U6179 (N_6179,N_3854,N_4121);
or U6180 (N_6180,N_4268,N_4262);
or U6181 (N_6181,N_4462,N_4983);
nand U6182 (N_6182,N_3748,N_4871);
nor U6183 (N_6183,N_3108,N_3445);
and U6184 (N_6184,N_3167,N_4384);
or U6185 (N_6185,N_4342,N_4852);
nand U6186 (N_6186,N_4870,N_4189);
or U6187 (N_6187,N_4838,N_4013);
or U6188 (N_6188,N_3907,N_2717);
and U6189 (N_6189,N_3799,N_2544);
nand U6190 (N_6190,N_4161,N_3092);
and U6191 (N_6191,N_3818,N_4729);
or U6192 (N_6192,N_3080,N_3845);
and U6193 (N_6193,N_3522,N_3959);
or U6194 (N_6194,N_4806,N_3944);
nand U6195 (N_6195,N_3617,N_4904);
nor U6196 (N_6196,N_2510,N_3810);
or U6197 (N_6197,N_4900,N_2818);
xnor U6198 (N_6198,N_3620,N_3879);
nor U6199 (N_6199,N_4911,N_3353);
nor U6200 (N_6200,N_4217,N_4037);
nor U6201 (N_6201,N_3121,N_4169);
and U6202 (N_6202,N_2696,N_4936);
and U6203 (N_6203,N_3568,N_3596);
or U6204 (N_6204,N_4143,N_4745);
nor U6205 (N_6205,N_3533,N_3994);
nor U6206 (N_6206,N_3475,N_3359);
and U6207 (N_6207,N_3605,N_4571);
nor U6208 (N_6208,N_4527,N_3181);
or U6209 (N_6209,N_2804,N_4292);
nand U6210 (N_6210,N_4559,N_4455);
nor U6211 (N_6211,N_2703,N_3068);
or U6212 (N_6212,N_3781,N_4545);
nand U6213 (N_6213,N_2831,N_4668);
xnor U6214 (N_6214,N_3942,N_4549);
nand U6215 (N_6215,N_2856,N_4273);
or U6216 (N_6216,N_3247,N_3500);
or U6217 (N_6217,N_4178,N_4636);
nor U6218 (N_6218,N_3024,N_2785);
nor U6219 (N_6219,N_4528,N_4958);
and U6220 (N_6220,N_4166,N_2872);
nor U6221 (N_6221,N_2726,N_4674);
or U6222 (N_6222,N_4847,N_3035);
nor U6223 (N_6223,N_2996,N_3729);
and U6224 (N_6224,N_3411,N_2765);
or U6225 (N_6225,N_3993,N_4448);
or U6226 (N_6226,N_4799,N_3089);
nand U6227 (N_6227,N_3408,N_3725);
nor U6228 (N_6228,N_4053,N_4701);
or U6229 (N_6229,N_3184,N_3294);
nand U6230 (N_6230,N_4231,N_3467);
and U6231 (N_6231,N_4064,N_3882);
or U6232 (N_6232,N_2877,N_4735);
or U6233 (N_6233,N_3425,N_4511);
nand U6234 (N_6234,N_3453,N_3161);
nand U6235 (N_6235,N_3322,N_3881);
nor U6236 (N_6236,N_4111,N_4249);
nand U6237 (N_6237,N_4067,N_4757);
nand U6238 (N_6238,N_2743,N_2861);
nor U6239 (N_6239,N_3542,N_3874);
nand U6240 (N_6240,N_4391,N_4501);
or U6241 (N_6241,N_3650,N_3299);
or U6242 (N_6242,N_3234,N_2826);
nand U6243 (N_6243,N_2929,N_2854);
and U6244 (N_6244,N_2509,N_4245);
or U6245 (N_6245,N_4420,N_3009);
or U6246 (N_6246,N_3335,N_4133);
and U6247 (N_6247,N_4553,N_2795);
xor U6248 (N_6248,N_4565,N_3175);
or U6249 (N_6249,N_4793,N_4988);
xor U6250 (N_6250,N_3219,N_4796);
or U6251 (N_6251,N_3446,N_3622);
and U6252 (N_6252,N_2984,N_2758);
nor U6253 (N_6253,N_3516,N_3258);
and U6254 (N_6254,N_4270,N_2711);
nand U6255 (N_6255,N_3809,N_3142);
and U6256 (N_6256,N_2590,N_4853);
nor U6257 (N_6257,N_4045,N_3645);
nor U6258 (N_6258,N_4772,N_3797);
and U6259 (N_6259,N_4062,N_3611);
and U6260 (N_6260,N_3657,N_2536);
nand U6261 (N_6261,N_4689,N_4724);
and U6262 (N_6262,N_3453,N_3838);
or U6263 (N_6263,N_4003,N_3845);
or U6264 (N_6264,N_2577,N_3055);
nor U6265 (N_6265,N_2728,N_4373);
nor U6266 (N_6266,N_3775,N_2747);
xor U6267 (N_6267,N_4051,N_4200);
nor U6268 (N_6268,N_3475,N_4066);
nor U6269 (N_6269,N_3764,N_2593);
nand U6270 (N_6270,N_3819,N_4158);
nand U6271 (N_6271,N_3268,N_3044);
nand U6272 (N_6272,N_2950,N_4885);
nor U6273 (N_6273,N_4563,N_3963);
nand U6274 (N_6274,N_3619,N_3595);
and U6275 (N_6275,N_3367,N_3829);
nor U6276 (N_6276,N_3644,N_4478);
nand U6277 (N_6277,N_3347,N_4165);
or U6278 (N_6278,N_4564,N_3124);
nor U6279 (N_6279,N_4385,N_4085);
nor U6280 (N_6280,N_3992,N_4492);
or U6281 (N_6281,N_4904,N_3689);
and U6282 (N_6282,N_4742,N_3440);
and U6283 (N_6283,N_4283,N_4732);
nor U6284 (N_6284,N_3833,N_3636);
and U6285 (N_6285,N_3371,N_3822);
xnor U6286 (N_6286,N_2745,N_3995);
nor U6287 (N_6287,N_3569,N_4915);
nor U6288 (N_6288,N_3602,N_4672);
nand U6289 (N_6289,N_3791,N_4722);
nor U6290 (N_6290,N_3547,N_3869);
nand U6291 (N_6291,N_3938,N_4136);
nand U6292 (N_6292,N_2671,N_4342);
xnor U6293 (N_6293,N_3280,N_2589);
and U6294 (N_6294,N_4142,N_2762);
nor U6295 (N_6295,N_2640,N_3851);
or U6296 (N_6296,N_3597,N_3632);
nor U6297 (N_6297,N_2782,N_3442);
nor U6298 (N_6298,N_3209,N_3808);
nor U6299 (N_6299,N_4837,N_3954);
and U6300 (N_6300,N_3169,N_3351);
nor U6301 (N_6301,N_3715,N_4027);
and U6302 (N_6302,N_4199,N_3117);
nand U6303 (N_6303,N_3835,N_3066);
nor U6304 (N_6304,N_3346,N_2641);
nor U6305 (N_6305,N_4994,N_3158);
nor U6306 (N_6306,N_3702,N_4327);
nor U6307 (N_6307,N_2795,N_3345);
and U6308 (N_6308,N_2876,N_4721);
or U6309 (N_6309,N_3321,N_3252);
nor U6310 (N_6310,N_4814,N_2728);
nor U6311 (N_6311,N_4874,N_4213);
or U6312 (N_6312,N_2868,N_3603);
or U6313 (N_6313,N_3158,N_2794);
and U6314 (N_6314,N_3963,N_3221);
nand U6315 (N_6315,N_4983,N_4211);
nor U6316 (N_6316,N_4221,N_4974);
xnor U6317 (N_6317,N_2821,N_2853);
nand U6318 (N_6318,N_4231,N_4991);
nand U6319 (N_6319,N_4694,N_4602);
nor U6320 (N_6320,N_3048,N_2606);
nor U6321 (N_6321,N_4623,N_3433);
and U6322 (N_6322,N_4265,N_3614);
or U6323 (N_6323,N_3176,N_2877);
and U6324 (N_6324,N_2528,N_3255);
nand U6325 (N_6325,N_2696,N_4080);
or U6326 (N_6326,N_4240,N_4280);
nand U6327 (N_6327,N_3792,N_3377);
or U6328 (N_6328,N_4364,N_4802);
and U6329 (N_6329,N_4454,N_2658);
and U6330 (N_6330,N_2977,N_4135);
or U6331 (N_6331,N_2621,N_3067);
or U6332 (N_6332,N_4808,N_4513);
xor U6333 (N_6333,N_4749,N_3720);
nor U6334 (N_6334,N_4624,N_2796);
nor U6335 (N_6335,N_2729,N_2867);
nand U6336 (N_6336,N_2534,N_4198);
nand U6337 (N_6337,N_4150,N_3474);
and U6338 (N_6338,N_4153,N_3446);
nor U6339 (N_6339,N_4853,N_3214);
nand U6340 (N_6340,N_3808,N_2991);
nand U6341 (N_6341,N_4240,N_3883);
or U6342 (N_6342,N_3060,N_3941);
nand U6343 (N_6343,N_3655,N_4240);
nor U6344 (N_6344,N_4795,N_2641);
or U6345 (N_6345,N_2578,N_3745);
or U6346 (N_6346,N_4913,N_3757);
nor U6347 (N_6347,N_4325,N_4583);
nand U6348 (N_6348,N_3745,N_3039);
and U6349 (N_6349,N_4515,N_3249);
or U6350 (N_6350,N_2816,N_2718);
xnor U6351 (N_6351,N_4670,N_3326);
nor U6352 (N_6352,N_3970,N_3109);
and U6353 (N_6353,N_3531,N_4821);
nor U6354 (N_6354,N_3316,N_4520);
and U6355 (N_6355,N_3045,N_4347);
xor U6356 (N_6356,N_2841,N_2566);
or U6357 (N_6357,N_4401,N_2986);
nor U6358 (N_6358,N_2638,N_4819);
and U6359 (N_6359,N_4956,N_3278);
and U6360 (N_6360,N_3114,N_2840);
xor U6361 (N_6361,N_3773,N_3919);
nand U6362 (N_6362,N_3408,N_4911);
nor U6363 (N_6363,N_3943,N_2787);
nand U6364 (N_6364,N_2664,N_3171);
and U6365 (N_6365,N_3799,N_3379);
and U6366 (N_6366,N_3149,N_2623);
and U6367 (N_6367,N_4884,N_3634);
nand U6368 (N_6368,N_2672,N_3543);
and U6369 (N_6369,N_4383,N_3274);
and U6370 (N_6370,N_4040,N_4292);
and U6371 (N_6371,N_4030,N_3785);
nor U6372 (N_6372,N_4420,N_2750);
or U6373 (N_6373,N_3985,N_3251);
nand U6374 (N_6374,N_3026,N_4880);
nor U6375 (N_6375,N_4583,N_3179);
nor U6376 (N_6376,N_4903,N_4617);
nor U6377 (N_6377,N_2912,N_3481);
and U6378 (N_6378,N_3982,N_2611);
or U6379 (N_6379,N_3685,N_3885);
nor U6380 (N_6380,N_3262,N_4183);
nand U6381 (N_6381,N_3097,N_2844);
and U6382 (N_6382,N_3726,N_4585);
and U6383 (N_6383,N_2551,N_2513);
and U6384 (N_6384,N_3534,N_3557);
and U6385 (N_6385,N_4570,N_3744);
nor U6386 (N_6386,N_4961,N_4565);
nand U6387 (N_6387,N_4879,N_3306);
or U6388 (N_6388,N_4071,N_2655);
or U6389 (N_6389,N_4791,N_3580);
nor U6390 (N_6390,N_2666,N_4752);
nand U6391 (N_6391,N_3159,N_4077);
nand U6392 (N_6392,N_4229,N_4981);
nand U6393 (N_6393,N_3542,N_4316);
nor U6394 (N_6394,N_3678,N_2596);
xor U6395 (N_6395,N_3124,N_3823);
or U6396 (N_6396,N_3080,N_3403);
nor U6397 (N_6397,N_3514,N_4259);
and U6398 (N_6398,N_3852,N_4655);
or U6399 (N_6399,N_3157,N_4867);
nor U6400 (N_6400,N_3298,N_3379);
and U6401 (N_6401,N_4116,N_4455);
and U6402 (N_6402,N_3119,N_4615);
xnor U6403 (N_6403,N_2655,N_3241);
nand U6404 (N_6404,N_4353,N_4999);
nor U6405 (N_6405,N_2958,N_4752);
nor U6406 (N_6406,N_4887,N_3036);
or U6407 (N_6407,N_3185,N_4969);
and U6408 (N_6408,N_3545,N_4882);
nand U6409 (N_6409,N_3682,N_3869);
or U6410 (N_6410,N_3461,N_3538);
and U6411 (N_6411,N_3820,N_4515);
or U6412 (N_6412,N_3590,N_3250);
nand U6413 (N_6413,N_4217,N_3292);
nand U6414 (N_6414,N_4699,N_3097);
and U6415 (N_6415,N_3199,N_4282);
and U6416 (N_6416,N_3442,N_3146);
and U6417 (N_6417,N_3064,N_3080);
or U6418 (N_6418,N_3969,N_2939);
or U6419 (N_6419,N_4023,N_3490);
and U6420 (N_6420,N_4871,N_4119);
and U6421 (N_6421,N_3918,N_3624);
nand U6422 (N_6422,N_2513,N_3021);
and U6423 (N_6423,N_4333,N_4702);
nor U6424 (N_6424,N_4030,N_3849);
and U6425 (N_6425,N_3541,N_4925);
nor U6426 (N_6426,N_3917,N_3012);
or U6427 (N_6427,N_2572,N_3422);
nand U6428 (N_6428,N_3525,N_4129);
and U6429 (N_6429,N_3497,N_4116);
nand U6430 (N_6430,N_4502,N_4347);
nand U6431 (N_6431,N_3202,N_4391);
nand U6432 (N_6432,N_2507,N_4394);
nor U6433 (N_6433,N_3414,N_4563);
nor U6434 (N_6434,N_3126,N_3761);
or U6435 (N_6435,N_3159,N_3698);
and U6436 (N_6436,N_3299,N_2787);
nor U6437 (N_6437,N_4213,N_4922);
nand U6438 (N_6438,N_2961,N_4909);
nand U6439 (N_6439,N_2599,N_4541);
and U6440 (N_6440,N_4178,N_3603);
nand U6441 (N_6441,N_3697,N_4445);
and U6442 (N_6442,N_3171,N_3933);
or U6443 (N_6443,N_4144,N_3907);
nand U6444 (N_6444,N_4398,N_3303);
nand U6445 (N_6445,N_2505,N_2667);
and U6446 (N_6446,N_2907,N_2837);
and U6447 (N_6447,N_4033,N_3160);
or U6448 (N_6448,N_3033,N_3743);
and U6449 (N_6449,N_3386,N_4986);
or U6450 (N_6450,N_3123,N_4961);
or U6451 (N_6451,N_2997,N_2600);
nand U6452 (N_6452,N_3858,N_3310);
nor U6453 (N_6453,N_2618,N_4859);
and U6454 (N_6454,N_4131,N_4606);
and U6455 (N_6455,N_4068,N_2571);
and U6456 (N_6456,N_3263,N_3127);
nand U6457 (N_6457,N_2954,N_3372);
and U6458 (N_6458,N_4990,N_3318);
nand U6459 (N_6459,N_2805,N_3574);
nand U6460 (N_6460,N_4423,N_2929);
nand U6461 (N_6461,N_3662,N_4300);
or U6462 (N_6462,N_4523,N_3107);
or U6463 (N_6463,N_4903,N_4226);
or U6464 (N_6464,N_4390,N_2587);
and U6465 (N_6465,N_3881,N_3697);
or U6466 (N_6466,N_4895,N_3358);
nor U6467 (N_6467,N_4765,N_4613);
or U6468 (N_6468,N_4427,N_3851);
nor U6469 (N_6469,N_2646,N_2849);
or U6470 (N_6470,N_2836,N_4441);
and U6471 (N_6471,N_2575,N_3371);
and U6472 (N_6472,N_4832,N_2510);
or U6473 (N_6473,N_2946,N_2593);
nor U6474 (N_6474,N_3816,N_3479);
or U6475 (N_6475,N_2725,N_3358);
or U6476 (N_6476,N_3704,N_2630);
nand U6477 (N_6477,N_4327,N_2791);
nand U6478 (N_6478,N_3196,N_4279);
and U6479 (N_6479,N_3179,N_3017);
or U6480 (N_6480,N_2873,N_4201);
nand U6481 (N_6481,N_2676,N_3119);
or U6482 (N_6482,N_2694,N_4759);
nand U6483 (N_6483,N_3883,N_3914);
nand U6484 (N_6484,N_3925,N_3794);
or U6485 (N_6485,N_2589,N_2982);
or U6486 (N_6486,N_4517,N_2524);
or U6487 (N_6487,N_2801,N_3414);
nand U6488 (N_6488,N_2981,N_3134);
xnor U6489 (N_6489,N_4435,N_4733);
or U6490 (N_6490,N_2984,N_3689);
or U6491 (N_6491,N_3315,N_4688);
nor U6492 (N_6492,N_2830,N_3064);
nand U6493 (N_6493,N_4574,N_3338);
nand U6494 (N_6494,N_4717,N_4130);
or U6495 (N_6495,N_3748,N_3929);
or U6496 (N_6496,N_2742,N_2718);
or U6497 (N_6497,N_4497,N_4002);
and U6498 (N_6498,N_3762,N_2960);
or U6499 (N_6499,N_4060,N_3381);
nand U6500 (N_6500,N_3800,N_4632);
or U6501 (N_6501,N_4223,N_4521);
xor U6502 (N_6502,N_4274,N_4670);
nand U6503 (N_6503,N_3397,N_3578);
and U6504 (N_6504,N_4404,N_2645);
xor U6505 (N_6505,N_4688,N_3809);
nor U6506 (N_6506,N_4436,N_4533);
nand U6507 (N_6507,N_3012,N_4291);
nand U6508 (N_6508,N_3609,N_4979);
or U6509 (N_6509,N_2929,N_3121);
nor U6510 (N_6510,N_3296,N_2738);
or U6511 (N_6511,N_3682,N_4787);
and U6512 (N_6512,N_4867,N_2743);
nor U6513 (N_6513,N_3186,N_2584);
or U6514 (N_6514,N_3279,N_3789);
and U6515 (N_6515,N_4473,N_3445);
or U6516 (N_6516,N_3560,N_3940);
and U6517 (N_6517,N_3083,N_3944);
xor U6518 (N_6518,N_3768,N_3722);
nor U6519 (N_6519,N_3015,N_4288);
nand U6520 (N_6520,N_3819,N_3151);
nor U6521 (N_6521,N_3648,N_3194);
xor U6522 (N_6522,N_3698,N_4831);
nand U6523 (N_6523,N_2521,N_3117);
or U6524 (N_6524,N_4610,N_4053);
nand U6525 (N_6525,N_4060,N_4614);
and U6526 (N_6526,N_2999,N_3472);
nor U6527 (N_6527,N_3964,N_4606);
nor U6528 (N_6528,N_4908,N_4281);
nor U6529 (N_6529,N_3072,N_4830);
xor U6530 (N_6530,N_4496,N_4985);
nor U6531 (N_6531,N_3708,N_3430);
or U6532 (N_6532,N_3773,N_2730);
or U6533 (N_6533,N_3591,N_4023);
nand U6534 (N_6534,N_2993,N_4719);
or U6535 (N_6535,N_3821,N_2775);
or U6536 (N_6536,N_3852,N_4651);
xor U6537 (N_6537,N_2735,N_2906);
nand U6538 (N_6538,N_4841,N_3878);
or U6539 (N_6539,N_3651,N_4045);
nand U6540 (N_6540,N_4061,N_3751);
nand U6541 (N_6541,N_4881,N_4904);
or U6542 (N_6542,N_4000,N_3794);
and U6543 (N_6543,N_4785,N_2707);
nand U6544 (N_6544,N_4414,N_3812);
or U6545 (N_6545,N_3874,N_3419);
and U6546 (N_6546,N_4966,N_3754);
or U6547 (N_6547,N_2801,N_2977);
xnor U6548 (N_6548,N_4577,N_4143);
nor U6549 (N_6549,N_2758,N_2930);
nand U6550 (N_6550,N_4125,N_3383);
nand U6551 (N_6551,N_3230,N_4169);
or U6552 (N_6552,N_2942,N_2818);
nor U6553 (N_6553,N_3717,N_4168);
nor U6554 (N_6554,N_2884,N_4371);
or U6555 (N_6555,N_3990,N_4127);
and U6556 (N_6556,N_2500,N_3732);
nor U6557 (N_6557,N_4100,N_2707);
and U6558 (N_6558,N_3386,N_3129);
nand U6559 (N_6559,N_4984,N_3981);
or U6560 (N_6560,N_2590,N_3909);
or U6561 (N_6561,N_2951,N_4623);
nor U6562 (N_6562,N_2594,N_3989);
and U6563 (N_6563,N_4333,N_3485);
and U6564 (N_6564,N_3883,N_3386);
or U6565 (N_6565,N_4631,N_3122);
nand U6566 (N_6566,N_3861,N_4699);
nor U6567 (N_6567,N_3197,N_4594);
nand U6568 (N_6568,N_2976,N_4762);
or U6569 (N_6569,N_3627,N_4865);
nor U6570 (N_6570,N_3727,N_3796);
or U6571 (N_6571,N_3584,N_3901);
nor U6572 (N_6572,N_4982,N_4248);
nand U6573 (N_6573,N_3016,N_4488);
nor U6574 (N_6574,N_2727,N_4431);
nor U6575 (N_6575,N_4131,N_4250);
and U6576 (N_6576,N_3889,N_3909);
or U6577 (N_6577,N_2995,N_3496);
nand U6578 (N_6578,N_4620,N_4224);
nand U6579 (N_6579,N_3666,N_3092);
or U6580 (N_6580,N_4163,N_4848);
nor U6581 (N_6581,N_2675,N_2691);
nor U6582 (N_6582,N_4794,N_4862);
nand U6583 (N_6583,N_3612,N_3404);
or U6584 (N_6584,N_4883,N_3024);
xnor U6585 (N_6585,N_3884,N_4095);
nand U6586 (N_6586,N_4276,N_2932);
nor U6587 (N_6587,N_3871,N_4276);
nand U6588 (N_6588,N_4470,N_2679);
nor U6589 (N_6589,N_4411,N_3832);
or U6590 (N_6590,N_2603,N_4727);
or U6591 (N_6591,N_3041,N_3392);
or U6592 (N_6592,N_4754,N_3812);
nand U6593 (N_6593,N_3058,N_4696);
or U6594 (N_6594,N_4360,N_4389);
nand U6595 (N_6595,N_4047,N_3024);
nand U6596 (N_6596,N_4082,N_3704);
or U6597 (N_6597,N_2703,N_4010);
and U6598 (N_6598,N_4822,N_4441);
nor U6599 (N_6599,N_2585,N_3475);
and U6600 (N_6600,N_4930,N_3374);
nand U6601 (N_6601,N_3433,N_3413);
nand U6602 (N_6602,N_4255,N_4439);
nor U6603 (N_6603,N_3962,N_4591);
nor U6604 (N_6604,N_3909,N_3803);
xor U6605 (N_6605,N_2693,N_3482);
and U6606 (N_6606,N_4975,N_2740);
nor U6607 (N_6607,N_3835,N_4123);
nor U6608 (N_6608,N_3040,N_4855);
and U6609 (N_6609,N_3085,N_4622);
or U6610 (N_6610,N_3815,N_2685);
nand U6611 (N_6611,N_4936,N_4685);
nor U6612 (N_6612,N_3465,N_4946);
nand U6613 (N_6613,N_2532,N_3817);
nor U6614 (N_6614,N_3630,N_4813);
nor U6615 (N_6615,N_4143,N_4898);
nor U6616 (N_6616,N_3581,N_4936);
nor U6617 (N_6617,N_4736,N_3087);
and U6618 (N_6618,N_3505,N_4773);
nand U6619 (N_6619,N_3681,N_2595);
or U6620 (N_6620,N_3660,N_2860);
nor U6621 (N_6621,N_2738,N_2743);
nand U6622 (N_6622,N_3901,N_4239);
and U6623 (N_6623,N_4384,N_4347);
or U6624 (N_6624,N_4036,N_2601);
xnor U6625 (N_6625,N_3430,N_3754);
or U6626 (N_6626,N_3009,N_3819);
nand U6627 (N_6627,N_4331,N_4252);
and U6628 (N_6628,N_3135,N_4386);
nor U6629 (N_6629,N_4974,N_3808);
and U6630 (N_6630,N_4434,N_4245);
or U6631 (N_6631,N_3179,N_2741);
nor U6632 (N_6632,N_2713,N_4049);
and U6633 (N_6633,N_4977,N_3487);
and U6634 (N_6634,N_4501,N_4261);
nor U6635 (N_6635,N_3005,N_4547);
nor U6636 (N_6636,N_3493,N_3259);
nor U6637 (N_6637,N_4428,N_2923);
and U6638 (N_6638,N_3923,N_4598);
nand U6639 (N_6639,N_4909,N_3232);
or U6640 (N_6640,N_3093,N_2539);
or U6641 (N_6641,N_3546,N_4186);
and U6642 (N_6642,N_4776,N_4074);
and U6643 (N_6643,N_3005,N_3187);
and U6644 (N_6644,N_3129,N_4576);
or U6645 (N_6645,N_2967,N_3386);
nor U6646 (N_6646,N_3336,N_2602);
and U6647 (N_6647,N_2764,N_2571);
nand U6648 (N_6648,N_3162,N_4049);
and U6649 (N_6649,N_4501,N_3958);
xor U6650 (N_6650,N_2550,N_2874);
or U6651 (N_6651,N_3193,N_4337);
nor U6652 (N_6652,N_4437,N_4899);
nand U6653 (N_6653,N_3640,N_2677);
nand U6654 (N_6654,N_3868,N_2680);
or U6655 (N_6655,N_3544,N_3183);
nand U6656 (N_6656,N_3659,N_4099);
nand U6657 (N_6657,N_3040,N_3370);
and U6658 (N_6658,N_4958,N_2912);
nor U6659 (N_6659,N_3788,N_4656);
nor U6660 (N_6660,N_3250,N_4786);
and U6661 (N_6661,N_3567,N_3407);
and U6662 (N_6662,N_2879,N_3314);
nand U6663 (N_6663,N_3814,N_3804);
nor U6664 (N_6664,N_3686,N_4502);
and U6665 (N_6665,N_3236,N_2571);
and U6666 (N_6666,N_4275,N_3305);
nand U6667 (N_6667,N_3004,N_3809);
and U6668 (N_6668,N_4410,N_3883);
and U6669 (N_6669,N_2691,N_4200);
and U6670 (N_6670,N_4026,N_2660);
nand U6671 (N_6671,N_4455,N_3413);
or U6672 (N_6672,N_4973,N_3654);
nor U6673 (N_6673,N_2752,N_4465);
and U6674 (N_6674,N_4511,N_3090);
nor U6675 (N_6675,N_4684,N_3922);
and U6676 (N_6676,N_3718,N_3875);
nand U6677 (N_6677,N_3973,N_3357);
and U6678 (N_6678,N_4374,N_4992);
or U6679 (N_6679,N_2625,N_3661);
or U6680 (N_6680,N_2912,N_2553);
nor U6681 (N_6681,N_4259,N_3197);
nand U6682 (N_6682,N_4891,N_3597);
nor U6683 (N_6683,N_3671,N_3420);
and U6684 (N_6684,N_2721,N_4955);
nand U6685 (N_6685,N_3730,N_4461);
or U6686 (N_6686,N_4708,N_4757);
nand U6687 (N_6687,N_3722,N_4040);
nor U6688 (N_6688,N_4580,N_3180);
or U6689 (N_6689,N_3864,N_2646);
and U6690 (N_6690,N_2732,N_3126);
nor U6691 (N_6691,N_3766,N_2615);
nor U6692 (N_6692,N_4003,N_4899);
nor U6693 (N_6693,N_4814,N_4790);
and U6694 (N_6694,N_3317,N_2822);
or U6695 (N_6695,N_4984,N_3141);
nand U6696 (N_6696,N_4057,N_2847);
and U6697 (N_6697,N_3795,N_3345);
and U6698 (N_6698,N_2943,N_4088);
and U6699 (N_6699,N_3939,N_4951);
or U6700 (N_6700,N_3177,N_3549);
xor U6701 (N_6701,N_3594,N_4825);
nor U6702 (N_6702,N_2800,N_4782);
nor U6703 (N_6703,N_4979,N_4404);
or U6704 (N_6704,N_3966,N_2908);
nand U6705 (N_6705,N_3223,N_4227);
and U6706 (N_6706,N_4169,N_3792);
xor U6707 (N_6707,N_4033,N_4089);
nor U6708 (N_6708,N_4389,N_3408);
nand U6709 (N_6709,N_3761,N_3232);
and U6710 (N_6710,N_4612,N_3305);
or U6711 (N_6711,N_2560,N_2808);
and U6712 (N_6712,N_3874,N_3983);
and U6713 (N_6713,N_4782,N_3386);
or U6714 (N_6714,N_4414,N_2561);
or U6715 (N_6715,N_3218,N_3202);
or U6716 (N_6716,N_4150,N_4887);
or U6717 (N_6717,N_3524,N_2753);
and U6718 (N_6718,N_4058,N_4282);
nand U6719 (N_6719,N_2934,N_4793);
nand U6720 (N_6720,N_4883,N_3069);
and U6721 (N_6721,N_4801,N_4227);
or U6722 (N_6722,N_4050,N_3098);
or U6723 (N_6723,N_4644,N_2998);
or U6724 (N_6724,N_4602,N_3018);
nand U6725 (N_6725,N_4338,N_4448);
xnor U6726 (N_6726,N_4311,N_4894);
xnor U6727 (N_6727,N_3049,N_4005);
or U6728 (N_6728,N_2755,N_3853);
nor U6729 (N_6729,N_4061,N_2594);
and U6730 (N_6730,N_3389,N_3822);
or U6731 (N_6731,N_3194,N_2780);
or U6732 (N_6732,N_4938,N_4312);
and U6733 (N_6733,N_3359,N_2796);
nor U6734 (N_6734,N_3978,N_3109);
or U6735 (N_6735,N_4595,N_3554);
and U6736 (N_6736,N_2592,N_2871);
nand U6737 (N_6737,N_3133,N_3112);
and U6738 (N_6738,N_3948,N_4562);
nor U6739 (N_6739,N_4854,N_3135);
nand U6740 (N_6740,N_4498,N_4133);
nand U6741 (N_6741,N_4323,N_3350);
and U6742 (N_6742,N_3694,N_3639);
nor U6743 (N_6743,N_3740,N_3614);
or U6744 (N_6744,N_4256,N_2593);
nand U6745 (N_6745,N_4532,N_2855);
or U6746 (N_6746,N_3219,N_4976);
nand U6747 (N_6747,N_2652,N_3524);
or U6748 (N_6748,N_2557,N_4412);
and U6749 (N_6749,N_4269,N_3751);
nor U6750 (N_6750,N_4675,N_4509);
nand U6751 (N_6751,N_4031,N_4099);
nor U6752 (N_6752,N_3047,N_3708);
and U6753 (N_6753,N_2606,N_3518);
nand U6754 (N_6754,N_3333,N_4662);
and U6755 (N_6755,N_4002,N_2753);
xnor U6756 (N_6756,N_3514,N_4993);
and U6757 (N_6757,N_3683,N_2861);
and U6758 (N_6758,N_3659,N_4619);
and U6759 (N_6759,N_4236,N_4208);
nand U6760 (N_6760,N_3774,N_4456);
and U6761 (N_6761,N_3038,N_2793);
or U6762 (N_6762,N_2602,N_3738);
xnor U6763 (N_6763,N_2874,N_3509);
nor U6764 (N_6764,N_4417,N_4503);
nand U6765 (N_6765,N_4358,N_3493);
or U6766 (N_6766,N_2716,N_4782);
nor U6767 (N_6767,N_2572,N_3081);
or U6768 (N_6768,N_3325,N_4126);
and U6769 (N_6769,N_3561,N_4010);
or U6770 (N_6770,N_3235,N_4716);
and U6771 (N_6771,N_4897,N_4286);
nor U6772 (N_6772,N_3320,N_3108);
and U6773 (N_6773,N_2583,N_2832);
and U6774 (N_6774,N_3444,N_3521);
nor U6775 (N_6775,N_2511,N_4527);
or U6776 (N_6776,N_4129,N_4060);
or U6777 (N_6777,N_2953,N_2952);
or U6778 (N_6778,N_2709,N_4365);
nor U6779 (N_6779,N_3053,N_4580);
and U6780 (N_6780,N_4513,N_2805);
or U6781 (N_6781,N_4746,N_3282);
and U6782 (N_6782,N_4407,N_4815);
or U6783 (N_6783,N_2933,N_3361);
and U6784 (N_6784,N_2769,N_3526);
nor U6785 (N_6785,N_4196,N_4727);
or U6786 (N_6786,N_3892,N_2610);
or U6787 (N_6787,N_3716,N_3948);
nor U6788 (N_6788,N_3601,N_4559);
and U6789 (N_6789,N_4973,N_3931);
and U6790 (N_6790,N_3917,N_4733);
nand U6791 (N_6791,N_3392,N_4429);
and U6792 (N_6792,N_3576,N_2654);
nor U6793 (N_6793,N_3285,N_4115);
or U6794 (N_6794,N_3433,N_4220);
xnor U6795 (N_6795,N_2678,N_3366);
nand U6796 (N_6796,N_4748,N_2768);
and U6797 (N_6797,N_3176,N_3223);
and U6798 (N_6798,N_3943,N_3665);
or U6799 (N_6799,N_2979,N_4278);
nand U6800 (N_6800,N_3929,N_2654);
and U6801 (N_6801,N_2668,N_3526);
nor U6802 (N_6802,N_3778,N_3356);
or U6803 (N_6803,N_4641,N_3465);
or U6804 (N_6804,N_4085,N_3446);
nand U6805 (N_6805,N_4921,N_3798);
or U6806 (N_6806,N_3632,N_3971);
or U6807 (N_6807,N_4539,N_3571);
and U6808 (N_6808,N_3859,N_3893);
nor U6809 (N_6809,N_2957,N_3456);
and U6810 (N_6810,N_4749,N_3607);
nand U6811 (N_6811,N_4528,N_3296);
and U6812 (N_6812,N_3899,N_3271);
nor U6813 (N_6813,N_3256,N_3236);
and U6814 (N_6814,N_3350,N_3821);
and U6815 (N_6815,N_2945,N_4612);
or U6816 (N_6816,N_4541,N_3692);
nor U6817 (N_6817,N_4898,N_4022);
nand U6818 (N_6818,N_3589,N_3205);
nor U6819 (N_6819,N_3861,N_2751);
or U6820 (N_6820,N_4169,N_3910);
nand U6821 (N_6821,N_4253,N_4876);
and U6822 (N_6822,N_4723,N_4675);
nor U6823 (N_6823,N_2769,N_2578);
and U6824 (N_6824,N_4658,N_2578);
nor U6825 (N_6825,N_3446,N_2546);
and U6826 (N_6826,N_3166,N_2728);
and U6827 (N_6827,N_3015,N_3494);
nor U6828 (N_6828,N_3973,N_4491);
nor U6829 (N_6829,N_2985,N_4630);
or U6830 (N_6830,N_2956,N_4182);
or U6831 (N_6831,N_4767,N_2907);
or U6832 (N_6832,N_4811,N_3660);
nor U6833 (N_6833,N_2884,N_4936);
and U6834 (N_6834,N_2814,N_3319);
nand U6835 (N_6835,N_3789,N_4379);
and U6836 (N_6836,N_3910,N_3908);
and U6837 (N_6837,N_3882,N_3581);
nor U6838 (N_6838,N_3813,N_4474);
or U6839 (N_6839,N_4909,N_4955);
nand U6840 (N_6840,N_3934,N_2784);
nand U6841 (N_6841,N_3787,N_2565);
nand U6842 (N_6842,N_3305,N_3253);
nand U6843 (N_6843,N_3602,N_4225);
or U6844 (N_6844,N_2819,N_4938);
or U6845 (N_6845,N_3597,N_4113);
and U6846 (N_6846,N_4081,N_4841);
nor U6847 (N_6847,N_4750,N_2549);
and U6848 (N_6848,N_3542,N_2755);
and U6849 (N_6849,N_3388,N_3320);
and U6850 (N_6850,N_3766,N_3327);
nor U6851 (N_6851,N_2844,N_3985);
nand U6852 (N_6852,N_2866,N_3666);
and U6853 (N_6853,N_2805,N_4325);
nand U6854 (N_6854,N_4943,N_3512);
and U6855 (N_6855,N_3793,N_4011);
or U6856 (N_6856,N_3298,N_3235);
nor U6857 (N_6857,N_3916,N_3914);
or U6858 (N_6858,N_2976,N_2714);
xnor U6859 (N_6859,N_4704,N_2791);
nand U6860 (N_6860,N_3557,N_4341);
nand U6861 (N_6861,N_3415,N_4767);
xor U6862 (N_6862,N_4700,N_2765);
nand U6863 (N_6863,N_3417,N_2501);
nand U6864 (N_6864,N_4108,N_4699);
nand U6865 (N_6865,N_4065,N_2752);
and U6866 (N_6866,N_4669,N_3161);
or U6867 (N_6867,N_3266,N_4432);
nor U6868 (N_6868,N_4012,N_3920);
or U6869 (N_6869,N_3110,N_3108);
nor U6870 (N_6870,N_4415,N_3234);
nor U6871 (N_6871,N_2511,N_3188);
nor U6872 (N_6872,N_3250,N_3268);
or U6873 (N_6873,N_2703,N_4372);
and U6874 (N_6874,N_3681,N_3094);
and U6875 (N_6875,N_2556,N_4657);
and U6876 (N_6876,N_4635,N_3327);
nor U6877 (N_6877,N_2503,N_3402);
nor U6878 (N_6878,N_4098,N_2993);
or U6879 (N_6879,N_4661,N_4551);
nand U6880 (N_6880,N_4109,N_3650);
and U6881 (N_6881,N_2981,N_3413);
and U6882 (N_6882,N_2881,N_3122);
and U6883 (N_6883,N_4332,N_4911);
nand U6884 (N_6884,N_4994,N_4318);
nor U6885 (N_6885,N_4719,N_4030);
or U6886 (N_6886,N_4411,N_4386);
nand U6887 (N_6887,N_2948,N_3884);
nor U6888 (N_6888,N_4933,N_3144);
and U6889 (N_6889,N_4310,N_3420);
nand U6890 (N_6890,N_4571,N_3420);
or U6891 (N_6891,N_4226,N_3415);
xnor U6892 (N_6892,N_4582,N_4323);
xnor U6893 (N_6893,N_3978,N_4780);
or U6894 (N_6894,N_4318,N_3631);
nor U6895 (N_6895,N_4007,N_4987);
nor U6896 (N_6896,N_2693,N_3656);
or U6897 (N_6897,N_2675,N_3672);
and U6898 (N_6898,N_3600,N_4091);
xor U6899 (N_6899,N_2651,N_3317);
or U6900 (N_6900,N_3530,N_3418);
nand U6901 (N_6901,N_4747,N_4852);
and U6902 (N_6902,N_4416,N_2740);
or U6903 (N_6903,N_3844,N_2769);
and U6904 (N_6904,N_3967,N_4057);
or U6905 (N_6905,N_2771,N_3933);
nand U6906 (N_6906,N_4747,N_4574);
or U6907 (N_6907,N_3400,N_4007);
nand U6908 (N_6908,N_4468,N_3388);
or U6909 (N_6909,N_3222,N_2687);
nand U6910 (N_6910,N_2978,N_2761);
or U6911 (N_6911,N_3330,N_3207);
or U6912 (N_6912,N_3654,N_2742);
nand U6913 (N_6913,N_3549,N_3718);
and U6914 (N_6914,N_4178,N_3989);
or U6915 (N_6915,N_3074,N_3076);
and U6916 (N_6916,N_3188,N_3527);
or U6917 (N_6917,N_4901,N_2504);
and U6918 (N_6918,N_2850,N_4520);
or U6919 (N_6919,N_3196,N_2791);
or U6920 (N_6920,N_3336,N_4185);
nand U6921 (N_6921,N_3932,N_2635);
nand U6922 (N_6922,N_4734,N_3683);
nand U6923 (N_6923,N_3044,N_3570);
xnor U6924 (N_6924,N_3758,N_2550);
and U6925 (N_6925,N_3852,N_2806);
or U6926 (N_6926,N_4319,N_4477);
and U6927 (N_6927,N_4616,N_4508);
and U6928 (N_6928,N_2971,N_4979);
and U6929 (N_6929,N_3020,N_3458);
and U6930 (N_6930,N_2673,N_4581);
and U6931 (N_6931,N_4823,N_3936);
nand U6932 (N_6932,N_3562,N_4137);
nand U6933 (N_6933,N_3111,N_2680);
and U6934 (N_6934,N_3684,N_4517);
xor U6935 (N_6935,N_4919,N_2804);
nor U6936 (N_6936,N_3705,N_3111);
and U6937 (N_6937,N_3793,N_2961);
or U6938 (N_6938,N_3712,N_4140);
nand U6939 (N_6939,N_3147,N_4621);
nor U6940 (N_6940,N_4520,N_4887);
nor U6941 (N_6941,N_3268,N_2762);
nor U6942 (N_6942,N_3367,N_2873);
nand U6943 (N_6943,N_4448,N_3723);
nand U6944 (N_6944,N_4631,N_3852);
and U6945 (N_6945,N_3524,N_3030);
nand U6946 (N_6946,N_4673,N_3522);
or U6947 (N_6947,N_2910,N_3142);
nor U6948 (N_6948,N_4509,N_3202);
nand U6949 (N_6949,N_4266,N_4863);
nand U6950 (N_6950,N_4429,N_4293);
nand U6951 (N_6951,N_3551,N_3669);
nand U6952 (N_6952,N_3938,N_4522);
nand U6953 (N_6953,N_3021,N_4474);
or U6954 (N_6954,N_3939,N_2679);
nor U6955 (N_6955,N_2528,N_3290);
or U6956 (N_6956,N_3083,N_4410);
nor U6957 (N_6957,N_4309,N_4679);
and U6958 (N_6958,N_2679,N_3125);
or U6959 (N_6959,N_4923,N_3700);
or U6960 (N_6960,N_4903,N_4418);
nor U6961 (N_6961,N_3701,N_4541);
nor U6962 (N_6962,N_2696,N_4196);
or U6963 (N_6963,N_3128,N_3955);
nor U6964 (N_6964,N_3060,N_4931);
and U6965 (N_6965,N_4543,N_3549);
nand U6966 (N_6966,N_3441,N_3198);
and U6967 (N_6967,N_4228,N_3120);
and U6968 (N_6968,N_2587,N_4852);
nor U6969 (N_6969,N_4604,N_2513);
nor U6970 (N_6970,N_4233,N_3216);
and U6971 (N_6971,N_3448,N_4752);
nor U6972 (N_6972,N_2867,N_4119);
xor U6973 (N_6973,N_4629,N_3141);
or U6974 (N_6974,N_3355,N_3283);
and U6975 (N_6975,N_3294,N_3478);
nor U6976 (N_6976,N_4691,N_4907);
and U6977 (N_6977,N_4883,N_2674);
and U6978 (N_6978,N_3436,N_3269);
or U6979 (N_6979,N_3468,N_2563);
or U6980 (N_6980,N_3767,N_2502);
nor U6981 (N_6981,N_3257,N_3920);
nor U6982 (N_6982,N_4629,N_2937);
or U6983 (N_6983,N_2793,N_2832);
and U6984 (N_6984,N_3930,N_3918);
and U6985 (N_6985,N_4020,N_3325);
and U6986 (N_6986,N_4139,N_2546);
nor U6987 (N_6987,N_4679,N_4696);
nand U6988 (N_6988,N_4518,N_3293);
nand U6989 (N_6989,N_3107,N_3585);
or U6990 (N_6990,N_3338,N_3254);
nor U6991 (N_6991,N_3900,N_3691);
or U6992 (N_6992,N_3703,N_2823);
xor U6993 (N_6993,N_2960,N_2536);
and U6994 (N_6994,N_4355,N_4741);
nand U6995 (N_6995,N_2809,N_3917);
and U6996 (N_6996,N_2668,N_3652);
or U6997 (N_6997,N_4510,N_4889);
nand U6998 (N_6998,N_2991,N_4430);
nor U6999 (N_6999,N_2963,N_3168);
or U7000 (N_7000,N_3947,N_4010);
or U7001 (N_7001,N_3760,N_2730);
or U7002 (N_7002,N_2564,N_4380);
nor U7003 (N_7003,N_3252,N_3760);
and U7004 (N_7004,N_4212,N_4960);
or U7005 (N_7005,N_3898,N_3130);
nand U7006 (N_7006,N_4338,N_4277);
nor U7007 (N_7007,N_2842,N_2531);
nand U7008 (N_7008,N_3775,N_4783);
and U7009 (N_7009,N_4249,N_4327);
nor U7010 (N_7010,N_3454,N_4198);
and U7011 (N_7011,N_3012,N_2853);
nor U7012 (N_7012,N_2917,N_4980);
or U7013 (N_7013,N_3568,N_3354);
or U7014 (N_7014,N_3583,N_2533);
and U7015 (N_7015,N_4647,N_3879);
xor U7016 (N_7016,N_3729,N_4119);
nor U7017 (N_7017,N_3081,N_4991);
nand U7018 (N_7018,N_2922,N_3628);
and U7019 (N_7019,N_4658,N_2507);
nor U7020 (N_7020,N_4385,N_3196);
nor U7021 (N_7021,N_2539,N_4646);
nor U7022 (N_7022,N_2995,N_3959);
and U7023 (N_7023,N_4589,N_3811);
and U7024 (N_7024,N_2925,N_4000);
xor U7025 (N_7025,N_3792,N_4374);
nor U7026 (N_7026,N_4269,N_2873);
nor U7027 (N_7027,N_2789,N_2895);
xor U7028 (N_7028,N_4048,N_4255);
nand U7029 (N_7029,N_3374,N_4199);
and U7030 (N_7030,N_3977,N_4613);
or U7031 (N_7031,N_2925,N_3816);
or U7032 (N_7032,N_2698,N_4811);
or U7033 (N_7033,N_4117,N_4809);
or U7034 (N_7034,N_4977,N_2616);
nand U7035 (N_7035,N_3531,N_2674);
xor U7036 (N_7036,N_3075,N_4217);
and U7037 (N_7037,N_3252,N_3254);
or U7038 (N_7038,N_4000,N_3612);
and U7039 (N_7039,N_4376,N_2835);
and U7040 (N_7040,N_2718,N_4735);
or U7041 (N_7041,N_4084,N_3823);
nor U7042 (N_7042,N_2957,N_4220);
nor U7043 (N_7043,N_4934,N_4210);
and U7044 (N_7044,N_3264,N_3496);
nand U7045 (N_7045,N_4878,N_3102);
nor U7046 (N_7046,N_4552,N_2624);
or U7047 (N_7047,N_4899,N_2666);
nand U7048 (N_7048,N_4141,N_3251);
nand U7049 (N_7049,N_2570,N_2741);
nor U7050 (N_7050,N_4099,N_3834);
or U7051 (N_7051,N_4106,N_2707);
and U7052 (N_7052,N_4242,N_4585);
nand U7053 (N_7053,N_4490,N_3666);
nand U7054 (N_7054,N_3555,N_2571);
nand U7055 (N_7055,N_2697,N_3600);
nand U7056 (N_7056,N_3334,N_4478);
and U7057 (N_7057,N_4634,N_2601);
nand U7058 (N_7058,N_2795,N_4987);
or U7059 (N_7059,N_2645,N_3836);
xor U7060 (N_7060,N_3812,N_2832);
nor U7061 (N_7061,N_3318,N_2968);
nand U7062 (N_7062,N_3557,N_2914);
or U7063 (N_7063,N_2936,N_2932);
nor U7064 (N_7064,N_3974,N_2983);
or U7065 (N_7065,N_3061,N_4315);
nor U7066 (N_7066,N_2989,N_4305);
or U7067 (N_7067,N_4845,N_3873);
or U7068 (N_7068,N_4172,N_4180);
or U7069 (N_7069,N_2986,N_3921);
and U7070 (N_7070,N_4981,N_3054);
nor U7071 (N_7071,N_2811,N_4430);
nand U7072 (N_7072,N_4805,N_3676);
or U7073 (N_7073,N_3319,N_2990);
nand U7074 (N_7074,N_3063,N_4126);
or U7075 (N_7075,N_3148,N_4841);
and U7076 (N_7076,N_2713,N_4738);
or U7077 (N_7077,N_3486,N_4323);
nand U7078 (N_7078,N_4635,N_3644);
nand U7079 (N_7079,N_4621,N_3024);
and U7080 (N_7080,N_4489,N_2636);
or U7081 (N_7081,N_3232,N_4578);
or U7082 (N_7082,N_3085,N_4076);
nand U7083 (N_7083,N_4603,N_3947);
nor U7084 (N_7084,N_4413,N_3487);
nand U7085 (N_7085,N_3844,N_4454);
and U7086 (N_7086,N_4706,N_4248);
nor U7087 (N_7087,N_4270,N_2582);
or U7088 (N_7088,N_4242,N_3994);
and U7089 (N_7089,N_4904,N_3663);
nor U7090 (N_7090,N_4783,N_3756);
or U7091 (N_7091,N_3547,N_4864);
nand U7092 (N_7092,N_4881,N_3274);
nor U7093 (N_7093,N_4271,N_2925);
and U7094 (N_7094,N_3862,N_3055);
or U7095 (N_7095,N_4299,N_2656);
and U7096 (N_7096,N_4871,N_4956);
and U7097 (N_7097,N_4947,N_4986);
and U7098 (N_7098,N_4595,N_4121);
and U7099 (N_7099,N_3399,N_4073);
or U7100 (N_7100,N_3915,N_4262);
nand U7101 (N_7101,N_3273,N_4041);
and U7102 (N_7102,N_2525,N_3838);
and U7103 (N_7103,N_3926,N_4524);
nor U7104 (N_7104,N_4378,N_3683);
nor U7105 (N_7105,N_4089,N_3452);
and U7106 (N_7106,N_4578,N_2547);
and U7107 (N_7107,N_3493,N_2853);
xor U7108 (N_7108,N_3534,N_3033);
nor U7109 (N_7109,N_2813,N_3689);
nand U7110 (N_7110,N_4913,N_2825);
or U7111 (N_7111,N_4927,N_3216);
nor U7112 (N_7112,N_4505,N_4317);
nand U7113 (N_7113,N_4199,N_4428);
or U7114 (N_7114,N_3900,N_3917);
nand U7115 (N_7115,N_4126,N_3352);
xor U7116 (N_7116,N_4034,N_3240);
and U7117 (N_7117,N_4076,N_4168);
or U7118 (N_7118,N_4334,N_4542);
and U7119 (N_7119,N_4029,N_4301);
nor U7120 (N_7120,N_3060,N_3491);
nand U7121 (N_7121,N_3799,N_3314);
or U7122 (N_7122,N_3252,N_3397);
and U7123 (N_7123,N_3984,N_3011);
nor U7124 (N_7124,N_2627,N_2625);
or U7125 (N_7125,N_3604,N_3187);
and U7126 (N_7126,N_3822,N_4844);
nand U7127 (N_7127,N_2830,N_2981);
and U7128 (N_7128,N_2695,N_2813);
or U7129 (N_7129,N_2734,N_3097);
nor U7130 (N_7130,N_4410,N_2912);
nor U7131 (N_7131,N_3076,N_4205);
nor U7132 (N_7132,N_3823,N_4938);
or U7133 (N_7133,N_4367,N_4506);
or U7134 (N_7134,N_3903,N_4532);
or U7135 (N_7135,N_3965,N_4722);
and U7136 (N_7136,N_4602,N_2752);
or U7137 (N_7137,N_3242,N_3258);
nor U7138 (N_7138,N_2619,N_3296);
and U7139 (N_7139,N_3202,N_3252);
and U7140 (N_7140,N_4339,N_3652);
and U7141 (N_7141,N_4649,N_4327);
nor U7142 (N_7142,N_4302,N_3461);
nand U7143 (N_7143,N_3853,N_2665);
nor U7144 (N_7144,N_3507,N_4885);
nor U7145 (N_7145,N_4422,N_4644);
xor U7146 (N_7146,N_2545,N_4245);
and U7147 (N_7147,N_4462,N_4149);
nand U7148 (N_7148,N_3749,N_4117);
or U7149 (N_7149,N_2573,N_3970);
nand U7150 (N_7150,N_3833,N_4721);
nand U7151 (N_7151,N_4997,N_3895);
and U7152 (N_7152,N_3341,N_4333);
and U7153 (N_7153,N_3602,N_2592);
nor U7154 (N_7154,N_3775,N_3698);
and U7155 (N_7155,N_3866,N_2968);
or U7156 (N_7156,N_3251,N_3277);
nor U7157 (N_7157,N_3698,N_3354);
nand U7158 (N_7158,N_3490,N_2865);
and U7159 (N_7159,N_3475,N_4720);
nand U7160 (N_7160,N_4269,N_4233);
or U7161 (N_7161,N_2913,N_3835);
and U7162 (N_7162,N_3145,N_4160);
and U7163 (N_7163,N_4835,N_3017);
nand U7164 (N_7164,N_4504,N_3017);
nor U7165 (N_7165,N_3813,N_2849);
xor U7166 (N_7166,N_2699,N_2760);
xnor U7167 (N_7167,N_3390,N_3709);
or U7168 (N_7168,N_4022,N_3578);
nor U7169 (N_7169,N_3446,N_3640);
and U7170 (N_7170,N_4767,N_3602);
or U7171 (N_7171,N_4805,N_4322);
nor U7172 (N_7172,N_3405,N_4880);
nand U7173 (N_7173,N_3592,N_4531);
or U7174 (N_7174,N_2575,N_4084);
xnor U7175 (N_7175,N_3881,N_4757);
xor U7176 (N_7176,N_2598,N_4970);
nor U7177 (N_7177,N_2518,N_3176);
nor U7178 (N_7178,N_4916,N_3907);
nor U7179 (N_7179,N_3524,N_3292);
nand U7180 (N_7180,N_4435,N_4157);
or U7181 (N_7181,N_4901,N_2805);
nor U7182 (N_7182,N_3550,N_4470);
and U7183 (N_7183,N_4865,N_3057);
and U7184 (N_7184,N_2760,N_4518);
nand U7185 (N_7185,N_4353,N_4665);
and U7186 (N_7186,N_4419,N_3552);
nor U7187 (N_7187,N_3083,N_2741);
and U7188 (N_7188,N_4620,N_3864);
and U7189 (N_7189,N_4555,N_2890);
nand U7190 (N_7190,N_3155,N_4412);
or U7191 (N_7191,N_3455,N_4667);
nor U7192 (N_7192,N_3773,N_4512);
or U7193 (N_7193,N_4776,N_4323);
nand U7194 (N_7194,N_2590,N_3256);
nor U7195 (N_7195,N_2624,N_4512);
nand U7196 (N_7196,N_3160,N_2807);
and U7197 (N_7197,N_2729,N_2667);
nor U7198 (N_7198,N_2633,N_4046);
nor U7199 (N_7199,N_3649,N_4877);
nor U7200 (N_7200,N_2929,N_3487);
or U7201 (N_7201,N_4255,N_4096);
nand U7202 (N_7202,N_4396,N_4824);
nor U7203 (N_7203,N_4587,N_3421);
nor U7204 (N_7204,N_2735,N_4414);
or U7205 (N_7205,N_2634,N_3179);
or U7206 (N_7206,N_3795,N_3143);
or U7207 (N_7207,N_4250,N_3299);
or U7208 (N_7208,N_4667,N_3957);
nand U7209 (N_7209,N_4466,N_4980);
nand U7210 (N_7210,N_3312,N_3616);
or U7211 (N_7211,N_3846,N_4275);
nand U7212 (N_7212,N_4854,N_4595);
and U7213 (N_7213,N_4190,N_2765);
and U7214 (N_7214,N_4343,N_3051);
nor U7215 (N_7215,N_3982,N_4184);
nand U7216 (N_7216,N_2563,N_3469);
or U7217 (N_7217,N_2993,N_4641);
or U7218 (N_7218,N_4619,N_3121);
or U7219 (N_7219,N_3138,N_4235);
and U7220 (N_7220,N_3691,N_2780);
nor U7221 (N_7221,N_4163,N_3191);
or U7222 (N_7222,N_4819,N_4057);
or U7223 (N_7223,N_3646,N_3686);
or U7224 (N_7224,N_4320,N_4749);
and U7225 (N_7225,N_3203,N_4652);
and U7226 (N_7226,N_4381,N_4266);
nor U7227 (N_7227,N_4415,N_4362);
nand U7228 (N_7228,N_2998,N_3068);
nor U7229 (N_7229,N_3522,N_3930);
and U7230 (N_7230,N_4007,N_2945);
nand U7231 (N_7231,N_3446,N_2994);
and U7232 (N_7232,N_3602,N_3220);
nand U7233 (N_7233,N_2527,N_3492);
nor U7234 (N_7234,N_4858,N_4559);
nand U7235 (N_7235,N_3882,N_4186);
and U7236 (N_7236,N_4547,N_4088);
nor U7237 (N_7237,N_2704,N_3563);
or U7238 (N_7238,N_3796,N_2931);
xnor U7239 (N_7239,N_4676,N_4435);
nor U7240 (N_7240,N_4876,N_4375);
nand U7241 (N_7241,N_4486,N_3308);
or U7242 (N_7242,N_4156,N_4593);
and U7243 (N_7243,N_2692,N_3568);
nor U7244 (N_7244,N_4444,N_2786);
xor U7245 (N_7245,N_3939,N_4964);
and U7246 (N_7246,N_2809,N_4107);
nand U7247 (N_7247,N_2567,N_4977);
nand U7248 (N_7248,N_3228,N_3041);
nand U7249 (N_7249,N_4080,N_3642);
and U7250 (N_7250,N_3022,N_4793);
nor U7251 (N_7251,N_3411,N_2539);
and U7252 (N_7252,N_3269,N_4949);
or U7253 (N_7253,N_4354,N_2862);
xor U7254 (N_7254,N_4771,N_3248);
and U7255 (N_7255,N_4219,N_2693);
nand U7256 (N_7256,N_4754,N_3587);
nand U7257 (N_7257,N_4244,N_2886);
and U7258 (N_7258,N_2681,N_4131);
xor U7259 (N_7259,N_3246,N_3031);
or U7260 (N_7260,N_3968,N_2823);
nand U7261 (N_7261,N_4465,N_3537);
nand U7262 (N_7262,N_3891,N_2762);
and U7263 (N_7263,N_2775,N_3178);
nor U7264 (N_7264,N_4926,N_4070);
or U7265 (N_7265,N_2897,N_3577);
nand U7266 (N_7266,N_3346,N_2845);
nor U7267 (N_7267,N_3054,N_4557);
nand U7268 (N_7268,N_3988,N_3071);
or U7269 (N_7269,N_4142,N_4438);
nand U7270 (N_7270,N_3575,N_4650);
and U7271 (N_7271,N_4235,N_3243);
nor U7272 (N_7272,N_2695,N_3413);
and U7273 (N_7273,N_3527,N_2791);
and U7274 (N_7274,N_3798,N_3893);
or U7275 (N_7275,N_3495,N_3983);
and U7276 (N_7276,N_3067,N_2889);
and U7277 (N_7277,N_2806,N_3032);
nand U7278 (N_7278,N_2831,N_4235);
nand U7279 (N_7279,N_3945,N_3559);
nor U7280 (N_7280,N_4087,N_4949);
nor U7281 (N_7281,N_4383,N_4478);
nand U7282 (N_7282,N_3947,N_3669);
or U7283 (N_7283,N_3063,N_3144);
nor U7284 (N_7284,N_3582,N_4431);
and U7285 (N_7285,N_4719,N_4095);
nand U7286 (N_7286,N_3384,N_3764);
and U7287 (N_7287,N_3272,N_4661);
and U7288 (N_7288,N_3324,N_3755);
xnor U7289 (N_7289,N_2787,N_4848);
or U7290 (N_7290,N_3699,N_3595);
or U7291 (N_7291,N_3440,N_3973);
and U7292 (N_7292,N_4631,N_4659);
nor U7293 (N_7293,N_4786,N_4037);
nand U7294 (N_7294,N_2510,N_2790);
nand U7295 (N_7295,N_4362,N_2557);
and U7296 (N_7296,N_2736,N_3561);
nor U7297 (N_7297,N_4993,N_3643);
nand U7298 (N_7298,N_2946,N_4046);
and U7299 (N_7299,N_4727,N_4776);
or U7300 (N_7300,N_2536,N_3373);
or U7301 (N_7301,N_3136,N_4753);
or U7302 (N_7302,N_2888,N_3974);
nor U7303 (N_7303,N_4949,N_3560);
or U7304 (N_7304,N_3769,N_3868);
or U7305 (N_7305,N_3920,N_3255);
nand U7306 (N_7306,N_4839,N_4379);
and U7307 (N_7307,N_2921,N_3349);
or U7308 (N_7308,N_3220,N_2971);
nor U7309 (N_7309,N_3431,N_4543);
and U7310 (N_7310,N_3285,N_3147);
and U7311 (N_7311,N_4940,N_4290);
nand U7312 (N_7312,N_2652,N_3984);
nor U7313 (N_7313,N_3430,N_3273);
and U7314 (N_7314,N_3796,N_2659);
nand U7315 (N_7315,N_4869,N_4058);
nand U7316 (N_7316,N_4507,N_2834);
or U7317 (N_7317,N_3584,N_3459);
nor U7318 (N_7318,N_4339,N_2633);
nand U7319 (N_7319,N_3750,N_3860);
and U7320 (N_7320,N_4405,N_4575);
nor U7321 (N_7321,N_2719,N_3499);
or U7322 (N_7322,N_3309,N_2874);
or U7323 (N_7323,N_4651,N_4865);
nor U7324 (N_7324,N_4323,N_4828);
or U7325 (N_7325,N_4574,N_3130);
nand U7326 (N_7326,N_3481,N_4593);
nand U7327 (N_7327,N_3908,N_4142);
and U7328 (N_7328,N_4498,N_4932);
nand U7329 (N_7329,N_4028,N_3682);
or U7330 (N_7330,N_3132,N_4028);
and U7331 (N_7331,N_3947,N_2576);
nand U7332 (N_7332,N_2516,N_3846);
and U7333 (N_7333,N_3634,N_2973);
nand U7334 (N_7334,N_4043,N_3034);
and U7335 (N_7335,N_4401,N_3897);
xor U7336 (N_7336,N_4070,N_4588);
and U7337 (N_7337,N_4847,N_3218);
or U7338 (N_7338,N_3815,N_4670);
and U7339 (N_7339,N_4015,N_3326);
nor U7340 (N_7340,N_2540,N_2807);
nand U7341 (N_7341,N_3886,N_3537);
or U7342 (N_7342,N_3840,N_3937);
or U7343 (N_7343,N_3341,N_3728);
nor U7344 (N_7344,N_2787,N_2966);
and U7345 (N_7345,N_3368,N_3310);
or U7346 (N_7346,N_3831,N_4798);
and U7347 (N_7347,N_3381,N_3165);
xor U7348 (N_7348,N_3753,N_3774);
and U7349 (N_7349,N_4564,N_3227);
nor U7350 (N_7350,N_4725,N_4131);
nand U7351 (N_7351,N_3830,N_3912);
nor U7352 (N_7352,N_2926,N_2558);
nor U7353 (N_7353,N_2739,N_3453);
and U7354 (N_7354,N_2880,N_4362);
or U7355 (N_7355,N_3678,N_2588);
nand U7356 (N_7356,N_4175,N_3342);
nor U7357 (N_7357,N_3424,N_3100);
or U7358 (N_7358,N_3928,N_4173);
nand U7359 (N_7359,N_3619,N_4424);
nand U7360 (N_7360,N_2636,N_4742);
and U7361 (N_7361,N_2746,N_4347);
xnor U7362 (N_7362,N_3306,N_3621);
or U7363 (N_7363,N_4312,N_4651);
nand U7364 (N_7364,N_3870,N_2934);
nand U7365 (N_7365,N_4257,N_3625);
nand U7366 (N_7366,N_4219,N_3285);
nor U7367 (N_7367,N_3400,N_4868);
or U7368 (N_7368,N_4200,N_4697);
nand U7369 (N_7369,N_3862,N_2944);
nand U7370 (N_7370,N_2767,N_4183);
nand U7371 (N_7371,N_3874,N_4682);
or U7372 (N_7372,N_4044,N_3516);
or U7373 (N_7373,N_4228,N_3009);
nand U7374 (N_7374,N_3864,N_4355);
nand U7375 (N_7375,N_3053,N_4985);
nand U7376 (N_7376,N_3850,N_4324);
and U7377 (N_7377,N_2772,N_3534);
nor U7378 (N_7378,N_2786,N_4823);
and U7379 (N_7379,N_4913,N_3490);
nor U7380 (N_7380,N_4156,N_4476);
or U7381 (N_7381,N_4423,N_4102);
nand U7382 (N_7382,N_4821,N_2889);
or U7383 (N_7383,N_4715,N_3008);
or U7384 (N_7384,N_4318,N_3308);
and U7385 (N_7385,N_4753,N_4367);
nor U7386 (N_7386,N_3517,N_3838);
nor U7387 (N_7387,N_2867,N_3627);
nor U7388 (N_7388,N_4308,N_4703);
nand U7389 (N_7389,N_4632,N_3275);
or U7390 (N_7390,N_3683,N_3756);
and U7391 (N_7391,N_4412,N_2809);
nand U7392 (N_7392,N_3034,N_2510);
nand U7393 (N_7393,N_3762,N_4004);
or U7394 (N_7394,N_3237,N_3455);
or U7395 (N_7395,N_3794,N_3679);
nor U7396 (N_7396,N_2706,N_4376);
and U7397 (N_7397,N_3932,N_3578);
and U7398 (N_7398,N_3676,N_4829);
nand U7399 (N_7399,N_4267,N_3717);
or U7400 (N_7400,N_4955,N_4934);
nand U7401 (N_7401,N_3879,N_4893);
or U7402 (N_7402,N_4443,N_4302);
xor U7403 (N_7403,N_3544,N_2592);
nand U7404 (N_7404,N_3882,N_4345);
and U7405 (N_7405,N_2961,N_3011);
and U7406 (N_7406,N_3422,N_4318);
and U7407 (N_7407,N_3406,N_3393);
and U7408 (N_7408,N_2581,N_3100);
nor U7409 (N_7409,N_4707,N_2911);
or U7410 (N_7410,N_4309,N_3754);
nand U7411 (N_7411,N_4491,N_3232);
nand U7412 (N_7412,N_2949,N_4553);
nand U7413 (N_7413,N_2943,N_2828);
and U7414 (N_7414,N_4832,N_3843);
nor U7415 (N_7415,N_3443,N_2653);
nor U7416 (N_7416,N_4592,N_3443);
nand U7417 (N_7417,N_3118,N_3641);
nor U7418 (N_7418,N_3085,N_4046);
nand U7419 (N_7419,N_3862,N_3347);
or U7420 (N_7420,N_4014,N_3094);
and U7421 (N_7421,N_3856,N_3186);
and U7422 (N_7422,N_3371,N_3779);
nor U7423 (N_7423,N_4593,N_4469);
or U7424 (N_7424,N_3774,N_4912);
or U7425 (N_7425,N_3419,N_3811);
nor U7426 (N_7426,N_4396,N_3925);
nor U7427 (N_7427,N_4782,N_2829);
nor U7428 (N_7428,N_4195,N_2694);
and U7429 (N_7429,N_3342,N_3481);
or U7430 (N_7430,N_2921,N_4914);
and U7431 (N_7431,N_2712,N_3757);
and U7432 (N_7432,N_3764,N_2628);
nand U7433 (N_7433,N_2611,N_3840);
nor U7434 (N_7434,N_2818,N_3084);
nand U7435 (N_7435,N_4986,N_4539);
or U7436 (N_7436,N_4815,N_2910);
xnor U7437 (N_7437,N_4757,N_3501);
and U7438 (N_7438,N_4611,N_4775);
nand U7439 (N_7439,N_3145,N_2959);
nand U7440 (N_7440,N_4217,N_3095);
and U7441 (N_7441,N_4384,N_4293);
and U7442 (N_7442,N_3109,N_4338);
nor U7443 (N_7443,N_3978,N_4762);
nand U7444 (N_7444,N_3604,N_2695);
nand U7445 (N_7445,N_3041,N_4831);
or U7446 (N_7446,N_2503,N_3732);
or U7447 (N_7447,N_3740,N_4614);
and U7448 (N_7448,N_3431,N_3338);
nor U7449 (N_7449,N_4076,N_3498);
nand U7450 (N_7450,N_4709,N_2521);
or U7451 (N_7451,N_3864,N_2633);
or U7452 (N_7452,N_3677,N_3214);
or U7453 (N_7453,N_2539,N_2602);
nand U7454 (N_7454,N_2818,N_4629);
and U7455 (N_7455,N_2587,N_3205);
nand U7456 (N_7456,N_2833,N_4000);
and U7457 (N_7457,N_3146,N_2826);
and U7458 (N_7458,N_4797,N_3706);
nand U7459 (N_7459,N_3964,N_4052);
or U7460 (N_7460,N_3543,N_3856);
nor U7461 (N_7461,N_3310,N_4348);
or U7462 (N_7462,N_4180,N_4524);
nor U7463 (N_7463,N_3436,N_3543);
nor U7464 (N_7464,N_2873,N_4991);
and U7465 (N_7465,N_4910,N_2967);
or U7466 (N_7466,N_4660,N_4566);
nand U7467 (N_7467,N_4076,N_3521);
nor U7468 (N_7468,N_3717,N_4055);
and U7469 (N_7469,N_4505,N_4350);
and U7470 (N_7470,N_4356,N_2636);
or U7471 (N_7471,N_4320,N_2632);
or U7472 (N_7472,N_4283,N_4257);
nand U7473 (N_7473,N_3368,N_3973);
and U7474 (N_7474,N_3640,N_3812);
and U7475 (N_7475,N_3331,N_3436);
and U7476 (N_7476,N_3562,N_3879);
and U7477 (N_7477,N_4836,N_3581);
or U7478 (N_7478,N_2581,N_4086);
and U7479 (N_7479,N_2878,N_4367);
xor U7480 (N_7480,N_2816,N_3446);
nand U7481 (N_7481,N_3829,N_4211);
or U7482 (N_7482,N_2891,N_2921);
or U7483 (N_7483,N_4014,N_4573);
nand U7484 (N_7484,N_3932,N_4868);
nand U7485 (N_7485,N_3185,N_2935);
nand U7486 (N_7486,N_4545,N_3765);
nor U7487 (N_7487,N_4986,N_4785);
or U7488 (N_7488,N_3748,N_4382);
or U7489 (N_7489,N_2608,N_4975);
nor U7490 (N_7490,N_4620,N_4133);
or U7491 (N_7491,N_3973,N_4636);
or U7492 (N_7492,N_4618,N_4510);
nand U7493 (N_7493,N_4089,N_2509);
nand U7494 (N_7494,N_2654,N_3689);
nand U7495 (N_7495,N_2659,N_2589);
xnor U7496 (N_7496,N_4300,N_3411);
or U7497 (N_7497,N_4683,N_3139);
or U7498 (N_7498,N_3408,N_4967);
nand U7499 (N_7499,N_4897,N_3807);
nand U7500 (N_7500,N_5511,N_5374);
nand U7501 (N_7501,N_6942,N_6614);
nor U7502 (N_7502,N_5873,N_6695);
and U7503 (N_7503,N_5618,N_6545);
nor U7504 (N_7504,N_6549,N_5451);
and U7505 (N_7505,N_6515,N_5611);
nor U7506 (N_7506,N_6211,N_7327);
or U7507 (N_7507,N_7286,N_6277);
nor U7508 (N_7508,N_6223,N_7044);
nand U7509 (N_7509,N_5169,N_5987);
or U7510 (N_7510,N_6326,N_6321);
nor U7511 (N_7511,N_6847,N_5978);
nor U7512 (N_7512,N_5926,N_6865);
nand U7513 (N_7513,N_7292,N_6180);
xor U7514 (N_7514,N_6711,N_5999);
nor U7515 (N_7515,N_7431,N_6876);
nand U7516 (N_7516,N_7251,N_7269);
nand U7517 (N_7517,N_5691,N_6388);
nand U7518 (N_7518,N_5966,N_5006);
nand U7519 (N_7519,N_6871,N_6690);
nand U7520 (N_7520,N_7266,N_5577);
nand U7521 (N_7521,N_7092,N_7473);
and U7522 (N_7522,N_5269,N_7201);
and U7523 (N_7523,N_6990,N_5233);
and U7524 (N_7524,N_5363,N_5876);
nor U7525 (N_7525,N_5840,N_5587);
or U7526 (N_7526,N_5834,N_7130);
or U7527 (N_7527,N_5854,N_5984);
or U7528 (N_7528,N_5317,N_6243);
nand U7529 (N_7529,N_7204,N_7028);
and U7530 (N_7530,N_6429,N_7448);
or U7531 (N_7531,N_5303,N_7158);
nor U7532 (N_7532,N_7335,N_6107);
and U7533 (N_7533,N_6616,N_5261);
or U7534 (N_7534,N_5575,N_6874);
nor U7535 (N_7535,N_7391,N_6664);
or U7536 (N_7536,N_6441,N_5730);
nor U7537 (N_7537,N_7396,N_5604);
nand U7538 (N_7538,N_7265,N_6597);
nor U7539 (N_7539,N_6879,N_6040);
and U7540 (N_7540,N_6662,N_5726);
and U7541 (N_7541,N_7351,N_6094);
and U7542 (N_7542,N_7123,N_7021);
nand U7543 (N_7543,N_6820,N_5260);
nand U7544 (N_7544,N_7227,N_5662);
nor U7545 (N_7545,N_7042,N_5743);
nor U7546 (N_7546,N_7104,N_5147);
and U7547 (N_7547,N_5073,N_6643);
xnor U7548 (N_7548,N_5150,N_6284);
or U7549 (N_7549,N_7062,N_7005);
and U7550 (N_7550,N_7152,N_5722);
or U7551 (N_7551,N_5787,N_5217);
nand U7552 (N_7552,N_6906,N_7154);
nand U7553 (N_7553,N_7127,N_7187);
and U7554 (N_7554,N_6862,N_5737);
nand U7555 (N_7555,N_6060,N_6057);
and U7556 (N_7556,N_5750,N_5461);
and U7557 (N_7557,N_7293,N_5431);
nor U7558 (N_7558,N_6384,N_7410);
nor U7559 (N_7559,N_6335,N_5181);
nor U7560 (N_7560,N_5045,N_5226);
nand U7561 (N_7561,N_6734,N_5323);
or U7562 (N_7562,N_5001,N_6934);
and U7563 (N_7563,N_5422,N_7339);
nand U7564 (N_7564,N_5000,N_5328);
or U7565 (N_7565,N_5453,N_5799);
nand U7566 (N_7566,N_6710,N_5128);
nor U7567 (N_7567,N_7031,N_6835);
and U7568 (N_7568,N_5164,N_5814);
and U7569 (N_7569,N_5078,N_6986);
and U7570 (N_7570,N_5187,N_7482);
nor U7571 (N_7571,N_6891,N_5507);
nor U7572 (N_7572,N_6632,N_6777);
or U7573 (N_7573,N_6880,N_5403);
nand U7574 (N_7574,N_6315,N_6764);
or U7575 (N_7575,N_7106,N_5468);
nand U7576 (N_7576,N_6207,N_6684);
and U7577 (N_7577,N_6016,N_6895);
nor U7578 (N_7578,N_5325,N_7372);
and U7579 (N_7579,N_5048,N_5306);
or U7580 (N_7580,N_6319,N_6945);
or U7581 (N_7581,N_6167,N_7144);
and U7582 (N_7582,N_5254,N_6842);
and U7583 (N_7583,N_5658,N_6964);
or U7584 (N_7584,N_5230,N_5247);
nor U7585 (N_7585,N_5767,N_7310);
nor U7586 (N_7586,N_6300,N_6754);
or U7587 (N_7587,N_7128,N_6355);
nand U7588 (N_7588,N_5483,N_5982);
and U7589 (N_7589,N_5019,N_7371);
nor U7590 (N_7590,N_7386,N_6745);
or U7591 (N_7591,N_7313,N_5257);
nand U7592 (N_7592,N_6806,N_6136);
nor U7593 (N_7593,N_5883,N_7132);
and U7594 (N_7594,N_6605,N_5887);
or U7595 (N_7595,N_5588,N_5253);
nand U7596 (N_7596,N_5290,N_6487);
or U7597 (N_7597,N_6323,N_5344);
nor U7598 (N_7598,N_5892,N_6656);
nor U7599 (N_7599,N_7491,N_7136);
or U7600 (N_7600,N_6314,N_5015);
nor U7601 (N_7601,N_7475,N_5139);
or U7602 (N_7602,N_6255,N_5090);
xor U7603 (N_7603,N_7043,N_6814);
nor U7604 (N_7604,N_7048,N_5042);
nand U7605 (N_7605,N_6125,N_5039);
or U7606 (N_7606,N_6655,N_5221);
and U7607 (N_7607,N_5336,N_5327);
and U7608 (N_7608,N_5936,N_5036);
and U7609 (N_7609,N_5003,N_6663);
and U7610 (N_7610,N_5734,N_6970);
and U7611 (N_7611,N_5439,N_6260);
nand U7612 (N_7612,N_7202,N_7484);
or U7613 (N_7613,N_5846,N_5447);
or U7614 (N_7614,N_5002,N_6090);
and U7615 (N_7615,N_5560,N_5717);
and U7616 (N_7616,N_7329,N_6619);
and U7617 (N_7617,N_7037,N_6088);
or U7618 (N_7618,N_6369,N_6360);
or U7619 (N_7619,N_7014,N_5277);
nor U7620 (N_7620,N_5410,N_5272);
or U7621 (N_7621,N_6095,N_6160);
and U7622 (N_7622,N_6954,N_5915);
and U7623 (N_7623,N_5592,N_6482);
nand U7624 (N_7624,N_6624,N_5478);
nand U7625 (N_7625,N_6770,N_7171);
or U7626 (N_7626,N_6784,N_6503);
nand U7627 (N_7627,N_5030,N_5929);
or U7628 (N_7628,N_7452,N_6174);
nor U7629 (N_7629,N_5205,N_6043);
nand U7630 (N_7630,N_5491,N_6254);
or U7631 (N_7631,N_6238,N_6123);
or U7632 (N_7632,N_6554,N_6608);
nor U7633 (N_7633,N_7065,N_6933);
nor U7634 (N_7634,N_5650,N_7487);
nand U7635 (N_7635,N_5867,N_7443);
nor U7636 (N_7636,N_6866,N_7451);
or U7637 (N_7637,N_5096,N_6112);
nand U7638 (N_7638,N_7141,N_5894);
nand U7639 (N_7639,N_6206,N_6885);
or U7640 (N_7640,N_5946,N_5416);
and U7641 (N_7641,N_5258,N_6807);
and U7642 (N_7642,N_7301,N_7314);
and U7643 (N_7643,N_5038,N_7343);
nand U7644 (N_7644,N_6298,N_7026);
or U7645 (N_7645,N_6898,N_6937);
or U7646 (N_7646,N_5341,N_5446);
nor U7647 (N_7647,N_7089,N_7226);
nand U7648 (N_7648,N_5681,N_5584);
or U7649 (N_7649,N_5084,N_6960);
and U7650 (N_7650,N_6737,N_7178);
nand U7651 (N_7651,N_5830,N_6020);
and U7652 (N_7652,N_5525,N_6295);
and U7653 (N_7653,N_6499,N_5527);
and U7654 (N_7654,N_6133,N_5660);
nor U7655 (N_7655,N_7366,N_7002);
or U7656 (N_7656,N_5385,N_5158);
nor U7657 (N_7657,N_7097,N_6634);
nand U7658 (N_7658,N_5295,N_6214);
and U7659 (N_7659,N_5364,N_6375);
or U7660 (N_7660,N_5063,N_5859);
or U7661 (N_7661,N_7462,N_6796);
and U7662 (N_7662,N_6542,N_6037);
nand U7663 (N_7663,N_5377,N_5811);
nor U7664 (N_7664,N_7398,N_6200);
xor U7665 (N_7665,N_5273,N_6669);
nand U7666 (N_7666,N_6069,N_5718);
and U7667 (N_7667,N_6956,N_6025);
or U7668 (N_7668,N_6142,N_5119);
or U7669 (N_7669,N_5842,N_5352);
or U7670 (N_7670,N_6989,N_6309);
nand U7671 (N_7671,N_6687,N_7342);
and U7672 (N_7672,N_7375,N_6121);
nand U7673 (N_7673,N_6537,N_7352);
or U7674 (N_7674,N_6002,N_6132);
nand U7675 (N_7675,N_6618,N_5764);
nor U7676 (N_7676,N_7060,N_5081);
and U7677 (N_7677,N_6638,N_5968);
and U7678 (N_7678,N_5311,N_5945);
or U7679 (N_7679,N_5329,N_6120);
or U7680 (N_7680,N_6282,N_6547);
and U7681 (N_7681,N_6527,N_6899);
nand U7682 (N_7682,N_7194,N_7019);
and U7683 (N_7683,N_6491,N_7205);
nand U7684 (N_7684,N_5398,N_7485);
nor U7685 (N_7685,N_6631,N_6299);
and U7686 (N_7686,N_5508,N_5499);
nor U7687 (N_7687,N_5298,N_5761);
nor U7688 (N_7688,N_5490,N_7453);
or U7689 (N_7689,N_5503,N_7274);
nand U7690 (N_7690,N_5620,N_7294);
nor U7691 (N_7691,N_7457,N_7146);
or U7692 (N_7692,N_5977,N_6803);
nor U7693 (N_7693,N_6209,N_7017);
and U7694 (N_7694,N_6595,N_5528);
nor U7695 (N_7695,N_6840,N_6253);
or U7696 (N_7696,N_6271,N_6064);
nand U7697 (N_7697,N_6078,N_7338);
nand U7698 (N_7698,N_6567,N_5095);
nand U7699 (N_7699,N_5760,N_5184);
nor U7700 (N_7700,N_6520,N_7032);
and U7701 (N_7701,N_5682,N_5808);
or U7702 (N_7702,N_6034,N_5395);
nor U7703 (N_7703,N_5440,N_6715);
nor U7704 (N_7704,N_5489,N_5732);
and U7705 (N_7705,N_5674,N_5635);
or U7706 (N_7706,N_6392,N_5880);
or U7707 (N_7707,N_5513,N_7221);
and U7708 (N_7708,N_6600,N_6359);
and U7709 (N_7709,N_5388,N_6403);
nor U7710 (N_7710,N_5529,N_6333);
or U7711 (N_7711,N_6424,N_6752);
or U7712 (N_7712,N_7413,N_6526);
or U7713 (N_7713,N_6967,N_6501);
and U7714 (N_7714,N_6483,N_5774);
and U7715 (N_7715,N_6158,N_6773);
nand U7716 (N_7716,N_6747,N_5343);
and U7717 (N_7717,N_5242,N_7206);
xnor U7718 (N_7718,N_5692,N_7216);
and U7719 (N_7719,N_5861,N_7483);
nand U7720 (N_7720,N_6717,N_5308);
nor U7721 (N_7721,N_6642,N_6370);
and U7722 (N_7722,N_6912,N_6210);
or U7723 (N_7723,N_5127,N_5467);
or U7724 (N_7724,N_5835,N_5871);
nand U7725 (N_7725,N_6026,N_6704);
and U7726 (N_7726,N_6406,N_6268);
nand U7727 (N_7727,N_6872,N_5683);
nand U7728 (N_7728,N_5536,N_5930);
or U7729 (N_7729,N_7155,N_7250);
nor U7730 (N_7730,N_6994,N_7015);
and U7731 (N_7731,N_5083,N_6224);
nor U7732 (N_7732,N_5051,N_6248);
nand U7733 (N_7733,N_5237,N_6193);
nor U7734 (N_7734,N_6725,N_6155);
nand U7735 (N_7735,N_5195,N_6412);
nand U7736 (N_7736,N_5183,N_5735);
or U7737 (N_7737,N_6466,N_6903);
or U7738 (N_7738,N_6336,N_5235);
or U7739 (N_7739,N_6213,N_6529);
or U7740 (N_7740,N_5879,N_7403);
and U7741 (N_7741,N_6073,N_5442);
and U7742 (N_7742,N_6053,N_5010);
nand U7743 (N_7743,N_6888,N_6293);
nor U7744 (N_7744,N_5839,N_6163);
nor U7745 (N_7745,N_6042,N_6505);
and U7746 (N_7746,N_5345,N_5408);
nand U7747 (N_7747,N_5309,N_6477);
nand U7748 (N_7748,N_5991,N_5227);
or U7749 (N_7749,N_6969,N_6910);
and U7750 (N_7750,N_7198,N_6237);
or U7751 (N_7751,N_7086,N_5144);
nor U7752 (N_7752,N_6489,N_5551);
nand U7753 (N_7753,N_5785,N_7302);
nor U7754 (N_7754,N_6099,N_7497);
nor U7755 (N_7755,N_7464,N_5379);
nor U7756 (N_7756,N_7259,N_6023);
and U7757 (N_7757,N_6114,N_6003);
nor U7758 (N_7758,N_6178,N_6444);
nor U7759 (N_7759,N_6636,N_5877);
nor U7760 (N_7760,N_5118,N_5104);
xor U7761 (N_7761,N_5625,N_7090);
and U7762 (N_7762,N_5980,N_5745);
nand U7763 (N_7763,N_5436,N_5292);
and U7764 (N_7764,N_6386,N_5054);
and U7765 (N_7765,N_6758,N_6781);
xnor U7766 (N_7766,N_5069,N_5133);
or U7767 (N_7767,N_7181,N_6014);
and U7768 (N_7768,N_7476,N_6630);
nor U7769 (N_7769,N_6522,N_7437);
or U7770 (N_7770,N_6726,N_5781);
nor U7771 (N_7771,N_7241,N_5220);
nor U7772 (N_7772,N_5448,N_6301);
nand U7773 (N_7773,N_5189,N_5917);
or U7774 (N_7774,N_6275,N_6379);
or U7775 (N_7775,N_5752,N_6322);
and U7776 (N_7776,N_5878,N_6571);
nor U7777 (N_7777,N_6346,N_7047);
nor U7778 (N_7778,N_6024,N_6744);
and U7779 (N_7779,N_6718,N_6154);
nor U7780 (N_7780,N_5178,N_6182);
nor U7781 (N_7781,N_5032,N_5517);
nand U7782 (N_7782,N_6714,N_5238);
nor U7783 (N_7783,N_7492,N_5041);
nor U7784 (N_7784,N_5202,N_7197);
and U7785 (N_7785,N_5893,N_6189);
nand U7786 (N_7786,N_6048,N_6805);
nand U7787 (N_7787,N_5070,N_6640);
nor U7788 (N_7788,N_7046,N_6713);
nor U7789 (N_7789,N_6348,N_6004);
nor U7790 (N_7790,N_7256,N_6201);
and U7791 (N_7791,N_5637,N_6497);
nor U7792 (N_7792,N_5291,N_6408);
and U7793 (N_7793,N_6813,N_6860);
nand U7794 (N_7794,N_6378,N_7298);
or U7795 (N_7795,N_5610,N_5225);
nor U7796 (N_7796,N_7125,N_5207);
nor U7797 (N_7797,N_5018,N_6649);
nor U7798 (N_7798,N_5182,N_5541);
and U7799 (N_7799,N_5145,N_6161);
nand U7800 (N_7800,N_6996,N_5952);
or U7801 (N_7801,N_5049,N_7499);
and U7802 (N_7802,N_6144,N_6918);
nand U7803 (N_7803,N_6347,N_5603);
nand U7804 (N_7804,N_6776,N_5149);
nor U7805 (N_7805,N_6442,N_6220);
nor U7806 (N_7806,N_6173,N_5697);
or U7807 (N_7807,N_6908,N_6476);
nand U7808 (N_7808,N_5004,N_5413);
nor U7809 (N_7809,N_6028,N_6274);
nor U7810 (N_7810,N_7049,N_5805);
nand U7811 (N_7811,N_5881,N_7107);
or U7812 (N_7812,N_7036,N_6997);
and U7813 (N_7813,N_6894,N_6485);
or U7814 (N_7814,N_6680,N_6637);
and U7815 (N_7815,N_6416,N_5969);
nor U7816 (N_7816,N_6881,N_5365);
nor U7817 (N_7817,N_7461,N_7323);
and U7818 (N_7818,N_7285,N_5792);
nand U7819 (N_7819,N_5671,N_6130);
and U7820 (N_7820,N_6588,N_6976);
and U7821 (N_7821,N_7405,N_7248);
nand U7822 (N_7822,N_5400,N_5862);
nand U7823 (N_7823,N_6286,N_6755);
nand U7824 (N_7824,N_5473,N_5330);
and U7825 (N_7825,N_6815,N_7385);
nand U7826 (N_7826,N_6399,N_6626);
and U7827 (N_7827,N_5535,N_5522);
nand U7828 (N_7828,N_5193,N_5652);
nand U7829 (N_7829,N_5627,N_6801);
nand U7830 (N_7830,N_7118,N_5825);
or U7831 (N_7831,N_5455,N_7460);
xnor U7832 (N_7832,N_5293,N_5180);
or U7833 (N_7833,N_7365,N_5066);
nor U7834 (N_7834,N_7361,N_7455);
and U7835 (N_7835,N_5602,N_6306);
nand U7836 (N_7836,N_7084,N_7219);
or U7837 (N_7837,N_5143,N_6615);
xnor U7838 (N_7838,N_5775,N_7394);
nor U7839 (N_7839,N_5838,N_7433);
or U7840 (N_7840,N_6905,N_7291);
and U7841 (N_7841,N_6580,N_6204);
and U7842 (N_7842,N_6904,N_5131);
nand U7843 (N_7843,N_6821,N_7055);
or U7844 (N_7844,N_5386,N_6592);
nand U7845 (N_7845,N_6622,N_6312);
and U7846 (N_7846,N_7126,N_6143);
nor U7847 (N_7847,N_7168,N_6019);
and U7848 (N_7848,N_6953,N_6682);
nor U7849 (N_7849,N_6457,N_6741);
or U7850 (N_7850,N_6096,N_6109);
nand U7851 (N_7851,N_5537,N_5393);
and U7852 (N_7852,N_5219,N_5313);
nor U7853 (N_7853,N_7209,N_6665);
and U7854 (N_7854,N_5411,N_7273);
nand U7855 (N_7855,N_5810,N_6766);
or U7856 (N_7856,N_5112,N_6454);
nor U7857 (N_7857,N_5074,N_5266);
or U7858 (N_7858,N_6500,N_7387);
nor U7859 (N_7859,N_5673,N_5705);
nand U7860 (N_7860,N_5462,N_6859);
and U7861 (N_7861,N_6077,N_5776);
nand U7862 (N_7862,N_6395,N_6443);
and U7863 (N_7863,N_6495,N_7199);
nor U7864 (N_7864,N_6239,N_5502);
or U7865 (N_7865,N_5639,N_5472);
nor U7866 (N_7866,N_5702,N_5744);
or U7867 (N_7867,N_5368,N_6550);
nor U7868 (N_7868,N_6971,N_7077);
nor U7869 (N_7869,N_6463,N_5264);
nor U7870 (N_7870,N_5210,N_5552);
nor U7871 (N_7871,N_5259,N_6291);
nand U7872 (N_7872,N_6452,N_5950);
or U7873 (N_7873,N_6707,N_6533);
and U7874 (N_7874,N_7353,N_5943);
nor U7875 (N_7875,N_5616,N_6345);
and U7876 (N_7876,N_6134,N_6594);
and U7877 (N_7877,N_7052,N_7010);
or U7878 (N_7878,N_7260,N_6846);
and U7879 (N_7879,N_6496,N_7271);
nand U7880 (N_7880,N_5695,N_6790);
or U7881 (N_7881,N_6011,N_6407);
and U7882 (N_7882,N_5457,N_6426);
and U7883 (N_7883,N_6599,N_7378);
nand U7884 (N_7884,N_6074,N_6930);
nand U7885 (N_7885,N_6218,N_7172);
nor U7886 (N_7886,N_7493,N_7196);
nor U7887 (N_7887,N_6892,N_7306);
nand U7888 (N_7888,N_5340,N_6516);
or U7889 (N_7889,N_7167,N_5392);
nand U7890 (N_7890,N_6280,N_6620);
nand U7891 (N_7891,N_5017,N_5645);
or U7892 (N_7892,N_5322,N_5800);
and U7893 (N_7893,N_6697,N_6196);
and U7894 (N_7894,N_6063,N_5085);
nor U7895 (N_7895,N_7442,N_7316);
nor U7896 (N_7896,N_6798,N_7094);
or U7897 (N_7897,N_7428,N_6514);
or U7898 (N_7898,N_5863,N_5741);
nand U7899 (N_7899,N_5141,N_5729);
or U7900 (N_7900,N_5583,N_7064);
nor U7901 (N_7901,N_6007,N_5086);
and U7902 (N_7902,N_5476,N_7389);
nand U7903 (N_7903,N_5585,N_7432);
and U7904 (N_7904,N_6907,N_5449);
or U7905 (N_7905,N_6445,N_6558);
nor U7906 (N_7906,N_6944,N_7018);
and U7907 (N_7907,N_6356,N_7025);
nor U7908 (N_7908,N_5044,N_6249);
or U7909 (N_7909,N_5430,N_6913);
nor U7910 (N_7910,N_5990,N_5464);
or U7911 (N_7911,N_7355,N_6297);
nand U7912 (N_7912,N_7082,N_6458);
nor U7913 (N_7913,N_5614,N_6749);
or U7914 (N_7914,N_5704,N_5031);
nand U7915 (N_7915,N_7217,N_7495);
nor U7916 (N_7916,N_7467,N_6968);
xor U7917 (N_7917,N_7284,N_5672);
nand U7918 (N_7918,N_5142,N_6357);
nand U7919 (N_7919,N_6082,N_7376);
nor U7920 (N_7920,N_7406,N_7423);
nor U7921 (N_7921,N_7169,N_5828);
nor U7922 (N_7922,N_5094,N_5716);
nand U7923 (N_7923,N_5168,N_6941);
or U7924 (N_7924,N_7441,N_5655);
nand U7925 (N_7925,N_6987,N_7332);
nand U7926 (N_7926,N_6308,N_5240);
and U7927 (N_7927,N_5299,N_5882);
and U7928 (N_7928,N_7268,N_5494);
nor U7929 (N_7929,N_5435,N_5140);
nor U7930 (N_7930,N_7034,N_6231);
and U7931 (N_7931,N_5832,N_7417);
nor U7932 (N_7932,N_6861,N_5562);
or U7933 (N_7933,N_6674,N_5179);
nor U7934 (N_7934,N_5441,N_6041);
nand U7935 (N_7935,N_5406,N_5617);
or U7936 (N_7936,N_6310,N_6389);
or U7937 (N_7937,N_5232,N_6760);
nand U7938 (N_7938,N_5058,N_6508);
nand U7939 (N_7939,N_6393,N_5263);
or U7940 (N_7940,N_6625,N_6320);
xnor U7941 (N_7941,N_7363,N_6118);
nand U7942 (N_7942,N_5394,N_6411);
nor U7943 (N_7943,N_6117,N_7211);
or U7944 (N_7944,N_5504,N_6546);
nor U7945 (N_7945,N_6948,N_6678);
nor U7946 (N_7946,N_6822,N_7496);
nor U7947 (N_7947,N_5381,N_6681);
and U7948 (N_7948,N_6113,N_5668);
xnor U7949 (N_7949,N_5715,N_6490);
and U7950 (N_7950,N_7192,N_5901);
and U7951 (N_7951,N_5712,N_6138);
nor U7952 (N_7952,N_5985,N_5474);
and U7953 (N_7953,N_6106,N_6606);
nor U7954 (N_7954,N_5278,N_5791);
or U7955 (N_7955,N_6676,N_6601);
nor U7956 (N_7956,N_7072,N_5523);
nor U7957 (N_7957,N_7232,N_6473);
and U7958 (N_7958,N_7345,N_6799);
nor U7959 (N_7959,N_5539,N_5068);
or U7960 (N_7960,N_6092,N_7066);
nand U7961 (N_7961,N_6165,N_6650);
and U7962 (N_7962,N_5818,N_5819);
nand U7963 (N_7963,N_6528,N_6050);
and U7964 (N_7964,N_6172,N_5955);
nand U7965 (N_7965,N_6363,N_6984);
and U7966 (N_7966,N_5699,N_6591);
and U7967 (N_7967,N_7304,N_5497);
and U7968 (N_7968,N_5564,N_6827);
nand U7969 (N_7969,N_7373,N_6602);
nand U7970 (N_7970,N_6938,N_5807);
and U7971 (N_7971,N_5275,N_5763);
nand U7972 (N_7972,N_5103,N_5559);
nor U7973 (N_7973,N_5013,N_5157);
or U7974 (N_7974,N_7145,N_6985);
and U7975 (N_7975,N_5318,N_5097);
or U7976 (N_7976,N_6148,N_6437);
or U7977 (N_7977,N_6646,N_5572);
and U7978 (N_7978,N_6877,N_6762);
nand U7979 (N_7979,N_6509,N_6022);
nand U7980 (N_7980,N_5209,N_5107);
nor U7981 (N_7981,N_5109,N_5267);
nand U7982 (N_7982,N_5664,N_5900);
nand U7983 (N_7983,N_6139,N_7098);
nor U7984 (N_7984,N_5475,N_6828);
or U7985 (N_7985,N_6573,N_6919);
nand U7986 (N_7986,N_5126,N_5850);
nand U7987 (N_7987,N_5029,N_5059);
nor U7988 (N_7988,N_6818,N_6839);
and U7989 (N_7989,N_7357,N_6285);
nand U7990 (N_7990,N_6791,N_5115);
and U7991 (N_7991,N_6787,N_5007);
or U7992 (N_7992,N_7262,N_5927);
nor U7993 (N_7993,N_6612,N_6332);
nor U7994 (N_7994,N_7380,N_5615);
nand U7995 (N_7995,N_7296,N_7390);
and U7996 (N_7996,N_7382,N_7057);
and U7997 (N_7997,N_5279,N_7008);
nand U7998 (N_7998,N_5953,N_7013);
nor U7999 (N_7999,N_5137,N_6883);
nor U8000 (N_8000,N_5480,N_5937);
and U8001 (N_8001,N_5315,N_7102);
and U8002 (N_8002,N_7307,N_7312);
nor U8003 (N_8003,N_6823,N_6551);
nor U8004 (N_8004,N_7012,N_7024);
or U8005 (N_8005,N_5353,N_6661);
nand U8006 (N_8006,N_5907,N_6893);
or U8007 (N_8007,N_7305,N_5573);
nor U8008 (N_8008,N_6519,N_7225);
nand U8009 (N_8009,N_7237,N_6140);
and U8010 (N_8010,N_5407,N_6977);
nor U8011 (N_8011,N_5922,N_7151);
nor U8012 (N_8012,N_6738,N_5111);
and U8013 (N_8013,N_5459,N_6763);
nor U8014 (N_8014,N_5548,N_5708);
nor U8015 (N_8015,N_7157,N_6447);
nand U8016 (N_8016,N_6152,N_7020);
xnor U8017 (N_8017,N_5338,N_5797);
and U8018 (N_8018,N_7139,N_6973);
and U8019 (N_8019,N_7040,N_6205);
or U8020 (N_8020,N_6598,N_5098);
nor U8021 (N_8021,N_5228,N_6383);
nand U8022 (N_8022,N_5771,N_7009);
and U8023 (N_8023,N_7319,N_5852);
or U8024 (N_8024,N_6236,N_7477);
nand U8025 (N_8025,N_6617,N_5721);
nor U8026 (N_8026,N_6400,N_6225);
nand U8027 (N_8027,N_7297,N_5890);
or U8028 (N_8028,N_7054,N_5727);
nor U8029 (N_8029,N_6721,N_7244);
or U8030 (N_8030,N_6156,N_5872);
nor U8031 (N_8031,N_5420,N_7404);
xnor U8032 (N_8032,N_5134,N_5638);
or U8033 (N_8033,N_6838,N_7137);
and U8034 (N_8034,N_5823,N_5809);
nor U8035 (N_8035,N_6890,N_6965);
nand U8036 (N_8036,N_5035,N_6208);
and U8037 (N_8037,N_7395,N_7222);
nand U8038 (N_8038,N_6812,N_7220);
or U8039 (N_8039,N_5376,N_7001);
and U8040 (N_8040,N_5661,N_6353);
and U8041 (N_8041,N_7401,N_6778);
and U8042 (N_8042,N_5864,N_6584);
nand U8043 (N_8043,N_7050,N_6263);
and U8044 (N_8044,N_7238,N_5912);
and U8045 (N_8045,N_7276,N_6826);
nand U8046 (N_8046,N_6469,N_5989);
nor U8047 (N_8047,N_7213,N_5153);
xnor U8048 (N_8048,N_6045,N_5798);
and U8049 (N_8049,N_5738,N_6267);
and U8050 (N_8050,N_6451,N_5689);
nand U8051 (N_8051,N_6867,N_7224);
nand U8052 (N_8052,N_5803,N_6170);
nor U8053 (N_8053,N_5324,N_5961);
nor U8054 (N_8054,N_6493,N_5064);
or U8055 (N_8055,N_6972,N_6951);
and U8056 (N_8056,N_7346,N_6334);
nand U8057 (N_8057,N_6484,N_5680);
nor U8058 (N_8058,N_5331,N_5428);
and U8059 (N_8059,N_6572,N_5065);
or U8060 (N_8060,N_7470,N_5486);
and U8061 (N_8061,N_7140,N_5091);
xnor U8062 (N_8062,N_5780,N_5556);
and U8063 (N_8063,N_5813,N_6756);
nand U8064 (N_8064,N_6868,N_5022);
and U8065 (N_8065,N_5117,N_5185);
or U8066 (N_8066,N_7325,N_7180);
nand U8067 (N_8067,N_6351,N_6974);
nor U8068 (N_8068,N_7096,N_6563);
nor U8069 (N_8069,N_5773,N_6185);
and U8070 (N_8070,N_5914,N_5283);
nor U8071 (N_8071,N_5579,N_5634);
nand U8072 (N_8072,N_5895,N_5021);
nand U8073 (N_8073,N_5762,N_5510);
and U8074 (N_8074,N_7191,N_6510);
and U8075 (N_8075,N_5768,N_6448);
and U8076 (N_8076,N_5700,N_7234);
nor U8077 (N_8077,N_7023,N_5362);
or U8078 (N_8078,N_6902,N_5747);
and U8079 (N_8079,N_6052,N_6012);
and U8080 (N_8080,N_5076,N_5108);
nand U8081 (N_8081,N_6853,N_6504);
nor U8082 (N_8082,N_5820,N_5518);
nor U8083 (N_8083,N_7480,N_6792);
nor U8084 (N_8084,N_5686,N_6819);
nand U8085 (N_8085,N_5897,N_5983);
nor U8086 (N_8086,N_7182,N_5597);
and U8087 (N_8087,N_5204,N_6647);
and U8088 (N_8088,N_6049,N_5199);
nor U8089 (N_8089,N_5632,N_5919);
nor U8090 (N_8090,N_6742,N_5728);
nand U8091 (N_8091,N_6186,N_5008);
nor U8092 (N_8092,N_5731,N_5101);
and U8093 (N_8093,N_5628,N_6540);
or U8094 (N_8094,N_5703,N_6759);
nor U8095 (N_8095,N_6376,N_7478);
and U8096 (N_8096,N_5793,N_6667);
and U8097 (N_8097,N_6513,N_5429);
or U8098 (N_8098,N_6044,N_6771);
nand U8099 (N_8099,N_5498,N_5815);
xor U8100 (N_8100,N_6410,N_7203);
nand U8101 (N_8101,N_5262,N_5057);
nand U8102 (N_8102,N_6946,N_7112);
or U8103 (N_8103,N_6330,N_5866);
nand U8104 (N_8104,N_5595,N_5976);
or U8105 (N_8105,N_6978,N_7035);
and U8106 (N_8106,N_7341,N_5460);
or U8107 (N_8107,N_7027,N_5171);
nor U8108 (N_8108,N_6212,N_7195);
or U8109 (N_8109,N_5921,N_7162);
nand U8110 (N_8110,N_7295,N_7113);
or U8111 (N_8111,N_5934,N_5294);
nand U8112 (N_8112,N_5357,N_6849);
and U8113 (N_8113,N_6732,N_6864);
or U8114 (N_8114,N_6350,N_6922);
nand U8115 (N_8115,N_6365,N_5623);
nand U8116 (N_8116,N_6679,N_6425);
and U8117 (N_8117,N_5174,N_6492);
nand U8118 (N_8118,N_7223,N_5896);
nor U8119 (N_8119,N_5212,N_6418);
nor U8120 (N_8120,N_7458,N_7481);
and U8121 (N_8121,N_6401,N_6164);
or U8122 (N_8122,N_6963,N_5028);
and U8123 (N_8123,N_5709,N_6845);
or U8124 (N_8124,N_5201,N_5544);
or U8125 (N_8125,N_7280,N_5037);
nand U8126 (N_8126,N_6992,N_6195);
or U8127 (N_8127,N_6349,N_6438);
nand U8128 (N_8128,N_5116,N_5928);
or U8129 (N_8129,N_7073,N_5740);
nor U8130 (N_8130,N_5102,N_5710);
and U8131 (N_8131,N_7445,N_5214);
and U8132 (N_8132,N_6887,N_6258);
nand U8133 (N_8133,N_6980,N_6067);
nand U8134 (N_8134,N_7421,N_5888);
nand U8135 (N_8135,N_6431,N_7088);
nand U8136 (N_8136,N_6241,N_5642);
nand U8137 (N_8137,N_5391,N_6900);
or U8138 (N_8138,N_6317,N_5995);
or U8139 (N_8139,N_6920,N_6623);
or U8140 (N_8140,N_6449,N_6229);
and U8141 (N_8141,N_6478,N_6290);
nor U8142 (N_8142,N_5444,N_6135);
nand U8143 (N_8143,N_5482,N_6372);
nand U8144 (N_8144,N_6076,N_6080);
nor U8145 (N_8145,N_7068,N_6583);
and U8146 (N_8146,N_5817,N_6047);
nor U8147 (N_8147,N_7184,N_5166);
nor U8148 (N_8148,N_5152,N_5733);
or U8149 (N_8149,N_5748,N_6786);
and U8150 (N_8150,N_7108,N_6103);
nor U8151 (N_8151,N_6396,N_6830);
nand U8152 (N_8152,N_5387,N_5821);
nor U8153 (N_8153,N_7183,N_6327);
and U8154 (N_8154,N_5337,N_5114);
xnor U8155 (N_8155,N_6785,N_6943);
or U8156 (N_8156,N_6541,N_6470);
nand U8157 (N_8157,N_7114,N_6228);
or U8158 (N_8158,N_5175,N_6761);
nand U8159 (N_8159,N_5574,N_6093);
and U8160 (N_8160,N_5519,N_7288);
and U8161 (N_8161,N_7349,N_6769);
nand U8162 (N_8162,N_5052,N_5146);
nor U8163 (N_8163,N_5676,N_6689);
nand U8164 (N_8164,N_5506,N_7333);
nor U8165 (N_8165,N_6137,N_7179);
nand U8166 (N_8166,N_6343,N_5794);
and U8167 (N_8167,N_5520,N_5868);
nand U8168 (N_8168,N_5567,N_7124);
nand U8169 (N_8169,N_6344,N_5050);
and U8170 (N_8170,N_5833,N_5218);
nor U8171 (N_8171,N_5378,N_5545);
nor U8172 (N_8172,N_6882,N_5644);
nor U8173 (N_8173,N_5654,N_5920);
nand U8174 (N_8174,N_7051,N_7091);
nor U8175 (N_8175,N_5766,N_5302);
and U8176 (N_8176,N_5211,N_6071);
or U8177 (N_8177,N_6816,N_7328);
and U8178 (N_8178,N_7186,N_6361);
nor U8179 (N_8179,N_6402,N_6352);
nor U8180 (N_8180,N_6565,N_7006);
nand U8181 (N_8181,N_6651,N_7315);
and U8182 (N_8182,N_7414,N_7120);
nand U8183 (N_8183,N_6728,N_7099);
and U8184 (N_8184,N_6247,N_5565);
nand U8185 (N_8185,N_6460,N_6753);
xnor U8186 (N_8186,N_6324,N_6686);
xnor U8187 (N_8187,N_7446,N_7427);
and U8188 (N_8188,N_7486,N_5350);
or U8189 (N_8189,N_5055,N_7240);
or U8190 (N_8190,N_5973,N_5099);
and U8191 (N_8191,N_6230,N_7116);
nand U8192 (N_8192,N_5493,N_6783);
and U8193 (N_8193,N_6518,N_7148);
nand U8194 (N_8194,N_6577,N_6793);
nor U8195 (N_8195,N_5960,N_5255);
nand U8196 (N_8196,N_6589,N_5034);
nand U8197 (N_8197,N_6265,N_5885);
nor U8198 (N_8198,N_6421,N_5678);
nor U8199 (N_8199,N_6952,N_6010);
and U8200 (N_8200,N_6671,N_7261);
or U8201 (N_8201,N_5570,N_5571);
nand U8202 (N_8202,N_5916,N_5549);
and U8203 (N_8203,N_5236,N_5425);
or U8204 (N_8204,N_7471,N_6288);
and U8205 (N_8205,N_5521,N_6439);
nor U8206 (N_8206,N_7450,N_5844);
nand U8207 (N_8207,N_6433,N_5012);
nor U8208 (N_8208,N_5383,N_6307);
and U8209 (N_8209,N_6245,N_5418);
and U8210 (N_8210,N_5860,N_7456);
and U8211 (N_8211,N_6127,N_7039);
nand U8212 (N_8212,N_7420,N_7425);
nand U8213 (N_8213,N_5186,N_6511);
or U8214 (N_8214,N_5904,N_6373);
or U8215 (N_8215,N_5959,N_6993);
nor U8216 (N_8216,N_7377,N_5359);
and U8217 (N_8217,N_5858,N_5138);
and U8218 (N_8218,N_7117,N_5016);
nand U8219 (N_8219,N_5077,N_5301);
nor U8220 (N_8220,N_5339,N_6159);
and U8221 (N_8221,N_5724,N_5371);
nand U8222 (N_8222,N_6455,N_5516);
and U8223 (N_8223,N_7360,N_7424);
nand U8224 (N_8224,N_5419,N_7103);
nand U8225 (N_8225,N_5663,N_7076);
or U8226 (N_8226,N_5122,N_5801);
or U8227 (N_8227,N_7449,N_5630);
or U8228 (N_8228,N_6557,N_7281);
nor U8229 (N_8229,N_5223,N_6696);
nand U8230 (N_8230,N_6896,N_5276);
nor U8231 (N_8231,N_6961,N_6145);
nand U8232 (N_8232,N_6731,N_6536);
and U8233 (N_8233,N_6579,N_7164);
nor U8234 (N_8234,N_7239,N_6975);
or U8235 (N_8235,N_6524,N_6413);
nor U8236 (N_8236,N_5974,N_7469);
nand U8237 (N_8237,N_6188,N_7093);
and U8238 (N_8238,N_7200,N_6187);
nand U8239 (N_8239,N_6162,N_5754);
nand U8240 (N_8240,N_5370,N_5454);
nand U8241 (N_8241,N_5646,N_5288);
or U8242 (N_8242,N_5723,N_7085);
nor U8243 (N_8243,N_5251,N_6305);
nor U8244 (N_8244,N_7246,N_5994);
or U8245 (N_8245,N_5105,N_6999);
xor U8246 (N_8246,N_7289,N_7218);
nand U8247 (N_8247,N_6098,N_7397);
nor U8248 (N_8248,N_6065,N_5765);
nor U8249 (N_8249,N_6436,N_5870);
and U8250 (N_8250,N_6036,N_5949);
or U8251 (N_8251,N_6700,N_5606);
nand U8252 (N_8252,N_5772,N_5910);
and U8253 (N_8253,N_5197,N_5213);
nand U8254 (N_8254,N_6194,N_7369);
nand U8255 (N_8255,N_6982,N_5932);
or U8256 (N_8256,N_5648,N_5659);
and U8257 (N_8257,N_5640,N_5831);
or U8258 (N_8258,N_5316,N_6001);
nor U8259 (N_8259,N_6936,N_5231);
nand U8260 (N_8260,N_5581,N_6250);
and U8261 (N_8261,N_6841,N_6834);
and U8262 (N_8262,N_7033,N_6459);
nor U8263 (N_8263,N_5532,N_7435);
nor U8264 (N_8264,N_5591,N_5694);
nand U8265 (N_8265,N_7159,N_5124);
or U8266 (N_8266,N_7069,N_6947);
nand U8267 (N_8267,N_5911,N_5026);
nand U8268 (N_8268,N_5531,N_5563);
or U8269 (N_8269,N_5389,N_7358);
xnor U8270 (N_8270,N_5080,N_6809);
nor U8271 (N_8271,N_6858,N_6017);
nand U8272 (N_8272,N_5837,N_6398);
and U8273 (N_8273,N_6108,N_6939);
nor U8274 (N_8274,N_7479,N_7340);
or U8275 (N_8275,N_7109,N_6627);
and U8276 (N_8276,N_6949,N_6578);
or U8277 (N_8277,N_5121,N_7174);
or U8278 (N_8278,N_5488,N_5206);
nor U8279 (N_8279,N_6153,N_5082);
nor U8280 (N_8280,N_5040,N_6279);
nor U8281 (N_8281,N_5120,N_7004);
and U8282 (N_8282,N_7067,N_5342);
nor U8283 (N_8283,N_6233,N_6068);
nand U8284 (N_8284,N_6240,N_7331);
nor U8285 (N_8285,N_5072,N_6935);
or U8286 (N_8286,N_5578,N_6046);
nand U8287 (N_8287,N_5268,N_6171);
and U8288 (N_8288,N_7257,N_7440);
nor U8289 (N_8289,N_5372,N_6775);
nor U8290 (N_8290,N_5992,N_7081);
nor U8291 (N_8291,N_6467,N_7160);
nand U8292 (N_8292,N_6184,N_5972);
nor U8293 (N_8293,N_6105,N_5234);
nor U8294 (N_8294,N_6797,N_5698);
nand U8295 (N_8295,N_6110,N_6727);
nand U8296 (N_8296,N_6435,N_5669);
nor U8297 (N_8297,N_5020,N_6199);
nand U8298 (N_8298,N_7279,N_6259);
nand U8299 (N_8299,N_6507,N_7247);
nand U8300 (N_8300,N_6596,N_6119);
and U8301 (N_8301,N_6202,N_7070);
or U8302 (N_8302,N_5161,N_7321);
and U8303 (N_8303,N_5918,N_6531);
nand U8304 (N_8304,N_6296,N_6672);
nor U8305 (N_8305,N_6430,N_5224);
and U8306 (N_8306,N_5426,N_5909);
or U8307 (N_8307,N_7030,N_6837);
nor U8308 (N_8308,N_5847,N_6278);
nand U8309 (N_8309,N_7275,N_5954);
and U8310 (N_8310,N_6488,N_7278);
nor U8311 (N_8311,N_5641,N_6633);
and U8312 (N_8312,N_6217,N_7233);
and U8313 (N_8313,N_5229,N_5613);
nand U8314 (N_8314,N_5382,N_5458);
nand U8315 (N_8315,N_7249,N_7255);
nor U8316 (N_8316,N_6081,N_7016);
nand U8317 (N_8317,N_5891,N_6854);
and U8318 (N_8318,N_6072,N_5110);
or U8319 (N_8319,N_7142,N_5216);
or U8320 (N_8320,N_5414,N_5100);
nand U8321 (N_8321,N_5390,N_5612);
nand U8322 (N_8322,N_6221,N_6169);
or U8323 (N_8323,N_5356,N_6708);
nor U8324 (N_8324,N_7119,N_5380);
nand U8325 (N_8325,N_5608,N_7263);
nor U8326 (N_8326,N_5033,N_5619);
or U8327 (N_8327,N_6486,N_7243);
nor U8328 (N_8328,N_6276,N_5993);
and U8329 (N_8329,N_6251,N_5555);
and U8330 (N_8330,N_6568,N_5176);
nor U8331 (N_8331,N_5605,N_5963);
or U8332 (N_8332,N_5874,N_7287);
or U8333 (N_8333,N_5759,N_6100);
and U8334 (N_8334,N_5304,N_5123);
or U8335 (N_8335,N_7110,N_5622);
nor U8336 (N_8336,N_5310,N_6191);
and U8337 (N_8337,N_7231,N_6654);
xor U8338 (N_8338,N_5636,N_5851);
nand U8339 (N_8339,N_6808,N_5170);
nor U8340 (N_8340,N_6699,N_7419);
or U8341 (N_8341,N_6039,N_5348);
and U8342 (N_8342,N_6059,N_6729);
or U8343 (N_8343,N_6962,N_7282);
nand U8344 (N_8344,N_5321,N_5777);
or U8345 (N_8345,N_5582,N_5043);
nor U8346 (N_8346,N_7011,N_7300);
or U8347 (N_8347,N_5530,N_5906);
and U8348 (N_8348,N_6252,N_5944);
or U8349 (N_8349,N_6215,N_5756);
or U8350 (N_8350,N_5543,N_7245);
xor U8351 (N_8351,N_5843,N_6915);
nor U8352 (N_8352,N_7320,N_5938);
or U8353 (N_8353,N_7254,N_6216);
and U8354 (N_8354,N_5163,N_6909);
or U8355 (N_8355,N_5550,N_5129);
and U8356 (N_8356,N_6367,N_6794);
nor U8357 (N_8357,N_6979,N_6855);
nand U8358 (N_8358,N_5784,N_5778);
nand U8359 (N_8359,N_5553,N_7207);
nand U8360 (N_8360,N_6628,N_6530);
nor U8361 (N_8361,N_7253,N_5841);
nor U8362 (N_8362,N_6450,N_6066);
nand U8363 (N_8363,N_6472,N_6955);
nand U8364 (N_8364,N_5540,N_6434);
nand U8365 (N_8365,N_6287,N_6087);
nor U8366 (N_8366,N_6765,N_6884);
or U8367 (N_8367,N_7463,N_5670);
nor U8368 (N_8368,N_6035,N_6283);
and U8369 (N_8369,N_6750,N_5789);
and U8370 (N_8370,N_7177,N_5524);
or U8371 (N_8371,N_5492,N_5713);
and U8372 (N_8372,N_6730,N_7359);
or U8373 (N_8373,N_5047,N_7143);
nor U8374 (N_8374,N_6456,N_6692);
nand U8375 (N_8375,N_5159,N_6397);
and U8376 (N_8376,N_5869,N_6033);
nand U8377 (N_8377,N_6512,N_6029);
nor U8378 (N_8378,N_6338,N_5667);
nor U8379 (N_8379,N_6724,N_6998);
nor U8380 (N_8380,N_5770,N_5739);
and U8381 (N_8381,N_5456,N_5665);
nand U8382 (N_8382,N_6141,N_6097);
and U8383 (N_8383,N_6498,N_5162);
and U8384 (N_8384,N_6523,N_7228);
or U8385 (N_8385,N_7415,N_6848);
or U8386 (N_8386,N_6873,N_7370);
nor U8387 (N_8387,N_5501,N_6691);
nor U8388 (N_8388,N_5297,N_6304);
nor U8389 (N_8389,N_6302,N_7029);
nand U8390 (N_8390,N_7063,N_6281);
nor U8391 (N_8391,N_6368,N_6932);
nor U8392 (N_8392,N_6222,N_6869);
nor U8393 (N_8393,N_6832,N_7400);
xor U8394 (N_8394,N_5450,N_6800);
or U8395 (N_8395,N_7383,N_5092);
or U8396 (N_8396,N_5423,N_5286);
or U8397 (N_8397,N_5445,N_5190);
nor U8398 (N_8398,N_5629,N_5647);
or U8399 (N_8399,N_5679,N_5208);
and U8400 (N_8400,N_6570,N_5979);
and U8401 (N_8401,N_6702,N_6405);
or U8402 (N_8402,N_7133,N_5557);
nand U8403 (N_8403,N_7264,N_6242);
and U8404 (N_8404,N_6789,N_5088);
and U8405 (N_8405,N_5725,N_6569);
nor U8406 (N_8406,N_6051,N_6603);
and U8407 (N_8407,N_5795,N_5132);
and U8408 (N_8408,N_6757,N_5305);
and U8409 (N_8409,N_6192,N_6709);
and U8410 (N_8410,N_7170,N_7212);
nor U8411 (N_8411,N_5215,N_5925);
nand U8412 (N_8412,N_6553,N_6703);
nor U8413 (N_8413,N_5586,N_6420);
or U8414 (N_8414,N_5688,N_5751);
nand U8415 (N_8415,N_5025,N_5427);
nor U8416 (N_8416,N_5600,N_5965);
or U8417 (N_8417,N_5913,N_6289);
nor U8418 (N_8418,N_7176,N_6878);
nor U8419 (N_8419,N_6124,N_6657);
and U8420 (N_8420,N_6788,N_6556);
nand U8421 (N_8421,N_6683,N_6648);
nor U8422 (N_8422,N_6629,N_5746);
and U8423 (N_8423,N_5479,N_6911);
or U8424 (N_8424,N_5354,N_7454);
or U8425 (N_8425,N_7402,N_7439);
xnor U8426 (N_8426,N_6733,N_6534);
nand U8427 (N_8427,N_7074,N_5346);
nor U8428 (N_8428,N_5677,N_7474);
or U8429 (N_8429,N_5487,N_7322);
nand U8430 (N_8430,N_6111,N_6219);
and U8431 (N_8431,N_7350,N_7083);
nor U8432 (N_8432,N_6341,N_7058);
and U8433 (N_8433,N_5009,N_5845);
or U8434 (N_8434,N_7235,N_5707);
nor U8435 (N_8435,N_6091,N_5804);
or U8436 (N_8436,N_6958,N_5534);
or U8437 (N_8437,N_6677,N_5154);
and U8438 (N_8438,N_7344,N_6804);
nand U8439 (N_8439,N_6535,N_6544);
and U8440 (N_8440,N_5437,N_6901);
nand U8441 (N_8441,N_7422,N_5786);
nor U8442 (N_8442,N_6889,N_6198);
nand U8443 (N_8443,N_6086,N_5505);
nor U8444 (N_8444,N_6561,N_7111);
xnor U8445 (N_8445,N_6916,N_6235);
and U8446 (N_8446,N_5369,N_6712);
and U8447 (N_8447,N_5471,N_6168);
nand U8448 (N_8448,N_7185,N_6521);
nand U8449 (N_8449,N_6560,N_7153);
and U8450 (N_8450,N_6924,N_5160);
nand U8451 (N_8451,N_5222,N_6641);
nand U8452 (N_8452,N_5593,N_6382);
nand U8453 (N_8453,N_6316,N_5156);
nor U8454 (N_8454,N_5964,N_7303);
nand U8455 (N_8455,N_5289,N_5826);
and U8456 (N_8456,N_7466,N_6716);
and U8457 (N_8457,N_5542,N_5666);
nor U8458 (N_8458,N_7100,N_6419);
or U8459 (N_8459,N_5720,N_6481);
and U8460 (N_8460,N_5024,N_5075);
or U8461 (N_8461,N_6391,N_5421);
nor U8462 (N_8462,N_6552,N_5355);
and U8463 (N_8463,N_5062,N_7393);
nand U8464 (N_8464,N_5349,N_7214);
and U8465 (N_8465,N_5796,N_5307);
nor U8466 (N_8466,N_7337,N_5701);
and U8467 (N_8467,N_5384,N_6748);
nor U8468 (N_8468,N_7138,N_6404);
nor U8469 (N_8469,N_5402,N_5265);
and U8470 (N_8470,N_5252,N_5599);
or U8471 (N_8471,N_6122,N_6723);
or U8472 (N_8472,N_5812,N_6272);
or U8473 (N_8473,N_6147,N_5849);
nor U8474 (N_8474,N_5687,N_7208);
or U8475 (N_8475,N_6246,N_6015);
nor U8476 (N_8476,N_6270,N_7252);
nor U8477 (N_8477,N_6381,N_5857);
and U8478 (N_8478,N_7230,N_5165);
nand U8479 (N_8479,N_5624,N_6190);
nor U8480 (N_8480,N_7190,N_6005);
and U8481 (N_8481,N_6423,N_5148);
nand U8482 (N_8482,N_6921,N_7444);
or U8483 (N_8483,N_5935,N_5643);
or U8484 (N_8484,N_7267,N_6494);
and U8485 (N_8485,N_6244,N_7436);
and U8486 (N_8486,N_6581,N_5089);
and U8487 (N_8487,N_6610,N_7368);
and U8488 (N_8488,N_7071,N_5250);
and U8489 (N_8489,N_5424,N_7334);
and U8490 (N_8490,N_5997,N_6377);
nand U8491 (N_8491,N_6390,N_6129);
nor U8492 (N_8492,N_6555,N_5975);
and U8493 (N_8493,N_6303,N_5865);
or U8494 (N_8494,N_5285,N_5246);
nand U8495 (N_8495,N_5434,N_5056);
nor U8496 (N_8496,N_5558,N_6009);
and U8497 (N_8497,N_5829,N_5988);
and U8498 (N_8498,N_6079,N_5477);
nor U8499 (N_8499,N_5939,N_6666);
nor U8500 (N_8500,N_7134,N_7272);
nand U8501 (N_8501,N_6675,N_5816);
nand U8502 (N_8502,N_6743,N_6432);
and U8503 (N_8503,N_5191,N_7290);
or U8504 (N_8504,N_5706,N_7242);
nand U8505 (N_8505,N_5690,N_7079);
and U8506 (N_8506,N_6380,N_7362);
and U8507 (N_8507,N_6795,N_5198);
nor U8508 (N_8508,N_7494,N_6030);
or U8509 (N_8509,N_7324,N_6102);
or U8510 (N_8510,N_6150,N_6101);
or U8511 (N_8511,N_6151,N_5693);
or U8512 (N_8512,N_6802,N_6929);
or U8513 (N_8513,N_5060,N_6746);
and U8514 (N_8514,N_6177,N_7367);
xnor U8515 (N_8515,N_6000,N_5769);
or U8516 (N_8516,N_5274,N_5757);
nor U8517 (N_8517,N_6018,N_7147);
nand U8518 (N_8518,N_6013,N_5898);
nand U8519 (N_8519,N_7348,N_5194);
nor U8520 (N_8520,N_6923,N_5320);
nand U8521 (N_8521,N_7330,N_5011);
or U8522 (N_8522,N_7156,N_7381);
xor U8523 (N_8523,N_5924,N_6917);
nor U8524 (N_8524,N_6075,N_6266);
nor U8525 (N_8525,N_6464,N_5884);
nand U8526 (N_8526,N_5125,N_7408);
and U8527 (N_8527,N_5956,N_6031);
nand U8528 (N_8528,N_7418,N_7129);
and U8529 (N_8529,N_5027,N_7163);
or U8530 (N_8530,N_7131,N_6851);
and U8531 (N_8531,N_7490,N_6604);
or U8532 (N_8532,N_7356,N_5399);
nand U8533 (N_8533,N_5902,N_5495);
and U8534 (N_8534,N_6698,N_7318);
and U8535 (N_8535,N_7041,N_5788);
nand U8536 (N_8536,N_5594,N_6203);
and U8537 (N_8537,N_7489,N_6364);
and U8538 (N_8538,N_7488,N_6027);
nand U8539 (N_8539,N_6706,N_6532);
and U8540 (N_8540,N_6256,N_5561);
or U8541 (N_8541,N_5496,N_5998);
nor U8542 (N_8542,N_5014,N_6468);
nor U8543 (N_8543,N_5281,N_6886);
nand U8544 (N_8544,N_5200,N_5326);
and U8545 (N_8545,N_6427,N_5241);
nand U8546 (N_8546,N_5855,N_5970);
and U8547 (N_8547,N_6621,N_5957);
and U8548 (N_8548,N_6264,N_5463);
and U8549 (N_8549,N_5554,N_5167);
or U8550 (N_8550,N_5940,N_7101);
and U8551 (N_8551,N_6311,N_6331);
and U8552 (N_8552,N_6337,N_7045);
nor U8553 (N_8553,N_5412,N_7459);
or U8554 (N_8554,N_6611,N_7175);
nor U8555 (N_8555,N_6940,N_5443);
nand U8556 (N_8556,N_5566,N_7007);
and U8557 (N_8557,N_7061,N_6957);
nand U8558 (N_8558,N_7105,N_6576);
and U8559 (N_8559,N_5319,N_5958);
or U8560 (N_8560,N_6325,N_5598);
nor U8561 (N_8561,N_6751,N_5942);
nand U8562 (N_8562,N_6115,N_6070);
or U8563 (N_8563,N_6639,N_6056);
nand U8564 (N_8564,N_7354,N_6318);
nor U8565 (N_8565,N_5967,N_6038);
or U8566 (N_8566,N_7309,N_6292);
nand U8567 (N_8567,N_6062,N_6340);
or U8568 (N_8568,N_6366,N_5270);
or U8569 (N_8569,N_6670,N_5758);
nor U8570 (N_8570,N_6294,N_6146);
nor U8571 (N_8571,N_7022,N_5546);
nand U8572 (N_8572,N_6768,N_6394);
and U8573 (N_8573,N_5509,N_5106);
nor U8574 (N_8574,N_6234,N_5905);
xor U8575 (N_8575,N_6564,N_6261);
or U8576 (N_8576,N_7270,N_7000);
nand U8577 (N_8577,N_5396,N_7122);
nor U8578 (N_8578,N_6668,N_7299);
nor U8579 (N_8579,N_7308,N_6104);
nor U8580 (N_8580,N_5373,N_6566);
nor U8581 (N_8581,N_6126,N_6548);
and U8582 (N_8582,N_6440,N_5569);
nand U8583 (N_8583,N_7412,N_6539);
nand U8584 (N_8584,N_5249,N_7258);
and U8585 (N_8585,N_6461,N_5248);
or U8586 (N_8586,N_5361,N_6824);
nand U8587 (N_8587,N_7115,N_6836);
or U8588 (N_8588,N_7392,N_5649);
and U8589 (N_8589,N_6857,N_7135);
and U8590 (N_8590,N_6685,N_5481);
or U8591 (N_8591,N_6694,N_6914);
and U8592 (N_8592,N_5484,N_7399);
nor U8593 (N_8593,N_5151,N_5332);
nand U8594 (N_8594,N_5245,N_6843);
and U8595 (N_8595,N_5282,N_5783);
or U8596 (N_8596,N_6181,N_5514);
nor U8597 (N_8597,N_5962,N_5889);
and U8598 (N_8598,N_6722,N_5196);
or U8599 (N_8599,N_6609,N_5755);
or U8600 (N_8600,N_6739,N_6525);
nand U8601 (N_8601,N_5470,N_6422);
nand U8602 (N_8602,N_6179,N_6659);
and U8603 (N_8603,N_6371,N_5284);
and U8604 (N_8604,N_6197,N_7311);
or U8605 (N_8605,N_6232,N_5335);
nor U8606 (N_8606,N_6635,N_5515);
or U8607 (N_8607,N_6474,N_5366);
nand U8608 (N_8608,N_5827,N_6875);
or U8609 (N_8609,N_6582,N_6262);
or U8610 (N_8610,N_7193,N_6083);
nand U8611 (N_8611,N_7087,N_5404);
or U8612 (N_8612,N_6362,N_6506);
or U8613 (N_8613,N_5300,N_6607);
nor U8614 (N_8614,N_7210,N_5192);
and U8615 (N_8615,N_6658,N_5824);
and U8616 (N_8616,N_6089,N_5432);
or U8617 (N_8617,N_6705,N_5947);
or U8618 (N_8618,N_6032,N_5631);
nor U8619 (N_8619,N_6701,N_6740);
nor U8620 (N_8620,N_5433,N_7166);
and U8621 (N_8621,N_5996,N_6810);
and U8622 (N_8622,N_6273,N_5188);
and U8623 (N_8623,N_5653,N_7053);
nor U8624 (N_8624,N_5296,N_7429);
xor U8625 (N_8625,N_5358,N_5971);
and U8626 (N_8626,N_5312,N_6959);
nand U8627 (N_8627,N_5256,N_5351);
nand U8628 (N_8628,N_6925,N_6085);
nand U8629 (N_8629,N_7434,N_6342);
or U8630 (N_8630,N_6981,N_7409);
and U8631 (N_8631,N_6950,N_7059);
nor U8632 (N_8632,N_7080,N_6774);
nand U8633 (N_8633,N_6517,N_6131);
nor U8634 (N_8634,N_5526,N_5375);
nor U8635 (N_8635,N_6850,N_5742);
nand U8636 (N_8636,N_6502,N_6735);
and U8637 (N_8637,N_7056,N_5547);
and U8638 (N_8638,N_6897,N_5244);
nand U8639 (N_8639,N_5243,N_5533);
nand U8640 (N_8640,N_5656,N_5347);
nand U8641 (N_8641,N_5856,N_6644);
nand U8642 (N_8642,N_7003,N_7095);
or U8643 (N_8643,N_5923,N_6313);
or U8644 (N_8644,N_6779,N_6931);
or U8645 (N_8645,N_6613,N_6465);
nor U8646 (N_8646,N_6574,N_6856);
or U8647 (N_8647,N_5875,N_5899);
and U8648 (N_8648,N_5886,N_6585);
nor U8649 (N_8649,N_6767,N_6825);
or U8650 (N_8650,N_7384,N_5753);
nor U8651 (N_8651,N_6462,N_5933);
nor U8652 (N_8652,N_5280,N_7379);
xor U8653 (N_8653,N_5172,N_6586);
and U8654 (N_8654,N_5005,N_5601);
and U8655 (N_8655,N_5113,N_6587);
nand U8656 (N_8656,N_5360,N_7078);
nor U8657 (N_8657,N_6480,N_5135);
or U8658 (N_8658,N_6991,N_7283);
nor U8659 (N_8659,N_6374,N_6227);
nand U8660 (N_8660,N_5287,N_7165);
or U8661 (N_8661,N_6084,N_5177);
nor U8662 (N_8662,N_7336,N_5417);
or U8663 (N_8663,N_6008,N_6183);
nand U8664 (N_8664,N_5596,N_6833);
and U8665 (N_8665,N_5685,N_6772);
nand U8666 (N_8666,N_5580,N_5607);
and U8667 (N_8667,N_6471,N_5609);
nand U8668 (N_8668,N_6058,N_5981);
and U8669 (N_8669,N_6428,N_5948);
nand U8670 (N_8670,N_5802,N_5067);
nor U8671 (N_8671,N_7149,N_7472);
and U8672 (N_8672,N_5239,N_7411);
nor U8673 (N_8673,N_6688,N_5908);
nor U8674 (N_8674,N_6176,N_6166);
xnor U8675 (N_8675,N_6446,N_5469);
or U8676 (N_8676,N_6055,N_7430);
or U8677 (N_8677,N_5931,N_5061);
nor U8678 (N_8678,N_6543,N_7161);
and U8679 (N_8679,N_7498,N_6645);
nand U8680 (N_8680,N_6780,N_6175);
and U8681 (N_8681,N_5790,N_7188);
and U8682 (N_8682,N_6409,N_5696);
and U8683 (N_8683,N_5749,N_6257);
or U8684 (N_8684,N_5711,N_7447);
and U8685 (N_8685,N_5271,N_5438);
and U8686 (N_8686,N_5651,N_5782);
nand U8687 (N_8687,N_5087,N_6116);
and U8688 (N_8688,N_5986,N_5951);
nor U8689 (N_8689,N_6653,N_6870);
or U8690 (N_8690,N_5136,N_7317);
nand U8691 (N_8691,N_5684,N_5576);
nor U8692 (N_8692,N_6693,N_5333);
or U8693 (N_8693,N_6475,N_5779);
nand U8694 (N_8694,N_6831,N_7416);
nor U8695 (N_8695,N_6479,N_6128);
and U8696 (N_8696,N_5409,N_6660);
or U8697 (N_8697,N_6852,N_5626);
nand U8698 (N_8698,N_7347,N_7236);
nor U8699 (N_8699,N_6054,N_6844);
nand U8700 (N_8700,N_5675,N_6415);
and U8701 (N_8701,N_5500,N_6414);
and U8702 (N_8702,N_6736,N_5941);
or U8703 (N_8703,N_6339,N_6328);
or U8704 (N_8704,N_6061,N_7121);
nor U8705 (N_8705,N_5822,N_7150);
or U8706 (N_8706,N_5397,N_7189);
nor U8707 (N_8707,N_5093,N_5903);
or U8708 (N_8708,N_6538,N_5130);
nand U8709 (N_8709,N_6995,N_5806);
or U8710 (N_8710,N_5853,N_6782);
nor U8711 (N_8711,N_5568,N_7173);
nor U8712 (N_8712,N_6983,N_5538);
nand U8713 (N_8713,N_5736,N_5633);
nand U8714 (N_8714,N_5334,N_6829);
and U8715 (N_8715,N_5155,N_5173);
nand U8716 (N_8716,N_6329,N_5589);
nand U8717 (N_8717,N_6966,N_7038);
nor U8718 (N_8718,N_6673,N_5590);
or U8719 (N_8719,N_5621,N_6354);
or U8720 (N_8720,N_6811,N_5657);
nand U8721 (N_8721,N_5415,N_6417);
nor U8722 (N_8722,N_6817,N_5053);
and U8723 (N_8723,N_5203,N_5314);
or U8724 (N_8724,N_6927,N_5401);
or U8725 (N_8725,N_7277,N_5046);
nor U8726 (N_8726,N_5512,N_5466);
nor U8727 (N_8727,N_6157,N_5071);
and U8728 (N_8728,N_6926,N_6453);
and U8729 (N_8729,N_7075,N_6358);
or U8730 (N_8730,N_6652,N_6149);
nor U8731 (N_8731,N_6720,N_6719);
nand U8732 (N_8732,N_6385,N_6021);
nand U8733 (N_8733,N_7426,N_7407);
nor U8734 (N_8734,N_5485,N_5719);
xnor U8735 (N_8735,N_6559,N_6226);
and U8736 (N_8736,N_6269,N_5079);
or U8737 (N_8737,N_5405,N_6988);
nor U8738 (N_8738,N_6928,N_5023);
and U8739 (N_8739,N_7465,N_6575);
or U8740 (N_8740,N_5836,N_5465);
and U8741 (N_8741,N_7229,N_7364);
or U8742 (N_8742,N_6590,N_6562);
nor U8743 (N_8743,N_6387,N_5714);
nand U8744 (N_8744,N_7215,N_6863);
nor U8745 (N_8745,N_7326,N_5367);
or U8746 (N_8746,N_6593,N_7438);
or U8747 (N_8747,N_6006,N_7374);
or U8748 (N_8748,N_7388,N_5452);
or U8749 (N_8749,N_5848,N_7468);
or U8750 (N_8750,N_5333,N_5215);
or U8751 (N_8751,N_5715,N_6441);
nand U8752 (N_8752,N_6714,N_6349);
nor U8753 (N_8753,N_5120,N_6783);
or U8754 (N_8754,N_6283,N_5215);
nand U8755 (N_8755,N_5263,N_7340);
nor U8756 (N_8756,N_5793,N_6095);
nand U8757 (N_8757,N_6999,N_5279);
nor U8758 (N_8758,N_5869,N_6446);
and U8759 (N_8759,N_5782,N_7303);
and U8760 (N_8760,N_6027,N_6496);
and U8761 (N_8761,N_5734,N_6139);
or U8762 (N_8762,N_7448,N_5520);
nand U8763 (N_8763,N_5828,N_6224);
xnor U8764 (N_8764,N_5144,N_6366);
or U8765 (N_8765,N_6190,N_6734);
and U8766 (N_8766,N_5060,N_6668);
or U8767 (N_8767,N_5493,N_7293);
and U8768 (N_8768,N_6521,N_5303);
nor U8769 (N_8769,N_6804,N_6120);
nor U8770 (N_8770,N_7483,N_5236);
nand U8771 (N_8771,N_6365,N_6118);
nor U8772 (N_8772,N_6938,N_6319);
and U8773 (N_8773,N_6007,N_6180);
and U8774 (N_8774,N_5539,N_7282);
or U8775 (N_8775,N_5901,N_6716);
or U8776 (N_8776,N_5834,N_7039);
nand U8777 (N_8777,N_6151,N_6047);
and U8778 (N_8778,N_5953,N_6268);
nand U8779 (N_8779,N_5546,N_5004);
and U8780 (N_8780,N_5995,N_5596);
nand U8781 (N_8781,N_6539,N_5818);
or U8782 (N_8782,N_7121,N_5974);
or U8783 (N_8783,N_5616,N_6473);
nand U8784 (N_8784,N_6583,N_6005);
nor U8785 (N_8785,N_5655,N_5916);
and U8786 (N_8786,N_5897,N_7496);
or U8787 (N_8787,N_7291,N_7378);
nor U8788 (N_8788,N_6058,N_6138);
and U8789 (N_8789,N_5075,N_5132);
xnor U8790 (N_8790,N_7040,N_5077);
nand U8791 (N_8791,N_6171,N_5334);
nand U8792 (N_8792,N_6443,N_6758);
nor U8793 (N_8793,N_5399,N_6276);
and U8794 (N_8794,N_5293,N_5552);
or U8795 (N_8795,N_6248,N_5702);
and U8796 (N_8796,N_6117,N_6944);
and U8797 (N_8797,N_6466,N_6624);
and U8798 (N_8798,N_5333,N_5055);
or U8799 (N_8799,N_5941,N_5687);
and U8800 (N_8800,N_5176,N_6560);
or U8801 (N_8801,N_6608,N_6905);
nor U8802 (N_8802,N_6034,N_5664);
nand U8803 (N_8803,N_5524,N_6256);
or U8804 (N_8804,N_5610,N_6850);
nand U8805 (N_8805,N_5886,N_5386);
nor U8806 (N_8806,N_6296,N_5353);
nand U8807 (N_8807,N_6933,N_6294);
and U8808 (N_8808,N_6555,N_6321);
nand U8809 (N_8809,N_7104,N_6589);
nand U8810 (N_8810,N_7006,N_6512);
and U8811 (N_8811,N_5691,N_6877);
or U8812 (N_8812,N_7452,N_6896);
nor U8813 (N_8813,N_6231,N_7079);
nand U8814 (N_8814,N_6633,N_6946);
or U8815 (N_8815,N_6253,N_6585);
or U8816 (N_8816,N_5433,N_6724);
nand U8817 (N_8817,N_5619,N_5741);
or U8818 (N_8818,N_6049,N_7208);
or U8819 (N_8819,N_5119,N_5835);
and U8820 (N_8820,N_5956,N_5613);
nand U8821 (N_8821,N_5906,N_5528);
or U8822 (N_8822,N_5000,N_6564);
or U8823 (N_8823,N_5500,N_5539);
nor U8824 (N_8824,N_6416,N_5020);
nor U8825 (N_8825,N_6308,N_5090);
nand U8826 (N_8826,N_6785,N_5851);
or U8827 (N_8827,N_5333,N_6353);
and U8828 (N_8828,N_5724,N_6986);
nor U8829 (N_8829,N_5289,N_5606);
nor U8830 (N_8830,N_6320,N_6928);
nand U8831 (N_8831,N_5801,N_7003);
and U8832 (N_8832,N_6606,N_5112);
nor U8833 (N_8833,N_6545,N_6104);
or U8834 (N_8834,N_5730,N_6082);
or U8835 (N_8835,N_6027,N_5640);
or U8836 (N_8836,N_5029,N_6660);
or U8837 (N_8837,N_6024,N_6601);
and U8838 (N_8838,N_5773,N_5962);
or U8839 (N_8839,N_6371,N_7137);
nor U8840 (N_8840,N_6223,N_7025);
nor U8841 (N_8841,N_6422,N_5380);
and U8842 (N_8842,N_5404,N_5218);
or U8843 (N_8843,N_7303,N_5839);
and U8844 (N_8844,N_7017,N_5101);
nand U8845 (N_8845,N_6157,N_6261);
or U8846 (N_8846,N_5475,N_5162);
and U8847 (N_8847,N_5504,N_5486);
nor U8848 (N_8848,N_6969,N_6074);
and U8849 (N_8849,N_7476,N_5744);
or U8850 (N_8850,N_5146,N_6333);
nand U8851 (N_8851,N_6382,N_6711);
and U8852 (N_8852,N_6073,N_5678);
and U8853 (N_8853,N_6515,N_6174);
nand U8854 (N_8854,N_6730,N_7092);
or U8855 (N_8855,N_5975,N_5229);
nand U8856 (N_8856,N_6259,N_5996);
and U8857 (N_8857,N_6703,N_6775);
nor U8858 (N_8858,N_5365,N_5813);
or U8859 (N_8859,N_6298,N_5719);
and U8860 (N_8860,N_7368,N_5058);
nand U8861 (N_8861,N_5918,N_6984);
or U8862 (N_8862,N_7054,N_5215);
nand U8863 (N_8863,N_6859,N_5865);
nor U8864 (N_8864,N_6803,N_5392);
nor U8865 (N_8865,N_6518,N_6284);
nand U8866 (N_8866,N_5258,N_6287);
nor U8867 (N_8867,N_5936,N_6800);
and U8868 (N_8868,N_7354,N_7020);
nand U8869 (N_8869,N_7240,N_6217);
nor U8870 (N_8870,N_7248,N_5401);
and U8871 (N_8871,N_6284,N_5089);
or U8872 (N_8872,N_6338,N_5427);
nor U8873 (N_8873,N_5800,N_6807);
or U8874 (N_8874,N_6116,N_6743);
and U8875 (N_8875,N_5625,N_5867);
and U8876 (N_8876,N_5386,N_6929);
or U8877 (N_8877,N_7024,N_5806);
nand U8878 (N_8878,N_6415,N_6289);
xnor U8879 (N_8879,N_6429,N_7327);
or U8880 (N_8880,N_5111,N_5397);
and U8881 (N_8881,N_5001,N_7059);
nand U8882 (N_8882,N_5812,N_5897);
or U8883 (N_8883,N_5523,N_5062);
and U8884 (N_8884,N_6354,N_5121);
and U8885 (N_8885,N_7464,N_6702);
and U8886 (N_8886,N_6123,N_6114);
or U8887 (N_8887,N_7135,N_5251);
or U8888 (N_8888,N_6482,N_6754);
nor U8889 (N_8889,N_5772,N_5076);
nor U8890 (N_8890,N_6469,N_6001);
and U8891 (N_8891,N_5717,N_6323);
nor U8892 (N_8892,N_6803,N_7294);
nor U8893 (N_8893,N_7300,N_5179);
nand U8894 (N_8894,N_5255,N_7033);
and U8895 (N_8895,N_7170,N_7469);
nor U8896 (N_8896,N_6035,N_6318);
or U8897 (N_8897,N_7152,N_6382);
and U8898 (N_8898,N_6425,N_5350);
or U8899 (N_8899,N_6268,N_7035);
and U8900 (N_8900,N_6080,N_6729);
or U8901 (N_8901,N_6724,N_5982);
or U8902 (N_8902,N_6426,N_7401);
xnor U8903 (N_8903,N_7021,N_6273);
nor U8904 (N_8904,N_6479,N_6607);
or U8905 (N_8905,N_7306,N_7235);
and U8906 (N_8906,N_6999,N_5995);
nor U8907 (N_8907,N_6700,N_5323);
xor U8908 (N_8908,N_6060,N_7368);
nand U8909 (N_8909,N_5408,N_7082);
or U8910 (N_8910,N_5555,N_6925);
and U8911 (N_8911,N_6308,N_5476);
nor U8912 (N_8912,N_6293,N_6458);
nand U8913 (N_8913,N_5769,N_7106);
and U8914 (N_8914,N_5790,N_6138);
or U8915 (N_8915,N_7152,N_5385);
or U8916 (N_8916,N_5563,N_6999);
or U8917 (N_8917,N_5332,N_6674);
nand U8918 (N_8918,N_7361,N_7128);
nor U8919 (N_8919,N_5786,N_6467);
nand U8920 (N_8920,N_5193,N_7462);
nand U8921 (N_8921,N_5968,N_5222);
and U8922 (N_8922,N_5271,N_6554);
and U8923 (N_8923,N_7030,N_5204);
or U8924 (N_8924,N_6170,N_5435);
and U8925 (N_8925,N_5985,N_7479);
or U8926 (N_8926,N_5854,N_5385);
nand U8927 (N_8927,N_6096,N_5676);
nor U8928 (N_8928,N_7459,N_5520);
nand U8929 (N_8929,N_6298,N_7229);
or U8930 (N_8930,N_5162,N_5579);
or U8931 (N_8931,N_6828,N_6290);
nor U8932 (N_8932,N_5175,N_5622);
and U8933 (N_8933,N_7142,N_7379);
or U8934 (N_8934,N_5325,N_5206);
and U8935 (N_8935,N_7255,N_6120);
and U8936 (N_8936,N_5183,N_7423);
or U8937 (N_8937,N_5306,N_6674);
or U8938 (N_8938,N_6470,N_6995);
nand U8939 (N_8939,N_5005,N_6653);
and U8940 (N_8940,N_5588,N_6583);
nand U8941 (N_8941,N_5387,N_6061);
nor U8942 (N_8942,N_6845,N_6995);
nor U8943 (N_8943,N_5553,N_6704);
or U8944 (N_8944,N_7029,N_7371);
or U8945 (N_8945,N_7298,N_5715);
or U8946 (N_8946,N_5538,N_6808);
or U8947 (N_8947,N_5139,N_6319);
nand U8948 (N_8948,N_6122,N_6682);
or U8949 (N_8949,N_5025,N_5053);
nand U8950 (N_8950,N_5380,N_5254);
and U8951 (N_8951,N_6743,N_6590);
nand U8952 (N_8952,N_5865,N_5948);
nand U8953 (N_8953,N_5803,N_6174);
nor U8954 (N_8954,N_7228,N_5482);
nor U8955 (N_8955,N_7105,N_6768);
nor U8956 (N_8956,N_7315,N_5138);
nor U8957 (N_8957,N_5004,N_7478);
nand U8958 (N_8958,N_7425,N_7166);
or U8959 (N_8959,N_6028,N_5078);
or U8960 (N_8960,N_6788,N_5076);
nand U8961 (N_8961,N_6992,N_6553);
and U8962 (N_8962,N_6849,N_5216);
nor U8963 (N_8963,N_7496,N_6373);
nor U8964 (N_8964,N_6834,N_5603);
or U8965 (N_8965,N_5874,N_6405);
or U8966 (N_8966,N_7345,N_6242);
and U8967 (N_8967,N_5545,N_6005);
and U8968 (N_8968,N_7140,N_6231);
nor U8969 (N_8969,N_5019,N_7495);
nand U8970 (N_8970,N_7422,N_5612);
nand U8971 (N_8971,N_6669,N_7093);
nand U8972 (N_8972,N_5474,N_6310);
nand U8973 (N_8973,N_6629,N_6455);
or U8974 (N_8974,N_5651,N_6076);
and U8975 (N_8975,N_5795,N_6273);
nand U8976 (N_8976,N_7392,N_7172);
or U8977 (N_8977,N_6138,N_6927);
or U8978 (N_8978,N_6528,N_6359);
and U8979 (N_8979,N_5357,N_5564);
nand U8980 (N_8980,N_5136,N_6657);
nor U8981 (N_8981,N_6520,N_6978);
nor U8982 (N_8982,N_5188,N_7154);
nor U8983 (N_8983,N_6240,N_6726);
and U8984 (N_8984,N_5211,N_6656);
nor U8985 (N_8985,N_5379,N_6696);
or U8986 (N_8986,N_5840,N_6668);
nor U8987 (N_8987,N_5084,N_6749);
nand U8988 (N_8988,N_5121,N_5838);
and U8989 (N_8989,N_5723,N_6116);
or U8990 (N_8990,N_5299,N_5626);
nor U8991 (N_8991,N_5520,N_6458);
nor U8992 (N_8992,N_6920,N_6428);
and U8993 (N_8993,N_7345,N_5221);
or U8994 (N_8994,N_5981,N_6345);
or U8995 (N_8995,N_5219,N_5445);
nor U8996 (N_8996,N_7013,N_5423);
nor U8997 (N_8997,N_6769,N_7496);
or U8998 (N_8998,N_7019,N_6873);
and U8999 (N_8999,N_7021,N_5327);
and U9000 (N_9000,N_7383,N_7044);
nor U9001 (N_9001,N_5945,N_5841);
or U9002 (N_9002,N_6404,N_6659);
nand U9003 (N_9003,N_5159,N_7324);
nand U9004 (N_9004,N_7419,N_6445);
nand U9005 (N_9005,N_6130,N_6492);
nand U9006 (N_9006,N_6731,N_5259);
and U9007 (N_9007,N_6688,N_6514);
xor U9008 (N_9008,N_5614,N_5873);
nor U9009 (N_9009,N_7290,N_6930);
nand U9010 (N_9010,N_6678,N_6460);
and U9011 (N_9011,N_5435,N_6567);
nor U9012 (N_9012,N_6956,N_7080);
and U9013 (N_9013,N_5498,N_7026);
nand U9014 (N_9014,N_6575,N_6684);
xor U9015 (N_9015,N_6163,N_5010);
or U9016 (N_9016,N_6498,N_6335);
nor U9017 (N_9017,N_5535,N_6690);
or U9018 (N_9018,N_6593,N_5830);
nor U9019 (N_9019,N_6620,N_7366);
nor U9020 (N_9020,N_7000,N_6757);
or U9021 (N_9021,N_6972,N_5067);
nor U9022 (N_9022,N_6852,N_5713);
nor U9023 (N_9023,N_6599,N_6206);
nor U9024 (N_9024,N_6095,N_6008);
and U9025 (N_9025,N_6204,N_6941);
or U9026 (N_9026,N_6197,N_5716);
or U9027 (N_9027,N_6505,N_7330);
nand U9028 (N_9028,N_6007,N_6682);
or U9029 (N_9029,N_7479,N_7379);
nor U9030 (N_9030,N_6439,N_6693);
xnor U9031 (N_9031,N_5334,N_7315);
or U9032 (N_9032,N_6516,N_6500);
nand U9033 (N_9033,N_6721,N_5934);
nor U9034 (N_9034,N_5196,N_5240);
nor U9035 (N_9035,N_6010,N_6446);
xor U9036 (N_9036,N_7357,N_5051);
or U9037 (N_9037,N_6880,N_6712);
nand U9038 (N_9038,N_5869,N_5901);
and U9039 (N_9039,N_6616,N_5833);
or U9040 (N_9040,N_6051,N_5838);
or U9041 (N_9041,N_5567,N_5035);
xor U9042 (N_9042,N_5710,N_7150);
nand U9043 (N_9043,N_7088,N_6367);
or U9044 (N_9044,N_6474,N_6998);
xnor U9045 (N_9045,N_5204,N_6450);
nand U9046 (N_9046,N_5969,N_6827);
or U9047 (N_9047,N_6304,N_5887);
nor U9048 (N_9048,N_5263,N_6600);
nand U9049 (N_9049,N_6676,N_5370);
nand U9050 (N_9050,N_5182,N_5349);
and U9051 (N_9051,N_7335,N_6489);
and U9052 (N_9052,N_6157,N_7338);
and U9053 (N_9053,N_6685,N_6881);
or U9054 (N_9054,N_5761,N_7443);
nor U9055 (N_9055,N_5522,N_6389);
nor U9056 (N_9056,N_7333,N_6477);
nand U9057 (N_9057,N_6710,N_5590);
or U9058 (N_9058,N_6237,N_5512);
or U9059 (N_9059,N_6443,N_5855);
nand U9060 (N_9060,N_6470,N_6245);
nand U9061 (N_9061,N_6903,N_5379);
or U9062 (N_9062,N_5106,N_6912);
nand U9063 (N_9063,N_5339,N_7397);
and U9064 (N_9064,N_7451,N_7463);
or U9065 (N_9065,N_5063,N_6296);
or U9066 (N_9066,N_6468,N_5745);
nand U9067 (N_9067,N_5211,N_6584);
nand U9068 (N_9068,N_5538,N_6444);
and U9069 (N_9069,N_5316,N_5644);
or U9070 (N_9070,N_6081,N_5052);
and U9071 (N_9071,N_6696,N_6292);
and U9072 (N_9072,N_6625,N_7067);
nand U9073 (N_9073,N_5303,N_6514);
nand U9074 (N_9074,N_6254,N_7420);
nor U9075 (N_9075,N_7376,N_5892);
or U9076 (N_9076,N_5996,N_6746);
nand U9077 (N_9077,N_6241,N_5457);
nor U9078 (N_9078,N_6158,N_6093);
and U9079 (N_9079,N_6570,N_6790);
xor U9080 (N_9080,N_6335,N_5808);
or U9081 (N_9081,N_5774,N_5260);
nand U9082 (N_9082,N_5728,N_5479);
and U9083 (N_9083,N_6554,N_5255);
and U9084 (N_9084,N_5834,N_7477);
nor U9085 (N_9085,N_7112,N_7487);
or U9086 (N_9086,N_7165,N_6094);
nand U9087 (N_9087,N_5203,N_6650);
or U9088 (N_9088,N_6028,N_7373);
and U9089 (N_9089,N_5943,N_6679);
nor U9090 (N_9090,N_6887,N_5852);
nand U9091 (N_9091,N_5213,N_6180);
nor U9092 (N_9092,N_5952,N_6133);
and U9093 (N_9093,N_6438,N_5022);
xnor U9094 (N_9094,N_5482,N_6746);
nor U9095 (N_9095,N_7097,N_7220);
or U9096 (N_9096,N_6791,N_5466);
nand U9097 (N_9097,N_7133,N_5171);
nand U9098 (N_9098,N_6028,N_5498);
and U9099 (N_9099,N_6490,N_6145);
and U9100 (N_9100,N_5118,N_5530);
and U9101 (N_9101,N_5224,N_5937);
nor U9102 (N_9102,N_6000,N_6690);
or U9103 (N_9103,N_6486,N_5078);
and U9104 (N_9104,N_6543,N_5744);
or U9105 (N_9105,N_6337,N_6563);
nor U9106 (N_9106,N_7402,N_7253);
nor U9107 (N_9107,N_5754,N_5936);
nand U9108 (N_9108,N_5366,N_5120);
nand U9109 (N_9109,N_6606,N_5105);
and U9110 (N_9110,N_6896,N_5161);
and U9111 (N_9111,N_5115,N_6669);
nor U9112 (N_9112,N_6958,N_5040);
and U9113 (N_9113,N_5639,N_5891);
and U9114 (N_9114,N_6529,N_7198);
xor U9115 (N_9115,N_7140,N_6805);
and U9116 (N_9116,N_6266,N_6654);
or U9117 (N_9117,N_6619,N_6138);
or U9118 (N_9118,N_6095,N_7124);
nor U9119 (N_9119,N_5864,N_5895);
nand U9120 (N_9120,N_7458,N_5471);
nand U9121 (N_9121,N_7421,N_7235);
nor U9122 (N_9122,N_6019,N_6162);
and U9123 (N_9123,N_5801,N_5710);
or U9124 (N_9124,N_5464,N_7372);
and U9125 (N_9125,N_6773,N_6276);
xnor U9126 (N_9126,N_5278,N_5673);
nor U9127 (N_9127,N_5737,N_6245);
nor U9128 (N_9128,N_6625,N_5409);
nor U9129 (N_9129,N_6056,N_5313);
nand U9130 (N_9130,N_5386,N_5825);
and U9131 (N_9131,N_5552,N_6029);
and U9132 (N_9132,N_5956,N_6234);
and U9133 (N_9133,N_5111,N_7166);
nand U9134 (N_9134,N_6153,N_5773);
nor U9135 (N_9135,N_5092,N_6871);
or U9136 (N_9136,N_5671,N_7385);
or U9137 (N_9137,N_5800,N_6186);
and U9138 (N_9138,N_5077,N_6072);
and U9139 (N_9139,N_6980,N_7394);
and U9140 (N_9140,N_5761,N_7161);
or U9141 (N_9141,N_6443,N_5812);
and U9142 (N_9142,N_6219,N_6115);
or U9143 (N_9143,N_5121,N_5398);
and U9144 (N_9144,N_7119,N_5850);
nor U9145 (N_9145,N_5254,N_7411);
and U9146 (N_9146,N_5925,N_6132);
or U9147 (N_9147,N_7284,N_7069);
and U9148 (N_9148,N_6794,N_6150);
nor U9149 (N_9149,N_6271,N_7441);
and U9150 (N_9150,N_6859,N_7382);
xor U9151 (N_9151,N_6602,N_5750);
nand U9152 (N_9152,N_6410,N_6837);
nor U9153 (N_9153,N_5368,N_6360);
or U9154 (N_9154,N_7248,N_5138);
and U9155 (N_9155,N_6544,N_6889);
and U9156 (N_9156,N_5082,N_6871);
or U9157 (N_9157,N_5202,N_5706);
and U9158 (N_9158,N_5590,N_6566);
and U9159 (N_9159,N_7338,N_5819);
and U9160 (N_9160,N_5734,N_6638);
nand U9161 (N_9161,N_5013,N_6804);
nand U9162 (N_9162,N_6150,N_6779);
and U9163 (N_9163,N_6084,N_7292);
or U9164 (N_9164,N_6562,N_5360);
nand U9165 (N_9165,N_7107,N_7385);
or U9166 (N_9166,N_6306,N_7055);
and U9167 (N_9167,N_5688,N_6650);
xnor U9168 (N_9168,N_6483,N_5894);
nor U9169 (N_9169,N_6695,N_5972);
and U9170 (N_9170,N_5701,N_6303);
nand U9171 (N_9171,N_6565,N_5961);
and U9172 (N_9172,N_6348,N_5714);
and U9173 (N_9173,N_6040,N_6530);
and U9174 (N_9174,N_6900,N_6177);
and U9175 (N_9175,N_6306,N_6241);
and U9176 (N_9176,N_6493,N_6495);
nor U9177 (N_9177,N_5969,N_5006);
or U9178 (N_9178,N_6118,N_6689);
and U9179 (N_9179,N_7045,N_5972);
and U9180 (N_9180,N_5163,N_5298);
nor U9181 (N_9181,N_7369,N_5074);
nand U9182 (N_9182,N_5182,N_5661);
or U9183 (N_9183,N_5786,N_6950);
or U9184 (N_9184,N_7307,N_5293);
and U9185 (N_9185,N_6034,N_6893);
nor U9186 (N_9186,N_5552,N_5738);
nor U9187 (N_9187,N_5187,N_5028);
nor U9188 (N_9188,N_5277,N_7267);
nor U9189 (N_9189,N_5538,N_6997);
nand U9190 (N_9190,N_7305,N_6772);
nand U9191 (N_9191,N_6612,N_5702);
nand U9192 (N_9192,N_5996,N_6121);
or U9193 (N_9193,N_5012,N_7268);
or U9194 (N_9194,N_5725,N_6230);
nand U9195 (N_9195,N_7378,N_7421);
or U9196 (N_9196,N_6830,N_6017);
nand U9197 (N_9197,N_5598,N_6182);
or U9198 (N_9198,N_5630,N_6647);
or U9199 (N_9199,N_5976,N_6697);
and U9200 (N_9200,N_5773,N_5289);
nor U9201 (N_9201,N_6326,N_7076);
nor U9202 (N_9202,N_5402,N_6449);
nor U9203 (N_9203,N_6768,N_7379);
or U9204 (N_9204,N_6701,N_5343);
or U9205 (N_9205,N_6086,N_5532);
nor U9206 (N_9206,N_5266,N_6208);
nand U9207 (N_9207,N_5702,N_7168);
or U9208 (N_9208,N_6433,N_6426);
or U9209 (N_9209,N_6936,N_7027);
and U9210 (N_9210,N_6948,N_6768);
nand U9211 (N_9211,N_5590,N_6635);
nor U9212 (N_9212,N_6089,N_7138);
or U9213 (N_9213,N_6844,N_7450);
and U9214 (N_9214,N_5602,N_6745);
or U9215 (N_9215,N_6198,N_7248);
nand U9216 (N_9216,N_5664,N_6259);
nor U9217 (N_9217,N_5307,N_6928);
and U9218 (N_9218,N_5489,N_5797);
nand U9219 (N_9219,N_7221,N_5313);
nand U9220 (N_9220,N_7404,N_5106);
or U9221 (N_9221,N_6346,N_5900);
nor U9222 (N_9222,N_6113,N_7379);
nand U9223 (N_9223,N_6867,N_7196);
or U9224 (N_9224,N_6604,N_6098);
nor U9225 (N_9225,N_5802,N_6381);
and U9226 (N_9226,N_6110,N_5472);
nor U9227 (N_9227,N_6963,N_6518);
or U9228 (N_9228,N_6427,N_5179);
nand U9229 (N_9229,N_7450,N_5927);
nand U9230 (N_9230,N_5137,N_5679);
nor U9231 (N_9231,N_5631,N_5822);
nor U9232 (N_9232,N_7335,N_5439);
and U9233 (N_9233,N_5556,N_5681);
or U9234 (N_9234,N_5690,N_7196);
or U9235 (N_9235,N_6322,N_5991);
nor U9236 (N_9236,N_5276,N_7310);
or U9237 (N_9237,N_6969,N_6866);
and U9238 (N_9238,N_7076,N_7360);
nand U9239 (N_9239,N_6110,N_5507);
nand U9240 (N_9240,N_6686,N_6985);
nor U9241 (N_9241,N_7178,N_7277);
nor U9242 (N_9242,N_5549,N_6720);
nor U9243 (N_9243,N_5360,N_6923);
xnor U9244 (N_9244,N_5652,N_5720);
nand U9245 (N_9245,N_5238,N_7334);
nor U9246 (N_9246,N_5865,N_5243);
and U9247 (N_9247,N_6403,N_5287);
and U9248 (N_9248,N_5837,N_5236);
or U9249 (N_9249,N_5156,N_6779);
or U9250 (N_9250,N_5440,N_5903);
and U9251 (N_9251,N_7161,N_5042);
nand U9252 (N_9252,N_6062,N_6519);
nand U9253 (N_9253,N_6161,N_7217);
or U9254 (N_9254,N_5996,N_6754);
nand U9255 (N_9255,N_7469,N_5130);
nand U9256 (N_9256,N_5522,N_7039);
or U9257 (N_9257,N_6954,N_7019);
or U9258 (N_9258,N_5051,N_5126);
nor U9259 (N_9259,N_5926,N_7314);
and U9260 (N_9260,N_5461,N_5404);
and U9261 (N_9261,N_7202,N_6733);
or U9262 (N_9262,N_5963,N_7333);
or U9263 (N_9263,N_5142,N_6798);
nand U9264 (N_9264,N_6689,N_5723);
nand U9265 (N_9265,N_6869,N_7380);
and U9266 (N_9266,N_6150,N_7238);
nand U9267 (N_9267,N_7445,N_6976);
or U9268 (N_9268,N_6809,N_5511);
nand U9269 (N_9269,N_6846,N_7360);
or U9270 (N_9270,N_6992,N_6904);
and U9271 (N_9271,N_5498,N_5486);
and U9272 (N_9272,N_6702,N_5973);
nand U9273 (N_9273,N_7424,N_7036);
or U9274 (N_9274,N_5502,N_5077);
nor U9275 (N_9275,N_7306,N_7022);
or U9276 (N_9276,N_7486,N_6336);
or U9277 (N_9277,N_7127,N_6656);
or U9278 (N_9278,N_5644,N_5107);
nand U9279 (N_9279,N_5668,N_7045);
nand U9280 (N_9280,N_5661,N_5094);
nand U9281 (N_9281,N_6249,N_6344);
or U9282 (N_9282,N_5014,N_5828);
nand U9283 (N_9283,N_5878,N_5374);
nand U9284 (N_9284,N_5436,N_7330);
nor U9285 (N_9285,N_7324,N_6295);
and U9286 (N_9286,N_6810,N_6535);
nand U9287 (N_9287,N_6878,N_5661);
or U9288 (N_9288,N_5288,N_6494);
and U9289 (N_9289,N_6106,N_5781);
nand U9290 (N_9290,N_5407,N_7097);
or U9291 (N_9291,N_6031,N_7362);
and U9292 (N_9292,N_7187,N_6510);
nand U9293 (N_9293,N_5301,N_6324);
nor U9294 (N_9294,N_7380,N_6049);
nand U9295 (N_9295,N_6818,N_6510);
nand U9296 (N_9296,N_5942,N_5895);
nand U9297 (N_9297,N_7017,N_5500);
and U9298 (N_9298,N_7275,N_5397);
and U9299 (N_9299,N_5721,N_5000);
nand U9300 (N_9300,N_6003,N_7135);
and U9301 (N_9301,N_7448,N_6248);
nor U9302 (N_9302,N_5397,N_7405);
or U9303 (N_9303,N_5325,N_5389);
or U9304 (N_9304,N_6747,N_6127);
or U9305 (N_9305,N_5264,N_6041);
nor U9306 (N_9306,N_7097,N_6923);
and U9307 (N_9307,N_7461,N_7474);
or U9308 (N_9308,N_7415,N_5655);
or U9309 (N_9309,N_6323,N_7134);
nor U9310 (N_9310,N_5770,N_6146);
nand U9311 (N_9311,N_5130,N_6379);
or U9312 (N_9312,N_5980,N_6829);
nor U9313 (N_9313,N_6058,N_7068);
nor U9314 (N_9314,N_5729,N_7395);
and U9315 (N_9315,N_6030,N_7313);
nor U9316 (N_9316,N_6264,N_5402);
and U9317 (N_9317,N_5435,N_6278);
nand U9318 (N_9318,N_5502,N_7264);
nor U9319 (N_9319,N_6825,N_6639);
xnor U9320 (N_9320,N_7250,N_5792);
and U9321 (N_9321,N_7312,N_5471);
nor U9322 (N_9322,N_5869,N_5693);
and U9323 (N_9323,N_5598,N_6468);
nand U9324 (N_9324,N_6770,N_7281);
nor U9325 (N_9325,N_6633,N_6459);
nor U9326 (N_9326,N_7135,N_5284);
nand U9327 (N_9327,N_5901,N_5102);
and U9328 (N_9328,N_6963,N_6198);
or U9329 (N_9329,N_6049,N_7287);
and U9330 (N_9330,N_5117,N_6411);
nor U9331 (N_9331,N_5603,N_6283);
and U9332 (N_9332,N_5978,N_7474);
or U9333 (N_9333,N_5469,N_6205);
nand U9334 (N_9334,N_6174,N_6326);
nand U9335 (N_9335,N_5525,N_6341);
xor U9336 (N_9336,N_7426,N_7267);
or U9337 (N_9337,N_5142,N_5685);
nand U9338 (N_9338,N_5686,N_5009);
nor U9339 (N_9339,N_6920,N_7312);
nand U9340 (N_9340,N_6239,N_5317);
nor U9341 (N_9341,N_6518,N_5103);
nor U9342 (N_9342,N_5713,N_5340);
xor U9343 (N_9343,N_7423,N_5914);
or U9344 (N_9344,N_6622,N_6561);
nor U9345 (N_9345,N_7372,N_5463);
and U9346 (N_9346,N_5170,N_7343);
and U9347 (N_9347,N_5923,N_6661);
nand U9348 (N_9348,N_6271,N_6395);
xor U9349 (N_9349,N_5710,N_7253);
nor U9350 (N_9350,N_5300,N_5239);
nor U9351 (N_9351,N_6128,N_6948);
or U9352 (N_9352,N_7403,N_7068);
or U9353 (N_9353,N_5229,N_5040);
or U9354 (N_9354,N_6527,N_5773);
nor U9355 (N_9355,N_6326,N_7317);
or U9356 (N_9356,N_6778,N_7450);
nand U9357 (N_9357,N_5164,N_6662);
xnor U9358 (N_9358,N_5734,N_5936);
nor U9359 (N_9359,N_6957,N_7188);
or U9360 (N_9360,N_5906,N_7277);
nand U9361 (N_9361,N_7061,N_6257);
and U9362 (N_9362,N_6674,N_5914);
and U9363 (N_9363,N_6648,N_5934);
nand U9364 (N_9364,N_5840,N_6174);
or U9365 (N_9365,N_5668,N_6124);
nand U9366 (N_9366,N_5857,N_7195);
nand U9367 (N_9367,N_5181,N_7340);
nand U9368 (N_9368,N_6661,N_5232);
or U9369 (N_9369,N_5684,N_6685);
and U9370 (N_9370,N_6596,N_7478);
and U9371 (N_9371,N_5704,N_5174);
nand U9372 (N_9372,N_5914,N_6597);
and U9373 (N_9373,N_5539,N_6700);
and U9374 (N_9374,N_6458,N_5052);
or U9375 (N_9375,N_5441,N_7458);
and U9376 (N_9376,N_7246,N_6367);
nand U9377 (N_9377,N_7442,N_5299);
or U9378 (N_9378,N_6744,N_6374);
or U9379 (N_9379,N_6597,N_6990);
or U9380 (N_9380,N_5602,N_5250);
nor U9381 (N_9381,N_5788,N_7076);
and U9382 (N_9382,N_6906,N_6314);
nor U9383 (N_9383,N_6544,N_5190);
and U9384 (N_9384,N_7312,N_5038);
or U9385 (N_9385,N_7109,N_6837);
and U9386 (N_9386,N_6918,N_5158);
and U9387 (N_9387,N_5323,N_6811);
or U9388 (N_9388,N_6496,N_5961);
nor U9389 (N_9389,N_5996,N_6273);
or U9390 (N_9390,N_6570,N_7195);
nand U9391 (N_9391,N_5482,N_6196);
nor U9392 (N_9392,N_5236,N_6799);
nor U9393 (N_9393,N_5701,N_6001);
or U9394 (N_9394,N_6140,N_6557);
or U9395 (N_9395,N_5732,N_5919);
and U9396 (N_9396,N_5924,N_6588);
nand U9397 (N_9397,N_7192,N_7452);
or U9398 (N_9398,N_6699,N_5020);
and U9399 (N_9399,N_7176,N_5124);
or U9400 (N_9400,N_5520,N_7379);
and U9401 (N_9401,N_7250,N_7094);
and U9402 (N_9402,N_6321,N_5783);
and U9403 (N_9403,N_6665,N_7268);
and U9404 (N_9404,N_5631,N_5324);
and U9405 (N_9405,N_6465,N_7246);
nand U9406 (N_9406,N_6875,N_6486);
nor U9407 (N_9407,N_6369,N_5360);
nand U9408 (N_9408,N_7340,N_5784);
xor U9409 (N_9409,N_5570,N_5836);
nor U9410 (N_9410,N_5837,N_7494);
nor U9411 (N_9411,N_5893,N_6223);
and U9412 (N_9412,N_5732,N_6051);
nand U9413 (N_9413,N_7190,N_6278);
nand U9414 (N_9414,N_6206,N_5863);
and U9415 (N_9415,N_5624,N_7358);
or U9416 (N_9416,N_6812,N_6411);
or U9417 (N_9417,N_7352,N_6320);
xnor U9418 (N_9418,N_6690,N_7325);
and U9419 (N_9419,N_7198,N_5431);
nand U9420 (N_9420,N_5626,N_5017);
or U9421 (N_9421,N_5204,N_6014);
or U9422 (N_9422,N_5435,N_6292);
or U9423 (N_9423,N_5442,N_6633);
nand U9424 (N_9424,N_5148,N_7070);
nor U9425 (N_9425,N_5707,N_5974);
and U9426 (N_9426,N_6253,N_6722);
or U9427 (N_9427,N_5559,N_5588);
nor U9428 (N_9428,N_7032,N_5636);
nand U9429 (N_9429,N_6630,N_5480);
and U9430 (N_9430,N_6029,N_5699);
nor U9431 (N_9431,N_6284,N_6696);
and U9432 (N_9432,N_5491,N_7134);
nand U9433 (N_9433,N_5601,N_5839);
nand U9434 (N_9434,N_7258,N_5531);
nand U9435 (N_9435,N_6654,N_6073);
nand U9436 (N_9436,N_6474,N_5652);
and U9437 (N_9437,N_6210,N_5673);
nand U9438 (N_9438,N_5976,N_6598);
or U9439 (N_9439,N_6959,N_6520);
and U9440 (N_9440,N_5109,N_6660);
or U9441 (N_9441,N_7446,N_5100);
xnor U9442 (N_9442,N_5229,N_5685);
and U9443 (N_9443,N_6002,N_6428);
nand U9444 (N_9444,N_6969,N_5148);
or U9445 (N_9445,N_5658,N_5529);
or U9446 (N_9446,N_6397,N_5470);
or U9447 (N_9447,N_5158,N_5606);
and U9448 (N_9448,N_6095,N_5094);
and U9449 (N_9449,N_5372,N_6132);
nand U9450 (N_9450,N_7147,N_5703);
nor U9451 (N_9451,N_7232,N_6206);
nand U9452 (N_9452,N_5915,N_5792);
and U9453 (N_9453,N_5662,N_6500);
or U9454 (N_9454,N_5822,N_7439);
nand U9455 (N_9455,N_6502,N_5557);
and U9456 (N_9456,N_6707,N_7065);
and U9457 (N_9457,N_6149,N_5840);
nand U9458 (N_9458,N_5281,N_5394);
nor U9459 (N_9459,N_7122,N_5122);
and U9460 (N_9460,N_7318,N_6285);
nor U9461 (N_9461,N_7464,N_5217);
nor U9462 (N_9462,N_6236,N_5631);
nor U9463 (N_9463,N_6195,N_5117);
nand U9464 (N_9464,N_6287,N_6625);
and U9465 (N_9465,N_7072,N_7117);
nand U9466 (N_9466,N_6813,N_7342);
nand U9467 (N_9467,N_5332,N_7424);
nor U9468 (N_9468,N_5521,N_5288);
nand U9469 (N_9469,N_7069,N_7359);
nand U9470 (N_9470,N_6876,N_5797);
nand U9471 (N_9471,N_6757,N_6758);
and U9472 (N_9472,N_6916,N_6405);
and U9473 (N_9473,N_5779,N_5849);
nor U9474 (N_9474,N_6889,N_6440);
or U9475 (N_9475,N_6477,N_7178);
xnor U9476 (N_9476,N_6748,N_5475);
nand U9477 (N_9477,N_6506,N_6446);
nor U9478 (N_9478,N_5598,N_6723);
and U9479 (N_9479,N_6761,N_6322);
and U9480 (N_9480,N_5886,N_7496);
and U9481 (N_9481,N_5010,N_6213);
or U9482 (N_9482,N_7344,N_5338);
nand U9483 (N_9483,N_5438,N_5146);
xnor U9484 (N_9484,N_5289,N_6262);
nor U9485 (N_9485,N_5833,N_6996);
nor U9486 (N_9486,N_5853,N_7133);
and U9487 (N_9487,N_7376,N_5031);
nand U9488 (N_9488,N_5211,N_6906);
nor U9489 (N_9489,N_6534,N_5534);
nand U9490 (N_9490,N_6916,N_5820);
nor U9491 (N_9491,N_6378,N_6827);
or U9492 (N_9492,N_5300,N_5796);
or U9493 (N_9493,N_5647,N_6407);
and U9494 (N_9494,N_7177,N_5087);
nor U9495 (N_9495,N_5551,N_6830);
nand U9496 (N_9496,N_5096,N_6729);
or U9497 (N_9497,N_6238,N_5692);
nand U9498 (N_9498,N_7061,N_6572);
nor U9499 (N_9499,N_5473,N_6129);
nand U9500 (N_9500,N_5753,N_7209);
nand U9501 (N_9501,N_6486,N_6644);
or U9502 (N_9502,N_7207,N_5908);
nand U9503 (N_9503,N_7029,N_6077);
and U9504 (N_9504,N_7451,N_5857);
or U9505 (N_9505,N_5179,N_7100);
and U9506 (N_9506,N_5143,N_5839);
nor U9507 (N_9507,N_6271,N_5768);
nand U9508 (N_9508,N_5809,N_5957);
and U9509 (N_9509,N_7381,N_6863);
or U9510 (N_9510,N_7494,N_7088);
nand U9511 (N_9511,N_5213,N_5018);
xnor U9512 (N_9512,N_6742,N_5035);
nand U9513 (N_9513,N_7459,N_6565);
nand U9514 (N_9514,N_6700,N_5188);
and U9515 (N_9515,N_5583,N_7129);
and U9516 (N_9516,N_6348,N_6147);
nand U9517 (N_9517,N_6243,N_7349);
nor U9518 (N_9518,N_6556,N_5543);
and U9519 (N_9519,N_7109,N_6438);
and U9520 (N_9520,N_6178,N_5022);
nor U9521 (N_9521,N_5781,N_6093);
nand U9522 (N_9522,N_5107,N_5228);
nor U9523 (N_9523,N_6512,N_5063);
nand U9524 (N_9524,N_5687,N_5824);
nand U9525 (N_9525,N_5546,N_7083);
nor U9526 (N_9526,N_6863,N_6110);
nand U9527 (N_9527,N_5357,N_6104);
and U9528 (N_9528,N_7018,N_5151);
nand U9529 (N_9529,N_5355,N_5655);
nor U9530 (N_9530,N_6269,N_5073);
or U9531 (N_9531,N_5382,N_7417);
nand U9532 (N_9532,N_7271,N_7465);
nand U9533 (N_9533,N_5892,N_5132);
and U9534 (N_9534,N_6427,N_6307);
and U9535 (N_9535,N_6761,N_6626);
and U9536 (N_9536,N_6050,N_5005);
nor U9537 (N_9537,N_5559,N_5788);
or U9538 (N_9538,N_7124,N_7309);
and U9539 (N_9539,N_5633,N_6626);
nand U9540 (N_9540,N_5449,N_5615);
nand U9541 (N_9541,N_5131,N_6296);
nand U9542 (N_9542,N_5395,N_6205);
or U9543 (N_9543,N_7128,N_5804);
and U9544 (N_9544,N_7375,N_5509);
nand U9545 (N_9545,N_6804,N_7248);
or U9546 (N_9546,N_6810,N_6549);
nor U9547 (N_9547,N_6813,N_5784);
or U9548 (N_9548,N_5474,N_6809);
and U9549 (N_9549,N_6759,N_6845);
and U9550 (N_9550,N_5601,N_7475);
or U9551 (N_9551,N_6883,N_5160);
nand U9552 (N_9552,N_6258,N_5269);
nand U9553 (N_9553,N_5474,N_5685);
or U9554 (N_9554,N_6471,N_6684);
nand U9555 (N_9555,N_7200,N_6561);
nand U9556 (N_9556,N_7414,N_7381);
xor U9557 (N_9557,N_5151,N_6238);
nand U9558 (N_9558,N_7124,N_7148);
or U9559 (N_9559,N_6409,N_7039);
nor U9560 (N_9560,N_5892,N_6653);
nor U9561 (N_9561,N_7424,N_5701);
nand U9562 (N_9562,N_6012,N_7496);
nand U9563 (N_9563,N_5342,N_7303);
and U9564 (N_9564,N_6363,N_6383);
nand U9565 (N_9565,N_6287,N_7439);
nand U9566 (N_9566,N_6906,N_5184);
nand U9567 (N_9567,N_5531,N_5586);
nand U9568 (N_9568,N_6606,N_5254);
nor U9569 (N_9569,N_6173,N_6194);
or U9570 (N_9570,N_5756,N_6899);
or U9571 (N_9571,N_5630,N_6952);
and U9572 (N_9572,N_7320,N_6276);
nor U9573 (N_9573,N_6707,N_7449);
nand U9574 (N_9574,N_5025,N_6983);
nand U9575 (N_9575,N_7382,N_5831);
nand U9576 (N_9576,N_5462,N_5447);
or U9577 (N_9577,N_5398,N_6265);
nor U9578 (N_9578,N_6566,N_6045);
xor U9579 (N_9579,N_5263,N_6728);
nand U9580 (N_9580,N_7003,N_5495);
nand U9581 (N_9581,N_6729,N_7105);
or U9582 (N_9582,N_6390,N_6937);
nand U9583 (N_9583,N_5728,N_6393);
or U9584 (N_9584,N_6201,N_5468);
and U9585 (N_9585,N_7369,N_6394);
or U9586 (N_9586,N_7074,N_5782);
and U9587 (N_9587,N_5140,N_5782);
and U9588 (N_9588,N_5793,N_5742);
nor U9589 (N_9589,N_5541,N_7430);
or U9590 (N_9590,N_5591,N_7382);
or U9591 (N_9591,N_5790,N_7086);
or U9592 (N_9592,N_6469,N_6122);
or U9593 (N_9593,N_6729,N_6423);
nand U9594 (N_9594,N_7161,N_7023);
and U9595 (N_9595,N_6768,N_7123);
or U9596 (N_9596,N_6518,N_5643);
nand U9597 (N_9597,N_6432,N_6407);
nor U9598 (N_9598,N_7071,N_5544);
and U9599 (N_9599,N_5133,N_5801);
and U9600 (N_9600,N_7408,N_7066);
nand U9601 (N_9601,N_5914,N_6314);
and U9602 (N_9602,N_7218,N_6505);
nand U9603 (N_9603,N_5802,N_5804);
or U9604 (N_9604,N_6559,N_5956);
or U9605 (N_9605,N_6621,N_6613);
nand U9606 (N_9606,N_5930,N_6015);
and U9607 (N_9607,N_7279,N_6198);
or U9608 (N_9608,N_6942,N_6743);
or U9609 (N_9609,N_5688,N_6518);
and U9610 (N_9610,N_7003,N_5889);
nand U9611 (N_9611,N_5082,N_6048);
and U9612 (N_9612,N_6591,N_6051);
nand U9613 (N_9613,N_7122,N_7388);
or U9614 (N_9614,N_5078,N_5995);
and U9615 (N_9615,N_5148,N_6282);
and U9616 (N_9616,N_5842,N_6303);
and U9617 (N_9617,N_5348,N_6056);
nand U9618 (N_9618,N_6414,N_5978);
nor U9619 (N_9619,N_5852,N_6435);
nor U9620 (N_9620,N_6257,N_5938);
xor U9621 (N_9621,N_6635,N_7318);
or U9622 (N_9622,N_7020,N_6579);
or U9623 (N_9623,N_7067,N_5832);
nand U9624 (N_9624,N_6248,N_5457);
or U9625 (N_9625,N_5102,N_5918);
nand U9626 (N_9626,N_7060,N_6197);
nand U9627 (N_9627,N_5198,N_6475);
and U9628 (N_9628,N_5134,N_6276);
or U9629 (N_9629,N_7145,N_6926);
and U9630 (N_9630,N_5209,N_5328);
nor U9631 (N_9631,N_5922,N_7099);
nand U9632 (N_9632,N_5603,N_5833);
nand U9633 (N_9633,N_7051,N_7078);
or U9634 (N_9634,N_6695,N_7115);
and U9635 (N_9635,N_6952,N_6125);
and U9636 (N_9636,N_7125,N_5136);
or U9637 (N_9637,N_7452,N_5090);
and U9638 (N_9638,N_5803,N_5452);
nand U9639 (N_9639,N_6132,N_5374);
nor U9640 (N_9640,N_7491,N_5863);
or U9641 (N_9641,N_7397,N_6197);
nand U9642 (N_9642,N_6075,N_6635);
or U9643 (N_9643,N_6501,N_6037);
xor U9644 (N_9644,N_6155,N_7482);
nor U9645 (N_9645,N_5547,N_7410);
and U9646 (N_9646,N_6494,N_5446);
or U9647 (N_9647,N_6305,N_5996);
xnor U9648 (N_9648,N_7155,N_5003);
nor U9649 (N_9649,N_6464,N_5947);
nand U9650 (N_9650,N_5213,N_5369);
and U9651 (N_9651,N_7392,N_6809);
or U9652 (N_9652,N_5010,N_5645);
and U9653 (N_9653,N_7005,N_6591);
or U9654 (N_9654,N_7201,N_6592);
or U9655 (N_9655,N_5724,N_6291);
nor U9656 (N_9656,N_6335,N_5538);
and U9657 (N_9657,N_5283,N_5194);
nor U9658 (N_9658,N_7231,N_6915);
nand U9659 (N_9659,N_6720,N_5085);
and U9660 (N_9660,N_5991,N_7441);
and U9661 (N_9661,N_5733,N_5385);
nor U9662 (N_9662,N_5415,N_7081);
and U9663 (N_9663,N_6128,N_6752);
and U9664 (N_9664,N_6576,N_5072);
nand U9665 (N_9665,N_7378,N_6714);
or U9666 (N_9666,N_6621,N_6860);
nand U9667 (N_9667,N_5631,N_7417);
or U9668 (N_9668,N_6429,N_5849);
or U9669 (N_9669,N_6243,N_7270);
or U9670 (N_9670,N_5682,N_6506);
nor U9671 (N_9671,N_7329,N_7075);
or U9672 (N_9672,N_7397,N_5137);
and U9673 (N_9673,N_6938,N_7170);
nor U9674 (N_9674,N_6971,N_6156);
and U9675 (N_9675,N_7259,N_7170);
and U9676 (N_9676,N_6168,N_5197);
and U9677 (N_9677,N_6267,N_7001);
or U9678 (N_9678,N_5525,N_7136);
or U9679 (N_9679,N_5099,N_5331);
nand U9680 (N_9680,N_5163,N_5623);
and U9681 (N_9681,N_7395,N_5220);
and U9682 (N_9682,N_5888,N_5105);
nor U9683 (N_9683,N_5057,N_6021);
nand U9684 (N_9684,N_5544,N_7404);
or U9685 (N_9685,N_6513,N_5945);
or U9686 (N_9686,N_6455,N_5283);
xor U9687 (N_9687,N_5925,N_5033);
or U9688 (N_9688,N_6749,N_6331);
or U9689 (N_9689,N_6113,N_6443);
nor U9690 (N_9690,N_5618,N_6573);
nor U9691 (N_9691,N_7218,N_6705);
and U9692 (N_9692,N_6382,N_6998);
and U9693 (N_9693,N_5252,N_5143);
or U9694 (N_9694,N_6487,N_5596);
and U9695 (N_9695,N_5499,N_6796);
and U9696 (N_9696,N_6724,N_5252);
nor U9697 (N_9697,N_6687,N_5645);
xnor U9698 (N_9698,N_5763,N_5005);
or U9699 (N_9699,N_6542,N_5510);
or U9700 (N_9700,N_5290,N_5718);
nor U9701 (N_9701,N_6450,N_5529);
nand U9702 (N_9702,N_6002,N_5439);
and U9703 (N_9703,N_7325,N_5217);
or U9704 (N_9704,N_7379,N_6680);
nor U9705 (N_9705,N_5385,N_5447);
nand U9706 (N_9706,N_6627,N_7175);
and U9707 (N_9707,N_7103,N_6043);
nand U9708 (N_9708,N_6970,N_5634);
and U9709 (N_9709,N_6595,N_5368);
or U9710 (N_9710,N_6938,N_5092);
nor U9711 (N_9711,N_6103,N_6414);
and U9712 (N_9712,N_5387,N_7286);
and U9713 (N_9713,N_7323,N_7280);
and U9714 (N_9714,N_5236,N_5093);
nand U9715 (N_9715,N_7241,N_5053);
nand U9716 (N_9716,N_5920,N_7222);
or U9717 (N_9717,N_5184,N_5150);
nor U9718 (N_9718,N_5969,N_7143);
nand U9719 (N_9719,N_5019,N_6502);
nand U9720 (N_9720,N_6367,N_7420);
nand U9721 (N_9721,N_7428,N_6399);
and U9722 (N_9722,N_6756,N_6064);
nor U9723 (N_9723,N_5026,N_7147);
nor U9724 (N_9724,N_5779,N_6574);
or U9725 (N_9725,N_6725,N_5321);
and U9726 (N_9726,N_5922,N_6625);
or U9727 (N_9727,N_7005,N_6255);
nor U9728 (N_9728,N_7080,N_6178);
nand U9729 (N_9729,N_6820,N_6379);
xor U9730 (N_9730,N_6069,N_6182);
or U9731 (N_9731,N_6376,N_6464);
and U9732 (N_9732,N_6901,N_6930);
nand U9733 (N_9733,N_5157,N_5951);
nand U9734 (N_9734,N_6137,N_7299);
or U9735 (N_9735,N_6300,N_5021);
or U9736 (N_9736,N_5951,N_5439);
or U9737 (N_9737,N_5091,N_5188);
or U9738 (N_9738,N_6495,N_6003);
nand U9739 (N_9739,N_6909,N_6324);
and U9740 (N_9740,N_5849,N_5850);
or U9741 (N_9741,N_5352,N_7237);
nor U9742 (N_9742,N_6714,N_6054);
and U9743 (N_9743,N_6860,N_5531);
nand U9744 (N_9744,N_7079,N_5100);
nand U9745 (N_9745,N_5885,N_7050);
xnor U9746 (N_9746,N_6046,N_6336);
and U9747 (N_9747,N_6997,N_5948);
and U9748 (N_9748,N_6409,N_7426);
and U9749 (N_9749,N_5791,N_5781);
xnor U9750 (N_9750,N_7149,N_6406);
nand U9751 (N_9751,N_6542,N_7358);
or U9752 (N_9752,N_5683,N_6418);
or U9753 (N_9753,N_6829,N_7017);
nor U9754 (N_9754,N_5616,N_7454);
nor U9755 (N_9755,N_5429,N_5041);
nand U9756 (N_9756,N_5882,N_6286);
nor U9757 (N_9757,N_7316,N_5952);
nand U9758 (N_9758,N_6433,N_7047);
nor U9759 (N_9759,N_6784,N_6205);
or U9760 (N_9760,N_5256,N_5137);
nor U9761 (N_9761,N_7382,N_5091);
nand U9762 (N_9762,N_5260,N_6522);
and U9763 (N_9763,N_5162,N_5727);
or U9764 (N_9764,N_5995,N_6106);
nor U9765 (N_9765,N_5794,N_6484);
nand U9766 (N_9766,N_7203,N_7283);
nand U9767 (N_9767,N_6214,N_5969);
or U9768 (N_9768,N_5803,N_6726);
and U9769 (N_9769,N_6544,N_5682);
nor U9770 (N_9770,N_6599,N_6109);
or U9771 (N_9771,N_7236,N_6216);
nor U9772 (N_9772,N_5405,N_6357);
nor U9773 (N_9773,N_7233,N_6168);
nand U9774 (N_9774,N_5704,N_6214);
nor U9775 (N_9775,N_6564,N_6759);
and U9776 (N_9776,N_7449,N_5848);
or U9777 (N_9777,N_5365,N_5301);
or U9778 (N_9778,N_7261,N_6335);
nor U9779 (N_9779,N_6811,N_7427);
nand U9780 (N_9780,N_7067,N_5237);
nand U9781 (N_9781,N_6395,N_6421);
nand U9782 (N_9782,N_6973,N_5267);
xnor U9783 (N_9783,N_7143,N_5780);
or U9784 (N_9784,N_7454,N_5501);
nor U9785 (N_9785,N_5810,N_7241);
xor U9786 (N_9786,N_7206,N_7432);
nand U9787 (N_9787,N_5770,N_5525);
nand U9788 (N_9788,N_6986,N_6645);
nor U9789 (N_9789,N_6024,N_5530);
nand U9790 (N_9790,N_6797,N_6779);
or U9791 (N_9791,N_5078,N_6020);
or U9792 (N_9792,N_5621,N_5277);
xnor U9793 (N_9793,N_5696,N_5976);
or U9794 (N_9794,N_5722,N_5215);
and U9795 (N_9795,N_6039,N_6636);
nand U9796 (N_9796,N_7200,N_6379);
xor U9797 (N_9797,N_5924,N_6118);
and U9798 (N_9798,N_6412,N_5769);
nor U9799 (N_9799,N_6038,N_6355);
or U9800 (N_9800,N_7393,N_5871);
nand U9801 (N_9801,N_6656,N_6047);
or U9802 (N_9802,N_6019,N_5387);
nor U9803 (N_9803,N_5356,N_5384);
or U9804 (N_9804,N_5072,N_5351);
or U9805 (N_9805,N_6381,N_5373);
nor U9806 (N_9806,N_6885,N_7099);
and U9807 (N_9807,N_5878,N_7191);
or U9808 (N_9808,N_5123,N_5773);
nor U9809 (N_9809,N_5680,N_5324);
nor U9810 (N_9810,N_5411,N_5474);
nand U9811 (N_9811,N_5164,N_6851);
and U9812 (N_9812,N_7037,N_6130);
and U9813 (N_9813,N_5772,N_5543);
and U9814 (N_9814,N_7218,N_6882);
nand U9815 (N_9815,N_6775,N_5647);
or U9816 (N_9816,N_6733,N_6051);
and U9817 (N_9817,N_7310,N_5035);
nand U9818 (N_9818,N_5255,N_7114);
and U9819 (N_9819,N_5418,N_5210);
and U9820 (N_9820,N_6471,N_5218);
nor U9821 (N_9821,N_7439,N_6708);
nor U9822 (N_9822,N_5598,N_6206);
xor U9823 (N_9823,N_7473,N_7023);
and U9824 (N_9824,N_5978,N_6388);
and U9825 (N_9825,N_5565,N_5518);
and U9826 (N_9826,N_5152,N_5643);
and U9827 (N_9827,N_6625,N_6665);
nand U9828 (N_9828,N_7298,N_6243);
or U9829 (N_9829,N_7299,N_7011);
or U9830 (N_9830,N_6420,N_7250);
or U9831 (N_9831,N_6644,N_7104);
or U9832 (N_9832,N_5600,N_7444);
nand U9833 (N_9833,N_6444,N_6249);
nand U9834 (N_9834,N_5935,N_5097);
nand U9835 (N_9835,N_5671,N_5323);
nor U9836 (N_9836,N_5010,N_6143);
and U9837 (N_9837,N_5978,N_7080);
and U9838 (N_9838,N_5452,N_6908);
or U9839 (N_9839,N_6866,N_5234);
and U9840 (N_9840,N_5983,N_7318);
nand U9841 (N_9841,N_7174,N_6077);
or U9842 (N_9842,N_6881,N_5562);
nor U9843 (N_9843,N_7359,N_6324);
and U9844 (N_9844,N_6729,N_5963);
nand U9845 (N_9845,N_6794,N_6194);
nand U9846 (N_9846,N_5039,N_5151);
nand U9847 (N_9847,N_7103,N_7047);
or U9848 (N_9848,N_5338,N_6624);
or U9849 (N_9849,N_5626,N_7400);
or U9850 (N_9850,N_5966,N_6241);
nand U9851 (N_9851,N_6700,N_7073);
nand U9852 (N_9852,N_6812,N_6847);
nor U9853 (N_9853,N_6052,N_6652);
nor U9854 (N_9854,N_6149,N_5432);
and U9855 (N_9855,N_5507,N_5984);
and U9856 (N_9856,N_5686,N_5602);
nor U9857 (N_9857,N_7033,N_5608);
or U9858 (N_9858,N_6825,N_7423);
nand U9859 (N_9859,N_6017,N_5845);
and U9860 (N_9860,N_6738,N_6702);
nor U9861 (N_9861,N_5802,N_6392);
and U9862 (N_9862,N_5085,N_5035);
nor U9863 (N_9863,N_5175,N_5193);
nand U9864 (N_9864,N_7412,N_6427);
or U9865 (N_9865,N_7494,N_5436);
and U9866 (N_9866,N_7004,N_5045);
nand U9867 (N_9867,N_7454,N_7085);
nor U9868 (N_9868,N_6280,N_5738);
nor U9869 (N_9869,N_5481,N_7016);
and U9870 (N_9870,N_5705,N_6460);
and U9871 (N_9871,N_7116,N_6975);
nand U9872 (N_9872,N_6558,N_5359);
nor U9873 (N_9873,N_5751,N_7208);
and U9874 (N_9874,N_5191,N_6461);
and U9875 (N_9875,N_6301,N_7484);
nor U9876 (N_9876,N_6137,N_6292);
or U9877 (N_9877,N_6977,N_6228);
nand U9878 (N_9878,N_5159,N_6130);
nand U9879 (N_9879,N_7219,N_5523);
or U9880 (N_9880,N_6909,N_5562);
nand U9881 (N_9881,N_5205,N_6621);
nor U9882 (N_9882,N_7148,N_5571);
nand U9883 (N_9883,N_6990,N_6364);
and U9884 (N_9884,N_6410,N_7476);
or U9885 (N_9885,N_5390,N_5829);
or U9886 (N_9886,N_7350,N_5904);
nor U9887 (N_9887,N_6645,N_6116);
and U9888 (N_9888,N_6242,N_7310);
nand U9889 (N_9889,N_6879,N_6888);
nand U9890 (N_9890,N_5271,N_7363);
or U9891 (N_9891,N_6555,N_6199);
nand U9892 (N_9892,N_6796,N_5556);
or U9893 (N_9893,N_7357,N_7204);
and U9894 (N_9894,N_5793,N_6619);
and U9895 (N_9895,N_7296,N_5306);
nor U9896 (N_9896,N_6401,N_6746);
and U9897 (N_9897,N_6347,N_5687);
or U9898 (N_9898,N_5079,N_5497);
or U9899 (N_9899,N_7376,N_6972);
and U9900 (N_9900,N_5154,N_5757);
or U9901 (N_9901,N_6046,N_5332);
nand U9902 (N_9902,N_5832,N_5839);
nor U9903 (N_9903,N_5897,N_5907);
or U9904 (N_9904,N_5905,N_5929);
or U9905 (N_9905,N_7430,N_5123);
or U9906 (N_9906,N_7049,N_7412);
and U9907 (N_9907,N_5689,N_5124);
nor U9908 (N_9908,N_6780,N_5253);
and U9909 (N_9909,N_6730,N_5003);
or U9910 (N_9910,N_5743,N_5713);
and U9911 (N_9911,N_6441,N_5345);
xnor U9912 (N_9912,N_6386,N_6846);
or U9913 (N_9913,N_6687,N_6636);
or U9914 (N_9914,N_7434,N_6248);
and U9915 (N_9915,N_7012,N_5108);
nor U9916 (N_9916,N_7365,N_5701);
xnor U9917 (N_9917,N_6412,N_6883);
nand U9918 (N_9918,N_5660,N_7230);
and U9919 (N_9919,N_5453,N_6579);
and U9920 (N_9920,N_5282,N_5768);
and U9921 (N_9921,N_5508,N_7177);
nor U9922 (N_9922,N_6557,N_5046);
and U9923 (N_9923,N_5820,N_5617);
nand U9924 (N_9924,N_6886,N_6910);
and U9925 (N_9925,N_5677,N_5532);
nand U9926 (N_9926,N_7458,N_5924);
xor U9927 (N_9927,N_5592,N_5573);
nand U9928 (N_9928,N_5985,N_7307);
nor U9929 (N_9929,N_6158,N_5515);
and U9930 (N_9930,N_5684,N_5593);
and U9931 (N_9931,N_6713,N_7211);
and U9932 (N_9932,N_5584,N_6788);
or U9933 (N_9933,N_5334,N_5309);
and U9934 (N_9934,N_6326,N_6853);
and U9935 (N_9935,N_7056,N_5040);
nor U9936 (N_9936,N_5385,N_6626);
or U9937 (N_9937,N_6020,N_6487);
nor U9938 (N_9938,N_5401,N_5791);
nor U9939 (N_9939,N_7021,N_6617);
nand U9940 (N_9940,N_6591,N_5374);
or U9941 (N_9941,N_5838,N_6410);
or U9942 (N_9942,N_6880,N_7219);
or U9943 (N_9943,N_6850,N_5123);
xnor U9944 (N_9944,N_5553,N_6915);
or U9945 (N_9945,N_6925,N_5059);
and U9946 (N_9946,N_7491,N_5189);
or U9947 (N_9947,N_5722,N_5379);
and U9948 (N_9948,N_6228,N_7194);
nor U9949 (N_9949,N_7255,N_5164);
nand U9950 (N_9950,N_5305,N_5404);
nand U9951 (N_9951,N_6665,N_6643);
and U9952 (N_9952,N_5146,N_7352);
nand U9953 (N_9953,N_5742,N_5671);
and U9954 (N_9954,N_6591,N_6958);
nor U9955 (N_9955,N_6870,N_7493);
and U9956 (N_9956,N_6808,N_6602);
nand U9957 (N_9957,N_6849,N_5336);
nand U9958 (N_9958,N_5474,N_6054);
nor U9959 (N_9959,N_6600,N_5464);
and U9960 (N_9960,N_6569,N_7163);
nor U9961 (N_9961,N_7227,N_7090);
nor U9962 (N_9962,N_7086,N_6460);
nand U9963 (N_9963,N_6149,N_5251);
or U9964 (N_9964,N_7245,N_6287);
nor U9965 (N_9965,N_5704,N_5106);
nand U9966 (N_9966,N_5730,N_5273);
nand U9967 (N_9967,N_5535,N_6856);
nor U9968 (N_9968,N_6692,N_5136);
or U9969 (N_9969,N_7435,N_5196);
and U9970 (N_9970,N_6718,N_7028);
and U9971 (N_9971,N_5216,N_6988);
and U9972 (N_9972,N_7422,N_5603);
nor U9973 (N_9973,N_5785,N_6899);
and U9974 (N_9974,N_6768,N_7224);
or U9975 (N_9975,N_7496,N_6076);
or U9976 (N_9976,N_7056,N_5854);
and U9977 (N_9977,N_6914,N_6869);
or U9978 (N_9978,N_6640,N_7356);
nand U9979 (N_9979,N_5186,N_6998);
nand U9980 (N_9980,N_6511,N_5054);
and U9981 (N_9981,N_5337,N_5084);
or U9982 (N_9982,N_6868,N_5898);
or U9983 (N_9983,N_5444,N_5587);
or U9984 (N_9984,N_5798,N_5597);
and U9985 (N_9985,N_5205,N_6350);
and U9986 (N_9986,N_6123,N_7363);
or U9987 (N_9987,N_5478,N_5186);
or U9988 (N_9988,N_6673,N_6358);
and U9989 (N_9989,N_5286,N_5197);
or U9990 (N_9990,N_5821,N_7063);
or U9991 (N_9991,N_6567,N_6224);
and U9992 (N_9992,N_5625,N_5773);
and U9993 (N_9993,N_5908,N_6149);
and U9994 (N_9994,N_6638,N_6865);
and U9995 (N_9995,N_6537,N_5507);
and U9996 (N_9996,N_6385,N_7146);
nand U9997 (N_9997,N_7367,N_6232);
or U9998 (N_9998,N_5377,N_6160);
nand U9999 (N_9999,N_5068,N_7461);
or UO_0 (O_0,N_7819,N_8485);
or UO_1 (O_1,N_8194,N_9160);
nor UO_2 (O_2,N_9432,N_7691);
or UO_3 (O_3,N_8325,N_9631);
nor UO_4 (O_4,N_7545,N_9413);
nand UO_5 (O_5,N_8370,N_8079);
nand UO_6 (O_6,N_9902,N_8430);
or UO_7 (O_7,N_8642,N_9658);
nor UO_8 (O_8,N_8948,N_8831);
nand UO_9 (O_9,N_9868,N_8421);
nor UO_10 (O_10,N_9044,N_8221);
or UO_11 (O_11,N_9789,N_7523);
and UO_12 (O_12,N_9155,N_7723);
nand UO_13 (O_13,N_8352,N_9786);
nand UO_14 (O_14,N_7813,N_9128);
or UO_15 (O_15,N_7538,N_9465);
nand UO_16 (O_16,N_7969,N_9643);
or UO_17 (O_17,N_9877,N_8181);
and UO_18 (O_18,N_9866,N_7880);
nand UO_19 (O_19,N_8660,N_8117);
nand UO_20 (O_20,N_9088,N_9520);
and UO_21 (O_21,N_7769,N_9619);
nand UO_22 (O_22,N_8164,N_8254);
and UO_23 (O_23,N_9648,N_7816);
and UO_24 (O_24,N_7830,N_8617);
nand UO_25 (O_25,N_7541,N_8032);
and UO_26 (O_26,N_8801,N_9672);
and UO_27 (O_27,N_8231,N_8108);
or UO_28 (O_28,N_9348,N_8057);
nand UO_29 (O_29,N_9264,N_9890);
nand UO_30 (O_30,N_7787,N_8677);
nand UO_31 (O_31,N_9669,N_7853);
or UO_32 (O_32,N_7936,N_8578);
nor UO_33 (O_33,N_7825,N_8227);
nand UO_34 (O_34,N_9375,N_8806);
and UO_35 (O_35,N_8982,N_7697);
nor UO_36 (O_36,N_8062,N_7924);
nor UO_37 (O_37,N_9070,N_7945);
nor UO_38 (O_38,N_8455,N_8726);
nand UO_39 (O_39,N_8196,N_8749);
or UO_40 (O_40,N_8741,N_8453);
nand UO_41 (O_41,N_9320,N_9365);
or UO_42 (O_42,N_8997,N_9286);
or UO_43 (O_43,N_9930,N_7535);
nand UO_44 (O_44,N_8050,N_9045);
nand UO_45 (O_45,N_9460,N_8454);
nand UO_46 (O_46,N_8715,N_9259);
nand UO_47 (O_47,N_8613,N_8844);
or UO_48 (O_48,N_8667,N_9006);
nor UO_49 (O_49,N_9040,N_8569);
nand UO_50 (O_50,N_8423,N_8022);
nand UO_51 (O_51,N_8949,N_8674);
nor UO_52 (O_52,N_8193,N_9493);
or UO_53 (O_53,N_7875,N_9411);
nor UO_54 (O_54,N_8826,N_7955);
and UO_55 (O_55,N_9826,N_9331);
and UO_56 (O_56,N_8870,N_8582);
or UO_57 (O_57,N_7514,N_9201);
or UO_58 (O_58,N_8590,N_8414);
nor UO_59 (O_59,N_9932,N_8863);
nor UO_60 (O_60,N_8415,N_8571);
nor UO_61 (O_61,N_8290,N_9087);
nor UO_62 (O_62,N_8872,N_9464);
and UO_63 (O_63,N_9858,N_8123);
xnor UO_64 (O_64,N_8085,N_9157);
and UO_65 (O_65,N_7999,N_9479);
nor UO_66 (O_66,N_8347,N_9692);
nor UO_67 (O_67,N_9033,N_9633);
nor UO_68 (O_68,N_8804,N_7504);
nand UO_69 (O_69,N_9846,N_8572);
nand UO_70 (O_70,N_9838,N_8541);
and UO_71 (O_71,N_8614,N_8862);
nor UO_72 (O_72,N_8697,N_8066);
nand UO_73 (O_73,N_9506,N_8373);
or UO_74 (O_74,N_9947,N_8452);
and UO_75 (O_75,N_7755,N_7569);
or UO_76 (O_76,N_8632,N_9207);
and UO_77 (O_77,N_8914,N_9165);
nand UO_78 (O_78,N_7991,N_7786);
nand UO_79 (O_79,N_7752,N_9483);
or UO_80 (O_80,N_9812,N_9974);
nor UO_81 (O_81,N_9314,N_8795);
nor UO_82 (O_82,N_8515,N_7624);
nor UO_83 (O_83,N_9120,N_9530);
or UO_84 (O_84,N_8887,N_8473);
and UO_85 (O_85,N_9030,N_9263);
and UO_86 (O_86,N_8670,N_9385);
and UO_87 (O_87,N_8885,N_8597);
or UO_88 (O_88,N_9579,N_9950);
xnor UO_89 (O_89,N_8889,N_8036);
and UO_90 (O_90,N_8437,N_7989);
and UO_91 (O_91,N_9687,N_9351);
or UO_92 (O_92,N_8777,N_8069);
and UO_93 (O_93,N_9934,N_8750);
and UO_94 (O_94,N_7930,N_8358);
nor UO_95 (O_95,N_9086,N_7548);
and UO_96 (O_96,N_8052,N_9970);
and UO_97 (O_97,N_7728,N_9377);
xor UO_98 (O_98,N_9136,N_9624);
nand UO_99 (O_99,N_9000,N_9834);
nor UO_100 (O_100,N_7790,N_8934);
nor UO_101 (O_101,N_9783,N_8110);
and UO_102 (O_102,N_8764,N_8360);
nand UO_103 (O_103,N_9913,N_9545);
nand UO_104 (O_104,N_9062,N_7658);
nor UO_105 (O_105,N_9374,N_8019);
nor UO_106 (O_106,N_8843,N_8270);
or UO_107 (O_107,N_7996,N_8903);
or UO_108 (O_108,N_9294,N_9336);
and UO_109 (O_109,N_7820,N_8609);
or UO_110 (O_110,N_9611,N_8368);
and UO_111 (O_111,N_7729,N_9049);
nand UO_112 (O_112,N_7946,N_8317);
nor UO_113 (O_113,N_8546,N_9043);
nand UO_114 (O_114,N_8707,N_8045);
and UO_115 (O_115,N_8217,N_8957);
or UO_116 (O_116,N_9205,N_8692);
and UO_117 (O_117,N_9435,N_8943);
or UO_118 (O_118,N_8257,N_9972);
nand UO_119 (O_119,N_9569,N_9050);
nor UO_120 (O_120,N_9880,N_9808);
xnor UO_121 (O_121,N_9038,N_9510);
or UO_122 (O_122,N_9738,N_8976);
and UO_123 (O_123,N_8895,N_9342);
and UO_124 (O_124,N_8098,N_9983);
nand UO_125 (O_125,N_8868,N_9380);
and UO_126 (O_126,N_8116,N_8979);
and UO_127 (O_127,N_9814,N_7603);
and UO_128 (O_128,N_7881,N_8179);
or UO_129 (O_129,N_9488,N_8854);
nand UO_130 (O_130,N_9558,N_8511);
or UO_131 (O_131,N_8133,N_8324);
or UO_132 (O_132,N_8721,N_7685);
nor UO_133 (O_133,N_9985,N_7968);
nand UO_134 (O_134,N_7859,N_9001);
or UO_135 (O_135,N_9756,N_8995);
or UO_136 (O_136,N_8812,N_8488);
or UO_137 (O_137,N_7808,N_8713);
nand UO_138 (O_138,N_9248,N_9338);
nor UO_139 (O_139,N_9570,N_9098);
nor UO_140 (O_140,N_9878,N_9412);
nor UO_141 (O_141,N_9709,N_7829);
nand UO_142 (O_142,N_9544,N_8813);
and UO_143 (O_143,N_9119,N_7674);
nor UO_144 (O_144,N_8586,N_8683);
nand UO_145 (O_145,N_8433,N_8260);
and UO_146 (O_146,N_8694,N_9613);
xnor UO_147 (O_147,N_9847,N_8836);
nand UO_148 (O_148,N_7975,N_8404);
or UO_149 (O_149,N_8576,N_9238);
nand UO_150 (O_150,N_8180,N_8418);
nor UO_151 (O_151,N_7725,N_9993);
nand UO_152 (O_152,N_7988,N_7689);
and UO_153 (O_153,N_9919,N_9796);
nor UO_154 (O_154,N_8672,N_8252);
nand UO_155 (O_155,N_9154,N_8969);
or UO_156 (O_156,N_8131,N_7977);
or UO_157 (O_157,N_9899,N_9221);
nor UO_158 (O_158,N_9256,N_7583);
and UO_159 (O_159,N_7534,N_9300);
or UO_160 (O_160,N_9478,N_9508);
and UO_161 (O_161,N_9711,N_7531);
or UO_162 (O_162,N_8309,N_9801);
and UO_163 (O_163,N_9287,N_9757);
nand UO_164 (O_164,N_7644,N_9935);
or UO_165 (O_165,N_7501,N_9228);
nand UO_166 (O_166,N_7507,N_8966);
or UO_167 (O_167,N_9410,N_7692);
nand UO_168 (O_168,N_8524,N_8395);
xnor UO_169 (O_169,N_7978,N_8145);
nand UO_170 (O_170,N_9112,N_9021);
nor UO_171 (O_171,N_7597,N_7879);
nand UO_172 (O_172,N_7715,N_9937);
or UO_173 (O_173,N_8607,N_9129);
nand UO_174 (O_174,N_8731,N_8356);
or UO_175 (O_175,N_7872,N_8086);
or UO_176 (O_176,N_7759,N_8757);
or UO_177 (O_177,N_7855,N_9197);
nor UO_178 (O_178,N_8702,N_9936);
nand UO_179 (O_179,N_9321,N_8323);
or UO_180 (O_180,N_8769,N_9524);
and UO_181 (O_181,N_7575,N_9952);
and UO_182 (O_182,N_7857,N_7610);
nor UO_183 (O_183,N_8880,N_8555);
nand UO_184 (O_184,N_8517,N_7647);
nor UO_185 (O_185,N_9209,N_8971);
nor UO_186 (O_186,N_7884,N_8648);
or UO_187 (O_187,N_8417,N_8581);
and UO_188 (O_188,N_9730,N_8779);
xnor UO_189 (O_189,N_7783,N_9311);
and UO_190 (O_190,N_8074,N_9056);
nor UO_191 (O_191,N_8160,N_9768);
or UO_192 (O_192,N_9054,N_7951);
or UO_193 (O_193,N_9004,N_9131);
or UO_194 (O_194,N_9518,N_9519);
or UO_195 (O_195,N_7745,N_7921);
nand UO_196 (O_196,N_7985,N_8816);
or UO_197 (O_197,N_9873,N_9299);
nand UO_198 (O_198,N_7874,N_7997);
xnor UO_199 (O_199,N_9270,N_9064);
and UO_200 (O_200,N_8424,N_8551);
nor UO_201 (O_201,N_8681,N_8600);
nor UO_202 (O_202,N_7672,N_8624);
nand UO_203 (O_203,N_8302,N_7664);
nor UO_204 (O_204,N_9130,N_7887);
nand UO_205 (O_205,N_8554,N_8748);
nor UO_206 (O_206,N_7681,N_8402);
nand UO_207 (O_207,N_8809,N_9760);
or UO_208 (O_208,N_7742,N_8587);
and UO_209 (O_209,N_8640,N_9785);
and UO_210 (O_210,N_8346,N_9398);
and UO_211 (O_211,N_8782,N_9068);
nor UO_212 (O_212,N_8530,N_8026);
nand UO_213 (O_213,N_7846,N_9978);
or UO_214 (O_214,N_8175,N_7952);
nor UO_215 (O_215,N_8172,N_9969);
and UO_216 (O_216,N_9470,N_8465);
nor UO_217 (O_217,N_9451,N_8710);
or UO_218 (O_218,N_8321,N_7770);
nor UO_219 (O_219,N_8449,N_7935);
and UO_220 (O_220,N_9604,N_8706);
and UO_221 (O_221,N_9487,N_9720);
nor UO_222 (O_222,N_9632,N_8818);
and UO_223 (O_223,N_7626,N_7910);
and UO_224 (O_224,N_8030,N_9162);
and UO_225 (O_225,N_7730,N_8040);
and UO_226 (O_226,N_9861,N_8932);
nor UO_227 (O_227,N_8186,N_9616);
and UO_228 (O_228,N_9822,N_9026);
and UO_229 (O_229,N_8407,N_9526);
nand UO_230 (O_230,N_9523,N_9968);
and UO_231 (O_231,N_9617,N_7915);
nand UO_232 (O_232,N_8192,N_8357);
and UO_233 (O_233,N_9436,N_7556);
or UO_234 (O_234,N_8082,N_9215);
nand UO_235 (O_235,N_8759,N_8850);
nor UO_236 (O_236,N_7718,N_8907);
and UO_237 (O_237,N_9053,N_8199);
nor UO_238 (O_238,N_9258,N_9325);
nor UO_239 (O_239,N_8183,N_8120);
nand UO_240 (O_240,N_8564,N_7596);
or UO_241 (O_241,N_7803,N_9614);
nand UO_242 (O_242,N_7850,N_9159);
and UO_243 (O_243,N_9859,N_8182);
or UO_244 (O_244,N_8408,N_9521);
or UO_245 (O_245,N_8558,N_9654);
or UO_246 (O_246,N_9670,N_7851);
or UO_247 (O_247,N_9942,N_8959);
nor UO_248 (O_248,N_8878,N_8915);
nand UO_249 (O_249,N_8393,N_8457);
nor UO_250 (O_250,N_7743,N_8251);
nor UO_251 (O_251,N_7923,N_8771);
xnor UO_252 (O_252,N_9513,N_8389);
nor UO_253 (O_253,N_9603,N_9772);
or UO_254 (O_254,N_7572,N_9090);
nand UO_255 (O_255,N_8262,N_8647);
nand UO_256 (O_256,N_7706,N_9010);
or UO_257 (O_257,N_9995,N_9875);
nor UO_258 (O_258,N_9565,N_8923);
or UO_259 (O_259,N_9057,N_8662);
nor UO_260 (O_260,N_8048,N_9369);
and UO_261 (O_261,N_8591,N_8666);
nand UO_262 (O_262,N_8925,N_8023);
nand UO_263 (O_263,N_7947,N_9431);
nand UO_264 (O_264,N_8964,N_8154);
nor UO_265 (O_265,N_9386,N_8051);
nand UO_266 (O_266,N_8920,N_8851);
nand UO_267 (O_267,N_7929,N_8960);
and UO_268 (O_268,N_7707,N_8785);
or UO_269 (O_269,N_7578,N_7905);
nor UO_270 (O_270,N_8810,N_8875);
and UO_271 (O_271,N_9237,N_9954);
and UO_272 (O_272,N_9231,N_7521);
nand UO_273 (O_273,N_8138,N_9511);
xor UO_274 (O_274,N_7721,N_9115);
or UO_275 (O_275,N_9929,N_8886);
nor UO_276 (O_276,N_8191,N_8800);
and UO_277 (O_277,N_9378,N_8746);
nor UO_278 (O_278,N_9623,N_8912);
nor UO_279 (O_279,N_7934,N_9168);
nor UO_280 (O_280,N_7637,N_9002);
nor UO_281 (O_281,N_9703,N_7640);
and UO_282 (O_282,N_9025,N_9618);
nor UO_283 (O_283,N_9099,N_7630);
nand UO_284 (O_284,N_7709,N_8918);
or UO_285 (O_285,N_8080,N_8874);
xor UO_286 (O_286,N_9288,N_7954);
nor UO_287 (O_287,N_8328,N_8763);
nor UO_288 (O_288,N_8282,N_9546);
nand UO_289 (O_289,N_9684,N_8815);
nor UO_290 (O_290,N_7878,N_7958);
or UO_291 (O_291,N_9484,N_7869);
or UO_292 (O_292,N_8207,N_8823);
or UO_293 (O_293,N_8313,N_9555);
nand UO_294 (O_294,N_7520,N_8780);
or UO_295 (O_295,N_8204,N_8708);
and UO_296 (O_296,N_9951,N_7741);
or UO_297 (O_297,N_9870,N_8367);
nor UO_298 (O_298,N_9240,N_7877);
nor UO_299 (O_299,N_8226,N_9172);
nand UO_300 (O_300,N_8723,N_8655);
nor UO_301 (O_301,N_9246,N_7839);
or UO_302 (O_302,N_9754,N_9339);
and UO_303 (O_303,N_8441,N_9071);
nor UO_304 (O_304,N_9980,N_8615);
nand UO_305 (O_305,N_9590,N_8950);
and UO_306 (O_306,N_7772,N_7841);
xor UO_307 (O_307,N_8503,N_8029);
and UO_308 (O_308,N_8289,N_8848);
nor UO_309 (O_309,N_9674,N_9559);
nand UO_310 (O_310,N_7619,N_8805);
and UO_311 (O_311,N_9492,N_9194);
nand UO_312 (O_312,N_8714,N_9975);
and UO_313 (O_313,N_9864,N_9457);
or UO_314 (O_314,N_9886,N_9047);
nor UO_315 (O_315,N_8059,N_8392);
or UO_316 (O_316,N_9609,N_7993);
nor UO_317 (O_317,N_9244,N_9897);
nor UO_318 (O_318,N_9312,N_9364);
or UO_319 (O_319,N_8263,N_7594);
or UO_320 (O_320,N_9399,N_7810);
or UO_321 (O_321,N_9835,N_7529);
and UO_322 (O_322,N_8743,N_9229);
nand UO_323 (O_323,N_8869,N_9769);
or UO_324 (O_324,N_8083,N_9179);
or UO_325 (O_325,N_8673,N_8386);
or UO_326 (O_326,N_9036,N_8579);
or UO_327 (O_327,N_8039,N_7606);
or UO_328 (O_328,N_9214,N_8988);
nand UO_329 (O_329,N_9096,N_9145);
xnor UO_330 (O_330,N_8222,N_8775);
nor UO_331 (O_331,N_8320,N_8447);
nor UO_332 (O_332,N_9607,N_8709);
nor UO_333 (O_333,N_9359,N_7982);
nand UO_334 (O_334,N_9466,N_8140);
nor UO_335 (O_335,N_9807,N_8876);
and UO_336 (O_336,N_8636,N_8926);
or UO_337 (O_337,N_9103,N_9236);
or UO_338 (O_338,N_9184,N_8371);
nor UO_339 (O_339,N_8213,N_8130);
or UO_340 (O_340,N_9111,N_8865);
or UO_341 (O_341,N_9798,N_9360);
nor UO_342 (O_342,N_9200,N_9502);
and UO_343 (O_343,N_9997,N_9211);
and UO_344 (O_344,N_9576,N_8456);
xnor UO_345 (O_345,N_8046,N_8671);
nor UO_346 (O_346,N_9713,N_9035);
or UO_347 (O_347,N_7774,N_7590);
or UO_348 (O_348,N_9437,N_9029);
nand UO_349 (O_349,N_8261,N_7611);
nor UO_350 (O_350,N_9811,N_9490);
nand UO_351 (O_351,N_7657,N_9525);
nand UO_352 (O_352,N_9243,N_9516);
and UO_353 (O_353,N_8475,N_9509);
nand UO_354 (O_354,N_7913,N_8291);
nand UO_355 (O_355,N_9589,N_9725);
and UO_356 (O_356,N_8119,N_9093);
nor UO_357 (O_357,N_9368,N_8300);
nor UO_358 (O_358,N_7828,N_8978);
and UO_359 (O_359,N_9220,N_8814);
nand UO_360 (O_360,N_9110,N_9885);
nand UO_361 (O_361,N_8333,N_9612);
nor UO_362 (O_362,N_9192,N_8519);
nand UO_363 (O_363,N_8202,N_9727);
nand UO_364 (O_364,N_9731,N_8256);
nor UO_365 (O_365,N_8722,N_9046);
or UO_366 (O_366,N_8442,N_8150);
or UO_367 (O_367,N_7612,N_9426);
or UO_368 (O_368,N_8124,N_9856);
nor UO_369 (O_369,N_7525,N_9055);
and UO_370 (O_370,N_7896,N_8195);
and UO_371 (O_371,N_9819,N_9733);
nor UO_372 (O_372,N_9548,N_7659);
and UO_373 (O_373,N_9923,N_9039);
nor UO_374 (O_374,N_7831,N_9247);
or UO_375 (O_375,N_9156,N_8450);
or UO_376 (O_376,N_9373,N_8244);
and UO_377 (O_377,N_9202,N_9125);
and UO_378 (O_378,N_9127,N_8625);
nand UO_379 (O_379,N_7651,N_7891);
and UO_380 (O_380,N_8893,N_8266);
xor UO_381 (O_381,N_8595,N_9764);
nand UO_382 (O_382,N_8902,N_8857);
nand UO_383 (O_383,N_7648,N_8536);
nand UO_384 (O_384,N_9906,N_9716);
nor UO_385 (O_385,N_7898,N_8072);
nand UO_386 (O_386,N_7971,N_8305);
nor UO_387 (O_387,N_8345,N_8992);
or UO_388 (O_388,N_7967,N_7508);
and UO_389 (O_389,N_8007,N_7843);
nor UO_390 (O_390,N_9638,N_9498);
nand UO_391 (O_391,N_9366,N_7581);
or UO_392 (O_392,N_7615,N_7515);
nand UO_393 (O_393,N_8834,N_8277);
nand UO_394 (O_394,N_7516,N_7738);
nand UO_395 (O_395,N_9898,N_8087);
nor UO_396 (O_396,N_8380,N_8152);
and UO_397 (O_397,N_9770,N_8512);
or UO_398 (O_398,N_9085,N_9344);
and UO_399 (O_399,N_8500,N_9960);
and UO_400 (O_400,N_7938,N_9126);
nand UO_401 (O_401,N_9271,N_9080);
nor UO_402 (O_402,N_8197,N_7795);
nand UO_403 (O_403,N_8544,N_9135);
nand UO_404 (O_404,N_9109,N_8972);
nor UO_405 (O_405,N_9013,N_8278);
nand UO_406 (O_406,N_9408,N_8526);
and UO_407 (O_407,N_8330,N_7974);
nand UO_408 (O_408,N_9625,N_8126);
or UO_409 (O_409,N_9134,N_9661);
and UO_410 (O_410,N_7732,N_9343);
or UO_411 (O_411,N_9362,N_7713);
or UO_412 (O_412,N_8911,N_9644);
or UO_413 (O_413,N_9938,N_9704);
and UO_414 (O_414,N_9356,N_7694);
xnor UO_415 (O_415,N_7608,N_7894);
and UO_416 (O_416,N_9636,N_8973);
or UO_417 (O_417,N_9973,N_8701);
nand UO_418 (O_418,N_7511,N_7798);
nor UO_419 (O_419,N_8020,N_9328);
nand UO_420 (O_420,N_7727,N_8686);
nand UO_421 (O_421,N_9139,N_8255);
nor UO_422 (O_422,N_8489,N_9438);
and UO_423 (O_423,N_8996,N_8467);
and UO_424 (O_424,N_9940,N_9924);
and UO_425 (O_425,N_7646,N_7797);
nor UO_426 (O_426,N_9788,N_8822);
xnor UO_427 (O_427,N_8965,N_9441);
or UO_428 (O_428,N_9901,N_8416);
nand UO_429 (O_429,N_7739,N_8700);
xor UO_430 (O_430,N_8766,N_8487);
nor UO_431 (O_431,N_9887,N_9204);
nor UO_432 (O_432,N_8419,N_8004);
nor UO_433 (O_433,N_9140,N_9007);
or UO_434 (O_434,N_9468,N_9815);
or UO_435 (O_435,N_9635,N_9371);
nand UO_436 (O_436,N_9630,N_8657);
nand UO_437 (O_437,N_9586,N_9537);
or UO_438 (O_438,N_9434,N_9967);
or UO_439 (O_439,N_8369,N_8012);
and UO_440 (O_440,N_9739,N_9305);
nor UO_441 (O_441,N_8101,N_7773);
or UO_442 (O_442,N_9800,N_8398);
nor UO_443 (O_443,N_9882,N_8977);
nor UO_444 (O_444,N_7925,N_9606);
and UO_445 (O_445,N_9051,N_9909);
and UO_446 (O_446,N_9844,N_8315);
nor UO_447 (O_447,N_8730,N_8054);
and UO_448 (O_448,N_9963,N_8651);
nand UO_449 (O_449,N_9186,N_8990);
nand UO_450 (O_450,N_9400,N_9907);
nor UO_451 (O_451,N_7963,N_7605);
or UO_452 (O_452,N_8445,N_9459);
nand UO_453 (O_453,N_9118,N_7660);
and UO_454 (O_454,N_7775,N_7570);
or UO_455 (O_455,N_7650,N_7909);
nor UO_456 (O_456,N_8668,N_9554);
nand UO_457 (O_457,N_7505,N_7865);
nor UO_458 (O_458,N_9745,N_9384);
nand UO_459 (O_459,N_8148,N_7542);
and UO_460 (O_460,N_9595,N_7994);
and UO_461 (O_461,N_7785,N_7622);
nand UO_462 (O_462,N_7842,N_7832);
and UO_463 (O_463,N_7631,N_7544);
nor UO_464 (O_464,N_9095,N_8570);
or UO_465 (O_465,N_8618,N_7838);
or UO_466 (O_466,N_8596,N_8219);
nor UO_467 (O_467,N_8711,N_7740);
nand UO_468 (O_468,N_9335,N_9620);
and UO_469 (O_469,N_9310,N_8236);
nor UO_470 (O_470,N_9597,N_8877);
nand UO_471 (O_471,N_8155,N_8983);
nand UO_472 (O_472,N_9181,N_9376);
nor UO_473 (O_473,N_9405,N_9023);
nand UO_474 (O_474,N_8669,N_7809);
or UO_475 (O_475,N_9361,N_7557);
nor UO_476 (O_476,N_7995,N_7661);
and UO_477 (O_477,N_8623,N_7771);
or UO_478 (O_478,N_9073,N_9628);
or UO_479 (O_479,N_8696,N_8353);
nand UO_480 (O_480,N_7766,N_9257);
nor UO_481 (O_481,N_9908,N_9164);
and UO_482 (O_482,N_9539,N_9991);
xnor UO_483 (O_483,N_9241,N_7502);
xnor UO_484 (O_484,N_9306,N_8755);
nand UO_485 (O_485,N_7673,N_7565);
nand UO_486 (O_486,N_8825,N_7509);
nand UO_487 (O_487,N_9170,N_7553);
nor UO_488 (O_488,N_8127,N_7807);
nand UO_489 (O_489,N_9825,N_8930);
or UO_490 (O_490,N_9301,N_8088);
and UO_491 (O_491,N_8507,N_9933);
nand UO_492 (O_492,N_8724,N_9146);
or UO_493 (O_493,N_9206,N_8017);
nand UO_494 (O_494,N_8234,N_7871);
nor UO_495 (O_495,N_7966,N_8153);
or UO_496 (O_496,N_8298,N_7562);
nor UO_497 (O_497,N_8936,N_8738);
nor UO_498 (O_498,N_8728,N_7802);
or UO_499 (O_499,N_9028,N_7675);
or UO_500 (O_500,N_9094,N_9699);
nand UO_501 (O_501,N_9250,N_9958);
nor UO_502 (O_502,N_9133,N_9702);
and UO_503 (O_503,N_9792,N_8604);
nand UO_504 (O_504,N_8499,N_8177);
or UO_505 (O_505,N_9462,N_8159);
or UO_506 (O_506,N_9210,N_8562);
or UO_507 (O_507,N_8841,N_9227);
and UO_508 (O_508,N_8856,N_9317);
and UO_509 (O_509,N_9686,N_9673);
or UO_510 (O_510,N_9076,N_7788);
or UO_511 (O_511,N_8549,N_8840);
nand UO_512 (O_512,N_7901,N_9793);
nand UO_513 (O_513,N_9842,N_9016);
nor UO_514 (O_514,N_9500,N_8747);
nand UO_515 (O_515,N_8426,N_9254);
nor UO_516 (O_516,N_9132,N_9665);
or UO_517 (O_517,N_8652,N_8808);
or UO_518 (O_518,N_9262,N_7762);
or UO_519 (O_519,N_9860,N_9218);
or UO_520 (O_520,N_8735,N_9728);
nor UO_521 (O_521,N_8705,N_8884);
nor UO_522 (O_522,N_8993,N_8171);
and UO_523 (O_523,N_9041,N_7749);
and UO_524 (O_524,N_9863,N_8946);
nand UO_525 (O_525,N_9444,N_7784);
nand UO_526 (O_526,N_7931,N_9276);
nand UO_527 (O_527,N_8751,N_8073);
nand UO_528 (O_528,N_9867,N_9697);
nor UO_529 (O_529,N_8961,N_9448);
and UO_530 (O_530,N_8921,N_8846);
or UO_531 (O_531,N_9552,N_8928);
nor UO_532 (O_532,N_9037,N_8077);
and UO_533 (O_533,N_9323,N_8508);
or UO_534 (O_534,N_7503,N_8361);
or UO_535 (O_535,N_8799,N_9627);
nor UO_536 (O_536,N_8143,N_8283);
and UO_537 (O_537,N_8390,N_9082);
or UO_538 (O_538,N_8975,N_9449);
nand UO_539 (O_539,N_8157,N_9580);
nor UO_540 (O_540,N_9979,N_8341);
nor UO_541 (O_541,N_9829,N_9587);
or UO_542 (O_542,N_9225,N_8092);
xor UO_543 (O_543,N_8537,N_8952);
or UO_544 (O_544,N_9629,N_8789);
nor UO_545 (O_545,N_8829,N_8016);
nand UO_546 (O_546,N_9163,N_8243);
and UO_547 (O_547,N_9660,N_9547);
and UO_548 (O_548,N_8327,N_8881);
nand UO_549 (O_549,N_8167,N_8067);
and UO_550 (O_550,N_8797,N_8363);
and UO_551 (O_551,N_8786,N_7777);
and UO_552 (O_552,N_7714,N_8680);
and UO_553 (O_553,N_8510,N_8435);
nand UO_554 (O_554,N_8462,N_9688);
xnor UO_555 (O_555,N_8529,N_7948);
and UO_556 (O_556,N_7889,N_9735);
or UO_557 (O_557,N_8432,N_8264);
nor UO_558 (O_558,N_7789,N_8448);
nor UO_559 (O_559,N_9759,N_9747);
or UO_560 (O_560,N_7911,N_7811);
nor UO_561 (O_561,N_8888,N_9066);
nor UO_562 (O_562,N_7903,N_8910);
nor UO_563 (O_563,N_9668,N_8477);
nand UO_564 (O_564,N_9199,N_7888);
or UO_565 (O_565,N_7680,N_7900);
and UO_566 (O_566,N_8334,N_8601);
and UO_567 (O_567,N_7890,N_9639);
nand UO_568 (O_568,N_8388,N_8314);
nor UO_569 (O_569,N_9529,N_8643);
and UO_570 (O_570,N_9151,N_7591);
nor UO_571 (O_571,N_9837,N_7733);
or UO_572 (O_572,N_9198,N_9647);
or UO_573 (O_573,N_9141,N_9795);
or UO_574 (O_574,N_9245,N_8210);
nand UO_575 (O_575,N_7964,N_7604);
nor UO_576 (O_576,N_7632,N_8917);
nor UO_577 (O_577,N_8584,N_7984);
or UO_578 (O_578,N_8994,N_8773);
and UO_579 (O_579,N_9994,N_9946);
nand UO_580 (O_580,N_9232,N_8693);
and UO_581 (O_581,N_9357,N_8233);
nor UO_582 (O_582,N_8156,N_7695);
nand UO_583 (O_583,N_7794,N_8761);
nor UO_584 (O_584,N_8890,N_9114);
nor UO_585 (O_585,N_7751,N_9077);
or UO_586 (O_586,N_7618,N_9920);
nand UO_587 (O_587,N_9396,N_8588);
nand UO_588 (O_588,N_8206,N_8550);
nand UO_589 (O_589,N_8332,N_8798);
or UO_590 (O_590,N_7633,N_9816);
nand UO_591 (O_591,N_8807,N_8650);
and UO_592 (O_592,N_8768,N_8531);
and UO_593 (O_593,N_7862,N_9032);
or UO_594 (O_594,N_7677,N_8945);
and UO_595 (O_595,N_9748,N_8349);
nand UO_596 (O_596,N_9542,N_7665);
nand UO_597 (O_597,N_9350,N_8703);
nand UO_598 (O_598,N_7750,N_8293);
nor UO_599 (O_599,N_8556,N_9273);
nand UO_600 (O_600,N_8383,N_7653);
nand UO_601 (O_601,N_7867,N_9515);
xnor UO_602 (O_602,N_7932,N_8299);
nand UO_603 (O_603,N_8901,N_7836);
or UO_604 (O_604,N_7598,N_8285);
nor UO_605 (O_605,N_9977,N_8989);
nand UO_606 (O_606,N_9100,N_9705);
and UO_607 (O_607,N_9446,N_9535);
nand UO_608 (O_608,N_8104,N_8762);
and UO_609 (O_609,N_8631,N_9471);
nand UO_610 (O_610,N_8866,N_9480);
nor UO_611 (O_611,N_9585,N_7649);
and UO_612 (O_612,N_9827,N_9501);
or UO_613 (O_613,N_8882,N_9927);
nand UO_614 (O_614,N_9767,N_9024);
nand UO_615 (O_615,N_8563,N_9905);
nand UO_616 (O_616,N_8348,N_7737);
and UO_617 (O_617,N_9575,N_9149);
and UO_618 (O_618,N_9388,N_8034);
and UO_619 (O_619,N_9761,N_8784);
or UO_620 (O_620,N_9653,N_9916);
and UO_621 (O_621,N_8420,N_9212);
nand UO_622 (O_622,N_9260,N_8144);
nand UO_623 (O_623,N_9828,N_8355);
nor UO_624 (O_624,N_7918,N_7628);
and UO_625 (O_625,N_8479,N_9831);
nand UO_626 (O_626,N_7579,N_8205);
or UO_627 (O_627,N_8224,N_9293);
nor UO_628 (O_628,N_8845,N_8329);
and UO_629 (O_629,N_7748,N_8891);
or UO_630 (O_630,N_8474,N_7536);
nand UO_631 (O_631,N_8401,N_8575);
nand UO_632 (O_632,N_8661,N_9602);
and UO_633 (O_633,N_9690,N_7614);
and UO_634 (O_634,N_7708,N_9019);
and UO_635 (O_635,N_8927,N_8365);
nand UO_636 (O_636,N_9564,N_8005);
nand UO_637 (O_637,N_9183,N_9251);
nand UO_638 (O_638,N_8174,N_9591);
and UO_639 (O_639,N_9742,N_9532);
and UO_640 (O_640,N_8543,N_7652);
or UO_641 (O_641,N_8533,N_9671);
or UO_642 (O_642,N_9261,N_8203);
or UO_643 (O_643,N_8385,N_9721);
nand UO_644 (O_644,N_9889,N_8338);
and UO_645 (O_645,N_9896,N_8476);
nor UO_646 (O_646,N_7519,N_7686);
nand UO_647 (O_647,N_8792,N_8781);
nand UO_648 (O_648,N_9349,N_8494);
nand UO_649 (O_649,N_9418,N_7655);
or UO_650 (O_650,N_8469,N_9497);
nand UO_651 (O_651,N_7584,N_9551);
nor UO_652 (O_652,N_9401,N_8359);
nor UO_653 (O_653,N_9871,N_9284);
or UO_654 (O_654,N_8468,N_8937);
or UO_655 (O_655,N_8986,N_8163);
xor UO_656 (O_656,N_8439,N_9430);
or UO_657 (O_657,N_9178,N_8904);
nand UO_658 (O_658,N_9346,N_9774);
or UO_659 (O_659,N_7796,N_8606);
and UO_660 (O_660,N_9707,N_8405);
nand UO_661 (O_661,N_9458,N_8319);
and UO_662 (O_662,N_9990,N_7960);
nor UO_663 (O_663,N_9689,N_8436);
nand UO_664 (O_664,N_9474,N_8162);
and UO_665 (O_665,N_9475,N_8791);
nor UO_666 (O_666,N_7928,N_9113);
or UO_667 (O_667,N_7601,N_9461);
or UO_668 (O_668,N_8336,N_7779);
and UO_669 (O_669,N_8232,N_7566);
and UO_670 (O_670,N_8170,N_8387);
nor UO_671 (O_671,N_8688,N_8819);
and UO_672 (O_672,N_8049,N_8568);
and UO_673 (O_673,N_8318,N_8852);
nor UO_674 (O_674,N_9781,N_8400);
nor UO_675 (O_675,N_7817,N_9961);
or UO_676 (O_676,N_8727,N_7981);
and UO_677 (O_677,N_9666,N_8342);
nor UO_678 (O_678,N_7746,N_8128);
nor UO_679 (O_679,N_9283,N_8113);
nand UO_680 (O_680,N_9315,N_9645);
and UO_681 (O_681,N_7616,N_8010);
nor UO_682 (O_682,N_8842,N_7588);
or UO_683 (O_683,N_8275,N_8835);
nor UO_684 (O_684,N_9802,N_9712);
or UO_685 (O_685,N_7679,N_8495);
or UO_686 (O_686,N_9239,N_7818);
and UO_687 (O_687,N_8107,N_9297);
or UO_688 (O_688,N_8292,N_8042);
nor UO_689 (O_689,N_8114,N_9917);
or UO_690 (O_690,N_7688,N_8391);
and UO_691 (O_691,N_9715,N_8559);
nand UO_692 (O_692,N_8486,N_7973);
or UO_693 (O_693,N_8991,N_8754);
nor UO_694 (O_694,N_7764,N_9988);
and UO_695 (O_695,N_9732,N_9662);
or UO_696 (O_696,N_9531,N_8038);
xor UO_697 (O_697,N_7722,N_9425);
nand UO_698 (O_698,N_8610,N_9018);
and UO_699 (O_699,N_8987,N_9031);
or UO_700 (O_700,N_7720,N_7950);
nor UO_701 (O_701,N_8247,N_8281);
nand UO_702 (O_702,N_8633,N_8058);
or UO_703 (O_703,N_9762,N_9295);
nor UO_704 (O_704,N_7571,N_8654);
nor UO_705 (O_705,N_9048,N_9779);
nor UO_706 (O_706,N_7654,N_9622);
nor UO_707 (O_707,N_9810,N_9402);
nand UO_708 (O_708,N_8044,N_9177);
or UO_709 (O_709,N_8793,N_8406);
nand UO_710 (O_710,N_7801,N_7866);
nand UO_711 (O_711,N_8523,N_7833);
nand UO_712 (O_712,N_8268,N_8068);
or UO_713 (O_713,N_7671,N_9152);
nand UO_714 (O_714,N_9148,N_7962);
nand UO_715 (O_715,N_9175,N_8364);
nor UO_716 (O_716,N_9698,N_9117);
nor UO_717 (O_717,N_8956,N_9588);
xor UO_718 (O_718,N_9121,N_9876);
nor UO_719 (O_719,N_9663,N_9803);
nor UO_720 (O_720,N_7847,N_7821);
nor UO_721 (O_721,N_8573,N_7780);
nand UO_722 (O_722,N_9536,N_7669);
and UO_723 (O_723,N_8734,N_8322);
or UO_724 (O_724,N_8099,N_9701);
or UO_725 (O_725,N_9065,N_7678);
nor UO_726 (O_726,N_8297,N_9921);
nor UO_727 (O_727,N_8827,N_8060);
nand UO_728 (O_728,N_8002,N_9944);
nand UO_729 (O_729,N_8699,N_9052);
or UO_730 (O_730,N_9646,N_9626);
nor UO_731 (O_731,N_8774,N_7574);
and UO_732 (O_732,N_7893,N_9749);
or UO_733 (O_733,N_9189,N_8542);
nor UO_734 (O_734,N_7667,N_8303);
nand UO_735 (O_735,N_8464,N_7563);
and UO_736 (O_736,N_9476,N_9584);
nor UO_737 (O_737,N_8312,N_8967);
or UO_738 (O_738,N_8422,N_9034);
nand UO_739 (O_739,N_7705,N_8970);
and UO_740 (O_740,N_8250,N_8944);
or UO_741 (O_741,N_8384,N_8308);
and UO_742 (O_742,N_7899,N_8644);
nand UO_743 (O_743,N_9664,N_8228);
and UO_744 (O_744,N_7953,N_9928);
or UO_745 (O_745,N_8962,N_9903);
nand UO_746 (O_746,N_9419,N_8245);
and UO_747 (O_747,N_8855,N_7805);
or UO_748 (O_748,N_9758,N_8620);
nand UO_749 (O_749,N_9428,N_9824);
or UO_750 (O_750,N_8169,N_7768);
nor UO_751 (O_751,N_9818,N_7592);
nand UO_752 (O_752,N_9423,N_8847);
nand UO_753 (O_753,N_9443,N_7927);
nor UO_754 (O_754,N_9427,N_8307);
and UO_755 (O_755,N_9285,N_8354);
or UO_756 (O_756,N_8602,N_8294);
and UO_757 (O_757,N_9850,N_9656);
and UO_758 (O_758,N_9447,N_8223);
nand UO_759 (O_759,N_9755,N_9962);
nor UO_760 (O_760,N_8557,N_9679);
or UO_761 (O_761,N_9718,N_8397);
or UO_762 (O_762,N_9302,N_9677);
nor UO_763 (O_763,N_8035,N_8892);
and UO_764 (O_764,N_9081,N_9931);
nand UO_765 (O_765,N_8919,N_8425);
nand UO_766 (O_766,N_8378,N_8853);
and UO_767 (O_767,N_8350,N_9852);
or UO_768 (O_768,N_8151,N_8492);
nor UO_769 (O_769,N_9600,N_8820);
and UO_770 (O_770,N_9574,N_8428);
nor UO_771 (O_771,N_9641,N_7559);
nor UO_772 (O_772,N_8076,N_8985);
and UO_773 (O_773,N_9797,N_9776);
and UO_774 (O_774,N_9253,N_8024);
nor UO_775 (O_775,N_9594,N_9652);
and UO_776 (O_776,N_9097,N_8259);
and UO_777 (O_777,N_8679,N_8608);
and UO_778 (O_778,N_8136,N_8665);
nand UO_779 (O_779,N_8220,N_9404);
nor UO_780 (O_780,N_7848,N_7763);
nor UO_781 (O_781,N_8941,N_8013);
nand UO_782 (O_782,N_9020,N_9442);
and UO_783 (O_783,N_8253,N_7532);
or UO_784 (O_784,N_9719,N_9481);
or UO_785 (O_785,N_8628,N_9414);
or UO_786 (O_786,N_8211,N_9463);
nand UO_787 (O_787,N_9406,N_7602);
and UO_788 (O_788,N_8121,N_8567);
xor UO_789 (O_789,N_7864,N_8411);
or UO_790 (O_790,N_8132,N_9265);
or UO_791 (O_791,N_7776,N_9538);
and UO_792 (O_792,N_9123,N_8134);
or UO_793 (O_793,N_7710,N_8335);
nor UO_794 (O_794,N_9840,N_8984);
and UO_795 (O_795,N_9289,N_8362);
nor UO_796 (O_796,N_9387,N_7568);
or UO_797 (O_797,N_9753,N_8241);
nor UO_798 (O_798,N_7698,N_9454);
nor UO_799 (O_799,N_7663,N_9394);
nor UO_800 (O_800,N_7550,N_9266);
xnor UO_801 (O_801,N_9252,N_9042);
and UO_802 (O_802,N_7957,N_9563);
or UO_803 (O_803,N_8998,N_9469);
or UO_804 (O_804,N_9496,N_9486);
nor UO_805 (O_805,N_9445,N_8725);
nor UO_806 (O_806,N_8466,N_9409);
nand UO_807 (O_807,N_7757,N_8015);
or UO_808 (O_808,N_7854,N_9195);
or UO_809 (O_809,N_7765,N_9292);
or UO_810 (O_810,N_8176,N_9452);
or UO_811 (O_811,N_9242,N_9334);
and UO_812 (O_812,N_8753,N_9341);
or UO_813 (O_813,N_8188,N_8443);
nand UO_814 (O_814,N_9503,N_8939);
nor UO_815 (O_815,N_9188,N_7636);
nor UO_816 (O_816,N_9267,N_8288);
or UO_817 (O_817,N_8663,N_9274);
nor UO_818 (O_818,N_7704,N_8122);
nor UO_819 (O_819,N_8561,N_7690);
nand UO_820 (O_820,N_8158,N_9193);
nor UO_821 (O_821,N_9955,N_9173);
or UO_822 (O_822,N_8276,N_9766);
and UO_823 (O_823,N_9683,N_9966);
and UO_824 (O_824,N_9790,N_8838);
nand UO_825 (O_825,N_8803,N_9736);
nor UO_826 (O_826,N_8135,N_7815);
and UO_827 (O_827,N_7662,N_8238);
or UO_828 (O_828,N_9308,N_8871);
and UO_829 (O_829,N_9182,N_8097);
and UO_830 (O_830,N_9830,N_7682);
nor UO_831 (O_831,N_9541,N_7524);
or UO_832 (O_832,N_9091,N_8790);
xnor UO_833 (O_833,N_9420,N_8802);
or UO_834 (O_834,N_8619,N_9354);
nand UO_835 (O_835,N_7883,N_7760);
or UO_836 (O_836,N_9397,N_9379);
and UO_837 (O_837,N_9696,N_9682);
and UO_838 (O_838,N_9167,N_8214);
or UO_839 (O_839,N_9809,N_7800);
or UO_840 (O_840,N_8311,N_9190);
nand UO_841 (O_841,N_8593,N_7937);
or UO_842 (O_842,N_9655,N_7965);
nor UO_843 (O_843,N_8041,N_8269);
and UO_844 (O_844,N_7623,N_8739);
nor UO_845 (O_845,N_8375,N_7849);
and UO_846 (O_846,N_8149,N_7500);
or UO_847 (O_847,N_7645,N_8778);
nand UO_848 (O_848,N_9608,N_9278);
and UO_849 (O_849,N_9005,N_9161);
nand UO_850 (O_850,N_9303,N_7546);
or UO_851 (O_851,N_7634,N_9680);
nand UO_852 (O_852,N_9869,N_8898);
nor UO_853 (O_853,N_8189,N_9560);
xor UO_854 (O_854,N_8955,N_9854);
nand UO_855 (O_855,N_8924,N_9403);
nand UO_856 (O_856,N_9417,N_8837);
or UO_857 (O_857,N_8444,N_9694);
nand UO_858 (O_858,N_8115,N_8758);
nand UO_859 (O_859,N_7522,N_8520);
or UO_860 (O_860,N_7517,N_8638);
or UO_861 (O_861,N_8237,N_8381);
nor UO_862 (O_862,N_9122,N_9491);
xor UO_863 (O_863,N_9996,N_8645);
nand UO_864 (O_864,N_9213,N_7527);
or UO_865 (O_865,N_9269,N_7702);
nor UO_866 (O_866,N_8821,N_9389);
nand UO_867 (O_867,N_7747,N_8756);
or UO_868 (O_868,N_9108,N_7639);
nor UO_869 (O_869,N_9453,N_7599);
nor UO_870 (O_870,N_9222,N_7629);
and UO_871 (O_871,N_8399,N_8429);
nor UO_872 (O_872,N_8980,N_8326);
nor UO_873 (O_873,N_7701,N_9561);
or UO_874 (O_874,N_9943,N_8343);
nand UO_875 (O_875,N_9473,N_9105);
nor UO_876 (O_876,N_7543,N_8745);
and UO_877 (O_877,N_8864,N_7756);
and UO_878 (O_878,N_7959,N_9507);
nand UO_879 (O_879,N_8859,N_9223);
or UO_880 (O_880,N_8267,N_8106);
nand UO_881 (O_881,N_9845,N_9279);
or UO_882 (O_882,N_9012,N_9918);
or UO_883 (O_883,N_8139,N_8105);
nand UO_884 (O_884,N_8374,N_8240);
nand UO_885 (O_885,N_9556,N_9651);
nor UO_886 (O_886,N_9067,N_7539);
nor UO_887 (O_887,N_9965,N_8146);
nor UO_888 (O_888,N_9467,N_7834);
nor UO_889 (O_889,N_9540,N_7858);
nand UO_890 (O_890,N_9894,N_8248);
nand UO_891 (O_891,N_9208,N_9717);
or UO_892 (O_892,N_9224,N_9567);
and UO_893 (O_893,N_8484,N_9577);
nand UO_894 (O_894,N_9922,N_8215);
and UO_895 (O_895,N_9775,N_9415);
or UO_896 (O_896,N_8216,N_7782);
or UO_897 (O_897,N_7656,N_8459);
nand UO_898 (O_898,N_7863,N_8413);
nor UO_899 (O_899,N_7642,N_9307);
or UO_900 (O_900,N_8412,N_8552);
nand UO_901 (O_901,N_7761,N_9782);
or UO_902 (O_902,N_7912,N_9640);
or UO_903 (O_903,N_9280,N_8472);
nand UO_904 (O_904,N_7844,N_9150);
and UO_905 (O_905,N_7949,N_8434);
nand UO_906 (O_906,N_8583,N_9272);
or UO_907 (O_907,N_7638,N_9984);
nand UO_908 (O_908,N_9550,N_8090);
nor UO_909 (O_909,N_8037,N_9853);
or UO_910 (O_910,N_9557,N_7990);
or UO_911 (O_911,N_9072,N_7902);
nand UO_912 (O_912,N_8137,N_9433);
nand UO_913 (O_913,N_7895,N_9060);
and UO_914 (O_914,N_8351,N_8212);
nand UO_915 (O_915,N_8929,N_9964);
or UO_916 (O_916,N_9784,N_9722);
nor UO_917 (O_917,N_7607,N_7814);
or UO_918 (O_918,N_7549,N_9706);
and UO_919 (O_919,N_7940,N_8776);
xnor UO_920 (O_920,N_8626,N_8230);
or UO_921 (O_921,N_7554,N_9358);
and UO_922 (O_922,N_9313,N_7767);
or UO_923 (O_923,N_8008,N_8788);
nor UO_924 (O_924,N_7943,N_7510);
and UO_925 (O_925,N_9841,N_8794);
nand UO_926 (O_926,N_7922,N_9857);
or UO_927 (O_927,N_9058,N_7987);
or UO_928 (O_928,N_8605,N_8879);
or UO_929 (O_929,N_8344,N_8141);
and UO_930 (O_930,N_8201,N_7916);
or UO_931 (O_931,N_7530,N_8372);
and UO_932 (O_932,N_8209,N_8639);
nor UO_933 (O_933,N_9450,N_9806);
or UO_934 (O_934,N_8103,N_7823);
or UO_935 (O_935,N_9605,N_9780);
nand UO_936 (O_936,N_9821,N_7696);
or UO_937 (O_937,N_7856,N_8916);
xnor UO_938 (O_938,N_9329,N_8938);
nand UO_939 (O_939,N_9571,N_8658);
nand UO_940 (O_940,N_7700,N_8239);
nor UO_941 (O_941,N_8521,N_8306);
or UO_942 (O_942,N_9714,N_8502);
nand UO_943 (O_943,N_7617,N_8646);
nor UO_944 (O_944,N_9763,N_8522);
nor UO_945 (O_945,N_9327,N_8873);
nor UO_946 (O_946,N_8506,N_8913);
nand UO_947 (O_947,N_8339,N_9883);
nor UO_948 (O_948,N_9799,N_9191);
or UO_949 (O_949,N_7876,N_8025);
nor UO_950 (O_950,N_9116,N_9533);
and UO_951 (O_951,N_9893,N_8947);
and UO_952 (O_952,N_8540,N_8704);
nand UO_953 (O_953,N_8168,N_8173);
or UO_954 (O_954,N_9710,N_9504);
or UO_955 (O_955,N_9953,N_9282);
or UO_956 (O_956,N_8954,N_9477);
and UO_957 (O_957,N_9708,N_7970);
and UO_958 (O_958,N_8974,N_8033);
nand UO_959 (O_959,N_9249,N_9495);
and UO_960 (O_960,N_9741,N_8752);
nor UO_961 (O_961,N_9976,N_9318);
and UO_962 (O_962,N_8102,N_8589);
nor UO_963 (O_963,N_9330,N_8166);
nor UO_964 (O_964,N_8999,N_8720);
nand UO_965 (O_965,N_7533,N_9291);
or UO_966 (O_966,N_8740,N_8208);
nor UO_967 (O_967,N_9176,N_8014);
nor UO_968 (O_968,N_7627,N_9008);
or UO_969 (O_969,N_7717,N_7758);
or UO_970 (O_970,N_9578,N_9794);
and UO_971 (O_971,N_9003,N_8064);
nor UO_972 (O_972,N_9971,N_9059);
or UO_973 (O_973,N_7744,N_8598);
and UO_974 (O_974,N_7870,N_9987);
nor UO_975 (O_975,N_7555,N_8009);
and UO_976 (O_976,N_9230,N_7684);
nor UO_977 (O_977,N_8594,N_7558);
and UO_978 (O_978,N_9744,N_9543);
or UO_979 (O_979,N_8483,N_8849);
and UO_980 (O_980,N_8498,N_8742);
or UO_981 (O_981,N_9171,N_9439);
nor UO_982 (O_982,N_9534,N_9676);
nor UO_983 (O_983,N_9180,N_7576);
nand UO_984 (O_984,N_8279,N_8094);
or UO_985 (O_985,N_8190,N_9862);
and UO_986 (O_986,N_9910,N_8185);
and UO_987 (O_987,N_7826,N_9572);
nand UO_988 (O_988,N_8470,N_9107);
and UO_989 (O_989,N_7573,N_8622);
nand UO_990 (O_990,N_9196,N_9657);
or UO_991 (O_991,N_9734,N_9836);
and UO_992 (O_992,N_9582,N_9549);
nor UO_993 (O_993,N_8310,N_8695);
and UO_994 (O_994,N_8147,N_7712);
nand UO_995 (O_995,N_9383,N_7582);
nor UO_996 (O_996,N_7693,N_9823);
and UO_997 (O_997,N_8118,N_9833);
nor UO_998 (O_998,N_9848,N_8899);
and UO_999 (O_999,N_8765,N_8028);
nor UO_1000 (O_1000,N_9912,N_9009);
or UO_1001 (O_1001,N_7972,N_9740);
and UO_1002 (O_1002,N_8684,N_9832);
nor UO_1003 (O_1003,N_9925,N_9872);
and UO_1004 (O_1004,N_8337,N_9022);
and UO_1005 (O_1005,N_7666,N_8585);
and UO_1006 (O_1006,N_9598,N_9895);
nor UO_1007 (O_1007,N_8718,N_8719);
nand UO_1008 (O_1008,N_8265,N_8897);
and UO_1009 (O_1009,N_8440,N_9353);
nand UO_1010 (O_1010,N_7724,N_9528);
nor UO_1011 (O_1011,N_9992,N_9281);
and UO_1012 (O_1012,N_7676,N_9981);
and UO_1013 (O_1013,N_9226,N_8772);
or UO_1014 (O_1014,N_8504,N_8198);
or UO_1015 (O_1015,N_9124,N_9234);
nor UO_1016 (O_1016,N_7840,N_8535);
nand UO_1017 (O_1017,N_8548,N_8047);
and UO_1018 (O_1018,N_8376,N_9174);
or UO_1019 (O_1019,N_8830,N_8480);
nor UO_1020 (O_1020,N_7587,N_8634);
nand UO_1021 (O_1021,N_7873,N_9277);
nor UO_1022 (O_1022,N_7998,N_7551);
nor UO_1023 (O_1023,N_9752,N_8547);
nand UO_1024 (O_1024,N_7683,N_7754);
nor UO_1025 (O_1025,N_9765,N_8817);
nand UO_1026 (O_1026,N_7845,N_7731);
nand UO_1027 (O_1027,N_9142,N_8839);
nor UO_1028 (O_1028,N_9078,N_8091);
xnor UO_1029 (O_1029,N_8165,N_9089);
or UO_1030 (O_1030,N_8496,N_8592);
nand UO_1031 (O_1031,N_8603,N_8574);
nand UO_1032 (O_1032,N_9678,N_8858);
nand UO_1033 (O_1033,N_8729,N_7822);
nand UO_1034 (O_1034,N_8272,N_8379);
and UO_1035 (O_1035,N_8770,N_8732);
nor UO_1036 (O_1036,N_9084,N_9407);
nand UO_1037 (O_1037,N_8501,N_8460);
nand UO_1038 (O_1038,N_9144,N_8883);
and UO_1039 (O_1039,N_8935,N_7812);
or UO_1040 (O_1040,N_9390,N_8478);
or UO_1041 (O_1041,N_8304,N_8438);
or UO_1042 (O_1042,N_8011,N_7827);
or UO_1043 (O_1043,N_9999,N_8482);
or UO_1044 (O_1044,N_7806,N_8095);
nor UO_1045 (O_1045,N_7736,N_9593);
nand UO_1046 (O_1046,N_9027,N_7917);
nor UO_1047 (O_1047,N_8063,N_9355);
or UO_1048 (O_1048,N_8366,N_7600);
nor UO_1049 (O_1049,N_8900,N_9517);
nor UO_1050 (O_1050,N_8675,N_9203);
or UO_1051 (O_1051,N_7781,N_9147);
nand UO_1052 (O_1052,N_9685,N_8394);
nor UO_1053 (O_1053,N_7613,N_8184);
or UO_1054 (O_1054,N_7716,N_8331);
and UO_1055 (O_1055,N_8963,N_7992);
and UO_1056 (O_1056,N_8698,N_9527);
or UO_1057 (O_1057,N_8340,N_9102);
nor UO_1058 (O_1058,N_9456,N_9659);
and UO_1059 (O_1059,N_7897,N_8509);
nor UO_1060 (O_1060,N_9615,N_8649);
and UO_1061 (O_1061,N_7835,N_8744);
nand UO_1062 (O_1062,N_9429,N_7609);
and UO_1063 (O_1063,N_8942,N_9482);
nor UO_1064 (O_1064,N_8685,N_8828);
nor UO_1065 (O_1065,N_9422,N_8532);
nand UO_1066 (O_1066,N_9143,N_9941);
nor UO_1067 (O_1067,N_9216,N_9332);
or UO_1068 (O_1068,N_7939,N_9153);
and UO_1069 (O_1069,N_8621,N_9839);
nand UO_1070 (O_1070,N_9998,N_9750);
and UO_1071 (O_1071,N_8641,N_8811);
and UO_1072 (O_1072,N_8111,N_9568);
nand UO_1073 (O_1073,N_9092,N_9695);
nor UO_1074 (O_1074,N_7793,N_9649);
xor UO_1075 (O_1075,N_9817,N_9014);
or UO_1076 (O_1076,N_9573,N_7885);
nand UO_1077 (O_1077,N_9723,N_8071);
and UO_1078 (O_1078,N_9642,N_7907);
or UO_1079 (O_1079,N_9138,N_7687);
or UO_1080 (O_1080,N_8951,N_8218);
and UO_1081 (O_1081,N_8061,N_8664);
and UO_1082 (O_1082,N_9391,N_7585);
xnor UO_1083 (O_1083,N_8656,N_7537);
nand UO_1084 (O_1084,N_8566,N_8659);
or UO_1085 (O_1085,N_9787,N_7595);
nor UO_1086 (O_1086,N_8678,N_8682);
nand UO_1087 (O_1087,N_8493,N_9914);
nor UO_1088 (O_1088,N_7906,N_8089);
nor UO_1089 (O_1089,N_9505,N_9185);
and UO_1090 (O_1090,N_8000,N_7560);
nand UO_1091 (O_1091,N_8242,N_7914);
xor UO_1092 (O_1092,N_9986,N_8676);
and UO_1093 (O_1093,N_9562,N_9989);
or UO_1094 (O_1094,N_9268,N_8953);
nor UO_1095 (O_1095,N_9820,N_7513);
and UO_1096 (O_1096,N_9512,N_9771);
nor UO_1097 (O_1097,N_9634,N_8043);
and UO_1098 (O_1098,N_7799,N_9304);
nand UO_1099 (O_1099,N_9849,N_9982);
or UO_1100 (O_1100,N_7540,N_9440);
xnor UO_1101 (O_1101,N_8093,N_7868);
and UO_1102 (O_1102,N_8287,N_8471);
and UO_1103 (O_1103,N_9751,N_7561);
and UO_1104 (O_1104,N_9345,N_9855);
nand UO_1105 (O_1105,N_7552,N_7526);
and UO_1106 (O_1106,N_7670,N_9874);
nor UO_1107 (O_1107,N_9939,N_8736);
nor UO_1108 (O_1108,N_9347,N_9911);
and UO_1109 (O_1109,N_8796,N_8627);
nand UO_1110 (O_1110,N_9553,N_7564);
or UO_1111 (O_1111,N_8860,N_7860);
nor UO_1112 (O_1112,N_8070,N_9395);
xor UO_1113 (O_1113,N_7920,N_9104);
nor UO_1114 (O_1114,N_8258,N_7753);
nor UO_1115 (O_1115,N_8931,N_9367);
nand UO_1116 (O_1116,N_9169,N_7734);
or UO_1117 (O_1117,N_7635,N_9322);
xor UO_1118 (O_1118,N_7589,N_7577);
nor UO_1119 (O_1119,N_9485,N_9381);
or UO_1120 (O_1120,N_8295,N_8427);
and UO_1121 (O_1121,N_8273,N_9948);
or UO_1122 (O_1122,N_7926,N_9233);
nand UO_1123 (O_1123,N_8021,N_8200);
xor UO_1124 (O_1124,N_9424,N_9421);
nand UO_1125 (O_1125,N_9737,N_7882);
nand UO_1126 (O_1126,N_9726,N_9219);
or UO_1127 (O_1127,N_9724,N_7886);
or UO_1128 (O_1128,N_9592,N_9945);
nor UO_1129 (O_1129,N_8129,N_9926);
and UO_1130 (O_1130,N_8096,N_8690);
and UO_1131 (O_1131,N_9499,N_8577);
nor UO_1132 (O_1132,N_7804,N_7837);
nand UO_1133 (O_1133,N_9382,N_7824);
nand UO_1134 (O_1134,N_9011,N_8056);
nand UO_1135 (O_1135,N_8560,N_9904);
or UO_1136 (O_1136,N_8187,N_7719);
or UO_1137 (O_1137,N_8767,N_8505);
or UO_1138 (O_1138,N_9746,N_8940);
and UO_1139 (O_1139,N_8409,N_8737);
and UO_1140 (O_1140,N_8787,N_8446);
or UO_1141 (O_1141,N_8274,N_7518);
or UO_1142 (O_1142,N_9494,N_8525);
nor UO_1143 (O_1143,N_9637,N_7625);
nand UO_1144 (O_1144,N_9363,N_9074);
and UO_1145 (O_1145,N_8461,N_7933);
or UO_1146 (O_1146,N_8081,N_7942);
nor UO_1147 (O_1147,N_9079,N_9187);
or UO_1148 (O_1148,N_7852,N_7567);
nand UO_1149 (O_1149,N_9393,N_8906);
nand UO_1150 (O_1150,N_8125,N_7892);
nand UO_1151 (O_1151,N_9956,N_8142);
or UO_1152 (O_1152,N_7593,N_8630);
or UO_1153 (O_1153,N_8580,N_8908);
and UO_1154 (O_1154,N_7586,N_8689);
or UO_1155 (O_1155,N_9743,N_9083);
nand UO_1156 (O_1156,N_8284,N_9777);
nand UO_1157 (O_1157,N_8513,N_7980);
and UO_1158 (O_1158,N_9392,N_9949);
nand UO_1159 (O_1159,N_9667,N_9851);
nor UO_1160 (O_1160,N_8382,N_8514);
and UO_1161 (O_1161,N_8084,N_9700);
nand UO_1162 (O_1162,N_8716,N_8031);
or UO_1163 (O_1163,N_9566,N_8824);
or UO_1164 (O_1164,N_9275,N_8490);
or UO_1165 (O_1165,N_9888,N_9352);
and UO_1166 (O_1166,N_9884,N_8109);
or UO_1167 (O_1167,N_8922,N_9813);
or UO_1168 (O_1168,N_8528,N_9372);
nor UO_1169 (O_1169,N_8545,N_9166);
or UO_1170 (O_1170,N_7983,N_9337);
and UO_1171 (O_1171,N_9106,N_7904);
nor UO_1172 (O_1172,N_9075,N_9881);
and UO_1173 (O_1173,N_8280,N_9455);
nor UO_1174 (O_1174,N_7919,N_9675);
or UO_1175 (O_1175,N_9773,N_9137);
or UO_1176 (O_1176,N_9805,N_7699);
nor UO_1177 (O_1177,N_9865,N_7528);
and UO_1178 (O_1178,N_8933,N_7735);
nand UO_1179 (O_1179,N_7643,N_7547);
nor UO_1180 (O_1180,N_7778,N_7986);
nand UO_1181 (O_1181,N_8377,N_9255);
nor UO_1182 (O_1182,N_9892,N_8458);
or UO_1183 (O_1183,N_8053,N_7703);
nor UO_1184 (O_1184,N_8861,N_8027);
nor UO_1185 (O_1185,N_8612,N_8896);
or UO_1186 (O_1186,N_8635,N_8316);
or UO_1187 (O_1187,N_8055,N_9298);
and UO_1188 (O_1188,N_7726,N_8161);
or UO_1189 (O_1189,N_8909,N_8712);
nor UO_1190 (O_1190,N_9069,N_9879);
nor UO_1191 (O_1191,N_9915,N_8653);
or UO_1192 (O_1192,N_8611,N_9522);
or UO_1193 (O_1193,N_8396,N_9235);
nor UO_1194 (O_1194,N_8271,N_8078);
and UO_1195 (O_1195,N_9101,N_9610);
or UO_1196 (O_1196,N_8497,N_8553);
or UO_1197 (O_1197,N_7580,N_8112);
and UO_1198 (O_1198,N_7512,N_8431);
xnor UO_1199 (O_1199,N_9778,N_8481);
nand UO_1200 (O_1200,N_7620,N_9472);
nand UO_1201 (O_1201,N_8958,N_7908);
nand UO_1202 (O_1202,N_7961,N_9957);
nand UO_1203 (O_1203,N_8833,N_7711);
and UO_1204 (O_1204,N_9015,N_9370);
nand UO_1205 (O_1205,N_8018,N_8687);
and UO_1206 (O_1206,N_9601,N_8867);
nand UO_1207 (O_1207,N_8832,N_8235);
and UO_1208 (O_1208,N_9599,N_9017);
and UO_1209 (O_1209,N_7668,N_9296);
nand UO_1210 (O_1210,N_9891,N_9316);
or UO_1211 (O_1211,N_8463,N_8296);
nand UO_1212 (O_1212,N_8783,N_9900);
nor UO_1213 (O_1213,N_8075,N_8760);
or UO_1214 (O_1214,N_8629,N_9489);
and UO_1215 (O_1215,N_8225,N_9843);
nor UO_1216 (O_1216,N_8006,N_8249);
nor UO_1217 (O_1217,N_7506,N_8981);
nor UO_1218 (O_1218,N_8733,N_8565);
xnor UO_1219 (O_1219,N_9158,N_9324);
nand UO_1220 (O_1220,N_9581,N_9804);
xnor UO_1221 (O_1221,N_9691,N_8100);
and UO_1222 (O_1222,N_7641,N_8178);
nand UO_1223 (O_1223,N_7979,N_8286);
and UO_1224 (O_1224,N_8599,N_7944);
or UO_1225 (O_1225,N_9791,N_8518);
or UO_1226 (O_1226,N_9681,N_8539);
and UO_1227 (O_1227,N_7976,N_9583);
nor UO_1228 (O_1228,N_8616,N_7791);
nor UO_1229 (O_1229,N_7941,N_8246);
and UO_1230 (O_1230,N_7956,N_8534);
nor UO_1231 (O_1231,N_9514,N_8229);
nand UO_1232 (O_1232,N_8065,N_8410);
and UO_1233 (O_1233,N_7861,N_7792);
nor UO_1234 (O_1234,N_8516,N_8905);
nor UO_1235 (O_1235,N_8894,N_9729);
nor UO_1236 (O_1236,N_9063,N_8968);
nand UO_1237 (O_1237,N_9326,N_9290);
nor UO_1238 (O_1238,N_9061,N_8717);
and UO_1239 (O_1239,N_9650,N_9621);
or UO_1240 (O_1240,N_8691,N_8637);
or UO_1241 (O_1241,N_9959,N_8451);
or UO_1242 (O_1242,N_8491,N_8003);
nor UO_1243 (O_1243,N_7621,N_8001);
nand UO_1244 (O_1244,N_9309,N_9693);
or UO_1245 (O_1245,N_8301,N_9596);
nor UO_1246 (O_1246,N_9217,N_8538);
and UO_1247 (O_1247,N_9340,N_9319);
nor UO_1248 (O_1248,N_9416,N_8403);
or UO_1249 (O_1249,N_9333,N_8527);
nand UO_1250 (O_1250,N_8386,N_7659);
or UO_1251 (O_1251,N_8093,N_9395);
nor UO_1252 (O_1252,N_9606,N_8075);
or UO_1253 (O_1253,N_8050,N_8454);
and UO_1254 (O_1254,N_9498,N_9165);
or UO_1255 (O_1255,N_9909,N_8467);
nor UO_1256 (O_1256,N_7775,N_8121);
or UO_1257 (O_1257,N_7796,N_9683);
nand UO_1258 (O_1258,N_7992,N_8322);
and UO_1259 (O_1259,N_7570,N_7730);
nor UO_1260 (O_1260,N_8859,N_8039);
nor UO_1261 (O_1261,N_8487,N_8101);
nand UO_1262 (O_1262,N_9150,N_9411);
nor UO_1263 (O_1263,N_9521,N_8158);
nor UO_1264 (O_1264,N_8169,N_9436);
and UO_1265 (O_1265,N_7907,N_7519);
and UO_1266 (O_1266,N_9325,N_9277);
nor UO_1267 (O_1267,N_8228,N_9610);
or UO_1268 (O_1268,N_8727,N_7728);
nor UO_1269 (O_1269,N_9174,N_8080);
or UO_1270 (O_1270,N_9326,N_8109);
nor UO_1271 (O_1271,N_8345,N_7565);
or UO_1272 (O_1272,N_9036,N_9277);
nor UO_1273 (O_1273,N_9606,N_9134);
or UO_1274 (O_1274,N_8336,N_9130);
and UO_1275 (O_1275,N_9383,N_7529);
and UO_1276 (O_1276,N_8334,N_8262);
or UO_1277 (O_1277,N_8831,N_8108);
or UO_1278 (O_1278,N_8089,N_7716);
nand UO_1279 (O_1279,N_8366,N_9822);
or UO_1280 (O_1280,N_9171,N_8934);
nand UO_1281 (O_1281,N_8424,N_8371);
and UO_1282 (O_1282,N_8494,N_8929);
or UO_1283 (O_1283,N_8267,N_8215);
and UO_1284 (O_1284,N_8319,N_7739);
and UO_1285 (O_1285,N_9462,N_8725);
and UO_1286 (O_1286,N_8714,N_9661);
or UO_1287 (O_1287,N_8083,N_8232);
or UO_1288 (O_1288,N_8862,N_7668);
or UO_1289 (O_1289,N_8412,N_8112);
nor UO_1290 (O_1290,N_7819,N_9625);
or UO_1291 (O_1291,N_8706,N_8515);
nand UO_1292 (O_1292,N_7610,N_9715);
nand UO_1293 (O_1293,N_9119,N_9412);
and UO_1294 (O_1294,N_8188,N_9085);
or UO_1295 (O_1295,N_8353,N_9894);
nand UO_1296 (O_1296,N_9662,N_8796);
and UO_1297 (O_1297,N_9173,N_9655);
nand UO_1298 (O_1298,N_8687,N_8177);
or UO_1299 (O_1299,N_7940,N_8727);
xor UO_1300 (O_1300,N_8889,N_8791);
or UO_1301 (O_1301,N_8434,N_8140);
nand UO_1302 (O_1302,N_9665,N_8803);
and UO_1303 (O_1303,N_9214,N_7820);
or UO_1304 (O_1304,N_9371,N_7621);
nor UO_1305 (O_1305,N_8037,N_7811);
and UO_1306 (O_1306,N_8876,N_7976);
nand UO_1307 (O_1307,N_9178,N_8290);
nor UO_1308 (O_1308,N_8449,N_8811);
nand UO_1309 (O_1309,N_9305,N_8654);
nand UO_1310 (O_1310,N_7785,N_8000);
nor UO_1311 (O_1311,N_8063,N_9872);
and UO_1312 (O_1312,N_9169,N_9899);
nor UO_1313 (O_1313,N_7740,N_9915);
nor UO_1314 (O_1314,N_9828,N_9470);
nor UO_1315 (O_1315,N_8098,N_9041);
nand UO_1316 (O_1316,N_9108,N_7830);
and UO_1317 (O_1317,N_8844,N_8681);
or UO_1318 (O_1318,N_9111,N_8076);
and UO_1319 (O_1319,N_9967,N_8306);
and UO_1320 (O_1320,N_9348,N_7787);
nand UO_1321 (O_1321,N_8551,N_9973);
or UO_1322 (O_1322,N_7781,N_9020);
and UO_1323 (O_1323,N_7770,N_9088);
or UO_1324 (O_1324,N_8789,N_8817);
or UO_1325 (O_1325,N_9040,N_9047);
nor UO_1326 (O_1326,N_9932,N_8546);
nand UO_1327 (O_1327,N_9706,N_8415);
nand UO_1328 (O_1328,N_9164,N_8564);
nand UO_1329 (O_1329,N_8925,N_9276);
and UO_1330 (O_1330,N_9268,N_9512);
and UO_1331 (O_1331,N_7918,N_7670);
nand UO_1332 (O_1332,N_9263,N_9803);
or UO_1333 (O_1333,N_7812,N_8641);
or UO_1334 (O_1334,N_8021,N_9598);
nor UO_1335 (O_1335,N_8790,N_8954);
nand UO_1336 (O_1336,N_8015,N_9223);
or UO_1337 (O_1337,N_8169,N_9410);
nor UO_1338 (O_1338,N_8666,N_9522);
nand UO_1339 (O_1339,N_9831,N_9199);
nor UO_1340 (O_1340,N_9386,N_7903);
and UO_1341 (O_1341,N_9466,N_9089);
nand UO_1342 (O_1342,N_8911,N_8198);
nor UO_1343 (O_1343,N_8296,N_8198);
and UO_1344 (O_1344,N_7517,N_8500);
and UO_1345 (O_1345,N_9775,N_7968);
xor UO_1346 (O_1346,N_9907,N_9611);
nand UO_1347 (O_1347,N_8105,N_9657);
nor UO_1348 (O_1348,N_7725,N_7898);
or UO_1349 (O_1349,N_8596,N_9168);
nand UO_1350 (O_1350,N_9387,N_9739);
or UO_1351 (O_1351,N_8852,N_8089);
nand UO_1352 (O_1352,N_9699,N_8499);
and UO_1353 (O_1353,N_8704,N_9434);
nand UO_1354 (O_1354,N_9957,N_9249);
and UO_1355 (O_1355,N_8360,N_9525);
and UO_1356 (O_1356,N_8321,N_7978);
and UO_1357 (O_1357,N_8097,N_8749);
and UO_1358 (O_1358,N_8217,N_7730);
and UO_1359 (O_1359,N_9118,N_7581);
nand UO_1360 (O_1360,N_7768,N_8278);
and UO_1361 (O_1361,N_8174,N_9535);
nand UO_1362 (O_1362,N_8903,N_8582);
and UO_1363 (O_1363,N_9287,N_9418);
nand UO_1364 (O_1364,N_8471,N_9050);
nor UO_1365 (O_1365,N_9815,N_8132);
and UO_1366 (O_1366,N_7597,N_8117);
or UO_1367 (O_1367,N_9184,N_8226);
and UO_1368 (O_1368,N_9941,N_9110);
nand UO_1369 (O_1369,N_9600,N_7548);
and UO_1370 (O_1370,N_8874,N_7610);
or UO_1371 (O_1371,N_7701,N_7885);
nand UO_1372 (O_1372,N_9926,N_9931);
xnor UO_1373 (O_1373,N_9180,N_7975);
and UO_1374 (O_1374,N_8645,N_9169);
or UO_1375 (O_1375,N_8878,N_8215);
or UO_1376 (O_1376,N_9622,N_8905);
or UO_1377 (O_1377,N_8085,N_8530);
and UO_1378 (O_1378,N_8100,N_9150);
nand UO_1379 (O_1379,N_8470,N_9925);
nand UO_1380 (O_1380,N_9346,N_8572);
nand UO_1381 (O_1381,N_8782,N_8966);
nand UO_1382 (O_1382,N_7965,N_9886);
nor UO_1383 (O_1383,N_8523,N_9306);
nor UO_1384 (O_1384,N_8289,N_9821);
or UO_1385 (O_1385,N_7925,N_9940);
nand UO_1386 (O_1386,N_7916,N_8623);
nor UO_1387 (O_1387,N_7982,N_8698);
or UO_1388 (O_1388,N_9790,N_7528);
nor UO_1389 (O_1389,N_7964,N_9095);
and UO_1390 (O_1390,N_8798,N_9223);
nand UO_1391 (O_1391,N_9535,N_9931);
and UO_1392 (O_1392,N_7948,N_9016);
or UO_1393 (O_1393,N_7909,N_8262);
and UO_1394 (O_1394,N_9991,N_9405);
or UO_1395 (O_1395,N_9470,N_9367);
or UO_1396 (O_1396,N_9818,N_9434);
nor UO_1397 (O_1397,N_9764,N_9723);
or UO_1398 (O_1398,N_8412,N_7849);
nor UO_1399 (O_1399,N_9341,N_8388);
xnor UO_1400 (O_1400,N_7920,N_8526);
nor UO_1401 (O_1401,N_9911,N_8943);
nand UO_1402 (O_1402,N_9099,N_8037);
nand UO_1403 (O_1403,N_9879,N_7932);
nor UO_1404 (O_1404,N_8946,N_7915);
and UO_1405 (O_1405,N_7676,N_9669);
or UO_1406 (O_1406,N_9672,N_9835);
or UO_1407 (O_1407,N_8591,N_7746);
and UO_1408 (O_1408,N_8572,N_9492);
or UO_1409 (O_1409,N_9837,N_9117);
nand UO_1410 (O_1410,N_7809,N_8705);
and UO_1411 (O_1411,N_9049,N_8163);
or UO_1412 (O_1412,N_8422,N_8799);
nand UO_1413 (O_1413,N_9778,N_8711);
or UO_1414 (O_1414,N_9398,N_9740);
and UO_1415 (O_1415,N_8156,N_9797);
nand UO_1416 (O_1416,N_9814,N_8444);
nor UO_1417 (O_1417,N_8691,N_9719);
nor UO_1418 (O_1418,N_7796,N_9446);
nor UO_1419 (O_1419,N_9418,N_9413);
and UO_1420 (O_1420,N_8196,N_7989);
nor UO_1421 (O_1421,N_9905,N_8040);
or UO_1422 (O_1422,N_9902,N_9352);
nand UO_1423 (O_1423,N_7893,N_9755);
nor UO_1424 (O_1424,N_9523,N_9350);
and UO_1425 (O_1425,N_7712,N_9435);
nor UO_1426 (O_1426,N_8792,N_8298);
and UO_1427 (O_1427,N_9222,N_9023);
nor UO_1428 (O_1428,N_9763,N_7507);
nor UO_1429 (O_1429,N_8915,N_7660);
or UO_1430 (O_1430,N_9884,N_8940);
and UO_1431 (O_1431,N_9906,N_9084);
nor UO_1432 (O_1432,N_9316,N_8529);
and UO_1433 (O_1433,N_8097,N_7625);
nand UO_1434 (O_1434,N_7912,N_8359);
and UO_1435 (O_1435,N_8085,N_8898);
nand UO_1436 (O_1436,N_8131,N_8232);
or UO_1437 (O_1437,N_9739,N_9947);
nor UO_1438 (O_1438,N_8182,N_8782);
xor UO_1439 (O_1439,N_9235,N_9494);
nor UO_1440 (O_1440,N_7524,N_8110);
nor UO_1441 (O_1441,N_9592,N_9324);
nor UO_1442 (O_1442,N_8639,N_8002);
or UO_1443 (O_1443,N_9027,N_8458);
and UO_1444 (O_1444,N_8203,N_9742);
and UO_1445 (O_1445,N_7607,N_7989);
and UO_1446 (O_1446,N_9609,N_8695);
and UO_1447 (O_1447,N_9893,N_8037);
and UO_1448 (O_1448,N_7973,N_8223);
and UO_1449 (O_1449,N_9689,N_9967);
nor UO_1450 (O_1450,N_7813,N_8294);
or UO_1451 (O_1451,N_9957,N_9745);
or UO_1452 (O_1452,N_9729,N_9977);
and UO_1453 (O_1453,N_8598,N_9947);
nand UO_1454 (O_1454,N_8712,N_9923);
and UO_1455 (O_1455,N_8034,N_8169);
nand UO_1456 (O_1456,N_7758,N_8090);
and UO_1457 (O_1457,N_7973,N_9942);
and UO_1458 (O_1458,N_9769,N_8254);
and UO_1459 (O_1459,N_7660,N_9413);
or UO_1460 (O_1460,N_8754,N_7759);
or UO_1461 (O_1461,N_8727,N_7948);
nand UO_1462 (O_1462,N_8851,N_8309);
or UO_1463 (O_1463,N_7853,N_8019);
or UO_1464 (O_1464,N_9486,N_8781);
and UO_1465 (O_1465,N_8910,N_8995);
or UO_1466 (O_1466,N_8355,N_9558);
nor UO_1467 (O_1467,N_8770,N_8865);
nor UO_1468 (O_1468,N_8984,N_8791);
or UO_1469 (O_1469,N_7671,N_8740);
or UO_1470 (O_1470,N_8009,N_8840);
xor UO_1471 (O_1471,N_7677,N_9314);
nand UO_1472 (O_1472,N_7883,N_8157);
nand UO_1473 (O_1473,N_8854,N_7679);
nor UO_1474 (O_1474,N_7520,N_8494);
and UO_1475 (O_1475,N_9169,N_8038);
nand UO_1476 (O_1476,N_8730,N_8117);
nor UO_1477 (O_1477,N_9570,N_9107);
and UO_1478 (O_1478,N_9021,N_8293);
nor UO_1479 (O_1479,N_8781,N_7839);
nand UO_1480 (O_1480,N_7822,N_9620);
nor UO_1481 (O_1481,N_9124,N_7696);
and UO_1482 (O_1482,N_8105,N_9520);
or UO_1483 (O_1483,N_9328,N_7982);
and UO_1484 (O_1484,N_8701,N_7514);
nand UO_1485 (O_1485,N_7836,N_7897);
or UO_1486 (O_1486,N_9937,N_9892);
and UO_1487 (O_1487,N_8352,N_7867);
nor UO_1488 (O_1488,N_9564,N_7999);
nor UO_1489 (O_1489,N_7717,N_9109);
and UO_1490 (O_1490,N_8141,N_9601);
or UO_1491 (O_1491,N_9712,N_9826);
nand UO_1492 (O_1492,N_8896,N_7800);
nor UO_1493 (O_1493,N_9447,N_7873);
and UO_1494 (O_1494,N_8358,N_8104);
nor UO_1495 (O_1495,N_7568,N_8921);
nand UO_1496 (O_1496,N_9830,N_8549);
or UO_1497 (O_1497,N_9629,N_9025);
and UO_1498 (O_1498,N_9661,N_8264);
nor UO_1499 (O_1499,N_8613,N_9328);
endmodule