module basic_1000_10000_1500_2_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5009,N_5010,N_5011,N_5012,N_5014,N_5018,N_5019,N_5020,N_5021,N_5022,N_5025,N_5028,N_5031,N_5033,N_5036,N_5038,N_5041,N_5043,N_5048,N_5049,N_5050,N_5051,N_5054,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5067,N_5068,N_5070,N_5072,N_5075,N_5076,N_5077,N_5079,N_5083,N_5085,N_5088,N_5090,N_5091,N_5092,N_5093,N_5095,N_5101,N_5102,N_5103,N_5105,N_5106,N_5109,N_5111,N_5112,N_5116,N_5117,N_5121,N_5124,N_5126,N_5129,N_5130,N_5131,N_5135,N_5136,N_5146,N_5147,N_5151,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5164,N_5165,N_5167,N_5168,N_5172,N_5176,N_5177,N_5180,N_5183,N_5185,N_5186,N_5187,N_5189,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5202,N_5203,N_5205,N_5206,N_5208,N_5209,N_5210,N_5211,N_5217,N_5218,N_5220,N_5222,N_5224,N_5227,N_5228,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5245,N_5246,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5256,N_5257,N_5258,N_5259,N_5260,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5269,N_5271,N_5272,N_5273,N_5274,N_5275,N_5278,N_5282,N_5284,N_5285,N_5287,N_5293,N_5294,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5304,N_5305,N_5308,N_5309,N_5310,N_5312,N_5314,N_5316,N_5317,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5328,N_5329,N_5331,N_5332,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5347,N_5348,N_5350,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5364,N_5365,N_5366,N_5369,N_5371,N_5372,N_5376,N_5377,N_5380,N_5382,N_5383,N_5387,N_5388,N_5390,N_5391,N_5392,N_5395,N_5396,N_5397,N_5398,N_5399,N_5402,N_5403,N_5404,N_5405,N_5406,N_5408,N_5410,N_5412,N_5414,N_5415,N_5416,N_5417,N_5419,N_5420,N_5422,N_5423,N_5424,N_5429,N_5431,N_5433,N_5436,N_5437,N_5440,N_5441,N_5442,N_5443,N_5444,N_5446,N_5447,N_5449,N_5450,N_5451,N_5452,N_5453,N_5456,N_5457,N_5460,N_5466,N_5467,N_5470,N_5471,N_5473,N_5475,N_5479,N_5483,N_5485,N_5487,N_5489,N_5493,N_5494,N_5495,N_5497,N_5499,N_5501,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5510,N_5511,N_5512,N_5516,N_5518,N_5519,N_5521,N_5524,N_5525,N_5528,N_5529,N_5530,N_5531,N_5532,N_5534,N_5535,N_5537,N_5539,N_5540,N_5542,N_5543,N_5544,N_5549,N_5551,N_5552,N_5553,N_5555,N_5556,N_5557,N_5560,N_5561,N_5563,N_5566,N_5567,N_5568,N_5569,N_5570,N_5574,N_5576,N_5579,N_5580,N_5582,N_5583,N_5585,N_5587,N_5590,N_5594,N_5595,N_5597,N_5600,N_5601,N_5603,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5624,N_5625,N_5626,N_5627,N_5628,N_5630,N_5632,N_5633,N_5634,N_5635,N_5639,N_5640,N_5642,N_5643,N_5645,N_5646,N_5648,N_5649,N_5651,N_5653,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5662,N_5667,N_5668,N_5669,N_5671,N_5672,N_5673,N_5674,N_5678,N_5680,N_5684,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5696,N_5697,N_5698,N_5700,N_5702,N_5704,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5714,N_5722,N_5724,N_5726,N_5727,N_5728,N_5730,N_5733,N_5734,N_5736,N_5740,N_5741,N_5743,N_5744,N_5745,N_5747,N_5748,N_5751,N_5752,N_5753,N_5754,N_5755,N_5762,N_5763,N_5765,N_5768,N_5770,N_5772,N_5773,N_5774,N_5775,N_5778,N_5779,N_5780,N_5784,N_5787,N_5789,N_5792,N_5793,N_5796,N_5797,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5807,N_5811,N_5812,N_5813,N_5814,N_5816,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5840,N_5841,N_5843,N_5844,N_5848,N_5849,N_5850,N_5851,N_5853,N_5855,N_5859,N_5861,N_5863,N_5864,N_5865,N_5867,N_5870,N_5872,N_5874,N_5875,N_5878,N_5879,N_5882,N_5883,N_5884,N_5885,N_5887,N_5889,N_5890,N_5891,N_5893,N_5894,N_5895,N_5896,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5909,N_5910,N_5912,N_5914,N_5915,N_5916,N_5917,N_5918,N_5920,N_5926,N_5927,N_5929,N_5935,N_5936,N_5937,N_5941,N_5942,N_5946,N_5949,N_5950,N_5951,N_5956,N_5958,N_5962,N_5964,N_5965,N_5966,N_5967,N_5970,N_5972,N_5974,N_5975,N_5976,N_5977,N_5978,N_5980,N_5982,N_5983,N_5985,N_5986,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5998,N_6004,N_6007,N_6008,N_6011,N_6013,N_6014,N_6015,N_6016,N_6020,N_6021,N_6022,N_6023,N_6024,N_6026,N_6027,N_6029,N_6032,N_6034,N_6035,N_6039,N_6041,N_6045,N_6048,N_6049,N_6050,N_6051,N_6052,N_6056,N_6057,N_6058,N_6059,N_6062,N_6063,N_6064,N_6065,N_6066,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6075,N_6076,N_6077,N_6078,N_6080,N_6082,N_6086,N_6087,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6099,N_6102,N_6103,N_6104,N_6106,N_6107,N_6108,N_6110,N_6112,N_6113,N_6115,N_6118,N_6121,N_6122,N_6123,N_6124,N_6125,N_6127,N_6129,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6139,N_6142,N_6143,N_6144,N_6146,N_6147,N_6148,N_6149,N_6151,N_6153,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6162,N_6164,N_6165,N_6167,N_6168,N_6169,N_6173,N_6174,N_6175,N_6176,N_6177,N_6179,N_6181,N_6182,N_6186,N_6187,N_6188,N_6189,N_6190,N_6192,N_6195,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6206,N_6209,N_6210,N_6212,N_6214,N_6216,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6230,N_6233,N_6235,N_6236,N_6237,N_6238,N_6239,N_6241,N_6244,N_6245,N_6247,N_6250,N_6251,N_6252,N_6255,N_6257,N_6258,N_6260,N_6262,N_6265,N_6266,N_6269,N_6270,N_6271,N_6273,N_6275,N_6276,N_6278,N_6280,N_6286,N_6287,N_6289,N_6290,N_6291,N_6294,N_6296,N_6302,N_6306,N_6307,N_6308,N_6310,N_6312,N_6313,N_6314,N_6316,N_6317,N_6318,N_6320,N_6321,N_6322,N_6325,N_6326,N_6328,N_6333,N_6334,N_6335,N_6336,N_6337,N_6340,N_6342,N_6344,N_6346,N_6352,N_6355,N_6356,N_6358,N_6359,N_6360,N_6363,N_6364,N_6365,N_6366,N_6370,N_6371,N_6373,N_6375,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6384,N_6386,N_6387,N_6388,N_6389,N_6390,N_6392,N_6393,N_6395,N_6396,N_6398,N_6399,N_6400,N_6401,N_6402,N_6405,N_6409,N_6410,N_6411,N_6414,N_6415,N_6417,N_6419,N_6421,N_6422,N_6423,N_6424,N_6429,N_6430,N_6431,N_6433,N_6434,N_6436,N_6437,N_6438,N_6439,N_6441,N_6443,N_6446,N_6449,N_6450,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6463,N_6466,N_6468,N_6469,N_6472,N_6473,N_6475,N_6477,N_6479,N_6480,N_6481,N_6483,N_6484,N_6488,N_6490,N_6493,N_6494,N_6495,N_6497,N_6498,N_6499,N_6501,N_6502,N_6503,N_6507,N_6510,N_6513,N_6515,N_6516,N_6517,N_6519,N_6520,N_6522,N_6523,N_6530,N_6531,N_6533,N_6534,N_6535,N_6538,N_6539,N_6540,N_6542,N_6543,N_6545,N_6546,N_6547,N_6549,N_6552,N_6553,N_6554,N_6555,N_6558,N_6559,N_6561,N_6562,N_6565,N_6569,N_6570,N_6573,N_6575,N_6576,N_6577,N_6578,N_6579,N_6581,N_6582,N_6584,N_6587,N_6591,N_6593,N_6594,N_6596,N_6597,N_6599,N_6600,N_6602,N_6603,N_6604,N_6605,N_6607,N_6608,N_6610,N_6612,N_6613,N_6617,N_6619,N_6623,N_6626,N_6627,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6636,N_6637,N_6640,N_6641,N_6643,N_6647,N_6648,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6660,N_6661,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6672,N_6673,N_6674,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6690,N_6691,N_6692,N_6693,N_6695,N_6696,N_6697,N_6700,N_6701,N_6702,N_6704,N_6705,N_6707,N_6708,N_6710,N_6711,N_6715,N_6718,N_6719,N_6722,N_6724,N_6727,N_6728,N_6729,N_6730,N_6732,N_6733,N_6734,N_6735,N_6737,N_6739,N_6740,N_6742,N_6745,N_6747,N_6748,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6767,N_6769,N_6770,N_6771,N_6772,N_6773,N_6775,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6786,N_6788,N_6789,N_6792,N_6793,N_6796,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6818,N_6820,N_6822,N_6823,N_6826,N_6827,N_6828,N_6830,N_6831,N_6834,N_6835,N_6836,N_6837,N_6838,N_6840,N_6841,N_6843,N_6847,N_6848,N_6851,N_6852,N_6853,N_6854,N_6855,N_6857,N_6858,N_6859,N_6860,N_6861,N_6863,N_6865,N_6866,N_6867,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6880,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6891,N_6893,N_6894,N_6896,N_6897,N_6899,N_6900,N_6903,N_6904,N_6906,N_6910,N_6914,N_6916,N_6920,N_6921,N_6923,N_6924,N_6927,N_6929,N_6930,N_6932,N_6935,N_6936,N_6937,N_6940,N_6942,N_6943,N_6944,N_6945,N_6947,N_6948,N_6949,N_6954,N_6956,N_6957,N_6959,N_6960,N_6961,N_6962,N_6964,N_6965,N_6966,N_6969,N_6970,N_6972,N_6976,N_6978,N_6982,N_6985,N_6987,N_6988,N_6989,N_6990,N_6992,N_6993,N_6994,N_6996,N_6997,N_6998,N_6999,N_7000,N_7004,N_7005,N_7009,N_7010,N_7012,N_7014,N_7016,N_7017,N_7018,N_7022,N_7026,N_7027,N_7028,N_7029,N_7031,N_7032,N_7033,N_7035,N_7036,N_7037,N_7038,N_7039,N_7045,N_7046,N_7048,N_7050,N_7053,N_7054,N_7056,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7068,N_7071,N_7072,N_7073,N_7075,N_7079,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7092,N_7093,N_7095,N_7096,N_7097,N_7098,N_7100,N_7101,N_7102,N_7103,N_7105,N_7106,N_7109,N_7111,N_7112,N_7113,N_7117,N_7118,N_7119,N_7121,N_7122,N_7123,N_7125,N_7126,N_7128,N_7130,N_7131,N_7133,N_7134,N_7139,N_7140,N_7141,N_7142,N_7143,N_7147,N_7148,N_7150,N_7151,N_7152,N_7153,N_7155,N_7159,N_7160,N_7162,N_7163,N_7165,N_7167,N_7168,N_7169,N_7172,N_7174,N_7175,N_7177,N_7178,N_7180,N_7183,N_7184,N_7185,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7198,N_7199,N_7201,N_7204,N_7205,N_7206,N_7209,N_7210,N_7212,N_7214,N_7216,N_7219,N_7220,N_7222,N_7226,N_7227,N_7230,N_7231,N_7232,N_7233,N_7235,N_7237,N_7238,N_7240,N_7241,N_7242,N_7244,N_7246,N_7247,N_7249,N_7251,N_7252,N_7254,N_7255,N_7258,N_7259,N_7260,N_7264,N_7266,N_7267,N_7268,N_7271,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7281,N_7282,N_7283,N_7286,N_7292,N_7294,N_7295,N_7297,N_7298,N_7299,N_7300,N_7302,N_7304,N_7305,N_7308,N_7310,N_7311,N_7313,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7322,N_7323,N_7325,N_7328,N_7329,N_7330,N_7331,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7340,N_7343,N_7344,N_7345,N_7346,N_7347,N_7352,N_7353,N_7354,N_7358,N_7359,N_7360,N_7361,N_7362,N_7365,N_7368,N_7371,N_7373,N_7374,N_7375,N_7376,N_7377,N_7379,N_7380,N_7381,N_7384,N_7387,N_7388,N_7390,N_7393,N_7394,N_7395,N_7396,N_7399,N_7400,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7410,N_7416,N_7417,N_7420,N_7421,N_7422,N_7423,N_7427,N_7428,N_7432,N_7435,N_7439,N_7441,N_7442,N_7443,N_7447,N_7449,N_7450,N_7452,N_7455,N_7457,N_7458,N_7459,N_7460,N_7461,N_7463,N_7464,N_7466,N_7467,N_7468,N_7469,N_7470,N_7473,N_7476,N_7478,N_7479,N_7480,N_7481,N_7483,N_7484,N_7486,N_7488,N_7492,N_7493,N_7494,N_7495,N_7498,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7513,N_7516,N_7517,N_7520,N_7522,N_7523,N_7526,N_7527,N_7530,N_7531,N_7532,N_7536,N_7537,N_7538,N_7540,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7550,N_7551,N_7552,N_7555,N_7556,N_7557,N_7559,N_7562,N_7563,N_7566,N_7567,N_7569,N_7571,N_7572,N_7573,N_7575,N_7577,N_7578,N_7579,N_7580,N_7582,N_7583,N_7585,N_7586,N_7588,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7598,N_7599,N_7601,N_7604,N_7605,N_7606,N_7607,N_7609,N_7611,N_7612,N_7615,N_7616,N_7617,N_7618,N_7620,N_7621,N_7622,N_7624,N_7626,N_7628,N_7629,N_7630,N_7631,N_7634,N_7637,N_7638,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7650,N_7651,N_7652,N_7653,N_7657,N_7658,N_7659,N_7660,N_7661,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7676,N_7678,N_7679,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7693,N_7695,N_7696,N_7697,N_7698,N_7699,N_7701,N_7702,N_7703,N_7704,N_7707,N_7709,N_7710,N_7712,N_7714,N_7715,N_7716,N_7717,N_7719,N_7720,N_7721,N_7724,N_7725,N_7727,N_7728,N_7729,N_7730,N_7732,N_7733,N_7734,N_7735,N_7737,N_7738,N_7739,N_7741,N_7747,N_7749,N_7750,N_7751,N_7752,N_7754,N_7756,N_7758,N_7759,N_7760,N_7762,N_7763,N_7764,N_7765,N_7766,N_7768,N_7769,N_7770,N_7772,N_7774,N_7776,N_7777,N_7779,N_7780,N_7781,N_7783,N_7785,N_7786,N_7787,N_7788,N_7790,N_7792,N_7794,N_7795,N_7799,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7808,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7818,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7829,N_7830,N_7833,N_7835,N_7836,N_7837,N_7838,N_7841,N_7842,N_7843,N_7845,N_7846,N_7848,N_7849,N_7850,N_7851,N_7853,N_7854,N_7856,N_7857,N_7858,N_7859,N_7860,N_7866,N_7869,N_7870,N_7873,N_7874,N_7875,N_7876,N_7880,N_7881,N_7883,N_7884,N_7885,N_7888,N_7890,N_7891,N_7894,N_7895,N_7897,N_7900,N_7901,N_7902,N_7903,N_7907,N_7910,N_7911,N_7912,N_7916,N_7919,N_7921,N_7922,N_7923,N_7924,N_7925,N_7928,N_7929,N_7931,N_7932,N_7933,N_7935,N_7937,N_7938,N_7939,N_7943,N_7945,N_7950,N_7951,N_7952,N_7953,N_7956,N_7961,N_7962,N_7963,N_7964,N_7970,N_7971,N_7973,N_7974,N_7975,N_7977,N_7978,N_7980,N_7981,N_7982,N_7983,N_7984,N_7987,N_7988,N_7989,N_7990,N_7993,N_7994,N_7995,N_7996,N_7999,N_8001,N_8003,N_8004,N_8006,N_8007,N_8011,N_8012,N_8013,N_8014,N_8016,N_8017,N_8018,N_8019,N_8021,N_8022,N_8027,N_8028,N_8029,N_8031,N_8032,N_8034,N_8036,N_8037,N_8038,N_8039,N_8043,N_8044,N_8046,N_8048,N_8049,N_8051,N_8052,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8062,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8072,N_8076,N_8077,N_8078,N_8081,N_8084,N_8085,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8094,N_8095,N_8096,N_8097,N_8100,N_8101,N_8102,N_8104,N_8105,N_8109,N_8110,N_8111,N_8116,N_8117,N_8118,N_8119,N_8123,N_8124,N_8127,N_8131,N_8134,N_8136,N_8137,N_8139,N_8145,N_8146,N_8147,N_8148,N_8149,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8164,N_8167,N_8168,N_8169,N_8170,N_8174,N_8176,N_8177,N_8179,N_8180,N_8181,N_8182,N_8183,N_8186,N_8187,N_8190,N_8193,N_8194,N_8198,N_8200,N_8201,N_8203,N_8206,N_8207,N_8208,N_8210,N_8211,N_8212,N_8216,N_8217,N_8218,N_8219,N_8222,N_8223,N_8227,N_8229,N_8230,N_8232,N_8233,N_8234,N_8235,N_8237,N_8238,N_8240,N_8241,N_8242,N_8244,N_8246,N_8247,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8257,N_8260,N_8261,N_8262,N_8265,N_8266,N_8268,N_8269,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8287,N_8288,N_8290,N_8291,N_8292,N_8295,N_8298,N_8300,N_8301,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8311,N_8312,N_8313,N_8315,N_8317,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8328,N_8331,N_8334,N_8336,N_8337,N_8338,N_8342,N_8345,N_8346,N_8348,N_8350,N_8351,N_8352,N_8354,N_8356,N_8357,N_8359,N_8360,N_8361,N_8362,N_8364,N_8365,N_8367,N_8368,N_8370,N_8371,N_8373,N_8374,N_8375,N_8377,N_8379,N_8380,N_8382,N_8384,N_8385,N_8387,N_8389,N_8390,N_8393,N_8395,N_8396,N_8397,N_8398,N_8401,N_8402,N_8403,N_8404,N_8407,N_8408,N_8409,N_8410,N_8411,N_8413,N_8414,N_8415,N_8416,N_8418,N_8419,N_8421,N_8422,N_8423,N_8425,N_8426,N_8429,N_8431,N_8432,N_8433,N_8434,N_8435,N_8437,N_8438,N_8441,N_8442,N_8443,N_8444,N_8445,N_8447,N_8450,N_8452,N_8457,N_8458,N_8459,N_8460,N_8462,N_8464,N_8465,N_8466,N_8468,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8486,N_8487,N_8488,N_8492,N_8496,N_8497,N_8498,N_8499,N_8503,N_8504,N_8505,N_8508,N_8510,N_8511,N_8512,N_8513,N_8515,N_8518,N_8519,N_8522,N_8524,N_8525,N_8526,N_8529,N_8533,N_8534,N_8536,N_8539,N_8541,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8552,N_8553,N_8554,N_8555,N_8558,N_8559,N_8560,N_8562,N_8564,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8576,N_8580,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8595,N_8596,N_8597,N_8599,N_8600,N_8602,N_8603,N_8605,N_8607,N_8608,N_8609,N_8610,N_8612,N_8617,N_8619,N_8620,N_8621,N_8622,N_8623,N_8625,N_8626,N_8629,N_8631,N_8632,N_8634,N_8635,N_8637,N_8638,N_8640,N_8641,N_8643,N_8644,N_8645,N_8646,N_8647,N_8650,N_8653,N_8655,N_8656,N_8658,N_8660,N_8661,N_8662,N_8663,N_8666,N_8667,N_8668,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8681,N_8682,N_8685,N_8686,N_8687,N_8688,N_8690,N_8691,N_8694,N_8697,N_8698,N_8700,N_8701,N_8703,N_8704,N_8705,N_8706,N_8707,N_8711,N_8712,N_8715,N_8716,N_8717,N_8719,N_8720,N_8721,N_8723,N_8724,N_8725,N_8726,N_8729,N_8732,N_8733,N_8734,N_8735,N_8736,N_8738,N_8740,N_8744,N_8745,N_8746,N_8748,N_8749,N_8751,N_8752,N_8753,N_8754,N_8759,N_8760,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8769,N_8771,N_8773,N_8774,N_8776,N_8777,N_8778,N_8780,N_8781,N_8783,N_8787,N_8788,N_8790,N_8791,N_8792,N_8793,N_8795,N_8796,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8806,N_8808,N_8809,N_8810,N_8812,N_8813,N_8815,N_8817,N_8818,N_8819,N_8820,N_8821,N_8827,N_8828,N_8829,N_8830,N_8831,N_8833,N_8835,N_8838,N_8840,N_8841,N_8843,N_8844,N_8847,N_8848,N_8850,N_8851,N_8853,N_8854,N_8855,N_8857,N_8858,N_8861,N_8866,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8891,N_8892,N_8893,N_8894,N_8896,N_8897,N_8899,N_8901,N_8902,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8923,N_8924,N_8929,N_8930,N_8932,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8944,N_8945,N_8947,N_8948,N_8951,N_8952,N_8953,N_8954,N_8955,N_8957,N_8959,N_8960,N_8961,N_8962,N_8964,N_8970,N_8971,N_8972,N_8975,N_8978,N_8979,N_8982,N_8984,N_8985,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8995,N_8996,N_8997,N_8998,N_9000,N_9004,N_9005,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9021,N_9022,N_9023,N_9025,N_9026,N_9027,N_9028,N_9030,N_9034,N_9038,N_9039,N_9040,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9052,N_9053,N_9054,N_9055,N_9057,N_9058,N_9059,N_9061,N_9062,N_9063,N_9064,N_9065,N_9067,N_9068,N_9069,N_9071,N_9072,N_9076,N_9078,N_9080,N_9082,N_9084,N_9087,N_9090,N_9091,N_9097,N_9098,N_9099,N_9101,N_9102,N_9103,N_9104,N_9107,N_9109,N_9110,N_9111,N_9112,N_9114,N_9116,N_9118,N_9121,N_9123,N_9124,N_9125,N_9129,N_9130,N_9133,N_9135,N_9136,N_9137,N_9138,N_9139,N_9141,N_9143,N_9144,N_9146,N_9147,N_9149,N_9150,N_9153,N_9155,N_9156,N_9161,N_9162,N_9163,N_9164,N_9169,N_9170,N_9171,N_9173,N_9177,N_9179,N_9181,N_9182,N_9183,N_9184,N_9188,N_9189,N_9190,N_9193,N_9195,N_9196,N_9199,N_9202,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9230,N_9231,N_9232,N_9234,N_9236,N_9239,N_9241,N_9242,N_9244,N_9245,N_9246,N_9250,N_9251,N_9252,N_9255,N_9256,N_9257,N_9258,N_9262,N_9263,N_9269,N_9270,N_9271,N_9274,N_9275,N_9278,N_9280,N_9281,N_9282,N_9286,N_9287,N_9288,N_9290,N_9291,N_9294,N_9295,N_9298,N_9300,N_9301,N_9303,N_9305,N_9306,N_9307,N_9310,N_9311,N_9314,N_9315,N_9316,N_9323,N_9325,N_9326,N_9327,N_9328,N_9330,N_9337,N_9338,N_9339,N_9340,N_9342,N_9343,N_9346,N_9347,N_9348,N_9351,N_9352,N_9354,N_9355,N_9356,N_9358,N_9359,N_9360,N_9361,N_9366,N_9367,N_9368,N_9370,N_9371,N_9374,N_9375,N_9381,N_9382,N_9383,N_9385,N_9386,N_9388,N_9389,N_9390,N_9392,N_9395,N_9396,N_9398,N_9399,N_9400,N_9401,N_9404,N_9405,N_9406,N_9407,N_9411,N_9413,N_9414,N_9415,N_9418,N_9420,N_9421,N_9422,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9431,N_9432,N_9433,N_9434,N_9436,N_9438,N_9439,N_9440,N_9441,N_9442,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9454,N_9455,N_9460,N_9461,N_9463,N_9466,N_9467,N_9470,N_9472,N_9474,N_9475,N_9477,N_9478,N_9481,N_9482,N_9483,N_9484,N_9486,N_9488,N_9489,N_9490,N_9493,N_9496,N_9497,N_9499,N_9500,N_9501,N_9502,N_9503,N_9505,N_9506,N_9511,N_9512,N_9513,N_9514,N_9515,N_9517,N_9518,N_9520,N_9523,N_9525,N_9528,N_9529,N_9532,N_9534,N_9535,N_9537,N_9540,N_9541,N_9546,N_9547,N_9548,N_9553,N_9554,N_9555,N_9556,N_9557,N_9559,N_9564,N_9566,N_9568,N_9569,N_9570,N_9571,N_9573,N_9576,N_9577,N_9578,N_9580,N_9581,N_9584,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9597,N_9599,N_9606,N_9608,N_9610,N_9611,N_9612,N_9613,N_9615,N_9616,N_9617,N_9619,N_9620,N_9622,N_9623,N_9624,N_9627,N_9628,N_9630,N_9633,N_9634,N_9636,N_9640,N_9641,N_9645,N_9646,N_9647,N_9649,N_9650,N_9652,N_9654,N_9657,N_9658,N_9659,N_9661,N_9663,N_9664,N_9667,N_9669,N_9670,N_9671,N_9674,N_9675,N_9676,N_9679,N_9682,N_9683,N_9686,N_9689,N_9690,N_9691,N_9693,N_9694,N_9695,N_9696,N_9697,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9709,N_9711,N_9712,N_9714,N_9716,N_9717,N_9718,N_9719,N_9721,N_9722,N_9723,N_9724,N_9725,N_9728,N_9730,N_9731,N_9732,N_9733,N_9734,N_9737,N_9738,N_9739,N_9740,N_9742,N_9743,N_9744,N_9747,N_9749,N_9751,N_9754,N_9757,N_9758,N_9759,N_9762,N_9763,N_9765,N_9768,N_9771,N_9772,N_9777,N_9778,N_9782,N_9785,N_9787,N_9788,N_9789,N_9790,N_9791,N_9793,N_9794,N_9796,N_9797,N_9798,N_9799,N_9801,N_9802,N_9806,N_9807,N_9808,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9823,N_9824,N_9826,N_9828,N_9829,N_9831,N_9834,N_9835,N_9837,N_9838,N_9839,N_9840,N_9841,N_9843,N_9844,N_9846,N_9847,N_9855,N_9856,N_9858,N_9860,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9888,N_9889,N_9892,N_9893,N_9895,N_9899,N_9900,N_9901,N_9903,N_9904,N_9905,N_9906,N_9908,N_9909,N_9911,N_9912,N_9915,N_9920,N_9921,N_9923,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9936,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9948,N_9950,N_9953,N_9954,N_9955,N_9958,N_9960,N_9961,N_9962,N_9964,N_9966,N_9970,N_9971,N_9974,N_9975,N_9977,N_9978,N_9981,N_9982,N_9983,N_9984,N_9987,N_9988,N_9989,N_9990,N_9991,N_9993,N_9995,N_9996,N_9998;
nor U0 (N_0,In_79,In_573);
and U1 (N_1,In_647,In_248);
nand U2 (N_2,In_178,In_36);
nand U3 (N_3,In_147,In_761);
nand U4 (N_4,In_87,In_665);
or U5 (N_5,In_332,In_957);
nor U6 (N_6,In_841,In_414);
and U7 (N_7,In_779,In_659);
and U8 (N_8,In_730,In_759);
or U9 (N_9,In_556,In_297);
or U10 (N_10,In_815,In_716);
and U11 (N_11,In_662,In_588);
or U12 (N_12,In_905,In_866);
and U13 (N_13,In_572,In_903);
nand U14 (N_14,In_997,In_243);
or U15 (N_15,In_3,In_879);
or U16 (N_16,In_485,In_198);
and U17 (N_17,In_606,In_436);
and U18 (N_18,In_531,In_520);
xor U19 (N_19,In_634,In_907);
nor U20 (N_20,In_686,In_702);
and U21 (N_21,In_868,In_182);
nor U22 (N_22,In_404,In_549);
nand U23 (N_23,In_145,In_741);
or U24 (N_24,In_77,In_101);
nor U25 (N_25,In_352,In_464);
and U26 (N_26,In_177,In_839);
nor U27 (N_27,In_433,In_583);
nand U28 (N_28,In_319,In_60);
nor U29 (N_29,In_74,In_943);
and U30 (N_30,In_481,In_607);
nor U31 (N_31,In_442,In_134);
and U32 (N_32,In_722,In_2);
or U33 (N_33,In_401,In_886);
or U34 (N_34,In_751,In_26);
nand U35 (N_35,In_110,In_192);
or U36 (N_36,In_174,In_435);
or U37 (N_37,In_407,In_270);
or U38 (N_38,In_652,In_561);
nor U39 (N_39,In_463,In_493);
and U40 (N_40,In_942,In_438);
or U41 (N_41,In_962,In_776);
xor U42 (N_42,In_506,In_940);
nand U43 (N_43,In_16,In_94);
xnor U44 (N_44,In_714,In_91);
nor U45 (N_45,In_509,In_15);
or U46 (N_46,In_650,In_807);
or U47 (N_47,In_181,In_837);
and U48 (N_48,In_928,In_673);
nor U49 (N_49,In_496,In_451);
or U50 (N_50,In_428,In_602);
and U51 (N_51,In_141,In_275);
nand U52 (N_52,In_516,In_191);
or U53 (N_53,In_582,In_971);
and U54 (N_54,In_621,In_551);
nor U55 (N_55,In_14,In_850);
or U56 (N_56,In_322,In_142);
and U57 (N_57,In_990,In_859);
nand U58 (N_58,In_711,In_749);
nor U59 (N_59,In_432,In_977);
or U60 (N_60,In_107,In_276);
nor U61 (N_61,In_236,In_614);
and U62 (N_62,In_186,In_871);
nand U63 (N_63,In_73,In_635);
and U64 (N_64,In_362,In_338);
and U65 (N_65,In_378,In_326);
or U66 (N_66,In_165,In_295);
or U67 (N_67,In_750,In_799);
and U68 (N_68,In_458,In_330);
xor U69 (N_69,In_305,In_980);
nand U70 (N_70,In_114,In_265);
and U71 (N_71,In_241,In_152);
or U72 (N_72,In_511,In_706);
nand U73 (N_73,In_715,In_22);
nor U74 (N_74,In_434,In_589);
nor U75 (N_75,In_400,In_742);
and U76 (N_76,In_317,In_563);
and U77 (N_77,In_160,In_535);
nor U78 (N_78,In_448,In_425);
nand U79 (N_79,In_772,In_704);
nor U80 (N_80,In_254,In_224);
and U81 (N_81,In_227,In_244);
or U82 (N_82,In_136,In_757);
nand U83 (N_83,In_45,In_479);
nor U84 (N_84,In_916,In_854);
or U85 (N_85,In_365,In_929);
nand U86 (N_86,In_67,In_148);
or U87 (N_87,In_84,In_180);
nor U88 (N_88,In_575,In_238);
nor U89 (N_89,In_791,In_974);
or U90 (N_90,In_351,In_814);
xnor U91 (N_91,In_620,In_695);
nor U92 (N_92,In_987,In_825);
nor U93 (N_93,In_623,In_83);
or U94 (N_94,In_547,In_294);
and U95 (N_95,In_112,In_934);
and U96 (N_96,In_840,In_342);
nand U97 (N_97,In_113,In_482);
xor U98 (N_98,In_334,In_590);
or U99 (N_99,In_372,In_768);
nand U100 (N_100,In_693,In_760);
or U101 (N_101,In_392,In_851);
and U102 (N_102,In_369,In_405);
xor U103 (N_103,In_502,In_116);
xnor U104 (N_104,In_619,In_975);
or U105 (N_105,In_890,In_259);
or U106 (N_106,In_288,In_228);
nand U107 (N_107,In_813,In_444);
nor U108 (N_108,In_808,In_472);
nand U109 (N_109,In_368,In_798);
nand U110 (N_110,In_431,In_568);
or U111 (N_111,In_40,In_735);
and U112 (N_112,In_324,In_403);
or U113 (N_113,In_230,In_34);
or U114 (N_114,In_52,In_654);
nor U115 (N_115,In_9,In_416);
nor U116 (N_116,In_505,In_501);
nand U117 (N_117,In_770,In_430);
and U118 (N_118,In_835,In_663);
nor U119 (N_119,In_781,In_7);
and U120 (N_120,In_225,In_679);
or U121 (N_121,In_950,In_47);
or U122 (N_122,In_540,In_98);
and U123 (N_123,In_27,In_769);
nor U124 (N_124,In_832,In_486);
nand U125 (N_125,In_63,In_255);
and U126 (N_126,In_353,In_137);
nor U127 (N_127,In_705,In_930);
or U128 (N_128,In_529,In_700);
nand U129 (N_129,In_775,In_193);
and U130 (N_130,In_144,In_592);
nand U131 (N_131,In_262,In_264);
nor U132 (N_132,In_133,In_280);
nand U133 (N_133,In_565,In_553);
nor U134 (N_134,In_956,In_739);
nand U135 (N_135,In_649,In_300);
or U136 (N_136,In_628,In_961);
nor U137 (N_137,In_97,In_901);
and U138 (N_138,In_530,In_536);
xnor U139 (N_139,In_398,In_158);
nor U140 (N_140,In_782,In_544);
nor U141 (N_141,In_828,In_963);
xor U142 (N_142,In_666,In_691);
xor U143 (N_143,In_201,In_797);
and U144 (N_144,In_682,In_44);
xor U145 (N_145,In_829,In_252);
nand U146 (N_146,In_972,In_296);
nor U147 (N_147,In_357,In_889);
nand U148 (N_148,In_584,In_811);
and U149 (N_149,In_371,In_450);
nand U150 (N_150,In_261,In_989);
or U151 (N_151,In_0,In_422);
nor U152 (N_152,In_690,In_877);
and U153 (N_153,In_429,In_893);
and U154 (N_154,In_370,In_75);
nand U155 (N_155,In_955,In_587);
or U156 (N_156,In_123,In_688);
or U157 (N_157,In_944,In_102);
nor U158 (N_158,In_612,In_643);
nor U159 (N_159,In_12,In_914);
nor U160 (N_160,In_564,In_831);
or U161 (N_161,In_591,In_793);
and U162 (N_162,In_172,In_289);
or U163 (N_163,In_211,In_683);
and U164 (N_164,In_862,In_718);
nor U165 (N_165,In_385,In_30);
nor U166 (N_166,In_473,In_888);
xor U167 (N_167,In_569,In_249);
and U168 (N_168,In_267,In_637);
and U169 (N_169,In_38,In_53);
xor U170 (N_170,In_915,In_651);
nor U171 (N_171,In_131,In_363);
nor U172 (N_172,In_155,In_283);
nor U173 (N_173,In_597,In_394);
nand U174 (N_174,In_106,In_303);
and U175 (N_175,In_272,In_696);
and U176 (N_176,In_812,In_323);
nand U177 (N_177,In_59,In_755);
nand U178 (N_178,In_870,In_164);
nand U179 (N_179,In_747,In_245);
or U180 (N_180,In_157,In_684);
nand U181 (N_181,In_388,In_848);
nor U182 (N_182,In_894,In_806);
nor U183 (N_183,In_256,In_156);
and U184 (N_184,In_846,In_960);
xnor U185 (N_185,In_550,In_393);
xnor U186 (N_186,In_910,In_132);
nor U187 (N_187,In_636,In_909);
or U188 (N_188,In_885,In_209);
nand U189 (N_189,In_118,In_308);
nor U190 (N_190,In_525,In_912);
or U191 (N_191,In_574,In_949);
and U192 (N_192,In_347,In_500);
nand U193 (N_193,In_250,In_712);
nor U194 (N_194,In_869,In_864);
or U195 (N_195,In_337,In_139);
and U196 (N_196,In_884,In_946);
and U197 (N_197,In_170,In_390);
nor U198 (N_198,In_710,In_307);
nor U199 (N_199,In_838,In_701);
xnor U200 (N_200,In_65,In_984);
or U201 (N_201,In_95,In_456);
nor U202 (N_202,In_212,In_459);
and U203 (N_203,In_736,In_924);
nand U204 (N_204,In_281,In_21);
nand U205 (N_205,In_268,In_465);
or U206 (N_206,In_253,In_821);
or U207 (N_207,In_855,In_534);
nor U208 (N_208,In_743,In_247);
or U209 (N_209,In_477,In_969);
or U210 (N_210,In_801,In_674);
nor U211 (N_211,In_417,In_626);
nor U212 (N_212,In_50,In_301);
or U213 (N_213,In_143,In_660);
xor U214 (N_214,In_271,In_35);
and U215 (N_215,In_708,In_533);
or U216 (N_216,In_827,In_366);
and U217 (N_217,In_555,In_891);
and U218 (N_218,In_518,In_542);
nor U219 (N_219,In_787,In_727);
nor U220 (N_220,In_108,In_777);
nor U221 (N_221,In_687,In_642);
xnor U222 (N_222,In_33,In_489);
and U223 (N_223,In_847,In_154);
nand U224 (N_224,In_599,In_938);
nand U225 (N_225,In_6,In_251);
or U226 (N_226,In_354,In_935);
or U227 (N_227,In_724,In_911);
xor U228 (N_228,In_291,In_857);
nor U229 (N_229,In_125,In_965);
nand U230 (N_230,In_664,In_558);
or U231 (N_231,In_183,In_699);
or U232 (N_232,In_382,In_188);
and U233 (N_233,In_217,In_629);
xor U234 (N_234,In_122,In_964);
and U235 (N_235,In_532,In_348);
or U236 (N_236,In_420,In_339);
nand U237 (N_237,In_557,In_878);
and U238 (N_238,In_552,In_215);
nor U239 (N_239,In_723,In_316);
or U240 (N_240,In_677,In_875);
nor U241 (N_241,In_277,In_387);
and U242 (N_242,In_852,In_640);
nor U243 (N_243,In_460,In_795);
and U244 (N_244,In_293,In_99);
nand U245 (N_245,In_344,In_287);
and U246 (N_246,In_207,In_395);
nand U247 (N_247,In_610,In_282);
and U248 (N_248,In_580,In_883);
or U249 (N_249,In_865,In_653);
and U250 (N_250,In_467,In_421);
or U251 (N_251,In_773,In_469);
xor U252 (N_252,In_483,In_921);
nand U253 (N_253,In_466,In_161);
nand U254 (N_254,In_830,In_672);
nor U255 (N_255,In_983,In_406);
nor U256 (N_256,In_546,In_680);
or U257 (N_257,In_982,In_31);
and U258 (N_258,In_601,In_266);
xnor U259 (N_259,In_927,In_25);
nand U260 (N_260,In_290,In_794);
or U261 (N_261,In_763,In_833);
nand U262 (N_262,In_457,In_853);
nand U263 (N_263,In_570,In_689);
nor U264 (N_264,In_976,In_163);
nor U265 (N_265,In_487,In_340);
nor U266 (N_266,In_758,In_816);
xor U267 (N_267,In_882,In_692);
and U268 (N_268,In_948,In_678);
nand U269 (N_269,In_917,In_605);
nor U270 (N_270,In_461,In_96);
xnor U271 (N_271,In_80,In_167);
nor U272 (N_272,In_311,In_1);
and U273 (N_273,In_202,In_159);
and U274 (N_274,In_81,In_959);
or U275 (N_275,In_146,In_299);
nor U276 (N_276,In_383,In_185);
nor U277 (N_277,In_541,In_203);
and U278 (N_278,In_992,In_970);
or U279 (N_279,In_545,In_127);
xor U280 (N_280,In_190,In_717);
or U281 (N_281,In_800,In_576);
and U282 (N_282,In_11,In_503);
or U283 (N_283,In_756,In_56);
nor U284 (N_284,In_313,In_269);
nand U285 (N_285,In_64,In_667);
nor U286 (N_286,In_104,In_5);
nor U287 (N_287,In_764,In_908);
nand U288 (N_288,In_967,In_343);
nand U289 (N_289,In_941,In_517);
and U290 (N_290,In_548,In_455);
and U291 (N_291,In_918,In_426);
or U292 (N_292,In_728,In_103);
xor U293 (N_293,In_611,In_199);
nor U294 (N_294,In_376,In_904);
nor U295 (N_295,In_792,In_805);
or U296 (N_296,In_658,In_887);
and U297 (N_297,In_115,In_998);
nand U298 (N_298,In_876,In_778);
or U299 (N_299,In_899,In_803);
or U300 (N_300,In_604,In_449);
and U301 (N_301,In_58,In_958);
or U302 (N_302,In_86,In_415);
and U303 (N_303,In_937,In_246);
or U304 (N_304,In_790,In_669);
or U305 (N_305,In_936,In_346);
nand U306 (N_306,In_412,In_932);
or U307 (N_307,In_187,In_522);
and U308 (N_308,In_93,In_423);
nor U309 (N_309,In_150,In_630);
and U310 (N_310,In_92,In_559);
xnor U311 (N_311,In_523,In_836);
nand U312 (N_312,In_437,In_418);
nand U313 (N_313,In_396,In_632);
and U314 (N_314,In_897,In_510);
nand U315 (N_315,In_61,In_320);
or U316 (N_316,In_89,In_48);
nor U317 (N_317,In_752,In_538);
nor U318 (N_318,In_719,In_234);
and U319 (N_319,In_381,In_685);
and U320 (N_320,In_208,In_740);
or U321 (N_321,In_82,In_8);
or U322 (N_322,In_386,In_856);
and U323 (N_323,In_298,In_923);
and U324 (N_324,In_492,In_384);
and U325 (N_325,In_738,In_46);
xor U326 (N_326,In_767,In_454);
nand U327 (N_327,In_746,In_744);
nand U328 (N_328,In_774,In_765);
and U329 (N_329,In_179,In_41);
or U330 (N_330,In_737,In_223);
and U331 (N_331,In_325,In_615);
and U332 (N_332,In_100,In_397);
nor U333 (N_333,In_951,In_895);
nand U334 (N_334,In_861,In_515);
xnor U335 (N_335,In_784,In_278);
nand U336 (N_336,In_913,In_221);
nand U337 (N_337,In_579,In_845);
nor U338 (N_338,In_600,In_72);
and U339 (N_339,In_419,In_257);
nand U340 (N_340,In_443,In_993);
and U341 (N_341,In_766,In_844);
and U342 (N_342,In_577,In_306);
and U343 (N_343,In_153,In_76);
nor U344 (N_344,In_554,In_631);
nor U345 (N_345,In_51,In_978);
and U346 (N_346,In_641,In_315);
nor U347 (N_347,In_380,In_843);
and U348 (N_348,In_860,In_117);
xor U349 (N_349,In_947,In_232);
nand U350 (N_350,In_331,In_90);
xor U351 (N_351,In_166,In_349);
or U352 (N_352,In_994,In_732);
nand U353 (N_353,In_18,In_988);
nand U354 (N_354,In_440,In_124);
nand U355 (N_355,In_820,In_312);
nand U356 (N_356,In_661,In_931);
and U357 (N_357,In_648,In_786);
or U358 (N_358,In_213,In_594);
and U359 (N_359,In_129,In_804);
nor U360 (N_360,In_603,In_194);
or U361 (N_361,In_881,In_608);
or U362 (N_362,In_411,In_952);
and U363 (N_363,In_379,In_66);
or U364 (N_364,In_586,In_214);
and U365 (N_365,In_328,In_788);
or U366 (N_366,In_309,In_70);
nand U367 (N_367,In_20,In_189);
and U368 (N_368,In_646,In_668);
nor U369 (N_369,In_655,In_842);
nor U370 (N_370,In_85,In_409);
and U371 (N_371,In_709,In_196);
nor U372 (N_372,In_355,In_476);
xnor U373 (N_373,In_622,In_240);
xnor U374 (N_374,In_771,In_336);
or U375 (N_375,In_880,In_242);
or U376 (N_376,In_900,In_32);
nor U377 (N_377,In_762,In_413);
nor U378 (N_378,In_780,In_210);
nor U379 (N_379,In_519,In_367);
and U380 (N_380,In_19,In_996);
nor U381 (N_381,In_57,In_452);
and U382 (N_382,In_17,In_872);
nor U383 (N_383,In_273,In_206);
and U384 (N_384,In_488,In_274);
or U385 (N_385,In_925,In_617);
or U386 (N_386,In_302,In_218);
or U387 (N_387,In_314,In_447);
or U388 (N_388,In_609,In_720);
nor U389 (N_389,In_135,In_318);
nand U390 (N_390,In_151,In_873);
or U391 (N_391,In_625,In_478);
nor U392 (N_392,In_919,In_898);
or U393 (N_393,In_480,In_475);
and U394 (N_394,In_356,In_507);
nand U395 (N_395,In_239,In_991);
and U396 (N_396,In_979,In_537);
nor U397 (N_397,In_494,In_754);
nand U398 (N_398,In_729,In_13);
and U399 (N_399,In_810,In_902);
and U400 (N_400,In_593,In_24);
nand U401 (N_401,In_205,In_725);
xor U402 (N_402,In_68,In_424);
or U403 (N_403,In_618,In_162);
and U404 (N_404,In_399,In_231);
nand U405 (N_405,In_524,In_539);
or U406 (N_406,In_470,In_310);
or U407 (N_407,In_327,In_638);
nand U408 (N_408,In_578,In_62);
nand U409 (N_409,In_981,In_748);
nor U410 (N_410,In_138,In_233);
nand U411 (N_411,In_945,In_200);
nor U412 (N_412,In_490,In_671);
xnor U413 (N_413,In_999,In_826);
or U414 (N_414,In_703,In_817);
and U415 (N_415,In_130,In_627);
nand U416 (N_416,In_235,In_676);
nand U417 (N_417,In_220,In_364);
and U418 (N_418,In_834,In_284);
nor U419 (N_419,In_391,In_49);
and U420 (N_420,In_954,In_818);
nand U421 (N_421,In_468,In_4);
or U422 (N_422,In_514,In_802);
nor U423 (N_423,In_119,In_721);
nand U424 (N_424,In_42,In_140);
nand U425 (N_425,In_939,In_726);
and U426 (N_426,In_731,In_995);
nand U427 (N_427,In_78,In_521);
nor U428 (N_428,In_528,In_69);
or U429 (N_429,In_508,In_753);
nor U430 (N_430,In_10,In_581);
nand U431 (N_431,In_849,In_335);
and U432 (N_432,In_585,In_734);
nand U433 (N_433,In_29,In_675);
nand U434 (N_434,In_410,In_341);
nor U435 (N_435,In_526,In_527);
nor U436 (N_436,In_920,In_613);
or U437 (N_437,In_986,In_789);
nor U438 (N_438,In_350,In_896);
nor U439 (N_439,In_906,In_513);
nand U440 (N_440,In_120,In_567);
and U441 (N_441,In_785,In_169);
or U442 (N_442,In_43,In_474);
nor U443 (N_443,In_111,In_745);
nand U444 (N_444,In_560,In_497);
nand U445 (N_445,In_633,In_656);
nor U446 (N_446,In_624,In_263);
or U447 (N_447,In_329,In_175);
xor U448 (N_448,In_858,In_204);
and U449 (N_449,In_373,In_408);
and U450 (N_450,In_926,In_23);
and U451 (N_451,In_616,In_359);
nor U452 (N_452,In_427,In_953);
or U453 (N_453,In_462,In_377);
nand U454 (N_454,In_698,In_237);
and U455 (N_455,In_445,In_543);
nand U456 (N_456,In_260,In_197);
and U457 (N_457,In_39,In_292);
nor U458 (N_458,In_176,In_491);
or U459 (N_459,In_446,In_985);
nor U460 (N_460,In_598,In_596);
nand U461 (N_461,In_226,In_304);
and U462 (N_462,In_863,In_571);
nand U463 (N_463,In_402,In_657);
nor U464 (N_464,In_819,In_933);
xnor U465 (N_465,In_874,In_713);
and U466 (N_466,In_822,In_173);
nor U467 (N_467,In_258,In_55);
nand U468 (N_468,In_498,In_219);
nand U469 (N_469,In_71,In_639);
or U470 (N_470,In_149,In_361);
xnor U471 (N_471,In_279,In_286);
nand U472 (N_472,In_88,In_922);
nor U473 (N_473,In_441,In_184);
xor U474 (N_474,In_109,In_499);
nand U475 (N_475,In_973,In_809);
nand U476 (N_476,In_229,In_823);
or U477 (N_477,In_453,In_681);
nand U478 (N_478,In_966,In_168);
and U479 (N_479,In_694,In_216);
and U480 (N_480,In_562,In_195);
nor U481 (N_481,In_471,In_644);
nand U482 (N_482,In_796,In_867);
nand U483 (N_483,In_824,In_439);
or U484 (N_484,In_566,In_892);
nand U485 (N_485,In_54,In_389);
or U486 (N_486,In_171,In_285);
nand U487 (N_487,In_121,In_783);
or U488 (N_488,In_321,In_670);
nand U489 (N_489,In_595,In_37);
nor U490 (N_490,In_375,In_222);
nor U491 (N_491,In_360,In_495);
nor U492 (N_492,In_733,In_645);
xor U493 (N_493,In_697,In_707);
or U494 (N_494,In_128,In_374);
and U495 (N_495,In_345,In_358);
xnor U496 (N_496,In_105,In_504);
and U497 (N_497,In_126,In_28);
and U498 (N_498,In_512,In_968);
xnor U499 (N_499,In_333,In_484);
nand U500 (N_500,In_579,In_93);
or U501 (N_501,In_64,In_651);
nand U502 (N_502,In_588,In_856);
nor U503 (N_503,In_816,In_99);
nand U504 (N_504,In_286,In_702);
and U505 (N_505,In_380,In_426);
nand U506 (N_506,In_510,In_831);
nand U507 (N_507,In_634,In_921);
nand U508 (N_508,In_790,In_542);
nand U509 (N_509,In_753,In_14);
or U510 (N_510,In_913,In_435);
or U511 (N_511,In_126,In_102);
or U512 (N_512,In_457,In_152);
and U513 (N_513,In_504,In_985);
nand U514 (N_514,In_36,In_971);
and U515 (N_515,In_130,In_584);
xor U516 (N_516,In_93,In_919);
and U517 (N_517,In_5,In_389);
nand U518 (N_518,In_168,In_58);
nand U519 (N_519,In_982,In_405);
nand U520 (N_520,In_627,In_32);
nor U521 (N_521,In_983,In_716);
xor U522 (N_522,In_940,In_532);
and U523 (N_523,In_609,In_269);
nand U524 (N_524,In_715,In_352);
or U525 (N_525,In_775,In_346);
or U526 (N_526,In_36,In_828);
and U527 (N_527,In_77,In_697);
nor U528 (N_528,In_772,In_970);
and U529 (N_529,In_818,In_59);
xor U530 (N_530,In_419,In_137);
and U531 (N_531,In_863,In_264);
and U532 (N_532,In_784,In_905);
nor U533 (N_533,In_116,In_615);
or U534 (N_534,In_790,In_370);
or U535 (N_535,In_420,In_535);
or U536 (N_536,In_733,In_22);
nor U537 (N_537,In_530,In_989);
or U538 (N_538,In_316,In_979);
or U539 (N_539,In_38,In_947);
nor U540 (N_540,In_822,In_824);
or U541 (N_541,In_904,In_285);
nand U542 (N_542,In_353,In_426);
nand U543 (N_543,In_271,In_149);
nor U544 (N_544,In_552,In_789);
xnor U545 (N_545,In_280,In_713);
nor U546 (N_546,In_493,In_22);
and U547 (N_547,In_473,In_425);
nand U548 (N_548,In_210,In_428);
or U549 (N_549,In_428,In_368);
nor U550 (N_550,In_695,In_164);
nand U551 (N_551,In_518,In_583);
nor U552 (N_552,In_821,In_171);
nor U553 (N_553,In_506,In_665);
and U554 (N_554,In_425,In_140);
nand U555 (N_555,In_636,In_139);
and U556 (N_556,In_398,In_466);
and U557 (N_557,In_836,In_635);
nand U558 (N_558,In_886,In_451);
and U559 (N_559,In_170,In_426);
nand U560 (N_560,In_821,In_720);
nand U561 (N_561,In_259,In_601);
or U562 (N_562,In_722,In_761);
nand U563 (N_563,In_940,In_15);
and U564 (N_564,In_80,In_808);
nand U565 (N_565,In_829,In_513);
or U566 (N_566,In_369,In_793);
nand U567 (N_567,In_75,In_803);
nand U568 (N_568,In_574,In_903);
xnor U569 (N_569,In_685,In_833);
or U570 (N_570,In_720,In_429);
nand U571 (N_571,In_916,In_70);
nor U572 (N_572,In_742,In_893);
or U573 (N_573,In_94,In_342);
nand U574 (N_574,In_307,In_321);
xor U575 (N_575,In_320,In_453);
nor U576 (N_576,In_952,In_878);
nand U577 (N_577,In_389,In_440);
and U578 (N_578,In_548,In_332);
and U579 (N_579,In_681,In_4);
nand U580 (N_580,In_50,In_306);
nand U581 (N_581,In_216,In_645);
nor U582 (N_582,In_939,In_972);
nand U583 (N_583,In_447,In_841);
or U584 (N_584,In_786,In_304);
and U585 (N_585,In_295,In_585);
or U586 (N_586,In_830,In_719);
nand U587 (N_587,In_198,In_850);
nor U588 (N_588,In_886,In_153);
and U589 (N_589,In_747,In_255);
nand U590 (N_590,In_108,In_99);
nor U591 (N_591,In_508,In_778);
nand U592 (N_592,In_444,In_906);
xor U593 (N_593,In_211,In_154);
or U594 (N_594,In_215,In_406);
nor U595 (N_595,In_239,In_175);
xor U596 (N_596,In_393,In_955);
xnor U597 (N_597,In_340,In_581);
nor U598 (N_598,In_242,In_902);
nand U599 (N_599,In_454,In_259);
nand U600 (N_600,In_335,In_733);
nand U601 (N_601,In_896,In_726);
or U602 (N_602,In_55,In_487);
nand U603 (N_603,In_842,In_897);
nor U604 (N_604,In_332,In_403);
or U605 (N_605,In_411,In_793);
and U606 (N_606,In_983,In_110);
nor U607 (N_607,In_715,In_707);
and U608 (N_608,In_144,In_261);
nor U609 (N_609,In_986,In_232);
and U610 (N_610,In_702,In_929);
xor U611 (N_611,In_176,In_108);
nor U612 (N_612,In_155,In_106);
xnor U613 (N_613,In_224,In_514);
or U614 (N_614,In_52,In_892);
or U615 (N_615,In_357,In_45);
xnor U616 (N_616,In_671,In_113);
and U617 (N_617,In_492,In_316);
nand U618 (N_618,In_652,In_700);
nand U619 (N_619,In_579,In_216);
nor U620 (N_620,In_777,In_994);
nand U621 (N_621,In_235,In_425);
and U622 (N_622,In_15,In_320);
nor U623 (N_623,In_611,In_366);
or U624 (N_624,In_171,In_691);
nor U625 (N_625,In_473,In_468);
and U626 (N_626,In_152,In_23);
nor U627 (N_627,In_986,In_971);
or U628 (N_628,In_915,In_164);
nand U629 (N_629,In_141,In_123);
nor U630 (N_630,In_47,In_576);
and U631 (N_631,In_856,In_65);
or U632 (N_632,In_715,In_740);
or U633 (N_633,In_617,In_436);
nor U634 (N_634,In_332,In_922);
xor U635 (N_635,In_145,In_350);
and U636 (N_636,In_733,In_135);
nor U637 (N_637,In_624,In_319);
and U638 (N_638,In_670,In_661);
nand U639 (N_639,In_739,In_46);
and U640 (N_640,In_141,In_76);
nor U641 (N_641,In_251,In_707);
or U642 (N_642,In_278,In_269);
nand U643 (N_643,In_498,In_549);
nand U644 (N_644,In_407,In_700);
or U645 (N_645,In_294,In_360);
and U646 (N_646,In_871,In_792);
xnor U647 (N_647,In_170,In_887);
nor U648 (N_648,In_274,In_968);
nand U649 (N_649,In_504,In_166);
xor U650 (N_650,In_758,In_138);
xor U651 (N_651,In_138,In_964);
nor U652 (N_652,In_655,In_576);
nand U653 (N_653,In_624,In_962);
nor U654 (N_654,In_614,In_451);
nand U655 (N_655,In_711,In_853);
or U656 (N_656,In_5,In_328);
nor U657 (N_657,In_486,In_973);
or U658 (N_658,In_586,In_681);
and U659 (N_659,In_635,In_770);
nor U660 (N_660,In_504,In_242);
nor U661 (N_661,In_589,In_850);
nor U662 (N_662,In_353,In_672);
and U663 (N_663,In_895,In_304);
nand U664 (N_664,In_160,In_582);
xnor U665 (N_665,In_647,In_88);
nand U666 (N_666,In_973,In_998);
or U667 (N_667,In_837,In_846);
nand U668 (N_668,In_525,In_930);
xor U669 (N_669,In_471,In_27);
or U670 (N_670,In_449,In_334);
nand U671 (N_671,In_698,In_401);
nand U672 (N_672,In_446,In_847);
nand U673 (N_673,In_811,In_86);
xor U674 (N_674,In_189,In_994);
nor U675 (N_675,In_785,In_391);
nand U676 (N_676,In_586,In_137);
nand U677 (N_677,In_12,In_670);
nand U678 (N_678,In_880,In_804);
nand U679 (N_679,In_82,In_52);
or U680 (N_680,In_483,In_791);
or U681 (N_681,In_177,In_646);
and U682 (N_682,In_360,In_47);
or U683 (N_683,In_426,In_919);
xnor U684 (N_684,In_361,In_279);
or U685 (N_685,In_447,In_991);
and U686 (N_686,In_536,In_405);
or U687 (N_687,In_155,In_952);
and U688 (N_688,In_18,In_46);
nand U689 (N_689,In_84,In_842);
or U690 (N_690,In_513,In_987);
or U691 (N_691,In_487,In_0);
or U692 (N_692,In_121,In_210);
nor U693 (N_693,In_71,In_223);
nand U694 (N_694,In_551,In_724);
or U695 (N_695,In_601,In_83);
and U696 (N_696,In_819,In_949);
and U697 (N_697,In_42,In_530);
or U698 (N_698,In_91,In_616);
and U699 (N_699,In_154,In_321);
and U700 (N_700,In_487,In_146);
nor U701 (N_701,In_618,In_355);
or U702 (N_702,In_844,In_341);
nor U703 (N_703,In_126,In_371);
and U704 (N_704,In_455,In_995);
and U705 (N_705,In_101,In_602);
nor U706 (N_706,In_764,In_782);
nor U707 (N_707,In_402,In_172);
and U708 (N_708,In_300,In_442);
and U709 (N_709,In_386,In_348);
nand U710 (N_710,In_156,In_720);
or U711 (N_711,In_861,In_154);
and U712 (N_712,In_957,In_311);
and U713 (N_713,In_370,In_332);
nand U714 (N_714,In_958,In_719);
and U715 (N_715,In_22,In_181);
and U716 (N_716,In_914,In_871);
nand U717 (N_717,In_740,In_35);
nand U718 (N_718,In_526,In_910);
and U719 (N_719,In_232,In_10);
or U720 (N_720,In_392,In_960);
nor U721 (N_721,In_122,In_367);
or U722 (N_722,In_972,In_24);
nand U723 (N_723,In_643,In_554);
nand U724 (N_724,In_290,In_171);
nor U725 (N_725,In_240,In_555);
nand U726 (N_726,In_766,In_670);
nor U727 (N_727,In_934,In_711);
and U728 (N_728,In_592,In_565);
or U729 (N_729,In_2,In_571);
and U730 (N_730,In_790,In_204);
xnor U731 (N_731,In_902,In_317);
xor U732 (N_732,In_923,In_869);
or U733 (N_733,In_248,In_55);
and U734 (N_734,In_598,In_394);
nor U735 (N_735,In_899,In_924);
nand U736 (N_736,In_706,In_167);
or U737 (N_737,In_130,In_601);
xor U738 (N_738,In_846,In_373);
nor U739 (N_739,In_643,In_310);
xor U740 (N_740,In_165,In_588);
or U741 (N_741,In_734,In_351);
or U742 (N_742,In_23,In_826);
or U743 (N_743,In_838,In_279);
nand U744 (N_744,In_821,In_236);
nand U745 (N_745,In_415,In_807);
or U746 (N_746,In_103,In_59);
nor U747 (N_747,In_849,In_480);
nand U748 (N_748,In_747,In_373);
and U749 (N_749,In_688,In_994);
nand U750 (N_750,In_587,In_707);
or U751 (N_751,In_779,In_874);
or U752 (N_752,In_366,In_203);
nor U753 (N_753,In_729,In_601);
and U754 (N_754,In_227,In_497);
nand U755 (N_755,In_749,In_532);
nor U756 (N_756,In_107,In_22);
nor U757 (N_757,In_800,In_603);
and U758 (N_758,In_290,In_591);
nor U759 (N_759,In_574,In_790);
nor U760 (N_760,In_647,In_673);
nor U761 (N_761,In_558,In_665);
or U762 (N_762,In_102,In_922);
nor U763 (N_763,In_703,In_936);
nor U764 (N_764,In_31,In_752);
or U765 (N_765,In_492,In_827);
or U766 (N_766,In_782,In_503);
or U767 (N_767,In_361,In_1);
nor U768 (N_768,In_100,In_934);
nand U769 (N_769,In_295,In_405);
nand U770 (N_770,In_384,In_822);
and U771 (N_771,In_495,In_749);
nand U772 (N_772,In_429,In_497);
or U773 (N_773,In_904,In_458);
and U774 (N_774,In_559,In_367);
or U775 (N_775,In_565,In_316);
nor U776 (N_776,In_987,In_762);
nor U777 (N_777,In_853,In_153);
or U778 (N_778,In_848,In_398);
nand U779 (N_779,In_60,In_639);
nor U780 (N_780,In_139,In_394);
and U781 (N_781,In_610,In_782);
or U782 (N_782,In_902,In_834);
and U783 (N_783,In_995,In_815);
xnor U784 (N_784,In_127,In_347);
nand U785 (N_785,In_270,In_964);
or U786 (N_786,In_307,In_647);
nand U787 (N_787,In_373,In_269);
and U788 (N_788,In_891,In_255);
nand U789 (N_789,In_181,In_239);
nand U790 (N_790,In_314,In_38);
nor U791 (N_791,In_778,In_912);
and U792 (N_792,In_394,In_392);
nand U793 (N_793,In_895,In_25);
and U794 (N_794,In_101,In_257);
nor U795 (N_795,In_91,In_250);
or U796 (N_796,In_289,In_819);
or U797 (N_797,In_309,In_430);
or U798 (N_798,In_713,In_807);
or U799 (N_799,In_356,In_754);
nor U800 (N_800,In_849,In_85);
xnor U801 (N_801,In_770,In_725);
nand U802 (N_802,In_991,In_962);
and U803 (N_803,In_862,In_546);
nand U804 (N_804,In_356,In_729);
nor U805 (N_805,In_306,In_823);
and U806 (N_806,In_620,In_189);
or U807 (N_807,In_588,In_514);
or U808 (N_808,In_541,In_810);
or U809 (N_809,In_325,In_963);
xor U810 (N_810,In_816,In_941);
xor U811 (N_811,In_982,In_857);
xnor U812 (N_812,In_984,In_409);
nor U813 (N_813,In_608,In_853);
nor U814 (N_814,In_886,In_391);
or U815 (N_815,In_229,In_200);
nand U816 (N_816,In_793,In_209);
xor U817 (N_817,In_913,In_901);
nand U818 (N_818,In_588,In_307);
and U819 (N_819,In_431,In_992);
and U820 (N_820,In_997,In_220);
nor U821 (N_821,In_216,In_262);
xor U822 (N_822,In_705,In_675);
nor U823 (N_823,In_383,In_510);
and U824 (N_824,In_804,In_239);
nor U825 (N_825,In_955,In_605);
or U826 (N_826,In_920,In_782);
nand U827 (N_827,In_592,In_575);
and U828 (N_828,In_252,In_581);
nand U829 (N_829,In_805,In_198);
nor U830 (N_830,In_279,In_432);
or U831 (N_831,In_856,In_22);
and U832 (N_832,In_189,In_790);
nor U833 (N_833,In_782,In_453);
nor U834 (N_834,In_183,In_770);
or U835 (N_835,In_567,In_610);
nand U836 (N_836,In_353,In_503);
nor U837 (N_837,In_266,In_188);
nor U838 (N_838,In_581,In_496);
nand U839 (N_839,In_752,In_889);
and U840 (N_840,In_389,In_945);
nor U841 (N_841,In_484,In_99);
or U842 (N_842,In_534,In_10);
nor U843 (N_843,In_19,In_401);
nand U844 (N_844,In_978,In_112);
or U845 (N_845,In_585,In_757);
nand U846 (N_846,In_535,In_419);
or U847 (N_847,In_169,In_193);
nor U848 (N_848,In_726,In_931);
and U849 (N_849,In_13,In_321);
nor U850 (N_850,In_870,In_628);
nand U851 (N_851,In_259,In_295);
nand U852 (N_852,In_58,In_724);
or U853 (N_853,In_803,In_579);
or U854 (N_854,In_918,In_313);
or U855 (N_855,In_86,In_495);
and U856 (N_856,In_171,In_962);
or U857 (N_857,In_591,In_76);
nor U858 (N_858,In_824,In_18);
and U859 (N_859,In_339,In_209);
xor U860 (N_860,In_696,In_200);
nor U861 (N_861,In_680,In_561);
nand U862 (N_862,In_350,In_679);
and U863 (N_863,In_176,In_625);
nand U864 (N_864,In_57,In_881);
or U865 (N_865,In_301,In_658);
xor U866 (N_866,In_272,In_340);
or U867 (N_867,In_93,In_774);
or U868 (N_868,In_709,In_310);
nand U869 (N_869,In_311,In_580);
nor U870 (N_870,In_595,In_199);
or U871 (N_871,In_205,In_606);
and U872 (N_872,In_85,In_357);
nor U873 (N_873,In_809,In_296);
nor U874 (N_874,In_582,In_685);
nand U875 (N_875,In_267,In_325);
and U876 (N_876,In_334,In_473);
nand U877 (N_877,In_149,In_741);
nand U878 (N_878,In_982,In_494);
and U879 (N_879,In_743,In_461);
nand U880 (N_880,In_475,In_900);
xor U881 (N_881,In_250,In_756);
and U882 (N_882,In_113,In_677);
nand U883 (N_883,In_737,In_194);
nor U884 (N_884,In_955,In_106);
nand U885 (N_885,In_439,In_441);
nor U886 (N_886,In_40,In_37);
nand U887 (N_887,In_810,In_333);
and U888 (N_888,In_343,In_784);
xor U889 (N_889,In_996,In_943);
and U890 (N_890,In_716,In_472);
and U891 (N_891,In_486,In_991);
and U892 (N_892,In_33,In_112);
or U893 (N_893,In_1,In_249);
nand U894 (N_894,In_858,In_372);
nor U895 (N_895,In_527,In_880);
nor U896 (N_896,In_911,In_471);
xnor U897 (N_897,In_848,In_661);
nand U898 (N_898,In_883,In_464);
nor U899 (N_899,In_898,In_821);
xor U900 (N_900,In_274,In_458);
and U901 (N_901,In_702,In_730);
nand U902 (N_902,In_365,In_418);
nand U903 (N_903,In_954,In_263);
or U904 (N_904,In_194,In_434);
xor U905 (N_905,In_543,In_143);
and U906 (N_906,In_827,In_43);
xnor U907 (N_907,In_949,In_611);
nand U908 (N_908,In_96,In_618);
and U909 (N_909,In_135,In_70);
nand U910 (N_910,In_925,In_507);
xor U911 (N_911,In_782,In_355);
or U912 (N_912,In_184,In_575);
nand U913 (N_913,In_519,In_200);
nor U914 (N_914,In_682,In_371);
nor U915 (N_915,In_99,In_480);
and U916 (N_916,In_369,In_945);
and U917 (N_917,In_976,In_264);
or U918 (N_918,In_608,In_223);
xnor U919 (N_919,In_91,In_446);
nand U920 (N_920,In_773,In_251);
nor U921 (N_921,In_128,In_320);
nor U922 (N_922,In_898,In_406);
and U923 (N_923,In_569,In_878);
or U924 (N_924,In_819,In_267);
nand U925 (N_925,In_899,In_444);
nor U926 (N_926,In_139,In_382);
nor U927 (N_927,In_237,In_448);
or U928 (N_928,In_764,In_216);
nand U929 (N_929,In_431,In_809);
and U930 (N_930,In_154,In_704);
nand U931 (N_931,In_192,In_326);
nand U932 (N_932,In_402,In_999);
and U933 (N_933,In_916,In_336);
and U934 (N_934,In_931,In_316);
and U935 (N_935,In_468,In_348);
and U936 (N_936,In_399,In_471);
or U937 (N_937,In_739,In_110);
and U938 (N_938,In_691,In_974);
and U939 (N_939,In_200,In_549);
nand U940 (N_940,In_229,In_598);
nor U941 (N_941,In_737,In_443);
or U942 (N_942,In_714,In_498);
nor U943 (N_943,In_319,In_516);
and U944 (N_944,In_827,In_939);
or U945 (N_945,In_400,In_756);
and U946 (N_946,In_250,In_532);
or U947 (N_947,In_337,In_232);
nand U948 (N_948,In_331,In_741);
and U949 (N_949,In_118,In_938);
and U950 (N_950,In_344,In_709);
and U951 (N_951,In_172,In_313);
and U952 (N_952,In_603,In_369);
or U953 (N_953,In_520,In_372);
nand U954 (N_954,In_877,In_764);
and U955 (N_955,In_608,In_96);
nor U956 (N_956,In_531,In_467);
nor U957 (N_957,In_510,In_242);
nand U958 (N_958,In_480,In_240);
nor U959 (N_959,In_480,In_426);
nand U960 (N_960,In_338,In_123);
nand U961 (N_961,In_426,In_76);
and U962 (N_962,In_237,In_921);
and U963 (N_963,In_436,In_443);
nand U964 (N_964,In_569,In_663);
and U965 (N_965,In_335,In_238);
or U966 (N_966,In_600,In_701);
nand U967 (N_967,In_344,In_796);
nor U968 (N_968,In_770,In_262);
nor U969 (N_969,In_634,In_506);
nor U970 (N_970,In_661,In_950);
or U971 (N_971,In_991,In_137);
and U972 (N_972,In_441,In_340);
and U973 (N_973,In_393,In_89);
nor U974 (N_974,In_858,In_548);
nor U975 (N_975,In_103,In_193);
xnor U976 (N_976,In_926,In_472);
and U977 (N_977,In_666,In_218);
nand U978 (N_978,In_615,In_975);
nand U979 (N_979,In_771,In_858);
nand U980 (N_980,In_664,In_388);
and U981 (N_981,In_943,In_991);
nor U982 (N_982,In_814,In_779);
nand U983 (N_983,In_298,In_602);
xor U984 (N_984,In_867,In_973);
nor U985 (N_985,In_487,In_328);
or U986 (N_986,In_512,In_604);
nor U987 (N_987,In_823,In_477);
or U988 (N_988,In_361,In_621);
or U989 (N_989,In_409,In_466);
and U990 (N_990,In_335,In_572);
and U991 (N_991,In_949,In_908);
and U992 (N_992,In_828,In_143);
nor U993 (N_993,In_57,In_233);
and U994 (N_994,In_408,In_359);
and U995 (N_995,In_172,In_204);
or U996 (N_996,In_66,In_694);
or U997 (N_997,In_894,In_842);
nor U998 (N_998,In_864,In_740);
xnor U999 (N_999,In_672,In_713);
and U1000 (N_1000,In_854,In_111);
nand U1001 (N_1001,In_8,In_579);
nor U1002 (N_1002,In_257,In_457);
nor U1003 (N_1003,In_570,In_434);
and U1004 (N_1004,In_648,In_908);
nand U1005 (N_1005,In_300,In_161);
and U1006 (N_1006,In_569,In_785);
or U1007 (N_1007,In_290,In_716);
nor U1008 (N_1008,In_68,In_565);
and U1009 (N_1009,In_634,In_110);
and U1010 (N_1010,In_935,In_759);
nor U1011 (N_1011,In_716,In_121);
nor U1012 (N_1012,In_587,In_22);
nand U1013 (N_1013,In_163,In_839);
and U1014 (N_1014,In_637,In_207);
nor U1015 (N_1015,In_995,In_419);
xor U1016 (N_1016,In_499,In_95);
and U1017 (N_1017,In_74,In_315);
or U1018 (N_1018,In_107,In_539);
and U1019 (N_1019,In_455,In_712);
nand U1020 (N_1020,In_99,In_487);
nand U1021 (N_1021,In_126,In_862);
nand U1022 (N_1022,In_97,In_702);
xnor U1023 (N_1023,In_157,In_521);
nand U1024 (N_1024,In_765,In_728);
or U1025 (N_1025,In_947,In_111);
nand U1026 (N_1026,In_511,In_347);
nand U1027 (N_1027,In_708,In_680);
nand U1028 (N_1028,In_481,In_686);
nor U1029 (N_1029,In_926,In_758);
or U1030 (N_1030,In_401,In_716);
and U1031 (N_1031,In_717,In_420);
and U1032 (N_1032,In_894,In_404);
nand U1033 (N_1033,In_556,In_489);
and U1034 (N_1034,In_393,In_264);
or U1035 (N_1035,In_268,In_305);
xnor U1036 (N_1036,In_851,In_745);
or U1037 (N_1037,In_682,In_340);
xor U1038 (N_1038,In_477,In_834);
nor U1039 (N_1039,In_573,In_813);
xor U1040 (N_1040,In_783,In_449);
xnor U1041 (N_1041,In_355,In_890);
or U1042 (N_1042,In_266,In_373);
nor U1043 (N_1043,In_254,In_187);
nor U1044 (N_1044,In_920,In_806);
nand U1045 (N_1045,In_441,In_532);
xor U1046 (N_1046,In_445,In_498);
and U1047 (N_1047,In_913,In_866);
xor U1048 (N_1048,In_833,In_836);
and U1049 (N_1049,In_229,In_371);
nand U1050 (N_1050,In_887,In_36);
nand U1051 (N_1051,In_746,In_926);
nor U1052 (N_1052,In_599,In_258);
and U1053 (N_1053,In_143,In_589);
nand U1054 (N_1054,In_918,In_181);
nor U1055 (N_1055,In_948,In_5);
nor U1056 (N_1056,In_103,In_459);
nor U1057 (N_1057,In_177,In_757);
nand U1058 (N_1058,In_927,In_848);
nand U1059 (N_1059,In_394,In_430);
nand U1060 (N_1060,In_37,In_665);
and U1061 (N_1061,In_545,In_177);
xnor U1062 (N_1062,In_60,In_70);
nor U1063 (N_1063,In_818,In_568);
nor U1064 (N_1064,In_641,In_518);
nand U1065 (N_1065,In_96,In_980);
nor U1066 (N_1066,In_169,In_112);
nor U1067 (N_1067,In_242,In_468);
and U1068 (N_1068,In_948,In_567);
or U1069 (N_1069,In_680,In_748);
or U1070 (N_1070,In_498,In_670);
nand U1071 (N_1071,In_150,In_143);
xnor U1072 (N_1072,In_417,In_527);
and U1073 (N_1073,In_801,In_658);
or U1074 (N_1074,In_990,In_312);
nor U1075 (N_1075,In_353,In_309);
or U1076 (N_1076,In_486,In_580);
and U1077 (N_1077,In_496,In_364);
nand U1078 (N_1078,In_293,In_569);
nor U1079 (N_1079,In_689,In_257);
nor U1080 (N_1080,In_874,In_548);
or U1081 (N_1081,In_728,In_380);
xor U1082 (N_1082,In_523,In_657);
nor U1083 (N_1083,In_534,In_327);
nand U1084 (N_1084,In_250,In_606);
or U1085 (N_1085,In_486,In_606);
nand U1086 (N_1086,In_241,In_592);
and U1087 (N_1087,In_594,In_212);
xor U1088 (N_1088,In_306,In_366);
or U1089 (N_1089,In_484,In_552);
and U1090 (N_1090,In_87,In_586);
and U1091 (N_1091,In_920,In_705);
nand U1092 (N_1092,In_831,In_375);
nor U1093 (N_1093,In_872,In_486);
and U1094 (N_1094,In_202,In_661);
xor U1095 (N_1095,In_477,In_276);
and U1096 (N_1096,In_680,In_80);
nand U1097 (N_1097,In_265,In_63);
and U1098 (N_1098,In_981,In_712);
and U1099 (N_1099,In_49,In_778);
nand U1100 (N_1100,In_57,In_330);
nor U1101 (N_1101,In_597,In_364);
and U1102 (N_1102,In_893,In_647);
and U1103 (N_1103,In_938,In_980);
nor U1104 (N_1104,In_123,In_742);
xnor U1105 (N_1105,In_981,In_124);
nor U1106 (N_1106,In_501,In_222);
nand U1107 (N_1107,In_427,In_644);
nor U1108 (N_1108,In_708,In_862);
nand U1109 (N_1109,In_177,In_795);
and U1110 (N_1110,In_19,In_506);
nor U1111 (N_1111,In_893,In_466);
or U1112 (N_1112,In_762,In_637);
nor U1113 (N_1113,In_332,In_967);
and U1114 (N_1114,In_478,In_885);
nor U1115 (N_1115,In_816,In_538);
nand U1116 (N_1116,In_189,In_93);
nor U1117 (N_1117,In_307,In_538);
and U1118 (N_1118,In_459,In_755);
nand U1119 (N_1119,In_850,In_424);
and U1120 (N_1120,In_430,In_781);
xor U1121 (N_1121,In_360,In_546);
nand U1122 (N_1122,In_923,In_824);
nand U1123 (N_1123,In_484,In_317);
and U1124 (N_1124,In_499,In_969);
nand U1125 (N_1125,In_858,In_196);
nand U1126 (N_1126,In_986,In_666);
nand U1127 (N_1127,In_982,In_399);
nand U1128 (N_1128,In_214,In_86);
and U1129 (N_1129,In_595,In_356);
nor U1130 (N_1130,In_579,In_44);
or U1131 (N_1131,In_433,In_311);
nand U1132 (N_1132,In_591,In_782);
xnor U1133 (N_1133,In_528,In_613);
or U1134 (N_1134,In_833,In_710);
nand U1135 (N_1135,In_70,In_827);
nor U1136 (N_1136,In_559,In_915);
and U1137 (N_1137,In_876,In_168);
xnor U1138 (N_1138,In_614,In_869);
or U1139 (N_1139,In_924,In_811);
or U1140 (N_1140,In_276,In_993);
and U1141 (N_1141,In_371,In_412);
nand U1142 (N_1142,In_484,In_407);
nand U1143 (N_1143,In_361,In_200);
or U1144 (N_1144,In_372,In_885);
and U1145 (N_1145,In_734,In_74);
nor U1146 (N_1146,In_101,In_549);
or U1147 (N_1147,In_944,In_10);
or U1148 (N_1148,In_495,In_184);
or U1149 (N_1149,In_660,In_806);
or U1150 (N_1150,In_208,In_894);
or U1151 (N_1151,In_187,In_805);
nand U1152 (N_1152,In_147,In_210);
nand U1153 (N_1153,In_531,In_882);
or U1154 (N_1154,In_265,In_231);
or U1155 (N_1155,In_422,In_711);
xor U1156 (N_1156,In_80,In_773);
nor U1157 (N_1157,In_50,In_861);
nor U1158 (N_1158,In_198,In_93);
and U1159 (N_1159,In_722,In_215);
or U1160 (N_1160,In_973,In_473);
nor U1161 (N_1161,In_486,In_133);
nand U1162 (N_1162,In_239,In_78);
nand U1163 (N_1163,In_602,In_280);
or U1164 (N_1164,In_285,In_565);
xor U1165 (N_1165,In_121,In_743);
and U1166 (N_1166,In_53,In_374);
nor U1167 (N_1167,In_849,In_223);
nor U1168 (N_1168,In_647,In_548);
nor U1169 (N_1169,In_345,In_103);
nor U1170 (N_1170,In_20,In_580);
nor U1171 (N_1171,In_730,In_267);
xor U1172 (N_1172,In_813,In_360);
and U1173 (N_1173,In_395,In_108);
nor U1174 (N_1174,In_708,In_360);
nor U1175 (N_1175,In_876,In_295);
and U1176 (N_1176,In_90,In_617);
or U1177 (N_1177,In_955,In_143);
xnor U1178 (N_1178,In_146,In_956);
and U1179 (N_1179,In_402,In_784);
or U1180 (N_1180,In_557,In_919);
xor U1181 (N_1181,In_832,In_315);
nor U1182 (N_1182,In_69,In_555);
nand U1183 (N_1183,In_674,In_12);
nor U1184 (N_1184,In_116,In_113);
nor U1185 (N_1185,In_685,In_850);
and U1186 (N_1186,In_380,In_348);
and U1187 (N_1187,In_635,In_123);
or U1188 (N_1188,In_904,In_373);
nor U1189 (N_1189,In_864,In_522);
or U1190 (N_1190,In_696,In_991);
xor U1191 (N_1191,In_68,In_84);
or U1192 (N_1192,In_681,In_774);
nand U1193 (N_1193,In_948,In_984);
nand U1194 (N_1194,In_119,In_297);
xnor U1195 (N_1195,In_479,In_385);
nand U1196 (N_1196,In_868,In_951);
or U1197 (N_1197,In_712,In_97);
nand U1198 (N_1198,In_778,In_989);
or U1199 (N_1199,In_52,In_352);
xor U1200 (N_1200,In_626,In_423);
nor U1201 (N_1201,In_616,In_285);
and U1202 (N_1202,In_93,In_825);
nor U1203 (N_1203,In_798,In_456);
xor U1204 (N_1204,In_744,In_591);
nor U1205 (N_1205,In_375,In_586);
nand U1206 (N_1206,In_170,In_191);
and U1207 (N_1207,In_376,In_125);
and U1208 (N_1208,In_597,In_354);
or U1209 (N_1209,In_23,In_765);
nand U1210 (N_1210,In_462,In_397);
nand U1211 (N_1211,In_353,In_487);
nand U1212 (N_1212,In_577,In_233);
or U1213 (N_1213,In_32,In_867);
nand U1214 (N_1214,In_609,In_959);
or U1215 (N_1215,In_802,In_185);
or U1216 (N_1216,In_470,In_745);
nand U1217 (N_1217,In_770,In_853);
xnor U1218 (N_1218,In_803,In_584);
and U1219 (N_1219,In_22,In_585);
xor U1220 (N_1220,In_0,In_979);
nand U1221 (N_1221,In_697,In_47);
nand U1222 (N_1222,In_464,In_763);
and U1223 (N_1223,In_865,In_1);
nand U1224 (N_1224,In_819,In_868);
and U1225 (N_1225,In_830,In_812);
or U1226 (N_1226,In_492,In_539);
nand U1227 (N_1227,In_269,In_323);
and U1228 (N_1228,In_377,In_77);
nor U1229 (N_1229,In_869,In_874);
nor U1230 (N_1230,In_146,In_785);
or U1231 (N_1231,In_197,In_371);
and U1232 (N_1232,In_311,In_84);
nand U1233 (N_1233,In_82,In_299);
nor U1234 (N_1234,In_80,In_322);
and U1235 (N_1235,In_232,In_95);
and U1236 (N_1236,In_56,In_515);
or U1237 (N_1237,In_292,In_640);
xnor U1238 (N_1238,In_808,In_246);
nand U1239 (N_1239,In_277,In_194);
xnor U1240 (N_1240,In_64,In_274);
or U1241 (N_1241,In_766,In_77);
xnor U1242 (N_1242,In_382,In_290);
nor U1243 (N_1243,In_828,In_754);
xnor U1244 (N_1244,In_913,In_357);
nor U1245 (N_1245,In_781,In_872);
and U1246 (N_1246,In_386,In_229);
nand U1247 (N_1247,In_805,In_657);
or U1248 (N_1248,In_217,In_336);
and U1249 (N_1249,In_297,In_734);
and U1250 (N_1250,In_45,In_142);
and U1251 (N_1251,In_925,In_335);
nand U1252 (N_1252,In_830,In_506);
nor U1253 (N_1253,In_861,In_183);
nor U1254 (N_1254,In_726,In_159);
nand U1255 (N_1255,In_81,In_499);
or U1256 (N_1256,In_83,In_693);
and U1257 (N_1257,In_222,In_739);
nor U1258 (N_1258,In_949,In_547);
or U1259 (N_1259,In_141,In_401);
and U1260 (N_1260,In_560,In_684);
nand U1261 (N_1261,In_134,In_364);
and U1262 (N_1262,In_222,In_250);
and U1263 (N_1263,In_428,In_564);
and U1264 (N_1264,In_548,In_667);
xor U1265 (N_1265,In_524,In_772);
and U1266 (N_1266,In_252,In_61);
and U1267 (N_1267,In_628,In_486);
and U1268 (N_1268,In_248,In_260);
nor U1269 (N_1269,In_786,In_445);
and U1270 (N_1270,In_735,In_401);
nor U1271 (N_1271,In_877,In_544);
nand U1272 (N_1272,In_956,In_572);
nor U1273 (N_1273,In_272,In_163);
or U1274 (N_1274,In_465,In_311);
and U1275 (N_1275,In_335,In_981);
nand U1276 (N_1276,In_566,In_534);
nand U1277 (N_1277,In_557,In_135);
nor U1278 (N_1278,In_94,In_519);
and U1279 (N_1279,In_919,In_516);
nor U1280 (N_1280,In_928,In_278);
nand U1281 (N_1281,In_405,In_166);
nand U1282 (N_1282,In_281,In_675);
nor U1283 (N_1283,In_341,In_572);
and U1284 (N_1284,In_944,In_282);
and U1285 (N_1285,In_629,In_591);
nor U1286 (N_1286,In_598,In_536);
and U1287 (N_1287,In_832,In_661);
xor U1288 (N_1288,In_58,In_173);
nor U1289 (N_1289,In_614,In_142);
and U1290 (N_1290,In_187,In_237);
nor U1291 (N_1291,In_387,In_624);
nand U1292 (N_1292,In_814,In_952);
nor U1293 (N_1293,In_376,In_279);
and U1294 (N_1294,In_403,In_813);
and U1295 (N_1295,In_425,In_147);
nand U1296 (N_1296,In_261,In_520);
nor U1297 (N_1297,In_127,In_798);
and U1298 (N_1298,In_540,In_551);
nor U1299 (N_1299,In_836,In_40);
and U1300 (N_1300,In_332,In_445);
nor U1301 (N_1301,In_409,In_407);
xnor U1302 (N_1302,In_277,In_923);
nor U1303 (N_1303,In_59,In_914);
and U1304 (N_1304,In_657,In_186);
or U1305 (N_1305,In_538,In_964);
or U1306 (N_1306,In_690,In_7);
xor U1307 (N_1307,In_329,In_600);
or U1308 (N_1308,In_617,In_750);
xor U1309 (N_1309,In_503,In_441);
and U1310 (N_1310,In_161,In_664);
and U1311 (N_1311,In_398,In_238);
or U1312 (N_1312,In_687,In_5);
nor U1313 (N_1313,In_883,In_589);
nand U1314 (N_1314,In_495,In_115);
xor U1315 (N_1315,In_49,In_600);
and U1316 (N_1316,In_17,In_454);
nor U1317 (N_1317,In_451,In_714);
and U1318 (N_1318,In_35,In_542);
nor U1319 (N_1319,In_945,In_791);
or U1320 (N_1320,In_721,In_466);
nor U1321 (N_1321,In_163,In_138);
or U1322 (N_1322,In_268,In_946);
and U1323 (N_1323,In_603,In_795);
nor U1324 (N_1324,In_954,In_889);
xnor U1325 (N_1325,In_265,In_391);
or U1326 (N_1326,In_451,In_67);
and U1327 (N_1327,In_709,In_64);
nor U1328 (N_1328,In_462,In_31);
nor U1329 (N_1329,In_765,In_819);
or U1330 (N_1330,In_806,In_364);
nor U1331 (N_1331,In_660,In_614);
or U1332 (N_1332,In_336,In_150);
nor U1333 (N_1333,In_948,In_101);
or U1334 (N_1334,In_36,In_550);
and U1335 (N_1335,In_357,In_555);
nand U1336 (N_1336,In_970,In_657);
nor U1337 (N_1337,In_828,In_556);
nand U1338 (N_1338,In_262,In_253);
or U1339 (N_1339,In_404,In_407);
nand U1340 (N_1340,In_408,In_48);
or U1341 (N_1341,In_139,In_997);
nor U1342 (N_1342,In_772,In_316);
or U1343 (N_1343,In_870,In_935);
and U1344 (N_1344,In_584,In_371);
nand U1345 (N_1345,In_280,In_710);
nor U1346 (N_1346,In_799,In_953);
nand U1347 (N_1347,In_968,In_163);
nand U1348 (N_1348,In_254,In_936);
and U1349 (N_1349,In_441,In_708);
xor U1350 (N_1350,In_35,In_444);
nor U1351 (N_1351,In_688,In_631);
and U1352 (N_1352,In_643,In_649);
and U1353 (N_1353,In_549,In_977);
nor U1354 (N_1354,In_140,In_336);
xnor U1355 (N_1355,In_186,In_51);
nand U1356 (N_1356,In_931,In_286);
nor U1357 (N_1357,In_877,In_104);
and U1358 (N_1358,In_29,In_391);
nor U1359 (N_1359,In_175,In_279);
nand U1360 (N_1360,In_992,In_566);
xor U1361 (N_1361,In_728,In_354);
nand U1362 (N_1362,In_680,In_885);
and U1363 (N_1363,In_905,In_51);
nand U1364 (N_1364,In_73,In_835);
nor U1365 (N_1365,In_612,In_844);
xnor U1366 (N_1366,In_577,In_227);
nand U1367 (N_1367,In_3,In_27);
nor U1368 (N_1368,In_398,In_445);
nand U1369 (N_1369,In_568,In_345);
xor U1370 (N_1370,In_810,In_61);
nand U1371 (N_1371,In_51,In_49);
or U1372 (N_1372,In_223,In_635);
and U1373 (N_1373,In_436,In_154);
nand U1374 (N_1374,In_177,In_242);
nand U1375 (N_1375,In_355,In_796);
nand U1376 (N_1376,In_122,In_154);
nor U1377 (N_1377,In_742,In_918);
and U1378 (N_1378,In_136,In_657);
and U1379 (N_1379,In_118,In_286);
nand U1380 (N_1380,In_21,In_662);
or U1381 (N_1381,In_77,In_700);
xnor U1382 (N_1382,In_532,In_325);
xor U1383 (N_1383,In_675,In_148);
nand U1384 (N_1384,In_489,In_469);
nor U1385 (N_1385,In_951,In_726);
xnor U1386 (N_1386,In_516,In_310);
xor U1387 (N_1387,In_795,In_906);
and U1388 (N_1388,In_159,In_519);
and U1389 (N_1389,In_112,In_608);
nor U1390 (N_1390,In_137,In_602);
or U1391 (N_1391,In_22,In_576);
and U1392 (N_1392,In_49,In_78);
and U1393 (N_1393,In_272,In_758);
or U1394 (N_1394,In_555,In_963);
and U1395 (N_1395,In_868,In_900);
nand U1396 (N_1396,In_229,In_31);
nor U1397 (N_1397,In_574,In_283);
and U1398 (N_1398,In_275,In_148);
nand U1399 (N_1399,In_347,In_351);
xnor U1400 (N_1400,In_548,In_352);
or U1401 (N_1401,In_926,In_660);
nand U1402 (N_1402,In_12,In_51);
nor U1403 (N_1403,In_354,In_568);
or U1404 (N_1404,In_231,In_697);
nand U1405 (N_1405,In_716,In_933);
and U1406 (N_1406,In_313,In_407);
nor U1407 (N_1407,In_27,In_386);
nand U1408 (N_1408,In_395,In_583);
and U1409 (N_1409,In_959,In_288);
xnor U1410 (N_1410,In_379,In_274);
nand U1411 (N_1411,In_916,In_567);
nand U1412 (N_1412,In_247,In_667);
nor U1413 (N_1413,In_672,In_377);
or U1414 (N_1414,In_582,In_90);
nor U1415 (N_1415,In_611,In_871);
or U1416 (N_1416,In_827,In_328);
nand U1417 (N_1417,In_249,In_530);
or U1418 (N_1418,In_232,In_244);
or U1419 (N_1419,In_638,In_794);
or U1420 (N_1420,In_720,In_56);
nand U1421 (N_1421,In_653,In_926);
or U1422 (N_1422,In_387,In_381);
and U1423 (N_1423,In_319,In_204);
or U1424 (N_1424,In_37,In_531);
and U1425 (N_1425,In_193,In_674);
and U1426 (N_1426,In_103,In_89);
or U1427 (N_1427,In_520,In_733);
nor U1428 (N_1428,In_466,In_389);
nand U1429 (N_1429,In_716,In_915);
xnor U1430 (N_1430,In_18,In_987);
or U1431 (N_1431,In_248,In_506);
nand U1432 (N_1432,In_61,In_721);
nor U1433 (N_1433,In_296,In_929);
nor U1434 (N_1434,In_339,In_137);
nand U1435 (N_1435,In_897,In_686);
or U1436 (N_1436,In_779,In_351);
nand U1437 (N_1437,In_278,In_808);
and U1438 (N_1438,In_792,In_330);
and U1439 (N_1439,In_551,In_397);
xnor U1440 (N_1440,In_240,In_83);
and U1441 (N_1441,In_80,In_952);
xnor U1442 (N_1442,In_345,In_150);
nand U1443 (N_1443,In_733,In_130);
nor U1444 (N_1444,In_599,In_769);
xor U1445 (N_1445,In_961,In_396);
nand U1446 (N_1446,In_991,In_154);
nor U1447 (N_1447,In_707,In_972);
nand U1448 (N_1448,In_708,In_784);
xnor U1449 (N_1449,In_580,In_56);
or U1450 (N_1450,In_14,In_679);
nand U1451 (N_1451,In_298,In_983);
nand U1452 (N_1452,In_477,In_712);
and U1453 (N_1453,In_673,In_572);
and U1454 (N_1454,In_855,In_946);
and U1455 (N_1455,In_792,In_359);
nand U1456 (N_1456,In_739,In_675);
nand U1457 (N_1457,In_700,In_235);
or U1458 (N_1458,In_857,In_674);
nor U1459 (N_1459,In_860,In_195);
or U1460 (N_1460,In_636,In_934);
nand U1461 (N_1461,In_70,In_507);
and U1462 (N_1462,In_234,In_109);
and U1463 (N_1463,In_874,In_41);
and U1464 (N_1464,In_688,In_236);
and U1465 (N_1465,In_513,In_156);
nor U1466 (N_1466,In_570,In_508);
nor U1467 (N_1467,In_422,In_449);
nor U1468 (N_1468,In_533,In_210);
xnor U1469 (N_1469,In_15,In_518);
xor U1470 (N_1470,In_788,In_29);
nor U1471 (N_1471,In_573,In_286);
and U1472 (N_1472,In_588,In_529);
nand U1473 (N_1473,In_224,In_953);
xnor U1474 (N_1474,In_420,In_737);
or U1475 (N_1475,In_391,In_801);
nand U1476 (N_1476,In_219,In_591);
or U1477 (N_1477,In_106,In_193);
nand U1478 (N_1478,In_895,In_958);
nor U1479 (N_1479,In_47,In_801);
and U1480 (N_1480,In_348,In_673);
nand U1481 (N_1481,In_410,In_783);
and U1482 (N_1482,In_361,In_738);
or U1483 (N_1483,In_734,In_437);
nand U1484 (N_1484,In_259,In_875);
or U1485 (N_1485,In_629,In_645);
and U1486 (N_1486,In_949,In_223);
nand U1487 (N_1487,In_37,In_967);
nor U1488 (N_1488,In_229,In_925);
nand U1489 (N_1489,In_314,In_641);
nor U1490 (N_1490,In_810,In_654);
or U1491 (N_1491,In_518,In_422);
nor U1492 (N_1492,In_622,In_204);
nand U1493 (N_1493,In_715,In_881);
xor U1494 (N_1494,In_851,In_923);
nor U1495 (N_1495,In_258,In_590);
nor U1496 (N_1496,In_715,In_446);
nor U1497 (N_1497,In_925,In_904);
nor U1498 (N_1498,In_476,In_149);
nand U1499 (N_1499,In_575,In_642);
or U1500 (N_1500,In_178,In_309);
nand U1501 (N_1501,In_460,In_407);
nand U1502 (N_1502,In_922,In_666);
and U1503 (N_1503,In_586,In_756);
nand U1504 (N_1504,In_423,In_951);
nand U1505 (N_1505,In_415,In_632);
nor U1506 (N_1506,In_17,In_552);
or U1507 (N_1507,In_793,In_797);
nor U1508 (N_1508,In_777,In_923);
or U1509 (N_1509,In_881,In_484);
and U1510 (N_1510,In_109,In_571);
or U1511 (N_1511,In_403,In_871);
xor U1512 (N_1512,In_186,In_844);
and U1513 (N_1513,In_673,In_894);
or U1514 (N_1514,In_301,In_133);
nand U1515 (N_1515,In_773,In_795);
nor U1516 (N_1516,In_197,In_589);
and U1517 (N_1517,In_384,In_886);
nor U1518 (N_1518,In_952,In_965);
nand U1519 (N_1519,In_600,In_254);
and U1520 (N_1520,In_622,In_810);
and U1521 (N_1521,In_666,In_967);
and U1522 (N_1522,In_909,In_217);
xor U1523 (N_1523,In_275,In_580);
or U1524 (N_1524,In_835,In_273);
nand U1525 (N_1525,In_583,In_324);
xnor U1526 (N_1526,In_626,In_821);
nor U1527 (N_1527,In_421,In_386);
and U1528 (N_1528,In_938,In_641);
nor U1529 (N_1529,In_531,In_54);
nor U1530 (N_1530,In_217,In_77);
and U1531 (N_1531,In_919,In_893);
nor U1532 (N_1532,In_894,In_255);
nand U1533 (N_1533,In_59,In_58);
nor U1534 (N_1534,In_618,In_223);
and U1535 (N_1535,In_906,In_792);
and U1536 (N_1536,In_118,In_616);
or U1537 (N_1537,In_431,In_873);
nor U1538 (N_1538,In_420,In_744);
nor U1539 (N_1539,In_797,In_606);
and U1540 (N_1540,In_905,In_260);
nor U1541 (N_1541,In_403,In_734);
or U1542 (N_1542,In_327,In_955);
or U1543 (N_1543,In_18,In_9);
or U1544 (N_1544,In_350,In_955);
nor U1545 (N_1545,In_399,In_356);
and U1546 (N_1546,In_481,In_860);
nand U1547 (N_1547,In_611,In_840);
and U1548 (N_1548,In_221,In_950);
and U1549 (N_1549,In_682,In_956);
and U1550 (N_1550,In_662,In_389);
nand U1551 (N_1551,In_595,In_559);
or U1552 (N_1552,In_843,In_634);
and U1553 (N_1553,In_572,In_7);
nand U1554 (N_1554,In_308,In_776);
and U1555 (N_1555,In_62,In_516);
and U1556 (N_1556,In_931,In_853);
and U1557 (N_1557,In_527,In_197);
nand U1558 (N_1558,In_760,In_403);
nand U1559 (N_1559,In_816,In_856);
nand U1560 (N_1560,In_712,In_399);
and U1561 (N_1561,In_34,In_920);
nor U1562 (N_1562,In_611,In_10);
nor U1563 (N_1563,In_399,In_140);
or U1564 (N_1564,In_788,In_654);
or U1565 (N_1565,In_308,In_890);
nand U1566 (N_1566,In_522,In_721);
and U1567 (N_1567,In_702,In_744);
and U1568 (N_1568,In_463,In_762);
nand U1569 (N_1569,In_619,In_673);
xor U1570 (N_1570,In_209,In_530);
xnor U1571 (N_1571,In_158,In_680);
nand U1572 (N_1572,In_761,In_540);
and U1573 (N_1573,In_614,In_253);
nand U1574 (N_1574,In_703,In_631);
xor U1575 (N_1575,In_645,In_54);
and U1576 (N_1576,In_722,In_224);
nor U1577 (N_1577,In_120,In_102);
and U1578 (N_1578,In_144,In_52);
or U1579 (N_1579,In_272,In_219);
nor U1580 (N_1580,In_447,In_723);
and U1581 (N_1581,In_783,In_557);
or U1582 (N_1582,In_811,In_192);
nor U1583 (N_1583,In_524,In_347);
nor U1584 (N_1584,In_36,In_653);
xnor U1585 (N_1585,In_626,In_215);
and U1586 (N_1586,In_810,In_242);
and U1587 (N_1587,In_322,In_670);
and U1588 (N_1588,In_90,In_571);
nor U1589 (N_1589,In_183,In_145);
or U1590 (N_1590,In_712,In_769);
nand U1591 (N_1591,In_518,In_313);
xor U1592 (N_1592,In_897,In_243);
nor U1593 (N_1593,In_374,In_22);
or U1594 (N_1594,In_809,In_840);
and U1595 (N_1595,In_596,In_107);
nor U1596 (N_1596,In_518,In_397);
and U1597 (N_1597,In_353,In_742);
nor U1598 (N_1598,In_900,In_244);
nand U1599 (N_1599,In_669,In_982);
nand U1600 (N_1600,In_360,In_574);
xor U1601 (N_1601,In_461,In_28);
xor U1602 (N_1602,In_176,In_938);
nand U1603 (N_1603,In_650,In_954);
nand U1604 (N_1604,In_888,In_78);
and U1605 (N_1605,In_356,In_183);
nand U1606 (N_1606,In_459,In_426);
nor U1607 (N_1607,In_806,In_211);
and U1608 (N_1608,In_604,In_705);
nor U1609 (N_1609,In_820,In_960);
or U1610 (N_1610,In_499,In_523);
and U1611 (N_1611,In_760,In_2);
nand U1612 (N_1612,In_118,In_110);
and U1613 (N_1613,In_961,In_809);
nor U1614 (N_1614,In_773,In_667);
and U1615 (N_1615,In_494,In_450);
nand U1616 (N_1616,In_204,In_547);
or U1617 (N_1617,In_237,In_670);
and U1618 (N_1618,In_10,In_694);
or U1619 (N_1619,In_993,In_411);
nor U1620 (N_1620,In_975,In_814);
nor U1621 (N_1621,In_962,In_992);
nand U1622 (N_1622,In_838,In_321);
or U1623 (N_1623,In_789,In_526);
nand U1624 (N_1624,In_404,In_653);
nand U1625 (N_1625,In_534,In_876);
nor U1626 (N_1626,In_847,In_537);
xnor U1627 (N_1627,In_109,In_783);
and U1628 (N_1628,In_865,In_558);
xnor U1629 (N_1629,In_352,In_246);
nor U1630 (N_1630,In_903,In_65);
or U1631 (N_1631,In_796,In_13);
and U1632 (N_1632,In_370,In_25);
nor U1633 (N_1633,In_915,In_969);
xor U1634 (N_1634,In_285,In_446);
nand U1635 (N_1635,In_896,In_362);
nor U1636 (N_1636,In_708,In_127);
nand U1637 (N_1637,In_872,In_422);
nand U1638 (N_1638,In_742,In_443);
and U1639 (N_1639,In_19,In_654);
nor U1640 (N_1640,In_667,In_623);
or U1641 (N_1641,In_881,In_551);
or U1642 (N_1642,In_659,In_900);
and U1643 (N_1643,In_164,In_815);
or U1644 (N_1644,In_33,In_197);
or U1645 (N_1645,In_46,In_898);
nand U1646 (N_1646,In_218,In_601);
and U1647 (N_1647,In_662,In_656);
xor U1648 (N_1648,In_970,In_188);
nand U1649 (N_1649,In_387,In_706);
nor U1650 (N_1650,In_189,In_416);
or U1651 (N_1651,In_230,In_766);
nor U1652 (N_1652,In_450,In_882);
or U1653 (N_1653,In_529,In_206);
nand U1654 (N_1654,In_505,In_292);
nand U1655 (N_1655,In_255,In_253);
nand U1656 (N_1656,In_609,In_313);
nand U1657 (N_1657,In_512,In_148);
or U1658 (N_1658,In_316,In_610);
nand U1659 (N_1659,In_837,In_116);
nor U1660 (N_1660,In_745,In_106);
xor U1661 (N_1661,In_605,In_132);
nor U1662 (N_1662,In_721,In_988);
xor U1663 (N_1663,In_36,In_916);
nand U1664 (N_1664,In_421,In_425);
xnor U1665 (N_1665,In_674,In_277);
nand U1666 (N_1666,In_828,In_39);
or U1667 (N_1667,In_25,In_101);
nand U1668 (N_1668,In_237,In_189);
nor U1669 (N_1669,In_449,In_241);
nand U1670 (N_1670,In_924,In_304);
nand U1671 (N_1671,In_774,In_968);
nand U1672 (N_1672,In_437,In_818);
nand U1673 (N_1673,In_387,In_337);
nor U1674 (N_1674,In_435,In_103);
nor U1675 (N_1675,In_208,In_603);
nand U1676 (N_1676,In_909,In_830);
nand U1677 (N_1677,In_29,In_49);
nor U1678 (N_1678,In_800,In_994);
nand U1679 (N_1679,In_380,In_325);
nor U1680 (N_1680,In_462,In_333);
nand U1681 (N_1681,In_452,In_518);
and U1682 (N_1682,In_16,In_581);
and U1683 (N_1683,In_287,In_664);
xor U1684 (N_1684,In_103,In_344);
nor U1685 (N_1685,In_27,In_94);
or U1686 (N_1686,In_893,In_836);
and U1687 (N_1687,In_519,In_972);
and U1688 (N_1688,In_311,In_838);
and U1689 (N_1689,In_526,In_191);
nor U1690 (N_1690,In_863,In_754);
nand U1691 (N_1691,In_812,In_775);
or U1692 (N_1692,In_248,In_735);
nand U1693 (N_1693,In_49,In_368);
nor U1694 (N_1694,In_163,In_809);
nand U1695 (N_1695,In_625,In_76);
nand U1696 (N_1696,In_363,In_184);
nor U1697 (N_1697,In_693,In_402);
xor U1698 (N_1698,In_497,In_879);
and U1699 (N_1699,In_308,In_681);
nand U1700 (N_1700,In_105,In_368);
and U1701 (N_1701,In_937,In_955);
or U1702 (N_1702,In_28,In_975);
nor U1703 (N_1703,In_913,In_413);
nor U1704 (N_1704,In_13,In_217);
and U1705 (N_1705,In_138,In_686);
and U1706 (N_1706,In_658,In_113);
and U1707 (N_1707,In_387,In_378);
nand U1708 (N_1708,In_183,In_731);
nor U1709 (N_1709,In_435,In_247);
and U1710 (N_1710,In_195,In_11);
and U1711 (N_1711,In_321,In_933);
and U1712 (N_1712,In_933,In_802);
or U1713 (N_1713,In_123,In_501);
nand U1714 (N_1714,In_842,In_337);
nand U1715 (N_1715,In_396,In_569);
nor U1716 (N_1716,In_67,In_574);
nand U1717 (N_1717,In_488,In_714);
nand U1718 (N_1718,In_61,In_366);
nand U1719 (N_1719,In_315,In_432);
nor U1720 (N_1720,In_549,In_89);
or U1721 (N_1721,In_980,In_856);
nand U1722 (N_1722,In_668,In_227);
and U1723 (N_1723,In_394,In_925);
nand U1724 (N_1724,In_778,In_967);
nor U1725 (N_1725,In_181,In_561);
and U1726 (N_1726,In_245,In_685);
nor U1727 (N_1727,In_460,In_279);
nand U1728 (N_1728,In_698,In_582);
nor U1729 (N_1729,In_662,In_960);
or U1730 (N_1730,In_280,In_980);
and U1731 (N_1731,In_192,In_786);
and U1732 (N_1732,In_702,In_708);
xor U1733 (N_1733,In_500,In_292);
and U1734 (N_1734,In_462,In_804);
nand U1735 (N_1735,In_554,In_241);
or U1736 (N_1736,In_599,In_31);
nor U1737 (N_1737,In_180,In_688);
xnor U1738 (N_1738,In_376,In_850);
or U1739 (N_1739,In_570,In_930);
and U1740 (N_1740,In_793,In_203);
nand U1741 (N_1741,In_287,In_478);
or U1742 (N_1742,In_985,In_569);
nand U1743 (N_1743,In_286,In_48);
nor U1744 (N_1744,In_610,In_725);
nand U1745 (N_1745,In_506,In_987);
and U1746 (N_1746,In_243,In_294);
nand U1747 (N_1747,In_760,In_595);
or U1748 (N_1748,In_451,In_748);
and U1749 (N_1749,In_619,In_14);
and U1750 (N_1750,In_390,In_201);
nor U1751 (N_1751,In_719,In_246);
nand U1752 (N_1752,In_831,In_326);
and U1753 (N_1753,In_554,In_595);
nor U1754 (N_1754,In_42,In_36);
nand U1755 (N_1755,In_973,In_113);
and U1756 (N_1756,In_152,In_516);
xor U1757 (N_1757,In_837,In_925);
nand U1758 (N_1758,In_324,In_669);
and U1759 (N_1759,In_388,In_8);
nor U1760 (N_1760,In_756,In_696);
and U1761 (N_1761,In_550,In_93);
nor U1762 (N_1762,In_777,In_188);
nor U1763 (N_1763,In_286,In_417);
nor U1764 (N_1764,In_330,In_147);
nor U1765 (N_1765,In_932,In_977);
and U1766 (N_1766,In_436,In_265);
nand U1767 (N_1767,In_592,In_200);
or U1768 (N_1768,In_55,In_747);
nor U1769 (N_1769,In_740,In_616);
or U1770 (N_1770,In_866,In_989);
nor U1771 (N_1771,In_708,In_331);
nor U1772 (N_1772,In_791,In_619);
nor U1773 (N_1773,In_534,In_159);
or U1774 (N_1774,In_703,In_633);
nand U1775 (N_1775,In_71,In_597);
nor U1776 (N_1776,In_978,In_765);
or U1777 (N_1777,In_455,In_531);
nand U1778 (N_1778,In_436,In_784);
or U1779 (N_1779,In_714,In_534);
nand U1780 (N_1780,In_392,In_832);
nor U1781 (N_1781,In_917,In_849);
and U1782 (N_1782,In_930,In_684);
nor U1783 (N_1783,In_413,In_830);
and U1784 (N_1784,In_800,In_511);
nor U1785 (N_1785,In_337,In_362);
nand U1786 (N_1786,In_107,In_154);
nand U1787 (N_1787,In_747,In_199);
nand U1788 (N_1788,In_968,In_157);
nand U1789 (N_1789,In_225,In_665);
or U1790 (N_1790,In_912,In_697);
and U1791 (N_1791,In_462,In_861);
or U1792 (N_1792,In_634,In_836);
or U1793 (N_1793,In_661,In_382);
nand U1794 (N_1794,In_95,In_118);
xor U1795 (N_1795,In_307,In_610);
nor U1796 (N_1796,In_169,In_223);
xor U1797 (N_1797,In_149,In_436);
nor U1798 (N_1798,In_714,In_937);
and U1799 (N_1799,In_181,In_321);
xor U1800 (N_1800,In_757,In_491);
or U1801 (N_1801,In_0,In_804);
nor U1802 (N_1802,In_171,In_240);
or U1803 (N_1803,In_664,In_574);
or U1804 (N_1804,In_39,In_232);
and U1805 (N_1805,In_514,In_441);
and U1806 (N_1806,In_193,In_414);
nor U1807 (N_1807,In_769,In_283);
or U1808 (N_1808,In_56,In_709);
nor U1809 (N_1809,In_872,In_676);
or U1810 (N_1810,In_542,In_97);
and U1811 (N_1811,In_242,In_996);
or U1812 (N_1812,In_556,In_45);
nand U1813 (N_1813,In_46,In_774);
nor U1814 (N_1814,In_369,In_918);
nor U1815 (N_1815,In_576,In_709);
or U1816 (N_1816,In_528,In_986);
nand U1817 (N_1817,In_275,In_409);
xor U1818 (N_1818,In_679,In_463);
nand U1819 (N_1819,In_793,In_195);
or U1820 (N_1820,In_678,In_971);
nand U1821 (N_1821,In_477,In_47);
nand U1822 (N_1822,In_445,In_142);
or U1823 (N_1823,In_884,In_760);
nor U1824 (N_1824,In_817,In_979);
nand U1825 (N_1825,In_913,In_265);
nor U1826 (N_1826,In_380,In_942);
and U1827 (N_1827,In_398,In_744);
xnor U1828 (N_1828,In_353,In_400);
and U1829 (N_1829,In_87,In_457);
nor U1830 (N_1830,In_330,In_913);
or U1831 (N_1831,In_656,In_263);
xor U1832 (N_1832,In_386,In_637);
or U1833 (N_1833,In_47,In_107);
and U1834 (N_1834,In_775,In_782);
and U1835 (N_1835,In_71,In_398);
nor U1836 (N_1836,In_530,In_276);
and U1837 (N_1837,In_681,In_463);
and U1838 (N_1838,In_294,In_780);
and U1839 (N_1839,In_649,In_526);
and U1840 (N_1840,In_650,In_173);
or U1841 (N_1841,In_420,In_891);
or U1842 (N_1842,In_550,In_774);
nor U1843 (N_1843,In_131,In_508);
nor U1844 (N_1844,In_94,In_372);
or U1845 (N_1845,In_471,In_891);
xor U1846 (N_1846,In_853,In_53);
nand U1847 (N_1847,In_753,In_398);
nor U1848 (N_1848,In_339,In_190);
nor U1849 (N_1849,In_14,In_329);
nand U1850 (N_1850,In_593,In_61);
nor U1851 (N_1851,In_175,In_152);
nor U1852 (N_1852,In_69,In_392);
or U1853 (N_1853,In_240,In_711);
or U1854 (N_1854,In_88,In_962);
nand U1855 (N_1855,In_864,In_233);
and U1856 (N_1856,In_684,In_854);
nand U1857 (N_1857,In_473,In_424);
nand U1858 (N_1858,In_875,In_26);
xnor U1859 (N_1859,In_157,In_321);
xnor U1860 (N_1860,In_742,In_585);
nand U1861 (N_1861,In_916,In_181);
nor U1862 (N_1862,In_642,In_670);
or U1863 (N_1863,In_892,In_180);
or U1864 (N_1864,In_414,In_897);
nand U1865 (N_1865,In_186,In_184);
nand U1866 (N_1866,In_365,In_842);
xnor U1867 (N_1867,In_467,In_396);
nand U1868 (N_1868,In_912,In_48);
nor U1869 (N_1869,In_207,In_312);
or U1870 (N_1870,In_734,In_314);
or U1871 (N_1871,In_121,In_672);
nand U1872 (N_1872,In_933,In_659);
nor U1873 (N_1873,In_131,In_481);
nand U1874 (N_1874,In_716,In_238);
nand U1875 (N_1875,In_531,In_317);
nand U1876 (N_1876,In_153,In_351);
and U1877 (N_1877,In_105,In_68);
nand U1878 (N_1878,In_143,In_757);
xor U1879 (N_1879,In_858,In_409);
or U1880 (N_1880,In_948,In_557);
xnor U1881 (N_1881,In_671,In_437);
nor U1882 (N_1882,In_353,In_839);
and U1883 (N_1883,In_593,In_142);
nor U1884 (N_1884,In_819,In_407);
nor U1885 (N_1885,In_781,In_864);
nor U1886 (N_1886,In_255,In_879);
nor U1887 (N_1887,In_374,In_227);
or U1888 (N_1888,In_724,In_330);
nor U1889 (N_1889,In_205,In_318);
nor U1890 (N_1890,In_108,In_470);
or U1891 (N_1891,In_769,In_64);
and U1892 (N_1892,In_844,In_230);
and U1893 (N_1893,In_780,In_746);
nor U1894 (N_1894,In_702,In_306);
xnor U1895 (N_1895,In_207,In_213);
nand U1896 (N_1896,In_617,In_192);
nor U1897 (N_1897,In_952,In_261);
or U1898 (N_1898,In_466,In_582);
nor U1899 (N_1899,In_472,In_170);
nor U1900 (N_1900,In_516,In_6);
and U1901 (N_1901,In_352,In_277);
nor U1902 (N_1902,In_687,In_664);
nor U1903 (N_1903,In_293,In_583);
or U1904 (N_1904,In_614,In_473);
or U1905 (N_1905,In_202,In_337);
nand U1906 (N_1906,In_645,In_5);
nor U1907 (N_1907,In_846,In_314);
nor U1908 (N_1908,In_937,In_283);
or U1909 (N_1909,In_133,In_462);
xor U1910 (N_1910,In_57,In_294);
xnor U1911 (N_1911,In_557,In_982);
nand U1912 (N_1912,In_665,In_193);
or U1913 (N_1913,In_509,In_262);
nand U1914 (N_1914,In_645,In_788);
nor U1915 (N_1915,In_920,In_470);
nor U1916 (N_1916,In_434,In_860);
or U1917 (N_1917,In_354,In_780);
or U1918 (N_1918,In_810,In_220);
or U1919 (N_1919,In_41,In_510);
and U1920 (N_1920,In_830,In_733);
xor U1921 (N_1921,In_328,In_245);
and U1922 (N_1922,In_247,In_113);
nand U1923 (N_1923,In_695,In_372);
and U1924 (N_1924,In_732,In_42);
or U1925 (N_1925,In_654,In_422);
or U1926 (N_1926,In_256,In_385);
nand U1927 (N_1927,In_678,In_366);
or U1928 (N_1928,In_553,In_754);
or U1929 (N_1929,In_507,In_16);
nand U1930 (N_1930,In_343,In_848);
or U1931 (N_1931,In_669,In_818);
or U1932 (N_1932,In_732,In_676);
nand U1933 (N_1933,In_728,In_147);
nand U1934 (N_1934,In_554,In_913);
nor U1935 (N_1935,In_520,In_968);
nand U1936 (N_1936,In_804,In_519);
xnor U1937 (N_1937,In_543,In_10);
nor U1938 (N_1938,In_178,In_819);
nor U1939 (N_1939,In_445,In_970);
nor U1940 (N_1940,In_713,In_761);
and U1941 (N_1941,In_678,In_170);
and U1942 (N_1942,In_810,In_25);
and U1943 (N_1943,In_655,In_377);
and U1944 (N_1944,In_406,In_824);
and U1945 (N_1945,In_596,In_403);
nand U1946 (N_1946,In_829,In_417);
and U1947 (N_1947,In_200,In_331);
nand U1948 (N_1948,In_632,In_490);
or U1949 (N_1949,In_727,In_261);
nor U1950 (N_1950,In_27,In_480);
xnor U1951 (N_1951,In_552,In_338);
and U1952 (N_1952,In_936,In_487);
nand U1953 (N_1953,In_794,In_217);
xnor U1954 (N_1954,In_267,In_75);
nand U1955 (N_1955,In_390,In_593);
nand U1956 (N_1956,In_307,In_18);
nor U1957 (N_1957,In_797,In_525);
nand U1958 (N_1958,In_758,In_632);
or U1959 (N_1959,In_159,In_846);
nand U1960 (N_1960,In_52,In_911);
nand U1961 (N_1961,In_387,In_32);
nand U1962 (N_1962,In_978,In_499);
xor U1963 (N_1963,In_676,In_160);
or U1964 (N_1964,In_664,In_651);
nor U1965 (N_1965,In_11,In_246);
or U1966 (N_1966,In_392,In_229);
and U1967 (N_1967,In_12,In_169);
nor U1968 (N_1968,In_44,In_657);
and U1969 (N_1969,In_173,In_882);
nand U1970 (N_1970,In_56,In_668);
and U1971 (N_1971,In_522,In_638);
nand U1972 (N_1972,In_834,In_799);
or U1973 (N_1973,In_227,In_718);
or U1974 (N_1974,In_39,In_13);
xnor U1975 (N_1975,In_167,In_921);
xnor U1976 (N_1976,In_525,In_485);
or U1977 (N_1977,In_172,In_457);
nor U1978 (N_1978,In_867,In_898);
nand U1979 (N_1979,In_352,In_468);
xnor U1980 (N_1980,In_17,In_78);
xor U1981 (N_1981,In_214,In_308);
nor U1982 (N_1982,In_224,In_592);
nor U1983 (N_1983,In_211,In_492);
nor U1984 (N_1984,In_219,In_67);
nor U1985 (N_1985,In_943,In_533);
and U1986 (N_1986,In_675,In_450);
nand U1987 (N_1987,In_582,In_502);
or U1988 (N_1988,In_247,In_446);
or U1989 (N_1989,In_775,In_588);
and U1990 (N_1990,In_406,In_253);
nor U1991 (N_1991,In_9,In_620);
and U1992 (N_1992,In_666,In_810);
and U1993 (N_1993,In_745,In_635);
nor U1994 (N_1994,In_117,In_153);
xor U1995 (N_1995,In_282,In_268);
or U1996 (N_1996,In_227,In_683);
nand U1997 (N_1997,In_120,In_88);
nand U1998 (N_1998,In_25,In_161);
and U1999 (N_1999,In_322,In_754);
or U2000 (N_2000,In_732,In_753);
and U2001 (N_2001,In_878,In_456);
xor U2002 (N_2002,In_167,In_68);
nand U2003 (N_2003,In_797,In_12);
xor U2004 (N_2004,In_199,In_665);
or U2005 (N_2005,In_807,In_60);
xnor U2006 (N_2006,In_260,In_650);
xor U2007 (N_2007,In_248,In_166);
and U2008 (N_2008,In_210,In_743);
or U2009 (N_2009,In_543,In_913);
nor U2010 (N_2010,In_600,In_639);
or U2011 (N_2011,In_287,In_687);
nand U2012 (N_2012,In_907,In_538);
and U2013 (N_2013,In_36,In_315);
or U2014 (N_2014,In_87,In_247);
nor U2015 (N_2015,In_995,In_849);
or U2016 (N_2016,In_437,In_793);
nor U2017 (N_2017,In_660,In_56);
xor U2018 (N_2018,In_389,In_922);
nand U2019 (N_2019,In_602,In_328);
and U2020 (N_2020,In_267,In_958);
and U2021 (N_2021,In_861,In_141);
xor U2022 (N_2022,In_665,In_704);
or U2023 (N_2023,In_133,In_17);
nor U2024 (N_2024,In_836,In_838);
xnor U2025 (N_2025,In_854,In_977);
or U2026 (N_2026,In_78,In_930);
and U2027 (N_2027,In_15,In_40);
xor U2028 (N_2028,In_644,In_935);
nand U2029 (N_2029,In_481,In_533);
nand U2030 (N_2030,In_867,In_908);
or U2031 (N_2031,In_649,In_21);
xor U2032 (N_2032,In_921,In_754);
and U2033 (N_2033,In_637,In_190);
or U2034 (N_2034,In_26,In_531);
or U2035 (N_2035,In_968,In_368);
nor U2036 (N_2036,In_795,In_464);
and U2037 (N_2037,In_889,In_579);
or U2038 (N_2038,In_973,In_764);
nand U2039 (N_2039,In_9,In_374);
nand U2040 (N_2040,In_512,In_311);
or U2041 (N_2041,In_742,In_48);
nand U2042 (N_2042,In_659,In_343);
nor U2043 (N_2043,In_179,In_354);
nand U2044 (N_2044,In_869,In_574);
and U2045 (N_2045,In_234,In_682);
nand U2046 (N_2046,In_806,In_726);
or U2047 (N_2047,In_850,In_769);
and U2048 (N_2048,In_757,In_47);
and U2049 (N_2049,In_35,In_130);
and U2050 (N_2050,In_892,In_903);
and U2051 (N_2051,In_470,In_899);
xor U2052 (N_2052,In_225,In_902);
nand U2053 (N_2053,In_433,In_380);
and U2054 (N_2054,In_311,In_989);
xnor U2055 (N_2055,In_264,In_16);
xnor U2056 (N_2056,In_725,In_640);
and U2057 (N_2057,In_896,In_113);
nor U2058 (N_2058,In_259,In_873);
nand U2059 (N_2059,In_66,In_569);
nand U2060 (N_2060,In_849,In_985);
xor U2061 (N_2061,In_542,In_146);
or U2062 (N_2062,In_48,In_164);
or U2063 (N_2063,In_828,In_435);
nand U2064 (N_2064,In_206,In_697);
or U2065 (N_2065,In_894,In_693);
and U2066 (N_2066,In_589,In_629);
xnor U2067 (N_2067,In_309,In_798);
or U2068 (N_2068,In_338,In_473);
xnor U2069 (N_2069,In_881,In_975);
nand U2070 (N_2070,In_664,In_63);
and U2071 (N_2071,In_112,In_347);
or U2072 (N_2072,In_721,In_574);
nand U2073 (N_2073,In_726,In_774);
and U2074 (N_2074,In_80,In_300);
nand U2075 (N_2075,In_988,In_390);
nand U2076 (N_2076,In_766,In_368);
and U2077 (N_2077,In_343,In_878);
nor U2078 (N_2078,In_284,In_751);
xnor U2079 (N_2079,In_535,In_913);
nor U2080 (N_2080,In_280,In_942);
xor U2081 (N_2081,In_282,In_565);
nand U2082 (N_2082,In_891,In_352);
and U2083 (N_2083,In_327,In_698);
and U2084 (N_2084,In_131,In_253);
and U2085 (N_2085,In_130,In_563);
or U2086 (N_2086,In_805,In_31);
nand U2087 (N_2087,In_401,In_74);
nand U2088 (N_2088,In_847,In_310);
and U2089 (N_2089,In_749,In_168);
nor U2090 (N_2090,In_231,In_936);
or U2091 (N_2091,In_365,In_611);
nand U2092 (N_2092,In_855,In_316);
and U2093 (N_2093,In_616,In_708);
nor U2094 (N_2094,In_350,In_982);
and U2095 (N_2095,In_817,In_878);
xnor U2096 (N_2096,In_863,In_773);
nor U2097 (N_2097,In_471,In_490);
or U2098 (N_2098,In_883,In_598);
nand U2099 (N_2099,In_403,In_415);
nand U2100 (N_2100,In_824,In_545);
nand U2101 (N_2101,In_649,In_773);
nor U2102 (N_2102,In_330,In_62);
nand U2103 (N_2103,In_738,In_280);
and U2104 (N_2104,In_999,In_859);
nor U2105 (N_2105,In_927,In_846);
nor U2106 (N_2106,In_981,In_400);
or U2107 (N_2107,In_488,In_733);
or U2108 (N_2108,In_510,In_875);
nand U2109 (N_2109,In_373,In_512);
or U2110 (N_2110,In_93,In_667);
or U2111 (N_2111,In_473,In_219);
nand U2112 (N_2112,In_732,In_155);
xnor U2113 (N_2113,In_382,In_41);
and U2114 (N_2114,In_501,In_893);
xnor U2115 (N_2115,In_889,In_76);
and U2116 (N_2116,In_39,In_387);
nor U2117 (N_2117,In_313,In_592);
or U2118 (N_2118,In_740,In_555);
nand U2119 (N_2119,In_593,In_65);
and U2120 (N_2120,In_980,In_818);
or U2121 (N_2121,In_726,In_165);
nor U2122 (N_2122,In_67,In_897);
nand U2123 (N_2123,In_896,In_647);
or U2124 (N_2124,In_988,In_95);
nor U2125 (N_2125,In_938,In_404);
and U2126 (N_2126,In_502,In_163);
nor U2127 (N_2127,In_124,In_685);
nand U2128 (N_2128,In_561,In_454);
nand U2129 (N_2129,In_494,In_354);
and U2130 (N_2130,In_13,In_771);
nand U2131 (N_2131,In_474,In_304);
and U2132 (N_2132,In_840,In_716);
nor U2133 (N_2133,In_395,In_239);
nor U2134 (N_2134,In_246,In_25);
nor U2135 (N_2135,In_178,In_363);
nor U2136 (N_2136,In_982,In_879);
and U2137 (N_2137,In_337,In_686);
or U2138 (N_2138,In_922,In_752);
or U2139 (N_2139,In_609,In_243);
xor U2140 (N_2140,In_931,In_991);
nand U2141 (N_2141,In_485,In_249);
or U2142 (N_2142,In_224,In_653);
or U2143 (N_2143,In_586,In_778);
nand U2144 (N_2144,In_157,In_31);
nor U2145 (N_2145,In_775,In_326);
xnor U2146 (N_2146,In_698,In_531);
and U2147 (N_2147,In_374,In_660);
xor U2148 (N_2148,In_608,In_247);
or U2149 (N_2149,In_165,In_608);
nor U2150 (N_2150,In_405,In_241);
and U2151 (N_2151,In_186,In_314);
nor U2152 (N_2152,In_866,In_302);
or U2153 (N_2153,In_252,In_541);
nor U2154 (N_2154,In_92,In_735);
nor U2155 (N_2155,In_461,In_276);
xor U2156 (N_2156,In_239,In_959);
nor U2157 (N_2157,In_458,In_427);
and U2158 (N_2158,In_945,In_466);
xnor U2159 (N_2159,In_448,In_581);
nand U2160 (N_2160,In_270,In_899);
or U2161 (N_2161,In_76,In_200);
nor U2162 (N_2162,In_14,In_153);
and U2163 (N_2163,In_727,In_48);
nand U2164 (N_2164,In_295,In_640);
or U2165 (N_2165,In_613,In_520);
nor U2166 (N_2166,In_459,In_959);
nor U2167 (N_2167,In_653,In_650);
and U2168 (N_2168,In_965,In_203);
nand U2169 (N_2169,In_212,In_101);
or U2170 (N_2170,In_864,In_528);
nand U2171 (N_2171,In_877,In_855);
or U2172 (N_2172,In_473,In_380);
nor U2173 (N_2173,In_380,In_746);
or U2174 (N_2174,In_393,In_156);
and U2175 (N_2175,In_31,In_914);
nor U2176 (N_2176,In_272,In_632);
and U2177 (N_2177,In_57,In_1);
nand U2178 (N_2178,In_63,In_317);
and U2179 (N_2179,In_282,In_993);
or U2180 (N_2180,In_683,In_886);
or U2181 (N_2181,In_753,In_487);
nand U2182 (N_2182,In_809,In_123);
or U2183 (N_2183,In_777,In_925);
xor U2184 (N_2184,In_862,In_162);
and U2185 (N_2185,In_402,In_293);
and U2186 (N_2186,In_796,In_227);
nand U2187 (N_2187,In_689,In_478);
and U2188 (N_2188,In_694,In_407);
or U2189 (N_2189,In_191,In_965);
or U2190 (N_2190,In_438,In_953);
or U2191 (N_2191,In_276,In_144);
nor U2192 (N_2192,In_469,In_124);
nand U2193 (N_2193,In_123,In_705);
and U2194 (N_2194,In_996,In_931);
or U2195 (N_2195,In_471,In_37);
and U2196 (N_2196,In_135,In_688);
nor U2197 (N_2197,In_500,In_70);
nor U2198 (N_2198,In_759,In_533);
nand U2199 (N_2199,In_551,In_891);
nor U2200 (N_2200,In_31,In_108);
nor U2201 (N_2201,In_344,In_368);
nor U2202 (N_2202,In_357,In_892);
xor U2203 (N_2203,In_68,In_547);
nor U2204 (N_2204,In_676,In_891);
nand U2205 (N_2205,In_113,In_946);
nor U2206 (N_2206,In_539,In_649);
nor U2207 (N_2207,In_39,In_948);
and U2208 (N_2208,In_152,In_875);
xor U2209 (N_2209,In_419,In_980);
and U2210 (N_2210,In_670,In_556);
or U2211 (N_2211,In_396,In_642);
and U2212 (N_2212,In_73,In_937);
xnor U2213 (N_2213,In_827,In_459);
xor U2214 (N_2214,In_747,In_142);
or U2215 (N_2215,In_706,In_560);
nand U2216 (N_2216,In_738,In_143);
nor U2217 (N_2217,In_270,In_514);
or U2218 (N_2218,In_80,In_989);
nand U2219 (N_2219,In_201,In_771);
or U2220 (N_2220,In_196,In_591);
nor U2221 (N_2221,In_397,In_424);
nand U2222 (N_2222,In_488,In_327);
or U2223 (N_2223,In_821,In_726);
nand U2224 (N_2224,In_836,In_112);
nor U2225 (N_2225,In_706,In_781);
nand U2226 (N_2226,In_24,In_393);
and U2227 (N_2227,In_819,In_926);
nor U2228 (N_2228,In_80,In_506);
and U2229 (N_2229,In_206,In_502);
or U2230 (N_2230,In_987,In_31);
xor U2231 (N_2231,In_834,In_194);
nand U2232 (N_2232,In_950,In_607);
nand U2233 (N_2233,In_854,In_307);
or U2234 (N_2234,In_89,In_430);
and U2235 (N_2235,In_792,In_103);
nand U2236 (N_2236,In_789,In_176);
nor U2237 (N_2237,In_875,In_364);
nand U2238 (N_2238,In_383,In_516);
and U2239 (N_2239,In_667,In_686);
or U2240 (N_2240,In_639,In_650);
and U2241 (N_2241,In_742,In_322);
xnor U2242 (N_2242,In_320,In_427);
nor U2243 (N_2243,In_376,In_24);
nand U2244 (N_2244,In_995,In_871);
and U2245 (N_2245,In_637,In_227);
or U2246 (N_2246,In_593,In_937);
or U2247 (N_2247,In_870,In_966);
xnor U2248 (N_2248,In_732,In_815);
or U2249 (N_2249,In_416,In_945);
or U2250 (N_2250,In_344,In_631);
or U2251 (N_2251,In_623,In_372);
nor U2252 (N_2252,In_152,In_974);
and U2253 (N_2253,In_369,In_188);
nand U2254 (N_2254,In_845,In_345);
and U2255 (N_2255,In_51,In_97);
nor U2256 (N_2256,In_865,In_2);
nor U2257 (N_2257,In_597,In_687);
or U2258 (N_2258,In_928,In_484);
and U2259 (N_2259,In_245,In_152);
nand U2260 (N_2260,In_745,In_113);
and U2261 (N_2261,In_488,In_907);
nor U2262 (N_2262,In_125,In_780);
nor U2263 (N_2263,In_983,In_601);
xnor U2264 (N_2264,In_646,In_474);
or U2265 (N_2265,In_269,In_376);
nand U2266 (N_2266,In_401,In_282);
or U2267 (N_2267,In_201,In_931);
nor U2268 (N_2268,In_665,In_852);
and U2269 (N_2269,In_368,In_216);
nor U2270 (N_2270,In_146,In_538);
xnor U2271 (N_2271,In_868,In_558);
and U2272 (N_2272,In_627,In_243);
nor U2273 (N_2273,In_965,In_769);
or U2274 (N_2274,In_215,In_610);
nor U2275 (N_2275,In_517,In_621);
nand U2276 (N_2276,In_438,In_120);
and U2277 (N_2277,In_522,In_12);
and U2278 (N_2278,In_661,In_128);
and U2279 (N_2279,In_107,In_100);
nand U2280 (N_2280,In_782,In_741);
nor U2281 (N_2281,In_312,In_126);
or U2282 (N_2282,In_918,In_916);
xor U2283 (N_2283,In_127,In_531);
or U2284 (N_2284,In_615,In_196);
nand U2285 (N_2285,In_503,In_746);
nor U2286 (N_2286,In_321,In_437);
nor U2287 (N_2287,In_843,In_435);
nand U2288 (N_2288,In_173,In_601);
and U2289 (N_2289,In_530,In_344);
and U2290 (N_2290,In_538,In_777);
nand U2291 (N_2291,In_633,In_892);
nor U2292 (N_2292,In_311,In_972);
nor U2293 (N_2293,In_353,In_711);
nand U2294 (N_2294,In_919,In_925);
or U2295 (N_2295,In_398,In_403);
and U2296 (N_2296,In_150,In_535);
nand U2297 (N_2297,In_271,In_234);
nand U2298 (N_2298,In_450,In_166);
or U2299 (N_2299,In_524,In_295);
nand U2300 (N_2300,In_757,In_607);
nor U2301 (N_2301,In_863,In_771);
or U2302 (N_2302,In_489,In_27);
nor U2303 (N_2303,In_966,In_386);
nand U2304 (N_2304,In_639,In_469);
nand U2305 (N_2305,In_114,In_275);
xnor U2306 (N_2306,In_187,In_329);
and U2307 (N_2307,In_743,In_325);
nor U2308 (N_2308,In_30,In_382);
nor U2309 (N_2309,In_947,In_172);
nor U2310 (N_2310,In_746,In_150);
or U2311 (N_2311,In_714,In_25);
nand U2312 (N_2312,In_964,In_261);
nor U2313 (N_2313,In_692,In_912);
or U2314 (N_2314,In_425,In_18);
and U2315 (N_2315,In_866,In_748);
xor U2316 (N_2316,In_820,In_862);
xor U2317 (N_2317,In_75,In_724);
or U2318 (N_2318,In_459,In_702);
and U2319 (N_2319,In_604,In_131);
and U2320 (N_2320,In_592,In_295);
or U2321 (N_2321,In_762,In_42);
and U2322 (N_2322,In_796,In_612);
and U2323 (N_2323,In_607,In_158);
and U2324 (N_2324,In_741,In_720);
and U2325 (N_2325,In_152,In_752);
nand U2326 (N_2326,In_268,In_410);
nand U2327 (N_2327,In_339,In_458);
nand U2328 (N_2328,In_29,In_199);
or U2329 (N_2329,In_48,In_626);
nor U2330 (N_2330,In_29,In_251);
or U2331 (N_2331,In_351,In_211);
and U2332 (N_2332,In_634,In_97);
nand U2333 (N_2333,In_385,In_752);
xor U2334 (N_2334,In_969,In_84);
or U2335 (N_2335,In_596,In_969);
nand U2336 (N_2336,In_452,In_447);
nor U2337 (N_2337,In_196,In_550);
nor U2338 (N_2338,In_184,In_526);
nor U2339 (N_2339,In_194,In_526);
and U2340 (N_2340,In_569,In_654);
and U2341 (N_2341,In_238,In_703);
nor U2342 (N_2342,In_351,In_910);
and U2343 (N_2343,In_617,In_352);
and U2344 (N_2344,In_454,In_325);
and U2345 (N_2345,In_674,In_759);
and U2346 (N_2346,In_346,In_331);
xnor U2347 (N_2347,In_315,In_271);
nor U2348 (N_2348,In_937,In_259);
or U2349 (N_2349,In_199,In_103);
or U2350 (N_2350,In_604,In_294);
or U2351 (N_2351,In_984,In_27);
nor U2352 (N_2352,In_69,In_607);
or U2353 (N_2353,In_216,In_395);
and U2354 (N_2354,In_764,In_294);
nand U2355 (N_2355,In_264,In_849);
and U2356 (N_2356,In_136,In_523);
nor U2357 (N_2357,In_817,In_16);
nor U2358 (N_2358,In_423,In_674);
nand U2359 (N_2359,In_128,In_950);
or U2360 (N_2360,In_653,In_323);
or U2361 (N_2361,In_650,In_418);
nand U2362 (N_2362,In_40,In_12);
nor U2363 (N_2363,In_594,In_955);
and U2364 (N_2364,In_735,In_174);
xor U2365 (N_2365,In_730,In_109);
nor U2366 (N_2366,In_375,In_449);
and U2367 (N_2367,In_235,In_483);
and U2368 (N_2368,In_182,In_117);
nand U2369 (N_2369,In_624,In_761);
nand U2370 (N_2370,In_951,In_648);
and U2371 (N_2371,In_192,In_936);
or U2372 (N_2372,In_332,In_914);
or U2373 (N_2373,In_828,In_163);
nor U2374 (N_2374,In_853,In_240);
nand U2375 (N_2375,In_784,In_432);
and U2376 (N_2376,In_871,In_161);
or U2377 (N_2377,In_899,In_369);
nor U2378 (N_2378,In_540,In_822);
or U2379 (N_2379,In_945,In_538);
nor U2380 (N_2380,In_135,In_498);
and U2381 (N_2381,In_59,In_157);
nor U2382 (N_2382,In_284,In_989);
xnor U2383 (N_2383,In_114,In_895);
or U2384 (N_2384,In_875,In_291);
or U2385 (N_2385,In_565,In_478);
and U2386 (N_2386,In_377,In_64);
nand U2387 (N_2387,In_971,In_309);
or U2388 (N_2388,In_20,In_936);
and U2389 (N_2389,In_998,In_632);
or U2390 (N_2390,In_87,In_236);
and U2391 (N_2391,In_434,In_148);
nand U2392 (N_2392,In_928,In_988);
nor U2393 (N_2393,In_184,In_463);
and U2394 (N_2394,In_248,In_311);
nand U2395 (N_2395,In_78,In_593);
xor U2396 (N_2396,In_74,In_670);
nor U2397 (N_2397,In_230,In_384);
nand U2398 (N_2398,In_459,In_635);
or U2399 (N_2399,In_918,In_619);
xor U2400 (N_2400,In_400,In_858);
and U2401 (N_2401,In_674,In_634);
and U2402 (N_2402,In_610,In_945);
or U2403 (N_2403,In_252,In_543);
nor U2404 (N_2404,In_494,In_83);
or U2405 (N_2405,In_903,In_101);
nor U2406 (N_2406,In_236,In_27);
nand U2407 (N_2407,In_364,In_836);
nor U2408 (N_2408,In_693,In_120);
xnor U2409 (N_2409,In_767,In_159);
xnor U2410 (N_2410,In_754,In_464);
xnor U2411 (N_2411,In_370,In_761);
or U2412 (N_2412,In_650,In_427);
nor U2413 (N_2413,In_90,In_591);
and U2414 (N_2414,In_183,In_141);
nor U2415 (N_2415,In_396,In_289);
or U2416 (N_2416,In_610,In_736);
and U2417 (N_2417,In_319,In_602);
nor U2418 (N_2418,In_518,In_332);
and U2419 (N_2419,In_522,In_26);
and U2420 (N_2420,In_460,In_471);
nor U2421 (N_2421,In_701,In_971);
and U2422 (N_2422,In_277,In_549);
nand U2423 (N_2423,In_91,In_797);
and U2424 (N_2424,In_170,In_324);
nand U2425 (N_2425,In_685,In_193);
or U2426 (N_2426,In_739,In_987);
or U2427 (N_2427,In_274,In_739);
and U2428 (N_2428,In_565,In_614);
nor U2429 (N_2429,In_285,In_333);
or U2430 (N_2430,In_422,In_490);
or U2431 (N_2431,In_701,In_989);
or U2432 (N_2432,In_693,In_327);
and U2433 (N_2433,In_840,In_934);
nor U2434 (N_2434,In_529,In_850);
nand U2435 (N_2435,In_107,In_353);
nor U2436 (N_2436,In_683,In_887);
xor U2437 (N_2437,In_453,In_279);
and U2438 (N_2438,In_740,In_587);
and U2439 (N_2439,In_862,In_928);
xor U2440 (N_2440,In_972,In_101);
nand U2441 (N_2441,In_683,In_688);
and U2442 (N_2442,In_949,In_781);
and U2443 (N_2443,In_853,In_300);
nor U2444 (N_2444,In_524,In_245);
or U2445 (N_2445,In_832,In_406);
nor U2446 (N_2446,In_209,In_314);
nand U2447 (N_2447,In_159,In_87);
and U2448 (N_2448,In_959,In_26);
or U2449 (N_2449,In_21,In_49);
nand U2450 (N_2450,In_510,In_376);
or U2451 (N_2451,In_809,In_898);
nor U2452 (N_2452,In_541,In_168);
nand U2453 (N_2453,In_993,In_288);
or U2454 (N_2454,In_262,In_609);
or U2455 (N_2455,In_970,In_957);
nand U2456 (N_2456,In_61,In_834);
and U2457 (N_2457,In_348,In_269);
nor U2458 (N_2458,In_42,In_278);
and U2459 (N_2459,In_517,In_120);
nand U2460 (N_2460,In_896,In_877);
or U2461 (N_2461,In_832,In_677);
xnor U2462 (N_2462,In_416,In_71);
nor U2463 (N_2463,In_936,In_877);
nand U2464 (N_2464,In_374,In_655);
and U2465 (N_2465,In_999,In_167);
and U2466 (N_2466,In_518,In_806);
or U2467 (N_2467,In_965,In_848);
nand U2468 (N_2468,In_703,In_802);
nor U2469 (N_2469,In_988,In_617);
nand U2470 (N_2470,In_806,In_971);
or U2471 (N_2471,In_972,In_919);
nand U2472 (N_2472,In_829,In_692);
nand U2473 (N_2473,In_375,In_127);
and U2474 (N_2474,In_362,In_608);
and U2475 (N_2475,In_460,In_85);
nor U2476 (N_2476,In_897,In_923);
and U2477 (N_2477,In_542,In_945);
nand U2478 (N_2478,In_470,In_770);
or U2479 (N_2479,In_308,In_452);
nor U2480 (N_2480,In_292,In_912);
nand U2481 (N_2481,In_751,In_676);
nand U2482 (N_2482,In_880,In_431);
and U2483 (N_2483,In_193,In_872);
and U2484 (N_2484,In_973,In_514);
and U2485 (N_2485,In_732,In_461);
or U2486 (N_2486,In_504,In_220);
nor U2487 (N_2487,In_576,In_571);
or U2488 (N_2488,In_142,In_666);
nand U2489 (N_2489,In_637,In_986);
and U2490 (N_2490,In_971,In_739);
and U2491 (N_2491,In_898,In_172);
xnor U2492 (N_2492,In_199,In_496);
and U2493 (N_2493,In_800,In_219);
or U2494 (N_2494,In_531,In_847);
or U2495 (N_2495,In_106,In_840);
nor U2496 (N_2496,In_318,In_67);
nor U2497 (N_2497,In_41,In_520);
xor U2498 (N_2498,In_728,In_158);
or U2499 (N_2499,In_344,In_415);
and U2500 (N_2500,In_908,In_873);
and U2501 (N_2501,In_633,In_508);
nor U2502 (N_2502,In_596,In_804);
xnor U2503 (N_2503,In_363,In_767);
nor U2504 (N_2504,In_211,In_966);
xnor U2505 (N_2505,In_477,In_313);
xor U2506 (N_2506,In_731,In_733);
nand U2507 (N_2507,In_652,In_178);
xnor U2508 (N_2508,In_226,In_602);
nor U2509 (N_2509,In_307,In_638);
nor U2510 (N_2510,In_989,In_168);
and U2511 (N_2511,In_329,In_124);
xnor U2512 (N_2512,In_473,In_699);
and U2513 (N_2513,In_882,In_907);
or U2514 (N_2514,In_793,In_688);
and U2515 (N_2515,In_446,In_303);
nor U2516 (N_2516,In_729,In_478);
nand U2517 (N_2517,In_394,In_369);
or U2518 (N_2518,In_772,In_242);
and U2519 (N_2519,In_303,In_437);
or U2520 (N_2520,In_722,In_521);
xnor U2521 (N_2521,In_407,In_711);
or U2522 (N_2522,In_491,In_352);
nor U2523 (N_2523,In_371,In_817);
nor U2524 (N_2524,In_324,In_334);
xnor U2525 (N_2525,In_372,In_760);
xor U2526 (N_2526,In_863,In_522);
nand U2527 (N_2527,In_283,In_644);
or U2528 (N_2528,In_80,In_823);
nand U2529 (N_2529,In_235,In_890);
and U2530 (N_2530,In_667,In_169);
and U2531 (N_2531,In_292,In_762);
and U2532 (N_2532,In_15,In_299);
nand U2533 (N_2533,In_984,In_521);
or U2534 (N_2534,In_974,In_76);
or U2535 (N_2535,In_500,In_893);
nor U2536 (N_2536,In_104,In_773);
nand U2537 (N_2537,In_421,In_598);
and U2538 (N_2538,In_574,In_411);
or U2539 (N_2539,In_438,In_937);
nand U2540 (N_2540,In_567,In_394);
and U2541 (N_2541,In_377,In_217);
or U2542 (N_2542,In_475,In_795);
nor U2543 (N_2543,In_685,In_946);
and U2544 (N_2544,In_940,In_842);
and U2545 (N_2545,In_112,In_555);
nor U2546 (N_2546,In_539,In_259);
and U2547 (N_2547,In_239,In_740);
or U2548 (N_2548,In_485,In_91);
and U2549 (N_2549,In_360,In_825);
nand U2550 (N_2550,In_812,In_156);
and U2551 (N_2551,In_261,In_789);
or U2552 (N_2552,In_852,In_188);
nand U2553 (N_2553,In_690,In_767);
nor U2554 (N_2554,In_387,In_312);
or U2555 (N_2555,In_19,In_431);
and U2556 (N_2556,In_559,In_106);
or U2557 (N_2557,In_822,In_316);
xnor U2558 (N_2558,In_589,In_802);
xnor U2559 (N_2559,In_719,In_564);
or U2560 (N_2560,In_929,In_992);
and U2561 (N_2561,In_955,In_694);
or U2562 (N_2562,In_851,In_101);
and U2563 (N_2563,In_664,In_454);
nor U2564 (N_2564,In_262,In_507);
or U2565 (N_2565,In_345,In_77);
and U2566 (N_2566,In_746,In_737);
nand U2567 (N_2567,In_571,In_808);
nand U2568 (N_2568,In_916,In_553);
and U2569 (N_2569,In_597,In_84);
nor U2570 (N_2570,In_8,In_391);
nor U2571 (N_2571,In_578,In_176);
nand U2572 (N_2572,In_936,In_433);
or U2573 (N_2573,In_866,In_503);
xnor U2574 (N_2574,In_557,In_116);
nand U2575 (N_2575,In_518,In_581);
or U2576 (N_2576,In_223,In_759);
or U2577 (N_2577,In_53,In_488);
or U2578 (N_2578,In_822,In_76);
nand U2579 (N_2579,In_637,In_831);
or U2580 (N_2580,In_977,In_856);
nor U2581 (N_2581,In_249,In_457);
nor U2582 (N_2582,In_212,In_432);
xnor U2583 (N_2583,In_783,In_779);
nor U2584 (N_2584,In_11,In_47);
or U2585 (N_2585,In_174,In_660);
or U2586 (N_2586,In_804,In_148);
and U2587 (N_2587,In_168,In_379);
or U2588 (N_2588,In_784,In_174);
nand U2589 (N_2589,In_376,In_849);
nand U2590 (N_2590,In_802,In_496);
nor U2591 (N_2591,In_147,In_184);
or U2592 (N_2592,In_988,In_421);
xor U2593 (N_2593,In_806,In_916);
or U2594 (N_2594,In_165,In_442);
or U2595 (N_2595,In_64,In_46);
xor U2596 (N_2596,In_533,In_448);
and U2597 (N_2597,In_91,In_185);
nand U2598 (N_2598,In_661,In_841);
nor U2599 (N_2599,In_753,In_314);
and U2600 (N_2600,In_663,In_572);
nand U2601 (N_2601,In_640,In_308);
nor U2602 (N_2602,In_268,In_879);
and U2603 (N_2603,In_781,In_277);
nor U2604 (N_2604,In_268,In_463);
or U2605 (N_2605,In_958,In_907);
xnor U2606 (N_2606,In_373,In_243);
nand U2607 (N_2607,In_969,In_722);
nor U2608 (N_2608,In_166,In_643);
and U2609 (N_2609,In_522,In_647);
nand U2610 (N_2610,In_407,In_684);
nand U2611 (N_2611,In_792,In_55);
or U2612 (N_2612,In_829,In_214);
nor U2613 (N_2613,In_447,In_213);
xnor U2614 (N_2614,In_408,In_946);
nor U2615 (N_2615,In_415,In_40);
nand U2616 (N_2616,In_20,In_296);
xnor U2617 (N_2617,In_289,In_520);
xnor U2618 (N_2618,In_421,In_819);
xor U2619 (N_2619,In_344,In_587);
xor U2620 (N_2620,In_749,In_336);
nor U2621 (N_2621,In_529,In_45);
nor U2622 (N_2622,In_112,In_443);
nand U2623 (N_2623,In_226,In_967);
nor U2624 (N_2624,In_550,In_976);
or U2625 (N_2625,In_806,In_794);
nor U2626 (N_2626,In_969,In_55);
nor U2627 (N_2627,In_472,In_245);
nor U2628 (N_2628,In_399,In_798);
or U2629 (N_2629,In_352,In_631);
nand U2630 (N_2630,In_770,In_793);
xnor U2631 (N_2631,In_827,In_808);
nand U2632 (N_2632,In_746,In_327);
or U2633 (N_2633,In_706,In_76);
and U2634 (N_2634,In_835,In_626);
or U2635 (N_2635,In_656,In_281);
nor U2636 (N_2636,In_347,In_699);
or U2637 (N_2637,In_392,In_264);
or U2638 (N_2638,In_961,In_824);
nor U2639 (N_2639,In_954,In_442);
and U2640 (N_2640,In_984,In_724);
and U2641 (N_2641,In_400,In_63);
xnor U2642 (N_2642,In_103,In_427);
and U2643 (N_2643,In_54,In_583);
nand U2644 (N_2644,In_109,In_223);
and U2645 (N_2645,In_584,In_32);
nor U2646 (N_2646,In_688,In_628);
and U2647 (N_2647,In_638,In_316);
and U2648 (N_2648,In_116,In_387);
xnor U2649 (N_2649,In_375,In_276);
nand U2650 (N_2650,In_824,In_496);
or U2651 (N_2651,In_39,In_824);
and U2652 (N_2652,In_598,In_131);
xor U2653 (N_2653,In_400,In_282);
or U2654 (N_2654,In_327,In_918);
xor U2655 (N_2655,In_523,In_782);
nand U2656 (N_2656,In_987,In_221);
nand U2657 (N_2657,In_759,In_128);
xor U2658 (N_2658,In_141,In_699);
or U2659 (N_2659,In_892,In_706);
nor U2660 (N_2660,In_204,In_538);
nand U2661 (N_2661,In_501,In_734);
or U2662 (N_2662,In_737,In_361);
or U2663 (N_2663,In_842,In_598);
nor U2664 (N_2664,In_886,In_329);
xnor U2665 (N_2665,In_804,In_406);
nor U2666 (N_2666,In_230,In_834);
nor U2667 (N_2667,In_225,In_249);
or U2668 (N_2668,In_406,In_313);
nor U2669 (N_2669,In_56,In_907);
nor U2670 (N_2670,In_931,In_414);
or U2671 (N_2671,In_739,In_132);
or U2672 (N_2672,In_743,In_695);
xor U2673 (N_2673,In_44,In_440);
and U2674 (N_2674,In_816,In_27);
or U2675 (N_2675,In_546,In_117);
nand U2676 (N_2676,In_553,In_877);
or U2677 (N_2677,In_765,In_298);
and U2678 (N_2678,In_29,In_296);
nor U2679 (N_2679,In_423,In_440);
and U2680 (N_2680,In_944,In_504);
nor U2681 (N_2681,In_57,In_542);
or U2682 (N_2682,In_834,In_240);
nor U2683 (N_2683,In_65,In_292);
nand U2684 (N_2684,In_636,In_570);
or U2685 (N_2685,In_416,In_732);
nand U2686 (N_2686,In_593,In_391);
nand U2687 (N_2687,In_803,In_561);
nor U2688 (N_2688,In_862,In_522);
xnor U2689 (N_2689,In_816,In_585);
nand U2690 (N_2690,In_905,In_548);
or U2691 (N_2691,In_247,In_986);
nor U2692 (N_2692,In_561,In_460);
nor U2693 (N_2693,In_913,In_72);
nand U2694 (N_2694,In_907,In_525);
xnor U2695 (N_2695,In_859,In_230);
nand U2696 (N_2696,In_400,In_448);
nand U2697 (N_2697,In_931,In_391);
or U2698 (N_2698,In_945,In_137);
or U2699 (N_2699,In_990,In_904);
or U2700 (N_2700,In_558,In_482);
or U2701 (N_2701,In_779,In_404);
and U2702 (N_2702,In_133,In_273);
nand U2703 (N_2703,In_626,In_496);
or U2704 (N_2704,In_382,In_322);
or U2705 (N_2705,In_426,In_614);
nand U2706 (N_2706,In_7,In_261);
or U2707 (N_2707,In_308,In_335);
nand U2708 (N_2708,In_887,In_650);
or U2709 (N_2709,In_743,In_923);
nor U2710 (N_2710,In_677,In_603);
or U2711 (N_2711,In_927,In_144);
and U2712 (N_2712,In_199,In_701);
and U2713 (N_2713,In_482,In_810);
and U2714 (N_2714,In_872,In_508);
nor U2715 (N_2715,In_130,In_774);
nand U2716 (N_2716,In_163,In_562);
nand U2717 (N_2717,In_186,In_716);
or U2718 (N_2718,In_340,In_8);
nand U2719 (N_2719,In_461,In_588);
or U2720 (N_2720,In_453,In_94);
nor U2721 (N_2721,In_95,In_551);
and U2722 (N_2722,In_857,In_511);
xnor U2723 (N_2723,In_725,In_84);
nor U2724 (N_2724,In_291,In_812);
nor U2725 (N_2725,In_856,In_764);
and U2726 (N_2726,In_962,In_74);
nor U2727 (N_2727,In_843,In_574);
nor U2728 (N_2728,In_81,In_378);
or U2729 (N_2729,In_621,In_883);
or U2730 (N_2730,In_443,In_740);
and U2731 (N_2731,In_63,In_234);
nor U2732 (N_2732,In_552,In_89);
and U2733 (N_2733,In_190,In_768);
nand U2734 (N_2734,In_618,In_825);
and U2735 (N_2735,In_386,In_930);
nor U2736 (N_2736,In_53,In_714);
nor U2737 (N_2737,In_682,In_888);
xor U2738 (N_2738,In_701,In_948);
nand U2739 (N_2739,In_595,In_913);
nor U2740 (N_2740,In_662,In_835);
and U2741 (N_2741,In_725,In_291);
nor U2742 (N_2742,In_387,In_383);
and U2743 (N_2743,In_45,In_678);
nor U2744 (N_2744,In_692,In_753);
nor U2745 (N_2745,In_308,In_221);
nor U2746 (N_2746,In_851,In_343);
and U2747 (N_2747,In_651,In_683);
nand U2748 (N_2748,In_141,In_126);
and U2749 (N_2749,In_279,In_328);
or U2750 (N_2750,In_685,In_144);
and U2751 (N_2751,In_904,In_144);
nand U2752 (N_2752,In_205,In_656);
or U2753 (N_2753,In_956,In_970);
nand U2754 (N_2754,In_629,In_368);
or U2755 (N_2755,In_609,In_628);
nand U2756 (N_2756,In_46,In_712);
nand U2757 (N_2757,In_325,In_312);
or U2758 (N_2758,In_942,In_101);
nand U2759 (N_2759,In_833,In_617);
nor U2760 (N_2760,In_231,In_120);
nor U2761 (N_2761,In_269,In_766);
xor U2762 (N_2762,In_262,In_663);
nor U2763 (N_2763,In_576,In_218);
xnor U2764 (N_2764,In_713,In_287);
or U2765 (N_2765,In_484,In_306);
and U2766 (N_2766,In_874,In_710);
xor U2767 (N_2767,In_89,In_102);
or U2768 (N_2768,In_250,In_634);
and U2769 (N_2769,In_13,In_856);
or U2770 (N_2770,In_685,In_389);
or U2771 (N_2771,In_199,In_533);
nand U2772 (N_2772,In_923,In_292);
or U2773 (N_2773,In_69,In_726);
xor U2774 (N_2774,In_574,In_735);
or U2775 (N_2775,In_870,In_309);
nand U2776 (N_2776,In_192,In_288);
nand U2777 (N_2777,In_68,In_924);
nand U2778 (N_2778,In_431,In_732);
and U2779 (N_2779,In_197,In_320);
xor U2780 (N_2780,In_366,In_424);
or U2781 (N_2781,In_308,In_874);
nor U2782 (N_2782,In_482,In_883);
nor U2783 (N_2783,In_240,In_523);
nand U2784 (N_2784,In_463,In_68);
and U2785 (N_2785,In_601,In_312);
or U2786 (N_2786,In_596,In_221);
nand U2787 (N_2787,In_814,In_608);
and U2788 (N_2788,In_921,In_116);
nand U2789 (N_2789,In_877,In_115);
or U2790 (N_2790,In_487,In_418);
nand U2791 (N_2791,In_156,In_671);
nand U2792 (N_2792,In_726,In_86);
nand U2793 (N_2793,In_570,In_993);
or U2794 (N_2794,In_730,In_539);
or U2795 (N_2795,In_370,In_526);
and U2796 (N_2796,In_461,In_584);
nand U2797 (N_2797,In_542,In_933);
and U2798 (N_2798,In_436,In_552);
nand U2799 (N_2799,In_688,In_386);
nor U2800 (N_2800,In_924,In_397);
and U2801 (N_2801,In_29,In_412);
nand U2802 (N_2802,In_149,In_774);
nor U2803 (N_2803,In_679,In_961);
nor U2804 (N_2804,In_103,In_797);
and U2805 (N_2805,In_630,In_789);
nand U2806 (N_2806,In_238,In_14);
nor U2807 (N_2807,In_143,In_923);
and U2808 (N_2808,In_807,In_306);
nand U2809 (N_2809,In_425,In_213);
or U2810 (N_2810,In_268,In_924);
nand U2811 (N_2811,In_467,In_852);
nor U2812 (N_2812,In_521,In_176);
nor U2813 (N_2813,In_15,In_206);
and U2814 (N_2814,In_858,In_278);
or U2815 (N_2815,In_988,In_370);
or U2816 (N_2816,In_215,In_756);
nor U2817 (N_2817,In_443,In_126);
xnor U2818 (N_2818,In_754,In_254);
or U2819 (N_2819,In_773,In_111);
and U2820 (N_2820,In_870,In_844);
nand U2821 (N_2821,In_540,In_108);
or U2822 (N_2822,In_642,In_669);
nand U2823 (N_2823,In_179,In_164);
nor U2824 (N_2824,In_406,In_476);
and U2825 (N_2825,In_489,In_951);
nor U2826 (N_2826,In_869,In_21);
nor U2827 (N_2827,In_811,In_229);
nand U2828 (N_2828,In_304,In_46);
nand U2829 (N_2829,In_909,In_557);
nand U2830 (N_2830,In_692,In_936);
nand U2831 (N_2831,In_360,In_752);
nor U2832 (N_2832,In_47,In_871);
nand U2833 (N_2833,In_892,In_971);
or U2834 (N_2834,In_42,In_891);
or U2835 (N_2835,In_44,In_465);
nand U2836 (N_2836,In_310,In_127);
and U2837 (N_2837,In_666,In_626);
xor U2838 (N_2838,In_947,In_922);
nand U2839 (N_2839,In_520,In_837);
nor U2840 (N_2840,In_750,In_275);
or U2841 (N_2841,In_93,In_663);
nor U2842 (N_2842,In_877,In_387);
and U2843 (N_2843,In_692,In_687);
nor U2844 (N_2844,In_214,In_498);
and U2845 (N_2845,In_171,In_752);
nor U2846 (N_2846,In_100,In_649);
xor U2847 (N_2847,In_388,In_381);
xnor U2848 (N_2848,In_224,In_410);
and U2849 (N_2849,In_167,In_406);
nand U2850 (N_2850,In_262,In_852);
or U2851 (N_2851,In_128,In_590);
or U2852 (N_2852,In_639,In_296);
nand U2853 (N_2853,In_951,In_432);
nor U2854 (N_2854,In_690,In_95);
or U2855 (N_2855,In_794,In_580);
or U2856 (N_2856,In_942,In_555);
or U2857 (N_2857,In_726,In_236);
nor U2858 (N_2858,In_619,In_611);
and U2859 (N_2859,In_87,In_118);
or U2860 (N_2860,In_445,In_345);
and U2861 (N_2861,In_285,In_216);
or U2862 (N_2862,In_204,In_60);
or U2863 (N_2863,In_346,In_621);
xnor U2864 (N_2864,In_747,In_60);
nand U2865 (N_2865,In_155,In_564);
nor U2866 (N_2866,In_345,In_318);
nor U2867 (N_2867,In_612,In_509);
or U2868 (N_2868,In_707,In_180);
nand U2869 (N_2869,In_324,In_367);
xnor U2870 (N_2870,In_943,In_732);
or U2871 (N_2871,In_973,In_699);
or U2872 (N_2872,In_70,In_154);
and U2873 (N_2873,In_22,In_794);
nand U2874 (N_2874,In_133,In_637);
and U2875 (N_2875,In_797,In_663);
nor U2876 (N_2876,In_749,In_218);
nor U2877 (N_2877,In_17,In_801);
and U2878 (N_2878,In_220,In_875);
nor U2879 (N_2879,In_297,In_367);
nand U2880 (N_2880,In_542,In_317);
nor U2881 (N_2881,In_127,In_326);
nand U2882 (N_2882,In_686,In_84);
and U2883 (N_2883,In_755,In_438);
nand U2884 (N_2884,In_610,In_196);
xnor U2885 (N_2885,In_344,In_381);
or U2886 (N_2886,In_393,In_645);
nand U2887 (N_2887,In_782,In_525);
or U2888 (N_2888,In_799,In_693);
and U2889 (N_2889,In_373,In_166);
nor U2890 (N_2890,In_666,In_565);
and U2891 (N_2891,In_717,In_711);
xnor U2892 (N_2892,In_901,In_857);
or U2893 (N_2893,In_871,In_138);
and U2894 (N_2894,In_256,In_38);
and U2895 (N_2895,In_877,In_186);
or U2896 (N_2896,In_244,In_33);
nor U2897 (N_2897,In_380,In_399);
nor U2898 (N_2898,In_639,In_897);
and U2899 (N_2899,In_68,In_326);
and U2900 (N_2900,In_67,In_822);
and U2901 (N_2901,In_926,In_353);
nand U2902 (N_2902,In_547,In_71);
nor U2903 (N_2903,In_527,In_492);
or U2904 (N_2904,In_640,In_47);
nor U2905 (N_2905,In_432,In_164);
xnor U2906 (N_2906,In_39,In_637);
or U2907 (N_2907,In_949,In_888);
or U2908 (N_2908,In_111,In_618);
and U2909 (N_2909,In_804,In_990);
or U2910 (N_2910,In_334,In_368);
nand U2911 (N_2911,In_574,In_145);
and U2912 (N_2912,In_758,In_548);
xor U2913 (N_2913,In_150,In_660);
nand U2914 (N_2914,In_175,In_594);
and U2915 (N_2915,In_709,In_276);
nand U2916 (N_2916,In_225,In_619);
nand U2917 (N_2917,In_61,In_605);
nand U2918 (N_2918,In_947,In_145);
or U2919 (N_2919,In_504,In_616);
nor U2920 (N_2920,In_149,In_46);
nor U2921 (N_2921,In_41,In_476);
nor U2922 (N_2922,In_991,In_438);
nand U2923 (N_2923,In_596,In_400);
and U2924 (N_2924,In_131,In_588);
and U2925 (N_2925,In_315,In_287);
and U2926 (N_2926,In_268,In_790);
or U2927 (N_2927,In_318,In_757);
nand U2928 (N_2928,In_563,In_41);
xor U2929 (N_2929,In_657,In_351);
nor U2930 (N_2930,In_532,In_389);
and U2931 (N_2931,In_477,In_915);
nand U2932 (N_2932,In_326,In_975);
nor U2933 (N_2933,In_143,In_409);
nand U2934 (N_2934,In_622,In_379);
and U2935 (N_2935,In_170,In_616);
nand U2936 (N_2936,In_738,In_329);
and U2937 (N_2937,In_384,In_964);
and U2938 (N_2938,In_511,In_773);
nor U2939 (N_2939,In_69,In_12);
or U2940 (N_2940,In_866,In_342);
or U2941 (N_2941,In_587,In_155);
or U2942 (N_2942,In_684,In_419);
and U2943 (N_2943,In_386,In_692);
nor U2944 (N_2944,In_142,In_797);
and U2945 (N_2945,In_911,In_29);
and U2946 (N_2946,In_962,In_698);
xnor U2947 (N_2947,In_427,In_95);
xnor U2948 (N_2948,In_823,In_307);
xor U2949 (N_2949,In_665,In_48);
and U2950 (N_2950,In_544,In_196);
nor U2951 (N_2951,In_99,In_418);
and U2952 (N_2952,In_960,In_476);
nand U2953 (N_2953,In_456,In_450);
nor U2954 (N_2954,In_176,In_925);
or U2955 (N_2955,In_562,In_819);
nand U2956 (N_2956,In_617,In_82);
nand U2957 (N_2957,In_26,In_127);
xor U2958 (N_2958,In_61,In_798);
or U2959 (N_2959,In_107,In_499);
or U2960 (N_2960,In_517,In_72);
nand U2961 (N_2961,In_472,In_761);
xnor U2962 (N_2962,In_353,In_303);
or U2963 (N_2963,In_961,In_954);
nor U2964 (N_2964,In_704,In_150);
nand U2965 (N_2965,In_51,In_902);
nor U2966 (N_2966,In_473,In_264);
xor U2967 (N_2967,In_6,In_436);
nor U2968 (N_2968,In_511,In_907);
nor U2969 (N_2969,In_819,In_790);
nand U2970 (N_2970,In_51,In_235);
nand U2971 (N_2971,In_100,In_113);
or U2972 (N_2972,In_199,In_925);
nor U2973 (N_2973,In_618,In_136);
or U2974 (N_2974,In_374,In_714);
nor U2975 (N_2975,In_315,In_745);
nand U2976 (N_2976,In_671,In_227);
nor U2977 (N_2977,In_949,In_383);
and U2978 (N_2978,In_848,In_312);
nand U2979 (N_2979,In_839,In_490);
nor U2980 (N_2980,In_320,In_464);
xor U2981 (N_2981,In_537,In_61);
and U2982 (N_2982,In_911,In_825);
xnor U2983 (N_2983,In_41,In_284);
xor U2984 (N_2984,In_309,In_49);
xnor U2985 (N_2985,In_719,In_792);
xnor U2986 (N_2986,In_264,In_502);
nand U2987 (N_2987,In_855,In_458);
and U2988 (N_2988,In_5,In_144);
xor U2989 (N_2989,In_195,In_221);
nand U2990 (N_2990,In_161,In_501);
and U2991 (N_2991,In_410,In_56);
and U2992 (N_2992,In_270,In_331);
nand U2993 (N_2993,In_26,In_926);
or U2994 (N_2994,In_56,In_879);
nand U2995 (N_2995,In_457,In_83);
nand U2996 (N_2996,In_146,In_379);
nand U2997 (N_2997,In_452,In_685);
or U2998 (N_2998,In_621,In_484);
and U2999 (N_2999,In_554,In_706);
nor U3000 (N_3000,In_103,In_55);
nand U3001 (N_3001,In_964,In_556);
nand U3002 (N_3002,In_45,In_182);
nor U3003 (N_3003,In_705,In_631);
nor U3004 (N_3004,In_482,In_679);
xnor U3005 (N_3005,In_177,In_618);
and U3006 (N_3006,In_95,In_383);
xor U3007 (N_3007,In_328,In_870);
xor U3008 (N_3008,In_702,In_537);
nor U3009 (N_3009,In_129,In_152);
xor U3010 (N_3010,In_850,In_98);
xnor U3011 (N_3011,In_420,In_275);
xnor U3012 (N_3012,In_707,In_473);
nand U3013 (N_3013,In_704,In_523);
nor U3014 (N_3014,In_238,In_92);
nand U3015 (N_3015,In_192,In_744);
nor U3016 (N_3016,In_399,In_93);
or U3017 (N_3017,In_282,In_193);
nand U3018 (N_3018,In_979,In_418);
nand U3019 (N_3019,In_767,In_431);
xor U3020 (N_3020,In_672,In_752);
and U3021 (N_3021,In_56,In_79);
nand U3022 (N_3022,In_771,In_534);
and U3023 (N_3023,In_870,In_310);
nor U3024 (N_3024,In_42,In_274);
and U3025 (N_3025,In_738,In_444);
nand U3026 (N_3026,In_124,In_828);
and U3027 (N_3027,In_679,In_699);
nand U3028 (N_3028,In_398,In_680);
nor U3029 (N_3029,In_911,In_688);
nand U3030 (N_3030,In_167,In_399);
or U3031 (N_3031,In_838,In_835);
or U3032 (N_3032,In_25,In_84);
nor U3033 (N_3033,In_283,In_884);
or U3034 (N_3034,In_979,In_743);
nor U3035 (N_3035,In_854,In_558);
and U3036 (N_3036,In_969,In_311);
nor U3037 (N_3037,In_641,In_612);
xnor U3038 (N_3038,In_63,In_328);
nor U3039 (N_3039,In_639,In_286);
nor U3040 (N_3040,In_938,In_133);
and U3041 (N_3041,In_534,In_204);
or U3042 (N_3042,In_540,In_623);
xor U3043 (N_3043,In_274,In_877);
nor U3044 (N_3044,In_761,In_940);
xor U3045 (N_3045,In_951,In_75);
nor U3046 (N_3046,In_883,In_967);
and U3047 (N_3047,In_707,In_61);
nor U3048 (N_3048,In_538,In_43);
and U3049 (N_3049,In_713,In_597);
nand U3050 (N_3050,In_388,In_356);
nor U3051 (N_3051,In_189,In_24);
and U3052 (N_3052,In_781,In_325);
or U3053 (N_3053,In_180,In_965);
and U3054 (N_3054,In_580,In_953);
nand U3055 (N_3055,In_692,In_858);
or U3056 (N_3056,In_602,In_590);
and U3057 (N_3057,In_131,In_767);
xor U3058 (N_3058,In_148,In_432);
nor U3059 (N_3059,In_746,In_113);
nor U3060 (N_3060,In_940,In_751);
and U3061 (N_3061,In_291,In_621);
or U3062 (N_3062,In_746,In_473);
nor U3063 (N_3063,In_573,In_451);
nand U3064 (N_3064,In_978,In_507);
nand U3065 (N_3065,In_764,In_917);
xor U3066 (N_3066,In_83,In_831);
nor U3067 (N_3067,In_402,In_457);
or U3068 (N_3068,In_446,In_588);
and U3069 (N_3069,In_863,In_463);
xnor U3070 (N_3070,In_65,In_423);
nor U3071 (N_3071,In_377,In_676);
nand U3072 (N_3072,In_830,In_286);
or U3073 (N_3073,In_234,In_568);
xor U3074 (N_3074,In_680,In_103);
nor U3075 (N_3075,In_342,In_702);
or U3076 (N_3076,In_229,In_911);
or U3077 (N_3077,In_920,In_107);
xor U3078 (N_3078,In_753,In_899);
nand U3079 (N_3079,In_140,In_176);
and U3080 (N_3080,In_602,In_889);
xnor U3081 (N_3081,In_144,In_168);
xnor U3082 (N_3082,In_423,In_351);
nor U3083 (N_3083,In_133,In_970);
or U3084 (N_3084,In_646,In_498);
nand U3085 (N_3085,In_698,In_18);
and U3086 (N_3086,In_168,In_952);
and U3087 (N_3087,In_455,In_108);
xor U3088 (N_3088,In_194,In_818);
nand U3089 (N_3089,In_409,In_521);
nor U3090 (N_3090,In_182,In_377);
nand U3091 (N_3091,In_150,In_58);
and U3092 (N_3092,In_82,In_306);
or U3093 (N_3093,In_882,In_159);
nor U3094 (N_3094,In_93,In_814);
and U3095 (N_3095,In_525,In_727);
nor U3096 (N_3096,In_137,In_160);
nor U3097 (N_3097,In_905,In_908);
nand U3098 (N_3098,In_941,In_784);
nor U3099 (N_3099,In_909,In_259);
nor U3100 (N_3100,In_155,In_947);
or U3101 (N_3101,In_601,In_626);
or U3102 (N_3102,In_547,In_725);
xnor U3103 (N_3103,In_129,In_547);
or U3104 (N_3104,In_642,In_772);
and U3105 (N_3105,In_402,In_558);
nand U3106 (N_3106,In_522,In_599);
nand U3107 (N_3107,In_366,In_935);
or U3108 (N_3108,In_477,In_607);
and U3109 (N_3109,In_227,In_188);
and U3110 (N_3110,In_971,In_85);
and U3111 (N_3111,In_115,In_579);
nand U3112 (N_3112,In_709,In_956);
xnor U3113 (N_3113,In_521,In_20);
xnor U3114 (N_3114,In_916,In_539);
xnor U3115 (N_3115,In_700,In_60);
nor U3116 (N_3116,In_210,In_367);
nand U3117 (N_3117,In_941,In_212);
or U3118 (N_3118,In_810,In_809);
or U3119 (N_3119,In_993,In_84);
nand U3120 (N_3120,In_272,In_23);
nor U3121 (N_3121,In_836,In_901);
nand U3122 (N_3122,In_622,In_41);
nor U3123 (N_3123,In_948,In_879);
and U3124 (N_3124,In_893,In_939);
or U3125 (N_3125,In_707,In_704);
or U3126 (N_3126,In_576,In_145);
and U3127 (N_3127,In_592,In_627);
xnor U3128 (N_3128,In_773,In_304);
nor U3129 (N_3129,In_12,In_42);
and U3130 (N_3130,In_677,In_820);
or U3131 (N_3131,In_628,In_543);
nor U3132 (N_3132,In_225,In_567);
xor U3133 (N_3133,In_159,In_682);
xnor U3134 (N_3134,In_188,In_371);
xor U3135 (N_3135,In_402,In_622);
xnor U3136 (N_3136,In_156,In_860);
or U3137 (N_3137,In_987,In_758);
and U3138 (N_3138,In_765,In_700);
nand U3139 (N_3139,In_912,In_345);
nand U3140 (N_3140,In_473,In_252);
nand U3141 (N_3141,In_874,In_20);
nand U3142 (N_3142,In_822,In_649);
or U3143 (N_3143,In_846,In_556);
xor U3144 (N_3144,In_6,In_346);
nor U3145 (N_3145,In_741,In_488);
xnor U3146 (N_3146,In_894,In_869);
nand U3147 (N_3147,In_339,In_588);
nor U3148 (N_3148,In_488,In_56);
or U3149 (N_3149,In_914,In_24);
xor U3150 (N_3150,In_769,In_100);
nand U3151 (N_3151,In_789,In_25);
nand U3152 (N_3152,In_661,In_699);
or U3153 (N_3153,In_156,In_689);
nand U3154 (N_3154,In_304,In_550);
nand U3155 (N_3155,In_659,In_110);
nor U3156 (N_3156,In_476,In_576);
and U3157 (N_3157,In_378,In_725);
xnor U3158 (N_3158,In_9,In_954);
or U3159 (N_3159,In_149,In_731);
nor U3160 (N_3160,In_944,In_58);
xor U3161 (N_3161,In_832,In_175);
nor U3162 (N_3162,In_308,In_200);
nand U3163 (N_3163,In_903,In_564);
nor U3164 (N_3164,In_4,In_168);
or U3165 (N_3165,In_184,In_980);
xor U3166 (N_3166,In_503,In_40);
nand U3167 (N_3167,In_234,In_445);
nor U3168 (N_3168,In_301,In_376);
nand U3169 (N_3169,In_344,In_159);
or U3170 (N_3170,In_680,In_851);
nand U3171 (N_3171,In_588,In_996);
nand U3172 (N_3172,In_484,In_726);
nor U3173 (N_3173,In_338,In_254);
and U3174 (N_3174,In_299,In_957);
nor U3175 (N_3175,In_517,In_819);
and U3176 (N_3176,In_426,In_401);
and U3177 (N_3177,In_570,In_657);
or U3178 (N_3178,In_171,In_72);
xnor U3179 (N_3179,In_690,In_618);
nand U3180 (N_3180,In_458,In_195);
or U3181 (N_3181,In_822,In_436);
and U3182 (N_3182,In_117,In_841);
xnor U3183 (N_3183,In_98,In_532);
nand U3184 (N_3184,In_555,In_262);
and U3185 (N_3185,In_860,In_879);
nand U3186 (N_3186,In_215,In_938);
nor U3187 (N_3187,In_122,In_709);
nand U3188 (N_3188,In_899,In_332);
and U3189 (N_3189,In_652,In_893);
and U3190 (N_3190,In_443,In_333);
xor U3191 (N_3191,In_566,In_217);
or U3192 (N_3192,In_117,In_411);
or U3193 (N_3193,In_921,In_837);
nand U3194 (N_3194,In_717,In_79);
and U3195 (N_3195,In_171,In_739);
xor U3196 (N_3196,In_666,In_692);
nand U3197 (N_3197,In_964,In_518);
or U3198 (N_3198,In_825,In_766);
nor U3199 (N_3199,In_894,In_503);
nor U3200 (N_3200,In_693,In_766);
and U3201 (N_3201,In_481,In_728);
or U3202 (N_3202,In_453,In_935);
or U3203 (N_3203,In_398,In_799);
and U3204 (N_3204,In_80,In_571);
nor U3205 (N_3205,In_795,In_529);
nor U3206 (N_3206,In_217,In_705);
nand U3207 (N_3207,In_373,In_441);
nand U3208 (N_3208,In_164,In_161);
and U3209 (N_3209,In_493,In_323);
nand U3210 (N_3210,In_457,In_102);
or U3211 (N_3211,In_688,In_855);
or U3212 (N_3212,In_336,In_388);
and U3213 (N_3213,In_401,In_989);
and U3214 (N_3214,In_714,In_959);
nand U3215 (N_3215,In_255,In_958);
nand U3216 (N_3216,In_258,In_507);
nand U3217 (N_3217,In_579,In_948);
nand U3218 (N_3218,In_223,In_932);
or U3219 (N_3219,In_973,In_400);
xor U3220 (N_3220,In_652,In_794);
and U3221 (N_3221,In_952,In_255);
or U3222 (N_3222,In_422,In_479);
xor U3223 (N_3223,In_760,In_338);
nor U3224 (N_3224,In_569,In_333);
nand U3225 (N_3225,In_457,In_2);
or U3226 (N_3226,In_905,In_944);
nand U3227 (N_3227,In_864,In_856);
nand U3228 (N_3228,In_709,In_987);
and U3229 (N_3229,In_162,In_111);
and U3230 (N_3230,In_298,In_535);
nand U3231 (N_3231,In_316,In_659);
and U3232 (N_3232,In_276,In_922);
nand U3233 (N_3233,In_379,In_474);
nand U3234 (N_3234,In_784,In_28);
and U3235 (N_3235,In_121,In_581);
nand U3236 (N_3236,In_861,In_502);
or U3237 (N_3237,In_571,In_215);
or U3238 (N_3238,In_924,In_464);
xor U3239 (N_3239,In_607,In_711);
or U3240 (N_3240,In_193,In_74);
and U3241 (N_3241,In_539,In_335);
or U3242 (N_3242,In_829,In_884);
and U3243 (N_3243,In_733,In_498);
xnor U3244 (N_3244,In_557,In_949);
and U3245 (N_3245,In_161,In_414);
nor U3246 (N_3246,In_429,In_546);
xnor U3247 (N_3247,In_293,In_676);
nand U3248 (N_3248,In_928,In_747);
nor U3249 (N_3249,In_263,In_141);
nand U3250 (N_3250,In_258,In_667);
nand U3251 (N_3251,In_337,In_258);
nand U3252 (N_3252,In_10,In_114);
xor U3253 (N_3253,In_220,In_183);
and U3254 (N_3254,In_720,In_106);
or U3255 (N_3255,In_927,In_344);
or U3256 (N_3256,In_758,In_349);
nor U3257 (N_3257,In_135,In_863);
and U3258 (N_3258,In_935,In_792);
and U3259 (N_3259,In_751,In_394);
nor U3260 (N_3260,In_60,In_77);
or U3261 (N_3261,In_835,In_289);
and U3262 (N_3262,In_808,In_181);
nand U3263 (N_3263,In_256,In_360);
or U3264 (N_3264,In_584,In_921);
nand U3265 (N_3265,In_918,In_781);
and U3266 (N_3266,In_973,In_370);
nor U3267 (N_3267,In_798,In_862);
nor U3268 (N_3268,In_368,In_913);
xor U3269 (N_3269,In_988,In_293);
or U3270 (N_3270,In_407,In_583);
xor U3271 (N_3271,In_940,In_106);
and U3272 (N_3272,In_603,In_135);
and U3273 (N_3273,In_632,In_792);
nand U3274 (N_3274,In_680,In_572);
nor U3275 (N_3275,In_713,In_612);
nand U3276 (N_3276,In_415,In_371);
nand U3277 (N_3277,In_36,In_168);
or U3278 (N_3278,In_337,In_903);
nand U3279 (N_3279,In_303,In_413);
and U3280 (N_3280,In_847,In_226);
nand U3281 (N_3281,In_966,In_524);
nand U3282 (N_3282,In_205,In_292);
nor U3283 (N_3283,In_763,In_553);
xnor U3284 (N_3284,In_119,In_424);
nand U3285 (N_3285,In_196,In_406);
and U3286 (N_3286,In_346,In_638);
nor U3287 (N_3287,In_580,In_825);
nand U3288 (N_3288,In_632,In_909);
nor U3289 (N_3289,In_661,In_84);
or U3290 (N_3290,In_948,In_798);
and U3291 (N_3291,In_541,In_604);
nand U3292 (N_3292,In_579,In_582);
or U3293 (N_3293,In_925,In_750);
nor U3294 (N_3294,In_502,In_665);
nand U3295 (N_3295,In_330,In_267);
nand U3296 (N_3296,In_903,In_217);
nor U3297 (N_3297,In_163,In_573);
or U3298 (N_3298,In_760,In_68);
nand U3299 (N_3299,In_725,In_922);
nor U3300 (N_3300,In_377,In_791);
nor U3301 (N_3301,In_606,In_665);
nand U3302 (N_3302,In_601,In_194);
nand U3303 (N_3303,In_508,In_826);
nand U3304 (N_3304,In_663,In_705);
nand U3305 (N_3305,In_121,In_103);
and U3306 (N_3306,In_126,In_835);
nand U3307 (N_3307,In_422,In_230);
nand U3308 (N_3308,In_703,In_317);
and U3309 (N_3309,In_989,In_929);
nor U3310 (N_3310,In_307,In_993);
nor U3311 (N_3311,In_437,In_635);
nand U3312 (N_3312,In_335,In_117);
and U3313 (N_3313,In_807,In_310);
or U3314 (N_3314,In_23,In_507);
or U3315 (N_3315,In_546,In_198);
or U3316 (N_3316,In_708,In_352);
xnor U3317 (N_3317,In_671,In_400);
nand U3318 (N_3318,In_393,In_805);
nor U3319 (N_3319,In_653,In_342);
or U3320 (N_3320,In_239,In_867);
nand U3321 (N_3321,In_846,In_577);
nand U3322 (N_3322,In_771,In_464);
or U3323 (N_3323,In_560,In_608);
nand U3324 (N_3324,In_862,In_363);
and U3325 (N_3325,In_658,In_602);
or U3326 (N_3326,In_202,In_948);
nand U3327 (N_3327,In_608,In_322);
nor U3328 (N_3328,In_599,In_660);
nand U3329 (N_3329,In_347,In_862);
nor U3330 (N_3330,In_399,In_150);
and U3331 (N_3331,In_130,In_4);
nor U3332 (N_3332,In_345,In_644);
xor U3333 (N_3333,In_516,In_513);
or U3334 (N_3334,In_765,In_164);
nor U3335 (N_3335,In_566,In_673);
nor U3336 (N_3336,In_88,In_24);
nor U3337 (N_3337,In_962,In_335);
nand U3338 (N_3338,In_747,In_320);
or U3339 (N_3339,In_699,In_794);
or U3340 (N_3340,In_990,In_642);
or U3341 (N_3341,In_380,In_591);
and U3342 (N_3342,In_671,In_357);
or U3343 (N_3343,In_530,In_54);
nor U3344 (N_3344,In_941,In_340);
nor U3345 (N_3345,In_139,In_735);
and U3346 (N_3346,In_90,In_675);
xor U3347 (N_3347,In_163,In_421);
or U3348 (N_3348,In_615,In_536);
or U3349 (N_3349,In_372,In_274);
nand U3350 (N_3350,In_66,In_692);
or U3351 (N_3351,In_569,In_260);
nand U3352 (N_3352,In_949,In_972);
and U3353 (N_3353,In_900,In_732);
or U3354 (N_3354,In_133,In_696);
xnor U3355 (N_3355,In_736,In_681);
or U3356 (N_3356,In_535,In_796);
or U3357 (N_3357,In_554,In_447);
nor U3358 (N_3358,In_881,In_230);
or U3359 (N_3359,In_8,In_86);
or U3360 (N_3360,In_977,In_258);
and U3361 (N_3361,In_184,In_979);
nor U3362 (N_3362,In_192,In_652);
nor U3363 (N_3363,In_745,In_875);
or U3364 (N_3364,In_354,In_209);
and U3365 (N_3365,In_35,In_826);
or U3366 (N_3366,In_688,In_433);
nand U3367 (N_3367,In_864,In_377);
or U3368 (N_3368,In_183,In_479);
nand U3369 (N_3369,In_735,In_207);
xor U3370 (N_3370,In_382,In_367);
xnor U3371 (N_3371,In_801,In_511);
nor U3372 (N_3372,In_602,In_0);
nand U3373 (N_3373,In_977,In_548);
nand U3374 (N_3374,In_804,In_640);
nor U3375 (N_3375,In_239,In_863);
or U3376 (N_3376,In_404,In_949);
and U3377 (N_3377,In_996,In_713);
nor U3378 (N_3378,In_466,In_516);
and U3379 (N_3379,In_341,In_760);
or U3380 (N_3380,In_757,In_464);
and U3381 (N_3381,In_421,In_139);
and U3382 (N_3382,In_840,In_192);
nor U3383 (N_3383,In_47,In_425);
and U3384 (N_3384,In_992,In_679);
xnor U3385 (N_3385,In_681,In_268);
or U3386 (N_3386,In_498,In_590);
and U3387 (N_3387,In_381,In_227);
nor U3388 (N_3388,In_663,In_854);
or U3389 (N_3389,In_864,In_334);
nor U3390 (N_3390,In_895,In_675);
nand U3391 (N_3391,In_246,In_763);
nor U3392 (N_3392,In_209,In_373);
nor U3393 (N_3393,In_402,In_942);
or U3394 (N_3394,In_838,In_477);
and U3395 (N_3395,In_105,In_954);
and U3396 (N_3396,In_829,In_473);
nand U3397 (N_3397,In_39,In_528);
nand U3398 (N_3398,In_198,In_409);
nor U3399 (N_3399,In_905,In_943);
nand U3400 (N_3400,In_251,In_249);
nand U3401 (N_3401,In_10,In_698);
nand U3402 (N_3402,In_571,In_962);
nand U3403 (N_3403,In_25,In_949);
or U3404 (N_3404,In_82,In_794);
nor U3405 (N_3405,In_948,In_235);
and U3406 (N_3406,In_116,In_93);
and U3407 (N_3407,In_662,In_545);
nand U3408 (N_3408,In_540,In_427);
or U3409 (N_3409,In_25,In_815);
nand U3410 (N_3410,In_796,In_124);
or U3411 (N_3411,In_948,In_803);
nor U3412 (N_3412,In_64,In_607);
and U3413 (N_3413,In_624,In_11);
and U3414 (N_3414,In_897,In_16);
xor U3415 (N_3415,In_895,In_367);
nor U3416 (N_3416,In_104,In_452);
xnor U3417 (N_3417,In_570,In_137);
nor U3418 (N_3418,In_106,In_19);
nand U3419 (N_3419,In_29,In_46);
nand U3420 (N_3420,In_974,In_964);
nand U3421 (N_3421,In_532,In_43);
or U3422 (N_3422,In_893,In_922);
nor U3423 (N_3423,In_653,In_441);
xor U3424 (N_3424,In_315,In_368);
nor U3425 (N_3425,In_307,In_505);
nor U3426 (N_3426,In_829,In_430);
nand U3427 (N_3427,In_331,In_51);
and U3428 (N_3428,In_978,In_924);
xor U3429 (N_3429,In_489,In_297);
or U3430 (N_3430,In_588,In_696);
and U3431 (N_3431,In_802,In_342);
or U3432 (N_3432,In_22,In_993);
xnor U3433 (N_3433,In_817,In_857);
nor U3434 (N_3434,In_745,In_472);
nor U3435 (N_3435,In_607,In_840);
and U3436 (N_3436,In_799,In_63);
xnor U3437 (N_3437,In_958,In_338);
or U3438 (N_3438,In_852,In_622);
nand U3439 (N_3439,In_956,In_66);
nand U3440 (N_3440,In_762,In_746);
and U3441 (N_3441,In_184,In_175);
nor U3442 (N_3442,In_784,In_821);
or U3443 (N_3443,In_319,In_570);
or U3444 (N_3444,In_858,In_264);
nand U3445 (N_3445,In_399,In_593);
or U3446 (N_3446,In_749,In_834);
nor U3447 (N_3447,In_270,In_308);
nor U3448 (N_3448,In_151,In_773);
or U3449 (N_3449,In_882,In_723);
nor U3450 (N_3450,In_123,In_734);
nand U3451 (N_3451,In_55,In_75);
and U3452 (N_3452,In_530,In_64);
or U3453 (N_3453,In_798,In_681);
nor U3454 (N_3454,In_91,In_927);
xnor U3455 (N_3455,In_710,In_310);
nor U3456 (N_3456,In_601,In_331);
nand U3457 (N_3457,In_820,In_857);
and U3458 (N_3458,In_531,In_956);
nor U3459 (N_3459,In_733,In_523);
nor U3460 (N_3460,In_60,In_414);
or U3461 (N_3461,In_679,In_65);
or U3462 (N_3462,In_36,In_283);
nor U3463 (N_3463,In_862,In_394);
nand U3464 (N_3464,In_31,In_784);
nand U3465 (N_3465,In_920,In_845);
or U3466 (N_3466,In_534,In_87);
and U3467 (N_3467,In_248,In_606);
or U3468 (N_3468,In_986,In_548);
and U3469 (N_3469,In_613,In_642);
or U3470 (N_3470,In_83,In_473);
and U3471 (N_3471,In_695,In_494);
and U3472 (N_3472,In_196,In_215);
nand U3473 (N_3473,In_32,In_519);
or U3474 (N_3474,In_747,In_596);
nor U3475 (N_3475,In_179,In_96);
nand U3476 (N_3476,In_347,In_398);
and U3477 (N_3477,In_686,In_263);
and U3478 (N_3478,In_828,In_763);
and U3479 (N_3479,In_482,In_774);
nor U3480 (N_3480,In_471,In_746);
nand U3481 (N_3481,In_964,In_590);
and U3482 (N_3482,In_127,In_62);
nand U3483 (N_3483,In_658,In_604);
and U3484 (N_3484,In_885,In_73);
and U3485 (N_3485,In_825,In_382);
nor U3486 (N_3486,In_842,In_92);
nand U3487 (N_3487,In_812,In_795);
nand U3488 (N_3488,In_514,In_31);
nor U3489 (N_3489,In_368,In_448);
nor U3490 (N_3490,In_500,In_622);
nand U3491 (N_3491,In_715,In_649);
or U3492 (N_3492,In_502,In_370);
or U3493 (N_3493,In_609,In_106);
and U3494 (N_3494,In_890,In_310);
nor U3495 (N_3495,In_753,In_62);
and U3496 (N_3496,In_358,In_114);
xnor U3497 (N_3497,In_18,In_476);
and U3498 (N_3498,In_650,In_870);
nor U3499 (N_3499,In_815,In_486);
nor U3500 (N_3500,In_721,In_157);
and U3501 (N_3501,In_864,In_646);
nand U3502 (N_3502,In_483,In_540);
nand U3503 (N_3503,In_345,In_756);
or U3504 (N_3504,In_788,In_615);
nand U3505 (N_3505,In_829,In_25);
or U3506 (N_3506,In_893,In_69);
or U3507 (N_3507,In_655,In_744);
xor U3508 (N_3508,In_208,In_788);
and U3509 (N_3509,In_152,In_317);
and U3510 (N_3510,In_198,In_225);
nand U3511 (N_3511,In_0,In_980);
nand U3512 (N_3512,In_228,In_780);
and U3513 (N_3513,In_401,In_920);
nor U3514 (N_3514,In_970,In_348);
nand U3515 (N_3515,In_548,In_186);
and U3516 (N_3516,In_674,In_574);
nand U3517 (N_3517,In_37,In_449);
or U3518 (N_3518,In_221,In_482);
nand U3519 (N_3519,In_401,In_296);
or U3520 (N_3520,In_526,In_473);
nor U3521 (N_3521,In_824,In_404);
or U3522 (N_3522,In_792,In_927);
nand U3523 (N_3523,In_400,In_426);
or U3524 (N_3524,In_981,In_329);
and U3525 (N_3525,In_26,In_862);
or U3526 (N_3526,In_117,In_898);
nor U3527 (N_3527,In_214,In_656);
or U3528 (N_3528,In_732,In_471);
and U3529 (N_3529,In_482,In_51);
nor U3530 (N_3530,In_861,In_874);
nand U3531 (N_3531,In_881,In_838);
xnor U3532 (N_3532,In_950,In_116);
or U3533 (N_3533,In_602,In_524);
nand U3534 (N_3534,In_135,In_890);
nand U3535 (N_3535,In_214,In_938);
or U3536 (N_3536,In_51,In_125);
and U3537 (N_3537,In_214,In_426);
nor U3538 (N_3538,In_802,In_919);
nand U3539 (N_3539,In_683,In_848);
nor U3540 (N_3540,In_263,In_539);
and U3541 (N_3541,In_559,In_70);
nand U3542 (N_3542,In_835,In_645);
xnor U3543 (N_3543,In_254,In_28);
or U3544 (N_3544,In_202,In_459);
and U3545 (N_3545,In_386,In_675);
nand U3546 (N_3546,In_502,In_597);
xnor U3547 (N_3547,In_523,In_410);
or U3548 (N_3548,In_390,In_177);
or U3549 (N_3549,In_528,In_230);
nor U3550 (N_3550,In_673,In_427);
or U3551 (N_3551,In_900,In_205);
and U3552 (N_3552,In_609,In_674);
and U3553 (N_3553,In_643,In_522);
xnor U3554 (N_3554,In_36,In_992);
nor U3555 (N_3555,In_968,In_182);
nand U3556 (N_3556,In_952,In_345);
nor U3557 (N_3557,In_686,In_920);
xor U3558 (N_3558,In_122,In_527);
nand U3559 (N_3559,In_824,In_918);
or U3560 (N_3560,In_987,In_827);
or U3561 (N_3561,In_579,In_360);
and U3562 (N_3562,In_723,In_676);
nand U3563 (N_3563,In_732,In_725);
nand U3564 (N_3564,In_877,In_762);
nand U3565 (N_3565,In_304,In_77);
xnor U3566 (N_3566,In_878,In_496);
nand U3567 (N_3567,In_299,In_359);
and U3568 (N_3568,In_14,In_552);
or U3569 (N_3569,In_388,In_260);
nor U3570 (N_3570,In_332,In_630);
and U3571 (N_3571,In_619,In_177);
or U3572 (N_3572,In_870,In_942);
and U3573 (N_3573,In_446,In_307);
and U3574 (N_3574,In_797,In_312);
or U3575 (N_3575,In_131,In_865);
nor U3576 (N_3576,In_467,In_627);
and U3577 (N_3577,In_487,In_558);
or U3578 (N_3578,In_263,In_709);
or U3579 (N_3579,In_129,In_75);
or U3580 (N_3580,In_639,In_271);
nor U3581 (N_3581,In_596,In_157);
nand U3582 (N_3582,In_878,In_375);
nand U3583 (N_3583,In_799,In_631);
and U3584 (N_3584,In_986,In_967);
or U3585 (N_3585,In_287,In_284);
xnor U3586 (N_3586,In_497,In_139);
and U3587 (N_3587,In_861,In_191);
xor U3588 (N_3588,In_988,In_724);
or U3589 (N_3589,In_450,In_235);
xnor U3590 (N_3590,In_713,In_291);
nand U3591 (N_3591,In_893,In_778);
and U3592 (N_3592,In_196,In_24);
xnor U3593 (N_3593,In_681,In_414);
or U3594 (N_3594,In_219,In_916);
and U3595 (N_3595,In_515,In_387);
and U3596 (N_3596,In_793,In_513);
and U3597 (N_3597,In_128,In_816);
or U3598 (N_3598,In_65,In_324);
or U3599 (N_3599,In_211,In_371);
nor U3600 (N_3600,In_937,In_675);
nor U3601 (N_3601,In_403,In_317);
or U3602 (N_3602,In_728,In_114);
xor U3603 (N_3603,In_923,In_908);
or U3604 (N_3604,In_886,In_845);
or U3605 (N_3605,In_462,In_167);
nor U3606 (N_3606,In_500,In_195);
nand U3607 (N_3607,In_107,In_136);
nand U3608 (N_3608,In_811,In_897);
or U3609 (N_3609,In_719,In_622);
or U3610 (N_3610,In_564,In_752);
nand U3611 (N_3611,In_314,In_662);
or U3612 (N_3612,In_270,In_114);
xor U3613 (N_3613,In_408,In_868);
and U3614 (N_3614,In_909,In_624);
or U3615 (N_3615,In_603,In_285);
nor U3616 (N_3616,In_826,In_387);
or U3617 (N_3617,In_803,In_245);
and U3618 (N_3618,In_335,In_996);
and U3619 (N_3619,In_126,In_576);
nand U3620 (N_3620,In_706,In_897);
nor U3621 (N_3621,In_575,In_532);
or U3622 (N_3622,In_750,In_641);
and U3623 (N_3623,In_321,In_774);
xnor U3624 (N_3624,In_933,In_509);
or U3625 (N_3625,In_906,In_885);
or U3626 (N_3626,In_622,In_897);
and U3627 (N_3627,In_112,In_838);
nor U3628 (N_3628,In_713,In_916);
nand U3629 (N_3629,In_407,In_140);
nor U3630 (N_3630,In_39,In_813);
or U3631 (N_3631,In_760,In_277);
nor U3632 (N_3632,In_450,In_226);
nand U3633 (N_3633,In_425,In_972);
and U3634 (N_3634,In_711,In_660);
or U3635 (N_3635,In_865,In_788);
or U3636 (N_3636,In_430,In_147);
nand U3637 (N_3637,In_743,In_569);
nand U3638 (N_3638,In_70,In_102);
and U3639 (N_3639,In_64,In_410);
nand U3640 (N_3640,In_514,In_155);
nor U3641 (N_3641,In_558,In_296);
or U3642 (N_3642,In_995,In_964);
or U3643 (N_3643,In_859,In_468);
or U3644 (N_3644,In_526,In_682);
and U3645 (N_3645,In_189,In_381);
nand U3646 (N_3646,In_47,In_700);
or U3647 (N_3647,In_17,In_76);
nand U3648 (N_3648,In_297,In_323);
and U3649 (N_3649,In_679,In_454);
nand U3650 (N_3650,In_941,In_959);
and U3651 (N_3651,In_826,In_753);
or U3652 (N_3652,In_985,In_853);
nor U3653 (N_3653,In_914,In_548);
nand U3654 (N_3654,In_642,In_265);
and U3655 (N_3655,In_996,In_248);
or U3656 (N_3656,In_530,In_341);
xnor U3657 (N_3657,In_720,In_188);
xor U3658 (N_3658,In_323,In_956);
and U3659 (N_3659,In_915,In_753);
or U3660 (N_3660,In_335,In_689);
and U3661 (N_3661,In_324,In_481);
nand U3662 (N_3662,In_615,In_95);
and U3663 (N_3663,In_493,In_869);
nand U3664 (N_3664,In_569,In_357);
or U3665 (N_3665,In_19,In_705);
or U3666 (N_3666,In_812,In_552);
xnor U3667 (N_3667,In_914,In_30);
xnor U3668 (N_3668,In_469,In_75);
or U3669 (N_3669,In_517,In_748);
or U3670 (N_3670,In_551,In_176);
nor U3671 (N_3671,In_980,In_381);
and U3672 (N_3672,In_350,In_140);
and U3673 (N_3673,In_569,In_359);
or U3674 (N_3674,In_197,In_328);
nand U3675 (N_3675,In_383,In_214);
nand U3676 (N_3676,In_958,In_36);
nand U3677 (N_3677,In_375,In_282);
xor U3678 (N_3678,In_934,In_593);
xnor U3679 (N_3679,In_280,In_766);
nor U3680 (N_3680,In_337,In_74);
and U3681 (N_3681,In_269,In_453);
and U3682 (N_3682,In_724,In_545);
nand U3683 (N_3683,In_776,In_20);
nand U3684 (N_3684,In_724,In_443);
nand U3685 (N_3685,In_468,In_922);
or U3686 (N_3686,In_255,In_991);
nor U3687 (N_3687,In_171,In_860);
xnor U3688 (N_3688,In_456,In_923);
nand U3689 (N_3689,In_223,In_583);
and U3690 (N_3690,In_907,In_716);
nor U3691 (N_3691,In_272,In_968);
xor U3692 (N_3692,In_495,In_812);
and U3693 (N_3693,In_841,In_955);
and U3694 (N_3694,In_371,In_161);
nand U3695 (N_3695,In_264,In_866);
nand U3696 (N_3696,In_98,In_807);
xnor U3697 (N_3697,In_301,In_787);
nand U3698 (N_3698,In_982,In_895);
xnor U3699 (N_3699,In_303,In_911);
and U3700 (N_3700,In_898,In_778);
nor U3701 (N_3701,In_483,In_742);
and U3702 (N_3702,In_413,In_819);
xor U3703 (N_3703,In_511,In_939);
nand U3704 (N_3704,In_794,In_889);
nand U3705 (N_3705,In_871,In_85);
nor U3706 (N_3706,In_353,In_129);
nor U3707 (N_3707,In_509,In_614);
nor U3708 (N_3708,In_350,In_739);
nand U3709 (N_3709,In_659,In_264);
or U3710 (N_3710,In_879,In_145);
nor U3711 (N_3711,In_89,In_581);
nor U3712 (N_3712,In_721,In_232);
and U3713 (N_3713,In_943,In_253);
and U3714 (N_3714,In_215,In_327);
nor U3715 (N_3715,In_151,In_911);
nand U3716 (N_3716,In_363,In_412);
nor U3717 (N_3717,In_919,In_815);
or U3718 (N_3718,In_868,In_96);
or U3719 (N_3719,In_998,In_780);
or U3720 (N_3720,In_500,In_17);
nor U3721 (N_3721,In_252,In_405);
nand U3722 (N_3722,In_998,In_63);
xnor U3723 (N_3723,In_594,In_571);
nand U3724 (N_3724,In_337,In_618);
and U3725 (N_3725,In_815,In_808);
nand U3726 (N_3726,In_815,In_234);
nor U3727 (N_3727,In_719,In_850);
or U3728 (N_3728,In_64,In_637);
nand U3729 (N_3729,In_798,In_178);
or U3730 (N_3730,In_858,In_961);
and U3731 (N_3731,In_144,In_27);
and U3732 (N_3732,In_450,In_991);
nor U3733 (N_3733,In_520,In_381);
nor U3734 (N_3734,In_302,In_552);
xnor U3735 (N_3735,In_527,In_5);
nand U3736 (N_3736,In_757,In_765);
or U3737 (N_3737,In_731,In_155);
xnor U3738 (N_3738,In_144,In_873);
xnor U3739 (N_3739,In_581,In_451);
and U3740 (N_3740,In_693,In_299);
and U3741 (N_3741,In_235,In_212);
xor U3742 (N_3742,In_286,In_683);
or U3743 (N_3743,In_18,In_743);
or U3744 (N_3744,In_783,In_740);
and U3745 (N_3745,In_8,In_716);
and U3746 (N_3746,In_424,In_524);
xnor U3747 (N_3747,In_457,In_759);
nor U3748 (N_3748,In_493,In_742);
and U3749 (N_3749,In_98,In_68);
or U3750 (N_3750,In_97,In_405);
nand U3751 (N_3751,In_314,In_427);
nand U3752 (N_3752,In_988,In_807);
and U3753 (N_3753,In_630,In_652);
nand U3754 (N_3754,In_397,In_235);
nor U3755 (N_3755,In_722,In_362);
or U3756 (N_3756,In_236,In_274);
nor U3757 (N_3757,In_2,In_191);
nor U3758 (N_3758,In_925,In_63);
or U3759 (N_3759,In_359,In_154);
nand U3760 (N_3760,In_760,In_883);
nand U3761 (N_3761,In_526,In_176);
nand U3762 (N_3762,In_696,In_803);
or U3763 (N_3763,In_32,In_755);
nor U3764 (N_3764,In_130,In_816);
or U3765 (N_3765,In_166,In_645);
or U3766 (N_3766,In_837,In_487);
or U3767 (N_3767,In_615,In_933);
nand U3768 (N_3768,In_710,In_41);
nand U3769 (N_3769,In_142,In_550);
and U3770 (N_3770,In_271,In_224);
nand U3771 (N_3771,In_819,In_671);
and U3772 (N_3772,In_353,In_950);
nand U3773 (N_3773,In_634,In_32);
nand U3774 (N_3774,In_900,In_75);
nor U3775 (N_3775,In_805,In_921);
nor U3776 (N_3776,In_698,In_383);
nor U3777 (N_3777,In_444,In_516);
xnor U3778 (N_3778,In_880,In_758);
and U3779 (N_3779,In_785,In_438);
nor U3780 (N_3780,In_868,In_585);
and U3781 (N_3781,In_807,In_568);
or U3782 (N_3782,In_167,In_510);
or U3783 (N_3783,In_221,In_723);
nor U3784 (N_3784,In_725,In_271);
nand U3785 (N_3785,In_709,In_689);
nor U3786 (N_3786,In_280,In_61);
xnor U3787 (N_3787,In_446,In_333);
or U3788 (N_3788,In_735,In_952);
nor U3789 (N_3789,In_189,In_348);
nand U3790 (N_3790,In_340,In_93);
nor U3791 (N_3791,In_553,In_407);
or U3792 (N_3792,In_446,In_748);
or U3793 (N_3793,In_291,In_130);
nor U3794 (N_3794,In_691,In_766);
or U3795 (N_3795,In_213,In_676);
nor U3796 (N_3796,In_827,In_608);
nor U3797 (N_3797,In_105,In_422);
nand U3798 (N_3798,In_232,In_673);
and U3799 (N_3799,In_194,In_941);
nand U3800 (N_3800,In_475,In_523);
nor U3801 (N_3801,In_816,In_712);
and U3802 (N_3802,In_255,In_823);
nand U3803 (N_3803,In_84,In_654);
nor U3804 (N_3804,In_169,In_127);
and U3805 (N_3805,In_788,In_87);
or U3806 (N_3806,In_97,In_95);
nor U3807 (N_3807,In_46,In_70);
and U3808 (N_3808,In_611,In_576);
and U3809 (N_3809,In_626,In_304);
nor U3810 (N_3810,In_647,In_136);
and U3811 (N_3811,In_534,In_452);
nor U3812 (N_3812,In_364,In_858);
and U3813 (N_3813,In_242,In_572);
nor U3814 (N_3814,In_730,In_996);
nand U3815 (N_3815,In_339,In_62);
nand U3816 (N_3816,In_160,In_621);
and U3817 (N_3817,In_91,In_59);
nor U3818 (N_3818,In_933,In_73);
nor U3819 (N_3819,In_768,In_367);
nand U3820 (N_3820,In_766,In_748);
nor U3821 (N_3821,In_722,In_624);
and U3822 (N_3822,In_557,In_809);
nand U3823 (N_3823,In_61,In_980);
and U3824 (N_3824,In_669,In_713);
or U3825 (N_3825,In_133,In_381);
and U3826 (N_3826,In_144,In_584);
nand U3827 (N_3827,In_292,In_234);
nor U3828 (N_3828,In_124,In_797);
nor U3829 (N_3829,In_338,In_164);
nor U3830 (N_3830,In_580,In_323);
nand U3831 (N_3831,In_743,In_577);
nand U3832 (N_3832,In_935,In_267);
and U3833 (N_3833,In_269,In_541);
nand U3834 (N_3834,In_675,In_541);
and U3835 (N_3835,In_435,In_332);
nor U3836 (N_3836,In_177,In_528);
or U3837 (N_3837,In_880,In_241);
and U3838 (N_3838,In_58,In_216);
nand U3839 (N_3839,In_924,In_840);
nand U3840 (N_3840,In_178,In_813);
nor U3841 (N_3841,In_98,In_332);
xor U3842 (N_3842,In_606,In_993);
nor U3843 (N_3843,In_461,In_470);
and U3844 (N_3844,In_216,In_610);
nor U3845 (N_3845,In_207,In_688);
xor U3846 (N_3846,In_370,In_260);
nor U3847 (N_3847,In_175,In_120);
and U3848 (N_3848,In_994,In_85);
nand U3849 (N_3849,In_279,In_166);
nor U3850 (N_3850,In_91,In_168);
or U3851 (N_3851,In_349,In_656);
or U3852 (N_3852,In_819,In_769);
or U3853 (N_3853,In_875,In_738);
nand U3854 (N_3854,In_733,In_560);
and U3855 (N_3855,In_631,In_415);
and U3856 (N_3856,In_147,In_558);
or U3857 (N_3857,In_911,In_832);
xor U3858 (N_3858,In_699,In_262);
and U3859 (N_3859,In_689,In_671);
nand U3860 (N_3860,In_953,In_546);
and U3861 (N_3861,In_89,In_418);
and U3862 (N_3862,In_433,In_321);
nor U3863 (N_3863,In_123,In_890);
or U3864 (N_3864,In_56,In_579);
and U3865 (N_3865,In_654,In_684);
and U3866 (N_3866,In_360,In_214);
and U3867 (N_3867,In_859,In_23);
xnor U3868 (N_3868,In_86,In_283);
nand U3869 (N_3869,In_991,In_814);
nor U3870 (N_3870,In_13,In_766);
nand U3871 (N_3871,In_71,In_913);
nand U3872 (N_3872,In_175,In_637);
or U3873 (N_3873,In_130,In_310);
xor U3874 (N_3874,In_954,In_895);
and U3875 (N_3875,In_790,In_511);
and U3876 (N_3876,In_716,In_237);
nor U3877 (N_3877,In_336,In_510);
and U3878 (N_3878,In_340,In_988);
nand U3879 (N_3879,In_691,In_426);
or U3880 (N_3880,In_870,In_586);
or U3881 (N_3881,In_77,In_212);
or U3882 (N_3882,In_966,In_987);
or U3883 (N_3883,In_914,In_769);
and U3884 (N_3884,In_447,In_587);
nor U3885 (N_3885,In_377,In_443);
and U3886 (N_3886,In_63,In_28);
or U3887 (N_3887,In_243,In_663);
nor U3888 (N_3888,In_945,In_792);
nand U3889 (N_3889,In_201,In_913);
nand U3890 (N_3890,In_693,In_647);
nand U3891 (N_3891,In_417,In_185);
nor U3892 (N_3892,In_249,In_59);
nand U3893 (N_3893,In_824,In_977);
and U3894 (N_3894,In_344,In_488);
and U3895 (N_3895,In_856,In_158);
nand U3896 (N_3896,In_178,In_877);
nand U3897 (N_3897,In_172,In_220);
and U3898 (N_3898,In_46,In_513);
nand U3899 (N_3899,In_603,In_872);
nand U3900 (N_3900,In_942,In_422);
and U3901 (N_3901,In_844,In_646);
nor U3902 (N_3902,In_897,In_544);
nand U3903 (N_3903,In_224,In_809);
or U3904 (N_3904,In_511,In_85);
nor U3905 (N_3905,In_189,In_632);
and U3906 (N_3906,In_651,In_405);
xnor U3907 (N_3907,In_324,In_69);
nor U3908 (N_3908,In_480,In_211);
nor U3909 (N_3909,In_739,In_951);
xnor U3910 (N_3910,In_755,In_111);
xnor U3911 (N_3911,In_79,In_83);
nor U3912 (N_3912,In_81,In_407);
nand U3913 (N_3913,In_228,In_229);
nand U3914 (N_3914,In_540,In_280);
nor U3915 (N_3915,In_748,In_668);
nand U3916 (N_3916,In_424,In_980);
or U3917 (N_3917,In_616,In_51);
nor U3918 (N_3918,In_713,In_427);
nor U3919 (N_3919,In_244,In_156);
or U3920 (N_3920,In_969,In_658);
nor U3921 (N_3921,In_152,In_136);
and U3922 (N_3922,In_26,In_432);
and U3923 (N_3923,In_373,In_171);
or U3924 (N_3924,In_734,In_418);
nand U3925 (N_3925,In_702,In_517);
xor U3926 (N_3926,In_977,In_428);
nor U3927 (N_3927,In_293,In_853);
nor U3928 (N_3928,In_511,In_927);
nand U3929 (N_3929,In_250,In_354);
xnor U3930 (N_3930,In_669,In_695);
and U3931 (N_3931,In_869,In_727);
nor U3932 (N_3932,In_622,In_594);
nand U3933 (N_3933,In_263,In_175);
nand U3934 (N_3934,In_699,In_11);
nand U3935 (N_3935,In_370,In_686);
and U3936 (N_3936,In_935,In_717);
nor U3937 (N_3937,In_433,In_616);
nor U3938 (N_3938,In_591,In_624);
nand U3939 (N_3939,In_268,In_447);
and U3940 (N_3940,In_577,In_710);
and U3941 (N_3941,In_940,In_385);
nor U3942 (N_3942,In_185,In_786);
nor U3943 (N_3943,In_633,In_975);
nand U3944 (N_3944,In_317,In_879);
xnor U3945 (N_3945,In_397,In_7);
or U3946 (N_3946,In_758,In_255);
and U3947 (N_3947,In_865,In_336);
xnor U3948 (N_3948,In_27,In_74);
nand U3949 (N_3949,In_48,In_215);
nor U3950 (N_3950,In_243,In_766);
and U3951 (N_3951,In_808,In_669);
and U3952 (N_3952,In_515,In_192);
nor U3953 (N_3953,In_240,In_796);
and U3954 (N_3954,In_57,In_261);
nor U3955 (N_3955,In_116,In_446);
nand U3956 (N_3956,In_417,In_178);
or U3957 (N_3957,In_237,In_212);
nor U3958 (N_3958,In_885,In_62);
or U3959 (N_3959,In_389,In_254);
and U3960 (N_3960,In_761,In_12);
nand U3961 (N_3961,In_43,In_394);
or U3962 (N_3962,In_748,In_740);
and U3963 (N_3963,In_650,In_763);
and U3964 (N_3964,In_331,In_180);
xor U3965 (N_3965,In_617,In_630);
nand U3966 (N_3966,In_396,In_544);
and U3967 (N_3967,In_620,In_121);
nor U3968 (N_3968,In_135,In_888);
nor U3969 (N_3969,In_238,In_235);
or U3970 (N_3970,In_419,In_93);
or U3971 (N_3971,In_705,In_14);
nor U3972 (N_3972,In_777,In_216);
nor U3973 (N_3973,In_340,In_325);
or U3974 (N_3974,In_627,In_204);
and U3975 (N_3975,In_776,In_988);
nand U3976 (N_3976,In_892,In_107);
xor U3977 (N_3977,In_755,In_227);
nor U3978 (N_3978,In_892,In_190);
and U3979 (N_3979,In_918,In_397);
nor U3980 (N_3980,In_691,In_747);
and U3981 (N_3981,In_372,In_658);
nand U3982 (N_3982,In_318,In_31);
and U3983 (N_3983,In_616,In_814);
or U3984 (N_3984,In_662,In_580);
and U3985 (N_3985,In_806,In_163);
nor U3986 (N_3986,In_31,In_531);
nand U3987 (N_3987,In_517,In_989);
and U3988 (N_3988,In_330,In_459);
nand U3989 (N_3989,In_616,In_297);
and U3990 (N_3990,In_953,In_509);
nor U3991 (N_3991,In_225,In_896);
nor U3992 (N_3992,In_252,In_118);
or U3993 (N_3993,In_982,In_829);
or U3994 (N_3994,In_154,In_591);
nor U3995 (N_3995,In_610,In_777);
nor U3996 (N_3996,In_100,In_665);
and U3997 (N_3997,In_965,In_34);
nand U3998 (N_3998,In_204,In_950);
and U3999 (N_3999,In_303,In_246);
or U4000 (N_4000,In_446,In_608);
or U4001 (N_4001,In_230,In_29);
or U4002 (N_4002,In_453,In_193);
and U4003 (N_4003,In_228,In_747);
xor U4004 (N_4004,In_416,In_659);
nand U4005 (N_4005,In_117,In_471);
or U4006 (N_4006,In_17,In_755);
nor U4007 (N_4007,In_219,In_117);
nor U4008 (N_4008,In_578,In_0);
nand U4009 (N_4009,In_286,In_558);
nor U4010 (N_4010,In_764,In_194);
xor U4011 (N_4011,In_65,In_880);
and U4012 (N_4012,In_350,In_797);
or U4013 (N_4013,In_249,In_288);
and U4014 (N_4014,In_29,In_60);
and U4015 (N_4015,In_323,In_159);
or U4016 (N_4016,In_122,In_26);
nand U4017 (N_4017,In_913,In_615);
and U4018 (N_4018,In_880,In_486);
nor U4019 (N_4019,In_573,In_116);
and U4020 (N_4020,In_496,In_309);
nor U4021 (N_4021,In_291,In_147);
nand U4022 (N_4022,In_190,In_170);
nor U4023 (N_4023,In_628,In_205);
nor U4024 (N_4024,In_279,In_13);
nor U4025 (N_4025,In_258,In_456);
nor U4026 (N_4026,In_530,In_66);
nand U4027 (N_4027,In_999,In_597);
nand U4028 (N_4028,In_3,In_788);
or U4029 (N_4029,In_907,In_862);
nand U4030 (N_4030,In_677,In_927);
nand U4031 (N_4031,In_819,In_629);
nor U4032 (N_4032,In_150,In_443);
and U4033 (N_4033,In_267,In_252);
nand U4034 (N_4034,In_759,In_200);
nand U4035 (N_4035,In_74,In_934);
nor U4036 (N_4036,In_744,In_715);
nor U4037 (N_4037,In_139,In_359);
nand U4038 (N_4038,In_963,In_824);
and U4039 (N_4039,In_376,In_649);
nor U4040 (N_4040,In_803,In_3);
nor U4041 (N_4041,In_271,In_273);
nor U4042 (N_4042,In_170,In_761);
nor U4043 (N_4043,In_783,In_289);
and U4044 (N_4044,In_529,In_922);
nor U4045 (N_4045,In_513,In_699);
nand U4046 (N_4046,In_367,In_7);
or U4047 (N_4047,In_104,In_919);
or U4048 (N_4048,In_623,In_582);
nand U4049 (N_4049,In_679,In_461);
and U4050 (N_4050,In_745,In_719);
and U4051 (N_4051,In_303,In_591);
nor U4052 (N_4052,In_959,In_401);
nor U4053 (N_4053,In_864,In_749);
or U4054 (N_4054,In_565,In_183);
and U4055 (N_4055,In_258,In_482);
or U4056 (N_4056,In_59,In_402);
or U4057 (N_4057,In_614,In_865);
and U4058 (N_4058,In_190,In_277);
or U4059 (N_4059,In_707,In_36);
or U4060 (N_4060,In_347,In_251);
nand U4061 (N_4061,In_367,In_177);
nor U4062 (N_4062,In_787,In_470);
nand U4063 (N_4063,In_878,In_931);
nand U4064 (N_4064,In_490,In_455);
xor U4065 (N_4065,In_977,In_790);
and U4066 (N_4066,In_36,In_969);
or U4067 (N_4067,In_670,In_671);
and U4068 (N_4068,In_366,In_586);
or U4069 (N_4069,In_837,In_411);
nand U4070 (N_4070,In_771,In_414);
or U4071 (N_4071,In_952,In_841);
nor U4072 (N_4072,In_956,In_123);
nand U4073 (N_4073,In_701,In_934);
or U4074 (N_4074,In_463,In_662);
and U4075 (N_4075,In_82,In_204);
and U4076 (N_4076,In_151,In_719);
nor U4077 (N_4077,In_121,In_754);
xor U4078 (N_4078,In_126,In_680);
xnor U4079 (N_4079,In_989,In_988);
nor U4080 (N_4080,In_85,In_379);
nand U4081 (N_4081,In_639,In_139);
xnor U4082 (N_4082,In_688,In_331);
and U4083 (N_4083,In_349,In_193);
and U4084 (N_4084,In_990,In_968);
nor U4085 (N_4085,In_119,In_467);
or U4086 (N_4086,In_108,In_322);
and U4087 (N_4087,In_572,In_51);
or U4088 (N_4088,In_885,In_676);
nor U4089 (N_4089,In_793,In_468);
or U4090 (N_4090,In_213,In_406);
nor U4091 (N_4091,In_871,In_80);
xor U4092 (N_4092,In_145,In_478);
nor U4093 (N_4093,In_614,In_897);
nand U4094 (N_4094,In_116,In_971);
nand U4095 (N_4095,In_264,In_270);
and U4096 (N_4096,In_817,In_900);
nor U4097 (N_4097,In_255,In_688);
nand U4098 (N_4098,In_570,In_202);
nand U4099 (N_4099,In_265,In_211);
nand U4100 (N_4100,In_974,In_322);
nand U4101 (N_4101,In_932,In_885);
nand U4102 (N_4102,In_497,In_280);
and U4103 (N_4103,In_453,In_382);
xor U4104 (N_4104,In_882,In_171);
and U4105 (N_4105,In_927,In_628);
nor U4106 (N_4106,In_151,In_247);
nor U4107 (N_4107,In_496,In_641);
nor U4108 (N_4108,In_589,In_750);
nand U4109 (N_4109,In_178,In_605);
or U4110 (N_4110,In_350,In_755);
nand U4111 (N_4111,In_583,In_116);
xnor U4112 (N_4112,In_888,In_617);
or U4113 (N_4113,In_289,In_801);
and U4114 (N_4114,In_463,In_870);
xnor U4115 (N_4115,In_972,In_436);
and U4116 (N_4116,In_401,In_603);
nand U4117 (N_4117,In_737,In_272);
nand U4118 (N_4118,In_443,In_127);
xnor U4119 (N_4119,In_219,In_170);
and U4120 (N_4120,In_153,In_845);
or U4121 (N_4121,In_475,In_599);
nor U4122 (N_4122,In_284,In_602);
nand U4123 (N_4123,In_122,In_492);
and U4124 (N_4124,In_903,In_787);
and U4125 (N_4125,In_561,In_720);
or U4126 (N_4126,In_637,In_822);
nor U4127 (N_4127,In_938,In_836);
or U4128 (N_4128,In_375,In_787);
and U4129 (N_4129,In_613,In_83);
and U4130 (N_4130,In_781,In_398);
nand U4131 (N_4131,In_709,In_440);
nor U4132 (N_4132,In_31,In_27);
nand U4133 (N_4133,In_389,In_171);
and U4134 (N_4134,In_42,In_308);
or U4135 (N_4135,In_8,In_622);
or U4136 (N_4136,In_255,In_307);
nor U4137 (N_4137,In_648,In_775);
nor U4138 (N_4138,In_623,In_73);
nand U4139 (N_4139,In_961,In_481);
or U4140 (N_4140,In_87,In_135);
nor U4141 (N_4141,In_797,In_598);
nand U4142 (N_4142,In_748,In_820);
nand U4143 (N_4143,In_960,In_916);
nand U4144 (N_4144,In_734,In_635);
and U4145 (N_4145,In_386,In_312);
and U4146 (N_4146,In_479,In_982);
and U4147 (N_4147,In_576,In_291);
nor U4148 (N_4148,In_489,In_689);
nand U4149 (N_4149,In_467,In_855);
and U4150 (N_4150,In_621,In_472);
and U4151 (N_4151,In_364,In_872);
nand U4152 (N_4152,In_598,In_943);
nand U4153 (N_4153,In_607,In_449);
nor U4154 (N_4154,In_905,In_521);
nor U4155 (N_4155,In_893,In_947);
xnor U4156 (N_4156,In_312,In_39);
or U4157 (N_4157,In_754,In_702);
and U4158 (N_4158,In_808,In_466);
and U4159 (N_4159,In_96,In_486);
or U4160 (N_4160,In_412,In_667);
and U4161 (N_4161,In_467,In_708);
or U4162 (N_4162,In_846,In_516);
and U4163 (N_4163,In_441,In_48);
or U4164 (N_4164,In_500,In_205);
nand U4165 (N_4165,In_625,In_577);
xor U4166 (N_4166,In_668,In_620);
and U4167 (N_4167,In_696,In_3);
nand U4168 (N_4168,In_657,In_753);
and U4169 (N_4169,In_159,In_56);
nor U4170 (N_4170,In_578,In_320);
nand U4171 (N_4171,In_832,In_552);
nand U4172 (N_4172,In_709,In_722);
nor U4173 (N_4173,In_894,In_290);
nor U4174 (N_4174,In_645,In_313);
nor U4175 (N_4175,In_979,In_320);
nand U4176 (N_4176,In_314,In_629);
or U4177 (N_4177,In_239,In_219);
or U4178 (N_4178,In_361,In_547);
nor U4179 (N_4179,In_397,In_599);
and U4180 (N_4180,In_446,In_534);
nor U4181 (N_4181,In_758,In_983);
and U4182 (N_4182,In_290,In_197);
nor U4183 (N_4183,In_394,In_55);
nand U4184 (N_4184,In_554,In_403);
nand U4185 (N_4185,In_995,In_288);
or U4186 (N_4186,In_426,In_176);
xor U4187 (N_4187,In_562,In_150);
and U4188 (N_4188,In_275,In_713);
and U4189 (N_4189,In_421,In_554);
or U4190 (N_4190,In_585,In_414);
nand U4191 (N_4191,In_480,In_269);
xor U4192 (N_4192,In_889,In_503);
nor U4193 (N_4193,In_447,In_851);
or U4194 (N_4194,In_631,In_663);
nand U4195 (N_4195,In_856,In_626);
or U4196 (N_4196,In_9,In_386);
nand U4197 (N_4197,In_631,In_911);
or U4198 (N_4198,In_562,In_873);
nand U4199 (N_4199,In_925,In_867);
and U4200 (N_4200,In_49,In_218);
nor U4201 (N_4201,In_178,In_506);
nor U4202 (N_4202,In_355,In_567);
and U4203 (N_4203,In_451,In_66);
and U4204 (N_4204,In_412,In_814);
nand U4205 (N_4205,In_401,In_29);
and U4206 (N_4206,In_197,In_768);
nand U4207 (N_4207,In_651,In_466);
and U4208 (N_4208,In_147,In_245);
nor U4209 (N_4209,In_867,In_407);
and U4210 (N_4210,In_409,In_708);
or U4211 (N_4211,In_24,In_760);
and U4212 (N_4212,In_78,In_447);
nor U4213 (N_4213,In_60,In_622);
nor U4214 (N_4214,In_124,In_704);
or U4215 (N_4215,In_128,In_385);
nand U4216 (N_4216,In_124,In_144);
and U4217 (N_4217,In_71,In_542);
or U4218 (N_4218,In_499,In_407);
and U4219 (N_4219,In_986,In_488);
nand U4220 (N_4220,In_950,In_326);
or U4221 (N_4221,In_754,In_95);
and U4222 (N_4222,In_19,In_947);
nand U4223 (N_4223,In_855,In_362);
and U4224 (N_4224,In_800,In_164);
nor U4225 (N_4225,In_919,In_115);
and U4226 (N_4226,In_961,In_464);
nor U4227 (N_4227,In_286,In_89);
and U4228 (N_4228,In_323,In_926);
nand U4229 (N_4229,In_847,In_245);
and U4230 (N_4230,In_161,In_490);
nand U4231 (N_4231,In_858,In_632);
nand U4232 (N_4232,In_119,In_341);
and U4233 (N_4233,In_305,In_761);
xnor U4234 (N_4234,In_395,In_270);
nand U4235 (N_4235,In_477,In_903);
nand U4236 (N_4236,In_72,In_56);
nand U4237 (N_4237,In_446,In_335);
or U4238 (N_4238,In_336,In_32);
nor U4239 (N_4239,In_806,In_309);
nand U4240 (N_4240,In_870,In_533);
or U4241 (N_4241,In_554,In_778);
and U4242 (N_4242,In_463,In_467);
and U4243 (N_4243,In_338,In_953);
nand U4244 (N_4244,In_941,In_43);
nand U4245 (N_4245,In_211,In_580);
nand U4246 (N_4246,In_593,In_921);
nor U4247 (N_4247,In_865,In_800);
nand U4248 (N_4248,In_260,In_996);
nor U4249 (N_4249,In_13,In_453);
xnor U4250 (N_4250,In_468,In_85);
nand U4251 (N_4251,In_599,In_385);
xnor U4252 (N_4252,In_408,In_156);
and U4253 (N_4253,In_672,In_52);
and U4254 (N_4254,In_840,In_147);
xor U4255 (N_4255,In_346,In_914);
nor U4256 (N_4256,In_691,In_42);
nor U4257 (N_4257,In_799,In_768);
nand U4258 (N_4258,In_478,In_119);
xor U4259 (N_4259,In_60,In_970);
nor U4260 (N_4260,In_993,In_672);
nand U4261 (N_4261,In_866,In_956);
xor U4262 (N_4262,In_84,In_892);
and U4263 (N_4263,In_500,In_312);
nand U4264 (N_4264,In_403,In_125);
xnor U4265 (N_4265,In_77,In_858);
nand U4266 (N_4266,In_617,In_346);
xnor U4267 (N_4267,In_972,In_535);
nand U4268 (N_4268,In_148,In_993);
nand U4269 (N_4269,In_650,In_612);
or U4270 (N_4270,In_421,In_248);
and U4271 (N_4271,In_168,In_203);
or U4272 (N_4272,In_362,In_221);
nor U4273 (N_4273,In_274,In_25);
nor U4274 (N_4274,In_519,In_322);
nor U4275 (N_4275,In_798,In_355);
nand U4276 (N_4276,In_389,In_521);
xor U4277 (N_4277,In_307,In_439);
and U4278 (N_4278,In_224,In_8);
xnor U4279 (N_4279,In_909,In_767);
or U4280 (N_4280,In_887,In_85);
nand U4281 (N_4281,In_401,In_658);
nor U4282 (N_4282,In_348,In_969);
nand U4283 (N_4283,In_387,In_722);
nand U4284 (N_4284,In_130,In_744);
nand U4285 (N_4285,In_430,In_408);
nand U4286 (N_4286,In_695,In_483);
or U4287 (N_4287,In_219,In_625);
and U4288 (N_4288,In_934,In_897);
and U4289 (N_4289,In_899,In_424);
xnor U4290 (N_4290,In_736,In_879);
and U4291 (N_4291,In_815,In_630);
or U4292 (N_4292,In_871,In_451);
and U4293 (N_4293,In_395,In_652);
nand U4294 (N_4294,In_658,In_974);
nand U4295 (N_4295,In_395,In_982);
and U4296 (N_4296,In_545,In_481);
and U4297 (N_4297,In_135,In_850);
or U4298 (N_4298,In_798,In_245);
nand U4299 (N_4299,In_383,In_902);
and U4300 (N_4300,In_887,In_639);
nand U4301 (N_4301,In_639,In_76);
xnor U4302 (N_4302,In_622,In_526);
xor U4303 (N_4303,In_110,In_569);
nor U4304 (N_4304,In_304,In_41);
and U4305 (N_4305,In_30,In_604);
or U4306 (N_4306,In_298,In_313);
nand U4307 (N_4307,In_931,In_958);
nor U4308 (N_4308,In_423,In_435);
xor U4309 (N_4309,In_105,In_842);
nor U4310 (N_4310,In_187,In_503);
and U4311 (N_4311,In_701,In_919);
xnor U4312 (N_4312,In_933,In_977);
nor U4313 (N_4313,In_439,In_914);
xnor U4314 (N_4314,In_663,In_9);
nand U4315 (N_4315,In_766,In_621);
nor U4316 (N_4316,In_675,In_723);
or U4317 (N_4317,In_235,In_568);
nand U4318 (N_4318,In_566,In_20);
or U4319 (N_4319,In_770,In_681);
nand U4320 (N_4320,In_244,In_460);
nand U4321 (N_4321,In_866,In_916);
xnor U4322 (N_4322,In_86,In_484);
nand U4323 (N_4323,In_367,In_258);
and U4324 (N_4324,In_304,In_637);
and U4325 (N_4325,In_330,In_608);
xnor U4326 (N_4326,In_448,In_106);
or U4327 (N_4327,In_761,In_737);
nor U4328 (N_4328,In_393,In_155);
nor U4329 (N_4329,In_438,In_760);
or U4330 (N_4330,In_945,In_678);
and U4331 (N_4331,In_134,In_880);
or U4332 (N_4332,In_514,In_700);
xor U4333 (N_4333,In_944,In_809);
xor U4334 (N_4334,In_627,In_355);
or U4335 (N_4335,In_371,In_386);
nand U4336 (N_4336,In_286,In_818);
nand U4337 (N_4337,In_82,In_538);
and U4338 (N_4338,In_709,In_611);
xor U4339 (N_4339,In_752,In_568);
and U4340 (N_4340,In_861,In_43);
and U4341 (N_4341,In_345,In_355);
and U4342 (N_4342,In_413,In_512);
nor U4343 (N_4343,In_36,In_795);
and U4344 (N_4344,In_645,In_634);
or U4345 (N_4345,In_550,In_559);
xnor U4346 (N_4346,In_714,In_872);
nand U4347 (N_4347,In_709,In_392);
nand U4348 (N_4348,In_643,In_457);
and U4349 (N_4349,In_878,In_363);
nor U4350 (N_4350,In_476,In_438);
xnor U4351 (N_4351,In_453,In_897);
and U4352 (N_4352,In_626,In_403);
and U4353 (N_4353,In_139,In_877);
and U4354 (N_4354,In_470,In_696);
nand U4355 (N_4355,In_313,In_910);
or U4356 (N_4356,In_7,In_648);
nor U4357 (N_4357,In_460,In_918);
or U4358 (N_4358,In_238,In_142);
nand U4359 (N_4359,In_594,In_125);
nand U4360 (N_4360,In_960,In_404);
or U4361 (N_4361,In_452,In_704);
xor U4362 (N_4362,In_926,In_210);
xor U4363 (N_4363,In_764,In_243);
and U4364 (N_4364,In_114,In_463);
and U4365 (N_4365,In_743,In_217);
and U4366 (N_4366,In_823,In_945);
or U4367 (N_4367,In_544,In_53);
and U4368 (N_4368,In_412,In_341);
or U4369 (N_4369,In_314,In_304);
and U4370 (N_4370,In_598,In_712);
nor U4371 (N_4371,In_701,In_564);
nor U4372 (N_4372,In_362,In_511);
nand U4373 (N_4373,In_788,In_583);
and U4374 (N_4374,In_592,In_550);
and U4375 (N_4375,In_416,In_678);
or U4376 (N_4376,In_227,In_964);
nor U4377 (N_4377,In_91,In_280);
nor U4378 (N_4378,In_208,In_503);
xnor U4379 (N_4379,In_724,In_352);
xnor U4380 (N_4380,In_556,In_983);
nand U4381 (N_4381,In_943,In_804);
xor U4382 (N_4382,In_982,In_905);
nand U4383 (N_4383,In_14,In_364);
or U4384 (N_4384,In_386,In_920);
nand U4385 (N_4385,In_572,In_316);
nor U4386 (N_4386,In_722,In_344);
xor U4387 (N_4387,In_203,In_433);
nor U4388 (N_4388,In_218,In_972);
or U4389 (N_4389,In_982,In_302);
nand U4390 (N_4390,In_137,In_609);
nand U4391 (N_4391,In_325,In_815);
xor U4392 (N_4392,In_560,In_326);
nand U4393 (N_4393,In_795,In_3);
nor U4394 (N_4394,In_403,In_870);
xor U4395 (N_4395,In_762,In_496);
xnor U4396 (N_4396,In_783,In_635);
or U4397 (N_4397,In_761,In_60);
xor U4398 (N_4398,In_56,In_618);
and U4399 (N_4399,In_82,In_559);
or U4400 (N_4400,In_739,In_419);
xnor U4401 (N_4401,In_391,In_11);
or U4402 (N_4402,In_294,In_350);
or U4403 (N_4403,In_553,In_615);
or U4404 (N_4404,In_201,In_838);
xor U4405 (N_4405,In_158,In_531);
xor U4406 (N_4406,In_897,In_563);
nor U4407 (N_4407,In_170,In_83);
or U4408 (N_4408,In_94,In_552);
and U4409 (N_4409,In_724,In_857);
xor U4410 (N_4410,In_134,In_898);
and U4411 (N_4411,In_495,In_524);
nand U4412 (N_4412,In_537,In_826);
and U4413 (N_4413,In_721,In_859);
nor U4414 (N_4414,In_820,In_146);
and U4415 (N_4415,In_331,In_382);
nand U4416 (N_4416,In_166,In_908);
xor U4417 (N_4417,In_945,In_804);
or U4418 (N_4418,In_193,In_392);
nor U4419 (N_4419,In_124,In_768);
nand U4420 (N_4420,In_134,In_414);
nor U4421 (N_4421,In_663,In_84);
or U4422 (N_4422,In_506,In_76);
nand U4423 (N_4423,In_731,In_538);
nand U4424 (N_4424,In_938,In_791);
nor U4425 (N_4425,In_911,In_643);
and U4426 (N_4426,In_988,In_725);
nand U4427 (N_4427,In_751,In_406);
and U4428 (N_4428,In_132,In_756);
or U4429 (N_4429,In_928,In_599);
nand U4430 (N_4430,In_963,In_392);
nor U4431 (N_4431,In_816,In_893);
nand U4432 (N_4432,In_40,In_875);
and U4433 (N_4433,In_933,In_57);
nor U4434 (N_4434,In_206,In_908);
and U4435 (N_4435,In_348,In_264);
nor U4436 (N_4436,In_432,In_401);
nor U4437 (N_4437,In_520,In_808);
and U4438 (N_4438,In_21,In_101);
nor U4439 (N_4439,In_256,In_550);
nor U4440 (N_4440,In_109,In_512);
or U4441 (N_4441,In_535,In_621);
and U4442 (N_4442,In_611,In_827);
or U4443 (N_4443,In_829,In_891);
nand U4444 (N_4444,In_345,In_530);
nand U4445 (N_4445,In_917,In_44);
and U4446 (N_4446,In_165,In_723);
nor U4447 (N_4447,In_888,In_105);
xnor U4448 (N_4448,In_909,In_116);
nor U4449 (N_4449,In_193,In_547);
or U4450 (N_4450,In_316,In_472);
nor U4451 (N_4451,In_778,In_372);
or U4452 (N_4452,In_353,In_733);
nor U4453 (N_4453,In_948,In_144);
and U4454 (N_4454,In_365,In_909);
or U4455 (N_4455,In_341,In_419);
nand U4456 (N_4456,In_842,In_747);
and U4457 (N_4457,In_188,In_760);
nand U4458 (N_4458,In_89,In_685);
xor U4459 (N_4459,In_732,In_848);
and U4460 (N_4460,In_533,In_866);
or U4461 (N_4461,In_643,In_840);
xor U4462 (N_4462,In_804,In_548);
nand U4463 (N_4463,In_498,In_71);
or U4464 (N_4464,In_817,In_284);
nor U4465 (N_4465,In_94,In_509);
or U4466 (N_4466,In_774,In_953);
and U4467 (N_4467,In_416,In_61);
or U4468 (N_4468,In_158,In_218);
and U4469 (N_4469,In_329,In_286);
and U4470 (N_4470,In_936,In_179);
nand U4471 (N_4471,In_828,In_939);
nand U4472 (N_4472,In_845,In_686);
nor U4473 (N_4473,In_739,In_481);
xnor U4474 (N_4474,In_553,In_913);
nand U4475 (N_4475,In_512,In_591);
or U4476 (N_4476,In_615,In_320);
xor U4477 (N_4477,In_780,In_29);
nor U4478 (N_4478,In_628,In_969);
nor U4479 (N_4479,In_357,In_926);
nand U4480 (N_4480,In_511,In_183);
and U4481 (N_4481,In_998,In_775);
nor U4482 (N_4482,In_939,In_538);
and U4483 (N_4483,In_248,In_415);
nand U4484 (N_4484,In_404,In_269);
xor U4485 (N_4485,In_626,In_591);
nor U4486 (N_4486,In_880,In_189);
or U4487 (N_4487,In_912,In_992);
and U4488 (N_4488,In_645,In_743);
and U4489 (N_4489,In_676,In_259);
and U4490 (N_4490,In_99,In_363);
nand U4491 (N_4491,In_239,In_213);
or U4492 (N_4492,In_392,In_528);
and U4493 (N_4493,In_441,In_664);
xnor U4494 (N_4494,In_492,In_191);
or U4495 (N_4495,In_450,In_34);
nor U4496 (N_4496,In_497,In_625);
nor U4497 (N_4497,In_433,In_880);
nand U4498 (N_4498,In_986,In_412);
nand U4499 (N_4499,In_436,In_355);
nand U4500 (N_4500,In_307,In_786);
nand U4501 (N_4501,In_469,In_85);
and U4502 (N_4502,In_331,In_535);
nand U4503 (N_4503,In_729,In_734);
nand U4504 (N_4504,In_397,In_579);
and U4505 (N_4505,In_831,In_24);
and U4506 (N_4506,In_174,In_899);
nand U4507 (N_4507,In_744,In_838);
nor U4508 (N_4508,In_848,In_596);
or U4509 (N_4509,In_650,In_7);
and U4510 (N_4510,In_465,In_801);
and U4511 (N_4511,In_593,In_661);
and U4512 (N_4512,In_433,In_947);
and U4513 (N_4513,In_137,In_638);
and U4514 (N_4514,In_288,In_374);
xor U4515 (N_4515,In_428,In_793);
nand U4516 (N_4516,In_656,In_630);
nor U4517 (N_4517,In_690,In_837);
and U4518 (N_4518,In_189,In_455);
nand U4519 (N_4519,In_270,In_256);
nand U4520 (N_4520,In_795,In_904);
nand U4521 (N_4521,In_287,In_974);
nand U4522 (N_4522,In_747,In_786);
and U4523 (N_4523,In_387,In_49);
nand U4524 (N_4524,In_41,In_509);
xnor U4525 (N_4525,In_531,In_807);
xnor U4526 (N_4526,In_653,In_878);
and U4527 (N_4527,In_700,In_405);
nand U4528 (N_4528,In_970,In_619);
and U4529 (N_4529,In_676,In_858);
or U4530 (N_4530,In_850,In_344);
nor U4531 (N_4531,In_24,In_375);
nand U4532 (N_4532,In_918,In_608);
and U4533 (N_4533,In_894,In_127);
and U4534 (N_4534,In_566,In_923);
and U4535 (N_4535,In_228,In_217);
or U4536 (N_4536,In_824,In_156);
nand U4537 (N_4537,In_510,In_75);
or U4538 (N_4538,In_525,In_756);
nand U4539 (N_4539,In_939,In_868);
nand U4540 (N_4540,In_395,In_95);
and U4541 (N_4541,In_951,In_581);
or U4542 (N_4542,In_402,In_428);
and U4543 (N_4543,In_476,In_167);
or U4544 (N_4544,In_215,In_154);
or U4545 (N_4545,In_138,In_600);
xnor U4546 (N_4546,In_155,In_339);
or U4547 (N_4547,In_764,In_921);
and U4548 (N_4548,In_901,In_278);
or U4549 (N_4549,In_542,In_961);
nor U4550 (N_4550,In_609,In_739);
nand U4551 (N_4551,In_749,In_228);
xor U4552 (N_4552,In_380,In_586);
xnor U4553 (N_4553,In_277,In_805);
nor U4554 (N_4554,In_919,In_993);
nor U4555 (N_4555,In_524,In_648);
nor U4556 (N_4556,In_249,In_451);
and U4557 (N_4557,In_599,In_393);
nor U4558 (N_4558,In_438,In_545);
xnor U4559 (N_4559,In_366,In_773);
and U4560 (N_4560,In_347,In_253);
nor U4561 (N_4561,In_966,In_801);
xor U4562 (N_4562,In_821,In_298);
nand U4563 (N_4563,In_817,In_176);
nor U4564 (N_4564,In_558,In_808);
nor U4565 (N_4565,In_600,In_401);
nand U4566 (N_4566,In_375,In_181);
nand U4567 (N_4567,In_52,In_689);
and U4568 (N_4568,In_945,In_647);
xnor U4569 (N_4569,In_326,In_953);
nand U4570 (N_4570,In_308,In_817);
and U4571 (N_4571,In_542,In_344);
and U4572 (N_4572,In_478,In_425);
xnor U4573 (N_4573,In_75,In_748);
nand U4574 (N_4574,In_950,In_376);
or U4575 (N_4575,In_6,In_920);
nor U4576 (N_4576,In_4,In_164);
nand U4577 (N_4577,In_496,In_144);
or U4578 (N_4578,In_119,In_488);
nand U4579 (N_4579,In_291,In_622);
or U4580 (N_4580,In_398,In_579);
or U4581 (N_4581,In_363,In_753);
and U4582 (N_4582,In_135,In_299);
xnor U4583 (N_4583,In_67,In_104);
nand U4584 (N_4584,In_847,In_246);
xnor U4585 (N_4585,In_0,In_709);
or U4586 (N_4586,In_582,In_925);
and U4587 (N_4587,In_468,In_934);
nor U4588 (N_4588,In_372,In_660);
or U4589 (N_4589,In_713,In_82);
or U4590 (N_4590,In_408,In_805);
xnor U4591 (N_4591,In_801,In_938);
nand U4592 (N_4592,In_186,In_674);
nand U4593 (N_4593,In_988,In_23);
or U4594 (N_4594,In_931,In_630);
nor U4595 (N_4595,In_586,In_261);
nor U4596 (N_4596,In_406,In_693);
nand U4597 (N_4597,In_480,In_746);
nor U4598 (N_4598,In_320,In_692);
nor U4599 (N_4599,In_173,In_592);
or U4600 (N_4600,In_930,In_884);
xnor U4601 (N_4601,In_838,In_288);
and U4602 (N_4602,In_49,In_320);
nand U4603 (N_4603,In_836,In_290);
or U4604 (N_4604,In_637,In_769);
nand U4605 (N_4605,In_655,In_154);
and U4606 (N_4606,In_19,In_998);
nor U4607 (N_4607,In_442,In_597);
and U4608 (N_4608,In_871,In_603);
xnor U4609 (N_4609,In_384,In_300);
nor U4610 (N_4610,In_207,In_847);
nor U4611 (N_4611,In_503,In_553);
nand U4612 (N_4612,In_213,In_166);
nand U4613 (N_4613,In_891,In_475);
nand U4614 (N_4614,In_814,In_80);
nand U4615 (N_4615,In_349,In_162);
or U4616 (N_4616,In_487,In_57);
nand U4617 (N_4617,In_119,In_349);
or U4618 (N_4618,In_18,In_340);
or U4619 (N_4619,In_229,In_838);
xnor U4620 (N_4620,In_894,In_230);
nor U4621 (N_4621,In_759,In_884);
and U4622 (N_4622,In_114,In_48);
and U4623 (N_4623,In_841,In_775);
or U4624 (N_4624,In_87,In_974);
and U4625 (N_4625,In_168,In_284);
nand U4626 (N_4626,In_230,In_310);
or U4627 (N_4627,In_204,In_267);
or U4628 (N_4628,In_137,In_849);
nor U4629 (N_4629,In_611,In_720);
nand U4630 (N_4630,In_791,In_454);
and U4631 (N_4631,In_234,In_851);
and U4632 (N_4632,In_460,In_354);
xnor U4633 (N_4633,In_324,In_934);
nand U4634 (N_4634,In_380,In_709);
nand U4635 (N_4635,In_859,In_88);
or U4636 (N_4636,In_770,In_298);
nand U4637 (N_4637,In_576,In_527);
nand U4638 (N_4638,In_602,In_267);
nor U4639 (N_4639,In_136,In_66);
and U4640 (N_4640,In_599,In_860);
or U4641 (N_4641,In_493,In_470);
and U4642 (N_4642,In_158,In_437);
and U4643 (N_4643,In_620,In_293);
nand U4644 (N_4644,In_16,In_383);
nand U4645 (N_4645,In_667,In_732);
and U4646 (N_4646,In_914,In_626);
nand U4647 (N_4647,In_785,In_642);
nand U4648 (N_4648,In_489,In_808);
or U4649 (N_4649,In_631,In_478);
and U4650 (N_4650,In_594,In_415);
nand U4651 (N_4651,In_115,In_704);
nand U4652 (N_4652,In_921,In_831);
nand U4653 (N_4653,In_191,In_507);
nor U4654 (N_4654,In_900,In_108);
and U4655 (N_4655,In_694,In_478);
and U4656 (N_4656,In_907,In_495);
nor U4657 (N_4657,In_95,In_64);
nor U4658 (N_4658,In_710,In_654);
and U4659 (N_4659,In_619,In_643);
or U4660 (N_4660,In_83,In_227);
nor U4661 (N_4661,In_876,In_652);
or U4662 (N_4662,In_989,In_544);
and U4663 (N_4663,In_457,In_300);
or U4664 (N_4664,In_219,In_846);
nor U4665 (N_4665,In_691,In_504);
nor U4666 (N_4666,In_373,In_995);
nand U4667 (N_4667,In_357,In_310);
nand U4668 (N_4668,In_84,In_886);
nand U4669 (N_4669,In_75,In_639);
and U4670 (N_4670,In_630,In_216);
or U4671 (N_4671,In_35,In_203);
nor U4672 (N_4672,In_391,In_392);
nand U4673 (N_4673,In_304,In_243);
xnor U4674 (N_4674,In_237,In_249);
and U4675 (N_4675,In_73,In_589);
and U4676 (N_4676,In_107,In_815);
nand U4677 (N_4677,In_813,In_44);
nand U4678 (N_4678,In_349,In_729);
and U4679 (N_4679,In_113,In_695);
xnor U4680 (N_4680,In_32,In_972);
nand U4681 (N_4681,In_490,In_384);
nand U4682 (N_4682,In_775,In_134);
and U4683 (N_4683,In_709,In_544);
nor U4684 (N_4684,In_932,In_616);
nor U4685 (N_4685,In_110,In_744);
or U4686 (N_4686,In_683,In_618);
or U4687 (N_4687,In_846,In_984);
nor U4688 (N_4688,In_681,In_606);
nand U4689 (N_4689,In_436,In_675);
and U4690 (N_4690,In_775,In_67);
or U4691 (N_4691,In_505,In_76);
and U4692 (N_4692,In_343,In_139);
or U4693 (N_4693,In_294,In_361);
nor U4694 (N_4694,In_503,In_254);
and U4695 (N_4695,In_720,In_878);
and U4696 (N_4696,In_146,In_221);
nand U4697 (N_4697,In_772,In_669);
or U4698 (N_4698,In_794,In_950);
nand U4699 (N_4699,In_977,In_899);
nand U4700 (N_4700,In_111,In_22);
nand U4701 (N_4701,In_917,In_437);
nor U4702 (N_4702,In_187,In_980);
or U4703 (N_4703,In_151,In_433);
nand U4704 (N_4704,In_740,In_811);
nand U4705 (N_4705,In_429,In_852);
nand U4706 (N_4706,In_228,In_765);
and U4707 (N_4707,In_539,In_89);
nand U4708 (N_4708,In_604,In_797);
or U4709 (N_4709,In_576,In_373);
or U4710 (N_4710,In_673,In_557);
and U4711 (N_4711,In_625,In_369);
nor U4712 (N_4712,In_671,In_655);
or U4713 (N_4713,In_915,In_587);
or U4714 (N_4714,In_610,In_121);
nor U4715 (N_4715,In_11,In_977);
nand U4716 (N_4716,In_257,In_124);
or U4717 (N_4717,In_379,In_247);
and U4718 (N_4718,In_107,In_968);
nand U4719 (N_4719,In_883,In_997);
nor U4720 (N_4720,In_462,In_823);
and U4721 (N_4721,In_721,In_256);
nor U4722 (N_4722,In_246,In_637);
or U4723 (N_4723,In_253,In_460);
nand U4724 (N_4724,In_804,In_8);
and U4725 (N_4725,In_506,In_330);
or U4726 (N_4726,In_431,In_220);
and U4727 (N_4727,In_87,In_981);
nand U4728 (N_4728,In_112,In_864);
and U4729 (N_4729,In_989,In_402);
and U4730 (N_4730,In_171,In_183);
nand U4731 (N_4731,In_345,In_633);
nor U4732 (N_4732,In_69,In_183);
or U4733 (N_4733,In_300,In_286);
nand U4734 (N_4734,In_62,In_203);
nor U4735 (N_4735,In_56,In_201);
nor U4736 (N_4736,In_152,In_450);
nor U4737 (N_4737,In_603,In_515);
or U4738 (N_4738,In_458,In_934);
nor U4739 (N_4739,In_594,In_665);
xor U4740 (N_4740,In_317,In_497);
nand U4741 (N_4741,In_92,In_538);
and U4742 (N_4742,In_150,In_967);
or U4743 (N_4743,In_319,In_800);
and U4744 (N_4744,In_405,In_799);
xnor U4745 (N_4745,In_869,In_137);
and U4746 (N_4746,In_920,In_13);
and U4747 (N_4747,In_850,In_34);
or U4748 (N_4748,In_864,In_372);
or U4749 (N_4749,In_511,In_715);
xor U4750 (N_4750,In_808,In_681);
nand U4751 (N_4751,In_858,In_903);
nor U4752 (N_4752,In_432,In_121);
and U4753 (N_4753,In_748,In_688);
nand U4754 (N_4754,In_723,In_343);
nor U4755 (N_4755,In_107,In_582);
and U4756 (N_4756,In_499,In_84);
xor U4757 (N_4757,In_979,In_759);
or U4758 (N_4758,In_417,In_210);
nand U4759 (N_4759,In_196,In_889);
nand U4760 (N_4760,In_927,In_265);
xnor U4761 (N_4761,In_886,In_69);
nand U4762 (N_4762,In_821,In_184);
and U4763 (N_4763,In_805,In_18);
xor U4764 (N_4764,In_880,In_593);
and U4765 (N_4765,In_724,In_555);
xor U4766 (N_4766,In_104,In_733);
or U4767 (N_4767,In_205,In_84);
or U4768 (N_4768,In_118,In_389);
nand U4769 (N_4769,In_407,In_188);
or U4770 (N_4770,In_308,In_169);
or U4771 (N_4771,In_146,In_415);
nor U4772 (N_4772,In_6,In_239);
nand U4773 (N_4773,In_528,In_674);
or U4774 (N_4774,In_793,In_470);
and U4775 (N_4775,In_364,In_819);
or U4776 (N_4776,In_759,In_374);
xor U4777 (N_4777,In_713,In_625);
nand U4778 (N_4778,In_670,In_130);
or U4779 (N_4779,In_655,In_776);
or U4780 (N_4780,In_646,In_874);
nor U4781 (N_4781,In_515,In_269);
or U4782 (N_4782,In_62,In_246);
and U4783 (N_4783,In_529,In_799);
nand U4784 (N_4784,In_154,In_413);
or U4785 (N_4785,In_310,In_3);
nand U4786 (N_4786,In_764,In_926);
xnor U4787 (N_4787,In_362,In_37);
and U4788 (N_4788,In_617,In_533);
or U4789 (N_4789,In_669,In_540);
or U4790 (N_4790,In_43,In_97);
nand U4791 (N_4791,In_713,In_541);
and U4792 (N_4792,In_892,In_924);
or U4793 (N_4793,In_632,In_159);
or U4794 (N_4794,In_447,In_626);
nand U4795 (N_4795,In_282,In_30);
and U4796 (N_4796,In_840,In_153);
or U4797 (N_4797,In_604,In_558);
and U4798 (N_4798,In_547,In_969);
or U4799 (N_4799,In_9,In_804);
or U4800 (N_4800,In_339,In_168);
nor U4801 (N_4801,In_714,In_787);
or U4802 (N_4802,In_753,In_608);
or U4803 (N_4803,In_533,In_353);
nor U4804 (N_4804,In_149,In_267);
nor U4805 (N_4805,In_338,In_69);
or U4806 (N_4806,In_278,In_314);
nand U4807 (N_4807,In_512,In_753);
and U4808 (N_4808,In_429,In_356);
nor U4809 (N_4809,In_471,In_48);
and U4810 (N_4810,In_567,In_345);
xor U4811 (N_4811,In_132,In_449);
nand U4812 (N_4812,In_983,In_262);
or U4813 (N_4813,In_955,In_641);
or U4814 (N_4814,In_886,In_270);
and U4815 (N_4815,In_263,In_770);
nor U4816 (N_4816,In_341,In_409);
nor U4817 (N_4817,In_406,In_477);
nand U4818 (N_4818,In_920,In_74);
nor U4819 (N_4819,In_243,In_471);
or U4820 (N_4820,In_676,In_36);
xnor U4821 (N_4821,In_558,In_941);
nand U4822 (N_4822,In_61,In_625);
and U4823 (N_4823,In_56,In_841);
xnor U4824 (N_4824,In_537,In_20);
or U4825 (N_4825,In_157,In_178);
xnor U4826 (N_4826,In_12,In_727);
or U4827 (N_4827,In_952,In_581);
nor U4828 (N_4828,In_818,In_219);
or U4829 (N_4829,In_981,In_847);
nand U4830 (N_4830,In_523,In_722);
xnor U4831 (N_4831,In_516,In_649);
nand U4832 (N_4832,In_628,In_166);
or U4833 (N_4833,In_471,In_400);
or U4834 (N_4834,In_311,In_810);
nor U4835 (N_4835,In_458,In_577);
or U4836 (N_4836,In_873,In_379);
or U4837 (N_4837,In_809,In_929);
nor U4838 (N_4838,In_339,In_115);
nor U4839 (N_4839,In_580,In_147);
xnor U4840 (N_4840,In_324,In_997);
xor U4841 (N_4841,In_933,In_885);
and U4842 (N_4842,In_79,In_723);
nor U4843 (N_4843,In_200,In_743);
nand U4844 (N_4844,In_935,In_737);
nand U4845 (N_4845,In_422,In_382);
or U4846 (N_4846,In_574,In_13);
xor U4847 (N_4847,In_627,In_99);
and U4848 (N_4848,In_585,In_211);
nand U4849 (N_4849,In_945,In_653);
or U4850 (N_4850,In_267,In_794);
xor U4851 (N_4851,In_792,In_915);
nor U4852 (N_4852,In_76,In_288);
or U4853 (N_4853,In_201,In_746);
and U4854 (N_4854,In_309,In_491);
and U4855 (N_4855,In_136,In_430);
nor U4856 (N_4856,In_192,In_293);
and U4857 (N_4857,In_276,In_896);
nor U4858 (N_4858,In_100,In_828);
and U4859 (N_4859,In_21,In_499);
nand U4860 (N_4860,In_372,In_810);
nor U4861 (N_4861,In_759,In_277);
and U4862 (N_4862,In_363,In_297);
nand U4863 (N_4863,In_686,In_112);
nand U4864 (N_4864,In_926,In_569);
nor U4865 (N_4865,In_892,In_63);
xnor U4866 (N_4866,In_631,In_50);
xor U4867 (N_4867,In_306,In_184);
nor U4868 (N_4868,In_416,In_250);
nand U4869 (N_4869,In_38,In_476);
xnor U4870 (N_4870,In_871,In_10);
or U4871 (N_4871,In_604,In_909);
and U4872 (N_4872,In_30,In_563);
nor U4873 (N_4873,In_538,In_511);
nand U4874 (N_4874,In_283,In_79);
xor U4875 (N_4875,In_506,In_423);
nor U4876 (N_4876,In_946,In_902);
and U4877 (N_4877,In_51,In_275);
nor U4878 (N_4878,In_572,In_630);
or U4879 (N_4879,In_305,In_10);
or U4880 (N_4880,In_432,In_657);
and U4881 (N_4881,In_58,In_41);
and U4882 (N_4882,In_819,In_117);
and U4883 (N_4883,In_621,In_550);
or U4884 (N_4884,In_588,In_889);
or U4885 (N_4885,In_296,In_690);
and U4886 (N_4886,In_167,In_468);
and U4887 (N_4887,In_452,In_488);
or U4888 (N_4888,In_515,In_63);
and U4889 (N_4889,In_181,In_255);
nor U4890 (N_4890,In_702,In_420);
and U4891 (N_4891,In_810,In_40);
or U4892 (N_4892,In_585,In_865);
nand U4893 (N_4893,In_1,In_357);
or U4894 (N_4894,In_219,In_456);
xnor U4895 (N_4895,In_741,In_936);
nand U4896 (N_4896,In_353,In_664);
nand U4897 (N_4897,In_230,In_576);
and U4898 (N_4898,In_846,In_311);
nand U4899 (N_4899,In_808,In_693);
nor U4900 (N_4900,In_151,In_196);
nor U4901 (N_4901,In_368,In_590);
and U4902 (N_4902,In_134,In_395);
nand U4903 (N_4903,In_794,In_698);
and U4904 (N_4904,In_618,In_489);
and U4905 (N_4905,In_483,In_572);
nand U4906 (N_4906,In_290,In_427);
nand U4907 (N_4907,In_1,In_454);
xnor U4908 (N_4908,In_637,In_147);
xor U4909 (N_4909,In_291,In_826);
or U4910 (N_4910,In_803,In_483);
and U4911 (N_4911,In_509,In_857);
nand U4912 (N_4912,In_675,In_672);
and U4913 (N_4913,In_310,In_479);
xor U4914 (N_4914,In_124,In_969);
nor U4915 (N_4915,In_864,In_957);
nand U4916 (N_4916,In_380,In_407);
or U4917 (N_4917,In_471,In_856);
nor U4918 (N_4918,In_372,In_295);
xnor U4919 (N_4919,In_228,In_929);
and U4920 (N_4920,In_821,In_156);
or U4921 (N_4921,In_866,In_732);
or U4922 (N_4922,In_557,In_465);
nand U4923 (N_4923,In_182,In_498);
xnor U4924 (N_4924,In_185,In_161);
or U4925 (N_4925,In_750,In_678);
nor U4926 (N_4926,In_925,In_842);
xor U4927 (N_4927,In_244,In_233);
or U4928 (N_4928,In_91,In_735);
or U4929 (N_4929,In_244,In_243);
nand U4930 (N_4930,In_190,In_614);
nand U4931 (N_4931,In_431,In_669);
nand U4932 (N_4932,In_43,In_216);
and U4933 (N_4933,In_186,In_867);
nor U4934 (N_4934,In_733,In_314);
and U4935 (N_4935,In_320,In_746);
nand U4936 (N_4936,In_527,In_477);
or U4937 (N_4937,In_657,In_309);
xor U4938 (N_4938,In_372,In_656);
xor U4939 (N_4939,In_431,In_998);
and U4940 (N_4940,In_505,In_370);
nor U4941 (N_4941,In_808,In_449);
nor U4942 (N_4942,In_313,In_957);
or U4943 (N_4943,In_420,In_976);
nor U4944 (N_4944,In_147,In_505);
or U4945 (N_4945,In_980,In_231);
and U4946 (N_4946,In_373,In_690);
xnor U4947 (N_4947,In_576,In_538);
nand U4948 (N_4948,In_216,In_965);
or U4949 (N_4949,In_66,In_996);
nand U4950 (N_4950,In_635,In_362);
and U4951 (N_4951,In_693,In_961);
nand U4952 (N_4952,In_812,In_302);
xor U4953 (N_4953,In_531,In_119);
or U4954 (N_4954,In_779,In_435);
and U4955 (N_4955,In_185,In_288);
and U4956 (N_4956,In_218,In_163);
nor U4957 (N_4957,In_956,In_817);
nor U4958 (N_4958,In_818,In_233);
or U4959 (N_4959,In_341,In_654);
xor U4960 (N_4960,In_600,In_839);
or U4961 (N_4961,In_813,In_267);
and U4962 (N_4962,In_843,In_220);
and U4963 (N_4963,In_266,In_827);
nor U4964 (N_4964,In_436,In_974);
and U4965 (N_4965,In_550,In_586);
or U4966 (N_4966,In_740,In_586);
nand U4967 (N_4967,In_964,In_927);
nand U4968 (N_4968,In_323,In_877);
xnor U4969 (N_4969,In_27,In_552);
nor U4970 (N_4970,In_154,In_576);
nor U4971 (N_4971,In_220,In_84);
and U4972 (N_4972,In_835,In_748);
and U4973 (N_4973,In_927,In_683);
xnor U4974 (N_4974,In_675,In_776);
nand U4975 (N_4975,In_74,In_229);
or U4976 (N_4976,In_92,In_685);
or U4977 (N_4977,In_981,In_235);
and U4978 (N_4978,In_710,In_790);
xor U4979 (N_4979,In_903,In_212);
xor U4980 (N_4980,In_385,In_163);
and U4981 (N_4981,In_62,In_624);
or U4982 (N_4982,In_122,In_272);
and U4983 (N_4983,In_779,In_529);
or U4984 (N_4984,In_460,In_186);
and U4985 (N_4985,In_391,In_806);
nand U4986 (N_4986,In_858,In_561);
nor U4987 (N_4987,In_446,In_816);
and U4988 (N_4988,In_704,In_969);
or U4989 (N_4989,In_717,In_901);
nor U4990 (N_4990,In_938,In_556);
nor U4991 (N_4991,In_595,In_279);
and U4992 (N_4992,In_707,In_373);
and U4993 (N_4993,In_892,In_855);
nand U4994 (N_4994,In_101,In_290);
nor U4995 (N_4995,In_562,In_250);
nand U4996 (N_4996,In_105,In_132);
nand U4997 (N_4997,In_156,In_838);
and U4998 (N_4998,In_140,In_797);
nand U4999 (N_4999,In_24,In_605);
nor U5000 (N_5000,N_3837,N_3257);
nand U5001 (N_5001,N_899,N_4029);
nand U5002 (N_5002,N_2536,N_878);
or U5003 (N_5003,N_2005,N_2934);
xnor U5004 (N_5004,N_1152,N_3614);
xnor U5005 (N_5005,N_4124,N_2882);
or U5006 (N_5006,N_3990,N_1034);
xor U5007 (N_5007,N_4403,N_2335);
xor U5008 (N_5008,N_1574,N_3073);
nand U5009 (N_5009,N_4069,N_437);
nand U5010 (N_5010,N_3610,N_65);
xnor U5011 (N_5011,N_2630,N_4825);
and U5012 (N_5012,N_4420,N_2166);
or U5013 (N_5013,N_317,N_2462);
nor U5014 (N_5014,N_2118,N_3928);
and U5015 (N_5015,N_1354,N_237);
nor U5016 (N_5016,N_3337,N_1584);
nor U5017 (N_5017,N_1198,N_1137);
and U5018 (N_5018,N_2999,N_2574);
xnor U5019 (N_5019,N_4841,N_4437);
nand U5020 (N_5020,N_1712,N_4577);
xor U5021 (N_5021,N_3214,N_2941);
nand U5022 (N_5022,N_4522,N_4008);
xor U5023 (N_5023,N_1104,N_2172);
nand U5024 (N_5024,N_2294,N_2647);
or U5025 (N_5025,N_1070,N_1081);
and U5026 (N_5026,N_2780,N_2827);
or U5027 (N_5027,N_812,N_1059);
nand U5028 (N_5028,N_4478,N_767);
nand U5029 (N_5029,N_4452,N_1901);
nand U5030 (N_5030,N_2487,N_1205);
or U5031 (N_5031,N_3889,N_35);
nand U5032 (N_5032,N_1167,N_3433);
or U5033 (N_5033,N_1475,N_770);
nor U5034 (N_5034,N_2627,N_4674);
and U5035 (N_5035,N_3576,N_2283);
and U5036 (N_5036,N_2730,N_3141);
and U5037 (N_5037,N_4222,N_738);
or U5038 (N_5038,N_4482,N_584);
or U5039 (N_5039,N_1272,N_1572);
nor U5040 (N_5040,N_1213,N_323);
or U5041 (N_5041,N_1490,N_1453);
and U5042 (N_5042,N_4473,N_1779);
and U5043 (N_5043,N_4949,N_604);
nor U5044 (N_5044,N_2579,N_659);
nand U5045 (N_5045,N_4719,N_4701);
nand U5046 (N_5046,N_345,N_4832);
or U5047 (N_5047,N_3356,N_4656);
nor U5048 (N_5048,N_4675,N_4599);
and U5049 (N_5049,N_1935,N_4773);
nand U5050 (N_5050,N_788,N_4147);
and U5051 (N_5051,N_315,N_3845);
xnor U5052 (N_5052,N_3276,N_4459);
nand U5053 (N_5053,N_577,N_2205);
nand U5054 (N_5054,N_4799,N_2901);
or U5055 (N_5055,N_1730,N_3014);
and U5056 (N_5056,N_2210,N_3184);
nor U5057 (N_5057,N_1688,N_3828);
nand U5058 (N_5058,N_4284,N_1865);
nand U5059 (N_5059,N_3999,N_470);
nor U5060 (N_5060,N_1384,N_1664);
nand U5061 (N_5061,N_1945,N_4234);
nand U5062 (N_5062,N_4047,N_1963);
xor U5063 (N_5063,N_2409,N_4537);
or U5064 (N_5064,N_2933,N_693);
and U5065 (N_5065,N_4692,N_3640);
and U5066 (N_5066,N_3705,N_4292);
and U5067 (N_5067,N_933,N_3065);
or U5068 (N_5068,N_610,N_2715);
and U5069 (N_5069,N_1208,N_1464);
nor U5070 (N_5070,N_3524,N_1260);
nand U5071 (N_5071,N_4135,N_1310);
and U5072 (N_5072,N_2719,N_2249);
or U5073 (N_5073,N_4689,N_3443);
or U5074 (N_5074,N_2452,N_3847);
or U5075 (N_5075,N_308,N_870);
nand U5076 (N_5076,N_612,N_4854);
xor U5077 (N_5077,N_1449,N_2662);
or U5078 (N_5078,N_3132,N_115);
nand U5079 (N_5079,N_1701,N_1146);
nor U5080 (N_5080,N_1643,N_4485);
or U5081 (N_5081,N_2717,N_4503);
or U5082 (N_5082,N_3967,N_3015);
nand U5083 (N_5083,N_965,N_732);
nor U5084 (N_5084,N_784,N_3961);
or U5085 (N_5085,N_566,N_680);
nand U5086 (N_5086,N_400,N_3632);
nand U5087 (N_5087,N_3700,N_1682);
or U5088 (N_5088,N_472,N_597);
nor U5089 (N_5089,N_3118,N_132);
and U5090 (N_5090,N_1617,N_140);
or U5091 (N_5091,N_1204,N_1436);
and U5092 (N_5092,N_4806,N_3223);
or U5093 (N_5093,N_1512,N_2638);
and U5094 (N_5094,N_3724,N_303);
nand U5095 (N_5095,N_3018,N_2553);
or U5096 (N_5096,N_519,N_4996);
nand U5097 (N_5097,N_1286,N_3788);
or U5098 (N_5098,N_4471,N_1559);
xnor U5099 (N_5099,N_3962,N_2509);
or U5100 (N_5100,N_1965,N_3309);
xor U5101 (N_5101,N_809,N_491);
and U5102 (N_5102,N_856,N_945);
nor U5103 (N_5103,N_1223,N_3075);
and U5104 (N_5104,N_1431,N_2112);
nand U5105 (N_5105,N_4308,N_1913);
xnor U5106 (N_5106,N_217,N_1823);
nand U5107 (N_5107,N_2423,N_2397);
nor U5108 (N_5108,N_4869,N_858);
nand U5109 (N_5109,N_1440,N_1822);
or U5110 (N_5110,N_3557,N_2142);
nand U5111 (N_5111,N_807,N_707);
nand U5112 (N_5112,N_2466,N_4794);
nand U5113 (N_5113,N_1888,N_2345);
and U5114 (N_5114,N_1615,N_1645);
and U5115 (N_5115,N_1777,N_3483);
nand U5116 (N_5116,N_4793,N_4247);
or U5117 (N_5117,N_2119,N_928);
nand U5118 (N_5118,N_1177,N_860);
nand U5119 (N_5119,N_4655,N_935);
nand U5120 (N_5120,N_329,N_2241);
nand U5121 (N_5121,N_2643,N_1616);
or U5122 (N_5122,N_1959,N_1073);
xnor U5123 (N_5123,N_660,N_2214);
nor U5124 (N_5124,N_558,N_1503);
nor U5125 (N_5125,N_1488,N_4067);
or U5126 (N_5126,N_4756,N_3471);
xnor U5127 (N_5127,N_740,N_3500);
and U5128 (N_5128,N_431,N_111);
nand U5129 (N_5129,N_3227,N_1504);
and U5130 (N_5130,N_350,N_999);
nor U5131 (N_5131,N_2239,N_275);
or U5132 (N_5132,N_3761,N_16);
and U5133 (N_5133,N_4850,N_17);
and U5134 (N_5134,N_782,N_1075);
and U5135 (N_5135,N_2012,N_2317);
nor U5136 (N_5136,N_316,N_2093);
and U5137 (N_5137,N_4628,N_2080);
xor U5138 (N_5138,N_3529,N_743);
and U5139 (N_5139,N_2282,N_994);
or U5140 (N_5140,N_2938,N_2301);
xor U5141 (N_5141,N_236,N_3365);
xnor U5142 (N_5142,N_3976,N_3985);
nor U5143 (N_5143,N_4753,N_2368);
nor U5144 (N_5144,N_1187,N_3499);
nor U5145 (N_5145,N_2331,N_3189);
or U5146 (N_5146,N_2690,N_3814);
or U5147 (N_5147,N_1719,N_3839);
xnor U5148 (N_5148,N_3736,N_4297);
or U5149 (N_5149,N_2923,N_3759);
or U5150 (N_5150,N_3032,N_2799);
nand U5151 (N_5151,N_2962,N_538);
and U5152 (N_5152,N_2890,N_1374);
and U5153 (N_5153,N_3507,N_4586);
nand U5154 (N_5154,N_3628,N_3397);
nand U5155 (N_5155,N_949,N_2569);
nor U5156 (N_5156,N_4136,N_4357);
xnor U5157 (N_5157,N_3563,N_4937);
xnor U5158 (N_5158,N_1882,N_3658);
xor U5159 (N_5159,N_2186,N_3644);
or U5160 (N_5160,N_1424,N_2144);
nor U5161 (N_5161,N_2967,N_1291);
or U5162 (N_5162,N_1898,N_434);
and U5163 (N_5163,N_1912,N_1125);
and U5164 (N_5164,N_1622,N_2013);
xor U5165 (N_5165,N_2953,N_849);
nand U5166 (N_5166,N_4477,N_4164);
xnor U5167 (N_5167,N_361,N_4945);
and U5168 (N_5168,N_2976,N_1557);
or U5169 (N_5169,N_1072,N_2160);
xnor U5170 (N_5170,N_4565,N_313);
nor U5171 (N_5171,N_4480,N_388);
nand U5172 (N_5172,N_1793,N_4249);
or U5173 (N_5173,N_4771,N_365);
and U5174 (N_5174,N_2918,N_1373);
nand U5175 (N_5175,N_967,N_3720);
xnor U5176 (N_5176,N_2386,N_1138);
nand U5177 (N_5177,N_3629,N_4368);
xnor U5178 (N_5178,N_4621,N_4940);
xnor U5179 (N_5179,N_4734,N_4143);
xor U5180 (N_5180,N_657,N_29);
xnor U5181 (N_5181,N_2695,N_3401);
nor U5182 (N_5182,N_4082,N_4351);
or U5183 (N_5183,N_2004,N_1709);
nor U5184 (N_5184,N_64,N_2649);
nand U5185 (N_5185,N_4422,N_370);
nand U5186 (N_5186,N_1438,N_3496);
or U5187 (N_5187,N_2064,N_271);
nor U5188 (N_5188,N_1606,N_4658);
nor U5189 (N_5189,N_4727,N_4105);
nor U5190 (N_5190,N_4294,N_263);
or U5191 (N_5191,N_2276,N_917);
nand U5192 (N_5192,N_1751,N_461);
or U5193 (N_5193,N_4810,N_1770);
or U5194 (N_5194,N_4010,N_3140);
and U5195 (N_5195,N_415,N_1519);
xnor U5196 (N_5196,N_4566,N_2861);
and U5197 (N_5197,N_2114,N_2833);
and U5198 (N_5198,N_4748,N_1983);
xnor U5199 (N_5199,N_2610,N_1928);
nor U5200 (N_5200,N_1218,N_2718);
xor U5201 (N_5201,N_4664,N_2231);
nand U5202 (N_5202,N_2990,N_2955);
nand U5203 (N_5203,N_290,N_4497);
or U5204 (N_5204,N_3957,N_4227);
nor U5205 (N_5205,N_2469,N_1571);
or U5206 (N_5206,N_2439,N_3183);
or U5207 (N_5207,N_105,N_3053);
nand U5208 (N_5208,N_4772,N_3);
nor U5209 (N_5209,N_4933,N_4316);
xnor U5210 (N_5210,N_1832,N_1895);
nor U5211 (N_5211,N_4663,N_4114);
xor U5212 (N_5212,N_1122,N_2903);
nand U5213 (N_5213,N_1129,N_71);
nand U5214 (N_5214,N_867,N_4398);
nor U5215 (N_5215,N_4571,N_4747);
and U5216 (N_5216,N_277,N_2107);
or U5217 (N_5217,N_387,N_4581);
nor U5218 (N_5218,N_3158,N_4838);
or U5219 (N_5219,N_1659,N_4768);
or U5220 (N_5220,N_2355,N_3717);
xnor U5221 (N_5221,N_3570,N_2503);
nor U5222 (N_5222,N_1466,N_1459);
nor U5223 (N_5223,N_3256,N_3777);
or U5224 (N_5224,N_3737,N_1479);
or U5225 (N_5225,N_372,N_4601);
nor U5226 (N_5226,N_3406,N_2778);
or U5227 (N_5227,N_4204,N_2607);
nor U5228 (N_5228,N_2473,N_3797);
nand U5229 (N_5229,N_3357,N_663);
nand U5230 (N_5230,N_487,N_1949);
nand U5231 (N_5231,N_866,N_4613);
nand U5232 (N_5232,N_3395,N_3941);
nand U5233 (N_5233,N_3911,N_686);
nand U5234 (N_5234,N_2742,N_3222);
or U5235 (N_5235,N_215,N_4019);
and U5236 (N_5236,N_2959,N_4597);
nand U5237 (N_5237,N_2325,N_4751);
and U5238 (N_5238,N_2372,N_3559);
and U5239 (N_5239,N_328,N_2480);
xor U5240 (N_5240,N_2703,N_4903);
xnor U5241 (N_5241,N_1242,N_1174);
xnor U5242 (N_5242,N_2958,N_4881);
and U5243 (N_5243,N_1710,N_1181);
and U5244 (N_5244,N_1210,N_4671);
or U5245 (N_5245,N_2248,N_2130);
or U5246 (N_5246,N_1604,N_2341);
and U5247 (N_5247,N_2075,N_2382);
xor U5248 (N_5248,N_3448,N_3179);
and U5249 (N_5249,N_3956,N_731);
and U5250 (N_5250,N_2942,N_2853);
nand U5251 (N_5251,N_1860,N_3565);
or U5252 (N_5252,N_1000,N_3601);
and U5253 (N_5253,N_2741,N_606);
and U5254 (N_5254,N_403,N_1406);
nand U5255 (N_5255,N_4836,N_854);
and U5256 (N_5256,N_2804,N_2099);
and U5257 (N_5257,N_3859,N_3177);
nor U5258 (N_5258,N_363,N_4786);
nand U5259 (N_5259,N_369,N_3329);
xnor U5260 (N_5260,N_3332,N_4044);
and U5261 (N_5261,N_4025,N_1350);
nand U5262 (N_5262,N_2582,N_3833);
nand U5263 (N_5263,N_2867,N_3208);
nand U5264 (N_5264,N_458,N_3168);
nor U5265 (N_5265,N_3259,N_2088);
or U5266 (N_5266,N_581,N_2187);
nand U5267 (N_5267,N_3299,N_3279);
and U5268 (N_5268,N_4667,N_3966);
nor U5269 (N_5269,N_2475,N_3339);
xor U5270 (N_5270,N_3454,N_4391);
nand U5271 (N_5271,N_4486,N_2623);
or U5272 (N_5272,N_2247,N_877);
nand U5273 (N_5273,N_926,N_379);
nand U5274 (N_5274,N_3322,N_2336);
and U5275 (N_5275,N_3829,N_1762);
or U5276 (N_5276,N_590,N_3661);
or U5277 (N_5277,N_3417,N_2222);
or U5278 (N_5278,N_1341,N_2000);
nand U5279 (N_5279,N_1325,N_3914);
nand U5280 (N_5280,N_2814,N_125);
nand U5281 (N_5281,N_2612,N_4139);
nor U5282 (N_5282,N_3145,N_4952);
nor U5283 (N_5283,N_4310,N_3897);
nor U5284 (N_5284,N_50,N_1165);
and U5285 (N_5285,N_2864,N_4737);
and U5286 (N_5286,N_547,N_2143);
or U5287 (N_5287,N_87,N_1747);
and U5288 (N_5288,N_1782,N_778);
nand U5289 (N_5289,N_182,N_2783);
nand U5290 (N_5290,N_811,N_1619);
nand U5291 (N_5291,N_2468,N_1514);
or U5292 (N_5292,N_2927,N_395);
or U5293 (N_5293,N_1744,N_2792);
or U5294 (N_5294,N_3115,N_3138);
or U5295 (N_5295,N_2197,N_256);
xnor U5296 (N_5296,N_2514,N_82);
and U5297 (N_5297,N_971,N_4875);
or U5298 (N_5298,N_2482,N_2847);
or U5299 (N_5299,N_4424,N_3019);
or U5300 (N_5300,N_2150,N_3306);
or U5301 (N_5301,N_245,N_1062);
or U5302 (N_5302,N_4347,N_3308);
nand U5303 (N_5303,N_1868,N_3623);
nor U5304 (N_5304,N_4358,N_489);
nor U5305 (N_5305,N_3776,N_2543);
or U5306 (N_5306,N_4785,N_4847);
nand U5307 (N_5307,N_3931,N_99);
and U5308 (N_5308,N_463,N_218);
nor U5309 (N_5309,N_1176,N_61);
and U5310 (N_5310,N_2800,N_3157);
and U5311 (N_5311,N_4997,N_2993);
and U5312 (N_5312,N_1361,N_3773);
nand U5313 (N_5313,N_1870,N_43);
nor U5314 (N_5314,N_102,N_432);
nor U5315 (N_5315,N_1605,N_4140);
and U5316 (N_5316,N_4913,N_4699);
or U5317 (N_5317,N_4987,N_1232);
and U5318 (N_5318,N_3281,N_1052);
and U5319 (N_5319,N_3811,N_638);
xnor U5320 (N_5320,N_1422,N_4556);
nor U5321 (N_5321,N_3770,N_4718);
and U5322 (N_5322,N_4231,N_739);
nor U5323 (N_5323,N_4740,N_1944);
nand U5324 (N_5324,N_2220,N_769);
or U5325 (N_5325,N_4916,N_2201);
nor U5326 (N_5326,N_327,N_4244);
xor U5327 (N_5327,N_1937,N_3134);
nand U5328 (N_5328,N_908,N_542);
nand U5329 (N_5329,N_4723,N_3298);
and U5330 (N_5330,N_2876,N_726);
and U5331 (N_5331,N_3642,N_4609);
nor U5332 (N_5332,N_4371,N_2292);
nor U5333 (N_5333,N_1791,N_268);
and U5334 (N_5334,N_3358,N_1840);
nand U5335 (N_5335,N_453,N_4220);
and U5336 (N_5336,N_647,N_734);
and U5337 (N_5337,N_2369,N_777);
nand U5338 (N_5338,N_2175,N_3836);
nand U5339 (N_5339,N_4962,N_909);
nand U5340 (N_5340,N_2635,N_3293);
nand U5341 (N_5341,N_3462,N_4661);
nor U5342 (N_5342,N_98,N_3671);
or U5343 (N_5343,N_1578,N_3783);
nor U5344 (N_5344,N_1078,N_3525);
nand U5345 (N_5345,N_4919,N_1362);
and U5346 (N_5346,N_2297,N_3230);
nand U5347 (N_5347,N_3943,N_3675);
nor U5348 (N_5348,N_540,N_600);
and U5349 (N_5349,N_2095,N_279);
nand U5350 (N_5350,N_3009,N_3917);
nand U5351 (N_5351,N_494,N_3772);
or U5352 (N_5352,N_1906,N_3561);
or U5353 (N_5353,N_1731,N_2495);
xnor U5354 (N_5354,N_2034,N_116);
and U5355 (N_5355,N_1769,N_2512);
and U5356 (N_5356,N_1432,N_2304);
nand U5357 (N_5357,N_2185,N_2165);
nand U5358 (N_5358,N_2094,N_2191);
or U5359 (N_5359,N_2489,N_3929);
nor U5360 (N_5360,N_1287,N_2318);
or U5361 (N_5361,N_2892,N_3185);
xor U5362 (N_5362,N_4390,N_110);
nor U5363 (N_5363,N_4091,N_3442);
nand U5364 (N_5364,N_741,N_1295);
and U5365 (N_5365,N_187,N_2436);
nand U5366 (N_5366,N_1396,N_3178);
and U5367 (N_5367,N_3674,N_2398);
nand U5368 (N_5368,N_4688,N_1494);
and U5369 (N_5369,N_733,N_1924);
nor U5370 (N_5370,N_4541,N_4319);
nor U5371 (N_5371,N_4846,N_2443);
and U5372 (N_5372,N_1943,N_2278);
and U5373 (N_5373,N_3342,N_4819);
and U5374 (N_5374,N_2878,N_3953);
and U5375 (N_5375,N_4595,N_1461);
or U5376 (N_5376,N_3960,N_4637);
nand U5377 (N_5377,N_7,N_2748);
xor U5378 (N_5378,N_2023,N_4160);
or U5379 (N_5379,N_4040,N_2155);
and U5380 (N_5380,N_512,N_4831);
nor U5381 (N_5381,N_1363,N_3954);
nand U5382 (N_5382,N_3469,N_1971);
nand U5383 (N_5383,N_3522,N_1752);
nand U5384 (N_5384,N_4145,N_417);
nand U5385 (N_5385,N_3219,N_3840);
nand U5386 (N_5386,N_2299,N_4990);
or U5387 (N_5387,N_2057,N_1544);
or U5388 (N_5388,N_1675,N_1127);
xor U5389 (N_5389,N_1936,N_4970);
nand U5390 (N_5390,N_4376,N_3351);
or U5391 (N_5391,N_1856,N_4254);
xnor U5392 (N_5392,N_477,N_1238);
or U5393 (N_5393,N_3531,N_2886);
and U5394 (N_5394,N_1917,N_756);
or U5395 (N_5395,N_4265,N_3434);
nand U5396 (N_5396,N_691,N_1566);
or U5397 (N_5397,N_3686,N_644);
nand U5398 (N_5398,N_4226,N_24);
and U5399 (N_5399,N_2755,N_456);
and U5400 (N_5400,N_685,N_3089);
or U5401 (N_5401,N_4245,N_2445);
nand U5402 (N_5402,N_153,N_3834);
nand U5403 (N_5403,N_4801,N_2073);
or U5404 (N_5404,N_4645,N_3461);
nand U5405 (N_5405,N_1324,N_2496);
nor U5406 (N_5406,N_4205,N_1050);
and U5407 (N_5407,N_3044,N_4968);
nor U5408 (N_5408,N_2828,N_4035);
and U5409 (N_5409,N_1261,N_338);
and U5410 (N_5410,N_1785,N_4063);
or U5411 (N_5411,N_4000,N_958);
and U5412 (N_5412,N_815,N_2928);
nand U5413 (N_5413,N_3647,N_2856);
nand U5414 (N_5414,N_1960,N_1946);
nor U5415 (N_5415,N_3768,N_4223);
or U5416 (N_5416,N_339,N_4153);
and U5417 (N_5417,N_1715,N_1666);
or U5418 (N_5418,N_3051,N_1554);
and U5419 (N_5419,N_3362,N_4752);
nor U5420 (N_5420,N_211,N_2120);
or U5421 (N_5421,N_2193,N_3654);
nor U5422 (N_5422,N_3988,N_3475);
xor U5423 (N_5423,N_3334,N_2361);
nor U5424 (N_5424,N_1357,N_2721);
and U5425 (N_5425,N_3918,N_2611);
xor U5426 (N_5426,N_1783,N_3584);
nor U5427 (N_5427,N_4083,N_2855);
nor U5428 (N_5428,N_3533,N_2428);
nand U5429 (N_5429,N_3937,N_2555);
nor U5430 (N_5430,N_1403,N_3894);
or U5431 (N_5431,N_3187,N_3304);
and U5432 (N_5432,N_2152,N_240);
nand U5433 (N_5433,N_2042,N_2133);
or U5434 (N_5434,N_694,N_2904);
nand U5435 (N_5435,N_3760,N_761);
and U5436 (N_5436,N_1425,N_262);
nand U5437 (N_5437,N_231,N_1650);
xnor U5438 (N_5438,N_4977,N_526);
nand U5439 (N_5439,N_1356,N_2052);
nand U5440 (N_5440,N_4030,N_4829);
nand U5441 (N_5441,N_396,N_2954);
and U5442 (N_5442,N_4602,N_2277);
and U5443 (N_5443,N_562,N_3486);
or U5444 (N_5444,N_92,N_4453);
and U5445 (N_5445,N_3341,N_3538);
nand U5446 (N_5446,N_3196,N_4094);
or U5447 (N_5447,N_2420,N_1728);
or U5448 (N_5448,N_1923,N_3203);
or U5449 (N_5449,N_3385,N_617);
nand U5450 (N_5450,N_1063,N_3239);
nand U5451 (N_5451,N_3478,N_783);
nand U5452 (N_5452,N_2309,N_3867);
nor U5453 (N_5453,N_1095,N_274);
and U5454 (N_5454,N_3904,N_1253);
nand U5455 (N_5455,N_3636,N_1290);
nor U5456 (N_5456,N_1005,N_3495);
nand U5457 (N_5457,N_3938,N_4394);
or U5458 (N_5458,N_853,N_2236);
and U5459 (N_5459,N_4588,N_3915);
and U5460 (N_5460,N_4028,N_1774);
nor U5461 (N_5461,N_1876,N_3896);
nor U5462 (N_5462,N_86,N_4134);
nor U5463 (N_5463,N_3913,N_615);
nor U5464 (N_5464,N_428,N_898);
and U5465 (N_5465,N_2421,N_3925);
and U5466 (N_5466,N_3266,N_1738);
xnor U5467 (N_5467,N_972,N_3311);
or U5468 (N_5468,N_826,N_2785);
nor U5469 (N_5469,N_2787,N_3541);
nand U5470 (N_5470,N_3481,N_3216);
or U5471 (N_5471,N_543,N_2001);
or U5472 (N_5472,N_1764,N_2889);
nor U5473 (N_5473,N_695,N_737);
nand U5474 (N_5474,N_4168,N_890);
and U5475 (N_5475,N_2877,N_4530);
or U5476 (N_5476,N_421,N_2259);
and U5477 (N_5477,N_4267,N_2530);
and U5478 (N_5478,N_4104,N_3922);
xor U5479 (N_5479,N_534,N_931);
nand U5480 (N_5480,N_4582,N_4781);
nand U5481 (N_5481,N_265,N_3399);
or U5482 (N_5482,N_1089,N_3986);
and U5483 (N_5483,N_1700,N_1333);
and U5484 (N_5484,N_3120,N_3662);
and U5485 (N_5485,N_4495,N_307);
nor U5486 (N_5486,N_1609,N_452);
nor U5487 (N_5487,N_4301,N_195);
xor U5488 (N_5488,N_4285,N_3111);
or U5489 (N_5489,N_2636,N_751);
nor U5490 (N_5490,N_1850,N_36);
and U5491 (N_5491,N_42,N_3046);
nor U5492 (N_5492,N_2275,N_3238);
or U5493 (N_5493,N_4434,N_305);
nor U5494 (N_5494,N_3676,N_3864);
or U5495 (N_5495,N_573,N_2279);
and U5496 (N_5496,N_306,N_682);
nor U5497 (N_5497,N_337,N_2104);
nor U5498 (N_5498,N_3635,N_4858);
and U5499 (N_5499,N_517,N_4715);
xor U5500 (N_5500,N_3430,N_2015);
and U5501 (N_5501,N_3368,N_1740);
nor U5502 (N_5502,N_572,N_4200);
nor U5503 (N_5503,N_4941,N_1112);
nand U5504 (N_5504,N_4921,N_4144);
nor U5505 (N_5505,N_1267,N_2298);
nor U5506 (N_5506,N_2658,N_1932);
or U5507 (N_5507,N_4364,N_885);
nor U5508 (N_5508,N_1014,N_1828);
nor U5509 (N_5509,N_2657,N_386);
nand U5510 (N_5510,N_4397,N_79);
and U5511 (N_5511,N_4444,N_3620);
nand U5512 (N_5512,N_40,N_205);
and U5513 (N_5513,N_3591,N_2977);
nand U5514 (N_5514,N_4171,N_3373);
or U5515 (N_5515,N_407,N_4998);
or U5516 (N_5516,N_112,N_1389);
and U5517 (N_5517,N_1395,N_4470);
and U5518 (N_5518,N_1629,N_4431);
or U5519 (N_5519,N_2809,N_4460);
nor U5520 (N_5520,N_3171,N_1343);
xor U5521 (N_5521,N_85,N_1694);
and U5522 (N_5522,N_1720,N_4065);
or U5523 (N_5523,N_4953,N_4629);
or U5524 (N_5524,N_2111,N_203);
nor U5525 (N_5525,N_4580,N_2830);
and U5526 (N_5526,N_1200,N_944);
xor U5527 (N_5527,N_1601,N_2791);
and U5528 (N_5528,N_156,N_390);
or U5529 (N_5529,N_633,N_3819);
nand U5530 (N_5530,N_2086,N_725);
or U5531 (N_5531,N_1550,N_3423);
nand U5532 (N_5532,N_648,N_2486);
or U5533 (N_5533,N_3100,N_2709);
nor U5534 (N_5534,N_76,N_3668);
nor U5535 (N_5535,N_4388,N_3148);
or U5536 (N_5536,N_2603,N_109);
nand U5537 (N_5537,N_2552,N_2138);
xor U5538 (N_5538,N_2507,N_609);
nand U5539 (N_5539,N_2429,N_522);
or U5540 (N_5540,N_155,N_2158);
xnor U5541 (N_5541,N_1886,N_2860);
or U5542 (N_5542,N_701,N_624);
and U5543 (N_5543,N_2314,N_2704);
nand U5544 (N_5544,N_3993,N_636);
nor U5545 (N_5545,N_3518,N_4163);
nand U5546 (N_5546,N_1680,N_1657);
xnor U5547 (N_5547,N_759,N_2441);
or U5548 (N_5548,N_1400,N_1017);
nand U5549 (N_5549,N_1008,N_3473);
and U5550 (N_5550,N_60,N_956);
and U5551 (N_5551,N_2379,N_1511);
nand U5552 (N_5552,N_4167,N_2625);
nand U5553 (N_5553,N_2344,N_869);
or U5554 (N_5554,N_1890,N_2364);
nor U5555 (N_5555,N_1244,N_3427);
nand U5556 (N_5556,N_3589,N_974);
and U5557 (N_5557,N_1185,N_3318);
and U5558 (N_5558,N_1801,N_4053);
and U5559 (N_5559,N_4592,N_2254);
nand U5560 (N_5560,N_3590,N_2671);
nor U5561 (N_5561,N_3240,N_2692);
or U5562 (N_5562,N_3117,N_3835);
nor U5563 (N_5563,N_3031,N_1330);
and U5564 (N_5564,N_1392,N_3103);
nand U5565 (N_5565,N_3684,N_399);
and U5566 (N_5566,N_1158,N_2675);
nand U5567 (N_5567,N_2432,N_4704);
and U5568 (N_5568,N_1849,N_3153);
and U5569 (N_5569,N_4488,N_3210);
and U5570 (N_5570,N_835,N_3599);
nand U5571 (N_5571,N_882,N_3274);
nor U5572 (N_5572,N_4341,N_1029);
nor U5573 (N_5573,N_673,N_3732);
or U5574 (N_5574,N_2682,N_3727);
nand U5575 (N_5575,N_259,N_2537);
nand U5576 (N_5576,N_2679,N_3998);
nand U5577 (N_5577,N_1972,N_744);
nor U5578 (N_5578,N_1240,N_1408);
nand U5579 (N_5579,N_1713,N_3394);
or U5580 (N_5580,N_170,N_4708);
and U5581 (N_5581,N_2266,N_3743);
and U5582 (N_5582,N_1069,N_3984);
and U5583 (N_5583,N_4074,N_1812);
nor U5584 (N_5584,N_1151,N_188);
nand U5585 (N_5585,N_2171,N_2985);
nor U5586 (N_5586,N_1968,N_1182);
nor U5587 (N_5587,N_1331,N_505);
nor U5588 (N_5588,N_995,N_2055);
nor U5589 (N_5589,N_2124,N_424);
nor U5590 (N_5590,N_4508,N_1588);
nor U5591 (N_5591,N_3798,N_3125);
nor U5592 (N_5592,N_3916,N_1626);
nand U5593 (N_5593,N_916,N_2674);
xor U5594 (N_5594,N_222,N_3463);
nor U5595 (N_5595,N_4789,N_4138);
or U5596 (N_5596,N_4430,N_3245);
or U5597 (N_5597,N_814,N_3526);
nor U5598 (N_5598,N_3508,N_3502);
and U5599 (N_5599,N_2881,N_1717);
nand U5600 (N_5600,N_1110,N_4295);
xnor U5601 (N_5601,N_4449,N_3086);
and U5602 (N_5602,N_189,N_4579);
and U5603 (N_5603,N_2914,N_2134);
nand U5604 (N_5604,N_2875,N_4625);
or U5605 (N_5605,N_4236,N_3096);
nand U5606 (N_5606,N_2378,N_634);
and U5607 (N_5607,N_1662,N_2296);
nor U5608 (N_5608,N_31,N_3067);
nand U5609 (N_5609,N_3688,N_210);
and U5610 (N_5610,N_3409,N_4766);
nor U5611 (N_5611,N_4131,N_4132);
nand U5612 (N_5612,N_1435,N_4092);
or U5613 (N_5613,N_4618,N_2713);
nand U5614 (N_5614,N_3716,N_1739);
xnor U5615 (N_5615,N_818,N_2587);
xnor U5616 (N_5616,N_1284,N_2237);
nand U5617 (N_5617,N_4273,N_874);
and U5618 (N_5618,N_1993,N_4323);
nor U5619 (N_5619,N_2026,N_2320);
or U5620 (N_5620,N_2438,N_2225);
nand U5621 (N_5621,N_3673,N_4755);
or U5622 (N_5622,N_1235,N_4476);
and U5623 (N_5623,N_2047,N_1545);
and U5624 (N_5624,N_3805,N_3173);
xnor U5625 (N_5625,N_1136,N_2992);
or U5626 (N_5626,N_1836,N_4077);
nor U5627 (N_5627,N_1241,N_4626);
nand U5628 (N_5628,N_2125,N_2170);
nor U5629 (N_5629,N_4839,N_2180);
and U5630 (N_5630,N_2663,N_4175);
xnor U5631 (N_5631,N_1687,N_1907);
nand U5632 (N_5632,N_1562,N_2040);
xor U5633 (N_5633,N_4352,N_478);
and U5634 (N_5634,N_242,N_4287);
and U5635 (N_5635,N_2032,N_4242);
xor U5636 (N_5636,N_2656,N_3886);
or U5637 (N_5637,N_208,N_2836);
and U5638 (N_5638,N_1214,N_1630);
nor U5639 (N_5639,N_4687,N_1327);
or U5640 (N_5640,N_4126,N_4884);
nor U5641 (N_5641,N_3013,N_3633);
nor U5642 (N_5642,N_1348,N_4991);
or U5643 (N_5643,N_2693,N_3622);
and U5644 (N_5644,N_251,N_1342);
or U5645 (N_5645,N_587,N_2128);
nor U5646 (N_5646,N_2906,N_1402);
or U5647 (N_5647,N_3939,N_4007);
or U5648 (N_5648,N_1203,N_1131);
nor U5649 (N_5649,N_1506,N_1821);
nand U5650 (N_5650,N_3320,N_200);
nand U5651 (N_5651,N_2091,N_2519);
nand U5652 (N_5652,N_4359,N_2872);
and U5653 (N_5653,N_3315,N_2773);
or U5654 (N_5654,N_4606,N_1939);
and U5655 (N_5655,N_199,N_3532);
and U5656 (N_5656,N_1285,N_3034);
nand U5657 (N_5657,N_4524,N_2017);
nor U5658 (N_5658,N_806,N_574);
or U5659 (N_5659,N_4012,N_1390);
nor U5660 (N_5660,N_3355,N_23);
and U5661 (N_5661,N_1930,N_67);
and U5662 (N_5662,N_4189,N_1142);
and U5663 (N_5663,N_2559,N_1359);
nor U5664 (N_5664,N_1743,N_2449);
or U5665 (N_5665,N_2739,N_3830);
or U5666 (N_5666,N_4759,N_493);
or U5667 (N_5667,N_4343,N_3021);
nand U5668 (N_5668,N_296,N_4710);
nor U5669 (N_5669,N_3745,N_1274);
or U5670 (N_5670,N_4446,N_121);
nor U5671 (N_5671,N_4712,N_1021);
nor U5672 (N_5672,N_4148,N_3254);
and U5673 (N_5673,N_4974,N_4534);
or U5674 (N_5674,N_1426,N_4899);
nor U5675 (N_5675,N_3807,N_4796);
and U5676 (N_5676,N_4426,N_2338);
or U5677 (N_5677,N_3907,N_1613);
xor U5678 (N_5678,N_1802,N_1117);
or U5679 (N_5679,N_1358,N_2911);
nand U5680 (N_5680,N_1257,N_619);
nand U5681 (N_5681,N_3560,N_1227);
nand U5682 (N_5682,N_3182,N_2151);
nand U5683 (N_5683,N_536,N_1088);
xor U5684 (N_5684,N_4023,N_2812);
or U5685 (N_5685,N_4467,N_1433);
or U5686 (N_5686,N_4883,N_4761);
and U5687 (N_5687,N_244,N_2148);
or U5688 (N_5688,N_2865,N_4560);
xnor U5689 (N_5689,N_3058,N_4238);
nor U5690 (N_5690,N_4356,N_59);
nor U5691 (N_5691,N_2465,N_2256);
nand U5692 (N_5692,N_2838,N_4963);
xor U5693 (N_5693,N_3088,N_1027);
or U5694 (N_5694,N_4237,N_1834);
nor U5695 (N_5695,N_1215,N_2769);
xnor U5696 (N_5696,N_1678,N_2744);
or U5697 (N_5697,N_1874,N_4169);
nor U5698 (N_5698,N_499,N_3392);
nor U5699 (N_5699,N_4109,N_3695);
and U5700 (N_5700,N_1065,N_3249);
or U5701 (N_5701,N_1987,N_4317);
or U5702 (N_5702,N_3832,N_4406);
nand U5703 (N_5703,N_269,N_3665);
and U5704 (N_5704,N_1827,N_2714);
xor U5705 (N_5705,N_888,N_4277);
xor U5706 (N_5706,N_4142,N_915);
nand U5707 (N_5707,N_2196,N_4325);
and U5708 (N_5708,N_1732,N_2633);
nand U5709 (N_5709,N_2442,N_3679);
nand U5710 (N_5710,N_19,N_3535);
or U5711 (N_5711,N_3350,N_1143);
or U5712 (N_5712,N_3952,N_964);
nor U5713 (N_5713,N_626,N_2252);
nor U5714 (N_5714,N_4835,N_294);
nor U5715 (N_5715,N_2784,N_3964);
or U5716 (N_5716,N_1094,N_1294);
and U5717 (N_5717,N_2194,N_1940);
or U5718 (N_5718,N_3992,N_1651);
and U5719 (N_5719,N_4086,N_2290);
xor U5720 (N_5720,N_4900,N_297);
or U5721 (N_5721,N_539,N_978);
or U5722 (N_5722,N_438,N_2550);
or U5723 (N_5723,N_3011,N_2467);
or U5724 (N_5724,N_4073,N_4049);
and U5725 (N_5725,N_1663,N_1207);
nand U5726 (N_5726,N_2200,N_12);
or U5727 (N_5727,N_1197,N_3813);
nor U5728 (N_5728,N_4218,N_135);
or U5729 (N_5729,N_159,N_2411);
nand U5730 (N_5730,N_49,N_2844);
nor U5731 (N_5731,N_2806,N_2154);
nand U5732 (N_5732,N_1019,N_1788);
nor U5733 (N_5733,N_514,N_755);
xor U5734 (N_5734,N_1201,N_1786);
and U5735 (N_5735,N_10,N_4157);
nand U5736 (N_5736,N_1194,N_3114);
or U5737 (N_5737,N_1863,N_4427);
nor U5738 (N_5738,N_1003,N_4392);
nand U5739 (N_5739,N_697,N_2726);
and U5740 (N_5740,N_4652,N_1170);
nor U5741 (N_5741,N_4213,N_1902);
nor U5742 (N_5742,N_621,N_3224);
nor U5743 (N_5743,N_537,N_3775);
or U5744 (N_5744,N_4496,N_4481);
nand U5745 (N_5745,N_1454,N_4484);
or U5746 (N_5746,N_2401,N_1498);
nand U5747 (N_5747,N_863,N_3137);
or U5748 (N_5748,N_4944,N_2337);
nand U5749 (N_5749,N_4880,N_2781);
or U5750 (N_5750,N_3010,N_1305);
nand U5751 (N_5751,N_4914,N_34);
xor U5752 (N_5752,N_1031,N_3188);
nand U5753 (N_5753,N_4409,N_829);
or U5754 (N_5754,N_3586,N_2324);
xnor U5755 (N_5755,N_3723,N_3817);
xor U5756 (N_5756,N_2746,N_3305);
nand U5757 (N_5757,N_4907,N_905);
nand U5758 (N_5758,N_702,N_3689);
nor U5759 (N_5759,N_2852,N_4059);
and U5760 (N_5760,N_4146,N_2848);
and U5761 (N_5761,N_2768,N_528);
nor U5762 (N_5762,N_3942,N_4985);
and U5763 (N_5763,N_4563,N_3476);
and U5764 (N_5764,N_1845,N_3016);
and U5765 (N_5765,N_918,N_4260);
nand U5766 (N_5766,N_3989,N_414);
nand U5767 (N_5767,N_2448,N_1439);
and U5768 (N_5768,N_3575,N_4078);
or U5769 (N_5769,N_1526,N_4425);
and U5770 (N_5770,N_2329,N_4110);
nand U5771 (N_5771,N_665,N_1159);
nor U5772 (N_5772,N_3124,N_4436);
or U5773 (N_5773,N_729,N_264);
nand U5774 (N_5774,N_2234,N_4917);
nor U5775 (N_5775,N_670,N_1387);
or U5776 (N_5776,N_4975,N_513);
nor U5777 (N_5777,N_3459,N_4217);
and U5778 (N_5778,N_4062,N_688);
or U5779 (N_5779,N_56,N_4248);
or U5780 (N_5780,N_2471,N_4526);
and U5781 (N_5781,N_4936,N_1707);
nand U5782 (N_5782,N_2092,N_649);
nand U5783 (N_5783,N_4454,N_4559);
and U5784 (N_5784,N_4641,N_3159);
nor U5785 (N_5785,N_1579,N_1456);
and U5786 (N_5786,N_1268,N_377);
nand U5787 (N_5787,N_4095,N_4149);
or U5788 (N_5788,N_2966,N_4107);
nor U5789 (N_5789,N_235,N_2770);
and U5790 (N_5790,N_1741,N_469);
xor U5791 (N_5791,N_1262,N_3504);
nor U5792 (N_5792,N_4889,N_4695);
nor U5793 (N_5793,N_557,N_2063);
nand U5794 (N_5794,N_4219,N_3881);
and U5795 (N_5795,N_1852,N_3513);
nand U5796 (N_5796,N_3510,N_3202);
nand U5797 (N_5797,N_1144,N_3959);
or U5798 (N_5798,N_4428,N_2062);
or U5799 (N_5799,N_2528,N_1635);
nor U5800 (N_5800,N_552,N_871);
and U5801 (N_5801,N_1116,N_2039);
nand U5802 (N_5802,N_3619,N_2202);
or U5803 (N_5803,N_37,N_3460);
nand U5804 (N_5804,N_1040,N_1683);
nand U5805 (N_5805,N_2366,N_4726);
and U5806 (N_5806,N_2660,N_3677);
xor U5807 (N_5807,N_4211,N_1150);
nor U5808 (N_5808,N_447,N_2316);
nor U5809 (N_5809,N_4697,N_530);
nand U5810 (N_5810,N_1022,N_405);
or U5811 (N_5811,N_2267,N_2044);
and U5812 (N_5812,N_803,N_2389);
or U5813 (N_5813,N_4060,N_2053);
nor U5814 (N_5814,N_2788,N_4894);
or U5815 (N_5815,N_1481,N_4011);
or U5816 (N_5816,N_823,N_4717);
xor U5817 (N_5817,N_950,N_4958);
or U5818 (N_5818,N_2568,N_3488);
or U5819 (N_5819,N_1508,N_4948);
or U5820 (N_5820,N_2826,N_4066);
nor U5821 (N_5821,N_654,N_364);
nand U5822 (N_5822,N_3888,N_3237);
or U5823 (N_5823,N_2767,N_2357);
and U5824 (N_5824,N_2190,N_4108);
xnor U5825 (N_5825,N_4572,N_1543);
nor U5826 (N_5826,N_4642,N_4291);
and U5827 (N_5827,N_504,N_3165);
nor U5828 (N_5828,N_4261,N_922);
and U5829 (N_5829,N_521,N_2618);
nand U5830 (N_5830,N_1696,N_2295);
nor U5831 (N_5831,N_3698,N_198);
nor U5832 (N_5832,N_3370,N_3936);
nand U5833 (N_5833,N_1698,N_4014);
or U5834 (N_5834,N_2963,N_334);
or U5835 (N_5835,N_810,N_1184);
and U5836 (N_5836,N_4298,N_3327);
or U5837 (N_5837,N_158,N_3754);
or U5838 (N_5838,N_3802,N_3078);
and U5839 (N_5839,N_2762,N_2686);
nor U5840 (N_5840,N_1561,N_332);
nand U5841 (N_5841,N_4500,N_4555);
and U5842 (N_5842,N_2716,N_3147);
nand U5843 (N_5843,N_4311,N_2300);
nand U5844 (N_5844,N_276,N_1458);
nand U5845 (N_5845,N_3301,N_2608);
nand U5846 (N_5846,N_1736,N_389);
nor U5847 (N_5847,N_808,N_4474);
or U5848 (N_5848,N_1894,N_2415);
nand U5849 (N_5849,N_1879,N_3098);
nand U5850 (N_5850,N_3604,N_2102);
nor U5851 (N_5851,N_2334,N_1045);
or U5852 (N_5852,N_1525,N_4593);
nor U5853 (N_5853,N_4728,N_1002);
nor U5854 (N_5854,N_3386,N_2027);
xnor U5855 (N_5855,N_4523,N_3369);
and U5856 (N_5856,N_4151,N_3919);
nor U5857 (N_5857,N_1472,N_655);
or U5858 (N_5858,N_3790,N_4009);
nand U5859 (N_5859,N_1135,N_1862);
or U5860 (N_5860,N_1597,N_3612);
xor U5861 (N_5861,N_2457,N_2727);
xor U5862 (N_5862,N_2418,N_2760);
nor U5863 (N_5863,N_194,N_3542);
nand U5864 (N_5864,N_1753,N_515);
nor U5865 (N_5865,N_416,N_2033);
nor U5866 (N_5866,N_2224,N_1042);
nor U5867 (N_5867,N_479,N_3645);
or U5868 (N_5868,N_2022,N_1805);
xor U5869 (N_5869,N_2352,N_4851);
and U5870 (N_5870,N_3102,N_3848);
nor U5871 (N_5871,N_2020,N_4589);
and U5872 (N_5872,N_3294,N_3806);
and U5873 (N_5873,N_1640,N_137);
xor U5874 (N_5874,N_3588,N_1569);
xnor U5875 (N_5875,N_4643,N_1703);
and U5876 (N_5876,N_343,N_589);
and U5877 (N_5877,N_765,N_2585);
nand U5878 (N_5878,N_2002,N_1180);
and U5879 (N_5879,N_1447,N_4366);
or U5880 (N_5880,N_2008,N_3820);
nand U5881 (N_5881,N_2917,N_130);
or U5882 (N_5882,N_2591,N_321);
nor U5883 (N_5883,N_535,N_3435);
nor U5884 (N_5884,N_700,N_3969);
or U5885 (N_5885,N_4904,N_705);
nand U5886 (N_5886,N_516,N_1884);
and U5887 (N_5887,N_868,N_2994);
or U5888 (N_5888,N_3898,N_4911);
or U5889 (N_5889,N_2213,N_3060);
or U5890 (N_5890,N_3353,N_4950);
nand U5891 (N_5891,N_748,N_3364);
nand U5892 (N_5892,N_1872,N_1480);
nor U5893 (N_5893,N_41,N_3932);
and U5894 (N_5894,N_4868,N_720);
nand U5895 (N_5895,N_1302,N_3949);
xor U5896 (N_5896,N_616,N_3062);
or U5897 (N_5897,N_5,N_1320);
xnor U5898 (N_5898,N_4472,N_2131);
and U5899 (N_5899,N_1243,N_937);
and U5900 (N_5900,N_3978,N_4202);
and U5901 (N_5901,N_2988,N_72);
nor U5902 (N_5902,N_687,N_4033);
and U5903 (N_5903,N_4137,N_689);
or U5904 (N_5904,N_3944,N_2998);
nand U5905 (N_5905,N_2174,N_4567);
and U5906 (N_5906,N_1420,N_2902);
or U5907 (N_5907,N_2268,N_1216);
or U5908 (N_5908,N_2588,N_3176);
xor U5909 (N_5909,N_3678,N_2408);
or U5910 (N_5910,N_2869,N_2182);
or U5911 (N_5911,N_2854,N_3634);
and U5912 (N_5912,N_4978,N_1871);
xnor U5913 (N_5913,N_4315,N_2491);
nand U5914 (N_5914,N_4973,N_1998);
and U5915 (N_5915,N_2394,N_2226);
and U5916 (N_5916,N_78,N_4745);
or U5917 (N_5917,N_1074,N_1591);
nor U5918 (N_5918,N_4349,N_2359);
or U5919 (N_5919,N_3968,N_4152);
xnor U5920 (N_5920,N_3095,N_2723);
and U5921 (N_5921,N_3757,N_3869);
nand U5922 (N_5922,N_3530,N_298);
or U5923 (N_5923,N_997,N_3468);
and U5924 (N_5924,N_2212,N_4300);
nand U5925 (N_5925,N_3260,N_2353);
or U5926 (N_5926,N_3035,N_1266);
nand U5927 (N_5927,N_3516,N_3261);
nand U5928 (N_5928,N_1660,N_1169);
or U5929 (N_5929,N_1502,N_549);
nand U5930 (N_5930,N_2219,N_3438);
nand U5931 (N_5931,N_1076,N_2211);
and U5932 (N_5932,N_4382,N_2272);
xor U5933 (N_5933,N_2669,N_3063);
nand U5934 (N_5934,N_4401,N_4912);
and U5935 (N_5935,N_2168,N_1708);
nor U5936 (N_5936,N_3740,N_1188);
nor U5937 (N_5937,N_4021,N_1217);
or U5938 (N_5938,N_4972,N_4113);
nor U5939 (N_5939,N_501,N_3323);
nor U5940 (N_5940,N_1878,N_1130);
nand U5941 (N_5941,N_2006,N_3755);
xnor U5942 (N_5942,N_2260,N_3275);
and U5943 (N_5943,N_2885,N_2895);
or U5944 (N_5944,N_2545,N_1910);
xnor U5945 (N_5945,N_3110,N_3882);
and U5946 (N_5946,N_289,N_2188);
and U5947 (N_5947,N_3352,N_4943);
or U5948 (N_5948,N_3231,N_2176);
nand U5949 (N_5949,N_3702,N_2808);
or U5950 (N_5950,N_2598,N_1303);
nand U5951 (N_5951,N_3070,N_977);
and U5952 (N_5952,N_4162,N_1478);
or U5953 (N_5953,N_3974,N_2971);
nand U5954 (N_5954,N_4767,N_4387);
nand U5955 (N_5955,N_1624,N_4788);
nor U5956 (N_5956,N_3808,N_2899);
nor U5957 (N_5957,N_1470,N_1301);
nor U5958 (N_5958,N_4054,N_2380);
nand U5959 (N_5959,N_1775,N_258);
nand U5960 (N_5960,N_3004,N_2839);
nor U5961 (N_5961,N_2446,N_2983);
nand U5962 (N_5962,N_2425,N_998);
and U5963 (N_5963,N_3980,N_2815);
nor U5964 (N_5964,N_3402,N_4342);
nor U5965 (N_5965,N_2945,N_3026);
xor U5966 (N_5966,N_4438,N_4507);
or U5967 (N_5967,N_2377,N_2245);
xor U5968 (N_5968,N_1423,N_178);
xor U5969 (N_5969,N_246,N_947);
xnor U5970 (N_5970,N_4122,N_961);
nor U5971 (N_5971,N_3343,N_846);
and U5972 (N_5972,N_3324,N_4221);
nor U5973 (N_5973,N_4551,N_2584);
nor U5974 (N_5974,N_1986,N_2233);
nand U5975 (N_5975,N_3630,N_2016);
nand U5976 (N_5976,N_4087,N_941);
nand U5977 (N_5977,N_4070,N_3174);
nor U5978 (N_5978,N_4770,N_3258);
or U5979 (N_5979,N_2265,N_3733);
xnor U5980 (N_5980,N_3887,N_3921);
xor U5981 (N_5981,N_4389,N_4648);
and U5982 (N_5982,N_4456,N_4557);
nor U5983 (N_5983,N_134,N_954);
and U5984 (N_5984,N_353,N_1228);
nor U5985 (N_5985,N_1444,N_325);
nand U5986 (N_5986,N_13,N_4289);
nor U5987 (N_5987,N_1607,N_2908);
nor U5988 (N_5988,N_1066,N_3080);
and U5989 (N_5989,N_1864,N_3972);
nor U5990 (N_5990,N_2599,N_2109);
or U5991 (N_5991,N_3466,N_1450);
nor U5992 (N_5992,N_292,N_2392);
or U5993 (N_5993,N_4711,N_3729);
nand U5994 (N_5994,N_3842,N_4195);
nor U5995 (N_5995,N_4830,N_3965);
and U5996 (N_5996,N_3398,N_1804);
or U5997 (N_5997,N_3912,N_1803);
nand U5998 (N_5998,N_1881,N_3205);
nand U5999 (N_5999,N_1553,N_4611);
or U6000 (N_6000,N_2422,N_2979);
nand U6001 (N_6001,N_3899,N_1369);
or U6002 (N_6002,N_1360,N_4333);
and U6003 (N_6003,N_1283,N_4681);
nand U6004 (N_6004,N_1556,N_2561);
or U6005 (N_6005,N_1515,N_4407);
and U6006 (N_6006,N_4306,N_2261);
nor U6007 (N_6007,N_3841,N_4657);
nor U6008 (N_6008,N_585,N_1382);
nand U6009 (N_6009,N_3849,N_4779);
nand U6010 (N_6010,N_3491,N_4076);
nor U6011 (N_6011,N_3388,N_1168);
nor U6012 (N_6012,N_3708,N_1018);
nand U6013 (N_6013,N_1632,N_2470);
nand U6014 (N_6014,N_3325,N_2078);
and U6015 (N_6015,N_4228,N_4857);
or U6016 (N_6016,N_2601,N_2540);
nand U6017 (N_6017,N_2360,N_4929);
and U6018 (N_6018,N_822,N_551);
or U6019 (N_6019,N_4532,N_3345);
nor U6020 (N_6020,N_2003,N_4493);
nor U6021 (N_6021,N_4763,N_485);
nor U6022 (N_6022,N_4615,N_441);
and U6023 (N_6023,N_1467,N_1211);
and U6024 (N_6024,N_4672,N_2145);
nor U6025 (N_6025,N_4384,N_3970);
or U6026 (N_6026,N_48,N_83);
and U6027 (N_6027,N_2173,N_3194);
nor U6028 (N_6028,N_798,N_440);
or U6029 (N_6029,N_247,N_4279);
nor U6030 (N_6030,N_439,N_880);
or U6031 (N_6031,N_3786,N_2087);
and U6032 (N_6032,N_3426,N_2943);
and U6033 (N_6033,N_2414,N_2706);
nand U6034 (N_6034,N_1255,N_2696);
and U6035 (N_6035,N_4742,N_4216);
nand U6036 (N_6036,N_3302,N_628);
and U6037 (N_6037,N_3617,N_2286);
or U6038 (N_6038,N_4512,N_4192);
nor U6039 (N_6039,N_2575,N_4612);
or U6040 (N_6040,N_3336,N_924);
nor U6041 (N_6041,N_1288,N_3554);
and U6042 (N_6042,N_1097,N_2461);
or U6043 (N_6043,N_4326,N_3407);
and U6044 (N_6044,N_845,N_2518);
nor U6045 (N_6045,N_4483,N_4372);
nand U6046 (N_6046,N_3545,N_3107);
or U6047 (N_6047,N_4631,N_1372);
nor U6048 (N_6048,N_2681,N_1817);
nand U6049 (N_6049,N_3211,N_4433);
nor U6050 (N_6050,N_2577,N_1920);
nor U6051 (N_6051,N_2284,N_4361);
xnor U6052 (N_6052,N_1225,N_3854);
nand U6053 (N_6053,N_2327,N_1830);
xor U6054 (N_6054,N_2766,N_2321);
nor U6055 (N_6055,N_3319,N_3515);
or U6056 (N_6056,N_1964,N_4305);
and U6057 (N_6057,N_2982,N_3810);
nor U6058 (N_6058,N_3025,N_3411);
and U6059 (N_6059,N_3045,N_3879);
xnor U6060 (N_6060,N_2402,N_413);
nor U6061 (N_6061,N_3479,N_1448);
nor U6062 (N_6062,N_3363,N_1304);
xor U6063 (N_6063,N_561,N_3764);
nand U6064 (N_6064,N_4435,N_2346);
or U6065 (N_6065,N_4544,N_1134);
and U6066 (N_6066,N_864,N_2481);
and U6067 (N_6067,N_4072,N_4405);
or U6068 (N_6068,N_502,N_371);
and U6069 (N_6069,N_1175,N_696);
nor U6070 (N_6070,N_1147,N_1321);
nor U6071 (N_6071,N_3375,N_1838);
nor U6072 (N_6072,N_719,N_988);
and U6073 (N_6073,N_4423,N_4018);
nor U6074 (N_6074,N_2560,N_1064);
nor U6075 (N_6075,N_4257,N_2358);
or U6076 (N_6076,N_3052,N_4573);
nor U6077 (N_6077,N_3493,N_2964);
and U6078 (N_6078,N_1226,N_2932);
and U6079 (N_6079,N_4253,N_1254);
xnor U6080 (N_6080,N_920,N_4015);
nand U6081 (N_6081,N_3082,N_4455);
nor U6082 (N_6082,N_4885,N_4373);
or U6083 (N_6083,N_2477,N_1190);
nand U6084 (N_6084,N_3002,N_3412);
or U6085 (N_6085,N_3105,N_4760);
or U6086 (N_6086,N_152,N_2348);
or U6087 (N_6087,N_887,N_3596);
and U6088 (N_6088,N_4198,N_1518);
nand U6089 (N_6089,N_1534,N_473);
nor U6090 (N_6090,N_1681,N_3742);
or U6091 (N_6091,N_3099,N_745);
and U6092 (N_6092,N_4946,N_1319);
nand U6093 (N_6093,N_2956,N_664);
nor U6094 (N_6094,N_2763,N_839);
or U6095 (N_6095,N_100,N_1493);
nand U6096 (N_6096,N_3690,N_1378);
or U6097 (N_6097,N_1355,N_282);
or U6098 (N_6098,N_1727,N_4971);
or U6099 (N_6099,N_1833,N_1648);
nand U6100 (N_6100,N_901,N_471);
nor U6101 (N_6101,N_2594,N_2051);
or U6102 (N_6102,N_3667,N_1451);
nor U6103 (N_6103,N_66,N_4630);
and U6104 (N_6104,N_2689,N_3543);
nand U6105 (N_6105,N_841,N_1391);
nand U6106 (N_6106,N_2654,N_2332);
nand U6107 (N_6107,N_1492,N_38);
nor U6108 (N_6108,N_2308,N_197);
or U6109 (N_6109,N_3858,N_3868);
or U6110 (N_6110,N_1366,N_4853);
nand U6111 (N_6111,N_1674,N_2511);
nor U6112 (N_6112,N_1589,N_4696);
nand U6113 (N_6113,N_671,N_136);
nand U6114 (N_6114,N_4487,N_139);
nand U6115 (N_6115,N_3655,N_3054);
or U6116 (N_6116,N_4784,N_2628);
xnor U6117 (N_6117,N_2969,N_4038);
and U6118 (N_6118,N_1484,N_1155);
nand U6119 (N_6119,N_1541,N_1404);
nand U6120 (N_6120,N_3263,N_2525);
or U6121 (N_6121,N_2312,N_69);
or U6122 (N_6122,N_2845,N_3374);
xnor U6123 (N_6123,N_3631,N_3416);
nor U6124 (N_6124,N_1798,N_3328);
nor U6125 (N_6125,N_1875,N_2049);
or U6126 (N_6126,N_548,N_2728);
nand U6127 (N_6127,N_1704,N_747);
nand U6128 (N_6128,N_3722,N_1776);
nor U6129 (N_6129,N_3226,N_921);
and U6130 (N_6130,N_2666,N_4375);
or U6131 (N_6131,N_2505,N_2743);
or U6132 (N_6132,N_3436,N_4691);
and U6133 (N_6133,N_2772,N_3404);
nor U6134 (N_6134,N_1340,N_455);
nand U6135 (N_6135,N_4809,N_1375);
nor U6136 (N_6136,N_4504,N_3213);
or U6137 (N_6137,N_2535,N_3523);
and U6138 (N_6138,N_873,N_3821);
or U6139 (N_6139,N_3996,N_3382);
nand U6140 (N_6140,N_90,N_1911);
or U6141 (N_6141,N_983,N_1047);
or U6142 (N_6142,N_4938,N_2968);
nand U6143 (N_6143,N_929,N_4731);
nand U6144 (N_6144,N_221,N_2072);
nor U6145 (N_6145,N_3453,N_4821);
nand U6146 (N_6146,N_4901,N_2322);
nand U6147 (N_6147,N_1985,N_4335);
nor U6148 (N_6148,N_3749,N_4190);
or U6149 (N_6149,N_4898,N_3546);
and U6150 (N_6150,N_2404,N_3769);
and U6151 (N_6151,N_2287,N_2622);
nand U6152 (N_6152,N_3963,N_2595);
nand U6153 (N_6153,N_228,N_844);
and U6154 (N_6154,N_3946,N_3680);
nor U6155 (N_6155,N_253,N_4462);
or U6156 (N_6156,N_3991,N_2604);
nand U6157 (N_6157,N_3703,N_3247);
and U6158 (N_6158,N_3648,N_1547);
xor U6159 (N_6159,N_2756,N_2546);
and U6160 (N_6160,N_2651,N_4490);
xnor U6161 (N_6161,N_2498,N_3997);
nor U6162 (N_6162,N_1132,N_47);
xnor U6163 (N_6163,N_546,N_3652);
xor U6164 (N_6164,N_532,N_3815);
xnor U6165 (N_6165,N_2305,N_3577);
nand U6166 (N_6166,N_3517,N_2729);
or U6167 (N_6167,N_138,N_2288);
nand U6168 (N_6168,N_1096,N_2405);
or U6169 (N_6169,N_4274,N_443);
nor U6170 (N_6170,N_4177,N_1486);
or U6171 (N_6171,N_3656,N_173);
or U6172 (N_6172,N_3951,N_1819);
nand U6173 (N_6173,N_3822,N_4492);
or U6174 (N_6174,N_4749,N_4048);
nor U6175 (N_6175,N_2831,N_4417);
or U6176 (N_6176,N_4525,N_3692);
or U6177 (N_6177,N_3494,N_2532);
nor U6178 (N_6178,N_207,N_2879);
or U6179 (N_6179,N_4776,N_3726);
and U6180 (N_6180,N_1611,N_912);
nor U6181 (N_6181,N_2698,N_4209);
nor U6182 (N_6182,N_1428,N_120);
nor U6183 (N_6183,N_1206,N_942);
and U6184 (N_6184,N_4307,N_3094);
or U6185 (N_6185,N_545,N_1263);
and U6186 (N_6186,N_1154,N_4993);
and U6187 (N_6187,N_3746,N_4324);
xnor U6188 (N_6188,N_295,N_320);
or U6189 (N_6189,N_1711,N_2038);
or U6190 (N_6190,N_1495,N_3550);
and U6191 (N_6191,N_2634,N_1086);
nand U6192 (N_6192,N_3360,N_3212);
nor U6193 (N_6193,N_3354,N_4210);
xor U6194 (N_6194,N_850,N_488);
and U6195 (N_6195,N_1010,N_622);
and U6196 (N_6196,N_233,N_2235);
and U6197 (N_6197,N_1580,N_1036);
or U6198 (N_6198,N_1725,N_1345);
or U6199 (N_6199,N_3241,N_2733);
and U6200 (N_6200,N_4080,N_1054);
and U6201 (N_6201,N_4058,N_3064);
nor U6202 (N_6202,N_322,N_4905);
or U6203 (N_6203,N_2694,N_4743);
or U6204 (N_6204,N_4873,N_118);
or U6205 (N_6205,N_992,N_391);
nor U6206 (N_6206,N_4969,N_2147);
and U6207 (N_6207,N_4813,N_3693);
nor U6208 (N_6208,N_1737,N_2794);
and U6209 (N_6209,N_366,N_2426);
or U6210 (N_6210,N_3977,N_3450);
or U6211 (N_6211,N_749,N_4725);
and U6212 (N_6212,N_4103,N_3666);
nand U6213 (N_6213,N_4790,N_2586);
nor U6214 (N_6214,N_3307,N_4172);
or U6215 (N_6215,N_451,N_2381);
nor U6216 (N_6216,N_4461,N_3851);
nor U6217 (N_6217,N_3221,N_2264);
nor U6218 (N_6218,N_4321,N_2554);
nand U6219 (N_6219,N_1754,N_2583);
nor U6220 (N_6220,N_161,N_4336);
xor U6221 (N_6221,N_2274,N_779);
nand U6222 (N_6222,N_3618,N_3626);
or U6223 (N_6223,N_1056,N_2333);
and U6224 (N_6224,N_3587,N_106);
nor U6225 (N_6225,N_1536,N_1057);
and U6226 (N_6226,N_1625,N_1799);
nor U6227 (N_6227,N_1980,N_2919);
and U6228 (N_6228,N_4233,N_2217);
and U6229 (N_6229,N_1351,N_4533);
and U6230 (N_6230,N_3958,N_1922);
or U6231 (N_6231,N_347,N_3314);
nand U6232 (N_6232,N_1309,N_2342);
nand U6233 (N_6233,N_2427,N_2935);
nand U6234 (N_6234,N_881,N_497);
xor U6235 (N_6235,N_4769,N_1760);
nor U6236 (N_6236,N_1957,N_1258);
nand U6237 (N_6237,N_2759,N_4051);
nand U6238 (N_6238,N_4055,N_302);
and U6239 (N_6239,N_2609,N_2285);
and U6240 (N_6240,N_3410,N_1891);
nor U6241 (N_6241,N_642,N_3048);
or U6242 (N_6242,N_3767,N_3225);
nor U6243 (N_6243,N_3204,N_4259);
nor U6244 (N_6244,N_529,N_1892);
nor U6245 (N_6245,N_2871,N_2311);
or U6246 (N_6246,N_556,N_2667);
nand U6247 (N_6247,N_4225,N_3119);
nand U6248 (N_6248,N_3800,N_876);
and U6249 (N_6249,N_1496,N_2557);
or U6250 (N_6250,N_57,N_1976);
nand U6251 (N_6251,N_851,N_3292);
xnor U6252 (N_6252,N_4554,N_2229);
xor U6253 (N_6253,N_3971,N_1442);
nand U6254 (N_6254,N_1256,N_2720);
nand U6255 (N_6255,N_2025,N_4680);
and U6256 (N_6256,N_3389,N_3762);
nand U6257 (N_6257,N_164,N_2617);
nand U6258 (N_6258,N_4955,N_2243);
xor U6259 (N_6259,N_3027,N_1489);
nand U6260 (N_6260,N_1593,N_260);
and U6261 (N_6261,N_1336,N_563);
nand U6262 (N_6262,N_3624,N_4345);
or U6263 (N_6263,N_3544,N_127);
or U6264 (N_6264,N_821,N_1264);
and U6265 (N_6265,N_3778,N_1316);
nand U6266 (N_6266,N_1421,N_430);
or U6267 (N_6267,N_2701,N_160);
nor U6268 (N_6268,N_3683,N_1531);
nor U6269 (N_6269,N_3852,N_3474);
nor U6270 (N_6270,N_4045,N_460);
nand U6271 (N_6271,N_2645,N_3396);
and U6272 (N_6272,N_641,N_1956);
nand U6273 (N_6273,N_1,N_4489);
nor U6274 (N_6274,N_1491,N_3751);
nand U6275 (N_6275,N_4700,N_2931);
nand U6276 (N_6276,N_2891,N_2508);
nand U6277 (N_6277,N_1524,N_2605);
nor U6278 (N_6278,N_1975,N_4529);
nor U6279 (N_6279,N_3994,N_959);
xnor U6280 (N_6280,N_2046,N_927);
or U6281 (N_6281,N_2843,N_678);
xor U6282 (N_6282,N_1610,N_1120);
nand U6283 (N_6283,N_3812,N_401);
nor U6284 (N_6284,N_3758,N_1672);
or U6285 (N_6285,N_3383,N_3371);
or U6286 (N_6286,N_2572,N_3569);
nor U6287 (N_6287,N_715,N_1237);
and U6288 (N_6288,N_2765,N_3853);
and U6289 (N_6289,N_1513,N_3763);
or U6290 (N_6290,N_4340,N_1035);
nor U6291 (N_6291,N_2097,N_4827);
nor U6292 (N_6292,N_1903,N_1252);
nor U6293 (N_6293,N_4334,N_1191);
nand U6294 (N_6294,N_4535,N_4120);
or U6295 (N_6295,N_3017,N_4256);
nand U6296 (N_6296,N_3826,N_3799);
and U6297 (N_6297,N_3598,N_4046);
xor U6298 (N_6298,N_248,N_1462);
nand U6299 (N_6299,N_2117,N_1538);
and U6300 (N_6300,N_4130,N_1800);
nor U6301 (N_6301,N_4016,N_4882);
nand U6302 (N_6302,N_4578,N_1904);
xor U6303 (N_6303,N_2835,N_790);
nand U6304 (N_6304,N_4594,N_1051);
nand U6305 (N_6305,N_1573,N_4797);
nand U6306 (N_6306,N_4005,N_4624);
nand U6307 (N_6307,N_4002,N_2208);
nor U6308 (N_6308,N_1551,N_14);
or U6309 (N_6309,N_1401,N_1289);
nor U6310 (N_6310,N_3246,N_4878);
or U6311 (N_6311,N_1621,N_168);
or U6312 (N_6312,N_4540,N_1352);
nand U6313 (N_6313,N_4251,N_794);
nor U6314 (N_6314,N_4552,N_1766);
and U6315 (N_6315,N_490,N_4339);
nand U6316 (N_6316,N_4951,N_101);
nor U6317 (N_6317,N_299,N_2374);
and U6318 (N_6318,N_3195,N_1835);
nor U6319 (N_6319,N_1140,N_4735);
or U6320 (N_6320,N_2837,N_4362);
and U6321 (N_6321,N_4886,N_2700);
xnor U6322 (N_6322,N_3861,N_261);
or U6323 (N_6323,N_310,N_4240);
nand U6324 (N_6324,N_4906,N_427);
nand U6325 (N_6325,N_495,N_2775);
and U6326 (N_6326,N_4516,N_4367);
or U6327 (N_6327,N_4668,N_3701);
or U6328 (N_6328,N_4024,N_1758);
or U6329 (N_6329,N_374,N_923);
and U6330 (N_6330,N_4320,N_2897);
nand U6331 (N_6331,N_3169,N_1473);
nand U6332 (N_6332,N_979,N_2506);
nand U6333 (N_6333,N_4288,N_1669);
and U6334 (N_6334,N_3312,N_3338);
nor U6335 (N_6335,N_742,N_4976);
and U6336 (N_6336,N_4498,N_704);
and U6337 (N_6337,N_2246,N_141);
nand U6338 (N_6338,N_2747,N_3514);
nand U6339 (N_6339,N_3785,N_1332);
nor U6340 (N_6340,N_4746,N_3458);
and U6341 (N_6341,N_1646,N_2823);
and U6342 (N_6342,N_3844,N_3093);
nand U6343 (N_6343,N_4934,N_1925);
or U6344 (N_6344,N_3753,N_4312);
or U6345 (N_6345,N_278,N_2734);
and U6346 (N_6346,N_2548,N_1156);
and U6347 (N_6347,N_4623,N_2129);
or U6348 (N_6348,N_3033,N_418);
and U6349 (N_6349,N_1516,N_2850);
and U6350 (N_6350,N_1585,N_2670);
or U6351 (N_6351,N_4337,N_4673);
or U6352 (N_6352,N_3432,N_1667);
nor U6353 (N_6353,N_4,N_4923);
nand U6354 (N_6354,N_576,N_1236);
or U6355 (N_6355,N_780,N_3581);
and U6356 (N_6356,N_3267,N_3164);
or U6357 (N_6357,N_2722,N_3186);
xor U6358 (N_6358,N_2567,N_4042);
nand U6359 (N_6359,N_468,N_2326);
and U6360 (N_6360,N_3663,N_919);
nand U6361 (N_6361,N_2456,N_4272);
nand U6362 (N_6362,N_511,N_3347);
nor U6363 (N_6363,N_1546,N_2596);
nor U6364 (N_6364,N_2944,N_4194);
nor U6365 (N_6365,N_627,N_2796);
and U6366 (N_6366,N_4187,N_3487);
and U6367 (N_6367,N_2406,N_3843);
nand U6368 (N_6368,N_2981,N_30);
nand U6369 (N_6369,N_1108,N_2492);
and U6370 (N_6370,N_836,N_4266);
nand U6371 (N_6371,N_2678,N_4617);
and U6372 (N_6372,N_948,N_1280);
and U6373 (N_6373,N_131,N_1501);
or U6374 (N_6374,N_4396,N_766);
nand U6375 (N_6375,N_3116,N_3505);
or U6376 (N_6376,N_148,N_1552);
nor U6377 (N_6377,N_957,N_1246);
or U6378 (N_6378,N_3139,N_594);
nand U6379 (N_6379,N_2253,N_980);
and U6380 (N_6380,N_397,N_1276);
or U6381 (N_6381,N_2672,N_3467);
or U6382 (N_6382,N_2070,N_1399);
nand U6383 (N_6383,N_1220,N_3490);
xnor U6384 (N_6384,N_3900,N_483);
or U6385 (N_6385,N_433,N_3779);
or U6386 (N_6386,N_4206,N_4199);
nor U6387 (N_6387,N_1831,N_2066);
nor U6388 (N_6388,N_3734,N_2789);
or U6389 (N_6389,N_3022,N_3232);
or U6390 (N_6390,N_481,N_450);
nand U6391 (N_6391,N_4848,N_830);
nand U6392 (N_6392,N_4402,N_4677);
nand U6393 (N_6393,N_893,N_1364);
nor U6394 (N_6394,N_46,N_2857);
or U6395 (N_6395,N_1482,N_4591);
nor U6396 (N_6396,N_1994,N_4604);
or U6397 (N_6397,N_3728,N_2642);
and U6398 (N_6398,N_4278,N_1292);
nor U6399 (N_6399,N_4506,N_564);
and U6400 (N_6400,N_4020,N_800);
nor U6401 (N_6401,N_1162,N_1025);
and U6402 (N_6402,N_1468,N_4574);
xnor U6403 (N_6403,N_1349,N_4027);
and U6404 (N_6404,N_77,N_1979);
and U6405 (N_6405,N_3568,N_3049);
or U6406 (N_6406,N_1734,N_1577);
xor U6407 (N_6407,N_793,N_955);
or U6408 (N_6408,N_1306,N_3878);
nor U6409 (N_6409,N_1966,N_1825);
nor U6410 (N_6410,N_3973,N_293);
or U6411 (N_6411,N_1749,N_2258);
nor U6412 (N_6412,N_2597,N_571);
nor U6413 (N_6413,N_3170,N_18);
and U6414 (N_6414,N_2793,N_2786);
nand U6415 (N_6415,N_4984,N_4056);
or U6416 (N_6416,N_3431,N_960);
nand U6417 (N_6417,N_1639,N_1767);
xnor U6418 (N_6418,N_1296,N_3036);
nand U6419 (N_6419,N_2149,N_583);
nor U6420 (N_6420,N_1858,N_3578);
nand U6421 (N_6421,N_3419,N_1581);
or U6422 (N_6422,N_1487,N_3084);
xor U6423 (N_6423,N_4281,N_3739);
nor U6424 (N_6424,N_3511,N_3030);
or U6425 (N_6425,N_4178,N_165);
xnor U6426 (N_6426,N_1847,N_3128);
nand U6427 (N_6427,N_789,N_4380);
nor U6428 (N_6428,N_1141,N_2653);
nor U6429 (N_6429,N_2403,N_2925);
nand U6430 (N_6430,N_4820,N_4378);
nand U6431 (N_6431,N_1763,N_3669);
nand U6432 (N_6432,N_2840,N_1883);
xnor U6433 (N_6433,N_1527,N_3707);
and U6434 (N_6434,N_2105,N_1603);
and U6435 (N_6435,N_1308,N_2619);
or U6436 (N_6436,N_1789,N_385);
and U6437 (N_6437,N_4705,N_2);
xor U6438 (N_6438,N_3081,N_2347);
nor U6439 (N_6439,N_484,N_2754);
nor U6440 (N_6440,N_4468,N_3122);
nor U6441 (N_6441,N_925,N_3979);
xnor U6442 (N_6442,N_367,N_639);
and U6443 (N_6443,N_1735,N_4774);
xnor U6444 (N_6444,N_1013,N_1270);
nand U6445 (N_6445,N_2440,N_1111);
nand U6446 (N_6446,N_1149,N_2947);
and U6447 (N_6447,N_184,N_1093);
nand U6448 (N_6448,N_503,N_4241);
nor U6449 (N_6449,N_1814,N_4686);
nor U6450 (N_6450,N_1397,N_2613);
xor U6451 (N_6451,N_1443,N_4659);
nor U6452 (N_6452,N_1307,N_2227);
and U6453 (N_6453,N_462,N_4208);
and U6454 (N_6454,N_4098,N_987);
and U6455 (N_6455,N_4662,N_1771);
or U6456 (N_6456,N_4440,N_304);
or U6457 (N_6457,N_2232,N_4893);
or U6458 (N_6458,N_2637,N_1385);
or U6459 (N_6459,N_2551,N_2707);
nor U6460 (N_6460,N_2819,N_3020);
nor U6461 (N_6461,N_352,N_601);
nor U6462 (N_6462,N_2323,N_3860);
nor U6463 (N_6463,N_1344,N_3824);
nor U6464 (N_6464,N_1001,N_1746);
or U6465 (N_6465,N_752,N_4910);
nand U6466 (N_6466,N_2164,N_1952);
and U6467 (N_6467,N_2821,N_754);
nor U6468 (N_6468,N_4992,N_4410);
nor U6469 (N_6469,N_288,N_3804);
and U6470 (N_6470,N_4112,N_2712);
nor U6471 (N_6471,N_4694,N_4031);
or U6472 (N_6472,N_1381,N_1087);
and U6473 (N_6473,N_2383,N_4787);
and U6474 (N_6474,N_1641,N_103);
or U6475 (N_6475,N_1560,N_3940);
and U6476 (N_6476,N_969,N_993);
or U6477 (N_6477,N_4647,N_2132);
and U6478 (N_6478,N_2303,N_3113);
or U6479 (N_6479,N_2883,N_3381);
nand U6480 (N_6480,N_951,N_2526);
nand U6481 (N_6481,N_4843,N_1465);
and U6482 (N_6482,N_1510,N_2021);
nor U6483 (N_6483,N_1796,N_2870);
nor U6484 (N_6484,N_2863,N_4676);
nand U6485 (N_6485,N_45,N_4161);
nor U6486 (N_6486,N_2230,N_393);
xor U6487 (N_6487,N_2393,N_861);
and U6488 (N_6488,N_3747,N_2513);
nor U6489 (N_6489,N_114,N_1528);
nand U6490 (N_6490,N_862,N_3485);
or U6491 (N_6491,N_768,N_4924);
nor U6492 (N_6492,N_4520,N_2413);
or U6493 (N_6493,N_1990,N_2089);
or U6494 (N_6494,N_775,N_796);
xnor U6495 (N_6495,N_602,N_1806);
or U6496 (N_6496,N_669,N_1889);
and U6497 (N_6497,N_3349,N_3265);
nand U6498 (N_6498,N_1020,N_4863);
or U6499 (N_6499,N_1673,N_4093);
nor U6500 (N_6500,N_333,N_465);
or U6501 (N_6501,N_341,N_454);
nor U6502 (N_6502,N_3271,N_3945);
or U6503 (N_6503,N_774,N_476);
and U6504 (N_6504,N_721,N_435);
nor U6505 (N_6505,N_2139,N_4639);
or U6506 (N_6506,N_4720,N_1417);
or U6507 (N_6507,N_1469,N_3930);
nor U6508 (N_6508,N_2801,N_1269);
nand U6509 (N_6509,N_2564,N_1602);
nand U6510 (N_6510,N_4116,N_2973);
or U6511 (N_6511,N_2520,N_2779);
or U6512 (N_6512,N_202,N_2035);
or U6513 (N_6513,N_2705,N_1171);
nand U6514 (N_6514,N_4791,N_3252);
and U6515 (N_6515,N_2751,N_1033);
or U6516 (N_6516,N_2435,N_3625);
and U6517 (N_6517,N_4457,N_4965);
and U6518 (N_6518,N_1418,N_3101);
nand U6519 (N_6519,N_2310,N_525);
or U6520 (N_6520,N_3066,N_4798);
nand U6521 (N_6521,N_3519,N_1583);
nand U6522 (N_6522,N_3330,N_3950);
nand U6523 (N_6523,N_718,N_1988);
nand U6524 (N_6524,N_730,N_1463);
nand U6525 (N_6525,N_2351,N_227);
nand U6526 (N_6526,N_544,N_3079);
nor U6527 (N_6527,N_3862,N_1043);
nand U6528 (N_6528,N_4239,N_3659);
nor U6529 (N_6529,N_4874,N_257);
nand U6530 (N_6530,N_2533,N_2343);
or U6531 (N_6531,N_3536,N_1068);
or U6532 (N_6532,N_1161,N_4370);
nand U6533 (N_6533,N_4864,N_3131);
xnor U6534 (N_6534,N_1962,N_2541);
and U6535 (N_6535,N_2464,N_3012);
nand U6536 (N_6536,N_201,N_3895);
or U6537 (N_6537,N_4679,N_4196);
and U6538 (N_6538,N_3947,N_4188);
or U6539 (N_6539,N_2896,N_1586);
or U6540 (N_6540,N_3047,N_4569);
nor U6541 (N_6541,N_2817,N_3870);
xnor U6542 (N_6542,N_1984,N_4915);
nand U6543 (N_6543,N_1452,N_3130);
nand U6544 (N_6544,N_52,N_3340);
nor U6545 (N_6545,N_3983,N_4721);
nand U6546 (N_6546,N_4583,N_4994);
or U6547 (N_6547,N_2184,N_4119);
nor U6548 (N_6548,N_1705,N_4429);
nand U6549 (N_6549,N_3333,N_1032);
or U6550 (N_6550,N_232,N_1665);
nor U6551 (N_6551,N_4587,N_2373);
nor U6552 (N_6552,N_255,N_575);
xor U6553 (N_6553,N_963,N_1961);
and U6554 (N_6554,N_662,N_1311);
xnor U6555 (N_6555,N_20,N_911);
nor U6556 (N_6556,N_2242,N_1745);
nand U6557 (N_6557,N_154,N_4125);
nand U6558 (N_6558,N_3437,N_2121);
and U6559 (N_6559,N_3242,N_1219);
nand U6560 (N_6560,N_3903,N_3981);
or U6561 (N_6561,N_2592,N_3422);
and U6562 (N_6562,N_3449,N_4724);
or U6563 (N_6563,N_340,N_1221);
xor U6564 (N_6564,N_4961,N_2500);
and U6565 (N_6565,N_2740,N_2753);
nor U6566 (N_6566,N_4494,N_1568);
nand U6567 (N_6567,N_183,N_3452);
or U6568 (N_6568,N_2476,N_3583);
nor U6569 (N_6569,N_3883,N_2157);
or U6570 (N_6570,N_1934,N_709);
and U6571 (N_6571,N_1259,N_4732);
or U6572 (N_6572,N_4369,N_1339);
nor U6573 (N_6573,N_2178,N_4895);
nand U6574 (N_6574,N_859,N_4713);
or U6575 (N_6575,N_4255,N_1164);
or U6576 (N_6576,N_3087,N_448);
or U6577 (N_6577,N_4849,N_4897);
or U6578 (N_6578,N_3909,N_3549);
or U6579 (N_6579,N_346,N_3376);
and U6580 (N_6580,N_53,N_667);
and U6581 (N_6581,N_832,N_3553);
xor U6582 (N_6582,N_4464,N_3646);
and U6583 (N_6583,N_4814,N_4318);
or U6584 (N_6584,N_1537,N_1202);
nor U6585 (N_6585,N_1716,N_1049);
nand U6586 (N_6586,N_4729,N_1231);
or U6587 (N_6587,N_1030,N_1160);
nand U6588 (N_6588,N_3697,N_943);
or U6589 (N_6589,N_632,N_1193);
or U6590 (N_6590,N_3926,N_3253);
nor U6591 (N_6591,N_422,N_2576);
nand U6592 (N_6592,N_3547,N_1153);
nand U6593 (N_6593,N_219,N_3792);
and U6594 (N_6594,N_254,N_2183);
or U6595 (N_6595,N_2437,N_4709);
or U6596 (N_6596,N_4224,N_4590);
nand U6597 (N_6597,N_757,N_2058);
nand U6598 (N_6598,N_349,N_1380);
nand U6599 (N_6599,N_4432,N_1277);
nand U6600 (N_6600,N_3891,N_1756);
nor U6601 (N_6601,N_2504,N_4331);
or U6602 (N_6602,N_1567,N_578);
or U6603 (N_6603,N_643,N_2558);
or U6604 (N_6604,N_143,N_239);
and U6605 (N_6605,N_4090,N_2458);
and U6606 (N_6606,N_3447,N_4328);
or U6607 (N_6607,N_1346,N_2921);
and U6608 (N_6608,N_249,N_910);
xor U6609 (N_6609,N_2650,N_2459);
and U6610 (N_6610,N_117,N_4803);
xnor U6611 (N_6611,N_1899,N_1592);
or U6612 (N_6612,N_2758,N_252);
or U6613 (N_6613,N_1455,N_3691);
or U6614 (N_6614,N_4207,N_735);
and U6615 (N_6615,N_3789,N_3771);
xnor U6616 (N_6616,N_4502,N_1250);
nand U6617 (N_6617,N_4262,N_1016);
nor U6618 (N_6618,N_1582,N_1298);
and U6619 (N_6619,N_3607,N_1841);
xor U6620 (N_6620,N_3766,N_4057);
or U6621 (N_6621,N_1102,N_3464);
nor U6622 (N_6622,N_2207,N_4386);
nor U6623 (N_6623,N_2146,N_209);
nor U6624 (N_6624,N_375,N_410);
and U6625 (N_6625,N_2106,N_11);
nor U6626 (N_6626,N_185,N_2195);
xnor U6627 (N_6627,N_4942,N_2661);
or U6628 (N_6628,N_2289,N_760);
nor U6629 (N_6629,N_1163,N_620);
and U6630 (N_6630,N_613,N_3796);
and U6631 (N_6631,N_3711,N_2810);
or U6632 (N_6632,N_28,N_3660);
nor U6633 (N_6633,N_690,N_3167);
nor U6634 (N_6634,N_2090,N_2024);
and U6635 (N_6635,N_4665,N_4079);
or U6636 (N_6636,N_330,N_2019);
nand U6637 (N_6637,N_1419,N_272);
and U6638 (N_6638,N_1810,N_4765);
nand U6639 (N_6639,N_1690,N_190);
nor U6640 (N_6640,N_1460,N_4908);
nand U6641 (N_6641,N_1921,N_3765);
xor U6642 (N_6642,N_4463,N_4778);
nand U6643 (N_6643,N_1477,N_2313);
or U6644 (N_6644,N_1866,N_1861);
and U6645 (N_6645,N_149,N_4890);
nand U6646 (N_6646,N_2499,N_2221);
or U6647 (N_6647,N_716,N_4003);
nand U6648 (N_6648,N_2076,N_2307);
nor U6649 (N_6649,N_4879,N_2687);
nand U6650 (N_6650,N_1485,N_1598);
nor U6651 (N_6651,N_4860,N_91);
or U6652 (N_6652,N_2255,N_398);
and U6653 (N_6653,N_799,N_3875);
and U6654 (N_6654,N_1954,N_2135);
nand U6655 (N_6655,N_3838,N_1587);
nor U6656 (N_6656,N_1249,N_2822);
nand U6657 (N_6657,N_1015,N_420);
and U6658 (N_6658,N_2387,N_991);
nor U6659 (N_6659,N_3393,N_4185);
nand U6660 (N_6660,N_2987,N_1313);
or U6661 (N_6661,N_4986,N_4598);
or U6662 (N_6662,N_3877,N_1178);
or U6663 (N_6663,N_1654,N_4872);
and U6664 (N_6664,N_611,N_3023);
and U6665 (N_6665,N_1061,N_3585);
nand U6666 (N_6666,N_4379,N_1999);
nor U6667 (N_6667,N_2218,N_2451);
and U6668 (N_6668,N_4129,N_2984);
xor U6669 (N_6669,N_4603,N_3880);
nor U6670 (N_6670,N_1273,N_3156);
nand U6671 (N_6671,N_3273,N_2915);
nor U6672 (N_6672,N_1109,N_2216);
or U6673 (N_6673,N_630,N_2455);
nor U6674 (N_6674,N_1718,N_123);
nor U6675 (N_6675,N_4935,N_1652);
and U6676 (N_6676,N_2367,N_1157);
xnor U6677 (N_6677,N_2396,N_1915);
nor U6678 (N_6678,N_3539,N_1041);
xor U6679 (N_6679,N_646,N_73);
and U6680 (N_6680,N_357,N_3890);
nor U6681 (N_6681,N_4174,N_2159);
nand U6682 (N_6682,N_2538,N_1761);
and U6683 (N_6683,N_2937,N_2068);
or U6684 (N_6684,N_2209,N_3893);
or U6685 (N_6685,N_2757,N_2067);
nor U6686 (N_6686,N_2989,N_4246);
or U6687 (N_6687,N_2490,N_4399);
and U6688 (N_6688,N_508,N_230);
nor U6689 (N_6689,N_938,N_1192);
nor U6690 (N_6690,N_4979,N_444);
nand U6691 (N_6691,N_852,N_4855);
or U6692 (N_6692,N_3297,N_2474);
and U6693 (N_6693,N_3520,N_1430);
and U6694 (N_6694,N_4154,N_4181);
and U6695 (N_6695,N_2257,N_2061);
nand U6696 (N_6696,N_4865,N_1787);
nor U6697 (N_6697,N_984,N_3512);
and U6698 (N_6698,N_2644,N_1067);
or U6699 (N_6699,N_4264,N_3028);
nor U6700 (N_6700,N_2350,N_677);
nand U6701 (N_6701,N_1507,N_446);
and U6702 (N_6702,N_2894,N_2790);
xor U6703 (N_6703,N_2898,N_3162);
nand U6704 (N_6704,N_3206,N_4632);
or U6705 (N_6705,N_39,N_464);
xor U6706 (N_6706,N_1724,N_1973);
xor U6707 (N_6707,N_1445,N_1107);
and U6708 (N_6708,N_354,N_2761);
and U6709 (N_6709,N_4706,N_2858);
nor U6710 (N_6710,N_204,N_2251);
nor U6711 (N_6711,N_907,N_4995);
nor U6712 (N_6712,N_4584,N_4669);
and U6713 (N_6713,N_1532,N_2007);
or U6714 (N_6714,N_3069,N_3657);
nor U6715 (N_6715,N_1323,N_1691);
nand U6716 (N_6716,N_1558,N_3855);
nor U6717 (N_6717,N_3975,N_95);
or U6718 (N_6718,N_763,N_2433);
and U6719 (N_6719,N_2009,N_1596);
or U6720 (N_6720,N_1570,N_857);
or U6721 (N_6721,N_753,N_580);
or U6722 (N_6722,N_1271,N_2029);
nand U6723 (N_6723,N_3446,N_952);
or U6724 (N_6724,N_4939,N_4441);
and U6725 (N_6725,N_524,N_2631);
xor U6726 (N_6726,N_1411,N_2664);
and U6727 (N_6727,N_3567,N_3857);
nand U6728 (N_6728,N_4805,N_359);
or U6729 (N_6729,N_1642,N_1300);
nor U6730 (N_6730,N_3077,N_147);
and U6731 (N_6731,N_3425,N_3142);
and U6732 (N_6732,N_2485,N_4651);
and U6733 (N_6733,N_650,N_2711);
and U6734 (N_6734,N_3316,N_2606);
nand U6735 (N_6735,N_4543,N_2807);
and U6736 (N_6736,N_608,N_3250);
nand U6737 (N_6737,N_595,N_3097);
and U6738 (N_6738,N_97,N_1842);
or U6739 (N_6739,N_1655,N_212);
or U6740 (N_6740,N_1908,N_4649);
nand U6741 (N_6741,N_2668,N_656);
xor U6742 (N_6742,N_55,N_3160);
xor U6743 (N_6743,N_3326,N_1813);
nand U6744 (N_6744,N_1317,N_213);
or U6745 (N_6745,N_1755,N_27);
or U6746 (N_6746,N_4562,N_2965);
or U6747 (N_6747,N_2750,N_2665);
nor U6748 (N_6748,N_51,N_3287);
nor U6749 (N_6749,N_2244,N_1873);
xor U6750 (N_6750,N_847,N_266);
nor U6751 (N_6751,N_1661,N_3884);
nor U6752 (N_6752,N_1026,N_225);
or U6753 (N_6753,N_582,N_1409);
or U6754 (N_6754,N_4439,N_1148);
nor U6755 (N_6755,N_736,N_3548);
xnor U6756 (N_6756,N_4106,N_708);
or U6757 (N_6757,N_1471,N_1887);
nand U6758 (N_6758,N_358,N_4270);
nand U6759 (N_6759,N_4258,N_402);
or U6760 (N_6760,N_4550,N_2215);
nand U6761 (N_6761,N_2407,N_2122);
nand U6762 (N_6762,N_80,N_2126);
and U6763 (N_6763,N_392,N_2868);
nand U6764 (N_6764,N_2578,N_4156);
or U6765 (N_6765,N_4707,N_404);
and U6766 (N_6766,N_129,N_2494);
and U6767 (N_6767,N_3042,N_4833);
or U6768 (N_6768,N_2416,N_2527);
or U6769 (N_6769,N_4111,N_2054);
or U6770 (N_6770,N_2074,N_4575);
nor U6771 (N_6771,N_449,N_4415);
nand U6772 (N_6772,N_335,N_4017);
nand U6773 (N_6773,N_1314,N_2802);
nor U6774 (N_6774,N_3650,N_4703);
or U6775 (N_6775,N_914,N_2547);
or U6776 (N_6776,N_1037,N_2580);
nor U6777 (N_6777,N_3509,N_906);
and U6778 (N_6778,N_4989,N_3482);
nor U6779 (N_6779,N_2640,N_1854);
nand U6780 (N_6780,N_3472,N_3284);
or U6781 (N_6781,N_4607,N_3041);
xnor U6782 (N_6782,N_668,N_4510);
xor U6783 (N_6783,N_1388,N_1071);
and U6784 (N_6784,N_2646,N_4404);
and U6785 (N_6785,N_3180,N_300);
and U6786 (N_6786,N_3201,N_312);
or U6787 (N_6787,N_2624,N_3540);
or U6788 (N_6788,N_1768,N_4182);
xnor U6789 (N_6789,N_1947,N_1931);
or U6790 (N_6790,N_2169,N_1656);
nand U6791 (N_6791,N_618,N_2291);
nor U6792 (N_6792,N_2655,N_4564);
and U6793 (N_6793,N_4353,N_3498);
xor U6794 (N_6794,N_4859,N_3441);
nor U6795 (N_6795,N_1996,N_1172);
nor U6796 (N_6796,N_4716,N_3104);
or U6797 (N_6797,N_2371,N_4549);
or U6798 (N_6798,N_568,N_3595);
nor U6799 (N_6799,N_3290,N_787);
nand U6800 (N_6800,N_3262,N_4346);
nand U6801 (N_6801,N_4926,N_1245);
nand U6802 (N_6802,N_1933,N_1522);
nor U6803 (N_6803,N_4927,N_2952);
nor U6804 (N_6804,N_4596,N_3603);
nor U6805 (N_6805,N_1053,N_1981);
nor U6806 (N_6806,N_4309,N_223);
xnor U6807 (N_6807,N_267,N_3295);
nor U6808 (N_6808,N_1809,N_32);
nor U6809 (N_6809,N_4690,N_3039);
nand U6810 (N_6810,N_3874,N_875);
and U6811 (N_6811,N_2060,N_4230);
and U6812 (N_6812,N_4355,N_1692);
and U6813 (N_6813,N_3133,N_4197);
xnor U6814 (N_6814,N_1637,N_1780);
and U6815 (N_6815,N_3244,N_4186);
or U6816 (N_6816,N_1028,N_3420);
and U6817 (N_6817,N_2270,N_4447);
or U6818 (N_6818,N_1113,N_1365);
nor U6819 (N_6819,N_1974,N_2228);
and U6820 (N_6820,N_4128,N_579);
xor U6821 (N_6821,N_1329,N_2565);
nand U6822 (N_6822,N_631,N_1846);
nor U6823 (N_6823,N_3750,N_4416);
nand U6824 (N_6824,N_1279,N_4068);
nand U6825 (N_6825,N_4383,N_593);
nor U6826 (N_6826,N_982,N_1977);
and U6827 (N_6827,N_1367,N_3457);
nand U6828 (N_6828,N_4870,N_412);
xnor U6829 (N_6829,N_3856,N_4620);
and U6830 (N_6830,N_1437,N_1521);
or U6831 (N_6831,N_3605,N_1229);
nand U6832 (N_6832,N_2922,N_1548);
and U6833 (N_6833,N_706,N_2113);
nand U6834 (N_6834,N_1539,N_2529);
or U6835 (N_6835,N_145,N_4089);
nor U6836 (N_6836,N_3794,N_2972);
xnor U6837 (N_6837,N_1212,N_4034);
nor U6838 (N_6838,N_3391,N_4650);
nor U6839 (N_6839,N_3129,N_2011);
and U6840 (N_6840,N_865,N_4812);
nor U6841 (N_6841,N_3781,N_4891);
or U6842 (N_6842,N_4102,N_1312);
and U6843 (N_6843,N_555,N_4215);
and U6844 (N_6844,N_4179,N_4693);
nand U6845 (N_6845,N_1101,N_2676);
xnor U6846 (N_6846,N_4888,N_1914);
nor U6847 (N_6847,N_640,N_4421);
or U6848 (N_6848,N_3303,N_3200);
nor U6849 (N_6849,N_2936,N_2874);
and U6850 (N_6850,N_3885,N_1576);
nor U6851 (N_6851,N_2412,N_1118);
nand U6852 (N_6852,N_3873,N_2103);
or U6853 (N_6853,N_3681,N_2820);
and U6854 (N_6854,N_2502,N_2900);
or U6855 (N_6855,N_1824,N_1685);
or U6856 (N_6856,N_3827,N_2162);
or U6857 (N_6857,N_3534,N_4925);
nor U6858 (N_6858,N_3725,N_523);
and U6859 (N_6859,N_553,N_4100);
or U6860 (N_6860,N_1880,N_3384);
xnor U6861 (N_6861,N_2123,N_4413);
or U6862 (N_6862,N_4043,N_1128);
and U6863 (N_6863,N_314,N_4816);
nand U6864 (N_6864,N_1410,N_2884);
xor U6865 (N_6865,N_727,N_2043);
or U6866 (N_6866,N_286,N_3787);
nor U6867 (N_6867,N_892,N_834);
and U6868 (N_6868,N_2699,N_1844);
or U6869 (N_6869,N_1055,N_1398);
xnor U6870 (N_6870,N_676,N_4118);
or U6871 (N_6871,N_2362,N_1867);
nand U6872 (N_6872,N_4332,N_658);
nand U6873 (N_6873,N_3291,N_4271);
nand U6874 (N_6874,N_1123,N_4619);
or U6875 (N_6875,N_128,N_968);
nand U6876 (N_6876,N_4191,N_3272);
nor U6877 (N_6877,N_3057,N_3537);
nand U6878 (N_6878,N_781,N_1080);
nor U6879 (N_6879,N_653,N_1100);
or U6880 (N_6880,N_442,N_4465);
and U6881 (N_6881,N_466,N_895);
or U6882 (N_6882,N_4576,N_1415);
and U6883 (N_6883,N_4739,N_4214);
nand U6884 (N_6884,N_1278,N_4412);
xor U6885 (N_6885,N_3609,N_4001);
and U6886 (N_6886,N_4918,N_4097);
nand U6887 (N_6887,N_4666,N_1765);
nor U6888 (N_6888,N_4037,N_1909);
and U6889 (N_6889,N_2447,N_2084);
nor U6890 (N_6890,N_3871,N_2037);
and U6891 (N_6891,N_2659,N_837);
or U6892 (N_6892,N_1706,N_1121);
or U6893 (N_6893,N_177,N_4183);
nor U6894 (N_6894,N_813,N_1955);
nor U6895 (N_6895,N_4815,N_1953);
nor U6896 (N_6896,N_1505,N_1023);
or U6897 (N_6897,N_4844,N_216);
or U6898 (N_6898,N_1697,N_2795);
nand U6899 (N_6899,N_683,N_3143);
or U6900 (N_6900,N_3424,N_1103);
nand U6901 (N_6901,N_2192,N_4553);
nor U6902 (N_6902,N_1106,N_1893);
and U6903 (N_6903,N_1222,N_1347);
and U6904 (N_6904,N_2280,N_4026);
and U6905 (N_6905,N_533,N_1265);
and U6906 (N_6906,N_1564,N_2929);
or U6907 (N_6907,N_2136,N_1729);
or U6908 (N_6908,N_4275,N_679);
nand U6909 (N_6909,N_4269,N_4448);
nand U6910 (N_6910,N_4290,N_2390);
nor U6911 (N_6911,N_4877,N_1942);
nor U6912 (N_6912,N_976,N_652);
or U6913 (N_6913,N_2752,N_1535);
or U6914 (N_6914,N_1376,N_4303);
and U6915 (N_6915,N_1183,N_592);
nand U6916 (N_6916,N_2363,N_4698);
nand U6917 (N_6917,N_4088,N_717);
and U6918 (N_6918,N_4964,N_3795);
or U6919 (N_6919,N_4327,N_2045);
and U6920 (N_6920,N_3641,N_88);
nor U6921 (N_6921,N_2920,N_2782);
xor U6922 (N_6922,N_2573,N_4644);
and U6923 (N_6923,N_1991,N_4518);
nor U6924 (N_6924,N_3348,N_1407);
nor U6925 (N_6925,N_2629,N_2602);
and U6926 (N_6926,N_4180,N_348);
and U6927 (N_6927,N_4982,N_1083);
and U6928 (N_6928,N_1671,N_1723);
or U6929 (N_6929,N_2648,N_344);
nand U6930 (N_6930,N_324,N_70);
or U6931 (N_6931,N_824,N_2829);
nor U6932 (N_6932,N_1699,N_3780);
nand U6933 (N_6933,N_883,N_699);
and U6934 (N_6934,N_360,N_2825);
nor U6935 (N_6935,N_3846,N_234);
nor U6936 (N_6936,N_4050,N_2684);
or U6937 (N_6937,N_2081,N_113);
and U6938 (N_6938,N_1612,N_2621);
or U6939 (N_6939,N_4542,N_3367);
or U6940 (N_6940,N_3497,N_3730);
nand U6941 (N_6941,N_1778,N_842);
nor U6942 (N_6942,N_2940,N_3191);
or U6943 (N_6943,N_1549,N_3709);
and U6944 (N_6944,N_4736,N_119);
and U6945 (N_6945,N_180,N_44);
nand U6946 (N_6946,N_192,N_3580);
or U6947 (N_6947,N_2115,N_482);
nand U6948 (N_6948,N_3470,N_3286);
nor U6949 (N_6949,N_3387,N_3331);
nor U6950 (N_6950,N_4052,N_2961);
or U6951 (N_6951,N_4683,N_1916);
and U6952 (N_6952,N_3451,N_2620);
and U6953 (N_6953,N_2483,N_4344);
xor U6954 (N_6954,N_3229,N_2273);
or U6955 (N_6955,N_206,N_3428);
and U6956 (N_6956,N_2450,N_804);
or U6957 (N_6957,N_4528,N_1733);
and U6958 (N_6958,N_2356,N_1383);
or U6959 (N_6959,N_4762,N_8);
nor U6960 (N_6960,N_2370,N_518);
nand U6961 (N_6961,N_3719,N_3346);
or U6962 (N_6962,N_889,N_1590);
and U6963 (N_6963,N_2926,N_2995);
nand U6964 (N_6964,N_1795,N_3653);
nor U6965 (N_6965,N_3366,N_4783);
nor U6966 (N_6966,N_599,N_588);
nand U6967 (N_6967,N_2444,N_1322);
or U6968 (N_6968,N_2340,N_3651);
nand U6969 (N_6969,N_567,N_1326);
xor U6970 (N_6970,N_368,N_4501);
or U6971 (N_6971,N_480,N_1189);
or U6972 (N_6972,N_4928,N_2980);
nor U6973 (N_6973,N_3615,N_510);
and U6974 (N_6974,N_3597,N_4654);
xnor U6975 (N_6975,N_3738,N_1896);
or U6976 (N_6976,N_2431,N_1529);
and U6977 (N_6977,N_1007,N_1039);
nor U6978 (N_6978,N_1807,N_2841);
nand U6979 (N_6979,N_2056,N_2590);
or U6980 (N_6980,N_1948,N_238);
nand U6981 (N_6981,N_1337,N_2488);
and U6982 (N_6982,N_4466,N_3699);
xnor U6983 (N_6983,N_179,N_1818);
and U6984 (N_6984,N_4600,N_4475);
nand U6985 (N_6985,N_122,N_764);
and U6986 (N_6986,N_4101,N_2179);
nand U6987 (N_6987,N_1877,N_3876);
and U6988 (N_6988,N_1631,N_355);
and U6989 (N_6989,N_2223,N_1079);
or U6990 (N_6990,N_635,N_3136);
or U6991 (N_6991,N_3920,N_2110);
nand U6992 (N_6992,N_107,N_2542);
and U6993 (N_6993,N_692,N_4393);
nor U6994 (N_6994,N_2913,N_4458);
nand U6995 (N_6995,N_58,N_4099);
nor U6996 (N_6996,N_3571,N_319);
nor U6997 (N_6997,N_2688,N_1978);
xor U6998 (N_6998,N_666,N_4636);
xnor U6999 (N_6999,N_3608,N_1048);
or U7000 (N_7000,N_4184,N_1595);
xor U7001 (N_7001,N_4374,N_4121);
nor U7002 (N_7002,N_1114,N_3572);
and U7003 (N_7003,N_4954,N_703);
nor U7004 (N_7004,N_1816,N_1427);
nor U7005 (N_7005,N_2085,N_710);
nand U7006 (N_7006,N_506,N_2997);
xor U7007 (N_7007,N_3731,N_3935);
nor U7008 (N_7008,N_2031,N_1133);
or U7009 (N_7009,N_4627,N_3579);
nor U7010 (N_7010,N_457,N_4862);
nor U7011 (N_7011,N_4513,N_4252);
nor U7012 (N_7012,N_2697,N_1679);
or U7013 (N_7013,N_2030,N_1334);
xor U7014 (N_7014,N_1555,N_4509);
nand U7015 (N_7015,N_986,N_4920);
and U7016 (N_7016,N_104,N_1497);
nor U7017 (N_7017,N_607,N_171);
or U7018 (N_7018,N_406,N_2725);
nand U7019 (N_7019,N_2912,N_3068);
xor U7020 (N_7020,N_2816,N_605);
nand U7021 (N_7021,N_3061,N_838);
nand U7022 (N_7022,N_2764,N_651);
or U7023 (N_7023,N_1837,N_2924);
nor U7024 (N_7024,N_1950,N_2137);
or U7025 (N_7025,N_1145,N_22);
or U7026 (N_7026,N_531,N_3408);
xor U7027 (N_7027,N_3217,N_2096);
xor U7028 (N_7028,N_4539,N_3501);
nand U7029 (N_7029,N_3682,N_3710);
nand U7030 (N_7030,N_2691,N_3455);
nand U7031 (N_7031,N_3359,N_1368);
or U7032 (N_7032,N_2478,N_1750);
nand U7033 (N_7033,N_4514,N_1634);
xor U7034 (N_7034,N_2153,N_2960);
and U7035 (N_7035,N_1386,N_672);
nor U7036 (N_7036,N_900,N_4408);
nand U7037 (N_7037,N_342,N_3477);
or U7038 (N_7038,N_273,N_33);
nand U7039 (N_7039,N_1594,N_2376);
nand U7040 (N_7040,N_3135,N_1377);
and U7041 (N_7041,N_2388,N_4338);
nand U7042 (N_7042,N_4545,N_1044);
xnor U7043 (N_7043,N_74,N_4702);
and U7044 (N_7044,N_2710,N_560);
nand U7045 (N_7045,N_3566,N_1233);
or U7046 (N_7046,N_1195,N_1509);
and U7047 (N_7047,N_3718,N_2069);
and U7048 (N_7048,N_2204,N_3040);
or U7049 (N_7049,N_2776,N_1434);
xnor U7050 (N_7050,N_4166,N_3558);
and U7051 (N_7051,N_496,N_214);
and U7052 (N_7052,N_939,N_2167);
or U7053 (N_7053,N_4956,N_1186);
or U7054 (N_7054,N_4115,N_4585);
nand U7055 (N_7055,N_4750,N_4823);
xor U7056 (N_7056,N_2460,N_4411);
xor U7057 (N_7057,N_1636,N_1060);
xnor U7058 (N_7058,N_1759,N_603);
or U7059 (N_7059,N_1224,N_4519);
nor U7060 (N_7060,N_1633,N_124);
nor U7061 (N_7061,N_786,N_1826);
nor U7062 (N_7062,N_1918,N_3289);
nand U7063 (N_7063,N_4170,N_287);
xnor U7064 (N_7064,N_1689,N_3527);
and U7065 (N_7065,N_3007,N_3910);
or U7066 (N_7066,N_3440,N_2986);
xnor U7067 (N_7067,N_2127,N_133);
nand U7068 (N_7068,N_1115,N_1638);
nor U7069 (N_7069,N_2907,N_4013);
nand U7070 (N_7070,N_772,N_2263);
xor U7071 (N_7071,N_3850,N_1474);
nand U7072 (N_7072,N_2556,N_311);
nand U7073 (N_7073,N_3236,N_3248);
xor U7074 (N_7074,N_817,N_4521);
nand U7075 (N_7075,N_157,N_1209);
and U7076 (N_7076,N_1997,N_4824);
nand U7077 (N_7077,N_2028,N_1919);
nand U7078 (N_7078,N_4967,N_2098);
or U7079 (N_7079,N_4633,N_1618);
or U7080 (N_7080,N_2240,N_797);
nand U7081 (N_7081,N_1982,N_4400);
nor U7082 (N_7082,N_3637,N_243);
or U7083 (N_7083,N_3296,N_3643);
nand U7084 (N_7084,N_785,N_2615);
nand U7085 (N_7085,N_2524,N_4293);
nand U7086 (N_7086,N_1281,N_990);
nor U7087 (N_7087,N_2497,N_934);
and U7088 (N_7088,N_4212,N_886);
and U7089 (N_7089,N_1647,N_4635);
nor U7090 (N_7090,N_2544,N_4738);
nor U7091 (N_7091,N_445,N_423);
nor U7092 (N_7092,N_2873,N_2685);
nor U7093 (N_7093,N_4807,N_4780);
nor U7094 (N_7094,N_3288,N_373);
nor U7095 (N_7095,N_4348,N_2626);
and U7096 (N_7096,N_1119,N_1196);
or U7097 (N_7097,N_4064,N_2862);
xor U7098 (N_7098,N_3390,N_1742);
and U7099 (N_7099,N_4276,N_1058);
xnor U7100 (N_7100,N_3056,N_825);
or U7101 (N_7101,N_2735,N_4451);
and U7102 (N_7102,N_1784,N_2395);
nor U7103 (N_7103,N_1085,N_4670);
and U7104 (N_7104,N_3418,N_4822);
xnor U7105 (N_7105,N_4117,N_3300);
nand U7106 (N_7106,N_2652,N_3083);
or U7107 (N_7107,N_4685,N_598);
nand U7108 (N_7108,N_879,N_4640);
or U7109 (N_7109,N_3735,N_1843);
or U7110 (N_7110,N_970,N_89);
and U7111 (N_7111,N_962,N_9);
nand U7112 (N_7112,N_897,N_3664);
or U7113 (N_7113,N_4268,N_4084);
and U7114 (N_7114,N_2732,N_4263);
or U7115 (N_7115,N_3639,N_3484);
or U7116 (N_7116,N_843,N_1869);
nand U7117 (N_7117,N_1772,N_4235);
nor U7118 (N_7118,N_2082,N_1929);
xnor U7119 (N_7119,N_3121,N_4845);
or U7120 (N_7120,N_975,N_792);
nand U7121 (N_7121,N_3378,N_1413);
nand U7122 (N_7122,N_3831,N_1293);
nor U7123 (N_7123,N_1082,N_2189);
xnor U7124 (N_7124,N_711,N_827);
nor U7125 (N_7125,N_1523,N_2430);
nand U7126 (N_7126,N_2677,N_4165);
or U7127 (N_7127,N_1853,N_163);
or U7128 (N_7128,N_2319,N_1370);
and U7129 (N_7129,N_459,N_3551);
nor U7130 (N_7130,N_674,N_3149);
nand U7131 (N_7131,N_1412,N_3161);
nor U7132 (N_7132,N_425,N_2108);
nor U7133 (N_7133,N_981,N_4155);
xnor U7134 (N_7134,N_802,N_698);
or U7135 (N_7135,N_2410,N_1627);
or U7136 (N_7136,N_3627,N_4071);
or U7137 (N_7137,N_3649,N_4546);
and U7138 (N_7138,N_3866,N_1992);
nand U7139 (N_7139,N_2302,N_1393);
or U7140 (N_7140,N_2059,N_4354);
or U7141 (N_7141,N_3074,N_142);
nand U7142 (N_7142,N_1483,N_146);
nand U7143 (N_7143,N_2774,N_2905);
nand U7144 (N_7144,N_4876,N_684);
and U7145 (N_7145,N_281,N_1318);
nor U7146 (N_7146,N_1282,N_4329);
nand U7147 (N_7147,N_224,N_4158);
and U7148 (N_7148,N_270,N_4568);
xor U7149 (N_7149,N_4682,N_3823);
xor U7150 (N_7150,N_2523,N_4479);
or U7151 (N_7151,N_2731,N_1012);
nand U7152 (N_7152,N_4730,N_1441);
and U7153 (N_7153,N_4377,N_4684);
nor U7154 (N_7154,N_591,N_1297);
or U7155 (N_7155,N_840,N_93);
nor U7156 (N_7156,N_474,N_3429);
nor U7157 (N_7157,N_3126,N_4922);
nand U7158 (N_7158,N_1676,N_3555);
nand U7159 (N_7159,N_541,N_3144);
nand U7160 (N_7160,N_1941,N_4443);
nand U7161 (N_7161,N_4826,N_1379);
nor U7162 (N_7162,N_1338,N_1792);
nor U7163 (N_7163,N_1575,N_2522);
or U7164 (N_7164,N_2177,N_1230);
and U7165 (N_7165,N_2375,N_2306);
xor U7166 (N_7166,N_3924,N_1794);
or U7167 (N_7167,N_2632,N_3006);
nor U7168 (N_7168,N_3361,N_4491);
and U7169 (N_7169,N_4947,N_1695);
or U7170 (N_7170,N_913,N_3782);
xor U7171 (N_7171,N_2834,N_2400);
and U7172 (N_7172,N_932,N_1247);
nor U7173 (N_7173,N_3923,N_4777);
and U7174 (N_7174,N_4282,N_3215);
nor U7175 (N_7175,N_3687,N_2600);
nor U7176 (N_7176,N_2349,N_4032);
nor U7177 (N_7177,N_1726,N_712);
nor U7178 (N_7178,N_2851,N_3199);
nand U7179 (N_7179,N_4811,N_4547);
nor U7180 (N_7180,N_2199,N_550);
nor U7181 (N_7181,N_4022,N_4176);
or U7182 (N_7182,N_4286,N_2970);
nor U7183 (N_7183,N_758,N_3892);
nor U7184 (N_7184,N_3335,N_3071);
nand U7185 (N_7185,N_166,N_527);
nand U7186 (N_7186,N_2563,N_4250);
nor U7187 (N_7187,N_3748,N_2250);
or U7188 (N_7188,N_3982,N_762);
nor U7189 (N_7189,N_2811,N_4302);
and U7190 (N_7190,N_4123,N_1429);
nand U7191 (N_7191,N_4834,N_4159);
or U7192 (N_7192,N_62,N_2549);
or U7193 (N_7193,N_3902,N_1900);
nor U7194 (N_7194,N_3218,N_3865);
nand U7195 (N_7195,N_4960,N_903);
or U7196 (N_7196,N_3562,N_2141);
or U7197 (N_7197,N_1248,N_714);
and U7198 (N_7198,N_3400,N_1859);
or U7199 (N_7199,N_162,N_1995);
xnor U7200 (N_7200,N_4757,N_2680);
or U7201 (N_7201,N_3175,N_196);
or U7202 (N_7202,N_2824,N_2453);
and U7203 (N_7203,N_3809,N_3251);
xnor U7204 (N_7204,N_2101,N_4828);
or U7205 (N_7205,N_3714,N_1927);
nand U7206 (N_7206,N_661,N_3207);
xor U7207 (N_7207,N_3694,N_2510);
nor U7208 (N_7208,N_1542,N_4818);
or U7209 (N_7209,N_3024,N_4966);
nand U7210 (N_7210,N_1820,N_1500);
nor U7211 (N_7211,N_3901,N_4852);
nor U7212 (N_7212,N_280,N_3685);
xnor U7213 (N_7213,N_3908,N_3001);
and U7214 (N_7214,N_4856,N_3220);
xnor U7215 (N_7215,N_4957,N_722);
or U7216 (N_7216,N_3415,N_3774);
and U7217 (N_7217,N_2365,N_2539);
nand U7218 (N_7218,N_1620,N_126);
and U7219 (N_7219,N_4775,N_3405);
and U7220 (N_7220,N_3492,N_3593);
nand U7221 (N_7221,N_4614,N_2708);
or U7222 (N_7222,N_3801,N_2996);
or U7223 (N_7223,N_356,N_1011);
nor U7224 (N_7224,N_629,N_3090);
and U7225 (N_7225,N_3233,N_3863);
or U7226 (N_7226,N_4538,N_2116);
nand U7227 (N_7227,N_1416,N_4638);
or U7228 (N_7228,N_3556,N_2950);
nor U7229 (N_7229,N_2515,N_376);
xnor U7230 (N_7230,N_2385,N_1405);
or U7231 (N_7231,N_833,N_301);
xor U7232 (N_7232,N_1686,N_2724);
nor U7233 (N_7233,N_4299,N_4932);
or U7234 (N_7234,N_3592,N_4660);
and U7235 (N_7235,N_2866,N_3108);
nand U7236 (N_7236,N_3421,N_1092);
and U7237 (N_7237,N_3465,N_1670);
nand U7238 (N_7238,N_3987,N_1989);
or U7239 (N_7239,N_25,N_2581);
nand U7240 (N_7240,N_4861,N_4243);
or U7241 (N_7241,N_3285,N_4322);
or U7242 (N_7242,N_4517,N_4414);
nor U7243 (N_7243,N_2797,N_4999);
and U7244 (N_7244,N_2749,N_2399);
or U7245 (N_7245,N_3198,N_559);
nor U7246 (N_7246,N_2434,N_2948);
and U7247 (N_7247,N_411,N_3872);
nor U7248 (N_7248,N_1077,N_3181);
nor U7249 (N_7249,N_801,N_2978);
or U7250 (N_7250,N_336,N_3008);
nor U7251 (N_7251,N_96,N_776);
nor U7252 (N_7252,N_2161,N_3906);
nor U7253 (N_7253,N_2771,N_2946);
nor U7254 (N_7254,N_4363,N_4610);
xnor U7255 (N_7255,N_4741,N_2472);
or U7256 (N_7256,N_2571,N_4004);
nand U7257 (N_7257,N_966,N_3313);
nor U7258 (N_7258,N_3818,N_429);
nor U7259 (N_7259,N_1234,N_728);
nor U7260 (N_7260,N_1315,N_1600);
or U7261 (N_7261,N_4782,N_2354);
nand U7262 (N_7262,N_4445,N_1628);
or U7263 (N_7263,N_2916,N_791);
nor U7264 (N_7264,N_4193,N_3280);
and U7265 (N_7265,N_1105,N_4804);
and U7266 (N_7266,N_3372,N_2887);
nand U7267 (N_7267,N_1563,N_3706);
xnor U7268 (N_7268,N_381,N_2566);
nand U7269 (N_7269,N_4061,N_1124);
nor U7270 (N_7270,N_2198,N_1815);
nand U7271 (N_7271,N_4548,N_2813);
and U7272 (N_7272,N_2702,N_4653);
nor U7273 (N_7273,N_3905,N_1533);
or U7274 (N_7274,N_2639,N_4616);
nor U7275 (N_7275,N_4536,N_2673);
and U7276 (N_7276,N_75,N_1446);
nand U7277 (N_7277,N_1239,N_3234);
or U7278 (N_7278,N_3317,N_4931);
nor U7279 (N_7279,N_507,N_54);
and U7280 (N_7280,N_3933,N_3055);
nor U7281 (N_7281,N_985,N_1371);
nor U7282 (N_7282,N_2463,N_4867);
nand U7283 (N_7283,N_3278,N_3696);
xor U7284 (N_7284,N_2683,N_1897);
xor U7285 (N_7285,N_614,N_291);
nor U7286 (N_7286,N_15,N_3282);
or U7287 (N_7287,N_193,N_3190);
nand U7288 (N_7288,N_4896,N_3197);
or U7289 (N_7289,N_3193,N_586);
nand U7290 (N_7290,N_4229,N_3050);
and U7291 (N_7291,N_4930,N_1099);
nand U7292 (N_7292,N_771,N_1857);
and U7293 (N_7293,N_169,N_2909);
nor U7294 (N_7294,N_4527,N_150);
or U7295 (N_7295,N_2951,N_2077);
nor U7296 (N_7296,N_819,N_3445);
and U7297 (N_7297,N_2269,N_3672);
or U7298 (N_7298,N_3413,N_4800);
xor U7299 (N_7299,N_2479,N_1623);
xnor U7300 (N_7300,N_3092,N_3444);
nor U7301 (N_7301,N_681,N_1517);
nor U7302 (N_7302,N_2050,N_1829);
and U7303 (N_7303,N_1173,N_498);
nand U7304 (N_7304,N_4605,N_2281);
or U7305 (N_7305,N_3582,N_3000);
nand U7306 (N_7306,N_902,N_1166);
and U7307 (N_7307,N_4646,N_2738);
nor U7308 (N_7308,N_4817,N_3192);
or U7309 (N_7309,N_3209,N_4081);
nand U7310 (N_7310,N_724,N_4304);
nor U7311 (N_7311,N_2910,N_3638);
xnor U7312 (N_7312,N_4096,N_3791);
nand U7313 (N_7313,N_4764,N_4499);
nor U7314 (N_7314,N_3744,N_383);
or U7315 (N_7315,N_1970,N_4866);
and U7316 (N_7316,N_1126,N_1540);
and U7317 (N_7317,N_3456,N_3803);
nand U7318 (N_7318,N_1938,N_220);
or U7319 (N_7319,N_1098,N_181);
nand U7320 (N_7320,N_3072,N_1091);
or U7321 (N_7321,N_2517,N_4280);
and U7322 (N_7322,N_84,N_2493);
and U7323 (N_7323,N_4419,N_2570);
and U7324 (N_7324,N_795,N_953);
nand U7325 (N_7325,N_492,N_68);
nor U7326 (N_7326,N_2777,N_4313);
nand U7327 (N_7327,N_2315,N_167);
and U7328 (N_7328,N_872,N_283);
nand U7329 (N_7329,N_4232,N_1722);
xnor U7330 (N_7330,N_3600,N_4871);
nor U7331 (N_7331,N_426,N_3321);
or U7332 (N_7332,N_1658,N_408);
and U7333 (N_7333,N_1024,N_750);
or U7334 (N_7334,N_2846,N_4722);
or U7335 (N_7335,N_3091,N_2805);
nor U7336 (N_7336,N_144,N_1714);
nor U7337 (N_7337,N_1721,N_4505);
or U7338 (N_7338,N_3228,N_4150);
nand U7339 (N_7339,N_3377,N_3573);
nand U7340 (N_7340,N_2589,N_1084);
or U7341 (N_7341,N_1394,N_1969);
nor U7342 (N_7342,N_3480,N_241);
nand U7343 (N_7343,N_1851,N_1951);
nor U7344 (N_7344,N_2893,N_4201);
or U7345 (N_7345,N_831,N_1644);
nor U7346 (N_7346,N_382,N_4758);
and U7347 (N_7347,N_1476,N_1781);
and U7348 (N_7348,N_596,N_3403);
nand U7349 (N_7349,N_3151,N_3155);
nor U7350 (N_7350,N_816,N_894);
and U7351 (N_7351,N_1905,N_3283);
or U7352 (N_7352,N_3109,N_4733);
nand U7353 (N_7353,N_380,N_3439);
and U7354 (N_7354,N_378,N_1677);
nand U7355 (N_7355,N_4127,N_1684);
nor U7356 (N_7356,N_2501,N_2293);
or U7357 (N_7357,N_6,N_175);
and U7358 (N_7358,N_940,N_3721);
nor U7359 (N_7359,N_250,N_3521);
nand U7360 (N_7360,N_1006,N_2957);
nand U7361 (N_7361,N_1885,N_820);
nand U7362 (N_7362,N_2417,N_3268);
nand U7363 (N_7363,N_326,N_3243);
or U7364 (N_7364,N_285,N_3793);
nand U7365 (N_7365,N_419,N_4531);
xor U7366 (N_7366,N_1848,N_351);
or U7367 (N_7367,N_3552,N_2888);
nor U7368 (N_7368,N_4988,N_2562);
or U7369 (N_7369,N_565,N_2880);
xnor U7370 (N_7370,N_63,N_3076);
nand U7371 (N_7371,N_884,N_2419);
nor U7372 (N_7372,N_4469,N_4754);
nand U7373 (N_7373,N_989,N_645);
and U7374 (N_7374,N_973,N_2100);
xor U7375 (N_7375,N_3380,N_2849);
and U7376 (N_7376,N_1328,N_1693);
nor U7377 (N_7377,N_2041,N_3085);
nand U7378 (N_7378,N_1139,N_4085);
nor U7379 (N_7379,N_3146,N_1839);
and U7380 (N_7380,N_4350,N_569);
nand U7381 (N_7381,N_3150,N_2206);
nand U7382 (N_7382,N_409,N_2203);
nor U7383 (N_7383,N_2974,N_3172);
xnor U7384 (N_7384,N_108,N_2745);
xor U7385 (N_7385,N_3602,N_1808);
xnor U7386 (N_7386,N_2484,N_4511);
or U7387 (N_7387,N_4983,N_4980);
nor U7388 (N_7388,N_896,N_891);
nand U7389 (N_7389,N_3756,N_2424);
nand U7390 (N_7390,N_637,N_4442);
or U7391 (N_7391,N_828,N_1009);
and U7392 (N_7392,N_2163,N_2516);
xor U7393 (N_7393,N_3574,N_4330);
or U7394 (N_7394,N_2614,N_3503);
or U7395 (N_7395,N_4714,N_3611);
nand U7396 (N_7396,N_3616,N_3712);
nand U7397 (N_7397,N_848,N_2083);
nor U7398 (N_7398,N_3005,N_3564);
nand U7399 (N_7399,N_4296,N_3059);
nand U7400 (N_7400,N_4981,N_746);
nor U7401 (N_7401,N_1335,N_2391);
and U7402 (N_7402,N_2454,N_4634);
nand U7403 (N_7403,N_2641,N_1275);
xor U7404 (N_7404,N_1926,N_1038);
and U7405 (N_7405,N_2531,N_3152);
or U7406 (N_7406,N_3934,N_186);
nand U7407 (N_7407,N_3235,N_4622);
or U7408 (N_7408,N_805,N_2014);
and U7409 (N_7409,N_3163,N_1199);
nand U7410 (N_7410,N_309,N_2018);
and U7411 (N_7411,N_2949,N_4902);
or U7412 (N_7412,N_226,N_2859);
and U7413 (N_7413,N_509,N_930);
and U7414 (N_7414,N_2181,N_1757);
nand U7415 (N_7415,N_3255,N_1608);
or U7416 (N_7416,N_2521,N_2593);
nand U7417 (N_7417,N_2991,N_3112);
nand U7418 (N_7418,N_2048,N_4283);
xor U7419 (N_7419,N_4887,N_3127);
and U7420 (N_7420,N_3613,N_1599);
nor U7421 (N_7421,N_3029,N_4385);
and U7422 (N_7422,N_4450,N_4075);
and U7423 (N_7423,N_2010,N_2616);
or U7424 (N_7424,N_3043,N_855);
xor U7425 (N_7425,N_467,N_2328);
nand U7426 (N_7426,N_4360,N_4133);
nor U7427 (N_7427,N_318,N_3784);
and U7428 (N_7428,N_1004,N_4041);
and U7429 (N_7429,N_3594,N_1353);
nand U7430 (N_7430,N_570,N_3816);
nor U7431 (N_7431,N_4909,N_4837);
nand U7432 (N_7432,N_3264,N_4173);
nand U7433 (N_7433,N_4381,N_2384);
and U7434 (N_7434,N_4744,N_4039);
or U7435 (N_7435,N_174,N_1046);
nand U7436 (N_7436,N_4141,N_4802);
or U7437 (N_7437,N_1530,N_4842);
and U7438 (N_7438,N_3037,N_4608);
nor U7439 (N_7439,N_3606,N_4515);
or U7440 (N_7440,N_3995,N_2798);
nor U7441 (N_7441,N_1773,N_1653);
nand U7442 (N_7442,N_2271,N_284);
or U7443 (N_7443,N_21,N_384);
xnor U7444 (N_7444,N_486,N_773);
nor U7445 (N_7445,N_1499,N_4036);
xor U7446 (N_7446,N_4561,N_4395);
xnor U7447 (N_7447,N_1251,N_0);
and U7448 (N_7448,N_2736,N_2534);
or U7449 (N_7449,N_3752,N_500);
or U7450 (N_7450,N_3154,N_3621);
or U7451 (N_7451,N_2036,N_623);
nor U7452 (N_7452,N_3414,N_3927);
nor U7453 (N_7453,N_675,N_4792);
and U7454 (N_7454,N_3277,N_1958);
and U7455 (N_7455,N_4678,N_1855);
and U7456 (N_7456,N_3955,N_3506);
nand U7457 (N_7457,N_4795,N_2818);
and U7458 (N_7458,N_4314,N_4418);
nor U7459 (N_7459,N_3106,N_4558);
or U7460 (N_7460,N_2238,N_3948);
and U7461 (N_7461,N_4365,N_2939);
nand U7462 (N_7462,N_723,N_3344);
nand U7463 (N_7463,N_713,N_172);
nor U7464 (N_7464,N_4203,N_904);
nor U7465 (N_7465,N_81,N_3123);
xor U7466 (N_7466,N_4959,N_1790);
nor U7467 (N_7467,N_2930,N_4840);
and U7468 (N_7468,N_436,N_2065);
nand U7469 (N_7469,N_3269,N_3741);
and U7470 (N_7470,N_2803,N_1702);
and U7471 (N_7471,N_3713,N_3003);
nor U7472 (N_7472,N_1967,N_1565);
nand U7473 (N_7473,N_4570,N_4006);
xnor U7474 (N_7474,N_2071,N_3310);
xor U7475 (N_7475,N_1520,N_3489);
and U7476 (N_7476,N_996,N_3038);
or U7477 (N_7477,N_1614,N_229);
or U7478 (N_7478,N_2140,N_3825);
xor U7479 (N_7479,N_2832,N_1797);
and U7480 (N_7480,N_936,N_2156);
or U7481 (N_7481,N_2262,N_176);
or U7482 (N_7482,N_1414,N_2079);
and U7483 (N_7483,N_362,N_2339);
or U7484 (N_7484,N_625,N_2737);
and U7485 (N_7485,N_4808,N_4892);
or U7486 (N_7486,N_3528,N_1811);
xor U7487 (N_7487,N_1668,N_331);
xnor U7488 (N_7488,N_3166,N_26);
nor U7489 (N_7489,N_3704,N_151);
nor U7490 (N_7490,N_1457,N_191);
or U7491 (N_7491,N_94,N_3270);
nand U7492 (N_7492,N_1299,N_3670);
nor U7493 (N_7493,N_394,N_2842);
and U7494 (N_7494,N_3379,N_1748);
nor U7495 (N_7495,N_1649,N_946);
nor U7496 (N_7496,N_475,N_520);
xnor U7497 (N_7497,N_1179,N_554);
nor U7498 (N_7498,N_2330,N_2975);
nand U7499 (N_7499,N_3715,N_1090);
or U7500 (N_7500,N_173,N_447);
and U7501 (N_7501,N_2031,N_2572);
and U7502 (N_7502,N_3288,N_1827);
and U7503 (N_7503,N_2375,N_4851);
nor U7504 (N_7504,N_3036,N_1185);
nor U7505 (N_7505,N_944,N_4487);
and U7506 (N_7506,N_1076,N_4548);
and U7507 (N_7507,N_2911,N_1679);
nor U7508 (N_7508,N_750,N_2468);
and U7509 (N_7509,N_1236,N_602);
and U7510 (N_7510,N_3920,N_3526);
nor U7511 (N_7511,N_2415,N_4156);
and U7512 (N_7512,N_4912,N_2724);
xnor U7513 (N_7513,N_493,N_321);
or U7514 (N_7514,N_899,N_3500);
xnor U7515 (N_7515,N_2865,N_370);
or U7516 (N_7516,N_1016,N_2347);
nor U7517 (N_7517,N_3112,N_456);
or U7518 (N_7518,N_822,N_1552);
or U7519 (N_7519,N_3285,N_828);
nor U7520 (N_7520,N_3735,N_1774);
and U7521 (N_7521,N_2709,N_4028);
and U7522 (N_7522,N_617,N_1764);
nor U7523 (N_7523,N_1909,N_563);
and U7524 (N_7524,N_3241,N_4925);
xor U7525 (N_7525,N_303,N_840);
nor U7526 (N_7526,N_4920,N_4474);
and U7527 (N_7527,N_537,N_1614);
nor U7528 (N_7528,N_2150,N_267);
and U7529 (N_7529,N_3620,N_3087);
or U7530 (N_7530,N_4899,N_270);
nor U7531 (N_7531,N_476,N_1745);
nor U7532 (N_7532,N_720,N_4260);
nand U7533 (N_7533,N_4228,N_409);
nor U7534 (N_7534,N_4596,N_4695);
or U7535 (N_7535,N_3893,N_2484);
nor U7536 (N_7536,N_2900,N_3509);
and U7537 (N_7537,N_2265,N_1966);
nor U7538 (N_7538,N_1300,N_3706);
nand U7539 (N_7539,N_3498,N_610);
nor U7540 (N_7540,N_1126,N_2498);
and U7541 (N_7541,N_3246,N_4582);
nor U7542 (N_7542,N_215,N_4390);
nor U7543 (N_7543,N_1528,N_4899);
and U7544 (N_7544,N_2704,N_4900);
or U7545 (N_7545,N_4424,N_1097);
or U7546 (N_7546,N_3742,N_1439);
and U7547 (N_7547,N_4343,N_1487);
nand U7548 (N_7548,N_1797,N_2777);
xor U7549 (N_7549,N_374,N_1236);
or U7550 (N_7550,N_4009,N_3080);
and U7551 (N_7551,N_2746,N_2394);
or U7552 (N_7552,N_1377,N_4421);
nand U7553 (N_7553,N_575,N_3063);
nand U7554 (N_7554,N_4561,N_2035);
nand U7555 (N_7555,N_1044,N_2927);
nand U7556 (N_7556,N_1886,N_498);
nand U7557 (N_7557,N_19,N_4035);
or U7558 (N_7558,N_765,N_4814);
nor U7559 (N_7559,N_70,N_2239);
xor U7560 (N_7560,N_330,N_3997);
or U7561 (N_7561,N_4747,N_1863);
nand U7562 (N_7562,N_4435,N_622);
or U7563 (N_7563,N_4979,N_599);
nand U7564 (N_7564,N_571,N_808);
nor U7565 (N_7565,N_1187,N_1093);
xor U7566 (N_7566,N_318,N_4442);
xnor U7567 (N_7567,N_4631,N_3173);
nor U7568 (N_7568,N_783,N_3837);
and U7569 (N_7569,N_1622,N_222);
or U7570 (N_7570,N_925,N_2010);
nand U7571 (N_7571,N_4295,N_318);
and U7572 (N_7572,N_2511,N_3936);
nor U7573 (N_7573,N_3216,N_1695);
or U7574 (N_7574,N_906,N_4611);
and U7575 (N_7575,N_4820,N_1203);
xnor U7576 (N_7576,N_3573,N_1212);
and U7577 (N_7577,N_1637,N_788);
nor U7578 (N_7578,N_1005,N_3419);
nor U7579 (N_7579,N_147,N_2665);
or U7580 (N_7580,N_4504,N_986);
xor U7581 (N_7581,N_2976,N_912);
or U7582 (N_7582,N_2778,N_2721);
or U7583 (N_7583,N_2618,N_3213);
nand U7584 (N_7584,N_4237,N_3052);
xnor U7585 (N_7585,N_4883,N_821);
and U7586 (N_7586,N_1909,N_2392);
or U7587 (N_7587,N_2156,N_4029);
and U7588 (N_7588,N_3832,N_2313);
and U7589 (N_7589,N_4201,N_57);
and U7590 (N_7590,N_233,N_786);
and U7591 (N_7591,N_74,N_686);
and U7592 (N_7592,N_925,N_942);
nor U7593 (N_7593,N_231,N_4859);
nand U7594 (N_7594,N_1786,N_1961);
nand U7595 (N_7595,N_708,N_3307);
and U7596 (N_7596,N_3127,N_3828);
and U7597 (N_7597,N_1994,N_1977);
and U7598 (N_7598,N_1043,N_3369);
or U7599 (N_7599,N_2080,N_895);
nand U7600 (N_7600,N_4980,N_1756);
or U7601 (N_7601,N_2610,N_277);
and U7602 (N_7602,N_4699,N_2736);
and U7603 (N_7603,N_2569,N_783);
or U7604 (N_7604,N_4007,N_1823);
nand U7605 (N_7605,N_2579,N_3667);
xnor U7606 (N_7606,N_3837,N_2289);
nand U7607 (N_7607,N_2610,N_2089);
and U7608 (N_7608,N_4012,N_860);
nand U7609 (N_7609,N_1465,N_3926);
xnor U7610 (N_7610,N_492,N_1576);
nand U7611 (N_7611,N_1053,N_2315);
nor U7612 (N_7612,N_4069,N_186);
nand U7613 (N_7613,N_3606,N_2119);
and U7614 (N_7614,N_1229,N_838);
nand U7615 (N_7615,N_3311,N_4482);
nor U7616 (N_7616,N_1332,N_3682);
xor U7617 (N_7617,N_2726,N_3893);
or U7618 (N_7618,N_889,N_3673);
nand U7619 (N_7619,N_1655,N_3946);
xnor U7620 (N_7620,N_3484,N_4061);
nor U7621 (N_7621,N_1646,N_799);
and U7622 (N_7622,N_3291,N_4361);
and U7623 (N_7623,N_2269,N_1917);
and U7624 (N_7624,N_2498,N_1131);
or U7625 (N_7625,N_4589,N_190);
nor U7626 (N_7626,N_912,N_424);
and U7627 (N_7627,N_3923,N_4163);
nand U7628 (N_7628,N_3865,N_2740);
nand U7629 (N_7629,N_1287,N_2507);
and U7630 (N_7630,N_3401,N_4701);
nor U7631 (N_7631,N_3887,N_2974);
nand U7632 (N_7632,N_4394,N_2370);
and U7633 (N_7633,N_3999,N_4846);
nor U7634 (N_7634,N_4211,N_3572);
or U7635 (N_7635,N_1859,N_177);
nand U7636 (N_7636,N_1312,N_1828);
nand U7637 (N_7637,N_96,N_1012);
and U7638 (N_7638,N_971,N_4646);
nand U7639 (N_7639,N_1731,N_508);
nand U7640 (N_7640,N_4873,N_3727);
and U7641 (N_7641,N_2880,N_4);
nand U7642 (N_7642,N_3164,N_1485);
or U7643 (N_7643,N_1616,N_183);
nand U7644 (N_7644,N_4086,N_321);
or U7645 (N_7645,N_1428,N_3072);
and U7646 (N_7646,N_3844,N_1971);
and U7647 (N_7647,N_1717,N_4221);
nand U7648 (N_7648,N_4372,N_2373);
and U7649 (N_7649,N_1141,N_33);
xor U7650 (N_7650,N_448,N_998);
and U7651 (N_7651,N_2534,N_2460);
or U7652 (N_7652,N_1466,N_2488);
or U7653 (N_7653,N_1692,N_3328);
or U7654 (N_7654,N_1363,N_1326);
or U7655 (N_7655,N_2438,N_2210);
nor U7656 (N_7656,N_4592,N_1722);
nor U7657 (N_7657,N_1868,N_341);
nor U7658 (N_7658,N_697,N_3644);
nor U7659 (N_7659,N_1826,N_3276);
nor U7660 (N_7660,N_3852,N_1495);
and U7661 (N_7661,N_4085,N_450);
and U7662 (N_7662,N_3925,N_789);
or U7663 (N_7663,N_4221,N_373);
or U7664 (N_7664,N_2235,N_5);
and U7665 (N_7665,N_3916,N_4154);
nand U7666 (N_7666,N_4355,N_1082);
nand U7667 (N_7667,N_4897,N_163);
or U7668 (N_7668,N_848,N_4307);
xnor U7669 (N_7669,N_2281,N_2293);
and U7670 (N_7670,N_395,N_4939);
xnor U7671 (N_7671,N_109,N_2904);
nor U7672 (N_7672,N_2233,N_1096);
nand U7673 (N_7673,N_4028,N_915);
nor U7674 (N_7674,N_2892,N_1774);
nor U7675 (N_7675,N_614,N_2805);
nand U7676 (N_7676,N_2728,N_200);
or U7677 (N_7677,N_711,N_910);
xor U7678 (N_7678,N_1779,N_1445);
and U7679 (N_7679,N_2071,N_3592);
xor U7680 (N_7680,N_1365,N_2251);
nand U7681 (N_7681,N_4529,N_3627);
nor U7682 (N_7682,N_2042,N_4061);
nand U7683 (N_7683,N_146,N_4479);
or U7684 (N_7684,N_3965,N_3061);
nand U7685 (N_7685,N_1512,N_1500);
nor U7686 (N_7686,N_4016,N_1116);
or U7687 (N_7687,N_1629,N_4823);
or U7688 (N_7688,N_4202,N_4504);
nand U7689 (N_7689,N_1815,N_4267);
nand U7690 (N_7690,N_1955,N_4044);
or U7691 (N_7691,N_458,N_3138);
xnor U7692 (N_7692,N_2504,N_1505);
or U7693 (N_7693,N_922,N_2089);
or U7694 (N_7694,N_1480,N_4047);
nor U7695 (N_7695,N_4774,N_3041);
or U7696 (N_7696,N_642,N_4903);
nand U7697 (N_7697,N_2592,N_1999);
and U7698 (N_7698,N_4414,N_2758);
and U7699 (N_7699,N_2895,N_2262);
and U7700 (N_7700,N_2947,N_4664);
and U7701 (N_7701,N_2373,N_2152);
nor U7702 (N_7702,N_4637,N_2118);
nor U7703 (N_7703,N_4365,N_2659);
nand U7704 (N_7704,N_1193,N_3083);
or U7705 (N_7705,N_865,N_1407);
nor U7706 (N_7706,N_4475,N_2597);
or U7707 (N_7707,N_1017,N_4154);
or U7708 (N_7708,N_2163,N_4546);
nor U7709 (N_7709,N_840,N_329);
nor U7710 (N_7710,N_669,N_3465);
xor U7711 (N_7711,N_2832,N_1049);
or U7712 (N_7712,N_3235,N_3453);
nor U7713 (N_7713,N_1500,N_4917);
or U7714 (N_7714,N_1726,N_3503);
and U7715 (N_7715,N_4407,N_2260);
nand U7716 (N_7716,N_1403,N_17);
nand U7717 (N_7717,N_2159,N_828);
or U7718 (N_7718,N_2240,N_2329);
nand U7719 (N_7719,N_399,N_4242);
nand U7720 (N_7720,N_4751,N_1575);
and U7721 (N_7721,N_4112,N_1297);
nand U7722 (N_7722,N_361,N_3059);
and U7723 (N_7723,N_3760,N_1313);
or U7724 (N_7724,N_3041,N_70);
nor U7725 (N_7725,N_578,N_4602);
xor U7726 (N_7726,N_3419,N_2735);
nand U7727 (N_7727,N_381,N_2022);
nand U7728 (N_7728,N_658,N_4957);
and U7729 (N_7729,N_1315,N_4620);
nor U7730 (N_7730,N_2184,N_3213);
or U7731 (N_7731,N_3283,N_727);
xnor U7732 (N_7732,N_550,N_911);
and U7733 (N_7733,N_2782,N_3385);
nand U7734 (N_7734,N_2208,N_3391);
nor U7735 (N_7735,N_2451,N_1886);
xor U7736 (N_7736,N_4509,N_2360);
or U7737 (N_7737,N_3285,N_2260);
nand U7738 (N_7738,N_3370,N_4085);
nor U7739 (N_7739,N_824,N_1648);
nand U7740 (N_7740,N_3987,N_4343);
xnor U7741 (N_7741,N_4379,N_307);
nor U7742 (N_7742,N_2871,N_3216);
and U7743 (N_7743,N_1609,N_2871);
xor U7744 (N_7744,N_3066,N_3852);
nor U7745 (N_7745,N_4179,N_3811);
xor U7746 (N_7746,N_3097,N_1663);
and U7747 (N_7747,N_3560,N_1899);
and U7748 (N_7748,N_4239,N_4663);
and U7749 (N_7749,N_1898,N_3561);
nand U7750 (N_7750,N_1730,N_3765);
or U7751 (N_7751,N_2097,N_2626);
or U7752 (N_7752,N_3619,N_1433);
xor U7753 (N_7753,N_3631,N_2839);
nand U7754 (N_7754,N_238,N_3025);
or U7755 (N_7755,N_3628,N_3823);
or U7756 (N_7756,N_1641,N_4695);
nand U7757 (N_7757,N_3531,N_2919);
nor U7758 (N_7758,N_1737,N_4951);
or U7759 (N_7759,N_4307,N_3290);
and U7760 (N_7760,N_917,N_2087);
nand U7761 (N_7761,N_1816,N_3408);
nor U7762 (N_7762,N_1922,N_3376);
and U7763 (N_7763,N_2293,N_644);
xor U7764 (N_7764,N_2732,N_4379);
and U7765 (N_7765,N_4683,N_2776);
xnor U7766 (N_7766,N_1478,N_3241);
xor U7767 (N_7767,N_2943,N_130);
or U7768 (N_7768,N_4930,N_3506);
and U7769 (N_7769,N_1040,N_4677);
and U7770 (N_7770,N_4077,N_4589);
nor U7771 (N_7771,N_3990,N_1685);
and U7772 (N_7772,N_1263,N_4418);
nand U7773 (N_7773,N_2363,N_2297);
xnor U7774 (N_7774,N_4906,N_1401);
nor U7775 (N_7775,N_3323,N_2056);
or U7776 (N_7776,N_4092,N_1898);
or U7777 (N_7777,N_2250,N_4566);
or U7778 (N_7778,N_1471,N_4094);
or U7779 (N_7779,N_2082,N_864);
or U7780 (N_7780,N_3890,N_3291);
nor U7781 (N_7781,N_3941,N_3926);
nor U7782 (N_7782,N_1510,N_1352);
xnor U7783 (N_7783,N_3055,N_3393);
or U7784 (N_7784,N_1973,N_177);
xnor U7785 (N_7785,N_3986,N_4383);
nand U7786 (N_7786,N_1373,N_1017);
xor U7787 (N_7787,N_3928,N_4155);
xor U7788 (N_7788,N_567,N_2660);
nand U7789 (N_7789,N_1031,N_2247);
nand U7790 (N_7790,N_4051,N_573);
nand U7791 (N_7791,N_718,N_4470);
nand U7792 (N_7792,N_822,N_2310);
xor U7793 (N_7793,N_929,N_357);
or U7794 (N_7794,N_4522,N_3219);
and U7795 (N_7795,N_902,N_4150);
or U7796 (N_7796,N_2402,N_2529);
or U7797 (N_7797,N_158,N_1626);
nor U7798 (N_7798,N_2672,N_3984);
nor U7799 (N_7799,N_3663,N_1925);
and U7800 (N_7800,N_897,N_2124);
or U7801 (N_7801,N_1133,N_3268);
and U7802 (N_7802,N_1071,N_3149);
and U7803 (N_7803,N_4732,N_2582);
nor U7804 (N_7804,N_419,N_750);
nand U7805 (N_7805,N_569,N_267);
nor U7806 (N_7806,N_4864,N_1906);
xnor U7807 (N_7807,N_2577,N_1741);
or U7808 (N_7808,N_1104,N_1578);
nand U7809 (N_7809,N_653,N_1984);
and U7810 (N_7810,N_2156,N_4928);
nand U7811 (N_7811,N_1533,N_4223);
or U7812 (N_7812,N_532,N_500);
nor U7813 (N_7813,N_1010,N_1504);
xnor U7814 (N_7814,N_3782,N_655);
and U7815 (N_7815,N_2225,N_4497);
and U7816 (N_7816,N_4457,N_1560);
nor U7817 (N_7817,N_4188,N_216);
nand U7818 (N_7818,N_3867,N_2136);
or U7819 (N_7819,N_2552,N_2302);
nand U7820 (N_7820,N_1235,N_1295);
nor U7821 (N_7821,N_4882,N_804);
nor U7822 (N_7822,N_2073,N_4874);
nor U7823 (N_7823,N_2992,N_1992);
xnor U7824 (N_7824,N_2451,N_1821);
nand U7825 (N_7825,N_1423,N_3869);
or U7826 (N_7826,N_978,N_2756);
or U7827 (N_7827,N_2709,N_755);
nand U7828 (N_7828,N_4056,N_3475);
nor U7829 (N_7829,N_4837,N_2474);
nor U7830 (N_7830,N_4257,N_2681);
nand U7831 (N_7831,N_117,N_2464);
and U7832 (N_7832,N_1319,N_4433);
and U7833 (N_7833,N_2678,N_4990);
xor U7834 (N_7834,N_858,N_2716);
nor U7835 (N_7835,N_3628,N_1013);
nand U7836 (N_7836,N_574,N_3204);
and U7837 (N_7837,N_849,N_3199);
xnor U7838 (N_7838,N_2535,N_14);
xnor U7839 (N_7839,N_1319,N_4772);
nand U7840 (N_7840,N_2138,N_3783);
xnor U7841 (N_7841,N_2772,N_854);
nor U7842 (N_7842,N_4958,N_2409);
nor U7843 (N_7843,N_2844,N_2966);
nand U7844 (N_7844,N_3746,N_2264);
xor U7845 (N_7845,N_510,N_3446);
and U7846 (N_7846,N_2325,N_2937);
and U7847 (N_7847,N_768,N_1284);
nor U7848 (N_7848,N_3341,N_4345);
nor U7849 (N_7849,N_2258,N_3572);
nand U7850 (N_7850,N_3239,N_220);
nand U7851 (N_7851,N_1666,N_3621);
xnor U7852 (N_7852,N_4704,N_2955);
and U7853 (N_7853,N_2683,N_3212);
xor U7854 (N_7854,N_2564,N_4787);
nor U7855 (N_7855,N_171,N_4598);
and U7856 (N_7856,N_1148,N_4895);
nor U7857 (N_7857,N_68,N_2090);
or U7858 (N_7858,N_4950,N_118);
xnor U7859 (N_7859,N_4928,N_1616);
nor U7860 (N_7860,N_19,N_3130);
and U7861 (N_7861,N_713,N_4973);
nor U7862 (N_7862,N_2880,N_3140);
nand U7863 (N_7863,N_1304,N_4778);
xor U7864 (N_7864,N_817,N_3271);
nand U7865 (N_7865,N_3209,N_170);
nor U7866 (N_7866,N_4740,N_2155);
or U7867 (N_7867,N_243,N_540);
nor U7868 (N_7868,N_4452,N_234);
nor U7869 (N_7869,N_1842,N_276);
nand U7870 (N_7870,N_2330,N_328);
and U7871 (N_7871,N_1600,N_1363);
and U7872 (N_7872,N_1345,N_2592);
nand U7873 (N_7873,N_4241,N_1015);
nand U7874 (N_7874,N_3251,N_2180);
and U7875 (N_7875,N_1443,N_66);
or U7876 (N_7876,N_1853,N_2380);
or U7877 (N_7877,N_3991,N_251);
or U7878 (N_7878,N_78,N_309);
or U7879 (N_7879,N_1810,N_1132);
or U7880 (N_7880,N_1406,N_4849);
and U7881 (N_7881,N_1672,N_3226);
nor U7882 (N_7882,N_991,N_3406);
nand U7883 (N_7883,N_4233,N_974);
nand U7884 (N_7884,N_1311,N_1694);
xor U7885 (N_7885,N_1946,N_3787);
nand U7886 (N_7886,N_2475,N_3978);
or U7887 (N_7887,N_949,N_4902);
or U7888 (N_7888,N_1626,N_2068);
nor U7889 (N_7889,N_4089,N_4762);
or U7890 (N_7890,N_4200,N_1501);
and U7891 (N_7891,N_3624,N_4100);
xnor U7892 (N_7892,N_411,N_2546);
or U7893 (N_7893,N_486,N_1247);
nor U7894 (N_7894,N_319,N_1966);
or U7895 (N_7895,N_1217,N_4473);
nand U7896 (N_7896,N_4279,N_1248);
nand U7897 (N_7897,N_4828,N_2538);
xnor U7898 (N_7898,N_1342,N_4713);
nor U7899 (N_7899,N_1557,N_4284);
and U7900 (N_7900,N_2607,N_1255);
nand U7901 (N_7901,N_4888,N_1129);
or U7902 (N_7902,N_217,N_1481);
and U7903 (N_7903,N_3662,N_1540);
and U7904 (N_7904,N_4528,N_4691);
and U7905 (N_7905,N_1230,N_3136);
and U7906 (N_7906,N_3343,N_3102);
nand U7907 (N_7907,N_2281,N_4088);
xor U7908 (N_7908,N_316,N_4197);
or U7909 (N_7909,N_3049,N_3640);
and U7910 (N_7910,N_944,N_2168);
nor U7911 (N_7911,N_1243,N_1387);
and U7912 (N_7912,N_4781,N_4904);
and U7913 (N_7913,N_1778,N_79);
and U7914 (N_7914,N_728,N_1683);
and U7915 (N_7915,N_4850,N_4530);
nor U7916 (N_7916,N_1190,N_4858);
nand U7917 (N_7917,N_1899,N_1618);
nor U7918 (N_7918,N_1435,N_2662);
and U7919 (N_7919,N_366,N_2717);
and U7920 (N_7920,N_1150,N_4691);
and U7921 (N_7921,N_2177,N_4320);
nand U7922 (N_7922,N_4820,N_3254);
and U7923 (N_7923,N_1606,N_629);
xor U7924 (N_7924,N_1535,N_2161);
xor U7925 (N_7925,N_771,N_3703);
nand U7926 (N_7926,N_1869,N_1862);
nand U7927 (N_7927,N_1663,N_3296);
xnor U7928 (N_7928,N_3555,N_4700);
or U7929 (N_7929,N_2494,N_4795);
and U7930 (N_7930,N_1291,N_3360);
or U7931 (N_7931,N_3634,N_893);
and U7932 (N_7932,N_2003,N_2492);
nand U7933 (N_7933,N_896,N_4268);
nor U7934 (N_7934,N_637,N_3094);
xor U7935 (N_7935,N_3926,N_801);
or U7936 (N_7936,N_96,N_368);
or U7937 (N_7937,N_1940,N_1612);
or U7938 (N_7938,N_1532,N_4720);
nand U7939 (N_7939,N_2924,N_3504);
nand U7940 (N_7940,N_272,N_2725);
nor U7941 (N_7941,N_86,N_2334);
and U7942 (N_7942,N_4937,N_4519);
or U7943 (N_7943,N_4898,N_3713);
or U7944 (N_7944,N_3686,N_165);
xnor U7945 (N_7945,N_2498,N_1892);
nor U7946 (N_7946,N_3151,N_2219);
and U7947 (N_7947,N_907,N_4859);
and U7948 (N_7948,N_4661,N_4217);
or U7949 (N_7949,N_1557,N_2552);
and U7950 (N_7950,N_3426,N_91);
nand U7951 (N_7951,N_447,N_949);
nor U7952 (N_7952,N_3419,N_2483);
or U7953 (N_7953,N_3671,N_592);
and U7954 (N_7954,N_3993,N_3626);
or U7955 (N_7955,N_4836,N_3970);
nor U7956 (N_7956,N_2974,N_4916);
nor U7957 (N_7957,N_3057,N_3958);
nor U7958 (N_7958,N_4097,N_3140);
xnor U7959 (N_7959,N_4963,N_4700);
xor U7960 (N_7960,N_3245,N_4242);
and U7961 (N_7961,N_4543,N_1837);
nor U7962 (N_7962,N_1137,N_2478);
or U7963 (N_7963,N_2293,N_4534);
or U7964 (N_7964,N_1639,N_1047);
and U7965 (N_7965,N_3781,N_1866);
nor U7966 (N_7966,N_3673,N_1693);
xor U7967 (N_7967,N_2442,N_2214);
nand U7968 (N_7968,N_2033,N_4050);
or U7969 (N_7969,N_1381,N_3686);
nor U7970 (N_7970,N_3744,N_196);
nor U7971 (N_7971,N_251,N_66);
nor U7972 (N_7972,N_4385,N_2022);
nor U7973 (N_7973,N_3559,N_4477);
nand U7974 (N_7974,N_1386,N_3759);
or U7975 (N_7975,N_3515,N_1665);
and U7976 (N_7976,N_381,N_1986);
or U7977 (N_7977,N_66,N_2500);
or U7978 (N_7978,N_430,N_1673);
and U7979 (N_7979,N_4460,N_3091);
and U7980 (N_7980,N_3958,N_2090);
and U7981 (N_7981,N_2453,N_865);
or U7982 (N_7982,N_2626,N_4487);
and U7983 (N_7983,N_1935,N_4712);
and U7984 (N_7984,N_4511,N_2824);
or U7985 (N_7985,N_1844,N_3041);
and U7986 (N_7986,N_306,N_367);
or U7987 (N_7987,N_4831,N_1395);
nand U7988 (N_7988,N_652,N_4125);
or U7989 (N_7989,N_2424,N_3884);
nand U7990 (N_7990,N_3644,N_4640);
nand U7991 (N_7991,N_2560,N_2562);
or U7992 (N_7992,N_1118,N_1732);
nor U7993 (N_7993,N_1721,N_3311);
nor U7994 (N_7994,N_3987,N_3768);
nor U7995 (N_7995,N_3395,N_1249);
nand U7996 (N_7996,N_3779,N_1725);
nand U7997 (N_7997,N_978,N_1648);
nand U7998 (N_7998,N_2986,N_1725);
nor U7999 (N_7999,N_4711,N_4085);
nor U8000 (N_8000,N_4811,N_3196);
nand U8001 (N_8001,N_3708,N_2224);
nor U8002 (N_8002,N_959,N_2878);
or U8003 (N_8003,N_1460,N_4426);
nand U8004 (N_8004,N_3468,N_3700);
xor U8005 (N_8005,N_2335,N_2714);
nand U8006 (N_8006,N_3644,N_1234);
nor U8007 (N_8007,N_3252,N_4342);
and U8008 (N_8008,N_2855,N_1560);
or U8009 (N_8009,N_123,N_4128);
and U8010 (N_8010,N_2166,N_2199);
xor U8011 (N_8011,N_2440,N_3879);
nand U8012 (N_8012,N_2554,N_2740);
nand U8013 (N_8013,N_3614,N_1584);
nor U8014 (N_8014,N_2269,N_652);
xor U8015 (N_8015,N_3910,N_1213);
or U8016 (N_8016,N_3137,N_3111);
xnor U8017 (N_8017,N_2765,N_3915);
nor U8018 (N_8018,N_1144,N_1202);
nand U8019 (N_8019,N_3395,N_3777);
xnor U8020 (N_8020,N_3773,N_1113);
xor U8021 (N_8021,N_2503,N_4379);
nor U8022 (N_8022,N_3286,N_1263);
or U8023 (N_8023,N_4286,N_4847);
nand U8024 (N_8024,N_3201,N_739);
and U8025 (N_8025,N_1126,N_1756);
and U8026 (N_8026,N_1619,N_3306);
nand U8027 (N_8027,N_2858,N_3738);
nand U8028 (N_8028,N_3964,N_726);
or U8029 (N_8029,N_2701,N_4650);
nor U8030 (N_8030,N_4825,N_3760);
nand U8031 (N_8031,N_2205,N_1509);
nand U8032 (N_8032,N_829,N_2769);
nor U8033 (N_8033,N_3575,N_13);
nor U8034 (N_8034,N_4186,N_446);
nor U8035 (N_8035,N_3581,N_4333);
nor U8036 (N_8036,N_1303,N_2943);
and U8037 (N_8037,N_273,N_277);
nor U8038 (N_8038,N_900,N_356);
nor U8039 (N_8039,N_1610,N_2644);
nor U8040 (N_8040,N_4926,N_2514);
or U8041 (N_8041,N_3368,N_1716);
nand U8042 (N_8042,N_4346,N_3397);
and U8043 (N_8043,N_2607,N_1992);
or U8044 (N_8044,N_1657,N_4212);
xor U8045 (N_8045,N_3762,N_4668);
nor U8046 (N_8046,N_1889,N_2596);
xor U8047 (N_8047,N_4415,N_4175);
xor U8048 (N_8048,N_709,N_846);
nand U8049 (N_8049,N_504,N_2860);
and U8050 (N_8050,N_1505,N_4046);
xor U8051 (N_8051,N_3031,N_2154);
or U8052 (N_8052,N_2023,N_2520);
nor U8053 (N_8053,N_1383,N_2433);
or U8054 (N_8054,N_4440,N_2028);
nand U8055 (N_8055,N_528,N_1574);
nor U8056 (N_8056,N_3353,N_475);
nand U8057 (N_8057,N_3766,N_4103);
nand U8058 (N_8058,N_3805,N_4158);
and U8059 (N_8059,N_397,N_3333);
or U8060 (N_8060,N_4156,N_1808);
or U8061 (N_8061,N_2346,N_27);
or U8062 (N_8062,N_4281,N_2437);
nor U8063 (N_8063,N_2909,N_4600);
xnor U8064 (N_8064,N_1785,N_3275);
and U8065 (N_8065,N_2979,N_2224);
or U8066 (N_8066,N_2094,N_128);
nand U8067 (N_8067,N_3291,N_87);
and U8068 (N_8068,N_2373,N_4585);
or U8069 (N_8069,N_3372,N_4040);
nand U8070 (N_8070,N_2533,N_4249);
and U8071 (N_8071,N_1272,N_3434);
nand U8072 (N_8072,N_150,N_4577);
and U8073 (N_8073,N_2941,N_634);
nor U8074 (N_8074,N_685,N_2072);
xor U8075 (N_8075,N_1516,N_3831);
or U8076 (N_8076,N_3580,N_3036);
nand U8077 (N_8077,N_1895,N_122);
nand U8078 (N_8078,N_2359,N_929);
nor U8079 (N_8079,N_3042,N_3558);
or U8080 (N_8080,N_2525,N_2287);
nor U8081 (N_8081,N_3626,N_561);
xor U8082 (N_8082,N_4153,N_1442);
xor U8083 (N_8083,N_3455,N_4515);
or U8084 (N_8084,N_3384,N_142);
xor U8085 (N_8085,N_3415,N_3428);
xor U8086 (N_8086,N_2565,N_426);
xor U8087 (N_8087,N_4966,N_438);
nand U8088 (N_8088,N_4400,N_2806);
and U8089 (N_8089,N_4582,N_4703);
nor U8090 (N_8090,N_900,N_4548);
nor U8091 (N_8091,N_1782,N_4865);
and U8092 (N_8092,N_1210,N_2222);
nand U8093 (N_8093,N_876,N_1402);
and U8094 (N_8094,N_972,N_3753);
nor U8095 (N_8095,N_3307,N_1327);
and U8096 (N_8096,N_3065,N_2599);
nand U8097 (N_8097,N_1600,N_4772);
nand U8098 (N_8098,N_2085,N_2413);
nor U8099 (N_8099,N_3937,N_4426);
and U8100 (N_8100,N_1292,N_4012);
xor U8101 (N_8101,N_1312,N_3463);
nor U8102 (N_8102,N_4136,N_4455);
nor U8103 (N_8103,N_4782,N_2675);
and U8104 (N_8104,N_1597,N_2799);
nor U8105 (N_8105,N_2741,N_3077);
nor U8106 (N_8106,N_4976,N_1572);
or U8107 (N_8107,N_1625,N_1536);
or U8108 (N_8108,N_2282,N_2040);
or U8109 (N_8109,N_2014,N_4397);
nor U8110 (N_8110,N_2988,N_2561);
or U8111 (N_8111,N_4017,N_2576);
and U8112 (N_8112,N_1251,N_3292);
nand U8113 (N_8113,N_249,N_1963);
and U8114 (N_8114,N_2999,N_70);
nand U8115 (N_8115,N_853,N_1439);
xnor U8116 (N_8116,N_3031,N_4875);
or U8117 (N_8117,N_3423,N_1045);
or U8118 (N_8118,N_1105,N_3097);
or U8119 (N_8119,N_4946,N_1347);
nand U8120 (N_8120,N_2005,N_2417);
xor U8121 (N_8121,N_2302,N_1169);
or U8122 (N_8122,N_1538,N_890);
nand U8123 (N_8123,N_4520,N_528);
nand U8124 (N_8124,N_1403,N_2215);
xnor U8125 (N_8125,N_4,N_468);
nor U8126 (N_8126,N_2021,N_4093);
or U8127 (N_8127,N_3665,N_3843);
nand U8128 (N_8128,N_2527,N_1663);
nand U8129 (N_8129,N_1160,N_2327);
or U8130 (N_8130,N_4102,N_3300);
nor U8131 (N_8131,N_3894,N_3035);
or U8132 (N_8132,N_1339,N_1354);
nor U8133 (N_8133,N_384,N_2014);
xnor U8134 (N_8134,N_1019,N_33);
or U8135 (N_8135,N_4526,N_4604);
xor U8136 (N_8136,N_695,N_3207);
or U8137 (N_8137,N_1364,N_1227);
xor U8138 (N_8138,N_708,N_4479);
and U8139 (N_8139,N_2663,N_2419);
or U8140 (N_8140,N_955,N_1312);
and U8141 (N_8141,N_1555,N_2251);
or U8142 (N_8142,N_2123,N_1427);
or U8143 (N_8143,N_3883,N_4964);
xor U8144 (N_8144,N_3008,N_3725);
nor U8145 (N_8145,N_80,N_227);
nand U8146 (N_8146,N_3385,N_2042);
or U8147 (N_8147,N_4682,N_3690);
nor U8148 (N_8148,N_4751,N_4357);
and U8149 (N_8149,N_3361,N_1263);
nand U8150 (N_8150,N_3167,N_4620);
and U8151 (N_8151,N_972,N_2812);
nor U8152 (N_8152,N_1032,N_2519);
nor U8153 (N_8153,N_74,N_3873);
or U8154 (N_8154,N_4930,N_891);
nor U8155 (N_8155,N_1743,N_3766);
and U8156 (N_8156,N_4395,N_396);
nor U8157 (N_8157,N_4869,N_106);
nor U8158 (N_8158,N_3149,N_2421);
and U8159 (N_8159,N_610,N_3334);
or U8160 (N_8160,N_2979,N_665);
xnor U8161 (N_8161,N_1653,N_3133);
nand U8162 (N_8162,N_3194,N_287);
xnor U8163 (N_8163,N_3374,N_614);
nor U8164 (N_8164,N_4709,N_3645);
or U8165 (N_8165,N_753,N_1719);
and U8166 (N_8166,N_103,N_3542);
and U8167 (N_8167,N_3798,N_3310);
nand U8168 (N_8168,N_130,N_3512);
or U8169 (N_8169,N_472,N_2333);
and U8170 (N_8170,N_2619,N_2193);
nand U8171 (N_8171,N_4448,N_1585);
nand U8172 (N_8172,N_1836,N_436);
or U8173 (N_8173,N_2206,N_2085);
nand U8174 (N_8174,N_4580,N_2159);
and U8175 (N_8175,N_4271,N_1093);
and U8176 (N_8176,N_2853,N_4211);
and U8177 (N_8177,N_3289,N_3286);
nor U8178 (N_8178,N_2035,N_4762);
or U8179 (N_8179,N_3448,N_1386);
or U8180 (N_8180,N_763,N_2549);
and U8181 (N_8181,N_220,N_575);
nor U8182 (N_8182,N_3737,N_50);
nor U8183 (N_8183,N_4166,N_3716);
nor U8184 (N_8184,N_4283,N_4332);
xnor U8185 (N_8185,N_2574,N_2792);
or U8186 (N_8186,N_755,N_3105);
nand U8187 (N_8187,N_4518,N_4801);
nor U8188 (N_8188,N_1880,N_1223);
nor U8189 (N_8189,N_3424,N_232);
and U8190 (N_8190,N_3856,N_413);
and U8191 (N_8191,N_4328,N_1672);
nor U8192 (N_8192,N_4861,N_2292);
nor U8193 (N_8193,N_1076,N_4685);
nand U8194 (N_8194,N_3230,N_1609);
nand U8195 (N_8195,N_2304,N_4294);
nor U8196 (N_8196,N_3636,N_1916);
nand U8197 (N_8197,N_4257,N_1215);
nand U8198 (N_8198,N_531,N_4009);
xor U8199 (N_8199,N_3462,N_3350);
nor U8200 (N_8200,N_3459,N_1601);
xnor U8201 (N_8201,N_4590,N_4200);
nand U8202 (N_8202,N_4838,N_387);
nand U8203 (N_8203,N_3795,N_487);
and U8204 (N_8204,N_3191,N_3282);
nor U8205 (N_8205,N_2976,N_553);
nand U8206 (N_8206,N_4503,N_4318);
nor U8207 (N_8207,N_3972,N_3894);
and U8208 (N_8208,N_2487,N_830);
nand U8209 (N_8209,N_791,N_4658);
and U8210 (N_8210,N_2110,N_3355);
or U8211 (N_8211,N_1702,N_367);
nor U8212 (N_8212,N_3845,N_3628);
nor U8213 (N_8213,N_3401,N_2918);
or U8214 (N_8214,N_3380,N_207);
nand U8215 (N_8215,N_4927,N_4959);
nor U8216 (N_8216,N_3540,N_3642);
nand U8217 (N_8217,N_1789,N_4980);
and U8218 (N_8218,N_2547,N_3427);
and U8219 (N_8219,N_4052,N_2195);
nor U8220 (N_8220,N_2433,N_1482);
nor U8221 (N_8221,N_480,N_4211);
and U8222 (N_8222,N_465,N_3271);
nand U8223 (N_8223,N_1365,N_1348);
xnor U8224 (N_8224,N_1398,N_1281);
or U8225 (N_8225,N_996,N_1077);
xnor U8226 (N_8226,N_1084,N_3892);
nand U8227 (N_8227,N_1221,N_4826);
nand U8228 (N_8228,N_3397,N_4650);
nor U8229 (N_8229,N_802,N_2952);
nor U8230 (N_8230,N_3269,N_4511);
xnor U8231 (N_8231,N_2416,N_1398);
and U8232 (N_8232,N_4668,N_4451);
nor U8233 (N_8233,N_1310,N_3523);
nor U8234 (N_8234,N_592,N_1143);
nand U8235 (N_8235,N_3447,N_138);
and U8236 (N_8236,N_2814,N_4110);
or U8237 (N_8237,N_253,N_4743);
nand U8238 (N_8238,N_4850,N_540);
nand U8239 (N_8239,N_2365,N_2887);
and U8240 (N_8240,N_2932,N_439);
nand U8241 (N_8241,N_3387,N_3749);
nor U8242 (N_8242,N_1876,N_797);
nor U8243 (N_8243,N_153,N_3008);
nor U8244 (N_8244,N_3063,N_2208);
and U8245 (N_8245,N_1482,N_1624);
nand U8246 (N_8246,N_2395,N_3931);
or U8247 (N_8247,N_4018,N_2060);
nand U8248 (N_8248,N_2870,N_1806);
nand U8249 (N_8249,N_3805,N_4044);
xnor U8250 (N_8250,N_827,N_2337);
nand U8251 (N_8251,N_3846,N_3183);
and U8252 (N_8252,N_4365,N_2136);
nand U8253 (N_8253,N_4621,N_628);
and U8254 (N_8254,N_1301,N_1847);
and U8255 (N_8255,N_1516,N_3788);
or U8256 (N_8256,N_4261,N_2070);
and U8257 (N_8257,N_1740,N_3210);
nand U8258 (N_8258,N_3418,N_502);
nand U8259 (N_8259,N_4864,N_1112);
or U8260 (N_8260,N_1529,N_4867);
nand U8261 (N_8261,N_4177,N_4683);
and U8262 (N_8262,N_4289,N_2493);
and U8263 (N_8263,N_193,N_1962);
nor U8264 (N_8264,N_4780,N_3783);
or U8265 (N_8265,N_482,N_3088);
and U8266 (N_8266,N_213,N_4514);
and U8267 (N_8267,N_3049,N_951);
nor U8268 (N_8268,N_4143,N_1457);
xnor U8269 (N_8269,N_3472,N_2151);
nor U8270 (N_8270,N_598,N_173);
or U8271 (N_8271,N_3099,N_177);
xnor U8272 (N_8272,N_3312,N_2856);
and U8273 (N_8273,N_2750,N_3700);
nor U8274 (N_8274,N_4293,N_1473);
or U8275 (N_8275,N_2138,N_3401);
nor U8276 (N_8276,N_1276,N_3275);
nand U8277 (N_8277,N_1640,N_1627);
nor U8278 (N_8278,N_1192,N_2543);
nor U8279 (N_8279,N_2023,N_2422);
and U8280 (N_8280,N_2140,N_222);
nand U8281 (N_8281,N_2739,N_270);
or U8282 (N_8282,N_629,N_1462);
nand U8283 (N_8283,N_3094,N_1771);
xnor U8284 (N_8284,N_435,N_1970);
or U8285 (N_8285,N_4934,N_331);
nor U8286 (N_8286,N_3689,N_2350);
xnor U8287 (N_8287,N_1182,N_4120);
and U8288 (N_8288,N_3071,N_3861);
nand U8289 (N_8289,N_3032,N_2926);
and U8290 (N_8290,N_4591,N_847);
nor U8291 (N_8291,N_4389,N_2367);
and U8292 (N_8292,N_91,N_2941);
or U8293 (N_8293,N_3496,N_385);
nand U8294 (N_8294,N_1832,N_841);
and U8295 (N_8295,N_2321,N_4646);
nor U8296 (N_8296,N_1303,N_4531);
nor U8297 (N_8297,N_1573,N_1333);
and U8298 (N_8298,N_4887,N_4504);
xnor U8299 (N_8299,N_979,N_1700);
nor U8300 (N_8300,N_1876,N_4422);
and U8301 (N_8301,N_4995,N_4382);
nand U8302 (N_8302,N_671,N_2847);
and U8303 (N_8303,N_3340,N_2060);
xor U8304 (N_8304,N_1764,N_1737);
or U8305 (N_8305,N_3437,N_1046);
or U8306 (N_8306,N_3689,N_4420);
nor U8307 (N_8307,N_1478,N_4150);
and U8308 (N_8308,N_3707,N_4419);
or U8309 (N_8309,N_3011,N_3741);
or U8310 (N_8310,N_4445,N_4695);
or U8311 (N_8311,N_3238,N_1536);
nand U8312 (N_8312,N_804,N_1090);
or U8313 (N_8313,N_2625,N_1361);
nor U8314 (N_8314,N_2228,N_1445);
nand U8315 (N_8315,N_4801,N_2063);
or U8316 (N_8316,N_2470,N_701);
and U8317 (N_8317,N_3621,N_564);
and U8318 (N_8318,N_764,N_2498);
nand U8319 (N_8319,N_1060,N_1044);
nor U8320 (N_8320,N_730,N_1693);
nand U8321 (N_8321,N_2133,N_2775);
or U8322 (N_8322,N_330,N_4564);
nor U8323 (N_8323,N_4985,N_1449);
nor U8324 (N_8324,N_1119,N_1694);
and U8325 (N_8325,N_4031,N_3561);
nand U8326 (N_8326,N_4953,N_2013);
xnor U8327 (N_8327,N_4902,N_3113);
and U8328 (N_8328,N_3630,N_4067);
nand U8329 (N_8329,N_2550,N_1034);
nand U8330 (N_8330,N_1959,N_3989);
or U8331 (N_8331,N_3447,N_2275);
nor U8332 (N_8332,N_698,N_4516);
nor U8333 (N_8333,N_746,N_2621);
nor U8334 (N_8334,N_3337,N_687);
nand U8335 (N_8335,N_3049,N_4405);
nor U8336 (N_8336,N_88,N_300);
nand U8337 (N_8337,N_4170,N_3502);
or U8338 (N_8338,N_466,N_1682);
or U8339 (N_8339,N_2958,N_1321);
and U8340 (N_8340,N_19,N_4661);
nand U8341 (N_8341,N_2980,N_4218);
or U8342 (N_8342,N_3112,N_3394);
nand U8343 (N_8343,N_1234,N_2413);
and U8344 (N_8344,N_1724,N_3635);
nand U8345 (N_8345,N_3839,N_1480);
or U8346 (N_8346,N_3712,N_3155);
nor U8347 (N_8347,N_2878,N_4067);
or U8348 (N_8348,N_3121,N_202);
or U8349 (N_8349,N_908,N_4380);
or U8350 (N_8350,N_4486,N_541);
and U8351 (N_8351,N_988,N_3740);
nor U8352 (N_8352,N_2560,N_1698);
and U8353 (N_8353,N_4642,N_4830);
nand U8354 (N_8354,N_3729,N_4649);
nor U8355 (N_8355,N_4879,N_3470);
nor U8356 (N_8356,N_4303,N_2573);
nand U8357 (N_8357,N_464,N_235);
and U8358 (N_8358,N_1594,N_2125);
xnor U8359 (N_8359,N_4049,N_2718);
nand U8360 (N_8360,N_2620,N_612);
nand U8361 (N_8361,N_4701,N_2546);
nand U8362 (N_8362,N_3562,N_136);
nor U8363 (N_8363,N_3527,N_104);
or U8364 (N_8364,N_2885,N_3928);
nand U8365 (N_8365,N_3786,N_1045);
and U8366 (N_8366,N_4485,N_88);
nor U8367 (N_8367,N_2267,N_3020);
nor U8368 (N_8368,N_755,N_2756);
nor U8369 (N_8369,N_915,N_1072);
nand U8370 (N_8370,N_3996,N_1507);
nor U8371 (N_8371,N_1022,N_1528);
and U8372 (N_8372,N_2415,N_1629);
nand U8373 (N_8373,N_1386,N_682);
nand U8374 (N_8374,N_2601,N_3726);
and U8375 (N_8375,N_1184,N_829);
and U8376 (N_8376,N_4532,N_2524);
xor U8377 (N_8377,N_393,N_2460);
or U8378 (N_8378,N_2166,N_2189);
or U8379 (N_8379,N_1836,N_2113);
or U8380 (N_8380,N_1324,N_4800);
nand U8381 (N_8381,N_3844,N_561);
nor U8382 (N_8382,N_3503,N_882);
and U8383 (N_8383,N_4212,N_3008);
and U8384 (N_8384,N_868,N_4179);
nor U8385 (N_8385,N_2377,N_279);
and U8386 (N_8386,N_2587,N_1363);
nand U8387 (N_8387,N_455,N_788);
nand U8388 (N_8388,N_3190,N_1231);
and U8389 (N_8389,N_2882,N_4352);
nand U8390 (N_8390,N_2236,N_1095);
nor U8391 (N_8391,N_2096,N_265);
nand U8392 (N_8392,N_1010,N_1906);
or U8393 (N_8393,N_518,N_3576);
and U8394 (N_8394,N_266,N_252);
xnor U8395 (N_8395,N_2836,N_4594);
or U8396 (N_8396,N_4992,N_172);
and U8397 (N_8397,N_2670,N_4572);
and U8398 (N_8398,N_1796,N_772);
nand U8399 (N_8399,N_4929,N_3358);
nor U8400 (N_8400,N_497,N_2564);
nor U8401 (N_8401,N_3853,N_3058);
and U8402 (N_8402,N_3622,N_4083);
or U8403 (N_8403,N_3676,N_2794);
nand U8404 (N_8404,N_3605,N_907);
xor U8405 (N_8405,N_1739,N_2129);
nand U8406 (N_8406,N_915,N_2725);
nand U8407 (N_8407,N_554,N_4117);
or U8408 (N_8408,N_905,N_4125);
or U8409 (N_8409,N_4343,N_299);
nor U8410 (N_8410,N_393,N_3311);
xnor U8411 (N_8411,N_2708,N_3088);
xor U8412 (N_8412,N_2837,N_3469);
and U8413 (N_8413,N_559,N_3451);
nand U8414 (N_8414,N_3515,N_2000);
xor U8415 (N_8415,N_3301,N_1301);
or U8416 (N_8416,N_3855,N_3188);
and U8417 (N_8417,N_4348,N_976);
nand U8418 (N_8418,N_8,N_420);
and U8419 (N_8419,N_4961,N_2943);
and U8420 (N_8420,N_2308,N_2412);
and U8421 (N_8421,N_254,N_4870);
nor U8422 (N_8422,N_2502,N_623);
or U8423 (N_8423,N_329,N_3549);
xnor U8424 (N_8424,N_4318,N_4591);
nand U8425 (N_8425,N_3122,N_4175);
and U8426 (N_8426,N_3470,N_3587);
and U8427 (N_8427,N_3812,N_2821);
and U8428 (N_8428,N_4187,N_3944);
nor U8429 (N_8429,N_3109,N_714);
nand U8430 (N_8430,N_2425,N_3493);
nand U8431 (N_8431,N_97,N_901);
nor U8432 (N_8432,N_2783,N_4093);
nand U8433 (N_8433,N_3196,N_3317);
or U8434 (N_8434,N_2625,N_2390);
nor U8435 (N_8435,N_2956,N_3841);
xnor U8436 (N_8436,N_3620,N_4762);
or U8437 (N_8437,N_4924,N_1188);
xnor U8438 (N_8438,N_3375,N_4394);
nand U8439 (N_8439,N_2284,N_4645);
and U8440 (N_8440,N_2471,N_568);
or U8441 (N_8441,N_2175,N_1736);
nand U8442 (N_8442,N_430,N_714);
nor U8443 (N_8443,N_591,N_920);
nand U8444 (N_8444,N_323,N_3347);
nor U8445 (N_8445,N_1497,N_441);
nand U8446 (N_8446,N_2360,N_4869);
and U8447 (N_8447,N_3790,N_3562);
nand U8448 (N_8448,N_1600,N_2183);
and U8449 (N_8449,N_1103,N_193);
xor U8450 (N_8450,N_2430,N_3915);
nor U8451 (N_8451,N_4869,N_2518);
xnor U8452 (N_8452,N_3734,N_1318);
and U8453 (N_8453,N_4651,N_1697);
nor U8454 (N_8454,N_1450,N_4802);
and U8455 (N_8455,N_517,N_4237);
nor U8456 (N_8456,N_3901,N_2479);
nor U8457 (N_8457,N_2961,N_4255);
nor U8458 (N_8458,N_2304,N_467);
or U8459 (N_8459,N_2809,N_4588);
nor U8460 (N_8460,N_3644,N_3943);
or U8461 (N_8461,N_2062,N_278);
and U8462 (N_8462,N_4000,N_3174);
and U8463 (N_8463,N_3688,N_253);
nor U8464 (N_8464,N_3824,N_1374);
and U8465 (N_8465,N_465,N_470);
or U8466 (N_8466,N_4254,N_463);
and U8467 (N_8467,N_1840,N_3912);
nand U8468 (N_8468,N_1096,N_3902);
nor U8469 (N_8469,N_1526,N_428);
nor U8470 (N_8470,N_554,N_1391);
or U8471 (N_8471,N_3654,N_3330);
nor U8472 (N_8472,N_4302,N_3917);
or U8473 (N_8473,N_3780,N_1678);
or U8474 (N_8474,N_2323,N_1914);
nor U8475 (N_8475,N_4873,N_2987);
nor U8476 (N_8476,N_1306,N_3384);
or U8477 (N_8477,N_579,N_2578);
and U8478 (N_8478,N_3347,N_3123);
nor U8479 (N_8479,N_1211,N_3632);
nor U8480 (N_8480,N_629,N_1433);
nor U8481 (N_8481,N_417,N_1166);
nor U8482 (N_8482,N_2738,N_3363);
or U8483 (N_8483,N_1568,N_954);
nand U8484 (N_8484,N_2620,N_3419);
and U8485 (N_8485,N_2489,N_4681);
or U8486 (N_8486,N_3331,N_3788);
or U8487 (N_8487,N_1445,N_2640);
nand U8488 (N_8488,N_2019,N_2778);
nor U8489 (N_8489,N_130,N_1078);
or U8490 (N_8490,N_2072,N_3858);
and U8491 (N_8491,N_4030,N_3935);
xor U8492 (N_8492,N_4585,N_1313);
nor U8493 (N_8493,N_779,N_996);
or U8494 (N_8494,N_1018,N_4629);
nor U8495 (N_8495,N_1567,N_112);
nor U8496 (N_8496,N_631,N_1690);
and U8497 (N_8497,N_1063,N_101);
or U8498 (N_8498,N_848,N_4414);
nor U8499 (N_8499,N_585,N_4812);
xor U8500 (N_8500,N_2618,N_2092);
and U8501 (N_8501,N_2209,N_1298);
nand U8502 (N_8502,N_3415,N_2526);
nand U8503 (N_8503,N_3610,N_2003);
nor U8504 (N_8504,N_4629,N_1361);
and U8505 (N_8505,N_4384,N_3175);
nand U8506 (N_8506,N_1253,N_3285);
nor U8507 (N_8507,N_2208,N_3581);
nor U8508 (N_8508,N_129,N_772);
and U8509 (N_8509,N_925,N_3452);
nor U8510 (N_8510,N_3784,N_488);
nor U8511 (N_8511,N_2936,N_302);
nand U8512 (N_8512,N_698,N_1963);
nand U8513 (N_8513,N_2846,N_682);
nand U8514 (N_8514,N_1728,N_3760);
or U8515 (N_8515,N_3436,N_3626);
nor U8516 (N_8516,N_1329,N_1946);
and U8517 (N_8517,N_2955,N_3602);
and U8518 (N_8518,N_4291,N_1702);
nand U8519 (N_8519,N_542,N_727);
nand U8520 (N_8520,N_2724,N_1968);
or U8521 (N_8521,N_2010,N_517);
xor U8522 (N_8522,N_1835,N_986);
or U8523 (N_8523,N_2145,N_2265);
or U8524 (N_8524,N_4569,N_2042);
nor U8525 (N_8525,N_3949,N_1671);
nor U8526 (N_8526,N_1776,N_2995);
or U8527 (N_8527,N_2480,N_1375);
and U8528 (N_8528,N_2805,N_3785);
nor U8529 (N_8529,N_4539,N_668);
nand U8530 (N_8530,N_991,N_1499);
nor U8531 (N_8531,N_3075,N_4371);
and U8532 (N_8532,N_3750,N_1521);
or U8533 (N_8533,N_4054,N_23);
and U8534 (N_8534,N_1927,N_224);
or U8535 (N_8535,N_460,N_2381);
and U8536 (N_8536,N_1828,N_4471);
nor U8537 (N_8537,N_2067,N_4315);
xnor U8538 (N_8538,N_263,N_2368);
and U8539 (N_8539,N_1259,N_3990);
or U8540 (N_8540,N_3494,N_4232);
nand U8541 (N_8541,N_72,N_1782);
and U8542 (N_8542,N_3733,N_1792);
xnor U8543 (N_8543,N_1555,N_3005);
or U8544 (N_8544,N_3157,N_3172);
xor U8545 (N_8545,N_3034,N_687);
and U8546 (N_8546,N_1424,N_4370);
xnor U8547 (N_8547,N_2782,N_1851);
or U8548 (N_8548,N_1780,N_4045);
or U8549 (N_8549,N_6,N_1981);
or U8550 (N_8550,N_3003,N_3797);
or U8551 (N_8551,N_404,N_2295);
and U8552 (N_8552,N_2665,N_1134);
nor U8553 (N_8553,N_4071,N_986);
xnor U8554 (N_8554,N_2213,N_4388);
xnor U8555 (N_8555,N_2031,N_350);
or U8556 (N_8556,N_735,N_4309);
and U8557 (N_8557,N_3975,N_3968);
xnor U8558 (N_8558,N_2248,N_3918);
nand U8559 (N_8559,N_1733,N_650);
xor U8560 (N_8560,N_3048,N_3501);
or U8561 (N_8561,N_3249,N_4921);
nor U8562 (N_8562,N_3053,N_1467);
or U8563 (N_8563,N_3540,N_4022);
nand U8564 (N_8564,N_4391,N_16);
nand U8565 (N_8565,N_252,N_2699);
nand U8566 (N_8566,N_2294,N_4265);
nor U8567 (N_8567,N_3465,N_4676);
and U8568 (N_8568,N_1022,N_4523);
and U8569 (N_8569,N_1118,N_2487);
nor U8570 (N_8570,N_1587,N_2690);
or U8571 (N_8571,N_2798,N_4106);
nor U8572 (N_8572,N_1416,N_3438);
or U8573 (N_8573,N_4211,N_2015);
nand U8574 (N_8574,N_1729,N_1175);
nor U8575 (N_8575,N_3327,N_388);
and U8576 (N_8576,N_216,N_3509);
or U8577 (N_8577,N_904,N_1489);
xor U8578 (N_8578,N_3843,N_286);
nor U8579 (N_8579,N_504,N_2694);
or U8580 (N_8580,N_1915,N_4631);
and U8581 (N_8581,N_164,N_4813);
nand U8582 (N_8582,N_3654,N_2693);
nor U8583 (N_8583,N_956,N_1650);
nand U8584 (N_8584,N_4,N_4495);
and U8585 (N_8585,N_54,N_186);
or U8586 (N_8586,N_4822,N_785);
or U8587 (N_8587,N_4207,N_62);
nor U8588 (N_8588,N_2181,N_2757);
nor U8589 (N_8589,N_3957,N_2579);
nand U8590 (N_8590,N_1645,N_3247);
xor U8591 (N_8591,N_238,N_308);
nor U8592 (N_8592,N_4001,N_3316);
and U8593 (N_8593,N_1422,N_4931);
nand U8594 (N_8594,N_1445,N_3494);
nand U8595 (N_8595,N_1696,N_3826);
and U8596 (N_8596,N_903,N_4224);
or U8597 (N_8597,N_425,N_476);
xnor U8598 (N_8598,N_4883,N_2275);
nand U8599 (N_8599,N_1780,N_2246);
and U8600 (N_8600,N_1718,N_4570);
nor U8601 (N_8601,N_56,N_4835);
nor U8602 (N_8602,N_3250,N_304);
nand U8603 (N_8603,N_969,N_522);
and U8604 (N_8604,N_2058,N_2131);
nor U8605 (N_8605,N_1144,N_2487);
and U8606 (N_8606,N_556,N_1736);
nor U8607 (N_8607,N_1761,N_2847);
and U8608 (N_8608,N_4887,N_2386);
or U8609 (N_8609,N_1326,N_1105);
and U8610 (N_8610,N_4851,N_134);
and U8611 (N_8611,N_2739,N_4319);
nor U8612 (N_8612,N_2075,N_2943);
or U8613 (N_8613,N_2779,N_3245);
xor U8614 (N_8614,N_4816,N_2198);
xnor U8615 (N_8615,N_4129,N_634);
or U8616 (N_8616,N_4241,N_3570);
and U8617 (N_8617,N_2729,N_1323);
or U8618 (N_8618,N_1648,N_4484);
nand U8619 (N_8619,N_1511,N_2339);
nor U8620 (N_8620,N_4602,N_2568);
or U8621 (N_8621,N_2986,N_1822);
xor U8622 (N_8622,N_482,N_841);
nand U8623 (N_8623,N_4670,N_3291);
nand U8624 (N_8624,N_2607,N_2599);
and U8625 (N_8625,N_3818,N_2178);
or U8626 (N_8626,N_3213,N_2242);
nor U8627 (N_8627,N_672,N_1258);
and U8628 (N_8628,N_3362,N_1214);
nor U8629 (N_8629,N_2023,N_654);
nor U8630 (N_8630,N_3030,N_1673);
nor U8631 (N_8631,N_4471,N_4653);
or U8632 (N_8632,N_245,N_3215);
nand U8633 (N_8633,N_2867,N_1095);
and U8634 (N_8634,N_2655,N_4486);
or U8635 (N_8635,N_2790,N_3873);
nand U8636 (N_8636,N_500,N_1890);
or U8637 (N_8637,N_4061,N_4611);
and U8638 (N_8638,N_4581,N_1063);
nor U8639 (N_8639,N_4728,N_196);
or U8640 (N_8640,N_2539,N_4380);
nor U8641 (N_8641,N_673,N_4924);
xnor U8642 (N_8642,N_191,N_2984);
nand U8643 (N_8643,N_825,N_281);
nand U8644 (N_8644,N_4485,N_869);
nor U8645 (N_8645,N_471,N_1292);
nand U8646 (N_8646,N_556,N_4796);
and U8647 (N_8647,N_2148,N_3508);
or U8648 (N_8648,N_3233,N_3312);
nor U8649 (N_8649,N_4544,N_2544);
nand U8650 (N_8650,N_1959,N_1410);
nor U8651 (N_8651,N_169,N_3169);
nor U8652 (N_8652,N_2137,N_918);
or U8653 (N_8653,N_258,N_3553);
xnor U8654 (N_8654,N_318,N_785);
nand U8655 (N_8655,N_1980,N_3386);
nor U8656 (N_8656,N_2104,N_3770);
nor U8657 (N_8657,N_2250,N_1337);
and U8658 (N_8658,N_164,N_117);
nor U8659 (N_8659,N_92,N_432);
or U8660 (N_8660,N_762,N_4100);
and U8661 (N_8661,N_4106,N_130);
nor U8662 (N_8662,N_3495,N_1015);
nor U8663 (N_8663,N_2474,N_106);
nor U8664 (N_8664,N_2075,N_4939);
nand U8665 (N_8665,N_4779,N_3173);
xor U8666 (N_8666,N_3131,N_2874);
or U8667 (N_8667,N_4558,N_3931);
or U8668 (N_8668,N_4940,N_2640);
and U8669 (N_8669,N_4642,N_1905);
or U8670 (N_8670,N_3605,N_1346);
or U8671 (N_8671,N_3191,N_3691);
or U8672 (N_8672,N_3522,N_1637);
nand U8673 (N_8673,N_1925,N_4725);
nand U8674 (N_8674,N_2876,N_169);
or U8675 (N_8675,N_2952,N_1638);
nand U8676 (N_8676,N_3406,N_2111);
or U8677 (N_8677,N_1037,N_93);
nand U8678 (N_8678,N_1906,N_1225);
nor U8679 (N_8679,N_4950,N_475);
nor U8680 (N_8680,N_1283,N_2935);
and U8681 (N_8681,N_1919,N_498);
or U8682 (N_8682,N_914,N_1653);
or U8683 (N_8683,N_3723,N_365);
xnor U8684 (N_8684,N_189,N_4106);
xor U8685 (N_8685,N_3039,N_3754);
nor U8686 (N_8686,N_1046,N_4653);
nand U8687 (N_8687,N_3057,N_4794);
nor U8688 (N_8688,N_4347,N_341);
or U8689 (N_8689,N_2895,N_4211);
or U8690 (N_8690,N_4907,N_4400);
or U8691 (N_8691,N_4813,N_3750);
nor U8692 (N_8692,N_2510,N_3423);
and U8693 (N_8693,N_277,N_3597);
nor U8694 (N_8694,N_3147,N_2102);
xor U8695 (N_8695,N_1792,N_128);
xor U8696 (N_8696,N_2823,N_1335);
nor U8697 (N_8697,N_2786,N_1467);
nor U8698 (N_8698,N_2512,N_4842);
and U8699 (N_8699,N_1612,N_1535);
and U8700 (N_8700,N_596,N_2487);
xnor U8701 (N_8701,N_446,N_4204);
nor U8702 (N_8702,N_3617,N_4509);
and U8703 (N_8703,N_1836,N_572);
or U8704 (N_8704,N_1388,N_1904);
nor U8705 (N_8705,N_2171,N_677);
and U8706 (N_8706,N_2786,N_679);
and U8707 (N_8707,N_4553,N_3112);
nand U8708 (N_8708,N_3749,N_1127);
or U8709 (N_8709,N_3091,N_1371);
and U8710 (N_8710,N_2462,N_3348);
nand U8711 (N_8711,N_996,N_171);
nor U8712 (N_8712,N_262,N_3606);
nor U8713 (N_8713,N_3021,N_4156);
nor U8714 (N_8714,N_2844,N_1534);
and U8715 (N_8715,N_3296,N_183);
nand U8716 (N_8716,N_4196,N_2353);
nand U8717 (N_8717,N_2978,N_2084);
nand U8718 (N_8718,N_4262,N_3567);
or U8719 (N_8719,N_2656,N_4619);
and U8720 (N_8720,N_3400,N_1254);
and U8721 (N_8721,N_110,N_1025);
nand U8722 (N_8722,N_3427,N_3514);
and U8723 (N_8723,N_807,N_1482);
nor U8724 (N_8724,N_4031,N_2097);
and U8725 (N_8725,N_1391,N_1351);
xnor U8726 (N_8726,N_4054,N_2917);
or U8727 (N_8727,N_79,N_3367);
xor U8728 (N_8728,N_1297,N_2934);
or U8729 (N_8729,N_1810,N_3510);
nand U8730 (N_8730,N_577,N_2569);
or U8731 (N_8731,N_4237,N_4566);
nand U8732 (N_8732,N_3147,N_3291);
nand U8733 (N_8733,N_968,N_4033);
nand U8734 (N_8734,N_802,N_1799);
or U8735 (N_8735,N_4527,N_3149);
nand U8736 (N_8736,N_4711,N_2822);
or U8737 (N_8737,N_218,N_295);
nand U8738 (N_8738,N_3501,N_2844);
or U8739 (N_8739,N_2674,N_3648);
nor U8740 (N_8740,N_163,N_117);
nand U8741 (N_8741,N_1256,N_1862);
nand U8742 (N_8742,N_27,N_3461);
nand U8743 (N_8743,N_725,N_992);
nand U8744 (N_8744,N_4688,N_3404);
xor U8745 (N_8745,N_1639,N_3988);
or U8746 (N_8746,N_3536,N_22);
or U8747 (N_8747,N_3297,N_3592);
or U8748 (N_8748,N_3257,N_4533);
or U8749 (N_8749,N_4601,N_968);
nor U8750 (N_8750,N_1080,N_115);
xor U8751 (N_8751,N_4077,N_2995);
nand U8752 (N_8752,N_186,N_881);
nand U8753 (N_8753,N_3387,N_4504);
or U8754 (N_8754,N_4949,N_4661);
or U8755 (N_8755,N_825,N_2877);
nor U8756 (N_8756,N_2160,N_1767);
nor U8757 (N_8757,N_3212,N_3015);
and U8758 (N_8758,N_1929,N_4760);
or U8759 (N_8759,N_1415,N_2397);
and U8760 (N_8760,N_1356,N_79);
xor U8761 (N_8761,N_3186,N_2195);
and U8762 (N_8762,N_1701,N_4977);
and U8763 (N_8763,N_352,N_3014);
and U8764 (N_8764,N_665,N_4570);
and U8765 (N_8765,N_376,N_1026);
and U8766 (N_8766,N_3498,N_211);
and U8767 (N_8767,N_917,N_2790);
or U8768 (N_8768,N_1378,N_3787);
nor U8769 (N_8769,N_176,N_3687);
or U8770 (N_8770,N_946,N_3359);
nor U8771 (N_8771,N_674,N_3534);
and U8772 (N_8772,N_4061,N_3873);
nor U8773 (N_8773,N_187,N_1915);
nor U8774 (N_8774,N_878,N_2500);
xnor U8775 (N_8775,N_632,N_224);
or U8776 (N_8776,N_2355,N_2518);
nand U8777 (N_8777,N_2124,N_781);
and U8778 (N_8778,N_360,N_2796);
or U8779 (N_8779,N_2153,N_119);
xnor U8780 (N_8780,N_4383,N_564);
nor U8781 (N_8781,N_4459,N_998);
or U8782 (N_8782,N_4206,N_4673);
nand U8783 (N_8783,N_1922,N_625);
and U8784 (N_8784,N_3270,N_4984);
nor U8785 (N_8785,N_3430,N_1953);
nand U8786 (N_8786,N_1699,N_1935);
xor U8787 (N_8787,N_1509,N_2110);
xnor U8788 (N_8788,N_3346,N_3206);
nor U8789 (N_8789,N_4200,N_3368);
and U8790 (N_8790,N_4532,N_2719);
and U8791 (N_8791,N_23,N_3914);
xor U8792 (N_8792,N_3389,N_2128);
xnor U8793 (N_8793,N_3549,N_1492);
or U8794 (N_8794,N_125,N_2627);
xor U8795 (N_8795,N_3315,N_4535);
or U8796 (N_8796,N_2296,N_3215);
or U8797 (N_8797,N_1815,N_3441);
or U8798 (N_8798,N_3316,N_598);
nand U8799 (N_8799,N_1748,N_2608);
and U8800 (N_8800,N_2991,N_4346);
and U8801 (N_8801,N_1301,N_1037);
and U8802 (N_8802,N_4285,N_3027);
or U8803 (N_8803,N_1831,N_1820);
or U8804 (N_8804,N_2649,N_3139);
and U8805 (N_8805,N_646,N_2048);
and U8806 (N_8806,N_3779,N_1902);
or U8807 (N_8807,N_262,N_3118);
nand U8808 (N_8808,N_92,N_1707);
or U8809 (N_8809,N_3280,N_2685);
and U8810 (N_8810,N_4895,N_2013);
or U8811 (N_8811,N_3325,N_2081);
and U8812 (N_8812,N_4038,N_2243);
nand U8813 (N_8813,N_4018,N_3496);
nor U8814 (N_8814,N_4645,N_563);
nand U8815 (N_8815,N_1566,N_4738);
and U8816 (N_8816,N_462,N_3627);
nand U8817 (N_8817,N_3980,N_636);
nand U8818 (N_8818,N_4607,N_4508);
and U8819 (N_8819,N_2130,N_3593);
or U8820 (N_8820,N_2794,N_2184);
nor U8821 (N_8821,N_1108,N_1365);
nand U8822 (N_8822,N_470,N_4417);
nor U8823 (N_8823,N_4691,N_1315);
nand U8824 (N_8824,N_2308,N_4156);
and U8825 (N_8825,N_731,N_334);
nand U8826 (N_8826,N_930,N_2821);
and U8827 (N_8827,N_1819,N_4039);
nand U8828 (N_8828,N_166,N_3298);
nand U8829 (N_8829,N_2768,N_97);
or U8830 (N_8830,N_805,N_460);
or U8831 (N_8831,N_3537,N_1155);
xor U8832 (N_8832,N_2786,N_4560);
and U8833 (N_8833,N_671,N_794);
or U8834 (N_8834,N_4972,N_4598);
and U8835 (N_8835,N_45,N_2613);
xor U8836 (N_8836,N_1913,N_4104);
nand U8837 (N_8837,N_4668,N_1421);
or U8838 (N_8838,N_3721,N_4455);
and U8839 (N_8839,N_3710,N_2942);
nand U8840 (N_8840,N_4985,N_3473);
or U8841 (N_8841,N_3901,N_1139);
and U8842 (N_8842,N_4351,N_2895);
nand U8843 (N_8843,N_702,N_489);
nand U8844 (N_8844,N_1464,N_477);
xnor U8845 (N_8845,N_746,N_4358);
and U8846 (N_8846,N_4561,N_1403);
and U8847 (N_8847,N_3712,N_93);
nor U8848 (N_8848,N_1149,N_3791);
nor U8849 (N_8849,N_1486,N_104);
xor U8850 (N_8850,N_2688,N_2338);
or U8851 (N_8851,N_879,N_1407);
nand U8852 (N_8852,N_844,N_2267);
nand U8853 (N_8853,N_709,N_4445);
or U8854 (N_8854,N_137,N_1692);
and U8855 (N_8855,N_2913,N_4213);
and U8856 (N_8856,N_2833,N_2305);
nand U8857 (N_8857,N_1127,N_4392);
and U8858 (N_8858,N_1660,N_1063);
nor U8859 (N_8859,N_4482,N_2560);
or U8860 (N_8860,N_204,N_2455);
nor U8861 (N_8861,N_3416,N_2942);
nor U8862 (N_8862,N_381,N_2922);
nand U8863 (N_8863,N_1249,N_3507);
nand U8864 (N_8864,N_729,N_273);
nand U8865 (N_8865,N_2521,N_4870);
and U8866 (N_8866,N_3403,N_524);
nor U8867 (N_8867,N_1784,N_2200);
or U8868 (N_8868,N_462,N_2153);
nand U8869 (N_8869,N_4311,N_3257);
or U8870 (N_8870,N_488,N_1635);
nand U8871 (N_8871,N_3624,N_177);
and U8872 (N_8872,N_816,N_4210);
or U8873 (N_8873,N_4322,N_1293);
and U8874 (N_8874,N_1437,N_2381);
and U8875 (N_8875,N_3865,N_1947);
nand U8876 (N_8876,N_3780,N_381);
nand U8877 (N_8877,N_3203,N_737);
nor U8878 (N_8878,N_38,N_4758);
nor U8879 (N_8879,N_3570,N_4351);
nand U8880 (N_8880,N_1499,N_2599);
nand U8881 (N_8881,N_3343,N_1307);
nor U8882 (N_8882,N_1451,N_2919);
nor U8883 (N_8883,N_2572,N_2243);
nand U8884 (N_8884,N_1434,N_3772);
nand U8885 (N_8885,N_4645,N_819);
nor U8886 (N_8886,N_700,N_1613);
nand U8887 (N_8887,N_1999,N_544);
nor U8888 (N_8888,N_1976,N_1391);
or U8889 (N_8889,N_2356,N_4344);
xnor U8890 (N_8890,N_4179,N_2941);
xor U8891 (N_8891,N_1191,N_4579);
and U8892 (N_8892,N_3393,N_1074);
or U8893 (N_8893,N_663,N_2712);
xor U8894 (N_8894,N_1500,N_107);
and U8895 (N_8895,N_1749,N_793);
xor U8896 (N_8896,N_3615,N_472);
nor U8897 (N_8897,N_1714,N_1129);
and U8898 (N_8898,N_143,N_469);
nor U8899 (N_8899,N_3707,N_264);
nor U8900 (N_8900,N_1356,N_4912);
nor U8901 (N_8901,N_3334,N_3631);
xor U8902 (N_8902,N_4452,N_4603);
or U8903 (N_8903,N_1112,N_3183);
nand U8904 (N_8904,N_1868,N_3573);
xnor U8905 (N_8905,N_4802,N_4041);
xor U8906 (N_8906,N_38,N_593);
and U8907 (N_8907,N_2180,N_3917);
nor U8908 (N_8908,N_2959,N_386);
nor U8909 (N_8909,N_4928,N_2229);
nor U8910 (N_8910,N_1605,N_2796);
nor U8911 (N_8911,N_4882,N_6);
or U8912 (N_8912,N_760,N_2853);
or U8913 (N_8913,N_169,N_3358);
or U8914 (N_8914,N_4401,N_1455);
or U8915 (N_8915,N_467,N_1701);
nand U8916 (N_8916,N_2982,N_799);
nor U8917 (N_8917,N_2759,N_2602);
and U8918 (N_8918,N_317,N_1155);
nor U8919 (N_8919,N_4609,N_3468);
nand U8920 (N_8920,N_1405,N_1823);
nand U8921 (N_8921,N_4210,N_4835);
nand U8922 (N_8922,N_1038,N_2204);
or U8923 (N_8923,N_3747,N_640);
and U8924 (N_8924,N_4942,N_1128);
and U8925 (N_8925,N_2958,N_2590);
xor U8926 (N_8926,N_2768,N_4224);
nor U8927 (N_8927,N_1790,N_2186);
or U8928 (N_8928,N_4017,N_1993);
and U8929 (N_8929,N_1899,N_4415);
or U8930 (N_8930,N_3315,N_1443);
xor U8931 (N_8931,N_4228,N_3228);
nor U8932 (N_8932,N_1715,N_3828);
or U8933 (N_8933,N_2862,N_3315);
nand U8934 (N_8934,N_4098,N_2162);
xor U8935 (N_8935,N_761,N_982);
and U8936 (N_8936,N_833,N_4555);
nor U8937 (N_8937,N_4894,N_2218);
and U8938 (N_8938,N_4455,N_2630);
or U8939 (N_8939,N_1761,N_1500);
nand U8940 (N_8940,N_935,N_1911);
and U8941 (N_8941,N_780,N_2618);
xnor U8942 (N_8942,N_418,N_4245);
xnor U8943 (N_8943,N_4564,N_3602);
and U8944 (N_8944,N_3821,N_2979);
and U8945 (N_8945,N_1205,N_1514);
or U8946 (N_8946,N_2078,N_365);
and U8947 (N_8947,N_3721,N_560);
xor U8948 (N_8948,N_4812,N_2666);
nor U8949 (N_8949,N_4503,N_2302);
nor U8950 (N_8950,N_1543,N_3612);
and U8951 (N_8951,N_4572,N_4871);
xor U8952 (N_8952,N_2423,N_1809);
nand U8953 (N_8953,N_908,N_2920);
nor U8954 (N_8954,N_3978,N_1131);
and U8955 (N_8955,N_1783,N_4376);
or U8956 (N_8956,N_2463,N_1728);
nand U8957 (N_8957,N_959,N_1992);
nor U8958 (N_8958,N_3303,N_1498);
nor U8959 (N_8959,N_2812,N_2959);
nor U8960 (N_8960,N_4695,N_1313);
nor U8961 (N_8961,N_1725,N_4523);
nor U8962 (N_8962,N_2252,N_56);
nand U8963 (N_8963,N_4727,N_2748);
nand U8964 (N_8964,N_3614,N_4939);
nand U8965 (N_8965,N_189,N_3631);
nand U8966 (N_8966,N_1964,N_1632);
and U8967 (N_8967,N_4228,N_3507);
xor U8968 (N_8968,N_4748,N_2824);
nor U8969 (N_8969,N_3079,N_4463);
nor U8970 (N_8970,N_4509,N_492);
nand U8971 (N_8971,N_3657,N_2507);
or U8972 (N_8972,N_4409,N_3024);
xnor U8973 (N_8973,N_2870,N_1133);
nand U8974 (N_8974,N_176,N_1860);
and U8975 (N_8975,N_672,N_145);
nand U8976 (N_8976,N_1302,N_2486);
nor U8977 (N_8977,N_1871,N_1580);
nor U8978 (N_8978,N_2782,N_2325);
or U8979 (N_8979,N_3132,N_2842);
or U8980 (N_8980,N_1985,N_3468);
nor U8981 (N_8981,N_3483,N_1917);
nor U8982 (N_8982,N_370,N_1616);
or U8983 (N_8983,N_404,N_2353);
nand U8984 (N_8984,N_1320,N_3482);
nor U8985 (N_8985,N_472,N_1556);
nor U8986 (N_8986,N_1034,N_1280);
nor U8987 (N_8987,N_2478,N_1012);
nor U8988 (N_8988,N_2354,N_301);
or U8989 (N_8989,N_4675,N_690);
and U8990 (N_8990,N_345,N_1116);
and U8991 (N_8991,N_3689,N_3987);
and U8992 (N_8992,N_1184,N_980);
or U8993 (N_8993,N_1833,N_2320);
or U8994 (N_8994,N_4958,N_3345);
nand U8995 (N_8995,N_1313,N_3327);
and U8996 (N_8996,N_3199,N_3381);
and U8997 (N_8997,N_3099,N_2356);
xor U8998 (N_8998,N_4285,N_1490);
or U8999 (N_8999,N_4358,N_784);
nand U9000 (N_9000,N_4622,N_4666);
nand U9001 (N_9001,N_3758,N_4156);
nor U9002 (N_9002,N_3436,N_2050);
and U9003 (N_9003,N_2684,N_3175);
and U9004 (N_9004,N_959,N_2033);
xor U9005 (N_9005,N_4758,N_4909);
xnor U9006 (N_9006,N_1599,N_1331);
nor U9007 (N_9007,N_4194,N_3089);
nor U9008 (N_9008,N_2079,N_630);
nor U9009 (N_9009,N_2226,N_1065);
nor U9010 (N_9010,N_145,N_2465);
and U9011 (N_9011,N_1572,N_3110);
xnor U9012 (N_9012,N_374,N_2874);
or U9013 (N_9013,N_1342,N_2713);
and U9014 (N_9014,N_4522,N_517);
or U9015 (N_9015,N_4476,N_200);
or U9016 (N_9016,N_2474,N_768);
and U9017 (N_9017,N_2594,N_3585);
xnor U9018 (N_9018,N_3937,N_2669);
nand U9019 (N_9019,N_3598,N_95);
or U9020 (N_9020,N_617,N_4621);
nor U9021 (N_9021,N_4474,N_1795);
nand U9022 (N_9022,N_1750,N_988);
xnor U9023 (N_9023,N_1749,N_3686);
nand U9024 (N_9024,N_1794,N_2529);
nor U9025 (N_9025,N_1351,N_941);
or U9026 (N_9026,N_4361,N_3755);
nand U9027 (N_9027,N_779,N_171);
xor U9028 (N_9028,N_3004,N_402);
nor U9029 (N_9029,N_4922,N_4216);
nor U9030 (N_9030,N_345,N_2798);
and U9031 (N_9031,N_2021,N_4363);
or U9032 (N_9032,N_4563,N_959);
nand U9033 (N_9033,N_3385,N_1759);
nor U9034 (N_9034,N_2504,N_2875);
nor U9035 (N_9035,N_3835,N_2765);
or U9036 (N_9036,N_2334,N_4392);
nor U9037 (N_9037,N_846,N_1068);
nor U9038 (N_9038,N_414,N_2722);
nand U9039 (N_9039,N_4149,N_4266);
nor U9040 (N_9040,N_469,N_2023);
nor U9041 (N_9041,N_2635,N_3216);
or U9042 (N_9042,N_119,N_588);
nor U9043 (N_9043,N_136,N_754);
nor U9044 (N_9044,N_76,N_4420);
and U9045 (N_9045,N_767,N_2823);
xnor U9046 (N_9046,N_3634,N_3986);
nor U9047 (N_9047,N_4163,N_637);
nand U9048 (N_9048,N_4347,N_3762);
and U9049 (N_9049,N_4382,N_439);
or U9050 (N_9050,N_564,N_1559);
and U9051 (N_9051,N_204,N_608);
nor U9052 (N_9052,N_365,N_176);
and U9053 (N_9053,N_3173,N_2883);
and U9054 (N_9054,N_1096,N_3547);
nand U9055 (N_9055,N_322,N_5);
nand U9056 (N_9056,N_4187,N_449);
or U9057 (N_9057,N_413,N_2838);
nor U9058 (N_9058,N_3854,N_2447);
and U9059 (N_9059,N_10,N_3855);
xor U9060 (N_9060,N_3863,N_1965);
and U9061 (N_9061,N_4632,N_4721);
or U9062 (N_9062,N_1078,N_3935);
and U9063 (N_9063,N_1365,N_4430);
nand U9064 (N_9064,N_2720,N_934);
nand U9065 (N_9065,N_4613,N_621);
xor U9066 (N_9066,N_4759,N_2832);
nand U9067 (N_9067,N_4996,N_793);
nand U9068 (N_9068,N_3914,N_2262);
nor U9069 (N_9069,N_1569,N_4804);
nand U9070 (N_9070,N_1859,N_4929);
or U9071 (N_9071,N_2207,N_4637);
nand U9072 (N_9072,N_4965,N_4716);
or U9073 (N_9073,N_2211,N_3482);
or U9074 (N_9074,N_2455,N_3240);
and U9075 (N_9075,N_3786,N_669);
and U9076 (N_9076,N_272,N_4212);
or U9077 (N_9077,N_3747,N_288);
nor U9078 (N_9078,N_1724,N_910);
nor U9079 (N_9079,N_2691,N_3887);
and U9080 (N_9080,N_1118,N_3418);
nand U9081 (N_9081,N_3398,N_4317);
nand U9082 (N_9082,N_1324,N_789);
xnor U9083 (N_9083,N_734,N_2103);
and U9084 (N_9084,N_1714,N_3865);
or U9085 (N_9085,N_1624,N_3618);
and U9086 (N_9086,N_1810,N_1330);
nand U9087 (N_9087,N_4260,N_4913);
nand U9088 (N_9088,N_1077,N_385);
and U9089 (N_9089,N_4679,N_1593);
nand U9090 (N_9090,N_3952,N_4053);
and U9091 (N_9091,N_3311,N_4866);
or U9092 (N_9092,N_1909,N_766);
nand U9093 (N_9093,N_4513,N_3736);
nand U9094 (N_9094,N_3332,N_3105);
nand U9095 (N_9095,N_2483,N_4407);
or U9096 (N_9096,N_1148,N_998);
or U9097 (N_9097,N_3730,N_3154);
nand U9098 (N_9098,N_2246,N_3129);
xnor U9099 (N_9099,N_809,N_1589);
or U9100 (N_9100,N_3503,N_978);
nand U9101 (N_9101,N_1925,N_3105);
and U9102 (N_9102,N_782,N_2166);
xor U9103 (N_9103,N_1521,N_115);
nand U9104 (N_9104,N_4453,N_97);
nand U9105 (N_9105,N_2417,N_4951);
or U9106 (N_9106,N_464,N_4776);
or U9107 (N_9107,N_741,N_4111);
and U9108 (N_9108,N_3075,N_1935);
nand U9109 (N_9109,N_1663,N_1500);
xor U9110 (N_9110,N_1,N_4993);
nor U9111 (N_9111,N_4376,N_1058);
or U9112 (N_9112,N_2398,N_2296);
nand U9113 (N_9113,N_760,N_1750);
or U9114 (N_9114,N_3754,N_1614);
and U9115 (N_9115,N_1503,N_157);
nand U9116 (N_9116,N_3071,N_794);
and U9117 (N_9117,N_2760,N_1985);
and U9118 (N_9118,N_4552,N_4530);
and U9119 (N_9119,N_4051,N_4564);
or U9120 (N_9120,N_1381,N_1389);
nand U9121 (N_9121,N_232,N_498);
nor U9122 (N_9122,N_395,N_219);
nand U9123 (N_9123,N_1374,N_3447);
nand U9124 (N_9124,N_2004,N_1026);
and U9125 (N_9125,N_2881,N_4024);
and U9126 (N_9126,N_505,N_4233);
and U9127 (N_9127,N_3326,N_1523);
and U9128 (N_9128,N_2908,N_4328);
and U9129 (N_9129,N_854,N_1936);
xnor U9130 (N_9130,N_3697,N_539);
nor U9131 (N_9131,N_1862,N_1324);
nand U9132 (N_9132,N_2626,N_1791);
and U9133 (N_9133,N_206,N_705);
nor U9134 (N_9134,N_2721,N_110);
nor U9135 (N_9135,N_4196,N_270);
nor U9136 (N_9136,N_4477,N_1644);
and U9137 (N_9137,N_2242,N_2807);
nand U9138 (N_9138,N_2682,N_1438);
nand U9139 (N_9139,N_4867,N_1756);
nand U9140 (N_9140,N_508,N_2327);
and U9141 (N_9141,N_4078,N_2648);
nand U9142 (N_9142,N_719,N_571);
nand U9143 (N_9143,N_3478,N_2398);
nor U9144 (N_9144,N_2844,N_3031);
nor U9145 (N_9145,N_4138,N_2945);
nand U9146 (N_9146,N_4385,N_325);
and U9147 (N_9147,N_3007,N_2365);
and U9148 (N_9148,N_1314,N_1206);
nand U9149 (N_9149,N_947,N_4551);
and U9150 (N_9150,N_1740,N_1186);
or U9151 (N_9151,N_574,N_3070);
and U9152 (N_9152,N_2955,N_3261);
nand U9153 (N_9153,N_4990,N_3674);
xnor U9154 (N_9154,N_2213,N_1357);
and U9155 (N_9155,N_4613,N_2725);
or U9156 (N_9156,N_4283,N_2752);
nand U9157 (N_9157,N_3833,N_3731);
or U9158 (N_9158,N_3468,N_1721);
or U9159 (N_9159,N_449,N_700);
and U9160 (N_9160,N_3942,N_4281);
nand U9161 (N_9161,N_4630,N_4907);
xnor U9162 (N_9162,N_625,N_2081);
xor U9163 (N_9163,N_789,N_2828);
xor U9164 (N_9164,N_2701,N_4078);
and U9165 (N_9165,N_1181,N_2846);
or U9166 (N_9166,N_2757,N_4932);
or U9167 (N_9167,N_2323,N_717);
xnor U9168 (N_9168,N_1792,N_2917);
nor U9169 (N_9169,N_383,N_3643);
or U9170 (N_9170,N_4909,N_3268);
or U9171 (N_9171,N_202,N_573);
nor U9172 (N_9172,N_2060,N_107);
and U9173 (N_9173,N_4586,N_2232);
nand U9174 (N_9174,N_1885,N_2973);
nand U9175 (N_9175,N_2967,N_3065);
and U9176 (N_9176,N_609,N_1215);
and U9177 (N_9177,N_2231,N_2721);
xor U9178 (N_9178,N_3232,N_3205);
xnor U9179 (N_9179,N_3284,N_4454);
xnor U9180 (N_9180,N_1379,N_2688);
or U9181 (N_9181,N_3961,N_2392);
nand U9182 (N_9182,N_415,N_518);
xnor U9183 (N_9183,N_3568,N_2403);
and U9184 (N_9184,N_4002,N_969);
and U9185 (N_9185,N_2128,N_4388);
nor U9186 (N_9186,N_4860,N_3818);
or U9187 (N_9187,N_787,N_2145);
nand U9188 (N_9188,N_1516,N_4784);
nand U9189 (N_9189,N_279,N_1877);
nand U9190 (N_9190,N_4205,N_4561);
xnor U9191 (N_9191,N_1251,N_3960);
or U9192 (N_9192,N_3983,N_220);
or U9193 (N_9193,N_648,N_1345);
or U9194 (N_9194,N_986,N_3742);
nand U9195 (N_9195,N_3803,N_4062);
nand U9196 (N_9196,N_1155,N_4006);
nand U9197 (N_9197,N_762,N_1626);
nor U9198 (N_9198,N_1739,N_1576);
and U9199 (N_9199,N_3924,N_2590);
xor U9200 (N_9200,N_3474,N_408);
or U9201 (N_9201,N_1061,N_3923);
nand U9202 (N_9202,N_1606,N_3063);
and U9203 (N_9203,N_1280,N_4558);
nand U9204 (N_9204,N_3003,N_2480);
and U9205 (N_9205,N_3372,N_3828);
xnor U9206 (N_9206,N_3955,N_2546);
nor U9207 (N_9207,N_1921,N_4914);
nand U9208 (N_9208,N_4002,N_3781);
nor U9209 (N_9209,N_4776,N_3077);
and U9210 (N_9210,N_915,N_4747);
nor U9211 (N_9211,N_3186,N_872);
nor U9212 (N_9212,N_3779,N_1840);
or U9213 (N_9213,N_4547,N_1699);
nand U9214 (N_9214,N_4955,N_911);
and U9215 (N_9215,N_440,N_2482);
nand U9216 (N_9216,N_4562,N_1912);
xor U9217 (N_9217,N_1144,N_2950);
or U9218 (N_9218,N_960,N_3242);
xnor U9219 (N_9219,N_1697,N_466);
or U9220 (N_9220,N_2240,N_4565);
xnor U9221 (N_9221,N_210,N_1850);
nor U9222 (N_9222,N_95,N_982);
xnor U9223 (N_9223,N_1982,N_3030);
xor U9224 (N_9224,N_366,N_4116);
or U9225 (N_9225,N_4801,N_1577);
nor U9226 (N_9226,N_1775,N_3333);
nor U9227 (N_9227,N_365,N_2477);
nand U9228 (N_9228,N_4020,N_4469);
and U9229 (N_9229,N_1808,N_1445);
xnor U9230 (N_9230,N_1295,N_1744);
nor U9231 (N_9231,N_3544,N_2049);
or U9232 (N_9232,N_830,N_2026);
xnor U9233 (N_9233,N_2643,N_4059);
or U9234 (N_9234,N_3434,N_799);
nor U9235 (N_9235,N_1165,N_1051);
and U9236 (N_9236,N_4517,N_2073);
nand U9237 (N_9237,N_1941,N_3764);
nand U9238 (N_9238,N_2190,N_3954);
nor U9239 (N_9239,N_1312,N_2940);
nor U9240 (N_9240,N_4024,N_4582);
or U9241 (N_9241,N_2425,N_4576);
nor U9242 (N_9242,N_201,N_1634);
and U9243 (N_9243,N_3010,N_3603);
and U9244 (N_9244,N_3226,N_1884);
nor U9245 (N_9245,N_2299,N_596);
and U9246 (N_9246,N_1509,N_4745);
xor U9247 (N_9247,N_1305,N_480);
nand U9248 (N_9248,N_1900,N_48);
nor U9249 (N_9249,N_1797,N_3372);
nor U9250 (N_9250,N_1889,N_4221);
or U9251 (N_9251,N_4139,N_4900);
xor U9252 (N_9252,N_2685,N_2262);
or U9253 (N_9253,N_2832,N_1120);
or U9254 (N_9254,N_73,N_4079);
xor U9255 (N_9255,N_4037,N_167);
or U9256 (N_9256,N_6,N_833);
xnor U9257 (N_9257,N_3179,N_4588);
and U9258 (N_9258,N_1761,N_3534);
and U9259 (N_9259,N_3395,N_1044);
nor U9260 (N_9260,N_1624,N_3948);
xnor U9261 (N_9261,N_315,N_4189);
and U9262 (N_9262,N_945,N_275);
and U9263 (N_9263,N_1347,N_302);
nor U9264 (N_9264,N_728,N_4674);
nand U9265 (N_9265,N_1399,N_457);
or U9266 (N_9266,N_3749,N_27);
nand U9267 (N_9267,N_3272,N_1805);
and U9268 (N_9268,N_1680,N_3155);
nor U9269 (N_9269,N_1338,N_248);
and U9270 (N_9270,N_2556,N_2147);
nand U9271 (N_9271,N_483,N_2167);
nand U9272 (N_9272,N_4526,N_2667);
or U9273 (N_9273,N_3271,N_3906);
nand U9274 (N_9274,N_3319,N_1600);
nand U9275 (N_9275,N_3203,N_3784);
or U9276 (N_9276,N_4455,N_412);
nor U9277 (N_9277,N_4302,N_145);
nand U9278 (N_9278,N_4865,N_2381);
xor U9279 (N_9279,N_1781,N_2846);
and U9280 (N_9280,N_3449,N_100);
nor U9281 (N_9281,N_4285,N_4318);
and U9282 (N_9282,N_4589,N_2280);
or U9283 (N_9283,N_2419,N_220);
nor U9284 (N_9284,N_1457,N_1070);
xnor U9285 (N_9285,N_823,N_4883);
and U9286 (N_9286,N_998,N_3833);
and U9287 (N_9287,N_877,N_3361);
xor U9288 (N_9288,N_738,N_735);
and U9289 (N_9289,N_3281,N_4703);
nor U9290 (N_9290,N_1142,N_1211);
nand U9291 (N_9291,N_3492,N_864);
xnor U9292 (N_9292,N_4164,N_4350);
and U9293 (N_9293,N_2620,N_1373);
nor U9294 (N_9294,N_4943,N_298);
nor U9295 (N_9295,N_1891,N_2140);
xor U9296 (N_9296,N_4074,N_3235);
and U9297 (N_9297,N_3581,N_2217);
nand U9298 (N_9298,N_266,N_675);
or U9299 (N_9299,N_3253,N_2775);
nand U9300 (N_9300,N_3049,N_2159);
or U9301 (N_9301,N_3991,N_2202);
nor U9302 (N_9302,N_1930,N_1153);
nand U9303 (N_9303,N_2122,N_1868);
nand U9304 (N_9304,N_17,N_4456);
xor U9305 (N_9305,N_4187,N_1329);
or U9306 (N_9306,N_3174,N_1880);
nor U9307 (N_9307,N_183,N_1751);
xor U9308 (N_9308,N_2168,N_1552);
or U9309 (N_9309,N_3636,N_1993);
and U9310 (N_9310,N_4451,N_3748);
and U9311 (N_9311,N_2332,N_2924);
or U9312 (N_9312,N_4844,N_3914);
or U9313 (N_9313,N_3730,N_1781);
or U9314 (N_9314,N_4435,N_3452);
xor U9315 (N_9315,N_2972,N_295);
nand U9316 (N_9316,N_2875,N_2859);
xor U9317 (N_9317,N_4527,N_3675);
xnor U9318 (N_9318,N_686,N_2723);
nand U9319 (N_9319,N_1311,N_4448);
or U9320 (N_9320,N_4829,N_3412);
or U9321 (N_9321,N_1102,N_3332);
and U9322 (N_9322,N_1019,N_967);
and U9323 (N_9323,N_2273,N_38);
nand U9324 (N_9324,N_4606,N_488);
and U9325 (N_9325,N_3475,N_4632);
nor U9326 (N_9326,N_2957,N_1426);
xnor U9327 (N_9327,N_2519,N_4850);
nand U9328 (N_9328,N_4177,N_10);
or U9329 (N_9329,N_3489,N_4913);
or U9330 (N_9330,N_3775,N_3464);
xor U9331 (N_9331,N_1689,N_3184);
nand U9332 (N_9332,N_4151,N_3290);
nand U9333 (N_9333,N_1541,N_3185);
nand U9334 (N_9334,N_4036,N_3374);
nor U9335 (N_9335,N_1519,N_2782);
and U9336 (N_9336,N_4156,N_3902);
nand U9337 (N_9337,N_1945,N_1794);
nor U9338 (N_9338,N_2158,N_3408);
nor U9339 (N_9339,N_3720,N_3067);
or U9340 (N_9340,N_1441,N_3815);
nand U9341 (N_9341,N_4664,N_458);
nand U9342 (N_9342,N_1347,N_3553);
nand U9343 (N_9343,N_4687,N_2320);
nor U9344 (N_9344,N_4858,N_3423);
and U9345 (N_9345,N_865,N_3391);
nor U9346 (N_9346,N_4354,N_3422);
nor U9347 (N_9347,N_3369,N_3231);
xnor U9348 (N_9348,N_3418,N_2117);
nor U9349 (N_9349,N_958,N_2431);
and U9350 (N_9350,N_3226,N_4214);
and U9351 (N_9351,N_2511,N_3806);
nor U9352 (N_9352,N_1889,N_2995);
nand U9353 (N_9353,N_113,N_2440);
nand U9354 (N_9354,N_3900,N_1382);
nor U9355 (N_9355,N_636,N_627);
nor U9356 (N_9356,N_4245,N_3273);
and U9357 (N_9357,N_664,N_3524);
or U9358 (N_9358,N_3272,N_712);
nor U9359 (N_9359,N_1339,N_744);
and U9360 (N_9360,N_385,N_2917);
and U9361 (N_9361,N_3397,N_153);
or U9362 (N_9362,N_2610,N_1406);
nor U9363 (N_9363,N_1015,N_2095);
nor U9364 (N_9364,N_4226,N_3450);
and U9365 (N_9365,N_2837,N_2253);
and U9366 (N_9366,N_188,N_3239);
nand U9367 (N_9367,N_4781,N_4909);
xnor U9368 (N_9368,N_472,N_623);
or U9369 (N_9369,N_2708,N_1873);
xnor U9370 (N_9370,N_668,N_2711);
nor U9371 (N_9371,N_1535,N_3376);
and U9372 (N_9372,N_457,N_2424);
and U9373 (N_9373,N_3940,N_4028);
nor U9374 (N_9374,N_1352,N_2664);
nand U9375 (N_9375,N_3562,N_4278);
xor U9376 (N_9376,N_475,N_4047);
xnor U9377 (N_9377,N_1277,N_1133);
and U9378 (N_9378,N_133,N_3285);
nand U9379 (N_9379,N_1037,N_4445);
or U9380 (N_9380,N_300,N_2956);
xor U9381 (N_9381,N_1564,N_3795);
and U9382 (N_9382,N_4588,N_3379);
and U9383 (N_9383,N_360,N_991);
nor U9384 (N_9384,N_4401,N_4383);
nor U9385 (N_9385,N_3047,N_2096);
and U9386 (N_9386,N_3162,N_688);
and U9387 (N_9387,N_3995,N_1657);
nor U9388 (N_9388,N_2817,N_3321);
and U9389 (N_9389,N_610,N_4370);
and U9390 (N_9390,N_3394,N_2319);
nand U9391 (N_9391,N_1765,N_2257);
nand U9392 (N_9392,N_3955,N_4690);
nand U9393 (N_9393,N_4479,N_4176);
or U9394 (N_9394,N_1846,N_4769);
xor U9395 (N_9395,N_4072,N_2537);
and U9396 (N_9396,N_1519,N_4787);
and U9397 (N_9397,N_1231,N_2913);
nand U9398 (N_9398,N_1489,N_302);
nand U9399 (N_9399,N_1101,N_3881);
xor U9400 (N_9400,N_3506,N_3637);
and U9401 (N_9401,N_1267,N_1142);
or U9402 (N_9402,N_4541,N_3598);
nor U9403 (N_9403,N_2725,N_2216);
or U9404 (N_9404,N_1442,N_3603);
and U9405 (N_9405,N_3868,N_295);
nor U9406 (N_9406,N_2649,N_4157);
nand U9407 (N_9407,N_4734,N_343);
nand U9408 (N_9408,N_1995,N_4027);
or U9409 (N_9409,N_1236,N_162);
xnor U9410 (N_9410,N_1559,N_2341);
nor U9411 (N_9411,N_1302,N_3240);
nor U9412 (N_9412,N_4781,N_3315);
nor U9413 (N_9413,N_1802,N_3197);
or U9414 (N_9414,N_1396,N_2912);
nand U9415 (N_9415,N_1573,N_919);
or U9416 (N_9416,N_2514,N_2618);
or U9417 (N_9417,N_3685,N_4179);
and U9418 (N_9418,N_1761,N_3674);
nand U9419 (N_9419,N_1416,N_4475);
or U9420 (N_9420,N_130,N_583);
and U9421 (N_9421,N_1487,N_2889);
or U9422 (N_9422,N_1221,N_491);
nand U9423 (N_9423,N_926,N_4936);
nand U9424 (N_9424,N_343,N_65);
and U9425 (N_9425,N_1749,N_4381);
xor U9426 (N_9426,N_4096,N_343);
xor U9427 (N_9427,N_2156,N_1921);
nor U9428 (N_9428,N_1595,N_2669);
and U9429 (N_9429,N_2273,N_4295);
or U9430 (N_9430,N_1211,N_4501);
xnor U9431 (N_9431,N_2485,N_1793);
nor U9432 (N_9432,N_3543,N_2985);
nor U9433 (N_9433,N_1656,N_3757);
and U9434 (N_9434,N_1020,N_4614);
or U9435 (N_9435,N_407,N_2621);
or U9436 (N_9436,N_2660,N_2110);
or U9437 (N_9437,N_4866,N_1884);
xnor U9438 (N_9438,N_228,N_3531);
nand U9439 (N_9439,N_1031,N_1097);
nand U9440 (N_9440,N_2507,N_570);
nor U9441 (N_9441,N_2111,N_2479);
or U9442 (N_9442,N_195,N_4468);
nor U9443 (N_9443,N_2803,N_3574);
or U9444 (N_9444,N_141,N_3769);
nand U9445 (N_9445,N_2074,N_3476);
and U9446 (N_9446,N_2558,N_1616);
xor U9447 (N_9447,N_3180,N_3469);
and U9448 (N_9448,N_775,N_1500);
or U9449 (N_9449,N_3947,N_482);
xor U9450 (N_9450,N_4843,N_1346);
or U9451 (N_9451,N_4444,N_35);
or U9452 (N_9452,N_463,N_2199);
and U9453 (N_9453,N_1587,N_1520);
nand U9454 (N_9454,N_4659,N_222);
or U9455 (N_9455,N_4039,N_16);
nand U9456 (N_9456,N_104,N_339);
or U9457 (N_9457,N_4380,N_1490);
nor U9458 (N_9458,N_2871,N_2158);
and U9459 (N_9459,N_1440,N_1817);
or U9460 (N_9460,N_3151,N_3948);
or U9461 (N_9461,N_3787,N_3936);
and U9462 (N_9462,N_4324,N_4268);
nand U9463 (N_9463,N_3224,N_8);
xor U9464 (N_9464,N_2090,N_3912);
nand U9465 (N_9465,N_75,N_1374);
xnor U9466 (N_9466,N_4627,N_999);
nand U9467 (N_9467,N_1603,N_4654);
xnor U9468 (N_9468,N_4809,N_1424);
nand U9469 (N_9469,N_120,N_1730);
xor U9470 (N_9470,N_2084,N_654);
nand U9471 (N_9471,N_1396,N_146);
nor U9472 (N_9472,N_3809,N_726);
or U9473 (N_9473,N_3934,N_4446);
and U9474 (N_9474,N_393,N_102);
or U9475 (N_9475,N_3592,N_4635);
or U9476 (N_9476,N_3219,N_1837);
nor U9477 (N_9477,N_2640,N_3648);
nand U9478 (N_9478,N_3427,N_4973);
nor U9479 (N_9479,N_4173,N_4076);
and U9480 (N_9480,N_4384,N_4746);
or U9481 (N_9481,N_1031,N_3617);
or U9482 (N_9482,N_1417,N_2388);
and U9483 (N_9483,N_3960,N_3572);
or U9484 (N_9484,N_1338,N_2523);
xor U9485 (N_9485,N_1156,N_4268);
or U9486 (N_9486,N_3299,N_158);
and U9487 (N_9487,N_525,N_2792);
or U9488 (N_9488,N_2684,N_2231);
nor U9489 (N_9489,N_458,N_1394);
and U9490 (N_9490,N_3163,N_748);
or U9491 (N_9491,N_955,N_1989);
xnor U9492 (N_9492,N_4417,N_2869);
xor U9493 (N_9493,N_1324,N_3081);
nand U9494 (N_9494,N_679,N_3577);
xor U9495 (N_9495,N_3082,N_1722);
or U9496 (N_9496,N_1132,N_4353);
xnor U9497 (N_9497,N_2368,N_2297);
nand U9498 (N_9498,N_1343,N_240);
and U9499 (N_9499,N_4713,N_4627);
xor U9500 (N_9500,N_74,N_2686);
and U9501 (N_9501,N_524,N_4587);
nand U9502 (N_9502,N_1765,N_2887);
or U9503 (N_9503,N_4415,N_2817);
nand U9504 (N_9504,N_2050,N_1589);
nor U9505 (N_9505,N_2161,N_4715);
nor U9506 (N_9506,N_1457,N_3619);
and U9507 (N_9507,N_284,N_900);
or U9508 (N_9508,N_2655,N_978);
and U9509 (N_9509,N_2713,N_2356);
and U9510 (N_9510,N_162,N_3045);
nor U9511 (N_9511,N_3807,N_732);
and U9512 (N_9512,N_2603,N_44);
and U9513 (N_9513,N_1558,N_459);
nor U9514 (N_9514,N_3202,N_4161);
and U9515 (N_9515,N_880,N_3943);
nor U9516 (N_9516,N_360,N_441);
or U9517 (N_9517,N_4115,N_4805);
xnor U9518 (N_9518,N_1833,N_622);
xor U9519 (N_9519,N_1846,N_1912);
nand U9520 (N_9520,N_2516,N_4968);
nor U9521 (N_9521,N_1637,N_3563);
or U9522 (N_9522,N_953,N_984);
or U9523 (N_9523,N_453,N_4059);
and U9524 (N_9524,N_2968,N_3437);
nor U9525 (N_9525,N_1370,N_642);
and U9526 (N_9526,N_1667,N_3815);
nor U9527 (N_9527,N_4372,N_3847);
nand U9528 (N_9528,N_186,N_1925);
and U9529 (N_9529,N_1044,N_122);
and U9530 (N_9530,N_4633,N_4524);
nor U9531 (N_9531,N_1305,N_2495);
or U9532 (N_9532,N_573,N_4971);
nor U9533 (N_9533,N_2179,N_961);
xor U9534 (N_9534,N_2015,N_2591);
and U9535 (N_9535,N_4111,N_4519);
nand U9536 (N_9536,N_3820,N_2867);
or U9537 (N_9537,N_4200,N_1595);
nand U9538 (N_9538,N_3462,N_511);
nor U9539 (N_9539,N_3535,N_4988);
nand U9540 (N_9540,N_1888,N_1586);
nand U9541 (N_9541,N_3657,N_436);
nor U9542 (N_9542,N_2065,N_2921);
nand U9543 (N_9543,N_4702,N_347);
and U9544 (N_9544,N_2995,N_493);
or U9545 (N_9545,N_1006,N_3209);
or U9546 (N_9546,N_4107,N_1848);
or U9547 (N_9547,N_3573,N_858);
and U9548 (N_9548,N_4871,N_4900);
nor U9549 (N_9549,N_3010,N_1555);
and U9550 (N_9550,N_4109,N_4873);
nand U9551 (N_9551,N_215,N_220);
nor U9552 (N_9552,N_280,N_855);
or U9553 (N_9553,N_909,N_4340);
nor U9554 (N_9554,N_31,N_519);
and U9555 (N_9555,N_966,N_144);
xor U9556 (N_9556,N_3638,N_3990);
or U9557 (N_9557,N_322,N_3849);
or U9558 (N_9558,N_66,N_2883);
nor U9559 (N_9559,N_4444,N_1664);
nor U9560 (N_9560,N_750,N_3483);
xnor U9561 (N_9561,N_4243,N_4013);
nand U9562 (N_9562,N_1709,N_3891);
and U9563 (N_9563,N_156,N_1419);
and U9564 (N_9564,N_2962,N_3848);
nor U9565 (N_9565,N_3757,N_4617);
and U9566 (N_9566,N_2528,N_4540);
or U9567 (N_9567,N_3499,N_1109);
nand U9568 (N_9568,N_3389,N_507);
nor U9569 (N_9569,N_3274,N_2005);
and U9570 (N_9570,N_1518,N_3650);
nor U9571 (N_9571,N_2371,N_2125);
or U9572 (N_9572,N_1777,N_2353);
nor U9573 (N_9573,N_1184,N_4616);
nor U9574 (N_9574,N_3549,N_172);
nor U9575 (N_9575,N_1705,N_1932);
xnor U9576 (N_9576,N_100,N_1211);
or U9577 (N_9577,N_2084,N_3850);
or U9578 (N_9578,N_2292,N_450);
or U9579 (N_9579,N_2979,N_3083);
or U9580 (N_9580,N_4856,N_2177);
or U9581 (N_9581,N_3652,N_3391);
nand U9582 (N_9582,N_1383,N_4252);
nor U9583 (N_9583,N_213,N_153);
nor U9584 (N_9584,N_654,N_2987);
and U9585 (N_9585,N_4506,N_4887);
or U9586 (N_9586,N_514,N_4180);
and U9587 (N_9587,N_3395,N_4784);
and U9588 (N_9588,N_4516,N_3953);
nor U9589 (N_9589,N_738,N_1391);
or U9590 (N_9590,N_2619,N_2638);
or U9591 (N_9591,N_2553,N_1713);
nor U9592 (N_9592,N_4048,N_1555);
nand U9593 (N_9593,N_3514,N_2338);
nand U9594 (N_9594,N_1679,N_1246);
xor U9595 (N_9595,N_3983,N_916);
nor U9596 (N_9596,N_2942,N_290);
xor U9597 (N_9597,N_1426,N_1768);
and U9598 (N_9598,N_768,N_4865);
nor U9599 (N_9599,N_4378,N_432);
or U9600 (N_9600,N_4974,N_4416);
and U9601 (N_9601,N_3214,N_628);
or U9602 (N_9602,N_4974,N_1005);
and U9603 (N_9603,N_1938,N_4658);
and U9604 (N_9604,N_3829,N_4947);
nand U9605 (N_9605,N_4183,N_1046);
nor U9606 (N_9606,N_1832,N_4180);
nor U9607 (N_9607,N_3288,N_529);
nand U9608 (N_9608,N_4004,N_1996);
and U9609 (N_9609,N_793,N_1834);
or U9610 (N_9610,N_33,N_891);
or U9611 (N_9611,N_2840,N_4839);
nor U9612 (N_9612,N_4939,N_1499);
nor U9613 (N_9613,N_2553,N_2126);
or U9614 (N_9614,N_2630,N_528);
nand U9615 (N_9615,N_3141,N_1538);
or U9616 (N_9616,N_4814,N_3386);
or U9617 (N_9617,N_3683,N_483);
xnor U9618 (N_9618,N_578,N_2710);
nand U9619 (N_9619,N_1070,N_322);
nor U9620 (N_9620,N_181,N_2869);
or U9621 (N_9621,N_2828,N_4175);
nand U9622 (N_9622,N_1138,N_542);
nand U9623 (N_9623,N_3432,N_3135);
nor U9624 (N_9624,N_3456,N_706);
and U9625 (N_9625,N_3789,N_1689);
nand U9626 (N_9626,N_2324,N_4290);
nand U9627 (N_9627,N_4579,N_3227);
nand U9628 (N_9628,N_655,N_4421);
nand U9629 (N_9629,N_652,N_2677);
nor U9630 (N_9630,N_4093,N_4266);
nand U9631 (N_9631,N_4755,N_941);
nand U9632 (N_9632,N_2969,N_3045);
or U9633 (N_9633,N_2198,N_1867);
nand U9634 (N_9634,N_3757,N_1033);
or U9635 (N_9635,N_3629,N_621);
nor U9636 (N_9636,N_1730,N_289);
or U9637 (N_9637,N_468,N_4946);
and U9638 (N_9638,N_2767,N_766);
and U9639 (N_9639,N_2463,N_4775);
nand U9640 (N_9640,N_324,N_1715);
nand U9641 (N_9641,N_4308,N_1691);
nor U9642 (N_9642,N_3620,N_4574);
and U9643 (N_9643,N_1746,N_4478);
nor U9644 (N_9644,N_2132,N_2178);
xor U9645 (N_9645,N_2307,N_3184);
nor U9646 (N_9646,N_1444,N_473);
and U9647 (N_9647,N_617,N_3610);
nor U9648 (N_9648,N_3011,N_589);
and U9649 (N_9649,N_4796,N_889);
or U9650 (N_9650,N_2724,N_4251);
or U9651 (N_9651,N_488,N_651);
nor U9652 (N_9652,N_3991,N_4265);
nand U9653 (N_9653,N_791,N_4514);
and U9654 (N_9654,N_4197,N_2877);
nor U9655 (N_9655,N_1372,N_4126);
nand U9656 (N_9656,N_2507,N_185);
nor U9657 (N_9657,N_1445,N_3181);
xor U9658 (N_9658,N_2189,N_4135);
nand U9659 (N_9659,N_4599,N_4153);
and U9660 (N_9660,N_1324,N_2900);
and U9661 (N_9661,N_1947,N_2714);
or U9662 (N_9662,N_3052,N_298);
nor U9663 (N_9663,N_1007,N_3512);
nand U9664 (N_9664,N_4120,N_3997);
xnor U9665 (N_9665,N_2927,N_3934);
nor U9666 (N_9666,N_4663,N_3511);
nor U9667 (N_9667,N_4653,N_833);
or U9668 (N_9668,N_2314,N_1215);
nor U9669 (N_9669,N_827,N_1515);
and U9670 (N_9670,N_3640,N_3464);
and U9671 (N_9671,N_4184,N_2264);
xor U9672 (N_9672,N_2072,N_1426);
nor U9673 (N_9673,N_1068,N_1558);
xnor U9674 (N_9674,N_98,N_4797);
nor U9675 (N_9675,N_828,N_4057);
xnor U9676 (N_9676,N_963,N_2570);
nand U9677 (N_9677,N_1723,N_807);
nor U9678 (N_9678,N_3663,N_3391);
nand U9679 (N_9679,N_3339,N_1426);
nand U9680 (N_9680,N_1915,N_4999);
xnor U9681 (N_9681,N_4627,N_2652);
nand U9682 (N_9682,N_4008,N_3271);
and U9683 (N_9683,N_4593,N_3774);
or U9684 (N_9684,N_3681,N_4520);
nor U9685 (N_9685,N_2549,N_1358);
nor U9686 (N_9686,N_1277,N_34);
nand U9687 (N_9687,N_1491,N_3423);
or U9688 (N_9688,N_3669,N_1785);
and U9689 (N_9689,N_2737,N_2372);
nand U9690 (N_9690,N_157,N_2572);
nor U9691 (N_9691,N_2543,N_483);
or U9692 (N_9692,N_244,N_2864);
xnor U9693 (N_9693,N_1227,N_1040);
nand U9694 (N_9694,N_2603,N_768);
nand U9695 (N_9695,N_2014,N_2326);
xnor U9696 (N_9696,N_1153,N_2199);
and U9697 (N_9697,N_2462,N_3148);
nor U9698 (N_9698,N_1243,N_753);
or U9699 (N_9699,N_30,N_1025);
nor U9700 (N_9700,N_2252,N_728);
or U9701 (N_9701,N_3682,N_3164);
nor U9702 (N_9702,N_148,N_541);
nor U9703 (N_9703,N_4732,N_1860);
and U9704 (N_9704,N_3388,N_3039);
xor U9705 (N_9705,N_4505,N_906);
nand U9706 (N_9706,N_1192,N_1051);
and U9707 (N_9707,N_2953,N_2966);
nand U9708 (N_9708,N_4102,N_2633);
xnor U9709 (N_9709,N_748,N_3747);
or U9710 (N_9710,N_4906,N_231);
nor U9711 (N_9711,N_4169,N_1828);
nor U9712 (N_9712,N_548,N_2770);
nor U9713 (N_9713,N_4086,N_1145);
or U9714 (N_9714,N_2075,N_4660);
nor U9715 (N_9715,N_503,N_1622);
and U9716 (N_9716,N_853,N_604);
or U9717 (N_9717,N_581,N_1761);
or U9718 (N_9718,N_2152,N_3548);
and U9719 (N_9719,N_3866,N_4236);
nor U9720 (N_9720,N_1749,N_2821);
and U9721 (N_9721,N_4991,N_828);
and U9722 (N_9722,N_4116,N_1501);
or U9723 (N_9723,N_99,N_3302);
and U9724 (N_9724,N_935,N_742);
nor U9725 (N_9725,N_2558,N_658);
nand U9726 (N_9726,N_2705,N_1016);
or U9727 (N_9727,N_3699,N_3198);
nand U9728 (N_9728,N_1888,N_750);
or U9729 (N_9729,N_4876,N_708);
or U9730 (N_9730,N_4994,N_3169);
or U9731 (N_9731,N_4928,N_3503);
or U9732 (N_9732,N_2198,N_524);
nor U9733 (N_9733,N_2566,N_1270);
nand U9734 (N_9734,N_3369,N_2812);
nand U9735 (N_9735,N_663,N_829);
nor U9736 (N_9736,N_1543,N_4658);
or U9737 (N_9737,N_1429,N_242);
nand U9738 (N_9738,N_3655,N_1543);
and U9739 (N_9739,N_571,N_2640);
xnor U9740 (N_9740,N_3420,N_3866);
nand U9741 (N_9741,N_178,N_3062);
or U9742 (N_9742,N_1432,N_4404);
or U9743 (N_9743,N_3887,N_704);
nor U9744 (N_9744,N_1993,N_3662);
nor U9745 (N_9745,N_4179,N_311);
xnor U9746 (N_9746,N_2931,N_1780);
and U9747 (N_9747,N_2536,N_639);
and U9748 (N_9748,N_1225,N_2721);
nand U9749 (N_9749,N_1247,N_2527);
nor U9750 (N_9750,N_2518,N_1700);
xnor U9751 (N_9751,N_1680,N_1134);
and U9752 (N_9752,N_4020,N_845);
and U9753 (N_9753,N_4301,N_3182);
or U9754 (N_9754,N_1697,N_917);
nor U9755 (N_9755,N_1057,N_41);
and U9756 (N_9756,N_2336,N_3403);
nor U9757 (N_9757,N_1650,N_4144);
xnor U9758 (N_9758,N_3803,N_198);
nor U9759 (N_9759,N_3046,N_4057);
and U9760 (N_9760,N_100,N_4497);
or U9761 (N_9761,N_2431,N_3552);
nor U9762 (N_9762,N_491,N_2);
and U9763 (N_9763,N_4092,N_1362);
xor U9764 (N_9764,N_576,N_3374);
and U9765 (N_9765,N_4846,N_2502);
xnor U9766 (N_9766,N_638,N_2330);
nor U9767 (N_9767,N_4891,N_245);
nor U9768 (N_9768,N_152,N_4787);
or U9769 (N_9769,N_3277,N_4545);
and U9770 (N_9770,N_2044,N_2523);
or U9771 (N_9771,N_4082,N_3753);
and U9772 (N_9772,N_2810,N_1599);
and U9773 (N_9773,N_2964,N_4540);
xnor U9774 (N_9774,N_624,N_2724);
nand U9775 (N_9775,N_4851,N_3533);
or U9776 (N_9776,N_4437,N_697);
nand U9777 (N_9777,N_855,N_2756);
nand U9778 (N_9778,N_718,N_3012);
nor U9779 (N_9779,N_157,N_1252);
nor U9780 (N_9780,N_1277,N_3229);
nand U9781 (N_9781,N_4998,N_1110);
nor U9782 (N_9782,N_161,N_3389);
nor U9783 (N_9783,N_2033,N_794);
or U9784 (N_9784,N_842,N_1277);
and U9785 (N_9785,N_4132,N_1963);
nand U9786 (N_9786,N_2883,N_3535);
and U9787 (N_9787,N_2501,N_1169);
nor U9788 (N_9788,N_514,N_3893);
or U9789 (N_9789,N_4898,N_4326);
nand U9790 (N_9790,N_4642,N_3641);
xnor U9791 (N_9791,N_1522,N_1752);
xor U9792 (N_9792,N_196,N_1719);
nand U9793 (N_9793,N_4281,N_482);
or U9794 (N_9794,N_660,N_1052);
nand U9795 (N_9795,N_4772,N_1798);
or U9796 (N_9796,N_1342,N_4856);
nand U9797 (N_9797,N_4867,N_3957);
nor U9798 (N_9798,N_3349,N_3816);
nand U9799 (N_9799,N_854,N_3034);
or U9800 (N_9800,N_317,N_3946);
nand U9801 (N_9801,N_2943,N_1044);
nand U9802 (N_9802,N_531,N_3310);
and U9803 (N_9803,N_1002,N_2223);
and U9804 (N_9804,N_726,N_1388);
or U9805 (N_9805,N_494,N_2224);
and U9806 (N_9806,N_2659,N_732);
nand U9807 (N_9807,N_2012,N_212);
or U9808 (N_9808,N_1930,N_4381);
or U9809 (N_9809,N_857,N_3895);
nor U9810 (N_9810,N_3394,N_3827);
and U9811 (N_9811,N_4992,N_3809);
nor U9812 (N_9812,N_3898,N_13);
or U9813 (N_9813,N_3260,N_2146);
nand U9814 (N_9814,N_1665,N_3575);
nand U9815 (N_9815,N_2242,N_277);
or U9816 (N_9816,N_2952,N_4729);
and U9817 (N_9817,N_3459,N_4077);
or U9818 (N_9818,N_578,N_352);
and U9819 (N_9819,N_1392,N_4253);
or U9820 (N_9820,N_4852,N_2444);
or U9821 (N_9821,N_1652,N_3958);
nand U9822 (N_9822,N_2836,N_3059);
nand U9823 (N_9823,N_4249,N_2654);
or U9824 (N_9824,N_4812,N_4050);
or U9825 (N_9825,N_1399,N_2995);
nand U9826 (N_9826,N_2326,N_438);
nand U9827 (N_9827,N_4920,N_77);
nor U9828 (N_9828,N_2535,N_4393);
or U9829 (N_9829,N_419,N_2466);
nor U9830 (N_9830,N_3608,N_4012);
nor U9831 (N_9831,N_3399,N_49);
nor U9832 (N_9832,N_2582,N_2143);
or U9833 (N_9833,N_1047,N_2418);
and U9834 (N_9834,N_1045,N_4020);
or U9835 (N_9835,N_1240,N_3720);
nor U9836 (N_9836,N_1901,N_605);
nor U9837 (N_9837,N_264,N_3268);
nand U9838 (N_9838,N_4747,N_833);
or U9839 (N_9839,N_3418,N_1760);
and U9840 (N_9840,N_3130,N_2534);
nand U9841 (N_9841,N_2103,N_2932);
nor U9842 (N_9842,N_3585,N_4728);
nand U9843 (N_9843,N_1405,N_3858);
or U9844 (N_9844,N_581,N_1925);
nor U9845 (N_9845,N_1960,N_3737);
xor U9846 (N_9846,N_2771,N_209);
nand U9847 (N_9847,N_705,N_2588);
or U9848 (N_9848,N_3100,N_3571);
nand U9849 (N_9849,N_3779,N_3940);
or U9850 (N_9850,N_3728,N_1727);
nand U9851 (N_9851,N_4080,N_4306);
and U9852 (N_9852,N_1324,N_1674);
and U9853 (N_9853,N_1036,N_3838);
nand U9854 (N_9854,N_4408,N_543);
nand U9855 (N_9855,N_4510,N_313);
or U9856 (N_9856,N_4044,N_3876);
nor U9857 (N_9857,N_2243,N_2988);
and U9858 (N_9858,N_3776,N_4257);
or U9859 (N_9859,N_4936,N_4451);
or U9860 (N_9860,N_4201,N_152);
nor U9861 (N_9861,N_2255,N_579);
nor U9862 (N_9862,N_4680,N_2058);
nand U9863 (N_9863,N_1868,N_1064);
nor U9864 (N_9864,N_1047,N_3008);
or U9865 (N_9865,N_3326,N_4178);
nor U9866 (N_9866,N_2632,N_4034);
or U9867 (N_9867,N_2504,N_3146);
and U9868 (N_9868,N_2098,N_2667);
or U9869 (N_9869,N_4524,N_828);
nor U9870 (N_9870,N_309,N_1009);
or U9871 (N_9871,N_970,N_2377);
and U9872 (N_9872,N_2401,N_4942);
nand U9873 (N_9873,N_2542,N_1956);
or U9874 (N_9874,N_3770,N_1173);
xnor U9875 (N_9875,N_1504,N_2948);
nand U9876 (N_9876,N_4481,N_4923);
and U9877 (N_9877,N_951,N_3608);
nand U9878 (N_9878,N_4771,N_1276);
or U9879 (N_9879,N_95,N_3597);
nor U9880 (N_9880,N_3805,N_3275);
or U9881 (N_9881,N_840,N_4594);
xnor U9882 (N_9882,N_1392,N_3638);
nor U9883 (N_9883,N_4923,N_4670);
and U9884 (N_9884,N_487,N_1942);
nand U9885 (N_9885,N_744,N_446);
or U9886 (N_9886,N_3922,N_258);
nand U9887 (N_9887,N_4835,N_1588);
nand U9888 (N_9888,N_3897,N_2396);
nor U9889 (N_9889,N_371,N_4047);
or U9890 (N_9890,N_751,N_1024);
and U9891 (N_9891,N_354,N_63);
xor U9892 (N_9892,N_4585,N_964);
and U9893 (N_9893,N_4806,N_3779);
and U9894 (N_9894,N_3887,N_4515);
and U9895 (N_9895,N_1800,N_570);
or U9896 (N_9896,N_1316,N_411);
or U9897 (N_9897,N_3412,N_1452);
and U9898 (N_9898,N_1796,N_2534);
or U9899 (N_9899,N_4920,N_3790);
nand U9900 (N_9900,N_3429,N_2880);
xnor U9901 (N_9901,N_4959,N_3462);
or U9902 (N_9902,N_4505,N_1733);
or U9903 (N_9903,N_3912,N_287);
xor U9904 (N_9904,N_679,N_2509);
or U9905 (N_9905,N_2124,N_2856);
nand U9906 (N_9906,N_3075,N_541);
or U9907 (N_9907,N_1492,N_2376);
nand U9908 (N_9908,N_4094,N_4689);
xor U9909 (N_9909,N_2092,N_269);
nand U9910 (N_9910,N_2029,N_4935);
nor U9911 (N_9911,N_235,N_495);
nand U9912 (N_9912,N_2700,N_2891);
nor U9913 (N_9913,N_4969,N_4389);
nor U9914 (N_9914,N_2773,N_4926);
or U9915 (N_9915,N_551,N_800);
nand U9916 (N_9916,N_4752,N_2134);
nand U9917 (N_9917,N_703,N_1307);
or U9918 (N_9918,N_343,N_2020);
or U9919 (N_9919,N_570,N_3406);
and U9920 (N_9920,N_4575,N_4038);
and U9921 (N_9921,N_3881,N_2119);
nand U9922 (N_9922,N_718,N_4415);
xor U9923 (N_9923,N_3979,N_1922);
nand U9924 (N_9924,N_3556,N_4756);
or U9925 (N_9925,N_1929,N_3076);
and U9926 (N_9926,N_232,N_4200);
or U9927 (N_9927,N_801,N_3438);
nand U9928 (N_9928,N_1856,N_3606);
and U9929 (N_9929,N_2710,N_204);
and U9930 (N_9930,N_3322,N_99);
nor U9931 (N_9931,N_1587,N_138);
and U9932 (N_9932,N_3352,N_4139);
and U9933 (N_9933,N_254,N_213);
nand U9934 (N_9934,N_2478,N_360);
nor U9935 (N_9935,N_815,N_2295);
or U9936 (N_9936,N_1554,N_2126);
nand U9937 (N_9937,N_3398,N_4893);
xnor U9938 (N_9938,N_3456,N_3731);
xor U9939 (N_9939,N_570,N_3883);
nand U9940 (N_9940,N_1346,N_3639);
or U9941 (N_9941,N_1977,N_4093);
and U9942 (N_9942,N_1038,N_4364);
and U9943 (N_9943,N_4618,N_2348);
nand U9944 (N_9944,N_3654,N_2216);
or U9945 (N_9945,N_4293,N_4053);
and U9946 (N_9946,N_226,N_363);
and U9947 (N_9947,N_1133,N_3210);
xnor U9948 (N_9948,N_2623,N_3558);
nor U9949 (N_9949,N_4021,N_409);
nor U9950 (N_9950,N_1895,N_2126);
or U9951 (N_9951,N_3526,N_4717);
nand U9952 (N_9952,N_2018,N_2587);
nand U9953 (N_9953,N_2892,N_3333);
xor U9954 (N_9954,N_36,N_1798);
xnor U9955 (N_9955,N_1618,N_2147);
or U9956 (N_9956,N_4938,N_272);
nand U9957 (N_9957,N_50,N_4154);
nand U9958 (N_9958,N_146,N_1488);
nand U9959 (N_9959,N_1536,N_2599);
or U9960 (N_9960,N_4034,N_1459);
nor U9961 (N_9961,N_1514,N_1552);
xor U9962 (N_9962,N_2912,N_4245);
xor U9963 (N_9963,N_2395,N_4471);
or U9964 (N_9964,N_518,N_2432);
xnor U9965 (N_9965,N_2134,N_1099);
and U9966 (N_9966,N_1059,N_2112);
and U9967 (N_9967,N_701,N_1511);
nand U9968 (N_9968,N_2084,N_3357);
nand U9969 (N_9969,N_2209,N_2421);
nor U9970 (N_9970,N_4873,N_975);
or U9971 (N_9971,N_797,N_4668);
nand U9972 (N_9972,N_1751,N_745);
xor U9973 (N_9973,N_225,N_3089);
and U9974 (N_9974,N_4874,N_4314);
nor U9975 (N_9975,N_3697,N_2056);
nand U9976 (N_9976,N_2061,N_3541);
nor U9977 (N_9977,N_4221,N_4543);
and U9978 (N_9978,N_2414,N_3023);
nor U9979 (N_9979,N_4254,N_2678);
and U9980 (N_9980,N_1251,N_4524);
xor U9981 (N_9981,N_3793,N_111);
and U9982 (N_9982,N_2901,N_4542);
nor U9983 (N_9983,N_2199,N_2395);
nor U9984 (N_9984,N_4834,N_1195);
and U9985 (N_9985,N_449,N_3085);
nor U9986 (N_9986,N_4784,N_4601);
nor U9987 (N_9987,N_124,N_1856);
xnor U9988 (N_9988,N_3443,N_2785);
or U9989 (N_9989,N_519,N_4438);
or U9990 (N_9990,N_1409,N_4839);
nand U9991 (N_9991,N_3679,N_1628);
and U9992 (N_9992,N_3196,N_626);
xor U9993 (N_9993,N_27,N_4159);
nor U9994 (N_9994,N_1573,N_4153);
and U9995 (N_9995,N_4962,N_1348);
xnor U9996 (N_9996,N_3901,N_2318);
nand U9997 (N_9997,N_1086,N_2888);
nor U9998 (N_9998,N_4934,N_1287);
nand U9999 (N_9999,N_4588,N_1868);
or UO_0 (O_0,N_6816,N_7467);
nor UO_1 (O_1,N_7153,N_5627);
nor UO_2 (O_2,N_9488,N_9102);
and UO_3 (O_3,N_6366,N_8100);
nor UO_4 (O_4,N_9287,N_6434);
and UO_5 (O_5,N_7227,N_8632);
nand UO_6 (O_6,N_7573,N_9069);
or UO_7 (O_7,N_9270,N_5936);
or UO_8 (O_8,N_5063,N_8954);
or UO_9 (O_9,N_8465,N_9346);
nor UO_10 (O_10,N_7068,N_8064);
or UO_11 (O_11,N_9882,N_9150);
and UO_12 (O_12,N_8760,N_8013);
nand UO_13 (O_13,N_8912,N_5266);
nor UO_14 (O_14,N_9414,N_7184);
and UO_15 (O_15,N_6668,N_7595);
nand UO_16 (O_16,N_5811,N_9062);
and UO_17 (O_17,N_9846,N_7278);
and UO_18 (O_18,N_8160,N_8681);
and UO_19 (O_19,N_8962,N_5338);
and UO_20 (O_20,N_8916,N_9923);
and UO_21 (O_21,N_7175,N_8303);
nand UO_22 (O_22,N_7634,N_6702);
nand UO_23 (O_23,N_6082,N_5222);
nand UO_24 (O_24,N_6266,N_8608);
nand UO_25 (O_25,N_5859,N_9098);
xor UO_26 (O_26,N_6454,N_8012);
nor UO_27 (O_27,N_7977,N_9440);
nor UO_28 (O_28,N_8667,N_6174);
nand UO_29 (O_29,N_8359,N_7860);
or UO_30 (O_30,N_5220,N_8476);
xor UO_31 (O_31,N_5658,N_7247);
xor UO_32 (O_32,N_6363,N_7204);
nor UO_33 (O_33,N_7295,N_9578);
and UO_34 (O_34,N_9646,N_9258);
nand UO_35 (O_35,N_5753,N_7297);
and UO_36 (O_36,N_9594,N_5927);
or UO_37 (O_37,N_8955,N_9004);
nor UO_38 (O_38,N_8726,N_9866);
and UO_39 (O_39,N_9693,N_7345);
or UO_40 (O_40,N_7260,N_9868);
nor UO_41 (O_41,N_9326,N_9557);
and UO_42 (O_42,N_5504,N_8414);
or UO_43 (O_43,N_5975,N_5704);
nor UO_44 (O_44,N_5180,N_8850);
or UO_45 (O_45,N_8157,N_5160);
nor UO_46 (O_46,N_8619,N_8818);
nand UO_47 (O_47,N_7360,N_6041);
xnor UO_48 (O_48,N_7543,N_7466);
nand UO_49 (O_49,N_6954,N_5521);
nand UO_50 (O_50,N_6704,N_5196);
and UO_51 (O_51,N_8136,N_5696);
or UO_52 (O_52,N_5730,N_5309);
xnor UO_53 (O_53,N_5208,N_6022);
nand UO_54 (O_54,N_9819,N_5534);
or UO_55 (O_55,N_5293,N_7660);
or UO_56 (O_56,N_6687,N_9931);
nand UO_57 (O_57,N_9768,N_7365);
nand UO_58 (O_58,N_8261,N_8801);
nand UO_59 (O_59,N_6949,N_5698);
or UO_60 (O_60,N_5914,N_9514);
and UO_61 (O_61,N_7172,N_7113);
xnor UO_62 (O_62,N_9147,N_8721);
nand UO_63 (O_63,N_8410,N_6480);
nor UO_64 (O_64,N_7575,N_5048);
nand UO_65 (O_65,N_5358,N_8092);
and UO_66 (O_66,N_6916,N_6197);
or UO_67 (O_67,N_5493,N_7045);
xnor UO_68 (O_68,N_9630,N_9058);
nand UO_69 (O_69,N_9815,N_6730);
nor UO_70 (O_70,N_8377,N_5605);
nand UO_71 (O_71,N_7048,N_8345);
or UO_72 (O_72,N_9009,N_5447);
or UO_73 (O_73,N_9785,N_6841);
nor UO_74 (O_74,N_7888,N_8066);
and UO_75 (O_75,N_6381,N_9177);
and UO_76 (O_76,N_6399,N_9411);
and UO_77 (O_77,N_5406,N_8483);
nand UO_78 (O_78,N_9811,N_6202);
or UO_79 (O_79,N_8282,N_5126);
and UO_80 (O_80,N_5672,N_7546);
nand UO_81 (O_81,N_8982,N_8798);
or UO_82 (O_82,N_7294,N_6377);
or UO_83 (O_83,N_5910,N_5072);
nor UO_84 (O_84,N_7323,N_5383);
nor UO_85 (O_85,N_5895,N_8533);
and UO_86 (O_86,N_8111,N_7579);
nor UO_87 (O_87,N_6539,N_8631);
or UO_88 (O_88,N_7273,N_8920);
nand UO_89 (O_89,N_5601,N_7628);
xor UO_90 (O_90,N_9528,N_5595);
and UO_91 (O_91,N_8174,N_9438);
or UO_92 (O_92,N_5989,N_7858);
or UO_93 (O_93,N_7079,N_5680);
nor UO_94 (O_94,N_5874,N_5779);
nand UO_95 (O_95,N_8244,N_5033);
nand UO_96 (O_96,N_5231,N_9219);
and UO_97 (O_97,N_6533,N_7845);
nand UO_98 (O_98,N_8919,N_7174);
nor UO_99 (O_99,N_5951,N_7953);
or UO_100 (O_100,N_8765,N_7838);
and UO_101 (O_101,N_8210,N_9130);
nand UO_102 (O_102,N_7824,N_7562);
and UO_103 (O_103,N_6674,N_7340);
nor UO_104 (O_104,N_5390,N_8892);
and UO_105 (O_105,N_9658,N_5246);
nand UO_106 (O_106,N_5070,N_8379);
or UO_107 (O_107,N_7028,N_5331);
nor UO_108 (O_108,N_8707,N_7016);
nor UO_109 (O_109,N_7932,N_6251);
or UO_110 (O_110,N_8062,N_9689);
and UO_111 (O_111,N_7058,N_5946);
nor UO_112 (O_112,N_9300,N_7551);
nand UO_113 (O_113,N_8078,N_8315);
or UO_114 (O_114,N_8588,N_8279);
nand UO_115 (O_115,N_7790,N_9490);
and UO_116 (O_116,N_7018,N_9104);
nand UO_117 (O_117,N_8081,N_9325);
or UO_118 (O_118,N_8591,N_5157);
nor UO_119 (O_119,N_7121,N_7631);
and UO_120 (O_120,N_7751,N_6190);
and UO_121 (O_121,N_7126,N_8418);
and UO_122 (O_122,N_6155,N_6906);
and UO_123 (O_123,N_9478,N_9645);
nor UO_124 (O_124,N_5064,N_7089);
nand UO_125 (O_125,N_6502,N_8233);
nor UO_126 (O_126,N_8799,N_7630);
nand UO_127 (O_127,N_5325,N_7830);
nor UO_128 (O_128,N_5422,N_6336);
and UO_129 (O_129,N_7646,N_7134);
xor UO_130 (O_130,N_8902,N_7480);
nand UO_131 (O_131,N_6770,N_7956);
nor UO_132 (O_132,N_5227,N_7428);
nand UO_133 (O_133,N_9535,N_7463);
and UO_134 (O_134,N_6523,N_6786);
nor UO_135 (O_135,N_9964,N_6573);
xnor UO_136 (O_136,N_7566,N_6810);
nand UO_137 (O_137,N_5796,N_6996);
nand UO_138 (O_138,N_7727,N_5117);
and UO_139 (O_139,N_6071,N_8580);
and UO_140 (O_140,N_9998,N_9371);
nor UO_141 (O_141,N_9196,N_8671);
and UO_142 (O_142,N_9877,N_7310);
xor UO_143 (O_143,N_6707,N_7210);
nor UO_144 (O_144,N_9782,N_7669);
nand UO_145 (O_145,N_7701,N_6520);
and UO_146 (O_146,N_6945,N_6782);
nor UO_147 (O_147,N_7168,N_5365);
xnor UO_148 (O_148,N_7689,N_5124);
and UO_149 (O_149,N_9840,N_8715);
and UO_150 (O_150,N_7479,N_9441);
nand UO_151 (O_151,N_9367,N_9970);
nor UO_152 (O_152,N_8384,N_6976);
or UO_153 (O_153,N_9719,N_7191);
or UO_154 (O_154,N_7283,N_8252);
xor UO_155 (O_155,N_9428,N_7009);
nand UO_156 (O_156,N_6552,N_9520);
or UO_157 (O_157,N_7155,N_8623);
nand UO_158 (O_158,N_9789,N_8457);
and UO_159 (O_159,N_6748,N_6441);
xor UO_160 (O_160,N_5566,N_5248);
and UO_161 (O_161,N_7642,N_5655);
nor UO_162 (O_162,N_7266,N_6603);
or UO_163 (O_163,N_7699,N_7907);
and UO_164 (O_164,N_8512,N_6402);
nand UO_165 (O_165,N_9424,N_6077);
and UO_166 (O_166,N_9422,N_5941);
and UO_167 (O_167,N_9568,N_7452);
nor UO_168 (O_168,N_5820,N_8658);
or UO_169 (O_169,N_9181,N_5702);
or UO_170 (O_170,N_8908,N_7607);
or UO_171 (O_171,N_7738,N_5660);
and UO_172 (O_172,N_8034,N_7785);
and UO_173 (O_173,N_9590,N_6873);
and UO_174 (O_174,N_7189,N_7133);
or UO_175 (O_175,N_5630,N_8971);
or UO_176 (O_176,N_5855,N_8529);
nand UO_177 (O_177,N_8978,N_7729);
nand UO_178 (O_178,N_5603,N_5904);
nand UO_179 (O_179,N_9257,N_9875);
nor UO_180 (O_180,N_6016,N_8290);
nor UO_181 (O_181,N_5861,N_6035);
nor UO_182 (O_182,N_7846,N_8725);
nand UO_183 (O_183,N_8177,N_8951);
and UO_184 (O_184,N_8438,N_9446);
nor UO_185 (O_185,N_9932,N_7866);
and UO_186 (O_186,N_9640,N_7734);
nand UO_187 (O_187,N_8989,N_9787);
and UO_188 (O_188,N_6461,N_6684);
nor UO_189 (O_189,N_8067,N_9118);
nor UO_190 (O_190,N_9691,N_6993);
and UO_191 (O_191,N_8472,N_5872);
and UO_192 (O_192,N_7443,N_7837);
or UO_193 (O_193,N_8685,N_6619);
or UO_194 (O_194,N_7987,N_6495);
xor UO_195 (O_195,N_9431,N_6013);
and UO_196 (O_196,N_8597,N_7447);
nor UO_197 (O_197,N_8621,N_6102);
and UO_198 (O_198,N_8170,N_8481);
or UO_199 (O_199,N_9682,N_8505);
nand UO_200 (O_200,N_9133,N_8873);
xnor UO_201 (O_201,N_8562,N_8168);
and UO_202 (O_202,N_8397,N_5743);
or UO_203 (O_203,N_7822,N_6239);
nor UO_204 (O_204,N_7921,N_6032);
nand UO_205 (O_205,N_9211,N_8149);
and UO_206 (O_206,N_5752,N_9224);
nor UO_207 (O_207,N_5025,N_5875);
and UO_208 (O_208,N_7770,N_9974);
and UO_209 (O_209,N_8464,N_8385);
nand UO_210 (O_210,N_7481,N_8637);
or UO_211 (O_211,N_7123,N_6419);
or UO_212 (O_212,N_7405,N_8566);
or UO_213 (O_213,N_7244,N_7939);
nand UO_214 (O_214,N_8497,N_8548);
nor UO_215 (O_215,N_5865,N_6459);
or UO_216 (O_216,N_5194,N_9844);
or UO_217 (O_217,N_6691,N_9045);
nor UO_218 (O_218,N_5242,N_8089);
and UO_219 (O_219,N_6739,N_8617);
nand UO_220 (O_220,N_6230,N_9936);
or UO_221 (O_221,N_7346,N_9401);
xor UO_222 (O_222,N_6838,N_7825);
nor UO_223 (O_223,N_8028,N_9777);
or UO_224 (O_224,N_8783,N_9399);
and UO_225 (O_225,N_6834,N_8599);
or UO_226 (O_226,N_6680,N_7591);
nor UO_227 (O_227,N_6617,N_5610);
nand UO_228 (O_228,N_7027,N_8361);
or UO_229 (O_229,N_7996,N_7690);
nand UO_230 (O_230,N_5744,N_8298);
nand UO_231 (O_231,N_6854,N_5669);
nor UO_232 (O_232,N_9569,N_9223);
xor UO_233 (O_233,N_9573,N_9989);
nor UO_234 (O_234,N_7150,N_6424);
or UO_235 (O_235,N_7781,N_8049);
nor UO_236 (O_236,N_9799,N_5021);
xor UO_237 (O_237,N_5091,N_5879);
nor UO_238 (O_238,N_8550,N_6964);
and UO_239 (O_239,N_6613,N_8589);
and UO_240 (O_240,N_6576,N_5028);
nor UO_241 (O_241,N_9048,N_7037);
and UO_242 (O_242,N_9671,N_9274);
xor UO_243 (O_243,N_5233,N_6558);
or UO_244 (O_244,N_8337,N_5312);
and UO_245 (O_245,N_7698,N_8346);
xnor UO_246 (O_246,N_9723,N_6132);
and UO_247 (O_247,N_5235,N_6870);
and UO_248 (O_248,N_5870,N_7508);
and UO_249 (O_249,N_6375,N_7313);
nor UO_250 (O_250,N_5092,N_8240);
nor UO_251 (O_251,N_9116,N_5396);
nor UO_252 (O_252,N_9135,N_9084);
nand UO_253 (O_253,N_9012,N_5199);
or UO_254 (O_254,N_7676,N_9697);
and UO_255 (O_255,N_7586,N_6373);
xor UO_256 (O_256,N_6051,N_8036);
or UO_257 (O_257,N_7792,N_7240);
or UO_258 (O_258,N_9008,N_8959);
nor UO_259 (O_259,N_5321,N_5835);
nor UO_260 (O_260,N_7118,N_9867);
nor UO_261 (O_261,N_6468,N_5186);
xnor UO_262 (O_262,N_9620,N_9080);
nand UO_263 (O_263,N_9195,N_8670);
or UO_264 (O_264,N_7687,N_8660);
xor UO_265 (O_265,N_8488,N_7311);
nor UO_266 (O_266,N_7710,N_9506);
nor UO_267 (O_267,N_9019,N_7299);
nor UO_268 (O_268,N_9930,N_6457);
nand UO_269 (O_269,N_8031,N_9014);
nor UO_270 (O_270,N_8146,N_5964);
nor UO_271 (O_271,N_8186,N_7571);
nor UO_272 (O_272,N_5797,N_9816);
and UO_273 (O_273,N_9835,N_6582);
nand UO_274 (O_274,N_9610,N_6073);
and UO_275 (O_275,N_8156,N_8937);
xnor UO_276 (O_276,N_7659,N_6852);
and UO_277 (O_277,N_6064,N_5451);
nor UO_278 (O_278,N_5361,N_5748);
nor UO_279 (O_279,N_5506,N_7811);
or UO_280 (O_280,N_6801,N_9797);
nand UO_281 (O_281,N_8435,N_9725);
xor UO_282 (O_282,N_9513,N_8241);
nor UO_283 (O_283,N_7072,N_8880);
or UO_284 (O_284,N_6660,N_7647);
nand UO_285 (O_285,N_7664,N_8368);
and UO_286 (O_286,N_8874,N_9255);
or UO_287 (O_287,N_5341,N_7952);
nor UO_288 (O_288,N_7139,N_9824);
xnor UO_289 (O_289,N_6020,N_6167);
nand UO_290 (O_290,N_9732,N_5116);
nor UO_291 (O_291,N_8077,N_8909);
or UO_292 (O_292,N_9123,N_7267);
nand UO_293 (O_293,N_5294,N_7601);
and UO_294 (O_294,N_8365,N_9540);
nand UO_295 (O_295,N_8705,N_7195);
nand UO_296 (O_296,N_6542,N_6235);
nand UO_297 (O_297,N_7362,N_7281);
and UO_298 (O_298,N_9872,N_5251);
nand UO_299 (O_299,N_5285,N_7693);
or UO_300 (O_300,N_6623,N_5228);
and UO_301 (O_301,N_5259,N_9209);
nor UO_302 (O_302,N_8322,N_6921);
and UO_303 (O_303,N_9920,N_6811);
and UO_304 (O_304,N_6608,N_8426);
or UO_305 (O_305,N_7022,N_8206);
and UO_306 (O_306,N_6878,N_5079);
nor UO_307 (O_307,N_9879,N_6820);
and UO_308 (O_308,N_5366,N_8331);
nor UO_309 (O_309,N_9025,N_8181);
and UO_310 (O_310,N_5237,N_5371);
or UO_311 (O_311,N_9337,N_5062);
or UO_312 (O_312,N_8574,N_9702);
or UO_313 (O_313,N_7109,N_7371);
and UO_314 (O_314,N_5773,N_8934);
or UO_315 (O_315,N_6380,N_7014);
nor UO_316 (O_316,N_7316,N_7842);
xnor UO_317 (O_317,N_5902,N_7820);
and UO_318 (O_318,N_8425,N_5844);
nor UO_319 (O_319,N_9153,N_7703);
nor UO_320 (O_320,N_5585,N_6165);
xnor UO_321 (O_321,N_9039,N_9064);
nor UO_322 (O_322,N_6118,N_5609);
or UO_323 (O_323,N_9017,N_7548);
or UO_324 (O_324,N_7626,N_7302);
and UO_325 (O_325,N_7459,N_6139);
and UO_326 (O_326,N_9612,N_6888);
xnor UO_327 (O_327,N_9584,N_8284);
and UO_328 (O_328,N_8524,N_5800);
nor UO_329 (O_329,N_8266,N_5621);
nor UO_330 (O_330,N_5250,N_9222);
nor UO_331 (O_331,N_5898,N_6559);
nor UO_332 (O_332,N_8444,N_5728);
or UO_333 (O_333,N_6683,N_8960);
and UO_334 (O_334,N_7783,N_6690);
or UO_335 (O_335,N_9420,N_7220);
and UO_336 (O_336,N_9475,N_6994);
nand UO_337 (O_337,N_6052,N_9581);
nand UO_338 (O_338,N_8947,N_5966);
nor UO_339 (O_339,N_6858,N_5801);
and UO_340 (O_340,N_9649,N_9751);
nor UO_341 (O_341,N_7377,N_9139);
or UO_342 (O_342,N_9455,N_6287);
and UO_343 (O_343,N_6876,N_8169);
nor UO_344 (O_344,N_8498,N_5398);
nor UO_345 (O_345,N_8992,N_7780);
nor UO_346 (O_346,N_9762,N_5831);
and UO_347 (O_347,N_8828,N_7230);
and UO_348 (O_348,N_8996,N_6761);
and UO_349 (O_349,N_5937,N_9873);
nand UO_350 (O_350,N_5135,N_7488);
xor UO_351 (O_351,N_8255,N_9742);
nor UO_352 (O_352,N_8964,N_8076);
nand UO_353 (O_353,N_9294,N_5734);
and UO_354 (O_354,N_6923,N_9954);
nor UO_355 (O_355,N_6688,N_8585);
nor UO_356 (O_356,N_8583,N_9097);
nand UO_357 (O_357,N_7937,N_7318);
nor UO_358 (O_358,N_5632,N_9040);
and UO_359 (O_359,N_7062,N_9885);
nand UO_360 (O_360,N_6224,N_9281);
and UO_361 (O_361,N_7730,N_9046);
and UO_362 (O_362,N_7216,N_8945);
and UO_363 (O_363,N_9463,N_6393);
nand UO_364 (O_364,N_5241,N_8222);
or UO_365 (O_365,N_5000,N_6312);
and UO_366 (O_366,N_9269,N_7233);
nor UO_367 (O_367,N_8938,N_6513);
xnor UO_368 (O_368,N_6788,N_7599);
or UO_369 (O_369,N_7531,N_8663);
and UO_370 (O_370,N_7504,N_9794);
and UO_371 (O_371,N_8265,N_8387);
and UO_372 (O_372,N_7159,N_5187);
nand UO_373 (O_373,N_5843,N_8198);
nand UO_374 (O_374,N_9731,N_5590);
nand UO_375 (O_375,N_7973,N_5007);
xor UO_376 (O_376,N_9156,N_9926);
and UO_377 (O_377,N_6449,N_5473);
and UO_378 (O_378,N_9328,N_9865);
xor UO_379 (O_379,N_6815,N_9734);
and UO_380 (O_380,N_6415,N_5083);
nor UO_381 (O_381,N_6370,N_9418);
or UO_382 (O_382,N_6134,N_7180);
nor UO_383 (O_383,N_7651,N_9173);
nand UO_384 (O_384,N_7328,N_9940);
and UO_385 (O_385,N_7806,N_8046);
nor UO_386 (O_386,N_8634,N_7582);
nand UO_387 (O_387,N_6848,N_9564);
nor UO_388 (O_388,N_6885,N_5697);
or UO_389 (O_389,N_7033,N_7795);
nand UO_390 (O_390,N_7298,N_5711);
nand UO_391 (O_391,N_7106,N_6396);
or UO_392 (O_392,N_7754,N_9306);
nand UO_393 (O_393,N_9072,N_6947);
or UO_394 (O_394,N_5105,N_7919);
and UO_395 (O_395,N_8159,N_6626);
nor UO_396 (O_396,N_7741,N_8833);
nand UO_397 (O_397,N_5284,N_6831);
nand UO_398 (O_398,N_9909,N_7352);
nand UO_399 (O_399,N_8351,N_8876);
nand UO_400 (O_400,N_9627,N_9503);
or UO_401 (O_401,N_6481,N_9398);
and UO_402 (O_402,N_8886,N_7388);
nand UO_403 (O_403,N_7308,N_8419);
nand UO_404 (O_404,N_8164,N_9733);
or UO_405 (O_405,N_7421,N_7881);
or UO_406 (O_406,N_8247,N_6836);
or UO_407 (O_407,N_5540,N_5298);
and UO_408 (O_408,N_6956,N_8942);
nor UO_409 (O_409,N_6443,N_5763);
and UO_410 (O_410,N_9461,N_8131);
xor UO_411 (O_411,N_5567,N_6531);
or UO_412 (O_412,N_6927,N_7193);
nor UO_413 (O_413,N_6200,N_8944);
nand UO_414 (O_414,N_8251,N_9555);
nor UO_415 (O_415,N_9928,N_7449);
nand UO_416 (O_416,N_9737,N_6673);
nand UO_417 (O_417,N_8382,N_8605);
nand UO_418 (O_418,N_6772,N_8118);
nand UO_419 (O_419,N_9899,N_7522);
and UO_420 (O_420,N_9218,N_8773);
or UO_421 (O_421,N_5706,N_5360);
nor UO_422 (O_422,N_9291,N_8291);
and UO_423 (O_423,N_7760,N_6837);
nand UO_424 (O_424,N_7334,N_9856);
nor UO_425 (O_425,N_6176,N_8858);
nand UO_426 (O_426,N_6732,N_5005);
nand UO_427 (O_427,N_9460,N_8877);
nand UO_428 (O_428,N_9624,N_9121);
and UO_429 (O_429,N_7503,N_7358);
or UO_430 (O_430,N_8907,N_7242);
and UO_431 (O_431,N_7151,N_9052);
nand UO_432 (O_432,N_7222,N_7841);
and UO_433 (O_433,N_8356,N_9798);
nand UO_434 (O_434,N_7201,N_7492);
nand UO_435 (O_435,N_8403,N_8396);
or UO_436 (O_436,N_9517,N_7890);
and UO_437 (O_437,N_9392,N_7359);
xnor UO_438 (O_438,N_9445,N_7199);
nor UO_439 (O_439,N_8037,N_5304);
and UO_440 (O_440,N_6605,N_6803);
xnor UO_441 (O_441,N_9988,N_9686);
nor UO_442 (O_442,N_6515,N_9245);
nor UO_443 (O_443,N_8620,N_9906);
nand UO_444 (O_444,N_9743,N_5615);
nand UO_445 (O_445,N_7686,N_6692);
and UO_446 (O_446,N_9747,N_5271);
and UO_447 (O_447,N_6965,N_6860);
and UO_448 (O_448,N_6302,N_6728);
xor UO_449 (O_449,N_5403,N_8995);
or UO_450 (O_450,N_6069,N_6045);
nor UO_451 (O_451,N_6059,N_5768);
nor UO_452 (O_452,N_7050,N_8571);
and UO_453 (O_453,N_9987,N_5348);
nor UO_454 (O_454,N_9484,N_9829);
and UO_455 (O_455,N_6522,N_8887);
nand UO_456 (O_456,N_8712,N_8504);
and UO_457 (O_457,N_5657,N_8421);
nand UO_458 (O_458,N_8534,N_7097);
and UO_459 (O_459,N_7563,N_8242);
nand UO_460 (O_460,N_8091,N_5172);
and UO_461 (O_461,N_5942,N_6737);
or UO_462 (O_462,N_8595,N_6483);
nand UO_463 (O_463,N_7988,N_7422);
and UO_464 (O_464,N_6561,N_7457);
or UO_465 (O_465,N_5799,N_8778);
and UO_466 (O_466,N_6809,N_8545);
and UO_467 (O_467,N_9466,N_7087);
and UO_468 (O_468,N_5700,N_5357);
and UO_469 (O_469,N_6484,N_5442);
and UO_470 (O_470,N_7836,N_7251);
or UO_471 (O_471,N_8269,N_6718);
and UO_472 (O_472,N_8102,N_7406);
nand UO_473 (O_473,N_6198,N_7098);
nor UO_474 (O_474,N_6318,N_9813);
or UO_475 (O_475,N_7556,N_8541);
nor UO_476 (O_476,N_6241,N_6494);
nand UO_477 (O_477,N_9107,N_7276);
nor UO_478 (O_478,N_7458,N_8044);
and UO_479 (O_479,N_5765,N_6631);
xor UO_480 (O_480,N_6247,N_9993);
nor UO_481 (O_481,N_7103,N_8364);
nor UO_482 (O_482,N_6612,N_8499);
or UO_483 (O_483,N_6106,N_5183);
nand UO_484 (O_484,N_6935,N_7483);
nand UO_485 (O_485,N_8626,N_7870);
nor UO_486 (O_486,N_6800,N_9990);
and UO_487 (O_487,N_9241,N_9028);
and UO_488 (O_488,N_5320,N_7125);
nor UO_489 (O_489,N_7526,N_9347);
nor UO_490 (O_490,N_7725,N_6417);
nor UO_491 (O_491,N_8007,N_6549);
xor UO_492 (O_492,N_9087,N_5467);
nor UO_493 (O_493,N_6168,N_7122);
nor UO_494 (O_494,N_6970,N_5616);
or UO_495 (O_495,N_7063,N_9101);
or UO_496 (O_496,N_6910,N_9796);
nand UO_497 (O_497,N_7671,N_8459);
nand UO_498 (O_498,N_8609,N_5095);
xnor UO_499 (O_499,N_9486,N_8979);
nor UO_500 (O_500,N_6076,N_7163);
or UO_501 (O_501,N_5234,N_6812);
nor UO_502 (O_502,N_8084,N_8313);
or UO_503 (O_503,N_9339,N_8711);
and UO_504 (O_504,N_7685,N_8319);
nor UO_505 (O_505,N_8336,N_9011);
nand UO_506 (O_506,N_6192,N_7071);
and UO_507 (O_507,N_5185,N_8753);
nor UO_508 (O_508,N_7259,N_5189);
nand UO_509 (O_509,N_7929,N_5878);
nor UO_510 (O_510,N_8065,N_7733);
and UO_511 (O_511,N_6769,N_7848);
and UO_512 (O_512,N_7765,N_7931);
or UO_513 (O_513,N_9884,N_5392);
and UO_514 (O_514,N_5470,N_7891);
nand UO_515 (O_515,N_5648,N_9700);
and UO_516 (O_516,N_8564,N_5296);
nor UO_517 (O_517,N_7407,N_7495);
or UO_518 (O_518,N_7381,N_8018);
and UO_519 (O_519,N_8482,N_7609);
nor UO_520 (O_520,N_7305,N_7682);
nand UO_521 (O_521,N_5009,N_8016);
or UO_522 (O_522,N_6569,N_8638);
nand UO_523 (O_523,N_5249,N_7612);
nand UO_524 (O_524,N_8466,N_5894);
and UO_525 (O_525,N_8948,N_7275);
and UO_526 (O_526,N_6705,N_9966);
nand UO_527 (O_527,N_8703,N_6510);
and UO_528 (O_528,N_5653,N_8894);
nor UO_529 (O_529,N_9566,N_9515);
xor UO_530 (O_530,N_9717,N_6460);
xnor UO_531 (O_531,N_7808,N_8127);
nand UO_532 (O_532,N_7214,N_8791);
or UO_533 (O_533,N_8087,N_9730);
or UO_534 (O_534,N_7982,N_8781);
nand UO_535 (O_535,N_5539,N_5337);
or UO_536 (O_536,N_7083,N_6669);
xor UO_537 (O_537,N_8200,N_7010);
nor UO_538 (O_538,N_7665,N_7702);
or UO_539 (O_539,N_6455,N_6903);
nor UO_540 (O_540,N_9388,N_7246);
nor UO_541 (O_541,N_5416,N_5507);
and UO_542 (O_542,N_9828,N_5935);
or UO_543 (O_543,N_9242,N_5038);
nand UO_544 (O_544,N_5301,N_7615);
nor UO_545 (O_545,N_9470,N_7320);
and UO_546 (O_546,N_5568,N_7788);
nand UO_547 (O_547,N_9207,N_7331);
or UO_548 (O_548,N_8939,N_8596);
or UO_549 (O_549,N_9950,N_9193);
xnor UO_550 (O_550,N_5625,N_8821);
nand UO_551 (O_551,N_8560,N_6227);
nor UO_552 (O_552,N_8249,N_8800);
and UO_553 (O_553,N_9905,N_9534);
nor UO_554 (O_554,N_6265,N_9316);
nor UO_555 (O_555,N_5441,N_7085);
nor UO_556 (O_556,N_6070,N_7593);
nand UO_557 (O_557,N_9007,N_8603);
xnor UO_558 (O_558,N_7786,N_9061);
nand UO_559 (O_559,N_9823,N_5553);
or UO_560 (O_560,N_9208,N_9305);
or UO_561 (O_561,N_6763,N_6754);
and UO_562 (O_562,N_9477,N_5466);
and UO_563 (O_563,N_8101,N_7622);
nor UO_564 (O_564,N_5832,N_5992);
nand UO_565 (O_565,N_9359,N_9370);
and UO_566 (O_566,N_9340,N_9068);
nor UO_567 (O_567,N_5054,N_5051);
xor UO_568 (O_568,N_7131,N_5058);
nand UO_569 (O_569,N_5343,N_9343);
nor UO_570 (O_570,N_9355,N_5377);
nand UO_571 (O_571,N_6212,N_6987);
and UO_572 (O_572,N_5359,N_9576);
nor UO_573 (O_573,N_8203,N_7417);
or UO_574 (O_574,N_9298,N_8841);
nand UO_575 (O_575,N_6024,N_5528);
or UO_576 (O_576,N_6430,N_6436);
and UO_577 (O_577,N_6049,N_8445);
nand UO_578 (O_578,N_9738,N_6137);
and UO_579 (O_579,N_9286,N_8370);
xor UO_580 (O_580,N_8473,N_6904);
or UO_581 (O_581,N_8323,N_8510);
nand UO_582 (O_582,N_5085,N_6113);
or UO_583 (O_583,N_9049,N_5130);
and UO_584 (O_584,N_6093,N_6555);
nor UO_585 (O_585,N_6160,N_8838);
xor UO_586 (O_586,N_5414,N_7088);
or UO_587 (O_587,N_9295,N_5275);
nor UO_588 (O_588,N_9413,N_9076);
nor UO_589 (O_589,N_5824,N_6216);
xnor UO_590 (O_590,N_9452,N_8229);
or UO_591 (O_591,N_5583,N_7794);
or UO_592 (O_592,N_5440,N_5970);
xor UO_593 (O_593,N_7818,N_7756);
xor UO_594 (O_594,N_7460,N_5308);
nand UO_595 (O_595,N_9876,N_7167);
or UO_596 (O_596,N_6278,N_6395);
or UO_597 (O_597,N_8508,N_8148);
nand UO_598 (O_598,N_6978,N_8576);
or UO_599 (O_599,N_5956,N_9330);
or UO_600 (O_600,N_9059,N_8694);
or UO_601 (O_601,N_6767,N_7857);
nand UO_602 (O_602,N_6665,N_6050);
and UO_603 (O_603,N_9511,N_8360);
or UO_604 (O_604,N_6914,N_5662);
and UO_605 (O_605,N_6727,N_6151);
and UO_606 (O_606,N_9838,N_7961);
or UO_607 (O_607,N_5101,N_5755);
or UO_608 (O_608,N_6115,N_6796);
nor UO_609 (O_609,N_7559,N_6210);
or UO_610 (O_610,N_7402,N_7319);
nand UO_611 (O_611,N_9955,N_8546);
nand UO_612 (O_612,N_9016,N_7537);
and UO_613 (O_613,N_9927,N_9758);
or UO_614 (O_614,N_5112,N_5770);
and UO_615 (O_615,N_7117,N_5570);
xnor UO_616 (O_616,N_7885,N_7494);
nand UO_617 (O_617,N_8227,N_8415);
or UO_618 (O_618,N_5689,N_5805);
or UO_619 (O_619,N_6144,N_5232);
nor UO_620 (O_620,N_9744,N_5151);
or UO_621 (O_621,N_9801,N_9396);
nor UO_622 (O_622,N_9676,N_8602);
nor UO_623 (O_623,N_9234,N_8348);
nand UO_624 (O_624,N_7752,N_5848);
or UO_625 (O_625,N_8350,N_6342);
and UO_626 (O_626,N_9615,N_8305);
xnor UO_627 (O_627,N_8698,N_7802);
nor UO_628 (O_628,N_6643,N_6636);
and UO_629 (O_629,N_5532,N_8641);
or UO_630 (O_630,N_9449,N_5710);
and UO_631 (O_631,N_8584,N_6493);
nand UO_632 (O_632,N_8970,N_9945);
or UO_633 (O_633,N_6775,N_5342);
or UO_634 (O_634,N_5443,N_6233);
nor UO_635 (O_635,N_5519,N_9361);
nor UO_636 (O_636,N_5851,N_5210);
nand UO_637 (O_637,N_8152,N_7911);
and UO_638 (O_638,N_7194,N_5693);
or UO_639 (O_639,N_5524,N_6306);
nand UO_640 (O_640,N_6276,N_7621);
or UO_641 (O_641,N_7643,N_8352);
nand UO_642 (O_642,N_5896,N_9124);
nor UO_643 (O_643,N_7111,N_7983);
nor UO_644 (O_644,N_8878,N_9709);
nand UO_645 (O_645,N_6999,N_6681);
or UO_646 (O_646,N_6063,N_8899);
or UO_647 (O_647,N_7017,N_9018);
or UO_648 (O_648,N_8769,N_9763);
nor UO_649 (O_649,N_9406,N_8374);
nand UO_650 (O_650,N_9228,N_8513);
nand UO_651 (O_651,N_7843,N_5917);
nand UO_652 (O_652,N_9454,N_6751);
nand UO_653 (O_653,N_9026,N_5651);
nor UO_654 (O_654,N_6188,N_7645);
and UO_655 (O_655,N_6438,N_5673);
nor UO_656 (O_656,N_6308,N_8984);
or UO_657 (O_657,N_6007,N_8808);
xnor UO_658 (O_658,N_8060,N_9817);
xor UO_659 (O_659,N_8104,N_7468);
nand UO_660 (O_660,N_9493,N_7572);
xnor UO_661 (O_661,N_5635,N_8301);
nor UO_662 (O_662,N_9704,N_8458);
and UO_663 (O_663,N_9580,N_6818);
nand UO_664 (O_664,N_5830,N_9903);
nor UO_665 (O_665,N_9395,N_8486);
or UO_666 (O_666,N_9650,N_9807);
nand UO_667 (O_667,N_7902,N_6654);
and UO_668 (O_668,N_7638,N_6969);
nand UO_669 (O_669,N_7557,N_5642);
and UO_670 (O_670,N_6099,N_7271);
or UO_671 (O_671,N_7816,N_9929);
nor UO_672 (O_672,N_5192,N_8278);
nor UO_673 (O_673,N_6781,N_8088);
nor UO_674 (O_674,N_6131,N_6516);
and UO_675 (O_675,N_8057,N_5336);
nor UO_676 (O_676,N_5240,N_5404);
and UO_677 (O_677,N_8806,N_9301);
or UO_678 (O_678,N_9975,N_6640);
nor UO_679 (O_679,N_5607,N_6547);
nor UO_680 (O_680,N_8777,N_5803);
xor UO_681 (O_681,N_6948,N_7673);
or UO_682 (O_682,N_8932,N_6034);
and UO_683 (O_683,N_8292,N_7854);
and UO_684 (O_684,N_6843,N_9654);
or UO_685 (O_685,N_8553,N_7598);
and UO_686 (O_686,N_9311,N_7903);
and UO_687 (O_687,N_7470,N_8719);
nor UO_688 (O_688,N_9164,N_8701);
nor UO_689 (O_689,N_9082,N_8429);
xnor UO_690 (O_690,N_9839,N_9263);
or UO_691 (O_691,N_9577,N_8940);
or UO_692 (O_692,N_6456,N_7205);
nand UO_693 (O_693,N_6206,N_8700);
or UO_694 (O_694,N_6122,N_8734);
and UO_695 (O_695,N_9290,N_6872);
xnor UO_696 (O_696,N_9772,N_6091);
or UO_697 (O_697,N_5893,N_5497);
and UO_698 (O_698,N_7964,N_6897);
nor UO_699 (O_699,N_8404,N_7416);
nand UO_700 (O_700,N_7721,N_9661);
nor UO_701 (O_701,N_5885,N_6661);
and UO_702 (O_702,N_8650,N_6095);
and UO_703 (O_703,N_5916,N_9942);
nor UO_704 (O_704,N_9962,N_8022);
or UO_705 (O_705,N_9670,N_8287);
nor UO_706 (O_706,N_6924,N_9354);
nor UO_707 (O_707,N_9659,N_6162);
nor UO_708 (O_708,N_9448,N_6296);
nor UO_709 (O_709,N_8235,N_6384);
nor UO_710 (O_710,N_8997,N_9111);
or UO_711 (O_711,N_8182,N_8134);
nand UO_712 (O_712,N_8554,N_5511);
xnor UO_713 (O_713,N_5487,N_8193);
and UO_714 (O_714,N_7823,N_6439);
xor UO_715 (O_715,N_5391,N_5245);
and UO_716 (O_716,N_7670,N_9718);
and UO_717 (O_717,N_7336,N_9114);
nand UO_718 (O_718,N_9053,N_7605);
nand UO_719 (O_719,N_8208,N_7577);
nor UO_720 (O_720,N_9368,N_7567);
nand UO_721 (O_721,N_8924,N_5382);
nand UO_722 (O_722,N_7719,N_9501);
or UO_723 (O_723,N_5475,N_9505);
or UO_724 (O_724,N_5812,N_8610);
nor UO_725 (O_725,N_8147,N_5129);
and UO_726 (O_726,N_6750,N_7827);
xor UO_727 (O_727,N_5884,N_6663);
nand UO_728 (O_728,N_7282,N_8810);
and UO_729 (O_729,N_9405,N_5537);
or UO_730 (O_730,N_5816,N_8961);
nor UO_731 (O_731,N_8762,N_9701);
or UO_732 (O_732,N_8295,N_8586);
xnor UO_733 (O_733,N_5792,N_7095);
nand UO_734 (O_734,N_5594,N_5972);
or UO_735 (O_735,N_6133,N_8544);
nand UO_736 (O_736,N_8212,N_7506);
nor UO_737 (O_737,N_8893,N_6437);
xor UO_738 (O_738,N_6755,N_9129);
nand UO_739 (O_739,N_7777,N_5419);
and UO_740 (O_740,N_8237,N_8433);
and UO_741 (O_741,N_8827,N_7709);
xnor UO_742 (O_742,N_7505,N_8647);
xnor UO_743 (O_743,N_6458,N_5317);
nand UO_744 (O_744,N_6762,N_6745);
nor UO_745 (O_745,N_9716,N_9754);
or UO_746 (O_746,N_9057,N_6793);
xor UO_747 (O_747,N_8462,N_5198);
and UO_748 (O_748,N_9657,N_8158);
xor UO_749 (O_749,N_6629,N_7812);
nand UO_750 (O_750,N_5899,N_6337);
nand UO_751 (O_751,N_5823,N_5102);
and UO_752 (O_752,N_9232,N_7678);
or UO_753 (O_753,N_6960,N_7813);
nor UO_754 (O_754,N_5980,N_5912);
nor UO_755 (O_755,N_6985,N_6696);
nor UO_756 (O_756,N_9915,N_6479);
and UO_757 (O_757,N_5269,N_6771);
and UO_758 (O_758,N_5516,N_9790);
or UO_759 (O_759,N_9137,N_8567);
or UO_760 (O_760,N_7241,N_5618);
nand UO_761 (O_761,N_8759,N_9679);
nor UO_762 (O_762,N_8881,N_9570);
nand UO_763 (O_763,N_9765,N_5453);
or UO_764 (O_764,N_7585,N_5077);
nor UO_765 (O_765,N_6779,N_5751);
and UO_766 (O_766,N_9722,N_7583);
nor UO_767 (O_767,N_9983,N_8803);
and UO_768 (O_768,N_7376,N_8543);
nor UO_769 (O_769,N_9358,N_7538);
and UO_770 (O_770,N_6807,N_5560);
and UO_771 (O_771,N_8549,N_6658);
nor UO_772 (O_772,N_7652,N_8475);
xor UO_773 (O_773,N_6466,N_9499);
nor UO_774 (O_774,N_9571,N_7799);
nor UO_775 (O_775,N_8570,N_5821);
or UO_776 (O_776,N_9889,N_8055);
nor UO_777 (O_777,N_9467,N_9711);
xor UO_778 (O_778,N_5709,N_9236);
nand UO_779 (O_779,N_5814,N_8573);
nand UO_780 (O_780,N_5900,N_8813);
nand UO_781 (O_781,N_5747,N_6475);
or UO_782 (O_782,N_8686,N_6094);
or UO_783 (O_783,N_6990,N_7196);
and UO_784 (O_784,N_5569,N_5412);
nand UO_785 (O_785,N_7206,N_8917);
or UO_786 (O_786,N_5978,N_6887);
nor UO_787 (O_787,N_8568,N_5159);
and UO_788 (O_788,N_6271,N_6072);
nor UO_789 (O_789,N_8117,N_8468);
or UO_790 (O_790,N_6822,N_5649);
and UO_791 (O_791,N_8006,N_6066);
nor UO_792 (O_792,N_8176,N_8230);
nand UO_793 (O_793,N_7763,N_8503);
or UO_794 (O_794,N_9814,N_9149);
nor UO_795 (O_795,N_7031,N_8552);
and UO_796 (O_796,N_7493,N_6238);
and UO_797 (O_797,N_8153,N_5988);
and UO_798 (O_798,N_8422,N_5217);
nor UO_799 (O_799,N_6014,N_9407);
and UO_800 (O_800,N_6778,N_6127);
xor UO_801 (O_801,N_8653,N_6290);
nor UO_802 (O_802,N_8051,N_5197);
xnor UO_803 (O_803,N_5993,N_7616);
and UO_804 (O_804,N_5692,N_6711);
or UO_805 (O_805,N_7826,N_8536);
nor UO_806 (O_806,N_9415,N_6599);
nor UO_807 (O_807,N_5690,N_8882);
xnor UO_808 (O_808,N_7096,N_5436);
or UO_809 (O_809,N_5236,N_8875);
nor UO_810 (O_810,N_8673,N_5850);
nand UO_811 (O_811,N_5745,N_9303);
xor UO_812 (O_812,N_8342,N_7476);
nand UO_813 (O_813,N_7766,N_5423);
or UO_814 (O_814,N_7277,N_6135);
nor UO_815 (O_815,N_7361,N_6998);
nand UO_816 (O_816,N_8930,N_6129);
or UO_817 (O_817,N_6894,N_6136);
nor UO_818 (O_818,N_6997,N_8434);
nor UO_819 (O_819,N_7712,N_8675);
or UO_820 (O_820,N_7086,N_6700);
nand UO_821 (O_821,N_5501,N_9695);
or UO_822 (O_822,N_6634,N_6936);
or UO_823 (O_823,N_7883,N_8285);
and UO_824 (O_824,N_9863,N_5287);
and UO_825 (O_825,N_7102,N_6753);
and UO_826 (O_826,N_6884,N_7875);
nor UO_827 (O_827,N_5863,N_7399);
or UO_828 (O_828,N_6245,N_7464);
nand UO_829 (O_829,N_7644,N_6175);
and UO_830 (O_830,N_8764,N_6637);
or UO_831 (O_831,N_7143,N_6189);
or UO_832 (O_832,N_8437,N_8752);
and UO_833 (O_833,N_6962,N_9525);
or UO_834 (O_834,N_6142,N_9869);
and UO_835 (O_835,N_7530,N_6228);
or UO_836 (O_836,N_7758,N_6657);
or UO_837 (O_837,N_8988,N_7304);
nand UO_838 (O_838,N_6108,N_7373);
nor UO_839 (O_839,N_8409,N_9843);
nor UO_840 (O_840,N_6957,N_7394);
or UO_841 (O_841,N_6886,N_7064);
and UO_842 (O_842,N_7596,N_6871);
or UO_843 (O_843,N_7592,N_7142);
and UO_844 (O_844,N_8957,N_5542);
nor UO_845 (O_845,N_6317,N_9169);
and UO_846 (O_846,N_8793,N_5252);
and UO_847 (O_847,N_5552,N_8795);
nor UO_848 (O_848,N_5195,N_8254);
nand UO_849 (O_849,N_7235,N_6534);
nor UO_850 (O_850,N_8207,N_7617);
xor UO_851 (O_851,N_6734,N_6411);
and UO_852 (O_852,N_6647,N_7667);
nand UO_853 (O_853,N_5399,N_8835);
xnor UO_854 (O_854,N_6929,N_8059);
and UO_855 (O_855,N_8871,N_8511);
and UO_856 (O_856,N_8910,N_9496);
nor UO_857 (O_857,N_5479,N_9162);
nor UO_858 (O_858,N_7183,N_7971);
or UO_859 (O_859,N_9497,N_7922);
or UO_860 (O_860,N_9288,N_6596);
xnor UO_861 (O_861,N_7951,N_6693);
or UO_862 (O_862,N_5551,N_7714);
or UO_863 (O_863,N_5345,N_7618);
nor UO_864 (O_864,N_7696,N_6857);
and UO_865 (O_865,N_8389,N_9382);
nand UO_866 (O_866,N_8043,N_6814);
or UO_867 (O_867,N_8058,N_8518);
or UO_868 (O_868,N_6802,N_5853);
xor UO_869 (O_869,N_6153,N_8749);
nor UO_870 (O_870,N_7547,N_7065);
or UO_871 (O_871,N_9617,N_9826);
or UO_872 (O_872,N_6604,N_8223);
nor UO_873 (O_873,N_6591,N_6314);
nor UO_874 (O_874,N_8751,N_5530);
nor UO_875 (O_875,N_7853,N_6499);
xor UO_876 (O_876,N_7980,N_5628);
or UO_877 (O_877,N_8891,N_5420);
nor UO_878 (O_878,N_8592,N_9421);
xor UO_879 (O_879,N_6252,N_7897);
nor UO_880 (O_880,N_8851,N_5976);
or UO_881 (O_881,N_6173,N_5789);
nor UO_882 (O_882,N_6148,N_5727);
or UO_883 (O_883,N_6322,N_9489);
or UO_884 (O_884,N_5415,N_5031);
xor UO_885 (O_885,N_8471,N_7185);
nand UO_886 (O_886,N_7322,N_6847);
xor UO_887 (O_887,N_5356,N_6359);
or UO_888 (O_888,N_9960,N_6701);
nand UO_889 (O_889,N_6409,N_5833);
nor UO_890 (O_890,N_6472,N_8038);
or UO_891 (O_891,N_6992,N_7594);
and UO_892 (O_892,N_8027,N_6386);
nor UO_893 (O_893,N_5549,N_6023);
xnor UO_894 (O_894,N_8935,N_9855);
or UO_895 (O_895,N_8154,N_7140);
xnor UO_896 (O_896,N_8442,N_9067);
or UO_897 (O_897,N_5754,N_9518);
nand UO_898 (O_898,N_8640,N_8268);
nand UO_899 (O_899,N_8004,N_8767);
nand UO_900 (O_900,N_6944,N_6490);
xnor UO_901 (O_901,N_7513,N_8052);
or UO_902 (O_902,N_7232,N_5297);
nor UO_903 (O_903,N_7536,N_9740);
nand UO_904 (O_904,N_5555,N_8216);
nand UO_905 (O_905,N_6587,N_6422);
or UO_906 (O_906,N_5780,N_7252);
nor UO_907 (O_907,N_5218,N_5376);
and UO_908 (O_908,N_9599,N_9958);
nor UO_909 (O_909,N_9327,N_5433);
or UO_910 (O_910,N_7046,N_5347);
nor UO_911 (O_911,N_8011,N_8447);
xnor UO_912 (O_912,N_8090,N_8262);
or UO_913 (O_913,N_6027,N_9512);
nor UO_914 (O_914,N_7916,N_9669);
and UO_915 (O_915,N_5278,N_5499);
or UO_916 (O_916,N_5043,N_9619);
xnor UO_917 (O_917,N_8238,N_8879);
and UO_918 (O_918,N_6421,N_8736);
xor UO_919 (O_919,N_5508,N_8496);
xor UO_920 (O_920,N_9472,N_6149);
nand UO_921 (O_921,N_5161,N_7732);
nor UO_922 (O_922,N_6335,N_8691);
and UO_923 (O_923,N_5543,N_6146);
nor UO_924 (O_924,N_7668,N_7728);
and UO_925 (O_925,N_7707,N_8869);
nand UO_926 (O_926,N_7869,N_9597);
and UO_927 (O_927,N_8776,N_6199);
nand UO_928 (O_928,N_8096,N_6269);
and UO_929 (O_929,N_8450,N_6029);
nand UO_930 (O_930,N_9847,N_6710);
and UO_931 (O_931,N_8371,N_9383);
and UO_932 (O_932,N_9971,N_8936);
nor UO_933 (O_933,N_5774,N_9862);
or UO_934 (O_934,N_5600,N_9978);
or UO_935 (O_935,N_6390,N_8183);
or UO_936 (O_936,N_5090,N_7084);
nor UO_937 (O_937,N_9593,N_6633);
and UO_938 (O_938,N_5146,N_6708);
nand UO_939 (O_939,N_5340,N_6757);
and UO_940 (O_940,N_6867,N_6828);
or UO_941 (O_941,N_7258,N_6423);
nand UO_942 (O_942,N_8901,N_7374);
nand UO_943 (O_943,N_9791,N_8661);
xnor UO_944 (O_944,N_7735,N_5067);
nand UO_945 (O_945,N_8717,N_7061);
or UO_946 (O_946,N_6209,N_6553);
xnor UO_947 (O_947,N_9806,N_6813);
nor UO_948 (O_948,N_9793,N_5503);
nand UO_949 (O_949,N_7924,N_6655);
nand UO_950 (O_950,N_6321,N_9389);
and UO_951 (O_951,N_5329,N_6159);
xnor UO_952 (O_952,N_6346,N_7004);
and UO_953 (O_953,N_5620,N_6062);
nor UO_954 (O_954,N_8474,N_6652);
xnor UO_955 (O_955,N_9616,N_8277);
or UO_956 (O_956,N_6431,N_5350);
or UO_957 (O_957,N_7540,N_7005);
nor UO_958 (O_958,N_6610,N_5991);
and UO_959 (O_959,N_6214,N_8668);
or UO_960 (O_960,N_6226,N_5656);
nand UO_961 (O_961,N_7901,N_7516);
nand UO_962 (O_962,N_5582,N_6740);
and UO_963 (O_963,N_7779,N_5452);
nand UO_964 (O_964,N_7995,N_7059);
nand UO_965 (O_965,N_9541,N_8644);
or UO_966 (O_966,N_9778,N_6358);
or UO_967 (O_967,N_9864,N_6546);
nand UO_968 (O_968,N_8334,N_7776);
nand UO_969 (O_969,N_9996,N_6827);
and UO_970 (O_970,N_6039,N_6378);
nor UO_971 (O_971,N_5512,N_9278);
or UO_972 (O_972,N_5708,N_9721);
nor UO_973 (O_973,N_8416,N_8321);
xor UO_974 (O_974,N_5920,N_9589);
or UO_975 (O_975,N_6900,N_7787);
nor UO_976 (O_976,N_5826,N_6225);
and UO_977 (O_977,N_6244,N_6747);
or UO_978 (O_978,N_8362,N_9034);
and UO_979 (O_979,N_9559,N_7439);
and UO_980 (O_980,N_5088,N_5012);
xor UO_981 (O_981,N_8431,N_8211);
nor UO_982 (O_982,N_9338,N_8194);
nand UO_983 (O_983,N_9647,N_9714);
nand UO_984 (O_984,N_9442,N_7993);
nand UO_985 (O_985,N_5168,N_5323);
nand UO_986 (O_986,N_9447,N_5829);
nor UO_987 (O_987,N_7035,N_6237);
nand UO_988 (O_988,N_9202,N_5316);
xor UO_989 (O_989,N_6401,N_9071);
or UO_990 (O_990,N_7873,N_9556);
and UO_991 (O_991,N_8201,N_9262);
nor UO_992 (O_992,N_5712,N_5369);
xnor UO_993 (O_993,N_9883,N_8487);
and UO_994 (O_994,N_6651,N_5674);
nand UO_995 (O_995,N_8607,N_7338);
and UO_996 (O_996,N_9623,N_8304);
and UO_997 (O_997,N_5267,N_6959);
xnor UO_998 (O_998,N_5147,N_9226);
nand UO_999 (O_999,N_8253,N_7420);
nor UO_1000 (O_1000,N_7396,N_5068);
or UO_1001 (O_1001,N_7849,N_6630);
nand UO_1002 (O_1002,N_6307,N_8367);
nor UO_1003 (O_1003,N_8484,N_6450);
nor UO_1004 (O_1004,N_8682,N_5918);
and UO_1005 (O_1005,N_7569,N_7910);
nand UO_1006 (O_1006,N_8539,N_6058);
and UO_1007 (O_1007,N_8913,N_9023);
xor UO_1008 (O_1008,N_5802,N_6932);
nor UO_1009 (O_1009,N_7254,N_8311);
or UO_1010 (O_1010,N_8423,N_8234);
or UO_1011 (O_1011,N_7815,N_8941);
or UO_1012 (O_1012,N_5495,N_8625);
xnor UO_1013 (O_1013,N_5985,N_9366);
or UO_1014 (O_1014,N_5556,N_7697);
nor UO_1015 (O_1015,N_7486,N_6719);
or UO_1016 (O_1016,N_5778,N_6891);
or UO_1017 (O_1017,N_5813,N_7933);
nor UO_1018 (O_1018,N_9934,N_5402);
and UO_1019 (O_1019,N_9179,N_6473);
or UO_1020 (O_1020,N_7880,N_8840);
and UO_1021 (O_1021,N_6262,N_9608);
nor UO_1022 (O_1022,N_5597,N_8039);
nor UO_1023 (O_1023,N_5990,N_7375);
nand UO_1024 (O_1024,N_7329,N_5983);
nor UO_1025 (O_1025,N_5014,N_8407);
or UO_1026 (O_1026,N_5263,N_9022);
and UO_1027 (O_1027,N_9190,N_8559);
nand UO_1028 (O_1028,N_7056,N_5405);
and UO_1029 (O_1029,N_5926,N_7762);
and UO_1030 (O_1030,N_9103,N_7900);
and UO_1031 (O_1031,N_6650,N_8137);
and UO_1032 (O_1032,N_5446,N_6497);
or UO_1033 (O_1033,N_7527,N_5154);
nand UO_1034 (O_1034,N_5211,N_8408);
and UO_1035 (O_1035,N_7264,N_7268);
xor UO_1036 (O_1036,N_5891,N_7945);
nor UO_1037 (O_1037,N_8032,N_6389);
and UO_1038 (O_1038,N_7450,N_5314);
xnor UO_1039 (O_1039,N_7704,N_5388);
and UO_1040 (O_1040,N_6008,N_8110);
or UO_1041 (O_1041,N_7147,N_6792);
nand UO_1042 (O_1042,N_6543,N_7160);
and UO_1043 (O_1043,N_9204,N_7925);
nand UO_1044 (O_1044,N_6722,N_9146);
nand UO_1045 (O_1045,N_7152,N_7928);
and UO_1046 (O_1046,N_6554,N_6223);
or UO_1047 (O_1047,N_9141,N_7053);
nand UO_1048 (O_1048,N_5457,N_5167);
or UO_1049 (O_1049,N_5165,N_6365);
nor UO_1050 (O_1050,N_5417,N_6320);
nor UO_1051 (O_1051,N_6577,N_9275);
or UO_1052 (O_1052,N_7249,N_8095);
and UO_1053 (O_1053,N_9231,N_5518);
or UO_1054 (O_1054,N_5050,N_9099);
or UO_1055 (O_1055,N_6826,N_9432);
or UO_1056 (O_1056,N_5203,N_6379);
or UO_1057 (O_1057,N_7974,N_5626);
or UO_1058 (O_1058,N_7212,N_5887);
or UO_1059 (O_1059,N_7523,N_5256);
nand UO_1060 (O_1060,N_7989,N_9109);
nand UO_1061 (O_1061,N_6157,N_5344);
and UO_1062 (O_1062,N_8792,N_8001);
and UO_1063 (O_1063,N_6835,N_9652);
and UO_1064 (O_1064,N_5155,N_7038);
xnor UO_1065 (O_1065,N_9712,N_9282);
nor UO_1066 (O_1066,N_5041,N_6086);
nand UO_1067 (O_1067,N_5429,N_7100);
nand UO_1068 (O_1068,N_6011,N_6859);
nand UO_1069 (O_1069,N_8021,N_5741);
or UO_1070 (O_1070,N_7178,N_8161);
nand UO_1071 (O_1071,N_5903,N_6581);
nand UO_1072 (O_1072,N_9948,N_8704);
nor UO_1073 (O_1073,N_9728,N_8190);
or UO_1074 (O_1074,N_7478,N_7737);
or UO_1075 (O_1075,N_6236,N_9374);
nand UO_1076 (O_1076,N_8354,N_8375);
nor UO_1077 (O_1077,N_7994,N_6270);
nor UO_1078 (O_1078,N_5206,N_7850);
nand UO_1079 (O_1079,N_7851,N_9537);
nor UO_1080 (O_1080,N_9161,N_7432);
or UO_1081 (O_1081,N_6477,N_8085);
or UO_1082 (O_1082,N_8746,N_9239);
nand UO_1083 (O_1083,N_9703,N_7578);
nor UO_1084 (O_1084,N_9271,N_6104);
nand UO_1085 (O_1085,N_6530,N_6107);
and UO_1086 (O_1086,N_6103,N_6463);
xnor UO_1087 (O_1087,N_5111,N_6328);
nand UO_1088 (O_1088,N_8357,N_7805);
nand UO_1089 (O_1089,N_6398,N_5410);
nor UO_1090 (O_1090,N_6877,N_8105);
or UO_1091 (O_1091,N_6724,N_7347);
or UO_1092 (O_1092,N_5262,N_8119);
nand UO_1093 (O_1093,N_5640,N_5671);
and UO_1094 (O_1094,N_5136,N_7484);
or UO_1095 (O_1095,N_9663,N_8729);
and UO_1096 (O_1096,N_5834,N_8123);
or UO_1097 (O_1097,N_8470,N_8395);
and UO_1098 (O_1098,N_6780,N_9425);
nand UO_1099 (O_1099,N_5694,N_8787);
nand UO_1100 (O_1100,N_8923,N_5804);
nand UO_1101 (O_1101,N_5890,N_8847);
and UO_1102 (O_1102,N_6648,N_5006);
xor UO_1103 (O_1103,N_5299,N_5579);
nor UO_1104 (O_1104,N_7209,N_6799);
and UO_1105 (O_1105,N_5882,N_7190);
or UO_1106 (O_1106,N_5643,N_8914);
nor UO_1107 (O_1107,N_7555,N_7981);
or UO_1108 (O_1108,N_9386,N_7801);
nand UO_1109 (O_1109,N_6742,N_9433);
xnor UO_1110 (O_1110,N_8280,N_6181);
and UO_1111 (O_1111,N_6593,N_6804);
nand UO_1112 (O_1112,N_8246,N_8745);
or UO_1113 (O_1113,N_6989,N_7119);
and UO_1114 (O_1114,N_9010,N_6883);
or UO_1115 (O_1115,N_9921,N_6861);
nand UO_1116 (O_1116,N_9888,N_9404);
xor UO_1117 (O_1117,N_8411,N_7188);
xnor UO_1118 (O_1118,N_6147,N_7999);
xor UO_1119 (O_1119,N_8844,N_7315);
nor UO_1120 (O_1120,N_7317,N_8492);
xor UO_1121 (O_1121,N_6578,N_8300);
nor UO_1122 (O_1122,N_9788,N_6433);
xor UO_1123 (O_1123,N_5949,N_6400);
and UO_1124 (O_1124,N_9694,N_7604);
or UO_1125 (O_1125,N_9000,N_9351);
nor UO_1126 (O_1126,N_8855,N_5901);
nand UO_1127 (O_1127,N_6653,N_7550);
nor UO_1128 (O_1128,N_9636,N_6893);
and UO_1129 (O_1129,N_6519,N_7237);
and UO_1130 (O_1130,N_9205,N_5726);
nand UO_1131 (O_1131,N_8325,N_6943);
nor UO_1132 (O_1132,N_7684,N_6783);
nand UO_1133 (O_1133,N_7716,N_6584);
and UO_1134 (O_1134,N_8870,N_6260);
or UO_1135 (O_1135,N_6641,N_7141);
nor UO_1136 (O_1136,N_9112,N_9400);
or UO_1137 (O_1137,N_5667,N_9982);
nand UO_1138 (O_1138,N_5431,N_9724);
nand UO_1139 (O_1139,N_9592,N_8187);
nand UO_1140 (O_1140,N_7354,N_6715);
and UO_1141 (O_1141,N_8402,N_5274);
or UO_1142 (O_1142,N_7715,N_9953);
nand UO_1143 (O_1143,N_7300,N_8738);
nor UO_1144 (O_1144,N_5258,N_5471);
nand UO_1145 (O_1145,N_9881,N_5202);
nor UO_1146 (O_1146,N_8328,N_5177);
xnor UO_1147 (O_1147,N_8678,N_7821);
xor UO_1148 (O_1148,N_6695,N_6121);
and UO_1149 (O_1149,N_8338,N_6875);
and UO_1150 (O_1150,N_6382,N_8953);
nor UO_1151 (O_1151,N_5740,N_6316);
nor UO_1152 (O_1152,N_6143,N_8109);
nand UO_1153 (O_1153,N_6602,N_7829);
xnor UO_1154 (O_1154,N_5587,N_9893);
or UO_1155 (O_1155,N_5328,N_5678);
nor UO_1156 (O_1156,N_8593,N_5093);
and UO_1157 (O_1157,N_6026,N_8306);
or UO_1158 (O_1158,N_8219,N_7469);
nand UO_1159 (O_1159,N_7368,N_6733);
and UO_1160 (O_1160,N_7461,N_8320);
nor UO_1161 (O_1161,N_9633,N_9199);
and UO_1162 (O_1162,N_9696,N_6087);
xnor UO_1163 (O_1163,N_9622,N_9256);
and UO_1164 (O_1164,N_5260,N_9055);
nor UO_1165 (O_1165,N_6255,N_9901);
or UO_1166 (O_1166,N_5193,N_8452);
and UO_1167 (O_1167,N_7395,N_9310);
nor UO_1168 (O_1168,N_8479,N_5974);
nand UO_1169 (O_1169,N_7975,N_6333);
and UO_1170 (O_1170,N_9170,N_9352);
or UO_1171 (O_1171,N_5238,N_7226);
nor UO_1172 (O_1172,N_8774,N_7039);
nor UO_1173 (O_1173,N_5372,N_9908);
nor UO_1174 (O_1174,N_8477,N_8815);
or UO_1175 (O_1175,N_8558,N_5239);
and UO_1176 (O_1176,N_8771,N_6429);
or UO_1177 (O_1177,N_6405,N_5822);
or UO_1178 (O_1178,N_9244,N_5733);
nor UO_1179 (O_1179,N_8139,N_9163);
or UO_1180 (O_1180,N_6048,N_9984);
and UO_1181 (O_1181,N_7935,N_8885);
or UO_1182 (O_1182,N_8622,N_8390);
or UO_1183 (O_1183,N_6656,N_5684);
and UO_1184 (O_1184,N_7912,N_9390);
and UO_1185 (O_1185,N_6078,N_8929);
and UO_1186 (O_1186,N_9206,N_9450);
nor UO_1187 (O_1187,N_7984,N_9641);
and UO_1188 (O_1188,N_6334,N_5075);
nor UO_1189 (O_1189,N_7588,N_8519);
xnor UO_1190 (O_1190,N_6092,N_7093);
xor UO_1191 (O_1191,N_6632,N_8072);
nand UO_1192 (O_1192,N_6326,N_9078);
or UO_1193 (O_1193,N_5645,N_5544);
nand UO_1194 (O_1194,N_6853,N_5339);
xor UO_1195 (O_1195,N_8572,N_6387);
nand UO_1196 (O_1196,N_8014,N_6823);
or UO_1197 (O_1197,N_5485,N_8048);
or UO_1198 (O_1198,N_6594,N_8676);
or UO_1199 (O_1199,N_9667,N_8780);
and UO_1200 (O_1200,N_5531,N_5001);
nand UO_1201 (O_1201,N_6360,N_6961);
and UO_1202 (O_1202,N_8068,N_8666);
nor UO_1203 (O_1203,N_9360,N_9548);
nand UO_1204 (O_1204,N_8854,N_8857);
and UO_1205 (O_1205,N_7990,N_7894);
and UO_1206 (O_1206,N_5060,N_7884);
nand UO_1207 (O_1207,N_7060,N_7661);
nor UO_1208 (O_1208,N_6535,N_7764);
or UO_1209 (O_1209,N_6966,N_8679);
nor UO_1210 (O_1210,N_6294,N_5424);
or UO_1211 (O_1211,N_6195,N_8288);
nand UO_1212 (O_1212,N_6575,N_5456);
and UO_1213 (O_1213,N_9171,N_9858);
or UO_1214 (O_1214,N_5883,N_7026);
nand UO_1215 (O_1215,N_9091,N_8312);
nor UO_1216 (O_1216,N_9434,N_7036);
xor UO_1217 (O_1217,N_9812,N_6388);
nand UO_1218 (O_1218,N_7387,N_9426);
nand UO_1219 (O_1219,N_6488,N_9841);
or UO_1220 (O_1220,N_9611,N_7112);
nor UO_1221 (O_1221,N_5460,N_5965);
nand UO_1222 (O_1222,N_5156,N_6760);
nand UO_1223 (O_1223,N_8515,N_5619);
nor UO_1224 (O_1224,N_7092,N_7739);
and UO_1225 (O_1225,N_8460,N_6865);
and UO_1226 (O_1226,N_9553,N_5036);
nand UO_1227 (O_1227,N_5633,N_8884);
nor UO_1228 (O_1228,N_9523,N_9944);
or UO_1229 (O_1229,N_8754,N_6682);
or UO_1230 (O_1230,N_9547,N_5019);
or UO_1231 (O_1231,N_6056,N_9136);
nand UO_1232 (O_1232,N_9874,N_6352);
or UO_1233 (O_1233,N_9880,N_6685);
nand UO_1234 (O_1234,N_6203,N_5049);
or UO_1235 (O_1235,N_7724,N_9674);
and UO_1236 (O_1236,N_9912,N_9047);
nor UO_1237 (O_1237,N_8830,N_5994);
or UO_1238 (O_1238,N_9821,N_5265);
and UO_1239 (O_1239,N_5529,N_6112);
or UO_1240 (O_1240,N_6607,N_5505);
nor UO_1241 (O_1241,N_5659,N_8744);
and UO_1242 (O_1242,N_9808,N_9184);
nor UO_1243 (O_1243,N_8820,N_7498);
and UO_1244 (O_1244,N_5535,N_6982);
nor UO_1245 (O_1245,N_8809,N_6021);
or UO_1246 (O_1246,N_5841,N_9125);
or UO_1247 (O_1247,N_5282,N_6182);
nand UO_1248 (O_1248,N_8029,N_8547);
nor UO_1249 (O_1249,N_7970,N_7400);
nor UO_1250 (O_1250,N_8656,N_8790);
and UO_1251 (O_1251,N_8872,N_5103);
nand UO_1252 (O_1252,N_7105,N_7978);
nor UO_1253 (O_1253,N_6392,N_8555);
nor UO_1254 (O_1254,N_9021,N_8662);
and UO_1255 (O_1255,N_8897,N_7803);
nand UO_1256 (O_1256,N_8019,N_8056);
nand UO_1257 (O_1257,N_6988,N_7943);
nor UO_1258 (O_1258,N_5772,N_8763);
nand UO_1259 (O_1259,N_7814,N_9451);
nand UO_1260 (O_1260,N_6562,N_7032);
or UO_1261 (O_1261,N_6597,N_6446);
or UO_1262 (O_1262,N_7950,N_8124);
and UO_1263 (O_1263,N_7231,N_8993);
nand UO_1264 (O_1264,N_8985,N_9834);
or UO_1265 (O_1265,N_8802,N_5707);
and UO_1266 (O_1266,N_8975,N_8987);
or UO_1267 (O_1267,N_7292,N_8866);
nor UO_1268 (O_1268,N_5836,N_6789);
xnor UO_1269 (O_1269,N_7750,N_8380);
and UO_1270 (O_1270,N_9759,N_6855);
nor UO_1271 (O_1271,N_5209,N_9699);
or UO_1272 (O_1272,N_6808,N_5483);
nand UO_1273 (O_1273,N_7435,N_9532);
nand UO_1274 (O_1274,N_7657,N_7410);
nor UO_1275 (O_1275,N_6930,N_9900);
nand UO_1276 (O_1276,N_6896,N_8281);
nand UO_1277 (O_1277,N_9182,N_5574);
nand UO_1278 (O_1278,N_5762,N_9690);
xnor UO_1279 (O_1279,N_7629,N_5300);
and UO_1280 (O_1280,N_6169,N_5807);
or UO_1281 (O_1281,N_9027,N_8587);
nor UO_1282 (O_1282,N_9189,N_5322);
and UO_1283 (O_1283,N_8590,N_5580);
nand UO_1284 (O_1284,N_5962,N_7509);
or UO_1285 (O_1285,N_6364,N_8317);
nand UO_1286 (O_1286,N_7029,N_5489);
nor UO_1287 (O_1287,N_5915,N_5724);
or UO_1288 (O_1288,N_5624,N_8740);
nand UO_1289 (O_1289,N_9943,N_6356);
or UO_1290 (O_1290,N_8180,N_7611);
nor UO_1291 (O_1291,N_6570,N_8861);
nand UO_1292 (O_1292,N_7520,N_6125);
or UO_1293 (O_1293,N_9063,N_5825);
and UO_1294 (O_1294,N_5909,N_7768);
xor UO_1295 (O_1295,N_7507,N_6075);
nor UO_1296 (O_1296,N_7380,N_7344);
nand UO_1297 (O_1297,N_8054,N_8155);
or UO_1298 (O_1298,N_6667,N_7390);
and UO_1299 (O_1299,N_9250,N_5397);
nor UO_1300 (O_1300,N_6545,N_8735);
nand UO_1301 (O_1301,N_8697,N_6729);
or UO_1302 (O_1302,N_9895,N_9230);
or UO_1303 (O_1303,N_8612,N_6759);
nor UO_1304 (O_1304,N_8991,N_8260);
nand UO_1305 (O_1305,N_8853,N_7552);
or UO_1306 (O_1306,N_8796,N_9664);
nor UO_1307 (O_1307,N_7337,N_7681);
nor UO_1308 (O_1308,N_7427,N_6840);
nand UO_1309 (O_1309,N_7255,N_5273);
and UO_1310 (O_1310,N_6874,N_8716);
nand UO_1311 (O_1311,N_9065,N_9144);
or UO_1312 (O_1312,N_6325,N_9315);
xor UO_1313 (O_1313,N_5864,N_5525);
nor UO_1314 (O_1314,N_7532,N_7075);
nor UO_1315 (O_1315,N_5998,N_8723);
and UO_1316 (O_1316,N_9683,N_7658);
nor UO_1317 (O_1317,N_8569,N_6057);
or UO_1318 (O_1318,N_6830,N_5257);
or UO_1319 (O_1319,N_9342,N_6940);
or UO_1320 (O_1320,N_7962,N_9991);
nor UO_1321 (O_1321,N_6972,N_5020);
nand UO_1322 (O_1322,N_8990,N_9554);
xor UO_1323 (O_1323,N_7054,N_7747);
nor UO_1324 (O_1324,N_7238,N_9500);
nor UO_1325 (O_1325,N_5310,N_6410);
nor UO_1326 (O_1326,N_9015,N_5950);
nand UO_1327 (O_1327,N_9155,N_5793);
and UO_1328 (O_1328,N_8831,N_6777);
xor UO_1329 (O_1329,N_7804,N_5576);
and UO_1330 (O_1330,N_8812,N_5977);
or UO_1331 (O_1331,N_5158,N_8600);
or UO_1332 (O_1332,N_9941,N_7162);
nor UO_1333 (O_1333,N_8672,N_6664);
and UO_1334 (O_1334,N_5840,N_6015);
nor UO_1335 (O_1335,N_8017,N_8643);
nand UO_1336 (O_1336,N_5787,N_6666);
nor UO_1337 (O_1337,N_5380,N_9911);
and UO_1338 (O_1338,N_5561,N_7874);
or UO_1339 (O_1339,N_8525,N_9090);
xnor UO_1340 (O_1340,N_8918,N_5408);
nor UO_1341 (O_1341,N_7695,N_7379);
and UO_1342 (O_1342,N_9870,N_8167);
nor UO_1343 (O_1343,N_7442,N_9933);
or UO_1344 (O_1344,N_9212,N_7769);
nor UO_1345 (O_1345,N_5061,N_6280);
nand UO_1346 (O_1346,N_6286,N_9860);
xnor UO_1347 (O_1347,N_6937,N_7923);
or UO_1348 (O_1348,N_5784,N_5205);
nor UO_1349 (O_1349,N_5224,N_7335);
and UO_1350 (O_1350,N_5264,N_6501);
and UO_1351 (O_1351,N_8526,N_5837);
nand UO_1352 (O_1352,N_8748,N_9739);
nor UO_1353 (O_1353,N_9481,N_6773);
nand UO_1354 (O_1354,N_9634,N_8817);
nor UO_1355 (O_1355,N_7286,N_9110);
nor UO_1356 (O_1356,N_7000,N_5691);
and UO_1357 (O_1357,N_6670,N_8307);
nor UO_1358 (O_1358,N_5646,N_9221);
xnor UO_1359 (O_1359,N_6250,N_9995);
nor UO_1360 (O_1360,N_8324,N_6179);
and UO_1361 (O_1361,N_8145,N_7012);
and UO_1362 (O_1362,N_8690,N_9356);
nor UO_1363 (O_1363,N_5668,N_5449);
nand UO_1364 (O_1364,N_7082,N_9030);
and UO_1365 (O_1365,N_6686,N_5437);
nor UO_1366 (O_1366,N_7325,N_7353);
xnor UO_1367 (O_1367,N_8003,N_9188);
nand UO_1368 (O_1368,N_8232,N_7393);
and UO_1369 (O_1369,N_9628,N_8398);
or UO_1370 (O_1370,N_6565,N_7165);
and UO_1371 (O_1371,N_6124,N_5109);
and UO_1372 (O_1372,N_9961,N_7219);
and UO_1373 (O_1373,N_8848,N_7590);
or UO_1374 (O_1374,N_6291,N_5450);
and UO_1375 (O_1375,N_6866,N_9143);
nand UO_1376 (O_1376,N_6784,N_8952);
and UO_1377 (O_1377,N_9892,N_8688);
nand UO_1378 (O_1378,N_5714,N_8432);
nand UO_1379 (O_1379,N_6600,N_7679);
nor UO_1380 (O_1380,N_5253,N_7148);
nor UO_1381 (O_1381,N_5557,N_7333);
or UO_1382 (O_1382,N_9436,N_5849);
or UO_1383 (O_1383,N_6186,N_5131);
xor UO_1384 (O_1384,N_9439,N_9183);
or UO_1385 (O_1385,N_5736,N_7606);
nand UO_1386 (O_1386,N_7653,N_5106);
nor UO_1387 (O_1387,N_5010,N_5967);
nand UO_1388 (O_1388,N_6498,N_8283);
and UO_1389 (O_1389,N_6257,N_8911);
or UO_1390 (O_1390,N_7895,N_9227);
and UO_1391 (O_1391,N_7688,N_6538);
nor UO_1392 (O_1392,N_6627,N_8441);
or UO_1393 (O_1393,N_8915,N_5059);
nor UO_1394 (O_1394,N_6177,N_5494);
nor UO_1395 (O_1395,N_6065,N_8724);
xor UO_1396 (O_1396,N_5634,N_7130);
nor UO_1397 (O_1397,N_8883,N_8998);
nor UO_1398 (O_1398,N_9757,N_9818);
nand UO_1399 (O_1399,N_9251,N_6756);
nand UO_1400 (O_1400,N_6310,N_6899);
or UO_1401 (O_1401,N_8116,N_8720);
and UO_1402 (O_1402,N_5002,N_9675);
nand UO_1403 (O_1403,N_7192,N_7101);
or UO_1404 (O_1404,N_7580,N_6156);
nand UO_1405 (O_1405,N_6579,N_8732);
or UO_1406 (O_1406,N_9038,N_7650);
nand UO_1407 (O_1407,N_7128,N_7169);
nand UO_1408 (O_1408,N_7403,N_6735);
nand UO_1409 (O_1409,N_5164,N_9613);
and UO_1410 (O_1410,N_9246,N_9044);
nand UO_1411 (O_1411,N_5004,N_8629);
nand UO_1412 (O_1412,N_8217,N_8522);
nor UO_1413 (O_1413,N_7749,N_8645);
nand UO_1414 (O_1414,N_6851,N_8443);
or UO_1415 (O_1415,N_7835,N_6371);
nor UO_1416 (O_1416,N_5395,N_7073);
and UO_1417 (O_1417,N_6942,N_9375);
xnor UO_1418 (O_1418,N_6258,N_6764);
or UO_1419 (O_1419,N_5305,N_5057);
or UO_1420 (O_1420,N_6222,N_9307);
nand UO_1421 (O_1421,N_5982,N_6469);
nor UO_1422 (O_1422,N_5121,N_9705);
xor UO_1423 (O_1423,N_8179,N_7384);
and UO_1424 (O_1424,N_8677,N_7544);
nand UO_1425 (O_1425,N_5022,N_8829);
nor UO_1426 (O_1426,N_8906,N_5018);
and UO_1427 (O_1427,N_8635,N_6201);
xor UO_1428 (O_1428,N_8094,N_7404);
or UO_1429 (O_1429,N_6355,N_5639);
nor UO_1430 (O_1430,N_6068,N_5003);
and UO_1431 (O_1431,N_7666,N_5606);
and UO_1432 (O_1432,N_6920,N_8646);
nand UO_1433 (O_1433,N_9252,N_8308);
or UO_1434 (O_1434,N_7833,N_9054);
nor UO_1435 (O_1435,N_8401,N_6004);
nor UO_1436 (O_1436,N_9591,N_7876);
and UO_1437 (O_1437,N_6313,N_8218);
xnor UO_1438 (O_1438,N_5332,N_7620);
nor UO_1439 (O_1439,N_7938,N_6863);
xor UO_1440 (O_1440,N_8896,N_8804);
nor UO_1441 (O_1441,N_9904,N_9981);
and UO_1442 (O_1442,N_9977,N_6340);
or UO_1443 (O_1443,N_5929,N_5563);
xor UO_1444 (O_1444,N_6164,N_5364);
or UO_1445 (O_1445,N_8706,N_5324);
and UO_1446 (O_1446,N_6697,N_6289);
nor UO_1447 (O_1447,N_7330,N_8582);
nand UO_1448 (O_1448,N_7859,N_9502);
nor UO_1449 (O_1449,N_9606,N_5272);
and UO_1450 (O_1450,N_9385,N_6517);
nor UO_1451 (O_1451,N_6540,N_8257);
nor UO_1452 (O_1452,N_9323,N_9529);
nand UO_1453 (O_1453,N_5775,N_6158);
or UO_1454 (O_1454,N_9220,N_7672);
and UO_1455 (O_1455,N_8788,N_9138);
or UO_1456 (O_1456,N_6090,N_9280);
nor UO_1457 (O_1457,N_7772,N_6752);
nor UO_1458 (O_1458,N_8819,N_7455);
nor UO_1459 (O_1459,N_7759,N_6344);
nand UO_1460 (O_1460,N_8069,N_9213);
nor UO_1461 (O_1461,N_9429,N_9546);
and UO_1462 (O_1462,N_5867,N_9314);
nand UO_1463 (O_1463,N_7517,N_7198);
and UO_1464 (O_1464,N_7683,N_5011);
and UO_1465 (O_1465,N_8972,N_5958);
nand UO_1466 (O_1466,N_9427,N_6672);
and UO_1467 (O_1467,N_9802,N_7637);
xor UO_1468 (O_1468,N_8655,N_5722);
nand UO_1469 (O_1469,N_8674,N_7545);
nor UO_1470 (O_1470,N_5076,N_9837);
nor UO_1471 (O_1471,N_8276,N_9210);
nand UO_1472 (O_1472,N_5444,N_5608);
nor UO_1473 (O_1473,N_7963,N_7641);
and UO_1474 (O_1474,N_9381,N_7177);
nand UO_1475 (O_1475,N_6880,N_7720);
or UO_1476 (O_1476,N_8687,N_6187);
nand UO_1477 (O_1477,N_7774,N_7441);
nor UO_1478 (O_1478,N_7066,N_6080);
xor UO_1479 (O_1479,N_9482,N_5510);
or UO_1480 (O_1480,N_5176,N_6123);
or UO_1481 (O_1481,N_5191,N_8766);
and UO_1482 (O_1482,N_6110,N_7510);
xor UO_1483 (O_1483,N_6414,N_5986);
or UO_1484 (O_1484,N_7624,N_9005);
and UO_1485 (O_1485,N_9483,N_5889);
xnor UO_1486 (O_1486,N_8393,N_6503);
xor UO_1487 (O_1487,N_6275,N_9831);
or UO_1488 (O_1488,N_5387,N_9474);
or UO_1489 (O_1489,N_8480,N_7423);
or UO_1490 (O_1490,N_8250,N_7274);
nor UO_1491 (O_1491,N_9820,N_7856);
and UO_1492 (O_1492,N_8097,N_6507);
nand UO_1493 (O_1493,N_6273,N_5617);
nand UO_1494 (O_1494,N_8413,N_7343);
and UO_1495 (O_1495,N_8733,N_7717);
or UO_1496 (O_1496,N_8373,N_7473);
nand UO_1497 (O_1497,N_9225,N_9749);
nor UO_1498 (O_1498,N_9886,N_9771);
nor UO_1499 (O_1499,N_8843,N_9348);
endmodule