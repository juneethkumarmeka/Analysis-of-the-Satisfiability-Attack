module basic_500_3000_500_15_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_199,In_186);
nand U1 (N_1,In_53,In_216);
or U2 (N_2,In_436,In_8);
nor U3 (N_3,In_138,In_289);
or U4 (N_4,In_373,In_204);
nor U5 (N_5,In_153,In_272);
nand U6 (N_6,In_476,In_181);
xnor U7 (N_7,In_228,In_420);
nor U8 (N_8,In_238,In_350);
or U9 (N_9,In_466,In_191);
and U10 (N_10,In_312,In_237);
and U11 (N_11,In_308,In_88);
nor U12 (N_12,In_254,In_14);
and U13 (N_13,In_295,In_323);
and U14 (N_14,In_86,In_257);
nor U15 (N_15,In_221,In_335);
nand U16 (N_16,In_403,In_61);
and U17 (N_17,In_177,In_215);
or U18 (N_18,In_438,In_42);
nand U19 (N_19,In_4,In_443);
xor U20 (N_20,In_28,In_454);
and U21 (N_21,In_102,In_149);
or U22 (N_22,In_366,In_266);
and U23 (N_23,In_162,In_133);
or U24 (N_24,In_161,In_406);
nand U25 (N_25,In_348,In_437);
nand U26 (N_26,In_417,In_452);
or U27 (N_27,In_176,In_194);
nor U28 (N_28,In_64,In_368);
or U29 (N_29,In_371,In_79);
nor U30 (N_30,In_74,In_475);
xnor U31 (N_31,In_93,In_392);
nand U32 (N_32,In_48,In_387);
xor U33 (N_33,In_151,In_72);
xor U34 (N_34,In_0,In_372);
xnor U35 (N_35,In_448,In_426);
or U36 (N_36,In_369,In_262);
and U37 (N_37,In_214,In_330);
or U38 (N_38,In_418,In_255);
nor U39 (N_39,In_349,In_124);
and U40 (N_40,In_139,In_423);
xor U41 (N_41,In_351,In_467);
nor U42 (N_42,In_311,In_44);
nor U43 (N_43,In_122,In_10);
or U44 (N_44,In_140,In_391);
xor U45 (N_45,In_20,In_337);
or U46 (N_46,In_256,In_469);
nor U47 (N_47,In_52,In_267);
or U48 (N_48,In_419,In_491);
or U49 (N_49,In_201,In_211);
xnor U50 (N_50,In_446,In_18);
nor U51 (N_51,In_333,In_1);
nand U52 (N_52,In_141,In_296);
xor U53 (N_53,In_409,In_269);
or U54 (N_54,In_261,In_229);
nor U55 (N_55,In_288,In_310);
xnor U56 (N_56,In_39,In_483);
and U57 (N_57,In_118,In_110);
or U58 (N_58,In_401,In_370);
or U59 (N_59,In_168,In_16);
and U60 (N_60,In_367,In_263);
or U61 (N_61,In_223,In_90);
and U62 (N_62,In_248,In_487);
or U63 (N_63,In_78,In_108);
or U64 (N_64,In_157,In_386);
xor U65 (N_65,In_200,In_384);
nor U66 (N_66,In_19,In_135);
xnor U67 (N_67,In_252,In_82);
nor U68 (N_68,In_111,In_481);
or U69 (N_69,In_407,In_51);
nor U70 (N_70,In_60,In_316);
or U71 (N_71,In_415,In_65);
or U72 (N_72,In_320,In_471);
nand U73 (N_73,In_318,In_359);
xnor U74 (N_74,In_66,In_94);
xnor U75 (N_75,In_499,In_291);
and U76 (N_76,In_179,In_188);
and U77 (N_77,In_245,In_395);
or U78 (N_78,In_461,In_21);
or U79 (N_79,In_101,In_339);
xor U80 (N_80,In_136,In_76);
xnor U81 (N_81,In_450,In_62);
xor U82 (N_82,In_422,In_260);
xor U83 (N_83,In_171,In_209);
nor U84 (N_84,In_128,In_159);
and U85 (N_85,In_63,In_428);
xnor U86 (N_86,In_219,In_71);
nand U87 (N_87,In_347,In_47);
nor U88 (N_88,In_217,In_435);
or U89 (N_89,In_441,In_379);
nand U90 (N_90,In_374,In_285);
or U91 (N_91,In_195,In_278);
and U92 (N_92,In_459,In_299);
and U93 (N_93,In_434,In_95);
and U94 (N_94,In_307,In_184);
xor U95 (N_95,In_105,In_125);
xor U96 (N_96,In_41,In_493);
and U97 (N_97,In_130,In_173);
and U98 (N_98,In_474,In_343);
and U99 (N_99,In_398,In_314);
xor U100 (N_100,In_489,In_45);
nor U101 (N_101,In_40,In_97);
xnor U102 (N_102,In_220,In_247);
and U103 (N_103,In_167,In_322);
nand U104 (N_104,In_99,In_77);
xor U105 (N_105,In_163,In_425);
or U106 (N_106,In_131,In_83);
nand U107 (N_107,In_399,In_146);
nand U108 (N_108,In_363,In_338);
or U109 (N_109,In_353,In_292);
and U110 (N_110,In_154,In_492);
and U111 (N_111,In_33,In_319);
nor U112 (N_112,In_43,In_210);
xor U113 (N_113,In_325,In_279);
or U114 (N_114,In_232,In_383);
xor U115 (N_115,In_54,In_123);
or U116 (N_116,In_31,In_37);
nor U117 (N_117,In_137,In_5);
and U118 (N_118,In_402,In_345);
nor U119 (N_119,In_277,In_439);
or U120 (N_120,In_429,In_119);
nand U121 (N_121,In_445,In_376);
xnor U122 (N_122,In_360,In_259);
xnor U123 (N_123,In_455,In_284);
nor U124 (N_124,In_300,In_96);
and U125 (N_125,In_282,In_462);
nor U126 (N_126,In_24,In_253);
nor U127 (N_127,In_227,In_497);
nor U128 (N_128,In_100,In_117);
nor U129 (N_129,In_241,In_30);
xor U130 (N_130,In_457,In_243);
and U131 (N_131,In_444,In_198);
nand U132 (N_132,In_341,In_364);
or U133 (N_133,In_165,In_470);
or U134 (N_134,In_283,In_104);
xor U135 (N_135,In_463,In_89);
nor U136 (N_136,In_84,In_273);
and U137 (N_137,In_116,In_327);
nor U138 (N_138,In_354,In_484);
xnor U139 (N_139,In_362,In_9);
nand U140 (N_140,In_158,In_189);
xnor U141 (N_141,In_17,In_197);
xor U142 (N_142,In_13,In_265);
xnor U143 (N_143,In_25,In_424);
and U144 (N_144,In_328,In_442);
xnor U145 (N_145,In_244,In_3);
and U146 (N_146,In_109,In_29);
xor U147 (N_147,In_495,In_212);
or U148 (N_148,In_496,In_239);
nor U149 (N_149,In_235,In_432);
nand U150 (N_150,In_98,In_485);
or U151 (N_151,In_150,In_358);
nor U152 (N_152,In_249,In_174);
or U153 (N_153,In_156,In_378);
and U154 (N_154,In_155,In_490);
xnor U155 (N_155,In_342,In_421);
nor U156 (N_156,In_275,In_482);
xor U157 (N_157,In_145,In_226);
and U158 (N_158,In_331,In_478);
or U159 (N_159,In_87,In_127);
and U160 (N_160,In_251,In_121);
nand U161 (N_161,In_207,In_166);
xor U162 (N_162,In_203,In_180);
xnor U163 (N_163,In_222,In_22);
or U164 (N_164,In_451,In_293);
xor U165 (N_165,In_479,In_202);
nor U166 (N_166,In_294,In_112);
nand U167 (N_167,In_6,In_58);
and U168 (N_168,In_23,In_144);
nand U169 (N_169,In_413,In_281);
nor U170 (N_170,In_309,In_147);
xor U171 (N_171,In_70,In_234);
nor U172 (N_172,In_393,In_356);
or U173 (N_173,In_185,In_304);
xor U174 (N_174,In_213,In_80);
xnor U175 (N_175,In_170,In_468);
xor U176 (N_176,In_225,In_405);
xor U177 (N_177,In_280,In_26);
nand U178 (N_178,In_274,In_132);
or U179 (N_179,In_134,In_175);
xor U180 (N_180,In_178,In_236);
and U181 (N_181,In_55,In_15);
xnor U182 (N_182,In_242,In_11);
and U183 (N_183,In_113,In_396);
nor U184 (N_184,In_50,In_12);
xnor U185 (N_185,In_196,In_143);
and U186 (N_186,In_91,In_306);
nand U187 (N_187,In_103,In_126);
xor U188 (N_188,In_381,In_321);
or U189 (N_189,In_460,In_488);
and U190 (N_190,In_59,In_107);
and U191 (N_191,In_164,In_187);
xnor U192 (N_192,In_447,In_38);
xnor U193 (N_193,In_301,In_240);
nor U194 (N_194,In_160,In_35);
or U195 (N_195,In_389,In_388);
nor U196 (N_196,In_286,In_303);
or U197 (N_197,In_271,In_494);
xor U198 (N_198,In_480,In_120);
or U199 (N_199,In_190,In_449);
and U200 (N_200,N_194,N_95);
xnor U201 (N_201,In_440,N_137);
nor U202 (N_202,N_68,N_170);
nor U203 (N_203,N_27,N_173);
or U204 (N_204,N_186,N_183);
nand U205 (N_205,N_19,In_313);
xor U206 (N_206,N_155,N_40);
xnor U207 (N_207,In_142,N_157);
nand U208 (N_208,N_49,In_169);
nand U209 (N_209,N_153,N_25);
nand U210 (N_210,In_290,N_181);
or U211 (N_211,N_160,In_465);
nand U212 (N_212,N_115,N_67);
or U213 (N_213,N_101,In_32);
nand U214 (N_214,In_148,N_116);
xor U215 (N_215,N_132,N_37);
nand U216 (N_216,N_79,N_3);
xnor U217 (N_217,N_80,N_171);
and U218 (N_218,N_145,N_59);
or U219 (N_219,N_6,N_131);
or U220 (N_220,N_121,In_208);
and U221 (N_221,N_70,In_412);
and U222 (N_222,In_56,N_164);
xnor U223 (N_223,In_410,N_48);
xor U224 (N_224,N_14,N_4);
nor U225 (N_225,N_129,In_377);
xor U226 (N_226,N_9,In_477);
nor U227 (N_227,In_473,N_133);
xor U228 (N_228,N_199,N_17);
nand U229 (N_229,In_129,In_464);
xnor U230 (N_230,In_224,N_106);
nand U231 (N_231,In_334,N_167);
nand U232 (N_232,In_264,N_74);
nand U233 (N_233,N_58,In_382);
xnor U234 (N_234,In_326,In_431);
and U235 (N_235,N_103,N_47);
nor U236 (N_236,N_120,N_166);
nor U237 (N_237,N_71,N_50);
nand U238 (N_238,N_161,N_124);
nand U239 (N_239,N_146,N_126);
and U240 (N_240,N_197,In_182);
xnor U241 (N_241,N_99,In_404);
nand U242 (N_242,In_411,N_43);
or U243 (N_243,In_430,N_162);
and U244 (N_244,N_119,N_158);
or U245 (N_245,In_268,N_125);
xnor U246 (N_246,N_75,In_375);
nor U247 (N_247,N_175,N_13);
nor U248 (N_248,In_400,N_92);
xor U249 (N_249,In_361,N_138);
xnor U250 (N_250,In_433,N_60);
xnor U251 (N_251,In_287,N_94);
nand U252 (N_252,N_107,In_458);
and U253 (N_253,N_191,N_130);
nor U254 (N_254,N_8,In_498);
nor U255 (N_255,N_35,In_380);
or U256 (N_256,In_357,N_118);
and U257 (N_257,N_51,N_108);
nor U258 (N_258,N_87,N_31);
nand U259 (N_259,N_1,N_54);
nor U260 (N_260,In_73,In_340);
xor U261 (N_261,In_57,N_76);
or U262 (N_262,N_149,N_140);
and U263 (N_263,In_346,N_179);
xor U264 (N_264,In_231,N_100);
nor U265 (N_265,N_172,In_336);
or U266 (N_266,N_5,N_89);
nand U267 (N_267,N_98,In_36);
or U268 (N_268,In_427,N_83);
or U269 (N_269,N_56,N_12);
and U270 (N_270,In_152,In_85);
or U271 (N_271,N_7,In_114);
nor U272 (N_272,In_486,N_23);
nor U273 (N_273,N_91,N_142);
nor U274 (N_274,In_27,N_163);
and U275 (N_275,N_93,N_69);
and U276 (N_276,In_69,In_218);
or U277 (N_277,N_128,N_84);
nand U278 (N_278,N_144,In_49);
xor U279 (N_279,N_127,N_32);
or U280 (N_280,N_36,N_177);
xnor U281 (N_281,N_196,N_97);
and U282 (N_282,N_53,N_198);
or U283 (N_283,N_152,In_183);
and U284 (N_284,N_110,N_45);
nor U285 (N_285,N_154,N_11);
or U286 (N_286,In_365,N_61);
nand U287 (N_287,N_55,N_187);
and U288 (N_288,In_193,In_302);
nand U289 (N_289,N_16,In_7);
xor U290 (N_290,N_148,In_258);
nand U291 (N_291,N_73,In_250);
or U292 (N_292,N_26,N_72);
nor U293 (N_293,N_182,In_298);
or U294 (N_294,In_34,N_165);
xnor U295 (N_295,N_190,N_192);
nand U296 (N_296,N_193,N_64);
xnor U297 (N_297,N_2,N_63);
xnor U298 (N_298,In_92,In_355);
xor U299 (N_299,N_176,N_159);
or U300 (N_300,In_397,N_147);
or U301 (N_301,N_85,N_136);
and U302 (N_302,In_453,N_29);
nand U303 (N_303,N_28,N_156);
and U304 (N_304,In_344,N_139);
nand U305 (N_305,N_112,N_188);
nor U306 (N_306,N_24,N_185);
nor U307 (N_307,In_46,In_394);
xnor U308 (N_308,N_114,In_2);
xor U309 (N_309,N_174,In_246);
or U310 (N_310,N_168,N_65);
nand U311 (N_311,In_324,In_315);
xor U312 (N_312,N_0,N_111);
nand U313 (N_313,N_195,In_205);
nand U314 (N_314,N_184,N_10);
or U315 (N_315,N_52,In_172);
nor U316 (N_316,N_122,In_276);
and U317 (N_317,In_270,N_77);
or U318 (N_318,N_34,N_42);
or U319 (N_319,In_329,In_106);
or U320 (N_320,N_90,In_390);
and U321 (N_321,N_96,N_151);
nor U322 (N_322,In_192,N_41);
nand U323 (N_323,In_472,N_178);
xnor U324 (N_324,N_134,In_408);
nor U325 (N_325,N_39,In_297);
xnor U326 (N_326,In_206,In_233);
nor U327 (N_327,In_416,N_20);
xnor U328 (N_328,N_82,N_109);
or U329 (N_329,N_113,In_456);
xor U330 (N_330,N_180,N_44);
and U331 (N_331,In_68,In_385);
or U332 (N_332,N_30,N_104);
or U333 (N_333,N_62,In_115);
nor U334 (N_334,N_81,N_86);
xnor U335 (N_335,N_66,N_141);
nor U336 (N_336,N_150,N_117);
or U337 (N_337,N_135,N_78);
and U338 (N_338,N_189,N_143);
and U339 (N_339,In_332,In_305);
xor U340 (N_340,N_33,N_123);
nor U341 (N_341,N_102,In_81);
or U342 (N_342,N_46,N_18);
xnor U343 (N_343,N_169,N_21);
xor U344 (N_344,In_317,N_15);
or U345 (N_345,N_38,N_105);
nor U346 (N_346,In_414,N_88);
xnor U347 (N_347,In_67,N_22);
nor U348 (N_348,N_57,In_352);
and U349 (N_349,In_230,In_75);
and U350 (N_350,In_67,N_110);
nand U351 (N_351,N_75,N_192);
nor U352 (N_352,N_166,N_57);
nand U353 (N_353,In_340,In_264);
and U354 (N_354,N_6,N_150);
xor U355 (N_355,N_107,In_397);
and U356 (N_356,N_63,N_71);
xor U357 (N_357,N_7,N_74);
and U358 (N_358,N_54,N_133);
xor U359 (N_359,N_80,In_473);
or U360 (N_360,N_20,N_193);
nand U361 (N_361,N_17,In_456);
nand U362 (N_362,N_102,In_390);
nor U363 (N_363,In_115,N_119);
nand U364 (N_364,N_166,N_82);
xor U365 (N_365,N_44,In_380);
and U366 (N_366,N_65,N_102);
nor U367 (N_367,In_81,N_97);
xnor U368 (N_368,N_69,N_14);
nand U369 (N_369,In_336,N_149);
xnor U370 (N_370,N_132,N_155);
or U371 (N_371,N_181,N_170);
or U372 (N_372,N_136,In_498);
and U373 (N_373,N_187,In_7);
nand U374 (N_374,In_336,N_171);
xnor U375 (N_375,N_43,N_47);
nor U376 (N_376,N_10,N_73);
nor U377 (N_377,In_472,N_141);
nand U378 (N_378,In_208,N_151);
xnor U379 (N_379,N_75,N_41);
or U380 (N_380,N_27,N_6);
or U381 (N_381,In_411,In_305);
nor U382 (N_382,N_87,N_129);
and U383 (N_383,In_404,N_100);
or U384 (N_384,N_155,N_109);
nor U385 (N_385,N_173,N_160);
and U386 (N_386,N_7,In_365);
and U387 (N_387,N_176,N_187);
or U388 (N_388,N_188,N_123);
and U389 (N_389,In_340,N_36);
nor U390 (N_390,N_146,N_85);
nor U391 (N_391,In_182,In_334);
and U392 (N_392,In_498,N_14);
xnor U393 (N_393,N_126,N_129);
nor U394 (N_394,N_20,In_92);
and U395 (N_395,In_416,N_182);
xor U396 (N_396,In_334,N_98);
and U397 (N_397,N_50,N_3);
or U398 (N_398,N_119,N_102);
and U399 (N_399,N_22,In_7);
or U400 (N_400,N_294,N_347);
nor U401 (N_401,N_328,N_284);
nand U402 (N_402,N_280,N_260);
and U403 (N_403,N_276,N_387);
xnor U404 (N_404,N_384,N_314);
xnor U405 (N_405,N_363,N_222);
and U406 (N_406,N_270,N_392);
nand U407 (N_407,N_228,N_268);
xor U408 (N_408,N_323,N_358);
nor U409 (N_409,N_214,N_297);
nand U410 (N_410,N_245,N_313);
nand U411 (N_411,N_310,N_200);
nand U412 (N_412,N_380,N_244);
or U413 (N_413,N_207,N_292);
nand U414 (N_414,N_286,N_259);
or U415 (N_415,N_386,N_394);
or U416 (N_416,N_360,N_203);
nand U417 (N_417,N_204,N_283);
and U418 (N_418,N_243,N_248);
nor U419 (N_419,N_212,N_338);
and U420 (N_420,N_215,N_218);
nand U421 (N_421,N_242,N_262);
nor U422 (N_422,N_235,N_217);
or U423 (N_423,N_226,N_255);
nor U424 (N_424,N_361,N_232);
nor U425 (N_425,N_306,N_397);
and U426 (N_426,N_389,N_377);
nand U427 (N_427,N_261,N_209);
nor U428 (N_428,N_330,N_354);
nand U429 (N_429,N_274,N_319);
or U430 (N_430,N_370,N_303);
nand U431 (N_431,N_351,N_369);
nand U432 (N_432,N_388,N_353);
xnor U433 (N_433,N_381,N_229);
nor U434 (N_434,N_374,N_329);
and U435 (N_435,N_246,N_339);
xnor U436 (N_436,N_201,N_266);
nor U437 (N_437,N_219,N_334);
and U438 (N_438,N_299,N_220);
and U439 (N_439,N_290,N_342);
xnor U440 (N_440,N_321,N_367);
nand U441 (N_441,N_337,N_375);
xnor U442 (N_442,N_288,N_293);
nand U443 (N_443,N_251,N_216);
and U444 (N_444,N_366,N_371);
xnor U445 (N_445,N_273,N_240);
nand U446 (N_446,N_281,N_233);
nand U447 (N_447,N_258,N_317);
and U448 (N_448,N_382,N_352);
or U449 (N_449,N_391,N_379);
or U450 (N_450,N_236,N_291);
and U451 (N_451,N_208,N_322);
xor U452 (N_452,N_239,N_385);
xor U453 (N_453,N_275,N_300);
xor U454 (N_454,N_238,N_265);
nor U455 (N_455,N_237,N_341);
nor U456 (N_456,N_287,N_223);
nor U457 (N_457,N_399,N_249);
nand U458 (N_458,N_250,N_348);
nor U459 (N_459,N_271,N_213);
xnor U460 (N_460,N_359,N_278);
nand U461 (N_461,N_315,N_234);
or U462 (N_462,N_316,N_365);
nor U463 (N_463,N_221,N_373);
nor U464 (N_464,N_254,N_307);
xnor U465 (N_465,N_231,N_202);
and U466 (N_466,N_205,N_269);
nand U467 (N_467,N_206,N_241);
or U468 (N_468,N_247,N_253);
nor U469 (N_469,N_390,N_343);
nand U470 (N_470,N_256,N_320);
or U471 (N_471,N_376,N_279);
and U472 (N_472,N_311,N_272);
and U473 (N_473,N_318,N_331);
nor U474 (N_474,N_383,N_356);
nor U475 (N_475,N_210,N_252);
xor U476 (N_476,N_302,N_308);
xor U477 (N_477,N_305,N_395);
and U478 (N_478,N_346,N_340);
or U479 (N_479,N_296,N_344);
xor U480 (N_480,N_224,N_349);
and U481 (N_481,N_324,N_398);
and U482 (N_482,N_230,N_267);
nor U483 (N_483,N_285,N_362);
or U484 (N_484,N_312,N_327);
nor U485 (N_485,N_378,N_282);
and U486 (N_486,N_350,N_396);
xnor U487 (N_487,N_357,N_335);
or U488 (N_488,N_372,N_301);
xnor U489 (N_489,N_309,N_325);
nor U490 (N_490,N_332,N_227);
or U491 (N_491,N_277,N_257);
nand U492 (N_492,N_289,N_298);
and U493 (N_493,N_263,N_264);
xor U494 (N_494,N_295,N_393);
xnor U495 (N_495,N_225,N_304);
nand U496 (N_496,N_345,N_333);
nand U497 (N_497,N_355,N_211);
or U498 (N_498,N_336,N_326);
and U499 (N_499,N_364,N_368);
or U500 (N_500,N_297,N_384);
and U501 (N_501,N_330,N_306);
or U502 (N_502,N_201,N_318);
or U503 (N_503,N_324,N_314);
nand U504 (N_504,N_284,N_395);
xnor U505 (N_505,N_266,N_214);
and U506 (N_506,N_315,N_369);
or U507 (N_507,N_278,N_301);
nor U508 (N_508,N_396,N_306);
and U509 (N_509,N_244,N_209);
or U510 (N_510,N_286,N_213);
nor U511 (N_511,N_324,N_304);
nor U512 (N_512,N_342,N_382);
nor U513 (N_513,N_262,N_307);
xnor U514 (N_514,N_270,N_303);
or U515 (N_515,N_371,N_311);
nor U516 (N_516,N_387,N_282);
and U517 (N_517,N_327,N_248);
xor U518 (N_518,N_287,N_252);
nand U519 (N_519,N_350,N_281);
and U520 (N_520,N_272,N_258);
nor U521 (N_521,N_260,N_215);
nor U522 (N_522,N_243,N_272);
nand U523 (N_523,N_211,N_231);
nand U524 (N_524,N_281,N_348);
nor U525 (N_525,N_373,N_266);
nor U526 (N_526,N_279,N_241);
xor U527 (N_527,N_360,N_353);
xor U528 (N_528,N_297,N_251);
nor U529 (N_529,N_293,N_205);
and U530 (N_530,N_360,N_381);
and U531 (N_531,N_249,N_248);
nand U532 (N_532,N_323,N_287);
nor U533 (N_533,N_267,N_282);
or U534 (N_534,N_302,N_394);
or U535 (N_535,N_268,N_298);
nand U536 (N_536,N_291,N_298);
nand U537 (N_537,N_253,N_351);
or U538 (N_538,N_204,N_216);
and U539 (N_539,N_268,N_223);
nand U540 (N_540,N_369,N_383);
and U541 (N_541,N_223,N_397);
or U542 (N_542,N_344,N_378);
or U543 (N_543,N_242,N_329);
xor U544 (N_544,N_328,N_229);
or U545 (N_545,N_203,N_288);
nand U546 (N_546,N_244,N_280);
xor U547 (N_547,N_283,N_399);
and U548 (N_548,N_322,N_347);
nand U549 (N_549,N_294,N_254);
xnor U550 (N_550,N_385,N_312);
nand U551 (N_551,N_228,N_216);
nand U552 (N_552,N_249,N_262);
nand U553 (N_553,N_354,N_272);
or U554 (N_554,N_385,N_255);
nand U555 (N_555,N_227,N_362);
nor U556 (N_556,N_237,N_381);
nand U557 (N_557,N_388,N_374);
xor U558 (N_558,N_255,N_374);
nand U559 (N_559,N_297,N_370);
or U560 (N_560,N_335,N_293);
nand U561 (N_561,N_359,N_232);
and U562 (N_562,N_296,N_368);
or U563 (N_563,N_349,N_201);
nor U564 (N_564,N_340,N_223);
nor U565 (N_565,N_231,N_225);
nand U566 (N_566,N_383,N_392);
nor U567 (N_567,N_296,N_350);
or U568 (N_568,N_251,N_339);
and U569 (N_569,N_231,N_220);
nand U570 (N_570,N_381,N_201);
nor U571 (N_571,N_269,N_353);
and U572 (N_572,N_258,N_281);
nor U573 (N_573,N_285,N_272);
and U574 (N_574,N_211,N_313);
nor U575 (N_575,N_246,N_265);
or U576 (N_576,N_302,N_351);
nor U577 (N_577,N_203,N_205);
and U578 (N_578,N_207,N_284);
or U579 (N_579,N_355,N_362);
and U580 (N_580,N_278,N_320);
and U581 (N_581,N_348,N_263);
or U582 (N_582,N_311,N_352);
nand U583 (N_583,N_376,N_303);
nor U584 (N_584,N_339,N_307);
or U585 (N_585,N_273,N_229);
xor U586 (N_586,N_384,N_321);
and U587 (N_587,N_223,N_236);
and U588 (N_588,N_267,N_314);
xor U589 (N_589,N_299,N_356);
or U590 (N_590,N_311,N_277);
nor U591 (N_591,N_261,N_219);
and U592 (N_592,N_236,N_257);
or U593 (N_593,N_271,N_214);
nand U594 (N_594,N_239,N_335);
nor U595 (N_595,N_239,N_398);
and U596 (N_596,N_320,N_323);
nor U597 (N_597,N_256,N_232);
or U598 (N_598,N_202,N_391);
nand U599 (N_599,N_240,N_226);
nor U600 (N_600,N_513,N_530);
or U601 (N_601,N_535,N_523);
xor U602 (N_602,N_419,N_548);
nand U603 (N_603,N_520,N_593);
nand U604 (N_604,N_441,N_572);
and U605 (N_605,N_594,N_425);
nor U606 (N_606,N_514,N_506);
or U607 (N_607,N_439,N_416);
xor U608 (N_608,N_407,N_564);
nor U609 (N_609,N_457,N_463);
and U610 (N_610,N_536,N_400);
and U611 (N_611,N_488,N_438);
xnor U612 (N_612,N_481,N_466);
and U613 (N_613,N_583,N_541);
nand U614 (N_614,N_467,N_571);
nand U615 (N_615,N_569,N_592);
nor U616 (N_616,N_544,N_537);
and U617 (N_617,N_597,N_462);
nor U618 (N_618,N_549,N_472);
nand U619 (N_619,N_505,N_598);
or U620 (N_620,N_582,N_404);
nor U621 (N_621,N_521,N_448);
xnor U622 (N_622,N_446,N_574);
or U623 (N_623,N_485,N_490);
and U624 (N_624,N_496,N_477);
and U625 (N_625,N_554,N_480);
nor U626 (N_626,N_487,N_581);
nand U627 (N_627,N_482,N_534);
or U628 (N_628,N_473,N_451);
and U629 (N_629,N_540,N_479);
nor U630 (N_630,N_423,N_561);
nor U631 (N_631,N_464,N_405);
or U632 (N_632,N_413,N_458);
and U633 (N_633,N_420,N_551);
and U634 (N_634,N_509,N_435);
or U635 (N_635,N_546,N_459);
and U636 (N_636,N_556,N_575);
xnor U637 (N_637,N_542,N_504);
nand U638 (N_638,N_460,N_492);
xnor U639 (N_639,N_494,N_427);
nor U640 (N_640,N_552,N_432);
nand U641 (N_641,N_595,N_570);
nor U642 (N_642,N_422,N_566);
and U643 (N_643,N_450,N_591);
and U644 (N_644,N_527,N_568);
or U645 (N_645,N_415,N_410);
and U646 (N_646,N_547,N_414);
nor U647 (N_647,N_498,N_495);
nand U648 (N_648,N_409,N_517);
nand U649 (N_649,N_456,N_412);
nand U650 (N_650,N_526,N_493);
xnor U651 (N_651,N_528,N_532);
and U652 (N_652,N_440,N_411);
nor U653 (N_653,N_401,N_565);
nor U654 (N_654,N_510,N_533);
xnor U655 (N_655,N_524,N_417);
nor U656 (N_656,N_471,N_406);
nor U657 (N_657,N_461,N_442);
nand U658 (N_658,N_543,N_508);
xor U659 (N_659,N_476,N_573);
xnor U660 (N_660,N_522,N_525);
and U661 (N_661,N_499,N_449);
or U662 (N_662,N_402,N_433);
and U663 (N_663,N_529,N_584);
and U664 (N_664,N_589,N_484);
xor U665 (N_665,N_444,N_428);
and U666 (N_666,N_576,N_587);
or U667 (N_667,N_585,N_501);
and U668 (N_668,N_599,N_486);
nand U669 (N_669,N_550,N_474);
nand U670 (N_670,N_553,N_512);
nand U671 (N_671,N_567,N_580);
nand U672 (N_672,N_586,N_500);
nor U673 (N_673,N_418,N_511);
nor U674 (N_674,N_579,N_560);
xnor U675 (N_675,N_515,N_539);
or U676 (N_676,N_483,N_545);
nand U677 (N_677,N_443,N_408);
nand U678 (N_678,N_577,N_531);
xor U679 (N_679,N_519,N_596);
xor U680 (N_680,N_558,N_489);
nand U681 (N_681,N_475,N_431);
xor U682 (N_682,N_454,N_465);
xnor U683 (N_683,N_452,N_445);
and U684 (N_684,N_455,N_562);
nand U685 (N_685,N_424,N_437);
or U686 (N_686,N_421,N_434);
nor U687 (N_687,N_426,N_502);
nand U688 (N_688,N_503,N_588);
nor U689 (N_689,N_563,N_470);
xnor U690 (N_690,N_469,N_468);
and U691 (N_691,N_518,N_429);
xnor U692 (N_692,N_590,N_478);
or U693 (N_693,N_436,N_403);
and U694 (N_694,N_491,N_557);
and U695 (N_695,N_447,N_453);
nand U696 (N_696,N_559,N_430);
xor U697 (N_697,N_516,N_538);
nand U698 (N_698,N_555,N_497);
or U699 (N_699,N_578,N_507);
xnor U700 (N_700,N_588,N_546);
nand U701 (N_701,N_401,N_479);
or U702 (N_702,N_442,N_434);
and U703 (N_703,N_498,N_419);
xnor U704 (N_704,N_480,N_491);
xnor U705 (N_705,N_511,N_445);
or U706 (N_706,N_420,N_565);
nand U707 (N_707,N_436,N_473);
or U708 (N_708,N_486,N_494);
xor U709 (N_709,N_424,N_484);
and U710 (N_710,N_420,N_583);
and U711 (N_711,N_486,N_566);
xnor U712 (N_712,N_478,N_510);
nand U713 (N_713,N_523,N_528);
xor U714 (N_714,N_484,N_400);
nand U715 (N_715,N_574,N_561);
or U716 (N_716,N_550,N_427);
nand U717 (N_717,N_428,N_474);
nand U718 (N_718,N_455,N_464);
or U719 (N_719,N_406,N_561);
xor U720 (N_720,N_508,N_527);
or U721 (N_721,N_599,N_419);
nor U722 (N_722,N_456,N_417);
xnor U723 (N_723,N_587,N_512);
and U724 (N_724,N_566,N_585);
nand U725 (N_725,N_515,N_434);
or U726 (N_726,N_411,N_530);
or U727 (N_727,N_540,N_434);
and U728 (N_728,N_590,N_577);
nand U729 (N_729,N_575,N_521);
and U730 (N_730,N_566,N_580);
and U731 (N_731,N_440,N_409);
xor U732 (N_732,N_408,N_538);
nor U733 (N_733,N_440,N_421);
nand U734 (N_734,N_417,N_452);
nor U735 (N_735,N_536,N_540);
or U736 (N_736,N_598,N_543);
and U737 (N_737,N_419,N_471);
xnor U738 (N_738,N_538,N_434);
xnor U739 (N_739,N_439,N_517);
and U740 (N_740,N_485,N_421);
and U741 (N_741,N_570,N_436);
nor U742 (N_742,N_424,N_544);
or U743 (N_743,N_493,N_511);
nand U744 (N_744,N_594,N_524);
or U745 (N_745,N_561,N_573);
and U746 (N_746,N_536,N_439);
xnor U747 (N_747,N_480,N_521);
and U748 (N_748,N_555,N_484);
nor U749 (N_749,N_420,N_545);
nor U750 (N_750,N_539,N_424);
and U751 (N_751,N_587,N_500);
and U752 (N_752,N_407,N_553);
nand U753 (N_753,N_402,N_521);
or U754 (N_754,N_466,N_549);
nor U755 (N_755,N_511,N_587);
and U756 (N_756,N_550,N_411);
and U757 (N_757,N_504,N_411);
xnor U758 (N_758,N_532,N_498);
xor U759 (N_759,N_421,N_534);
and U760 (N_760,N_434,N_568);
nor U761 (N_761,N_426,N_452);
and U762 (N_762,N_584,N_424);
nor U763 (N_763,N_558,N_414);
xor U764 (N_764,N_437,N_479);
nand U765 (N_765,N_500,N_410);
xnor U766 (N_766,N_433,N_430);
nor U767 (N_767,N_554,N_521);
nor U768 (N_768,N_452,N_478);
or U769 (N_769,N_577,N_417);
nor U770 (N_770,N_470,N_402);
and U771 (N_771,N_589,N_565);
nor U772 (N_772,N_563,N_457);
and U773 (N_773,N_491,N_443);
or U774 (N_774,N_576,N_536);
xor U775 (N_775,N_523,N_500);
and U776 (N_776,N_476,N_484);
nand U777 (N_777,N_428,N_552);
and U778 (N_778,N_439,N_434);
or U779 (N_779,N_495,N_597);
nand U780 (N_780,N_512,N_564);
or U781 (N_781,N_469,N_463);
nand U782 (N_782,N_466,N_483);
nor U783 (N_783,N_485,N_515);
nor U784 (N_784,N_442,N_502);
nor U785 (N_785,N_463,N_467);
xnor U786 (N_786,N_450,N_463);
and U787 (N_787,N_430,N_585);
or U788 (N_788,N_528,N_578);
or U789 (N_789,N_562,N_497);
or U790 (N_790,N_599,N_445);
or U791 (N_791,N_542,N_587);
xnor U792 (N_792,N_411,N_446);
or U793 (N_793,N_419,N_515);
nand U794 (N_794,N_439,N_534);
nor U795 (N_795,N_521,N_585);
xnor U796 (N_796,N_481,N_565);
or U797 (N_797,N_450,N_427);
nor U798 (N_798,N_439,N_503);
xnor U799 (N_799,N_536,N_501);
xor U800 (N_800,N_690,N_646);
xnor U801 (N_801,N_635,N_624);
or U802 (N_802,N_606,N_629);
and U803 (N_803,N_664,N_745);
or U804 (N_804,N_602,N_647);
or U805 (N_805,N_603,N_619);
or U806 (N_806,N_798,N_700);
nand U807 (N_807,N_654,N_702);
xnor U808 (N_808,N_668,N_652);
nor U809 (N_809,N_665,N_648);
or U810 (N_810,N_712,N_696);
and U811 (N_811,N_787,N_715);
nor U812 (N_812,N_760,N_734);
xor U813 (N_813,N_786,N_617);
xor U814 (N_814,N_722,N_643);
or U815 (N_815,N_601,N_615);
nor U816 (N_816,N_768,N_781);
or U817 (N_817,N_739,N_618);
nor U818 (N_818,N_782,N_737);
or U819 (N_819,N_772,N_795);
or U820 (N_820,N_637,N_735);
and U821 (N_821,N_677,N_680);
or U822 (N_822,N_756,N_688);
nor U823 (N_823,N_723,N_607);
and U824 (N_824,N_730,N_790);
nand U825 (N_825,N_655,N_764);
or U826 (N_826,N_758,N_775);
nand U827 (N_827,N_742,N_632);
xor U828 (N_828,N_639,N_683);
xor U829 (N_829,N_682,N_627);
xor U830 (N_830,N_649,N_681);
and U831 (N_831,N_699,N_642);
or U832 (N_832,N_721,N_779);
nor U833 (N_833,N_796,N_612);
nand U834 (N_834,N_622,N_773);
xor U835 (N_835,N_733,N_666);
nor U836 (N_836,N_670,N_713);
nor U837 (N_837,N_705,N_633);
nand U838 (N_838,N_678,N_759);
xnor U839 (N_839,N_708,N_727);
xnor U840 (N_840,N_650,N_761);
nand U841 (N_841,N_789,N_725);
xor U842 (N_842,N_740,N_620);
or U843 (N_843,N_684,N_778);
nand U844 (N_844,N_663,N_767);
nor U845 (N_845,N_638,N_608);
nor U846 (N_846,N_752,N_610);
nand U847 (N_847,N_728,N_776);
xor U848 (N_848,N_797,N_766);
and U849 (N_849,N_704,N_750);
nor U850 (N_850,N_634,N_792);
nor U851 (N_851,N_686,N_770);
or U852 (N_852,N_703,N_679);
xor U853 (N_853,N_777,N_724);
or U854 (N_854,N_657,N_671);
or U855 (N_855,N_757,N_799);
xor U856 (N_856,N_625,N_687);
nand U857 (N_857,N_611,N_673);
and U858 (N_858,N_613,N_784);
nor U859 (N_859,N_755,N_780);
xnor U860 (N_860,N_609,N_763);
nand U861 (N_861,N_707,N_689);
xnor U862 (N_862,N_626,N_714);
nor U863 (N_863,N_640,N_743);
and U864 (N_864,N_741,N_604);
xnor U865 (N_865,N_651,N_706);
nor U866 (N_866,N_660,N_645);
and U867 (N_867,N_658,N_711);
nor U868 (N_868,N_662,N_746);
xor U869 (N_869,N_605,N_697);
or U870 (N_870,N_726,N_674);
and U871 (N_871,N_791,N_623);
or U872 (N_872,N_691,N_628);
xnor U873 (N_873,N_718,N_736);
and U874 (N_874,N_692,N_636);
nor U875 (N_875,N_748,N_675);
nor U876 (N_876,N_631,N_695);
nor U877 (N_877,N_676,N_783);
nand U878 (N_878,N_765,N_716);
or U879 (N_879,N_698,N_753);
nor U880 (N_880,N_738,N_710);
xor U881 (N_881,N_794,N_720);
nor U882 (N_882,N_661,N_769);
and U883 (N_883,N_771,N_614);
or U884 (N_884,N_644,N_751);
nand U885 (N_885,N_709,N_717);
xor U886 (N_886,N_672,N_694);
xnor U887 (N_887,N_774,N_749);
xor U888 (N_888,N_754,N_667);
or U889 (N_889,N_600,N_732);
nand U890 (N_890,N_630,N_701);
nor U891 (N_891,N_788,N_762);
or U892 (N_892,N_793,N_621);
or U893 (N_893,N_731,N_693);
or U894 (N_894,N_653,N_641);
and U895 (N_895,N_719,N_747);
nand U896 (N_896,N_616,N_669);
or U897 (N_897,N_656,N_659);
or U898 (N_898,N_685,N_744);
xnor U899 (N_899,N_785,N_729);
nand U900 (N_900,N_650,N_769);
nand U901 (N_901,N_761,N_704);
or U902 (N_902,N_756,N_799);
nand U903 (N_903,N_601,N_700);
nor U904 (N_904,N_636,N_783);
nand U905 (N_905,N_781,N_751);
nor U906 (N_906,N_743,N_705);
nor U907 (N_907,N_683,N_771);
or U908 (N_908,N_669,N_765);
nand U909 (N_909,N_672,N_664);
xnor U910 (N_910,N_622,N_747);
or U911 (N_911,N_650,N_727);
and U912 (N_912,N_722,N_611);
xnor U913 (N_913,N_752,N_692);
or U914 (N_914,N_780,N_667);
and U915 (N_915,N_729,N_685);
nor U916 (N_916,N_705,N_799);
xor U917 (N_917,N_744,N_727);
and U918 (N_918,N_652,N_676);
xor U919 (N_919,N_606,N_729);
or U920 (N_920,N_642,N_778);
nand U921 (N_921,N_645,N_751);
or U922 (N_922,N_747,N_742);
xor U923 (N_923,N_674,N_635);
and U924 (N_924,N_793,N_619);
xnor U925 (N_925,N_713,N_796);
or U926 (N_926,N_686,N_764);
nor U927 (N_927,N_757,N_620);
xnor U928 (N_928,N_716,N_604);
nor U929 (N_929,N_660,N_753);
xnor U930 (N_930,N_745,N_705);
nor U931 (N_931,N_760,N_608);
and U932 (N_932,N_702,N_757);
and U933 (N_933,N_726,N_704);
and U934 (N_934,N_775,N_754);
and U935 (N_935,N_697,N_736);
and U936 (N_936,N_631,N_671);
nand U937 (N_937,N_770,N_793);
nor U938 (N_938,N_670,N_630);
xor U939 (N_939,N_706,N_664);
nor U940 (N_940,N_778,N_726);
and U941 (N_941,N_698,N_696);
or U942 (N_942,N_746,N_659);
or U943 (N_943,N_630,N_675);
xnor U944 (N_944,N_687,N_714);
xnor U945 (N_945,N_600,N_784);
nand U946 (N_946,N_665,N_756);
and U947 (N_947,N_634,N_760);
or U948 (N_948,N_786,N_601);
xnor U949 (N_949,N_753,N_679);
xor U950 (N_950,N_640,N_727);
xor U951 (N_951,N_667,N_695);
nor U952 (N_952,N_757,N_679);
xor U953 (N_953,N_601,N_748);
nand U954 (N_954,N_757,N_792);
or U955 (N_955,N_669,N_603);
nor U956 (N_956,N_790,N_717);
nand U957 (N_957,N_600,N_668);
nor U958 (N_958,N_777,N_706);
nand U959 (N_959,N_665,N_629);
nor U960 (N_960,N_730,N_648);
or U961 (N_961,N_628,N_732);
nand U962 (N_962,N_755,N_622);
and U963 (N_963,N_606,N_757);
and U964 (N_964,N_795,N_792);
nor U965 (N_965,N_671,N_695);
nor U966 (N_966,N_628,N_769);
nand U967 (N_967,N_709,N_780);
nor U968 (N_968,N_714,N_769);
nor U969 (N_969,N_754,N_745);
nor U970 (N_970,N_682,N_772);
nand U971 (N_971,N_799,N_781);
nand U972 (N_972,N_701,N_672);
or U973 (N_973,N_732,N_670);
nand U974 (N_974,N_608,N_652);
xor U975 (N_975,N_707,N_718);
and U976 (N_976,N_628,N_791);
nand U977 (N_977,N_772,N_715);
nand U978 (N_978,N_711,N_653);
nor U979 (N_979,N_746,N_641);
nand U980 (N_980,N_662,N_689);
and U981 (N_981,N_692,N_755);
nand U982 (N_982,N_633,N_712);
xnor U983 (N_983,N_624,N_773);
and U984 (N_984,N_741,N_619);
or U985 (N_985,N_775,N_798);
and U986 (N_986,N_724,N_632);
and U987 (N_987,N_628,N_762);
nand U988 (N_988,N_673,N_647);
and U989 (N_989,N_725,N_637);
and U990 (N_990,N_681,N_764);
xnor U991 (N_991,N_636,N_789);
nor U992 (N_992,N_788,N_668);
nor U993 (N_993,N_729,N_768);
xnor U994 (N_994,N_601,N_768);
nand U995 (N_995,N_717,N_799);
xnor U996 (N_996,N_787,N_798);
nand U997 (N_997,N_606,N_723);
xnor U998 (N_998,N_751,N_766);
xor U999 (N_999,N_749,N_772);
nand U1000 (N_1000,N_810,N_808);
xnor U1001 (N_1001,N_910,N_859);
nor U1002 (N_1002,N_868,N_879);
or U1003 (N_1003,N_811,N_894);
xor U1004 (N_1004,N_920,N_992);
and U1005 (N_1005,N_994,N_937);
nand U1006 (N_1006,N_861,N_829);
nor U1007 (N_1007,N_847,N_979);
nand U1008 (N_1008,N_941,N_821);
or U1009 (N_1009,N_932,N_851);
and U1010 (N_1010,N_940,N_918);
or U1011 (N_1011,N_883,N_885);
nand U1012 (N_1012,N_878,N_950);
or U1013 (N_1013,N_828,N_956);
and U1014 (N_1014,N_902,N_976);
nor U1015 (N_1015,N_857,N_969);
xnor U1016 (N_1016,N_930,N_949);
nand U1017 (N_1017,N_884,N_826);
or U1018 (N_1018,N_998,N_844);
nand U1019 (N_1019,N_849,N_960);
nor U1020 (N_1020,N_995,N_934);
nand U1021 (N_1021,N_993,N_974);
nor U1022 (N_1022,N_882,N_899);
and U1023 (N_1023,N_822,N_863);
and U1024 (N_1024,N_886,N_888);
nor U1025 (N_1025,N_957,N_825);
nand U1026 (N_1026,N_819,N_905);
or U1027 (N_1027,N_947,N_893);
nor U1028 (N_1028,N_964,N_996);
and U1029 (N_1029,N_848,N_989);
nor U1030 (N_1030,N_911,N_831);
or U1031 (N_1031,N_967,N_985);
and U1032 (N_1032,N_954,N_933);
xnor U1033 (N_1033,N_870,N_841);
nand U1034 (N_1034,N_850,N_951);
xor U1035 (N_1035,N_890,N_919);
and U1036 (N_1036,N_914,N_921);
or U1037 (N_1037,N_897,N_896);
xor U1038 (N_1038,N_970,N_815);
or U1039 (N_1039,N_975,N_952);
and U1040 (N_1040,N_820,N_982);
or U1041 (N_1041,N_824,N_809);
or U1042 (N_1042,N_986,N_832);
nor U1043 (N_1043,N_855,N_968);
xnor U1044 (N_1044,N_805,N_927);
nor U1045 (N_1045,N_802,N_917);
nand U1046 (N_1046,N_959,N_997);
and U1047 (N_1047,N_906,N_991);
xor U1048 (N_1048,N_833,N_843);
nor U1049 (N_1049,N_830,N_891);
or U1050 (N_1050,N_887,N_889);
nor U1051 (N_1051,N_984,N_901);
and U1052 (N_1052,N_963,N_912);
nand U1053 (N_1053,N_904,N_942);
nand U1054 (N_1054,N_945,N_856);
nor U1055 (N_1055,N_909,N_871);
nand U1056 (N_1056,N_922,N_931);
nor U1057 (N_1057,N_987,N_898);
nand U1058 (N_1058,N_842,N_845);
or U1059 (N_1059,N_846,N_938);
or U1060 (N_1060,N_983,N_840);
nor U1061 (N_1061,N_836,N_962);
and U1062 (N_1062,N_999,N_862);
or U1063 (N_1063,N_981,N_980);
nor U1064 (N_1064,N_880,N_874);
or U1065 (N_1065,N_972,N_966);
nor U1066 (N_1066,N_953,N_804);
or U1067 (N_1067,N_939,N_903);
nor U1068 (N_1068,N_924,N_816);
nor U1069 (N_1069,N_867,N_835);
and U1070 (N_1070,N_900,N_936);
nor U1071 (N_1071,N_869,N_818);
and U1072 (N_1072,N_971,N_907);
or U1073 (N_1073,N_946,N_803);
xnor U1074 (N_1074,N_823,N_814);
and U1075 (N_1075,N_943,N_923);
nor U1076 (N_1076,N_955,N_853);
xnor U1077 (N_1077,N_961,N_834);
nand U1078 (N_1078,N_812,N_876);
nor U1079 (N_1079,N_860,N_852);
nand U1080 (N_1080,N_875,N_895);
nand U1081 (N_1081,N_838,N_929);
xnor U1082 (N_1082,N_977,N_928);
nand U1083 (N_1083,N_866,N_978);
nor U1084 (N_1084,N_872,N_935);
nand U1085 (N_1085,N_913,N_965);
nand U1086 (N_1086,N_948,N_839);
or U1087 (N_1087,N_817,N_892);
nand U1088 (N_1088,N_864,N_837);
and U1089 (N_1089,N_877,N_827);
xor U1090 (N_1090,N_973,N_807);
nand U1091 (N_1091,N_801,N_873);
or U1092 (N_1092,N_865,N_990);
nor U1093 (N_1093,N_988,N_800);
xnor U1094 (N_1094,N_958,N_858);
xor U1095 (N_1095,N_915,N_813);
nor U1096 (N_1096,N_806,N_854);
nor U1097 (N_1097,N_881,N_926);
or U1098 (N_1098,N_916,N_908);
and U1099 (N_1099,N_944,N_925);
and U1100 (N_1100,N_962,N_833);
and U1101 (N_1101,N_872,N_829);
nand U1102 (N_1102,N_973,N_959);
xor U1103 (N_1103,N_989,N_819);
nor U1104 (N_1104,N_996,N_951);
or U1105 (N_1105,N_912,N_976);
nand U1106 (N_1106,N_946,N_961);
nor U1107 (N_1107,N_811,N_872);
nand U1108 (N_1108,N_856,N_841);
nor U1109 (N_1109,N_891,N_989);
and U1110 (N_1110,N_908,N_819);
nor U1111 (N_1111,N_993,N_954);
or U1112 (N_1112,N_880,N_946);
nand U1113 (N_1113,N_820,N_884);
nand U1114 (N_1114,N_931,N_839);
nor U1115 (N_1115,N_941,N_877);
nor U1116 (N_1116,N_871,N_820);
and U1117 (N_1117,N_814,N_944);
nor U1118 (N_1118,N_979,N_830);
xnor U1119 (N_1119,N_981,N_953);
xnor U1120 (N_1120,N_849,N_898);
nand U1121 (N_1121,N_908,N_889);
nand U1122 (N_1122,N_895,N_905);
xor U1123 (N_1123,N_903,N_879);
xnor U1124 (N_1124,N_993,N_944);
and U1125 (N_1125,N_995,N_970);
and U1126 (N_1126,N_885,N_918);
and U1127 (N_1127,N_890,N_845);
or U1128 (N_1128,N_927,N_875);
nor U1129 (N_1129,N_849,N_824);
nand U1130 (N_1130,N_807,N_953);
nand U1131 (N_1131,N_929,N_911);
nand U1132 (N_1132,N_906,N_890);
nor U1133 (N_1133,N_977,N_950);
nor U1134 (N_1134,N_822,N_862);
nor U1135 (N_1135,N_942,N_929);
xnor U1136 (N_1136,N_816,N_881);
xnor U1137 (N_1137,N_979,N_883);
nand U1138 (N_1138,N_959,N_974);
and U1139 (N_1139,N_882,N_908);
xor U1140 (N_1140,N_926,N_822);
nor U1141 (N_1141,N_873,N_961);
nand U1142 (N_1142,N_926,N_868);
xnor U1143 (N_1143,N_812,N_924);
nor U1144 (N_1144,N_968,N_967);
or U1145 (N_1145,N_906,N_992);
or U1146 (N_1146,N_992,N_873);
or U1147 (N_1147,N_877,N_982);
and U1148 (N_1148,N_934,N_843);
xnor U1149 (N_1149,N_804,N_982);
and U1150 (N_1150,N_999,N_847);
nand U1151 (N_1151,N_832,N_865);
nor U1152 (N_1152,N_859,N_975);
nor U1153 (N_1153,N_980,N_842);
xnor U1154 (N_1154,N_918,N_904);
and U1155 (N_1155,N_959,N_878);
or U1156 (N_1156,N_950,N_851);
and U1157 (N_1157,N_812,N_870);
nor U1158 (N_1158,N_879,N_872);
and U1159 (N_1159,N_865,N_853);
nand U1160 (N_1160,N_960,N_944);
nor U1161 (N_1161,N_997,N_921);
and U1162 (N_1162,N_858,N_906);
nand U1163 (N_1163,N_993,N_832);
nor U1164 (N_1164,N_840,N_862);
nand U1165 (N_1165,N_836,N_818);
xnor U1166 (N_1166,N_932,N_958);
xor U1167 (N_1167,N_927,N_831);
or U1168 (N_1168,N_879,N_914);
or U1169 (N_1169,N_938,N_901);
and U1170 (N_1170,N_981,N_889);
nor U1171 (N_1171,N_884,N_985);
or U1172 (N_1172,N_990,N_879);
or U1173 (N_1173,N_831,N_914);
xnor U1174 (N_1174,N_868,N_929);
nor U1175 (N_1175,N_933,N_951);
or U1176 (N_1176,N_853,N_958);
nand U1177 (N_1177,N_866,N_886);
and U1178 (N_1178,N_805,N_923);
nand U1179 (N_1179,N_856,N_989);
nor U1180 (N_1180,N_908,N_984);
nor U1181 (N_1181,N_928,N_827);
nand U1182 (N_1182,N_917,N_961);
nor U1183 (N_1183,N_898,N_817);
or U1184 (N_1184,N_870,N_816);
or U1185 (N_1185,N_952,N_916);
and U1186 (N_1186,N_854,N_936);
nand U1187 (N_1187,N_961,N_893);
nand U1188 (N_1188,N_818,N_817);
xor U1189 (N_1189,N_914,N_842);
and U1190 (N_1190,N_964,N_952);
nand U1191 (N_1191,N_993,N_923);
nand U1192 (N_1192,N_828,N_898);
xor U1193 (N_1193,N_914,N_807);
xnor U1194 (N_1194,N_950,N_805);
nor U1195 (N_1195,N_937,N_941);
nand U1196 (N_1196,N_847,N_955);
and U1197 (N_1197,N_826,N_944);
nand U1198 (N_1198,N_812,N_819);
xor U1199 (N_1199,N_985,N_855);
nor U1200 (N_1200,N_1199,N_1056);
nor U1201 (N_1201,N_1111,N_1063);
or U1202 (N_1202,N_1147,N_1191);
and U1203 (N_1203,N_1082,N_1070);
nor U1204 (N_1204,N_1169,N_1156);
or U1205 (N_1205,N_1061,N_1188);
and U1206 (N_1206,N_1010,N_1112);
nor U1207 (N_1207,N_1189,N_1001);
nor U1208 (N_1208,N_1119,N_1183);
or U1209 (N_1209,N_1033,N_1076);
or U1210 (N_1210,N_1013,N_1058);
and U1211 (N_1211,N_1159,N_1027);
or U1212 (N_1212,N_1190,N_1011);
and U1213 (N_1213,N_1185,N_1150);
and U1214 (N_1214,N_1025,N_1115);
nor U1215 (N_1215,N_1129,N_1122);
nand U1216 (N_1216,N_1073,N_1134);
nand U1217 (N_1217,N_1036,N_1162);
or U1218 (N_1218,N_1142,N_1153);
nor U1219 (N_1219,N_1087,N_1178);
and U1220 (N_1220,N_1007,N_1106);
nor U1221 (N_1221,N_1154,N_1037);
and U1222 (N_1222,N_1155,N_1044);
and U1223 (N_1223,N_1175,N_1004);
nor U1224 (N_1224,N_1020,N_1074);
xnor U1225 (N_1225,N_1014,N_1019);
nand U1226 (N_1226,N_1127,N_1021);
nand U1227 (N_1227,N_1006,N_1091);
xor U1228 (N_1228,N_1015,N_1085);
and U1229 (N_1229,N_1008,N_1078);
nor U1230 (N_1230,N_1077,N_1138);
and U1231 (N_1231,N_1103,N_1145);
xor U1232 (N_1232,N_1046,N_1184);
nand U1233 (N_1233,N_1179,N_1053);
and U1234 (N_1234,N_1090,N_1079);
nand U1235 (N_1235,N_1124,N_1132);
nand U1236 (N_1236,N_1003,N_1167);
or U1237 (N_1237,N_1170,N_1110);
nand U1238 (N_1238,N_1196,N_1049);
nor U1239 (N_1239,N_1118,N_1052);
xnor U1240 (N_1240,N_1104,N_1114);
and U1241 (N_1241,N_1038,N_1163);
or U1242 (N_1242,N_1113,N_1080);
nand U1243 (N_1243,N_1095,N_1187);
and U1244 (N_1244,N_1055,N_1140);
and U1245 (N_1245,N_1030,N_1093);
nor U1246 (N_1246,N_1041,N_1068);
nor U1247 (N_1247,N_1084,N_1094);
xnor U1248 (N_1248,N_1071,N_1133);
nor U1249 (N_1249,N_1128,N_1157);
and U1250 (N_1250,N_1005,N_1017);
nand U1251 (N_1251,N_1048,N_1139);
nor U1252 (N_1252,N_1125,N_1009);
or U1253 (N_1253,N_1149,N_1016);
nand U1254 (N_1254,N_1034,N_1018);
or U1255 (N_1255,N_1192,N_1160);
and U1256 (N_1256,N_1051,N_1059);
xnor U1257 (N_1257,N_1097,N_1144);
nand U1258 (N_1258,N_1035,N_1126);
or U1259 (N_1259,N_1174,N_1064);
nand U1260 (N_1260,N_1172,N_1152);
or U1261 (N_1261,N_1107,N_1171);
nand U1262 (N_1262,N_1148,N_1083);
and U1263 (N_1263,N_1062,N_1177);
xnor U1264 (N_1264,N_1026,N_1193);
or U1265 (N_1265,N_1173,N_1135);
or U1266 (N_1266,N_1143,N_1065);
nand U1267 (N_1267,N_1194,N_1197);
nor U1268 (N_1268,N_1101,N_1031);
and U1269 (N_1269,N_1168,N_1002);
or U1270 (N_1270,N_1120,N_1088);
and U1271 (N_1271,N_1102,N_1050);
or U1272 (N_1272,N_1166,N_1039);
nor U1273 (N_1273,N_1105,N_1131);
and U1274 (N_1274,N_1047,N_1000);
xor U1275 (N_1275,N_1069,N_1032);
nand U1276 (N_1276,N_1158,N_1057);
or U1277 (N_1277,N_1181,N_1060);
and U1278 (N_1278,N_1198,N_1141);
xor U1279 (N_1279,N_1180,N_1116);
nand U1280 (N_1280,N_1137,N_1151);
xnor U1281 (N_1281,N_1075,N_1023);
and U1282 (N_1282,N_1043,N_1024);
nor U1283 (N_1283,N_1054,N_1022);
or U1284 (N_1284,N_1045,N_1067);
and U1285 (N_1285,N_1098,N_1042);
xor U1286 (N_1286,N_1195,N_1100);
nand U1287 (N_1287,N_1176,N_1028);
and U1288 (N_1288,N_1092,N_1161);
nor U1289 (N_1289,N_1109,N_1123);
xor U1290 (N_1290,N_1086,N_1121);
and U1291 (N_1291,N_1182,N_1089);
xor U1292 (N_1292,N_1146,N_1117);
or U1293 (N_1293,N_1096,N_1066);
xor U1294 (N_1294,N_1029,N_1099);
nand U1295 (N_1295,N_1165,N_1040);
nand U1296 (N_1296,N_1012,N_1164);
nand U1297 (N_1297,N_1130,N_1072);
or U1298 (N_1298,N_1186,N_1136);
or U1299 (N_1299,N_1108,N_1081);
xnor U1300 (N_1300,N_1138,N_1021);
xor U1301 (N_1301,N_1162,N_1067);
or U1302 (N_1302,N_1019,N_1082);
or U1303 (N_1303,N_1120,N_1017);
nor U1304 (N_1304,N_1087,N_1026);
xor U1305 (N_1305,N_1089,N_1043);
and U1306 (N_1306,N_1145,N_1009);
or U1307 (N_1307,N_1182,N_1118);
xnor U1308 (N_1308,N_1069,N_1057);
and U1309 (N_1309,N_1043,N_1126);
xnor U1310 (N_1310,N_1084,N_1182);
and U1311 (N_1311,N_1186,N_1160);
or U1312 (N_1312,N_1099,N_1032);
nand U1313 (N_1313,N_1126,N_1168);
nand U1314 (N_1314,N_1003,N_1015);
nand U1315 (N_1315,N_1058,N_1039);
nor U1316 (N_1316,N_1096,N_1043);
nand U1317 (N_1317,N_1192,N_1196);
or U1318 (N_1318,N_1195,N_1125);
nor U1319 (N_1319,N_1090,N_1104);
or U1320 (N_1320,N_1028,N_1039);
or U1321 (N_1321,N_1053,N_1000);
nand U1322 (N_1322,N_1033,N_1080);
xnor U1323 (N_1323,N_1035,N_1121);
and U1324 (N_1324,N_1006,N_1103);
xnor U1325 (N_1325,N_1126,N_1173);
xnor U1326 (N_1326,N_1064,N_1168);
or U1327 (N_1327,N_1099,N_1022);
xnor U1328 (N_1328,N_1162,N_1107);
nor U1329 (N_1329,N_1141,N_1163);
and U1330 (N_1330,N_1102,N_1023);
and U1331 (N_1331,N_1073,N_1065);
nor U1332 (N_1332,N_1077,N_1125);
or U1333 (N_1333,N_1028,N_1159);
xor U1334 (N_1334,N_1196,N_1036);
nor U1335 (N_1335,N_1080,N_1007);
or U1336 (N_1336,N_1091,N_1078);
xor U1337 (N_1337,N_1092,N_1006);
and U1338 (N_1338,N_1075,N_1191);
nand U1339 (N_1339,N_1176,N_1045);
or U1340 (N_1340,N_1111,N_1056);
xor U1341 (N_1341,N_1060,N_1074);
or U1342 (N_1342,N_1021,N_1108);
nor U1343 (N_1343,N_1008,N_1091);
nor U1344 (N_1344,N_1122,N_1078);
nand U1345 (N_1345,N_1043,N_1174);
or U1346 (N_1346,N_1128,N_1040);
nand U1347 (N_1347,N_1001,N_1185);
nor U1348 (N_1348,N_1019,N_1115);
nor U1349 (N_1349,N_1139,N_1108);
or U1350 (N_1350,N_1022,N_1166);
nor U1351 (N_1351,N_1066,N_1081);
nor U1352 (N_1352,N_1168,N_1087);
or U1353 (N_1353,N_1110,N_1095);
and U1354 (N_1354,N_1142,N_1000);
xnor U1355 (N_1355,N_1030,N_1198);
nand U1356 (N_1356,N_1172,N_1179);
nor U1357 (N_1357,N_1118,N_1046);
nor U1358 (N_1358,N_1187,N_1054);
nor U1359 (N_1359,N_1049,N_1162);
nor U1360 (N_1360,N_1007,N_1120);
xnor U1361 (N_1361,N_1079,N_1125);
and U1362 (N_1362,N_1025,N_1154);
nor U1363 (N_1363,N_1124,N_1028);
xnor U1364 (N_1364,N_1023,N_1029);
or U1365 (N_1365,N_1076,N_1064);
and U1366 (N_1366,N_1063,N_1098);
xnor U1367 (N_1367,N_1147,N_1132);
xnor U1368 (N_1368,N_1074,N_1182);
nor U1369 (N_1369,N_1182,N_1145);
nor U1370 (N_1370,N_1060,N_1042);
xor U1371 (N_1371,N_1073,N_1004);
or U1372 (N_1372,N_1172,N_1170);
nand U1373 (N_1373,N_1128,N_1090);
xnor U1374 (N_1374,N_1102,N_1161);
nand U1375 (N_1375,N_1011,N_1117);
xor U1376 (N_1376,N_1066,N_1106);
nand U1377 (N_1377,N_1194,N_1017);
nand U1378 (N_1378,N_1024,N_1097);
nor U1379 (N_1379,N_1192,N_1069);
or U1380 (N_1380,N_1120,N_1039);
xor U1381 (N_1381,N_1127,N_1184);
nor U1382 (N_1382,N_1110,N_1194);
nand U1383 (N_1383,N_1180,N_1108);
nand U1384 (N_1384,N_1172,N_1197);
xor U1385 (N_1385,N_1067,N_1006);
nand U1386 (N_1386,N_1176,N_1041);
xor U1387 (N_1387,N_1033,N_1137);
and U1388 (N_1388,N_1066,N_1061);
or U1389 (N_1389,N_1127,N_1112);
xnor U1390 (N_1390,N_1176,N_1199);
nand U1391 (N_1391,N_1071,N_1197);
or U1392 (N_1392,N_1082,N_1119);
nand U1393 (N_1393,N_1198,N_1158);
nor U1394 (N_1394,N_1066,N_1014);
and U1395 (N_1395,N_1155,N_1166);
nand U1396 (N_1396,N_1067,N_1102);
xnor U1397 (N_1397,N_1163,N_1148);
xnor U1398 (N_1398,N_1060,N_1016);
nand U1399 (N_1399,N_1126,N_1023);
nand U1400 (N_1400,N_1360,N_1211);
nor U1401 (N_1401,N_1374,N_1258);
or U1402 (N_1402,N_1201,N_1383);
or U1403 (N_1403,N_1330,N_1262);
and U1404 (N_1404,N_1265,N_1340);
nand U1405 (N_1405,N_1333,N_1342);
or U1406 (N_1406,N_1396,N_1299);
xnor U1407 (N_1407,N_1274,N_1208);
nand U1408 (N_1408,N_1324,N_1369);
or U1409 (N_1409,N_1388,N_1259);
or U1410 (N_1410,N_1241,N_1243);
nand U1411 (N_1411,N_1361,N_1332);
nand U1412 (N_1412,N_1257,N_1203);
and U1413 (N_1413,N_1313,N_1267);
xor U1414 (N_1414,N_1338,N_1215);
nand U1415 (N_1415,N_1232,N_1287);
or U1416 (N_1416,N_1235,N_1285);
and U1417 (N_1417,N_1291,N_1379);
and U1418 (N_1418,N_1389,N_1331);
or U1419 (N_1419,N_1254,N_1205);
nand U1420 (N_1420,N_1206,N_1376);
xnor U1421 (N_1421,N_1349,N_1230);
nor U1422 (N_1422,N_1371,N_1236);
nor U1423 (N_1423,N_1398,N_1326);
nand U1424 (N_1424,N_1357,N_1352);
xor U1425 (N_1425,N_1377,N_1202);
nand U1426 (N_1426,N_1283,N_1221);
xor U1427 (N_1427,N_1271,N_1229);
nand U1428 (N_1428,N_1214,N_1218);
or U1429 (N_1429,N_1225,N_1204);
nand U1430 (N_1430,N_1370,N_1347);
xor U1431 (N_1431,N_1343,N_1295);
or U1432 (N_1432,N_1270,N_1336);
and U1433 (N_1433,N_1284,N_1269);
nor U1434 (N_1434,N_1216,N_1255);
or U1435 (N_1435,N_1280,N_1384);
xnor U1436 (N_1436,N_1226,N_1334);
nor U1437 (N_1437,N_1391,N_1213);
or U1438 (N_1438,N_1368,N_1309);
nor U1439 (N_1439,N_1301,N_1387);
and U1440 (N_1440,N_1231,N_1282);
nor U1441 (N_1441,N_1293,N_1339);
nor U1442 (N_1442,N_1253,N_1292);
or U1443 (N_1443,N_1308,N_1328);
nand U1444 (N_1444,N_1341,N_1335);
and U1445 (N_1445,N_1363,N_1234);
nand U1446 (N_1446,N_1264,N_1397);
or U1447 (N_1447,N_1224,N_1382);
nor U1448 (N_1448,N_1298,N_1260);
or U1449 (N_1449,N_1385,N_1277);
nand U1450 (N_1450,N_1325,N_1305);
and U1451 (N_1451,N_1312,N_1296);
or U1452 (N_1452,N_1300,N_1256);
xor U1453 (N_1453,N_1276,N_1275);
and U1454 (N_1454,N_1210,N_1302);
nand U1455 (N_1455,N_1273,N_1367);
or U1456 (N_1456,N_1237,N_1307);
and U1457 (N_1457,N_1245,N_1322);
and U1458 (N_1458,N_1329,N_1288);
nand U1459 (N_1459,N_1294,N_1355);
nor U1460 (N_1460,N_1266,N_1217);
and U1461 (N_1461,N_1278,N_1219);
xnor U1462 (N_1462,N_1320,N_1344);
nor U1463 (N_1463,N_1303,N_1392);
nand U1464 (N_1464,N_1372,N_1381);
nor U1465 (N_1465,N_1317,N_1318);
nand U1466 (N_1466,N_1263,N_1358);
or U1467 (N_1467,N_1261,N_1227);
nor U1468 (N_1468,N_1321,N_1390);
nand U1469 (N_1469,N_1378,N_1200);
nor U1470 (N_1470,N_1223,N_1399);
and U1471 (N_1471,N_1290,N_1356);
nor U1472 (N_1472,N_1314,N_1286);
nand U1473 (N_1473,N_1346,N_1393);
nand U1474 (N_1474,N_1362,N_1310);
xor U1475 (N_1475,N_1375,N_1327);
xnor U1476 (N_1476,N_1297,N_1351);
xor U1477 (N_1477,N_1315,N_1323);
nor U1478 (N_1478,N_1238,N_1242);
nor U1479 (N_1479,N_1289,N_1239);
and U1480 (N_1480,N_1373,N_1395);
or U1481 (N_1481,N_1251,N_1348);
and U1482 (N_1482,N_1247,N_1350);
xnor U1483 (N_1483,N_1268,N_1359);
nand U1484 (N_1484,N_1380,N_1345);
xor U1485 (N_1485,N_1304,N_1209);
or U1486 (N_1486,N_1281,N_1366);
and U1487 (N_1487,N_1220,N_1279);
nand U1488 (N_1488,N_1252,N_1248);
or U1489 (N_1489,N_1337,N_1354);
nor U1490 (N_1490,N_1365,N_1306);
and U1491 (N_1491,N_1353,N_1246);
xnor U1492 (N_1492,N_1394,N_1250);
xor U1493 (N_1493,N_1319,N_1386);
or U1494 (N_1494,N_1212,N_1249);
nor U1495 (N_1495,N_1240,N_1207);
xnor U1496 (N_1496,N_1228,N_1244);
nand U1497 (N_1497,N_1316,N_1364);
and U1498 (N_1498,N_1272,N_1233);
nand U1499 (N_1499,N_1222,N_1311);
and U1500 (N_1500,N_1223,N_1288);
xnor U1501 (N_1501,N_1329,N_1266);
and U1502 (N_1502,N_1268,N_1263);
nand U1503 (N_1503,N_1221,N_1312);
and U1504 (N_1504,N_1333,N_1252);
or U1505 (N_1505,N_1256,N_1268);
xor U1506 (N_1506,N_1310,N_1247);
nor U1507 (N_1507,N_1360,N_1210);
nand U1508 (N_1508,N_1260,N_1342);
xor U1509 (N_1509,N_1367,N_1309);
and U1510 (N_1510,N_1230,N_1267);
xor U1511 (N_1511,N_1305,N_1242);
or U1512 (N_1512,N_1235,N_1363);
and U1513 (N_1513,N_1251,N_1276);
and U1514 (N_1514,N_1336,N_1231);
or U1515 (N_1515,N_1369,N_1312);
or U1516 (N_1516,N_1274,N_1397);
nand U1517 (N_1517,N_1386,N_1286);
nor U1518 (N_1518,N_1293,N_1360);
or U1519 (N_1519,N_1238,N_1355);
nor U1520 (N_1520,N_1306,N_1395);
xnor U1521 (N_1521,N_1312,N_1295);
nand U1522 (N_1522,N_1252,N_1210);
nand U1523 (N_1523,N_1350,N_1268);
nor U1524 (N_1524,N_1269,N_1391);
or U1525 (N_1525,N_1290,N_1267);
nand U1526 (N_1526,N_1226,N_1248);
nor U1527 (N_1527,N_1394,N_1387);
nor U1528 (N_1528,N_1325,N_1331);
nor U1529 (N_1529,N_1234,N_1378);
or U1530 (N_1530,N_1283,N_1206);
and U1531 (N_1531,N_1230,N_1202);
nand U1532 (N_1532,N_1232,N_1234);
nand U1533 (N_1533,N_1302,N_1200);
or U1534 (N_1534,N_1359,N_1248);
nand U1535 (N_1535,N_1320,N_1225);
xor U1536 (N_1536,N_1338,N_1264);
nand U1537 (N_1537,N_1352,N_1220);
and U1538 (N_1538,N_1373,N_1338);
xnor U1539 (N_1539,N_1257,N_1322);
or U1540 (N_1540,N_1348,N_1302);
or U1541 (N_1541,N_1375,N_1348);
xor U1542 (N_1542,N_1368,N_1244);
nand U1543 (N_1543,N_1395,N_1360);
nor U1544 (N_1544,N_1341,N_1222);
nor U1545 (N_1545,N_1269,N_1247);
and U1546 (N_1546,N_1238,N_1277);
and U1547 (N_1547,N_1264,N_1299);
nand U1548 (N_1548,N_1256,N_1396);
xnor U1549 (N_1549,N_1319,N_1213);
nand U1550 (N_1550,N_1239,N_1213);
nor U1551 (N_1551,N_1251,N_1387);
and U1552 (N_1552,N_1210,N_1319);
xor U1553 (N_1553,N_1305,N_1399);
and U1554 (N_1554,N_1328,N_1257);
xnor U1555 (N_1555,N_1264,N_1274);
xor U1556 (N_1556,N_1351,N_1383);
and U1557 (N_1557,N_1223,N_1228);
nand U1558 (N_1558,N_1280,N_1371);
nand U1559 (N_1559,N_1283,N_1395);
nor U1560 (N_1560,N_1272,N_1347);
or U1561 (N_1561,N_1281,N_1345);
or U1562 (N_1562,N_1294,N_1321);
and U1563 (N_1563,N_1228,N_1260);
xor U1564 (N_1564,N_1271,N_1300);
nor U1565 (N_1565,N_1332,N_1209);
and U1566 (N_1566,N_1365,N_1374);
or U1567 (N_1567,N_1279,N_1322);
and U1568 (N_1568,N_1201,N_1380);
and U1569 (N_1569,N_1275,N_1289);
nand U1570 (N_1570,N_1221,N_1295);
nor U1571 (N_1571,N_1233,N_1369);
nand U1572 (N_1572,N_1207,N_1239);
xor U1573 (N_1573,N_1213,N_1374);
or U1574 (N_1574,N_1359,N_1217);
nand U1575 (N_1575,N_1368,N_1251);
or U1576 (N_1576,N_1389,N_1271);
xnor U1577 (N_1577,N_1203,N_1328);
or U1578 (N_1578,N_1264,N_1321);
xor U1579 (N_1579,N_1276,N_1330);
nor U1580 (N_1580,N_1243,N_1211);
nand U1581 (N_1581,N_1238,N_1201);
xnor U1582 (N_1582,N_1269,N_1367);
or U1583 (N_1583,N_1245,N_1338);
xor U1584 (N_1584,N_1354,N_1341);
or U1585 (N_1585,N_1397,N_1236);
nand U1586 (N_1586,N_1246,N_1374);
or U1587 (N_1587,N_1323,N_1316);
nand U1588 (N_1588,N_1386,N_1373);
nand U1589 (N_1589,N_1200,N_1262);
or U1590 (N_1590,N_1313,N_1354);
xnor U1591 (N_1591,N_1319,N_1257);
xor U1592 (N_1592,N_1373,N_1276);
nand U1593 (N_1593,N_1349,N_1327);
xnor U1594 (N_1594,N_1219,N_1201);
and U1595 (N_1595,N_1389,N_1303);
and U1596 (N_1596,N_1297,N_1230);
nor U1597 (N_1597,N_1242,N_1325);
or U1598 (N_1598,N_1340,N_1214);
and U1599 (N_1599,N_1377,N_1258);
or U1600 (N_1600,N_1557,N_1574);
xnor U1601 (N_1601,N_1404,N_1530);
nand U1602 (N_1602,N_1582,N_1413);
xnor U1603 (N_1603,N_1570,N_1412);
nor U1604 (N_1604,N_1426,N_1512);
nor U1605 (N_1605,N_1478,N_1408);
nand U1606 (N_1606,N_1499,N_1553);
xor U1607 (N_1607,N_1568,N_1581);
xor U1608 (N_1608,N_1435,N_1470);
nand U1609 (N_1609,N_1474,N_1416);
or U1610 (N_1610,N_1531,N_1491);
or U1611 (N_1611,N_1538,N_1479);
or U1612 (N_1612,N_1493,N_1497);
nand U1613 (N_1613,N_1539,N_1540);
or U1614 (N_1614,N_1431,N_1502);
nor U1615 (N_1615,N_1584,N_1503);
xnor U1616 (N_1616,N_1496,N_1547);
nand U1617 (N_1617,N_1505,N_1415);
and U1618 (N_1618,N_1549,N_1575);
or U1619 (N_1619,N_1508,N_1562);
nand U1620 (N_1620,N_1556,N_1514);
nor U1621 (N_1621,N_1564,N_1545);
xnor U1622 (N_1622,N_1509,N_1518);
nand U1623 (N_1623,N_1465,N_1536);
nand U1624 (N_1624,N_1537,N_1550);
xor U1625 (N_1625,N_1421,N_1488);
and U1626 (N_1626,N_1551,N_1469);
or U1627 (N_1627,N_1464,N_1513);
xor U1628 (N_1628,N_1472,N_1487);
nor U1629 (N_1629,N_1592,N_1458);
xor U1630 (N_1630,N_1429,N_1593);
nand U1631 (N_1631,N_1579,N_1427);
and U1632 (N_1632,N_1495,N_1520);
xnor U1633 (N_1633,N_1554,N_1437);
xnor U1634 (N_1634,N_1566,N_1444);
and U1635 (N_1635,N_1489,N_1462);
and U1636 (N_1636,N_1451,N_1494);
nand U1637 (N_1637,N_1477,N_1484);
nor U1638 (N_1638,N_1596,N_1482);
nand U1639 (N_1639,N_1403,N_1559);
nor U1640 (N_1640,N_1485,N_1442);
nor U1641 (N_1641,N_1527,N_1500);
xnor U1642 (N_1642,N_1468,N_1585);
or U1643 (N_1643,N_1449,N_1511);
nand U1644 (N_1644,N_1587,N_1519);
nand U1645 (N_1645,N_1591,N_1534);
nor U1646 (N_1646,N_1565,N_1409);
nand U1647 (N_1647,N_1483,N_1523);
nand U1648 (N_1648,N_1586,N_1590);
and U1649 (N_1649,N_1419,N_1561);
nor U1650 (N_1650,N_1422,N_1441);
xnor U1651 (N_1651,N_1490,N_1480);
and U1652 (N_1652,N_1595,N_1434);
and U1653 (N_1653,N_1457,N_1571);
xor U1654 (N_1654,N_1414,N_1443);
nand U1655 (N_1655,N_1417,N_1439);
and U1656 (N_1656,N_1572,N_1418);
and U1657 (N_1657,N_1507,N_1406);
nor U1658 (N_1658,N_1525,N_1460);
nor U1659 (N_1659,N_1510,N_1576);
nor U1660 (N_1660,N_1552,N_1411);
or U1661 (N_1661,N_1467,N_1446);
nand U1662 (N_1662,N_1501,N_1448);
nand U1663 (N_1663,N_1425,N_1498);
xnor U1664 (N_1664,N_1577,N_1473);
or U1665 (N_1665,N_1588,N_1533);
and U1666 (N_1666,N_1459,N_1521);
nor U1667 (N_1667,N_1567,N_1445);
xnor U1668 (N_1668,N_1528,N_1420);
nor U1669 (N_1669,N_1455,N_1453);
nand U1670 (N_1670,N_1516,N_1555);
nand U1671 (N_1671,N_1517,N_1532);
xor U1672 (N_1672,N_1546,N_1529);
and U1673 (N_1673,N_1436,N_1447);
xor U1674 (N_1674,N_1504,N_1526);
and U1675 (N_1675,N_1463,N_1430);
nand U1676 (N_1676,N_1589,N_1405);
nand U1677 (N_1677,N_1548,N_1524);
and U1678 (N_1678,N_1428,N_1410);
nor U1679 (N_1679,N_1580,N_1456);
xor U1680 (N_1680,N_1438,N_1407);
or U1681 (N_1681,N_1558,N_1573);
xnor U1682 (N_1682,N_1452,N_1535);
or U1683 (N_1683,N_1599,N_1515);
or U1684 (N_1684,N_1583,N_1433);
xor U1685 (N_1685,N_1544,N_1542);
or U1686 (N_1686,N_1506,N_1424);
or U1687 (N_1687,N_1400,N_1563);
nand U1688 (N_1688,N_1440,N_1466);
xnor U1689 (N_1689,N_1481,N_1486);
nand U1690 (N_1690,N_1569,N_1454);
and U1691 (N_1691,N_1450,N_1492);
nor U1692 (N_1692,N_1401,N_1476);
nand U1693 (N_1693,N_1560,N_1432);
and U1694 (N_1694,N_1475,N_1578);
and U1695 (N_1695,N_1423,N_1541);
and U1696 (N_1696,N_1402,N_1461);
nand U1697 (N_1697,N_1594,N_1598);
nor U1698 (N_1698,N_1543,N_1597);
nand U1699 (N_1699,N_1471,N_1522);
and U1700 (N_1700,N_1498,N_1504);
xnor U1701 (N_1701,N_1429,N_1514);
nor U1702 (N_1702,N_1556,N_1500);
nor U1703 (N_1703,N_1413,N_1486);
nor U1704 (N_1704,N_1559,N_1597);
xnor U1705 (N_1705,N_1587,N_1400);
nor U1706 (N_1706,N_1533,N_1464);
nand U1707 (N_1707,N_1559,N_1507);
or U1708 (N_1708,N_1434,N_1497);
nand U1709 (N_1709,N_1480,N_1487);
or U1710 (N_1710,N_1537,N_1560);
or U1711 (N_1711,N_1518,N_1535);
nor U1712 (N_1712,N_1451,N_1419);
xnor U1713 (N_1713,N_1522,N_1411);
and U1714 (N_1714,N_1546,N_1591);
and U1715 (N_1715,N_1465,N_1587);
xor U1716 (N_1716,N_1471,N_1524);
and U1717 (N_1717,N_1444,N_1574);
or U1718 (N_1718,N_1400,N_1455);
nand U1719 (N_1719,N_1584,N_1438);
nor U1720 (N_1720,N_1541,N_1532);
nor U1721 (N_1721,N_1410,N_1500);
nor U1722 (N_1722,N_1505,N_1451);
nor U1723 (N_1723,N_1402,N_1547);
nand U1724 (N_1724,N_1483,N_1496);
xnor U1725 (N_1725,N_1413,N_1478);
nand U1726 (N_1726,N_1497,N_1579);
and U1727 (N_1727,N_1538,N_1565);
or U1728 (N_1728,N_1589,N_1515);
xor U1729 (N_1729,N_1519,N_1569);
or U1730 (N_1730,N_1441,N_1421);
and U1731 (N_1731,N_1548,N_1483);
nor U1732 (N_1732,N_1450,N_1405);
or U1733 (N_1733,N_1442,N_1471);
nor U1734 (N_1734,N_1513,N_1437);
xor U1735 (N_1735,N_1564,N_1491);
nor U1736 (N_1736,N_1596,N_1578);
and U1737 (N_1737,N_1407,N_1440);
and U1738 (N_1738,N_1593,N_1507);
or U1739 (N_1739,N_1514,N_1473);
or U1740 (N_1740,N_1402,N_1434);
nand U1741 (N_1741,N_1440,N_1511);
nand U1742 (N_1742,N_1452,N_1451);
xor U1743 (N_1743,N_1599,N_1457);
xnor U1744 (N_1744,N_1450,N_1538);
nor U1745 (N_1745,N_1461,N_1442);
xnor U1746 (N_1746,N_1593,N_1564);
nand U1747 (N_1747,N_1592,N_1542);
nor U1748 (N_1748,N_1514,N_1422);
nand U1749 (N_1749,N_1429,N_1503);
and U1750 (N_1750,N_1575,N_1531);
nand U1751 (N_1751,N_1500,N_1530);
xor U1752 (N_1752,N_1584,N_1542);
nand U1753 (N_1753,N_1444,N_1428);
nor U1754 (N_1754,N_1541,N_1413);
or U1755 (N_1755,N_1480,N_1489);
nand U1756 (N_1756,N_1462,N_1580);
xor U1757 (N_1757,N_1523,N_1560);
nand U1758 (N_1758,N_1561,N_1467);
nand U1759 (N_1759,N_1556,N_1411);
nand U1760 (N_1760,N_1519,N_1580);
and U1761 (N_1761,N_1513,N_1424);
or U1762 (N_1762,N_1475,N_1592);
nor U1763 (N_1763,N_1576,N_1445);
nand U1764 (N_1764,N_1493,N_1562);
and U1765 (N_1765,N_1552,N_1518);
nand U1766 (N_1766,N_1570,N_1591);
xnor U1767 (N_1767,N_1498,N_1415);
nand U1768 (N_1768,N_1561,N_1509);
xnor U1769 (N_1769,N_1498,N_1576);
nor U1770 (N_1770,N_1571,N_1558);
xnor U1771 (N_1771,N_1430,N_1487);
xor U1772 (N_1772,N_1466,N_1545);
nor U1773 (N_1773,N_1593,N_1555);
and U1774 (N_1774,N_1471,N_1578);
nand U1775 (N_1775,N_1416,N_1460);
nand U1776 (N_1776,N_1469,N_1533);
nand U1777 (N_1777,N_1569,N_1598);
and U1778 (N_1778,N_1484,N_1586);
xor U1779 (N_1779,N_1428,N_1577);
xor U1780 (N_1780,N_1474,N_1496);
nor U1781 (N_1781,N_1587,N_1428);
xor U1782 (N_1782,N_1437,N_1561);
nand U1783 (N_1783,N_1478,N_1420);
xnor U1784 (N_1784,N_1400,N_1424);
or U1785 (N_1785,N_1407,N_1443);
xor U1786 (N_1786,N_1436,N_1565);
and U1787 (N_1787,N_1523,N_1510);
and U1788 (N_1788,N_1562,N_1492);
xor U1789 (N_1789,N_1597,N_1573);
or U1790 (N_1790,N_1523,N_1459);
nand U1791 (N_1791,N_1411,N_1510);
xor U1792 (N_1792,N_1574,N_1504);
nand U1793 (N_1793,N_1433,N_1567);
nor U1794 (N_1794,N_1530,N_1470);
and U1795 (N_1795,N_1486,N_1434);
or U1796 (N_1796,N_1557,N_1500);
nand U1797 (N_1797,N_1593,N_1528);
nand U1798 (N_1798,N_1538,N_1447);
and U1799 (N_1799,N_1505,N_1404);
xnor U1800 (N_1800,N_1604,N_1698);
nand U1801 (N_1801,N_1607,N_1793);
nor U1802 (N_1802,N_1752,N_1614);
nor U1803 (N_1803,N_1675,N_1726);
nand U1804 (N_1804,N_1662,N_1703);
or U1805 (N_1805,N_1684,N_1668);
xnor U1806 (N_1806,N_1782,N_1620);
and U1807 (N_1807,N_1742,N_1762);
or U1808 (N_1808,N_1695,N_1720);
nor U1809 (N_1809,N_1729,N_1718);
nand U1810 (N_1810,N_1640,N_1738);
or U1811 (N_1811,N_1725,N_1716);
nor U1812 (N_1812,N_1658,N_1778);
nor U1813 (N_1813,N_1717,N_1615);
nor U1814 (N_1814,N_1643,N_1753);
and U1815 (N_1815,N_1637,N_1669);
nor U1816 (N_1816,N_1736,N_1722);
nor U1817 (N_1817,N_1727,N_1653);
and U1818 (N_1818,N_1734,N_1665);
and U1819 (N_1819,N_1747,N_1744);
nand U1820 (N_1820,N_1699,N_1602);
nor U1821 (N_1821,N_1619,N_1706);
nor U1822 (N_1822,N_1644,N_1608);
xor U1823 (N_1823,N_1701,N_1693);
nand U1824 (N_1824,N_1764,N_1783);
and U1825 (N_1825,N_1690,N_1775);
or U1826 (N_1826,N_1745,N_1618);
or U1827 (N_1827,N_1623,N_1768);
xor U1828 (N_1828,N_1642,N_1645);
and U1829 (N_1829,N_1700,N_1677);
nor U1830 (N_1830,N_1621,N_1622);
nand U1831 (N_1831,N_1664,N_1611);
and U1832 (N_1832,N_1647,N_1633);
and U1833 (N_1833,N_1617,N_1624);
nor U1834 (N_1834,N_1648,N_1650);
nor U1835 (N_1835,N_1681,N_1603);
nor U1836 (N_1836,N_1606,N_1777);
or U1837 (N_1837,N_1794,N_1679);
or U1838 (N_1838,N_1638,N_1678);
xnor U1839 (N_1839,N_1613,N_1692);
xor U1840 (N_1840,N_1760,N_1799);
or U1841 (N_1841,N_1723,N_1763);
nand U1842 (N_1842,N_1773,N_1661);
nand U1843 (N_1843,N_1691,N_1771);
xnor U1844 (N_1844,N_1672,N_1770);
nand U1845 (N_1845,N_1656,N_1707);
xor U1846 (N_1846,N_1733,N_1766);
or U1847 (N_1847,N_1758,N_1715);
and U1848 (N_1848,N_1781,N_1756);
nand U1849 (N_1849,N_1680,N_1641);
xor U1850 (N_1850,N_1765,N_1780);
nor U1851 (N_1851,N_1676,N_1787);
nor U1852 (N_1852,N_1731,N_1772);
and U1853 (N_1853,N_1712,N_1746);
nor U1854 (N_1854,N_1612,N_1688);
and U1855 (N_1855,N_1797,N_1735);
or U1856 (N_1856,N_1790,N_1769);
xnor U1857 (N_1857,N_1711,N_1697);
or U1858 (N_1858,N_1748,N_1635);
xnor U1859 (N_1859,N_1687,N_1646);
nor U1860 (N_1860,N_1774,N_1761);
xnor U1861 (N_1861,N_1728,N_1719);
nor U1862 (N_1862,N_1696,N_1755);
nor U1863 (N_1863,N_1632,N_1751);
xnor U1864 (N_1864,N_1791,N_1673);
nor U1865 (N_1865,N_1610,N_1659);
and U1866 (N_1866,N_1710,N_1627);
xor U1867 (N_1867,N_1737,N_1657);
nor U1868 (N_1868,N_1709,N_1743);
xor U1869 (N_1869,N_1601,N_1702);
xor U1870 (N_1870,N_1651,N_1685);
xor U1871 (N_1871,N_1667,N_1795);
xor U1872 (N_1872,N_1630,N_1750);
nor U1873 (N_1873,N_1605,N_1713);
nor U1874 (N_1874,N_1721,N_1704);
and U1875 (N_1875,N_1759,N_1798);
xnor U1876 (N_1876,N_1626,N_1796);
or U1877 (N_1877,N_1767,N_1776);
nor U1878 (N_1878,N_1724,N_1705);
and U1879 (N_1879,N_1749,N_1739);
and U1880 (N_1880,N_1784,N_1740);
nand U1881 (N_1881,N_1694,N_1654);
or U1882 (N_1882,N_1741,N_1785);
nand U1883 (N_1883,N_1666,N_1682);
or U1884 (N_1884,N_1786,N_1663);
xnor U1885 (N_1885,N_1639,N_1789);
nand U1886 (N_1886,N_1625,N_1636);
and U1887 (N_1887,N_1779,N_1788);
and U1888 (N_1888,N_1649,N_1600);
nor U1889 (N_1889,N_1754,N_1730);
nor U1890 (N_1890,N_1634,N_1670);
xor U1891 (N_1891,N_1674,N_1652);
nor U1892 (N_1892,N_1792,N_1683);
or U1893 (N_1893,N_1689,N_1660);
nor U1894 (N_1894,N_1628,N_1629);
nand U1895 (N_1895,N_1708,N_1671);
nand U1896 (N_1896,N_1732,N_1686);
xnor U1897 (N_1897,N_1714,N_1631);
nor U1898 (N_1898,N_1616,N_1655);
and U1899 (N_1899,N_1609,N_1757);
nor U1900 (N_1900,N_1737,N_1779);
and U1901 (N_1901,N_1657,N_1776);
and U1902 (N_1902,N_1700,N_1694);
nor U1903 (N_1903,N_1730,N_1792);
nor U1904 (N_1904,N_1736,N_1655);
and U1905 (N_1905,N_1758,N_1634);
or U1906 (N_1906,N_1624,N_1711);
nand U1907 (N_1907,N_1763,N_1776);
nor U1908 (N_1908,N_1662,N_1613);
xnor U1909 (N_1909,N_1778,N_1649);
nand U1910 (N_1910,N_1626,N_1631);
nand U1911 (N_1911,N_1652,N_1684);
and U1912 (N_1912,N_1785,N_1674);
and U1913 (N_1913,N_1793,N_1749);
and U1914 (N_1914,N_1623,N_1722);
nand U1915 (N_1915,N_1770,N_1794);
xnor U1916 (N_1916,N_1789,N_1666);
nand U1917 (N_1917,N_1653,N_1666);
or U1918 (N_1918,N_1669,N_1790);
xnor U1919 (N_1919,N_1779,N_1735);
or U1920 (N_1920,N_1640,N_1614);
and U1921 (N_1921,N_1602,N_1669);
nand U1922 (N_1922,N_1712,N_1621);
nor U1923 (N_1923,N_1605,N_1685);
and U1924 (N_1924,N_1712,N_1626);
nor U1925 (N_1925,N_1741,N_1655);
nor U1926 (N_1926,N_1688,N_1692);
nor U1927 (N_1927,N_1635,N_1722);
or U1928 (N_1928,N_1601,N_1682);
or U1929 (N_1929,N_1701,N_1656);
or U1930 (N_1930,N_1760,N_1640);
or U1931 (N_1931,N_1675,N_1682);
and U1932 (N_1932,N_1756,N_1793);
nor U1933 (N_1933,N_1691,N_1671);
nor U1934 (N_1934,N_1635,N_1612);
nand U1935 (N_1935,N_1618,N_1765);
or U1936 (N_1936,N_1647,N_1743);
xnor U1937 (N_1937,N_1705,N_1712);
nor U1938 (N_1938,N_1638,N_1631);
and U1939 (N_1939,N_1700,N_1637);
or U1940 (N_1940,N_1713,N_1648);
nand U1941 (N_1941,N_1737,N_1633);
and U1942 (N_1942,N_1680,N_1763);
or U1943 (N_1943,N_1657,N_1721);
xor U1944 (N_1944,N_1697,N_1670);
nor U1945 (N_1945,N_1672,N_1671);
xnor U1946 (N_1946,N_1723,N_1740);
nor U1947 (N_1947,N_1684,N_1661);
nand U1948 (N_1948,N_1773,N_1746);
and U1949 (N_1949,N_1772,N_1777);
xor U1950 (N_1950,N_1624,N_1673);
nor U1951 (N_1951,N_1650,N_1704);
xnor U1952 (N_1952,N_1620,N_1660);
nor U1953 (N_1953,N_1705,N_1720);
nor U1954 (N_1954,N_1715,N_1705);
or U1955 (N_1955,N_1787,N_1721);
and U1956 (N_1956,N_1630,N_1610);
nand U1957 (N_1957,N_1680,N_1644);
xnor U1958 (N_1958,N_1677,N_1719);
xor U1959 (N_1959,N_1737,N_1733);
nand U1960 (N_1960,N_1678,N_1773);
nand U1961 (N_1961,N_1634,N_1666);
nor U1962 (N_1962,N_1656,N_1603);
xor U1963 (N_1963,N_1720,N_1621);
and U1964 (N_1964,N_1733,N_1779);
xor U1965 (N_1965,N_1731,N_1680);
xnor U1966 (N_1966,N_1701,N_1686);
nand U1967 (N_1967,N_1779,N_1755);
and U1968 (N_1968,N_1783,N_1640);
nand U1969 (N_1969,N_1736,N_1702);
nor U1970 (N_1970,N_1687,N_1761);
xnor U1971 (N_1971,N_1657,N_1711);
nor U1972 (N_1972,N_1600,N_1774);
nor U1973 (N_1973,N_1752,N_1647);
xnor U1974 (N_1974,N_1763,N_1742);
xor U1975 (N_1975,N_1659,N_1753);
or U1976 (N_1976,N_1650,N_1674);
xor U1977 (N_1977,N_1720,N_1657);
nand U1978 (N_1978,N_1658,N_1642);
or U1979 (N_1979,N_1734,N_1649);
nor U1980 (N_1980,N_1742,N_1741);
nor U1981 (N_1981,N_1615,N_1667);
xor U1982 (N_1982,N_1704,N_1737);
and U1983 (N_1983,N_1600,N_1724);
xnor U1984 (N_1984,N_1744,N_1717);
xor U1985 (N_1985,N_1642,N_1611);
nand U1986 (N_1986,N_1716,N_1758);
or U1987 (N_1987,N_1637,N_1646);
nor U1988 (N_1988,N_1604,N_1648);
xor U1989 (N_1989,N_1642,N_1698);
xnor U1990 (N_1990,N_1715,N_1734);
and U1991 (N_1991,N_1746,N_1692);
or U1992 (N_1992,N_1721,N_1668);
and U1993 (N_1993,N_1669,N_1758);
nand U1994 (N_1994,N_1764,N_1614);
or U1995 (N_1995,N_1632,N_1655);
and U1996 (N_1996,N_1601,N_1786);
nor U1997 (N_1997,N_1622,N_1717);
or U1998 (N_1998,N_1729,N_1680);
xor U1999 (N_1999,N_1691,N_1790);
nor U2000 (N_2000,N_1981,N_1914);
nor U2001 (N_2001,N_1877,N_1922);
xor U2002 (N_2002,N_1955,N_1898);
nand U2003 (N_2003,N_1863,N_1856);
nand U2004 (N_2004,N_1990,N_1968);
or U2005 (N_2005,N_1857,N_1829);
nor U2006 (N_2006,N_1805,N_1943);
xor U2007 (N_2007,N_1889,N_1906);
and U2008 (N_2008,N_1984,N_1939);
xor U2009 (N_2009,N_1995,N_1975);
or U2010 (N_2010,N_1989,N_1985);
nor U2011 (N_2011,N_1897,N_1954);
and U2012 (N_2012,N_1841,N_1960);
and U2013 (N_2013,N_1813,N_1896);
or U2014 (N_2014,N_1997,N_1959);
nor U2015 (N_2015,N_1957,N_1835);
nor U2016 (N_2016,N_1903,N_1900);
or U2017 (N_2017,N_1840,N_1883);
nand U2018 (N_2018,N_1811,N_1938);
nor U2019 (N_2019,N_1942,N_1801);
xor U2020 (N_2020,N_1983,N_1916);
xor U2021 (N_2021,N_1923,N_1929);
nand U2022 (N_2022,N_1918,N_1937);
nor U2023 (N_2023,N_1845,N_1988);
nand U2024 (N_2024,N_1904,N_1850);
or U2025 (N_2025,N_1927,N_1825);
or U2026 (N_2026,N_1982,N_1854);
or U2027 (N_2027,N_1996,N_1969);
xnor U2028 (N_2028,N_1860,N_1820);
and U2029 (N_2029,N_1974,N_1991);
nor U2030 (N_2030,N_1928,N_1999);
xor U2031 (N_2031,N_1902,N_1802);
xor U2032 (N_2032,N_1882,N_1930);
nand U2033 (N_2033,N_1800,N_1888);
or U2034 (N_2034,N_1915,N_1879);
or U2035 (N_2035,N_1891,N_1893);
nor U2036 (N_2036,N_1876,N_1839);
nand U2037 (N_2037,N_1807,N_1947);
nor U2038 (N_2038,N_1972,N_1907);
and U2039 (N_2039,N_1842,N_1998);
or U2040 (N_2040,N_1932,N_1818);
and U2041 (N_2041,N_1867,N_1936);
or U2042 (N_2042,N_1980,N_1886);
xor U2043 (N_2043,N_1961,N_1884);
nand U2044 (N_2044,N_1912,N_1806);
or U2045 (N_2045,N_1865,N_1837);
nor U2046 (N_2046,N_1803,N_1862);
and U2047 (N_2047,N_1941,N_1987);
nor U2048 (N_2048,N_1855,N_1951);
or U2049 (N_2049,N_1872,N_1852);
and U2050 (N_2050,N_1965,N_1919);
xnor U2051 (N_2051,N_1973,N_1821);
or U2052 (N_2052,N_1828,N_1817);
and U2053 (N_2053,N_1926,N_1869);
xnor U2054 (N_2054,N_1958,N_1940);
nor U2055 (N_2055,N_1962,N_1830);
nor U2056 (N_2056,N_1808,N_1868);
xnor U2057 (N_2057,N_1831,N_1870);
or U2058 (N_2058,N_1910,N_1809);
or U2059 (N_2059,N_1881,N_1953);
or U2060 (N_2060,N_1946,N_1812);
and U2061 (N_2061,N_1956,N_1895);
nand U2062 (N_2062,N_1866,N_1949);
xnor U2063 (N_2063,N_1966,N_1851);
or U2064 (N_2064,N_1925,N_1992);
nor U2065 (N_2065,N_1899,N_1933);
nand U2066 (N_2066,N_1950,N_1846);
xnor U2067 (N_2067,N_1977,N_1834);
and U2068 (N_2068,N_1901,N_1843);
and U2069 (N_2069,N_1909,N_1978);
xnor U2070 (N_2070,N_1993,N_1848);
xnor U2071 (N_2071,N_1967,N_1948);
xnor U2072 (N_2072,N_1836,N_1894);
nor U2073 (N_2073,N_1924,N_1952);
or U2074 (N_2074,N_1964,N_1804);
nand U2075 (N_2075,N_1885,N_1847);
or U2076 (N_2076,N_1832,N_1810);
nand U2077 (N_2077,N_1890,N_1861);
or U2078 (N_2078,N_1822,N_1931);
and U2079 (N_2079,N_1911,N_1963);
xor U2080 (N_2080,N_1874,N_1849);
and U2081 (N_2081,N_1908,N_1853);
and U2082 (N_2082,N_1838,N_1816);
nor U2083 (N_2083,N_1875,N_1880);
or U2084 (N_2084,N_1892,N_1819);
xnor U2085 (N_2085,N_1858,N_1844);
or U2086 (N_2086,N_1935,N_1833);
xnor U2087 (N_2087,N_1878,N_1994);
and U2088 (N_2088,N_1920,N_1887);
nand U2089 (N_2089,N_1971,N_1944);
xnor U2090 (N_2090,N_1827,N_1979);
nor U2091 (N_2091,N_1976,N_1864);
or U2092 (N_2092,N_1859,N_1824);
nor U2093 (N_2093,N_1921,N_1871);
xnor U2094 (N_2094,N_1826,N_1905);
and U2095 (N_2095,N_1815,N_1917);
nand U2096 (N_2096,N_1934,N_1873);
xor U2097 (N_2097,N_1986,N_1823);
or U2098 (N_2098,N_1970,N_1913);
nor U2099 (N_2099,N_1945,N_1814);
nor U2100 (N_2100,N_1974,N_1993);
nor U2101 (N_2101,N_1949,N_1867);
or U2102 (N_2102,N_1969,N_1856);
and U2103 (N_2103,N_1905,N_1870);
xnor U2104 (N_2104,N_1927,N_1821);
xor U2105 (N_2105,N_1987,N_1823);
nor U2106 (N_2106,N_1904,N_1916);
nor U2107 (N_2107,N_1912,N_1875);
xor U2108 (N_2108,N_1899,N_1852);
nor U2109 (N_2109,N_1969,N_1939);
and U2110 (N_2110,N_1879,N_1907);
xnor U2111 (N_2111,N_1849,N_1998);
nand U2112 (N_2112,N_1880,N_1879);
nor U2113 (N_2113,N_1837,N_1957);
and U2114 (N_2114,N_1950,N_1988);
xor U2115 (N_2115,N_1801,N_1850);
xor U2116 (N_2116,N_1955,N_1813);
xor U2117 (N_2117,N_1936,N_1978);
xnor U2118 (N_2118,N_1940,N_1804);
nand U2119 (N_2119,N_1965,N_1983);
and U2120 (N_2120,N_1839,N_1937);
nor U2121 (N_2121,N_1988,N_1981);
or U2122 (N_2122,N_1834,N_1837);
xor U2123 (N_2123,N_1947,N_1841);
nor U2124 (N_2124,N_1842,N_1910);
and U2125 (N_2125,N_1922,N_1971);
xor U2126 (N_2126,N_1938,N_1974);
and U2127 (N_2127,N_1912,N_1855);
or U2128 (N_2128,N_1931,N_1802);
nor U2129 (N_2129,N_1806,N_1844);
xor U2130 (N_2130,N_1881,N_1910);
xnor U2131 (N_2131,N_1952,N_1959);
and U2132 (N_2132,N_1803,N_1821);
xnor U2133 (N_2133,N_1929,N_1933);
or U2134 (N_2134,N_1900,N_1922);
nand U2135 (N_2135,N_1850,N_1837);
nand U2136 (N_2136,N_1947,N_1885);
and U2137 (N_2137,N_1933,N_1948);
or U2138 (N_2138,N_1919,N_1805);
and U2139 (N_2139,N_1919,N_1818);
nand U2140 (N_2140,N_1956,N_1873);
and U2141 (N_2141,N_1898,N_1827);
and U2142 (N_2142,N_1956,N_1865);
nand U2143 (N_2143,N_1870,N_1879);
nor U2144 (N_2144,N_1925,N_1934);
xor U2145 (N_2145,N_1922,N_1800);
nand U2146 (N_2146,N_1988,N_1887);
or U2147 (N_2147,N_1973,N_1849);
nand U2148 (N_2148,N_1905,N_1973);
nand U2149 (N_2149,N_1918,N_1807);
or U2150 (N_2150,N_1949,N_1833);
and U2151 (N_2151,N_1923,N_1804);
xnor U2152 (N_2152,N_1911,N_1908);
nor U2153 (N_2153,N_1818,N_1821);
xnor U2154 (N_2154,N_1817,N_1912);
and U2155 (N_2155,N_1936,N_1844);
xor U2156 (N_2156,N_1899,N_1884);
xnor U2157 (N_2157,N_1871,N_1940);
or U2158 (N_2158,N_1984,N_1870);
xnor U2159 (N_2159,N_1838,N_1804);
nand U2160 (N_2160,N_1814,N_1903);
and U2161 (N_2161,N_1863,N_1861);
and U2162 (N_2162,N_1818,N_1930);
and U2163 (N_2163,N_1873,N_1932);
xnor U2164 (N_2164,N_1854,N_1912);
nand U2165 (N_2165,N_1817,N_1898);
and U2166 (N_2166,N_1896,N_1877);
nand U2167 (N_2167,N_1975,N_1996);
nand U2168 (N_2168,N_1875,N_1873);
nand U2169 (N_2169,N_1996,N_1961);
nand U2170 (N_2170,N_1878,N_1973);
nor U2171 (N_2171,N_1832,N_1879);
nor U2172 (N_2172,N_1930,N_1947);
or U2173 (N_2173,N_1856,N_1877);
nand U2174 (N_2174,N_1889,N_1962);
or U2175 (N_2175,N_1995,N_1958);
xnor U2176 (N_2176,N_1909,N_1923);
xnor U2177 (N_2177,N_1953,N_1938);
nand U2178 (N_2178,N_1896,N_1873);
xor U2179 (N_2179,N_1877,N_1812);
or U2180 (N_2180,N_1855,N_1969);
nand U2181 (N_2181,N_1818,N_1879);
and U2182 (N_2182,N_1807,N_1840);
nor U2183 (N_2183,N_1982,N_1984);
nor U2184 (N_2184,N_1861,N_1820);
xor U2185 (N_2185,N_1919,N_1929);
xor U2186 (N_2186,N_1838,N_1852);
xor U2187 (N_2187,N_1943,N_1816);
xor U2188 (N_2188,N_1924,N_1975);
and U2189 (N_2189,N_1872,N_1905);
or U2190 (N_2190,N_1949,N_1895);
or U2191 (N_2191,N_1818,N_1867);
xor U2192 (N_2192,N_1811,N_1931);
nand U2193 (N_2193,N_1887,N_1998);
nor U2194 (N_2194,N_1971,N_1943);
nand U2195 (N_2195,N_1963,N_1852);
and U2196 (N_2196,N_1913,N_1991);
xor U2197 (N_2197,N_1977,N_1957);
xor U2198 (N_2198,N_1817,N_1848);
nor U2199 (N_2199,N_1825,N_1930);
and U2200 (N_2200,N_2017,N_2088);
nor U2201 (N_2201,N_2117,N_2010);
nand U2202 (N_2202,N_2182,N_2173);
or U2203 (N_2203,N_2176,N_2107);
or U2204 (N_2204,N_2085,N_2067);
or U2205 (N_2205,N_2160,N_2167);
xnor U2206 (N_2206,N_2188,N_2004);
nand U2207 (N_2207,N_2022,N_2080);
and U2208 (N_2208,N_2081,N_2034);
nand U2209 (N_2209,N_2174,N_2123);
nor U2210 (N_2210,N_2165,N_2073);
xor U2211 (N_2211,N_2156,N_2185);
nor U2212 (N_2212,N_2166,N_2133);
nand U2213 (N_2213,N_2039,N_2001);
or U2214 (N_2214,N_2051,N_2075);
nor U2215 (N_2215,N_2105,N_2198);
or U2216 (N_2216,N_2020,N_2037);
and U2217 (N_2217,N_2016,N_2029);
and U2218 (N_2218,N_2122,N_2152);
and U2219 (N_2219,N_2153,N_2045);
nor U2220 (N_2220,N_2097,N_2128);
or U2221 (N_2221,N_2145,N_2148);
and U2222 (N_2222,N_2026,N_2106);
nand U2223 (N_2223,N_2030,N_2099);
nor U2224 (N_2224,N_2191,N_2177);
nor U2225 (N_2225,N_2157,N_2008);
xor U2226 (N_2226,N_2007,N_2102);
xor U2227 (N_2227,N_2072,N_2052);
nor U2228 (N_2228,N_2086,N_2044);
or U2229 (N_2229,N_2035,N_2094);
or U2230 (N_2230,N_2028,N_2129);
or U2231 (N_2231,N_2084,N_2048);
nand U2232 (N_2232,N_2135,N_2083);
xnor U2233 (N_2233,N_2125,N_2141);
or U2234 (N_2234,N_2127,N_2015);
nor U2235 (N_2235,N_2151,N_2070);
and U2236 (N_2236,N_2064,N_2025);
and U2237 (N_2237,N_2013,N_2058);
or U2238 (N_2238,N_2056,N_2074);
or U2239 (N_2239,N_2047,N_2131);
nor U2240 (N_2240,N_2071,N_2042);
and U2241 (N_2241,N_2012,N_2104);
nor U2242 (N_2242,N_2009,N_2187);
and U2243 (N_2243,N_2053,N_2114);
or U2244 (N_2244,N_2049,N_2168);
nand U2245 (N_2245,N_2065,N_2118);
or U2246 (N_2246,N_2190,N_2093);
nor U2247 (N_2247,N_2055,N_2040);
nor U2248 (N_2248,N_2124,N_2103);
nand U2249 (N_2249,N_2003,N_2021);
and U2250 (N_2250,N_2046,N_2041);
or U2251 (N_2251,N_2054,N_2147);
nor U2252 (N_2252,N_2090,N_2197);
and U2253 (N_2253,N_2139,N_2199);
and U2254 (N_2254,N_2130,N_2179);
nor U2255 (N_2255,N_2100,N_2171);
xnor U2256 (N_2256,N_2180,N_2134);
nand U2257 (N_2257,N_2050,N_2120);
nor U2258 (N_2258,N_2032,N_2043);
nor U2259 (N_2259,N_2061,N_2178);
nor U2260 (N_2260,N_2110,N_2169);
nor U2261 (N_2261,N_2138,N_2091);
xor U2262 (N_2262,N_2079,N_2066);
and U2263 (N_2263,N_2150,N_2140);
nand U2264 (N_2264,N_2121,N_2101);
xor U2265 (N_2265,N_2158,N_2143);
or U2266 (N_2266,N_2126,N_2144);
nor U2267 (N_2267,N_2115,N_2024);
and U2268 (N_2268,N_2186,N_2059);
nor U2269 (N_2269,N_2132,N_2108);
and U2270 (N_2270,N_2057,N_2027);
xnor U2271 (N_2271,N_2078,N_2112);
xnor U2272 (N_2272,N_2089,N_2060);
nor U2273 (N_2273,N_2006,N_2155);
nand U2274 (N_2274,N_2095,N_2000);
or U2275 (N_2275,N_2069,N_2076);
nor U2276 (N_2276,N_2113,N_2068);
nor U2277 (N_2277,N_2011,N_2005);
or U2278 (N_2278,N_2137,N_2014);
and U2279 (N_2279,N_2194,N_2175);
nor U2280 (N_2280,N_2096,N_2136);
xor U2281 (N_2281,N_2098,N_2163);
and U2282 (N_2282,N_2195,N_2149);
xnor U2283 (N_2283,N_2062,N_2192);
nand U2284 (N_2284,N_2116,N_2087);
nor U2285 (N_2285,N_2142,N_2193);
nand U2286 (N_2286,N_2183,N_2170);
or U2287 (N_2287,N_2184,N_2196);
nor U2288 (N_2288,N_2038,N_2036);
and U2289 (N_2289,N_2092,N_2161);
xnor U2290 (N_2290,N_2162,N_2109);
nand U2291 (N_2291,N_2018,N_2031);
xor U2292 (N_2292,N_2119,N_2023);
or U2293 (N_2293,N_2063,N_2002);
xnor U2294 (N_2294,N_2019,N_2164);
xor U2295 (N_2295,N_2172,N_2033);
xor U2296 (N_2296,N_2111,N_2082);
or U2297 (N_2297,N_2159,N_2146);
and U2298 (N_2298,N_2181,N_2189);
xor U2299 (N_2299,N_2077,N_2154);
nor U2300 (N_2300,N_2160,N_2071);
xnor U2301 (N_2301,N_2007,N_2171);
nor U2302 (N_2302,N_2185,N_2169);
or U2303 (N_2303,N_2174,N_2143);
and U2304 (N_2304,N_2173,N_2198);
nor U2305 (N_2305,N_2139,N_2134);
or U2306 (N_2306,N_2026,N_2021);
nor U2307 (N_2307,N_2142,N_2124);
xnor U2308 (N_2308,N_2069,N_2009);
nand U2309 (N_2309,N_2014,N_2111);
nand U2310 (N_2310,N_2027,N_2170);
and U2311 (N_2311,N_2055,N_2143);
nor U2312 (N_2312,N_2052,N_2132);
xor U2313 (N_2313,N_2096,N_2121);
and U2314 (N_2314,N_2019,N_2179);
and U2315 (N_2315,N_2041,N_2146);
and U2316 (N_2316,N_2097,N_2079);
nor U2317 (N_2317,N_2074,N_2002);
nand U2318 (N_2318,N_2145,N_2116);
xnor U2319 (N_2319,N_2152,N_2176);
nand U2320 (N_2320,N_2117,N_2182);
nand U2321 (N_2321,N_2085,N_2043);
xor U2322 (N_2322,N_2172,N_2131);
xor U2323 (N_2323,N_2165,N_2009);
xnor U2324 (N_2324,N_2038,N_2142);
xor U2325 (N_2325,N_2136,N_2112);
nor U2326 (N_2326,N_2175,N_2111);
nor U2327 (N_2327,N_2090,N_2140);
nor U2328 (N_2328,N_2080,N_2174);
and U2329 (N_2329,N_2151,N_2191);
and U2330 (N_2330,N_2160,N_2133);
xor U2331 (N_2331,N_2126,N_2116);
nand U2332 (N_2332,N_2159,N_2078);
nand U2333 (N_2333,N_2075,N_2139);
and U2334 (N_2334,N_2048,N_2039);
or U2335 (N_2335,N_2106,N_2028);
xnor U2336 (N_2336,N_2051,N_2019);
xnor U2337 (N_2337,N_2027,N_2034);
nand U2338 (N_2338,N_2170,N_2084);
and U2339 (N_2339,N_2091,N_2016);
or U2340 (N_2340,N_2173,N_2145);
xor U2341 (N_2341,N_2114,N_2131);
or U2342 (N_2342,N_2044,N_2026);
nand U2343 (N_2343,N_2013,N_2039);
or U2344 (N_2344,N_2059,N_2014);
xor U2345 (N_2345,N_2062,N_2083);
and U2346 (N_2346,N_2065,N_2143);
and U2347 (N_2347,N_2193,N_2018);
nor U2348 (N_2348,N_2162,N_2174);
or U2349 (N_2349,N_2111,N_2108);
or U2350 (N_2350,N_2182,N_2184);
nand U2351 (N_2351,N_2104,N_2005);
xor U2352 (N_2352,N_2036,N_2069);
nand U2353 (N_2353,N_2122,N_2096);
xnor U2354 (N_2354,N_2066,N_2091);
nor U2355 (N_2355,N_2182,N_2187);
or U2356 (N_2356,N_2130,N_2172);
nand U2357 (N_2357,N_2154,N_2005);
or U2358 (N_2358,N_2047,N_2092);
and U2359 (N_2359,N_2191,N_2045);
nand U2360 (N_2360,N_2055,N_2060);
nand U2361 (N_2361,N_2021,N_2119);
or U2362 (N_2362,N_2078,N_2077);
nand U2363 (N_2363,N_2043,N_2128);
nand U2364 (N_2364,N_2090,N_2076);
xor U2365 (N_2365,N_2033,N_2008);
xor U2366 (N_2366,N_2034,N_2057);
nand U2367 (N_2367,N_2053,N_2062);
nor U2368 (N_2368,N_2114,N_2176);
and U2369 (N_2369,N_2085,N_2129);
nor U2370 (N_2370,N_2062,N_2112);
xor U2371 (N_2371,N_2177,N_2195);
nor U2372 (N_2372,N_2008,N_2123);
and U2373 (N_2373,N_2130,N_2021);
or U2374 (N_2374,N_2072,N_2194);
xnor U2375 (N_2375,N_2187,N_2046);
nand U2376 (N_2376,N_2183,N_2172);
and U2377 (N_2377,N_2097,N_2043);
and U2378 (N_2378,N_2067,N_2176);
or U2379 (N_2379,N_2004,N_2002);
and U2380 (N_2380,N_2188,N_2046);
nand U2381 (N_2381,N_2076,N_2048);
or U2382 (N_2382,N_2128,N_2000);
xnor U2383 (N_2383,N_2184,N_2001);
xor U2384 (N_2384,N_2176,N_2106);
nand U2385 (N_2385,N_2082,N_2127);
nor U2386 (N_2386,N_2102,N_2088);
nor U2387 (N_2387,N_2008,N_2110);
nor U2388 (N_2388,N_2055,N_2164);
and U2389 (N_2389,N_2102,N_2182);
nand U2390 (N_2390,N_2125,N_2102);
nor U2391 (N_2391,N_2168,N_2111);
or U2392 (N_2392,N_2039,N_2044);
or U2393 (N_2393,N_2115,N_2137);
xor U2394 (N_2394,N_2179,N_2191);
nand U2395 (N_2395,N_2043,N_2088);
and U2396 (N_2396,N_2070,N_2181);
nand U2397 (N_2397,N_2067,N_2154);
nor U2398 (N_2398,N_2059,N_2011);
and U2399 (N_2399,N_2095,N_2172);
and U2400 (N_2400,N_2386,N_2337);
or U2401 (N_2401,N_2294,N_2293);
or U2402 (N_2402,N_2332,N_2308);
nor U2403 (N_2403,N_2322,N_2343);
xor U2404 (N_2404,N_2315,N_2301);
or U2405 (N_2405,N_2360,N_2388);
or U2406 (N_2406,N_2346,N_2350);
nor U2407 (N_2407,N_2354,N_2238);
nor U2408 (N_2408,N_2200,N_2280);
or U2409 (N_2409,N_2230,N_2314);
nand U2410 (N_2410,N_2362,N_2275);
or U2411 (N_2411,N_2368,N_2390);
or U2412 (N_2412,N_2380,N_2222);
nand U2413 (N_2413,N_2252,N_2313);
xor U2414 (N_2414,N_2374,N_2338);
or U2415 (N_2415,N_2299,N_2377);
xnor U2416 (N_2416,N_2334,N_2341);
nand U2417 (N_2417,N_2273,N_2209);
xnor U2418 (N_2418,N_2364,N_2292);
xnor U2419 (N_2419,N_2210,N_2361);
nand U2420 (N_2420,N_2353,N_2286);
and U2421 (N_2421,N_2305,N_2223);
and U2422 (N_2422,N_2216,N_2336);
xor U2423 (N_2423,N_2318,N_2225);
or U2424 (N_2424,N_2381,N_2249);
or U2425 (N_2425,N_2247,N_2309);
and U2426 (N_2426,N_2207,N_2234);
nor U2427 (N_2427,N_2300,N_2291);
nor U2428 (N_2428,N_2373,N_2269);
nor U2429 (N_2429,N_2383,N_2329);
nand U2430 (N_2430,N_2363,N_2296);
nor U2431 (N_2431,N_2370,N_2260);
xnor U2432 (N_2432,N_2358,N_2297);
or U2433 (N_2433,N_2344,N_2250);
nand U2434 (N_2434,N_2226,N_2303);
xor U2435 (N_2435,N_2352,N_2319);
nand U2436 (N_2436,N_2239,N_2317);
nand U2437 (N_2437,N_2320,N_2257);
xnor U2438 (N_2438,N_2212,N_2202);
or U2439 (N_2439,N_2399,N_2262);
xnor U2440 (N_2440,N_2235,N_2393);
nor U2441 (N_2441,N_2316,N_2342);
or U2442 (N_2442,N_2295,N_2227);
and U2443 (N_2443,N_2274,N_2345);
or U2444 (N_2444,N_2288,N_2371);
nor U2445 (N_2445,N_2214,N_2276);
nand U2446 (N_2446,N_2351,N_2347);
nor U2447 (N_2447,N_2339,N_2271);
or U2448 (N_2448,N_2365,N_2289);
nor U2449 (N_2449,N_2233,N_2311);
and U2450 (N_2450,N_2281,N_2391);
or U2451 (N_2451,N_2228,N_2253);
nor U2452 (N_2452,N_2265,N_2256);
or U2453 (N_2453,N_2355,N_2201);
nand U2454 (N_2454,N_2213,N_2392);
and U2455 (N_2455,N_2323,N_2325);
or U2456 (N_2456,N_2298,N_2387);
xor U2457 (N_2457,N_2282,N_2217);
or U2458 (N_2458,N_2397,N_2335);
xor U2459 (N_2459,N_2221,N_2330);
and U2460 (N_2460,N_2204,N_2307);
and U2461 (N_2461,N_2268,N_2278);
xor U2462 (N_2462,N_2236,N_2272);
and U2463 (N_2463,N_2333,N_2283);
and U2464 (N_2464,N_2266,N_2264);
and U2465 (N_2465,N_2378,N_2395);
nand U2466 (N_2466,N_2287,N_2220);
xnor U2467 (N_2467,N_2348,N_2331);
nand U2468 (N_2468,N_2254,N_2394);
or U2469 (N_2469,N_2321,N_2328);
nand U2470 (N_2470,N_2205,N_2219);
xor U2471 (N_2471,N_2243,N_2246);
or U2472 (N_2472,N_2208,N_2284);
xnor U2473 (N_2473,N_2259,N_2306);
and U2474 (N_2474,N_2327,N_2385);
or U2475 (N_2475,N_2375,N_2324);
nor U2476 (N_2476,N_2224,N_2251);
xor U2477 (N_2477,N_2240,N_2237);
or U2478 (N_2478,N_2267,N_2367);
nand U2479 (N_2479,N_2203,N_2244);
xor U2480 (N_2480,N_2263,N_2326);
nand U2481 (N_2481,N_2242,N_2270);
nor U2482 (N_2482,N_2232,N_2245);
xor U2483 (N_2483,N_2372,N_2277);
and U2484 (N_2484,N_2379,N_2382);
and U2485 (N_2485,N_2229,N_2279);
xnor U2486 (N_2486,N_2215,N_2231);
nor U2487 (N_2487,N_2359,N_2356);
or U2488 (N_2488,N_2349,N_2211);
nand U2489 (N_2489,N_2218,N_2376);
or U2490 (N_2490,N_2357,N_2248);
nand U2491 (N_2491,N_2389,N_2261);
xor U2492 (N_2492,N_2285,N_2312);
or U2493 (N_2493,N_2398,N_2310);
or U2494 (N_2494,N_2366,N_2384);
or U2495 (N_2495,N_2255,N_2396);
nand U2496 (N_2496,N_2369,N_2241);
xor U2497 (N_2497,N_2206,N_2290);
or U2498 (N_2498,N_2258,N_2304);
xnor U2499 (N_2499,N_2302,N_2340);
xor U2500 (N_2500,N_2291,N_2263);
nor U2501 (N_2501,N_2220,N_2204);
and U2502 (N_2502,N_2244,N_2283);
or U2503 (N_2503,N_2256,N_2291);
and U2504 (N_2504,N_2321,N_2209);
and U2505 (N_2505,N_2258,N_2399);
and U2506 (N_2506,N_2350,N_2384);
or U2507 (N_2507,N_2297,N_2324);
nor U2508 (N_2508,N_2228,N_2306);
and U2509 (N_2509,N_2274,N_2311);
nor U2510 (N_2510,N_2325,N_2363);
nor U2511 (N_2511,N_2242,N_2299);
xnor U2512 (N_2512,N_2214,N_2337);
nor U2513 (N_2513,N_2229,N_2240);
and U2514 (N_2514,N_2347,N_2392);
xnor U2515 (N_2515,N_2359,N_2210);
or U2516 (N_2516,N_2379,N_2283);
nand U2517 (N_2517,N_2236,N_2351);
xor U2518 (N_2518,N_2332,N_2206);
xor U2519 (N_2519,N_2333,N_2275);
and U2520 (N_2520,N_2366,N_2323);
xnor U2521 (N_2521,N_2202,N_2219);
or U2522 (N_2522,N_2210,N_2343);
or U2523 (N_2523,N_2297,N_2300);
or U2524 (N_2524,N_2212,N_2363);
nor U2525 (N_2525,N_2214,N_2310);
and U2526 (N_2526,N_2356,N_2333);
and U2527 (N_2527,N_2225,N_2272);
xnor U2528 (N_2528,N_2235,N_2273);
nand U2529 (N_2529,N_2287,N_2211);
or U2530 (N_2530,N_2376,N_2306);
xor U2531 (N_2531,N_2258,N_2353);
or U2532 (N_2532,N_2397,N_2323);
nand U2533 (N_2533,N_2338,N_2235);
or U2534 (N_2534,N_2271,N_2200);
or U2535 (N_2535,N_2313,N_2334);
nor U2536 (N_2536,N_2289,N_2342);
nor U2537 (N_2537,N_2257,N_2306);
xnor U2538 (N_2538,N_2255,N_2377);
xor U2539 (N_2539,N_2200,N_2241);
nor U2540 (N_2540,N_2379,N_2251);
and U2541 (N_2541,N_2392,N_2344);
and U2542 (N_2542,N_2366,N_2282);
nor U2543 (N_2543,N_2239,N_2213);
nand U2544 (N_2544,N_2337,N_2270);
and U2545 (N_2545,N_2365,N_2301);
nor U2546 (N_2546,N_2249,N_2289);
nand U2547 (N_2547,N_2242,N_2356);
nand U2548 (N_2548,N_2255,N_2391);
xnor U2549 (N_2549,N_2372,N_2324);
xnor U2550 (N_2550,N_2341,N_2217);
and U2551 (N_2551,N_2202,N_2375);
and U2552 (N_2552,N_2358,N_2241);
nand U2553 (N_2553,N_2247,N_2371);
and U2554 (N_2554,N_2225,N_2208);
or U2555 (N_2555,N_2389,N_2235);
and U2556 (N_2556,N_2347,N_2238);
nor U2557 (N_2557,N_2352,N_2272);
xnor U2558 (N_2558,N_2399,N_2334);
and U2559 (N_2559,N_2346,N_2367);
nor U2560 (N_2560,N_2277,N_2276);
or U2561 (N_2561,N_2256,N_2334);
or U2562 (N_2562,N_2292,N_2272);
nand U2563 (N_2563,N_2282,N_2273);
nor U2564 (N_2564,N_2395,N_2315);
or U2565 (N_2565,N_2353,N_2306);
nor U2566 (N_2566,N_2239,N_2241);
nor U2567 (N_2567,N_2255,N_2236);
and U2568 (N_2568,N_2392,N_2336);
xnor U2569 (N_2569,N_2279,N_2246);
nand U2570 (N_2570,N_2237,N_2246);
or U2571 (N_2571,N_2359,N_2243);
nor U2572 (N_2572,N_2366,N_2231);
nand U2573 (N_2573,N_2303,N_2356);
nand U2574 (N_2574,N_2235,N_2262);
nand U2575 (N_2575,N_2302,N_2217);
xor U2576 (N_2576,N_2387,N_2327);
or U2577 (N_2577,N_2356,N_2345);
xor U2578 (N_2578,N_2244,N_2312);
nor U2579 (N_2579,N_2237,N_2261);
xnor U2580 (N_2580,N_2258,N_2295);
xnor U2581 (N_2581,N_2204,N_2242);
nor U2582 (N_2582,N_2350,N_2200);
or U2583 (N_2583,N_2330,N_2309);
nand U2584 (N_2584,N_2283,N_2215);
nand U2585 (N_2585,N_2240,N_2246);
and U2586 (N_2586,N_2350,N_2275);
xor U2587 (N_2587,N_2252,N_2255);
nor U2588 (N_2588,N_2284,N_2280);
nand U2589 (N_2589,N_2317,N_2262);
or U2590 (N_2590,N_2227,N_2356);
xor U2591 (N_2591,N_2222,N_2371);
xor U2592 (N_2592,N_2333,N_2342);
xnor U2593 (N_2593,N_2242,N_2284);
nand U2594 (N_2594,N_2304,N_2238);
nor U2595 (N_2595,N_2233,N_2201);
nor U2596 (N_2596,N_2251,N_2246);
nor U2597 (N_2597,N_2200,N_2317);
nor U2598 (N_2598,N_2367,N_2331);
or U2599 (N_2599,N_2356,N_2258);
or U2600 (N_2600,N_2442,N_2500);
nand U2601 (N_2601,N_2559,N_2493);
xor U2602 (N_2602,N_2553,N_2562);
nand U2603 (N_2603,N_2534,N_2456);
and U2604 (N_2604,N_2517,N_2549);
and U2605 (N_2605,N_2418,N_2461);
and U2606 (N_2606,N_2505,N_2573);
nor U2607 (N_2607,N_2544,N_2536);
or U2608 (N_2608,N_2514,N_2574);
xnor U2609 (N_2609,N_2581,N_2464);
and U2610 (N_2610,N_2492,N_2498);
xnor U2611 (N_2611,N_2524,N_2585);
and U2612 (N_2612,N_2484,N_2474);
nand U2613 (N_2613,N_2413,N_2402);
and U2614 (N_2614,N_2589,N_2576);
and U2615 (N_2615,N_2421,N_2583);
or U2616 (N_2616,N_2482,N_2508);
and U2617 (N_2617,N_2566,N_2584);
or U2618 (N_2618,N_2494,N_2506);
nor U2619 (N_2619,N_2444,N_2588);
nor U2620 (N_2620,N_2570,N_2441);
xor U2621 (N_2621,N_2522,N_2507);
and U2622 (N_2622,N_2422,N_2569);
nand U2623 (N_2623,N_2543,N_2470);
or U2624 (N_2624,N_2460,N_2410);
nor U2625 (N_2625,N_2438,N_2480);
and U2626 (N_2626,N_2586,N_2533);
or U2627 (N_2627,N_2490,N_2530);
nand U2628 (N_2628,N_2459,N_2556);
or U2629 (N_2629,N_2511,N_2405);
and U2630 (N_2630,N_2582,N_2451);
nor U2631 (N_2631,N_2516,N_2579);
xnor U2632 (N_2632,N_2551,N_2535);
or U2633 (N_2633,N_2593,N_2590);
nand U2634 (N_2634,N_2479,N_2434);
or U2635 (N_2635,N_2497,N_2538);
and U2636 (N_2636,N_2412,N_2564);
nand U2637 (N_2637,N_2489,N_2599);
and U2638 (N_2638,N_2546,N_2427);
nand U2639 (N_2639,N_2515,N_2430);
nand U2640 (N_2640,N_2528,N_2469);
nor U2641 (N_2641,N_2597,N_2414);
nor U2642 (N_2642,N_2453,N_2567);
nand U2643 (N_2643,N_2446,N_2529);
and U2644 (N_2644,N_2445,N_2554);
nor U2645 (N_2645,N_2443,N_2425);
and U2646 (N_2646,N_2495,N_2488);
nand U2647 (N_2647,N_2423,N_2548);
or U2648 (N_2648,N_2435,N_2407);
or U2649 (N_2649,N_2424,N_2431);
nor U2650 (N_2650,N_2577,N_2555);
nor U2651 (N_2651,N_2478,N_2416);
nand U2652 (N_2652,N_2518,N_2452);
and U2653 (N_2653,N_2578,N_2447);
and U2654 (N_2654,N_2448,N_2545);
nand U2655 (N_2655,N_2513,N_2429);
or U2656 (N_2656,N_2542,N_2531);
nand U2657 (N_2657,N_2419,N_2592);
and U2658 (N_2658,N_2400,N_2510);
xnor U2659 (N_2659,N_2501,N_2472);
xnor U2660 (N_2660,N_2415,N_2466);
nor U2661 (N_2661,N_2468,N_2454);
and U2662 (N_2662,N_2409,N_2455);
or U2663 (N_2663,N_2557,N_2580);
nand U2664 (N_2664,N_2532,N_2475);
xor U2665 (N_2665,N_2572,N_2449);
and U2666 (N_2666,N_2575,N_2526);
xnor U2667 (N_2667,N_2433,N_2439);
or U2668 (N_2668,N_2420,N_2591);
and U2669 (N_2669,N_2417,N_2561);
and U2670 (N_2670,N_2568,N_2560);
nand U2671 (N_2671,N_2457,N_2499);
and U2672 (N_2672,N_2558,N_2408);
xnor U2673 (N_2673,N_2440,N_2401);
and U2674 (N_2674,N_2403,N_2594);
nand U2675 (N_2675,N_2523,N_2502);
nand U2676 (N_2676,N_2476,N_2477);
nor U2677 (N_2677,N_2437,N_2487);
and U2678 (N_2678,N_2552,N_2547);
nand U2679 (N_2679,N_2436,N_2527);
nand U2680 (N_2680,N_2571,N_2458);
xnor U2681 (N_2681,N_2596,N_2509);
nor U2682 (N_2682,N_2483,N_2406);
nand U2683 (N_2683,N_2537,N_2565);
nand U2684 (N_2684,N_2550,N_2473);
and U2685 (N_2685,N_2450,N_2504);
xor U2686 (N_2686,N_2404,N_2595);
xor U2687 (N_2687,N_2598,N_2503);
and U2688 (N_2688,N_2521,N_2481);
and U2689 (N_2689,N_2467,N_2432);
nand U2690 (N_2690,N_2520,N_2471);
xor U2691 (N_2691,N_2465,N_2463);
nor U2692 (N_2692,N_2519,N_2540);
xnor U2693 (N_2693,N_2491,N_2539);
xor U2694 (N_2694,N_2485,N_2462);
xor U2695 (N_2695,N_2512,N_2563);
or U2696 (N_2696,N_2486,N_2411);
and U2697 (N_2697,N_2428,N_2426);
and U2698 (N_2698,N_2525,N_2587);
nor U2699 (N_2699,N_2541,N_2496);
or U2700 (N_2700,N_2432,N_2487);
or U2701 (N_2701,N_2477,N_2571);
nor U2702 (N_2702,N_2427,N_2558);
xor U2703 (N_2703,N_2441,N_2515);
nand U2704 (N_2704,N_2423,N_2436);
xor U2705 (N_2705,N_2501,N_2560);
or U2706 (N_2706,N_2527,N_2583);
or U2707 (N_2707,N_2404,N_2588);
nor U2708 (N_2708,N_2403,N_2596);
and U2709 (N_2709,N_2587,N_2407);
xor U2710 (N_2710,N_2554,N_2547);
xor U2711 (N_2711,N_2424,N_2455);
or U2712 (N_2712,N_2431,N_2405);
and U2713 (N_2713,N_2435,N_2483);
xnor U2714 (N_2714,N_2496,N_2413);
or U2715 (N_2715,N_2410,N_2589);
nand U2716 (N_2716,N_2581,N_2541);
nand U2717 (N_2717,N_2485,N_2428);
or U2718 (N_2718,N_2463,N_2493);
and U2719 (N_2719,N_2420,N_2528);
or U2720 (N_2720,N_2535,N_2431);
and U2721 (N_2721,N_2540,N_2470);
nand U2722 (N_2722,N_2450,N_2401);
or U2723 (N_2723,N_2538,N_2478);
nand U2724 (N_2724,N_2499,N_2544);
or U2725 (N_2725,N_2558,N_2435);
or U2726 (N_2726,N_2461,N_2465);
or U2727 (N_2727,N_2569,N_2428);
and U2728 (N_2728,N_2560,N_2546);
xnor U2729 (N_2729,N_2563,N_2545);
xor U2730 (N_2730,N_2542,N_2551);
nand U2731 (N_2731,N_2459,N_2438);
nand U2732 (N_2732,N_2479,N_2592);
nand U2733 (N_2733,N_2493,N_2478);
and U2734 (N_2734,N_2487,N_2577);
or U2735 (N_2735,N_2401,N_2575);
xor U2736 (N_2736,N_2588,N_2466);
xnor U2737 (N_2737,N_2408,N_2432);
nand U2738 (N_2738,N_2526,N_2480);
xor U2739 (N_2739,N_2495,N_2497);
xnor U2740 (N_2740,N_2456,N_2531);
and U2741 (N_2741,N_2441,N_2445);
xor U2742 (N_2742,N_2480,N_2527);
and U2743 (N_2743,N_2403,N_2493);
nor U2744 (N_2744,N_2486,N_2536);
and U2745 (N_2745,N_2466,N_2403);
and U2746 (N_2746,N_2583,N_2506);
nor U2747 (N_2747,N_2512,N_2470);
nor U2748 (N_2748,N_2450,N_2594);
xor U2749 (N_2749,N_2440,N_2461);
xor U2750 (N_2750,N_2446,N_2400);
nor U2751 (N_2751,N_2479,N_2459);
nand U2752 (N_2752,N_2477,N_2413);
and U2753 (N_2753,N_2400,N_2460);
xor U2754 (N_2754,N_2522,N_2576);
nand U2755 (N_2755,N_2568,N_2573);
and U2756 (N_2756,N_2479,N_2416);
xnor U2757 (N_2757,N_2487,N_2484);
nor U2758 (N_2758,N_2514,N_2479);
nor U2759 (N_2759,N_2459,N_2517);
or U2760 (N_2760,N_2549,N_2482);
and U2761 (N_2761,N_2517,N_2471);
nor U2762 (N_2762,N_2590,N_2468);
nor U2763 (N_2763,N_2470,N_2419);
and U2764 (N_2764,N_2437,N_2405);
and U2765 (N_2765,N_2523,N_2576);
and U2766 (N_2766,N_2588,N_2586);
xnor U2767 (N_2767,N_2541,N_2402);
or U2768 (N_2768,N_2537,N_2521);
and U2769 (N_2769,N_2599,N_2567);
nor U2770 (N_2770,N_2517,N_2442);
or U2771 (N_2771,N_2448,N_2555);
and U2772 (N_2772,N_2490,N_2473);
and U2773 (N_2773,N_2548,N_2537);
nor U2774 (N_2774,N_2435,N_2518);
xor U2775 (N_2775,N_2424,N_2541);
nand U2776 (N_2776,N_2475,N_2564);
and U2777 (N_2777,N_2410,N_2473);
nor U2778 (N_2778,N_2461,N_2510);
and U2779 (N_2779,N_2481,N_2441);
xor U2780 (N_2780,N_2586,N_2517);
nand U2781 (N_2781,N_2489,N_2420);
and U2782 (N_2782,N_2427,N_2526);
or U2783 (N_2783,N_2420,N_2429);
nor U2784 (N_2784,N_2480,N_2577);
and U2785 (N_2785,N_2515,N_2526);
or U2786 (N_2786,N_2500,N_2458);
xor U2787 (N_2787,N_2538,N_2441);
nand U2788 (N_2788,N_2466,N_2420);
or U2789 (N_2789,N_2571,N_2518);
and U2790 (N_2790,N_2448,N_2538);
xor U2791 (N_2791,N_2412,N_2471);
or U2792 (N_2792,N_2516,N_2481);
nor U2793 (N_2793,N_2460,N_2424);
or U2794 (N_2794,N_2407,N_2549);
xor U2795 (N_2795,N_2555,N_2550);
xnor U2796 (N_2796,N_2482,N_2480);
xnor U2797 (N_2797,N_2452,N_2539);
xnor U2798 (N_2798,N_2473,N_2576);
or U2799 (N_2799,N_2449,N_2501);
nor U2800 (N_2800,N_2698,N_2625);
or U2801 (N_2801,N_2778,N_2685);
nor U2802 (N_2802,N_2709,N_2741);
or U2803 (N_2803,N_2676,N_2603);
nand U2804 (N_2804,N_2660,N_2728);
xor U2805 (N_2805,N_2679,N_2792);
nor U2806 (N_2806,N_2730,N_2621);
nor U2807 (N_2807,N_2678,N_2705);
xnor U2808 (N_2808,N_2729,N_2703);
xor U2809 (N_2809,N_2769,N_2617);
or U2810 (N_2810,N_2734,N_2752);
nand U2811 (N_2811,N_2682,N_2736);
nor U2812 (N_2812,N_2650,N_2756);
nand U2813 (N_2813,N_2718,N_2794);
and U2814 (N_2814,N_2751,N_2661);
xor U2815 (N_2815,N_2616,N_2680);
nor U2816 (N_2816,N_2608,N_2717);
and U2817 (N_2817,N_2737,N_2768);
xor U2818 (N_2818,N_2649,N_2712);
or U2819 (N_2819,N_2619,N_2665);
nand U2820 (N_2820,N_2706,N_2771);
nor U2821 (N_2821,N_2600,N_2732);
xnor U2822 (N_2822,N_2711,N_2677);
nor U2823 (N_2823,N_2644,N_2633);
or U2824 (N_2824,N_2776,N_2782);
and U2825 (N_2825,N_2713,N_2797);
and U2826 (N_2826,N_2683,N_2690);
xor U2827 (N_2827,N_2610,N_2708);
and U2828 (N_2828,N_2646,N_2761);
xnor U2829 (N_2829,N_2758,N_2601);
or U2830 (N_2830,N_2618,N_2669);
or U2831 (N_2831,N_2742,N_2727);
xnor U2832 (N_2832,N_2673,N_2726);
nand U2833 (N_2833,N_2658,N_2607);
xnor U2834 (N_2834,N_2614,N_2749);
or U2835 (N_2835,N_2642,N_2605);
and U2836 (N_2836,N_2700,N_2606);
and U2837 (N_2837,N_2710,N_2755);
or U2838 (N_2838,N_2716,N_2604);
xnor U2839 (N_2839,N_2784,N_2641);
nand U2840 (N_2840,N_2788,N_2662);
and U2841 (N_2841,N_2671,N_2747);
nor U2842 (N_2842,N_2655,N_2627);
or U2843 (N_2843,N_2651,N_2656);
nor U2844 (N_2844,N_2659,N_2670);
and U2845 (N_2845,N_2681,N_2623);
nor U2846 (N_2846,N_2626,N_2615);
and U2847 (N_2847,N_2786,N_2643);
nor U2848 (N_2848,N_2745,N_2657);
nor U2849 (N_2849,N_2781,N_2789);
and U2850 (N_2850,N_2611,N_2757);
and U2851 (N_2851,N_2620,N_2739);
nand U2852 (N_2852,N_2720,N_2696);
nor U2853 (N_2853,N_2707,N_2686);
and U2854 (N_2854,N_2750,N_2687);
xnor U2855 (N_2855,N_2692,N_2780);
nor U2856 (N_2856,N_2631,N_2640);
xnor U2857 (N_2857,N_2715,N_2722);
or U2858 (N_2858,N_2672,N_2675);
and U2859 (N_2859,N_2721,N_2652);
nor U2860 (N_2860,N_2637,N_2763);
nand U2861 (N_2861,N_2663,N_2759);
nand U2862 (N_2862,N_2791,N_2684);
nor U2863 (N_2863,N_2785,N_2733);
and U2864 (N_2864,N_2629,N_2787);
xnor U2865 (N_2865,N_2754,N_2795);
nand U2866 (N_2866,N_2622,N_2770);
xnor U2867 (N_2867,N_2635,N_2779);
and U2868 (N_2868,N_2798,N_2743);
nand U2869 (N_2869,N_2777,N_2699);
nor U2870 (N_2870,N_2762,N_2725);
nand U2871 (N_2871,N_2697,N_2790);
or U2872 (N_2872,N_2793,N_2735);
nor U2873 (N_2873,N_2738,N_2764);
or U2874 (N_2874,N_2613,N_2731);
nand U2875 (N_2875,N_2602,N_2773);
nor U2876 (N_2876,N_2689,N_2695);
and U2877 (N_2877,N_2630,N_2799);
nor U2878 (N_2878,N_2639,N_2767);
nand U2879 (N_2879,N_2609,N_2654);
and U2880 (N_2880,N_2702,N_2667);
nand U2881 (N_2881,N_2666,N_2638);
and U2882 (N_2882,N_2647,N_2648);
and U2883 (N_2883,N_2704,N_2664);
xnor U2884 (N_2884,N_2693,N_2740);
and U2885 (N_2885,N_2634,N_2760);
xnor U2886 (N_2886,N_2694,N_2783);
nand U2887 (N_2887,N_2691,N_2753);
nor U2888 (N_2888,N_2748,N_2636);
nand U2889 (N_2889,N_2772,N_2774);
xnor U2890 (N_2890,N_2645,N_2714);
nor U2891 (N_2891,N_2724,N_2701);
xor U2892 (N_2892,N_2719,N_2688);
xor U2893 (N_2893,N_2775,N_2765);
nand U2894 (N_2894,N_2723,N_2628);
nor U2895 (N_2895,N_2624,N_2674);
or U2896 (N_2896,N_2766,N_2612);
and U2897 (N_2897,N_2653,N_2632);
and U2898 (N_2898,N_2668,N_2744);
or U2899 (N_2899,N_2746,N_2796);
xnor U2900 (N_2900,N_2658,N_2764);
nor U2901 (N_2901,N_2763,N_2601);
xor U2902 (N_2902,N_2751,N_2773);
nand U2903 (N_2903,N_2677,N_2750);
nor U2904 (N_2904,N_2644,N_2645);
xor U2905 (N_2905,N_2618,N_2656);
xor U2906 (N_2906,N_2602,N_2704);
nor U2907 (N_2907,N_2696,N_2735);
nor U2908 (N_2908,N_2724,N_2732);
and U2909 (N_2909,N_2615,N_2643);
nor U2910 (N_2910,N_2686,N_2668);
and U2911 (N_2911,N_2605,N_2623);
nor U2912 (N_2912,N_2627,N_2703);
or U2913 (N_2913,N_2762,N_2780);
nand U2914 (N_2914,N_2758,N_2783);
or U2915 (N_2915,N_2669,N_2765);
xor U2916 (N_2916,N_2750,N_2641);
nand U2917 (N_2917,N_2602,N_2650);
nand U2918 (N_2918,N_2612,N_2693);
nor U2919 (N_2919,N_2734,N_2652);
nand U2920 (N_2920,N_2757,N_2646);
and U2921 (N_2921,N_2707,N_2623);
or U2922 (N_2922,N_2601,N_2655);
xnor U2923 (N_2923,N_2630,N_2693);
nor U2924 (N_2924,N_2753,N_2741);
nor U2925 (N_2925,N_2634,N_2757);
and U2926 (N_2926,N_2723,N_2636);
or U2927 (N_2927,N_2657,N_2710);
nor U2928 (N_2928,N_2704,N_2605);
nand U2929 (N_2929,N_2778,N_2725);
nand U2930 (N_2930,N_2745,N_2649);
and U2931 (N_2931,N_2644,N_2677);
or U2932 (N_2932,N_2655,N_2670);
nor U2933 (N_2933,N_2643,N_2721);
or U2934 (N_2934,N_2643,N_2630);
nor U2935 (N_2935,N_2636,N_2611);
nor U2936 (N_2936,N_2650,N_2777);
xnor U2937 (N_2937,N_2713,N_2695);
nand U2938 (N_2938,N_2692,N_2609);
xor U2939 (N_2939,N_2749,N_2619);
or U2940 (N_2940,N_2643,N_2706);
nand U2941 (N_2941,N_2653,N_2731);
xnor U2942 (N_2942,N_2718,N_2648);
nor U2943 (N_2943,N_2788,N_2698);
and U2944 (N_2944,N_2615,N_2667);
and U2945 (N_2945,N_2798,N_2789);
nor U2946 (N_2946,N_2776,N_2617);
xor U2947 (N_2947,N_2657,N_2653);
and U2948 (N_2948,N_2731,N_2642);
nand U2949 (N_2949,N_2719,N_2779);
nor U2950 (N_2950,N_2654,N_2776);
or U2951 (N_2951,N_2651,N_2707);
nand U2952 (N_2952,N_2723,N_2724);
or U2953 (N_2953,N_2611,N_2643);
or U2954 (N_2954,N_2659,N_2772);
xnor U2955 (N_2955,N_2749,N_2764);
xor U2956 (N_2956,N_2762,N_2789);
xnor U2957 (N_2957,N_2654,N_2734);
or U2958 (N_2958,N_2769,N_2707);
xnor U2959 (N_2959,N_2789,N_2684);
nor U2960 (N_2960,N_2773,N_2758);
or U2961 (N_2961,N_2737,N_2700);
xnor U2962 (N_2962,N_2637,N_2625);
nor U2963 (N_2963,N_2711,N_2624);
and U2964 (N_2964,N_2796,N_2619);
and U2965 (N_2965,N_2707,N_2682);
nor U2966 (N_2966,N_2796,N_2651);
or U2967 (N_2967,N_2670,N_2741);
nand U2968 (N_2968,N_2795,N_2664);
or U2969 (N_2969,N_2703,N_2655);
and U2970 (N_2970,N_2711,N_2633);
xor U2971 (N_2971,N_2604,N_2664);
and U2972 (N_2972,N_2735,N_2794);
and U2973 (N_2973,N_2644,N_2675);
xor U2974 (N_2974,N_2710,N_2668);
nand U2975 (N_2975,N_2683,N_2636);
xor U2976 (N_2976,N_2601,N_2759);
and U2977 (N_2977,N_2740,N_2704);
nand U2978 (N_2978,N_2709,N_2635);
nand U2979 (N_2979,N_2756,N_2781);
xor U2980 (N_2980,N_2677,N_2770);
xor U2981 (N_2981,N_2617,N_2645);
and U2982 (N_2982,N_2641,N_2762);
nor U2983 (N_2983,N_2667,N_2663);
nor U2984 (N_2984,N_2723,N_2777);
nand U2985 (N_2985,N_2684,N_2623);
or U2986 (N_2986,N_2712,N_2728);
nor U2987 (N_2987,N_2652,N_2666);
or U2988 (N_2988,N_2691,N_2614);
nor U2989 (N_2989,N_2639,N_2707);
xor U2990 (N_2990,N_2614,N_2605);
and U2991 (N_2991,N_2679,N_2704);
xor U2992 (N_2992,N_2624,N_2602);
xor U2993 (N_2993,N_2614,N_2745);
xor U2994 (N_2994,N_2686,N_2750);
nand U2995 (N_2995,N_2691,N_2710);
xor U2996 (N_2996,N_2742,N_2654);
nor U2997 (N_2997,N_2791,N_2777);
xor U2998 (N_2998,N_2612,N_2718);
or U2999 (N_2999,N_2759,N_2679);
nor UO_0 (O_0,N_2816,N_2818);
and UO_1 (O_1,N_2843,N_2848);
nor UO_2 (O_2,N_2869,N_2917);
nor UO_3 (O_3,N_2859,N_2940);
and UO_4 (O_4,N_2860,N_2933);
or UO_5 (O_5,N_2811,N_2889);
nand UO_6 (O_6,N_2906,N_2960);
and UO_7 (O_7,N_2950,N_2946);
and UO_8 (O_8,N_2814,N_2943);
xor UO_9 (O_9,N_2885,N_2934);
and UO_10 (O_10,N_2912,N_2966);
nand UO_11 (O_11,N_2981,N_2810);
or UO_12 (O_12,N_2967,N_2945);
xnor UO_13 (O_13,N_2897,N_2931);
nand UO_14 (O_14,N_2991,N_2990);
xor UO_15 (O_15,N_2987,N_2831);
xnor UO_16 (O_16,N_2833,N_2850);
xor UO_17 (O_17,N_2999,N_2876);
or UO_18 (O_18,N_2823,N_2863);
and UO_19 (O_19,N_2985,N_2997);
and UO_20 (O_20,N_2805,N_2941);
xor UO_21 (O_21,N_2838,N_2832);
and UO_22 (O_22,N_2830,N_2845);
or UO_23 (O_23,N_2924,N_2898);
or UO_24 (O_24,N_2836,N_2888);
nor UO_25 (O_25,N_2929,N_2938);
nor UO_26 (O_26,N_2879,N_2948);
nor UO_27 (O_27,N_2854,N_2802);
nor UO_28 (O_28,N_2914,N_2902);
or UO_29 (O_29,N_2839,N_2891);
and UO_30 (O_30,N_2865,N_2826);
xor UO_31 (O_31,N_2951,N_2974);
and UO_32 (O_32,N_2834,N_2947);
nor UO_33 (O_33,N_2872,N_2837);
xor UO_34 (O_34,N_2904,N_2909);
xor UO_35 (O_35,N_2827,N_2886);
and UO_36 (O_36,N_2870,N_2989);
nor UO_37 (O_37,N_2862,N_2982);
xor UO_38 (O_38,N_2952,N_2942);
and UO_39 (O_39,N_2846,N_2925);
nand UO_40 (O_40,N_2923,N_2883);
and UO_41 (O_41,N_2986,N_2922);
nor UO_42 (O_42,N_2857,N_2841);
nand UO_43 (O_43,N_2901,N_2988);
and UO_44 (O_44,N_2820,N_2899);
or UO_45 (O_45,N_2961,N_2969);
nand UO_46 (O_46,N_2822,N_2955);
or UO_47 (O_47,N_2962,N_2896);
and UO_48 (O_48,N_2949,N_2927);
or UO_49 (O_49,N_2829,N_2873);
xnor UO_50 (O_50,N_2964,N_2882);
xnor UO_51 (O_51,N_2919,N_2858);
nand UO_52 (O_52,N_2847,N_2852);
and UO_53 (O_53,N_2932,N_2861);
xnor UO_54 (O_54,N_2894,N_2815);
nor UO_55 (O_55,N_2812,N_2842);
xor UO_56 (O_56,N_2871,N_2813);
nor UO_57 (O_57,N_2995,N_2851);
and UO_58 (O_58,N_2980,N_2939);
xor UO_59 (O_59,N_2890,N_2868);
nand UO_60 (O_60,N_2910,N_2992);
xnor UO_61 (O_61,N_2973,N_2887);
and UO_62 (O_62,N_2903,N_2803);
nor UO_63 (O_63,N_2908,N_2840);
or UO_64 (O_64,N_2957,N_2998);
or UO_65 (O_65,N_2920,N_2975);
and UO_66 (O_66,N_2996,N_2972);
nor UO_67 (O_67,N_2911,N_2935);
nor UO_68 (O_68,N_2963,N_2970);
nor UO_69 (O_69,N_2855,N_2937);
or UO_70 (O_70,N_2884,N_2892);
nand UO_71 (O_71,N_2874,N_2956);
nor UO_72 (O_72,N_2953,N_2828);
or UO_73 (O_73,N_2926,N_2844);
or UO_74 (O_74,N_2856,N_2976);
nand UO_75 (O_75,N_2809,N_2893);
nand UO_76 (O_76,N_2979,N_2959);
nand UO_77 (O_77,N_2907,N_2867);
nor UO_78 (O_78,N_2881,N_2954);
and UO_79 (O_79,N_2877,N_2808);
nor UO_80 (O_80,N_2994,N_2978);
nor UO_81 (O_81,N_2807,N_2968);
or UO_82 (O_82,N_2977,N_2993);
xnor UO_83 (O_83,N_2821,N_2824);
or UO_84 (O_84,N_2817,N_2971);
or UO_85 (O_85,N_2866,N_2918);
or UO_86 (O_86,N_2895,N_2905);
xor UO_87 (O_87,N_2864,N_2984);
and UO_88 (O_88,N_2958,N_2916);
nand UO_89 (O_89,N_2944,N_2800);
nor UO_90 (O_90,N_2965,N_2936);
nand UO_91 (O_91,N_2801,N_2825);
nand UO_92 (O_92,N_2849,N_2930);
xnor UO_93 (O_93,N_2913,N_2928);
nor UO_94 (O_94,N_2921,N_2853);
xor UO_95 (O_95,N_2835,N_2878);
nor UO_96 (O_96,N_2804,N_2983);
nand UO_97 (O_97,N_2915,N_2900);
and UO_98 (O_98,N_2819,N_2806);
or UO_99 (O_99,N_2880,N_2875);
nor UO_100 (O_100,N_2875,N_2838);
xnor UO_101 (O_101,N_2827,N_2901);
and UO_102 (O_102,N_2918,N_2941);
and UO_103 (O_103,N_2921,N_2819);
and UO_104 (O_104,N_2847,N_2992);
or UO_105 (O_105,N_2973,N_2909);
or UO_106 (O_106,N_2843,N_2884);
or UO_107 (O_107,N_2995,N_2947);
xor UO_108 (O_108,N_2865,N_2901);
nand UO_109 (O_109,N_2817,N_2827);
xor UO_110 (O_110,N_2809,N_2819);
nor UO_111 (O_111,N_2843,N_2999);
nand UO_112 (O_112,N_2928,N_2885);
xor UO_113 (O_113,N_2837,N_2807);
nor UO_114 (O_114,N_2980,N_2894);
and UO_115 (O_115,N_2981,N_2997);
xnor UO_116 (O_116,N_2832,N_2907);
nand UO_117 (O_117,N_2831,N_2979);
or UO_118 (O_118,N_2956,N_2848);
nand UO_119 (O_119,N_2885,N_2823);
xor UO_120 (O_120,N_2898,N_2862);
nand UO_121 (O_121,N_2941,N_2946);
xor UO_122 (O_122,N_2866,N_2909);
and UO_123 (O_123,N_2944,N_2927);
xor UO_124 (O_124,N_2872,N_2814);
and UO_125 (O_125,N_2887,N_2922);
and UO_126 (O_126,N_2801,N_2892);
and UO_127 (O_127,N_2982,N_2872);
nor UO_128 (O_128,N_2998,N_2894);
and UO_129 (O_129,N_2833,N_2872);
xnor UO_130 (O_130,N_2808,N_2949);
xor UO_131 (O_131,N_2902,N_2845);
xnor UO_132 (O_132,N_2947,N_2806);
and UO_133 (O_133,N_2958,N_2970);
and UO_134 (O_134,N_2975,N_2845);
xnor UO_135 (O_135,N_2870,N_2968);
nor UO_136 (O_136,N_2806,N_2833);
nor UO_137 (O_137,N_2910,N_2956);
or UO_138 (O_138,N_2884,N_2832);
nor UO_139 (O_139,N_2928,N_2901);
xor UO_140 (O_140,N_2987,N_2995);
or UO_141 (O_141,N_2916,N_2856);
nand UO_142 (O_142,N_2957,N_2850);
nor UO_143 (O_143,N_2895,N_2870);
and UO_144 (O_144,N_2888,N_2868);
nor UO_145 (O_145,N_2940,N_2908);
and UO_146 (O_146,N_2968,N_2943);
or UO_147 (O_147,N_2818,N_2988);
nor UO_148 (O_148,N_2817,N_2899);
nand UO_149 (O_149,N_2863,N_2834);
xnor UO_150 (O_150,N_2900,N_2970);
and UO_151 (O_151,N_2802,N_2962);
xor UO_152 (O_152,N_2907,N_2865);
nor UO_153 (O_153,N_2828,N_2900);
nand UO_154 (O_154,N_2826,N_2816);
and UO_155 (O_155,N_2961,N_2835);
nand UO_156 (O_156,N_2801,N_2879);
or UO_157 (O_157,N_2938,N_2817);
nor UO_158 (O_158,N_2921,N_2968);
and UO_159 (O_159,N_2977,N_2878);
or UO_160 (O_160,N_2880,N_2888);
or UO_161 (O_161,N_2843,N_2979);
or UO_162 (O_162,N_2975,N_2945);
and UO_163 (O_163,N_2813,N_2821);
and UO_164 (O_164,N_2976,N_2878);
or UO_165 (O_165,N_2816,N_2963);
xnor UO_166 (O_166,N_2920,N_2991);
or UO_167 (O_167,N_2846,N_2926);
nor UO_168 (O_168,N_2929,N_2924);
xor UO_169 (O_169,N_2847,N_2838);
nand UO_170 (O_170,N_2979,N_2895);
and UO_171 (O_171,N_2849,N_2963);
nand UO_172 (O_172,N_2959,N_2985);
xnor UO_173 (O_173,N_2901,N_2938);
and UO_174 (O_174,N_2975,N_2824);
nor UO_175 (O_175,N_2982,N_2932);
and UO_176 (O_176,N_2942,N_2917);
nand UO_177 (O_177,N_2997,N_2983);
xnor UO_178 (O_178,N_2978,N_2856);
or UO_179 (O_179,N_2861,N_2805);
xor UO_180 (O_180,N_2905,N_2911);
xnor UO_181 (O_181,N_2941,N_2961);
and UO_182 (O_182,N_2884,N_2805);
nor UO_183 (O_183,N_2955,N_2953);
and UO_184 (O_184,N_2808,N_2831);
or UO_185 (O_185,N_2818,N_2862);
nand UO_186 (O_186,N_2888,N_2957);
xnor UO_187 (O_187,N_2845,N_2843);
or UO_188 (O_188,N_2846,N_2809);
or UO_189 (O_189,N_2934,N_2826);
nand UO_190 (O_190,N_2874,N_2811);
xnor UO_191 (O_191,N_2936,N_2898);
nor UO_192 (O_192,N_2954,N_2804);
or UO_193 (O_193,N_2832,N_2866);
nand UO_194 (O_194,N_2959,N_2902);
and UO_195 (O_195,N_2982,N_2810);
nand UO_196 (O_196,N_2978,N_2936);
xor UO_197 (O_197,N_2869,N_2894);
nor UO_198 (O_198,N_2934,N_2902);
xnor UO_199 (O_199,N_2891,N_2878);
and UO_200 (O_200,N_2987,N_2822);
or UO_201 (O_201,N_2846,N_2828);
nand UO_202 (O_202,N_2815,N_2853);
and UO_203 (O_203,N_2908,N_2922);
nand UO_204 (O_204,N_2888,N_2807);
xor UO_205 (O_205,N_2931,N_2886);
nor UO_206 (O_206,N_2877,N_2983);
and UO_207 (O_207,N_2914,N_2805);
nand UO_208 (O_208,N_2995,N_2953);
or UO_209 (O_209,N_2822,N_2997);
xnor UO_210 (O_210,N_2850,N_2867);
xnor UO_211 (O_211,N_2988,N_2864);
and UO_212 (O_212,N_2888,N_2850);
xnor UO_213 (O_213,N_2872,N_2978);
and UO_214 (O_214,N_2900,N_2918);
and UO_215 (O_215,N_2959,N_2940);
nor UO_216 (O_216,N_2939,N_2844);
nand UO_217 (O_217,N_2831,N_2982);
nand UO_218 (O_218,N_2934,N_2819);
xnor UO_219 (O_219,N_2938,N_2809);
xor UO_220 (O_220,N_2992,N_2887);
nand UO_221 (O_221,N_2804,N_2992);
and UO_222 (O_222,N_2971,N_2954);
and UO_223 (O_223,N_2979,N_2837);
or UO_224 (O_224,N_2939,N_2841);
nand UO_225 (O_225,N_2975,N_2815);
and UO_226 (O_226,N_2972,N_2891);
nor UO_227 (O_227,N_2829,N_2848);
and UO_228 (O_228,N_2866,N_2898);
and UO_229 (O_229,N_2920,N_2978);
nor UO_230 (O_230,N_2971,N_2855);
and UO_231 (O_231,N_2882,N_2980);
nand UO_232 (O_232,N_2859,N_2953);
nor UO_233 (O_233,N_2861,N_2841);
nor UO_234 (O_234,N_2817,N_2948);
nand UO_235 (O_235,N_2916,N_2802);
xnor UO_236 (O_236,N_2994,N_2930);
nand UO_237 (O_237,N_2833,N_2925);
nand UO_238 (O_238,N_2979,N_2860);
nand UO_239 (O_239,N_2907,N_2993);
nand UO_240 (O_240,N_2865,N_2988);
and UO_241 (O_241,N_2901,N_2891);
and UO_242 (O_242,N_2961,N_2816);
nor UO_243 (O_243,N_2910,N_2961);
nor UO_244 (O_244,N_2890,N_2938);
nor UO_245 (O_245,N_2843,N_2874);
nor UO_246 (O_246,N_2877,N_2902);
xnor UO_247 (O_247,N_2948,N_2923);
nand UO_248 (O_248,N_2827,N_2954);
and UO_249 (O_249,N_2897,N_2993);
xor UO_250 (O_250,N_2945,N_2884);
nor UO_251 (O_251,N_2810,N_2876);
xnor UO_252 (O_252,N_2937,N_2957);
nor UO_253 (O_253,N_2961,N_2836);
nand UO_254 (O_254,N_2854,N_2857);
nand UO_255 (O_255,N_2873,N_2954);
or UO_256 (O_256,N_2889,N_2925);
nand UO_257 (O_257,N_2911,N_2831);
or UO_258 (O_258,N_2899,N_2915);
or UO_259 (O_259,N_2868,N_2833);
nand UO_260 (O_260,N_2894,N_2872);
nand UO_261 (O_261,N_2882,N_2892);
and UO_262 (O_262,N_2892,N_2874);
and UO_263 (O_263,N_2993,N_2991);
xnor UO_264 (O_264,N_2844,N_2813);
and UO_265 (O_265,N_2907,N_2961);
or UO_266 (O_266,N_2945,N_2921);
nor UO_267 (O_267,N_2959,N_2870);
nor UO_268 (O_268,N_2901,N_2833);
nand UO_269 (O_269,N_2804,N_2987);
nand UO_270 (O_270,N_2878,N_2935);
and UO_271 (O_271,N_2952,N_2801);
xor UO_272 (O_272,N_2929,N_2999);
or UO_273 (O_273,N_2967,N_2892);
or UO_274 (O_274,N_2909,N_2919);
and UO_275 (O_275,N_2839,N_2824);
nor UO_276 (O_276,N_2894,N_2907);
and UO_277 (O_277,N_2807,N_2884);
xor UO_278 (O_278,N_2870,N_2954);
or UO_279 (O_279,N_2927,N_2914);
nand UO_280 (O_280,N_2969,N_2945);
nand UO_281 (O_281,N_2983,N_2875);
nand UO_282 (O_282,N_2924,N_2835);
or UO_283 (O_283,N_2806,N_2807);
nand UO_284 (O_284,N_2826,N_2840);
and UO_285 (O_285,N_2823,N_2806);
nand UO_286 (O_286,N_2823,N_2828);
xnor UO_287 (O_287,N_2820,N_2942);
nor UO_288 (O_288,N_2872,N_2831);
and UO_289 (O_289,N_2899,N_2810);
xor UO_290 (O_290,N_2851,N_2891);
nor UO_291 (O_291,N_2948,N_2910);
nor UO_292 (O_292,N_2852,N_2884);
xor UO_293 (O_293,N_2821,N_2923);
or UO_294 (O_294,N_2955,N_2851);
nor UO_295 (O_295,N_2889,N_2977);
or UO_296 (O_296,N_2976,N_2864);
xnor UO_297 (O_297,N_2878,N_2865);
nor UO_298 (O_298,N_2805,N_2923);
and UO_299 (O_299,N_2986,N_2817);
and UO_300 (O_300,N_2993,N_2860);
nor UO_301 (O_301,N_2944,N_2804);
nor UO_302 (O_302,N_2838,N_2883);
nand UO_303 (O_303,N_2839,N_2908);
or UO_304 (O_304,N_2852,N_2812);
xor UO_305 (O_305,N_2822,N_2893);
and UO_306 (O_306,N_2865,N_2816);
and UO_307 (O_307,N_2972,N_2945);
xor UO_308 (O_308,N_2931,N_2800);
nand UO_309 (O_309,N_2867,N_2956);
and UO_310 (O_310,N_2835,N_2985);
or UO_311 (O_311,N_2839,N_2995);
or UO_312 (O_312,N_2981,N_2826);
nor UO_313 (O_313,N_2986,N_2987);
xor UO_314 (O_314,N_2981,N_2909);
nor UO_315 (O_315,N_2903,N_2800);
or UO_316 (O_316,N_2917,N_2979);
nand UO_317 (O_317,N_2852,N_2909);
nand UO_318 (O_318,N_2800,N_2909);
or UO_319 (O_319,N_2961,N_2916);
nor UO_320 (O_320,N_2816,N_2947);
nor UO_321 (O_321,N_2982,N_2850);
xnor UO_322 (O_322,N_2939,N_2902);
nor UO_323 (O_323,N_2980,N_2996);
and UO_324 (O_324,N_2857,N_2950);
or UO_325 (O_325,N_2801,N_2857);
xnor UO_326 (O_326,N_2918,N_2981);
xnor UO_327 (O_327,N_2969,N_2892);
nor UO_328 (O_328,N_2957,N_2893);
nand UO_329 (O_329,N_2926,N_2856);
nor UO_330 (O_330,N_2967,N_2815);
nand UO_331 (O_331,N_2921,N_2809);
xnor UO_332 (O_332,N_2864,N_2987);
nor UO_333 (O_333,N_2975,N_2904);
and UO_334 (O_334,N_2948,N_2874);
nand UO_335 (O_335,N_2902,N_2883);
or UO_336 (O_336,N_2828,N_2925);
xnor UO_337 (O_337,N_2822,N_2973);
xnor UO_338 (O_338,N_2827,N_2953);
nor UO_339 (O_339,N_2885,N_2883);
or UO_340 (O_340,N_2913,N_2801);
or UO_341 (O_341,N_2969,N_2902);
nor UO_342 (O_342,N_2850,N_2981);
nand UO_343 (O_343,N_2885,N_2952);
nor UO_344 (O_344,N_2907,N_2887);
nand UO_345 (O_345,N_2966,N_2837);
xnor UO_346 (O_346,N_2818,N_2982);
or UO_347 (O_347,N_2933,N_2941);
nor UO_348 (O_348,N_2842,N_2966);
nor UO_349 (O_349,N_2896,N_2928);
and UO_350 (O_350,N_2819,N_2945);
nor UO_351 (O_351,N_2827,N_2855);
or UO_352 (O_352,N_2857,N_2907);
xor UO_353 (O_353,N_2874,N_2974);
nand UO_354 (O_354,N_2847,N_2829);
or UO_355 (O_355,N_2815,N_2954);
nor UO_356 (O_356,N_2992,N_2867);
nor UO_357 (O_357,N_2919,N_2914);
and UO_358 (O_358,N_2966,N_2955);
or UO_359 (O_359,N_2881,N_2864);
nand UO_360 (O_360,N_2928,N_2868);
xnor UO_361 (O_361,N_2838,N_2981);
xnor UO_362 (O_362,N_2957,N_2837);
or UO_363 (O_363,N_2924,N_2848);
nand UO_364 (O_364,N_2853,N_2903);
and UO_365 (O_365,N_2891,N_2874);
xor UO_366 (O_366,N_2822,N_2948);
nor UO_367 (O_367,N_2880,N_2892);
or UO_368 (O_368,N_2953,N_2826);
nor UO_369 (O_369,N_2804,N_2940);
and UO_370 (O_370,N_2826,N_2887);
nand UO_371 (O_371,N_2983,N_2925);
or UO_372 (O_372,N_2941,N_2996);
nand UO_373 (O_373,N_2904,N_2858);
or UO_374 (O_374,N_2919,N_2978);
or UO_375 (O_375,N_2954,N_2983);
xnor UO_376 (O_376,N_2956,N_2803);
nor UO_377 (O_377,N_2841,N_2945);
and UO_378 (O_378,N_2908,N_2918);
and UO_379 (O_379,N_2844,N_2856);
or UO_380 (O_380,N_2848,N_2839);
nor UO_381 (O_381,N_2916,N_2937);
nand UO_382 (O_382,N_2962,N_2983);
and UO_383 (O_383,N_2824,N_2953);
or UO_384 (O_384,N_2839,N_2811);
xor UO_385 (O_385,N_2985,N_2823);
or UO_386 (O_386,N_2896,N_2930);
nand UO_387 (O_387,N_2998,N_2880);
or UO_388 (O_388,N_2848,N_2913);
and UO_389 (O_389,N_2907,N_2874);
nor UO_390 (O_390,N_2973,N_2975);
nand UO_391 (O_391,N_2982,N_2863);
nand UO_392 (O_392,N_2982,N_2909);
nor UO_393 (O_393,N_2831,N_2960);
or UO_394 (O_394,N_2845,N_2835);
and UO_395 (O_395,N_2857,N_2800);
or UO_396 (O_396,N_2946,N_2981);
nor UO_397 (O_397,N_2861,N_2948);
xnor UO_398 (O_398,N_2931,N_2979);
or UO_399 (O_399,N_2850,N_2880);
or UO_400 (O_400,N_2944,N_2972);
and UO_401 (O_401,N_2963,N_2815);
nand UO_402 (O_402,N_2877,N_2951);
nor UO_403 (O_403,N_2855,N_2804);
or UO_404 (O_404,N_2999,N_2837);
and UO_405 (O_405,N_2946,N_2872);
or UO_406 (O_406,N_2930,N_2972);
xnor UO_407 (O_407,N_2854,N_2937);
xnor UO_408 (O_408,N_2816,N_2860);
or UO_409 (O_409,N_2822,N_2832);
xnor UO_410 (O_410,N_2972,N_2880);
nor UO_411 (O_411,N_2892,N_2943);
and UO_412 (O_412,N_2838,N_2916);
nor UO_413 (O_413,N_2973,N_2821);
and UO_414 (O_414,N_2973,N_2985);
and UO_415 (O_415,N_2883,N_2987);
nor UO_416 (O_416,N_2963,N_2931);
or UO_417 (O_417,N_2903,N_2966);
or UO_418 (O_418,N_2924,N_2992);
and UO_419 (O_419,N_2915,N_2946);
and UO_420 (O_420,N_2907,N_2856);
nand UO_421 (O_421,N_2979,N_2923);
nor UO_422 (O_422,N_2909,N_2849);
or UO_423 (O_423,N_2975,N_2928);
or UO_424 (O_424,N_2958,N_2883);
or UO_425 (O_425,N_2882,N_2814);
nor UO_426 (O_426,N_2887,N_2807);
nor UO_427 (O_427,N_2905,N_2801);
xnor UO_428 (O_428,N_2800,N_2956);
nor UO_429 (O_429,N_2947,N_2960);
and UO_430 (O_430,N_2997,N_2956);
and UO_431 (O_431,N_2923,N_2888);
nor UO_432 (O_432,N_2886,N_2803);
xor UO_433 (O_433,N_2955,N_2862);
xnor UO_434 (O_434,N_2864,N_2892);
xnor UO_435 (O_435,N_2952,N_2951);
nor UO_436 (O_436,N_2839,N_2948);
and UO_437 (O_437,N_2956,N_2842);
nand UO_438 (O_438,N_2972,N_2877);
or UO_439 (O_439,N_2861,N_2828);
nand UO_440 (O_440,N_2955,N_2920);
nor UO_441 (O_441,N_2876,N_2838);
and UO_442 (O_442,N_2812,N_2902);
xor UO_443 (O_443,N_2901,N_2850);
nor UO_444 (O_444,N_2837,N_2959);
nand UO_445 (O_445,N_2833,N_2845);
and UO_446 (O_446,N_2846,N_2903);
nand UO_447 (O_447,N_2917,N_2834);
nor UO_448 (O_448,N_2854,N_2942);
nor UO_449 (O_449,N_2841,N_2984);
and UO_450 (O_450,N_2987,N_2921);
nand UO_451 (O_451,N_2972,N_2804);
or UO_452 (O_452,N_2810,N_2875);
nand UO_453 (O_453,N_2883,N_2938);
and UO_454 (O_454,N_2825,N_2890);
and UO_455 (O_455,N_2976,N_2845);
and UO_456 (O_456,N_2950,N_2904);
or UO_457 (O_457,N_2815,N_2817);
or UO_458 (O_458,N_2890,N_2810);
or UO_459 (O_459,N_2955,N_2988);
and UO_460 (O_460,N_2960,N_2987);
xor UO_461 (O_461,N_2921,N_2893);
nand UO_462 (O_462,N_2953,N_2976);
nor UO_463 (O_463,N_2930,N_2940);
or UO_464 (O_464,N_2964,N_2836);
xnor UO_465 (O_465,N_2927,N_2877);
nand UO_466 (O_466,N_2979,N_2972);
nand UO_467 (O_467,N_2863,N_2827);
nand UO_468 (O_468,N_2821,N_2979);
nor UO_469 (O_469,N_2840,N_2877);
xnor UO_470 (O_470,N_2966,N_2849);
and UO_471 (O_471,N_2963,N_2987);
and UO_472 (O_472,N_2872,N_2898);
or UO_473 (O_473,N_2916,N_2927);
and UO_474 (O_474,N_2968,N_2812);
xnor UO_475 (O_475,N_2970,N_2949);
nand UO_476 (O_476,N_2899,N_2945);
nor UO_477 (O_477,N_2913,N_2897);
nor UO_478 (O_478,N_2938,N_2930);
nand UO_479 (O_479,N_2958,N_2821);
nor UO_480 (O_480,N_2816,N_2936);
and UO_481 (O_481,N_2804,N_2977);
or UO_482 (O_482,N_2899,N_2866);
or UO_483 (O_483,N_2807,N_2843);
xnor UO_484 (O_484,N_2998,N_2814);
nand UO_485 (O_485,N_2966,N_2902);
and UO_486 (O_486,N_2942,N_2880);
xor UO_487 (O_487,N_2842,N_2938);
and UO_488 (O_488,N_2940,N_2905);
nand UO_489 (O_489,N_2864,N_2934);
nor UO_490 (O_490,N_2802,N_2922);
nor UO_491 (O_491,N_2863,N_2824);
or UO_492 (O_492,N_2848,N_2827);
xnor UO_493 (O_493,N_2849,N_2921);
xor UO_494 (O_494,N_2805,N_2866);
or UO_495 (O_495,N_2964,N_2838);
nand UO_496 (O_496,N_2876,N_2912);
xnor UO_497 (O_497,N_2937,N_2952);
nor UO_498 (O_498,N_2879,N_2935);
and UO_499 (O_499,N_2825,N_2829);
endmodule