module basic_750_5000_1000_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_572,In_428);
xnor U1 (N_1,In_425,In_203);
and U2 (N_2,In_448,In_537);
or U3 (N_3,In_71,In_671);
xor U4 (N_4,In_343,In_417);
xnor U5 (N_5,In_541,In_69);
and U6 (N_6,In_597,In_515);
and U7 (N_7,In_124,In_204);
nand U8 (N_8,In_227,In_30);
or U9 (N_9,In_578,In_216);
and U10 (N_10,In_443,In_586);
nor U11 (N_11,In_238,In_290);
xnor U12 (N_12,In_126,In_280);
xor U13 (N_13,In_478,In_392);
nor U14 (N_14,In_451,In_195);
or U15 (N_15,In_221,In_624);
or U16 (N_16,In_147,In_271);
nand U17 (N_17,In_42,In_437);
and U18 (N_18,In_207,In_731);
nand U19 (N_19,In_288,In_678);
xor U20 (N_20,In_401,In_329);
nand U21 (N_21,In_130,In_587);
xnor U22 (N_22,In_63,In_67);
and U23 (N_23,In_418,In_676);
nor U24 (N_24,In_60,In_420);
or U25 (N_25,In_562,In_354);
xnor U26 (N_26,In_146,In_361);
nand U27 (N_27,In_426,In_727);
xnor U28 (N_28,In_114,In_157);
and U29 (N_29,In_315,In_513);
nor U30 (N_30,In_364,In_480);
nor U31 (N_31,In_331,In_270);
nor U32 (N_32,In_400,In_273);
nor U33 (N_33,In_10,In_345);
and U34 (N_34,In_222,In_319);
xor U35 (N_35,In_390,In_557);
xnor U36 (N_36,In_320,In_46);
and U37 (N_37,In_610,In_163);
or U38 (N_38,In_430,In_25);
and U39 (N_39,In_29,In_566);
nand U40 (N_40,In_675,In_249);
and U41 (N_41,In_258,In_447);
xnor U42 (N_42,In_623,In_733);
or U43 (N_43,In_110,In_301);
or U44 (N_44,In_24,In_252);
and U45 (N_45,In_398,In_213);
xor U46 (N_46,In_720,In_441);
nor U47 (N_47,In_17,In_602);
nand U48 (N_48,In_19,In_322);
nor U49 (N_49,In_326,In_618);
nor U50 (N_50,In_520,In_479);
nand U51 (N_51,In_214,In_483);
or U52 (N_52,In_427,In_306);
xor U53 (N_53,In_487,In_554);
nor U54 (N_54,In_715,In_149);
or U55 (N_55,In_607,In_158);
nor U56 (N_56,In_89,In_583);
and U57 (N_57,In_416,In_95);
nand U58 (N_58,In_482,In_540);
nand U59 (N_59,In_576,In_160);
nor U60 (N_60,In_517,In_674);
and U61 (N_61,In_497,In_358);
and U62 (N_62,In_429,In_709);
and U63 (N_63,In_355,In_710);
or U64 (N_64,In_645,In_380);
nand U65 (N_65,In_615,In_558);
or U66 (N_66,In_542,In_712);
or U67 (N_67,In_632,In_634);
xnor U68 (N_68,In_27,In_510);
or U69 (N_69,In_279,In_545);
nor U70 (N_70,In_12,In_412);
xnor U71 (N_71,In_198,In_184);
or U72 (N_72,In_611,In_434);
nor U73 (N_73,In_38,In_350);
nand U74 (N_74,In_155,In_525);
xnor U75 (N_75,In_100,In_643);
nor U76 (N_76,In_310,In_594);
or U77 (N_77,In_599,In_263);
or U78 (N_78,In_706,In_440);
xor U79 (N_79,In_685,In_14);
and U80 (N_80,In_405,In_508);
xor U81 (N_81,In_116,In_352);
and U82 (N_82,In_551,In_743);
or U83 (N_83,In_395,In_43);
and U84 (N_84,In_229,In_389);
nor U85 (N_85,In_255,In_553);
and U86 (N_86,In_664,In_749);
nand U87 (N_87,In_708,In_650);
and U88 (N_88,In_208,In_555);
nand U89 (N_89,In_449,In_682);
nand U90 (N_90,In_248,In_103);
xor U91 (N_91,In_563,In_236);
nor U92 (N_92,In_346,In_212);
nand U93 (N_93,In_704,In_128);
or U94 (N_94,In_588,In_86);
xnor U95 (N_95,In_174,In_18);
nor U96 (N_96,In_596,In_409);
xnor U97 (N_97,In_591,In_64);
nand U98 (N_98,In_717,In_382);
nand U99 (N_99,In_393,In_442);
xnor U100 (N_100,In_61,In_237);
nand U101 (N_101,In_431,In_359);
nor U102 (N_102,In_692,In_215);
and U103 (N_103,In_565,In_538);
xor U104 (N_104,In_651,In_250);
nand U105 (N_105,In_580,In_220);
nand U106 (N_106,In_22,In_402);
nor U107 (N_107,In_115,In_690);
xnor U108 (N_108,In_104,In_622);
nand U109 (N_109,In_458,In_694);
nor U110 (N_110,In_106,In_432);
xor U111 (N_111,In_687,In_461);
or U112 (N_112,In_88,In_261);
nand U113 (N_113,In_272,In_492);
or U114 (N_114,In_330,In_721);
nand U115 (N_115,In_728,In_481);
nor U116 (N_116,In_544,In_183);
xor U117 (N_117,In_136,In_714);
nor U118 (N_118,In_631,In_683);
nor U119 (N_119,In_150,In_85);
xnor U120 (N_120,In_57,In_524);
nand U121 (N_121,In_499,In_502);
or U122 (N_122,In_351,In_713);
and U123 (N_123,In_747,In_152);
xnor U124 (N_124,In_112,In_16);
or U125 (N_125,In_96,In_72);
and U126 (N_126,In_403,In_275);
xnor U127 (N_127,In_323,In_700);
xnor U128 (N_128,In_247,In_699);
nand U129 (N_129,In_87,In_530);
xnor U130 (N_130,In_298,In_48);
xor U131 (N_131,In_410,In_388);
or U132 (N_132,In_450,In_598);
or U133 (N_133,In_91,In_219);
and U134 (N_134,In_180,In_534);
or U135 (N_135,In_295,In_745);
xor U136 (N_136,In_696,In_469);
xnor U137 (N_137,In_304,In_44);
or U138 (N_138,In_669,In_338);
and U139 (N_139,In_28,In_702);
nand U140 (N_140,In_670,In_209);
nor U141 (N_141,In_285,In_202);
xor U142 (N_142,In_74,In_582);
nor U143 (N_143,In_101,In_4);
nor U144 (N_144,In_467,In_665);
nand U145 (N_145,In_569,In_471);
nand U146 (N_146,In_653,In_80);
or U147 (N_147,In_404,In_484);
nor U148 (N_148,In_567,In_577);
or U149 (N_149,In_59,In_318);
and U150 (N_150,In_644,In_140);
and U151 (N_151,In_648,In_438);
and U152 (N_152,In_627,In_739);
xnor U153 (N_153,In_83,In_287);
nor U154 (N_154,In_600,In_34);
nor U155 (N_155,In_433,In_111);
nor U156 (N_156,In_79,In_585);
nor U157 (N_157,In_139,In_374);
nand U158 (N_158,In_546,In_603);
and U159 (N_159,In_415,In_617);
and U160 (N_160,In_168,In_496);
nor U161 (N_161,In_197,In_143);
and U162 (N_162,In_133,In_532);
nor U163 (N_163,In_439,In_668);
nor U164 (N_164,In_408,In_62);
nor U165 (N_165,In_454,In_284);
nand U166 (N_166,In_93,In_226);
and U167 (N_167,In_719,In_381);
and U168 (N_168,In_21,In_657);
xnor U169 (N_169,In_200,In_453);
nand U170 (N_170,In_205,In_550);
and U171 (N_171,In_192,In_309);
nand U172 (N_172,In_135,In_641);
nor U173 (N_173,In_182,In_424);
nand U174 (N_174,In_47,In_729);
and U175 (N_175,In_9,In_573);
and U176 (N_176,In_262,In_691);
and U177 (N_177,In_0,In_512);
or U178 (N_178,In_385,In_194);
or U179 (N_179,In_356,In_52);
xor U180 (N_180,In_742,In_341);
nand U181 (N_181,In_638,In_593);
or U182 (N_182,In_604,In_397);
xor U183 (N_183,In_501,In_628);
nor U184 (N_184,In_463,In_196);
nor U185 (N_185,In_373,In_734);
and U186 (N_186,In_23,In_37);
nor U187 (N_187,In_489,In_276);
nand U188 (N_188,In_514,In_148);
or U189 (N_189,In_107,In_7);
or U190 (N_190,In_39,In_460);
nor U191 (N_191,In_187,In_575);
nand U192 (N_192,In_190,In_137);
xor U193 (N_193,In_490,In_84);
or U194 (N_194,In_521,In_141);
xor U195 (N_195,In_286,In_457);
or U196 (N_196,In_58,In_477);
nand U197 (N_197,In_156,In_169);
nor U198 (N_198,In_711,In_475);
nand U199 (N_199,In_268,In_109);
nand U200 (N_200,In_120,In_97);
xor U201 (N_201,In_297,In_741);
xnor U202 (N_202,In_680,In_703);
nand U203 (N_203,In_144,In_661);
xnor U204 (N_204,In_244,In_166);
nand U205 (N_205,In_102,In_142);
and U206 (N_206,In_667,In_383);
nand U207 (N_207,In_239,In_462);
nand U208 (N_208,In_649,In_289);
xnor U209 (N_209,In_199,In_518);
and U210 (N_210,In_179,In_172);
and U211 (N_211,In_105,In_716);
nor U212 (N_212,In_185,In_231);
and U213 (N_213,In_53,In_488);
xor U214 (N_214,In_684,In_344);
or U215 (N_215,In_317,In_459);
nor U216 (N_216,In_595,In_436);
nand U217 (N_217,In_73,In_642);
xnor U218 (N_218,In_363,In_165);
xor U219 (N_219,In_178,In_151);
and U220 (N_220,In_293,In_125);
or U221 (N_221,In_737,In_570);
nor U222 (N_222,In_294,In_673);
nand U223 (N_223,In_693,In_311);
nand U224 (N_224,In_689,In_500);
or U225 (N_225,In_305,In_206);
xor U226 (N_226,In_366,In_35);
and U227 (N_227,In_347,In_51);
nor U228 (N_228,In_620,In_686);
nand U229 (N_229,In_254,In_260);
xnor U230 (N_230,In_2,In_571);
nand U231 (N_231,In_523,In_626);
nand U232 (N_232,In_740,In_253);
xor U233 (N_233,In_94,In_324);
or U234 (N_234,In_472,In_65);
or U235 (N_235,In_186,In_606);
and U236 (N_236,In_49,In_108);
xnor U237 (N_237,In_579,In_362);
nor U238 (N_238,In_99,In_493);
or U239 (N_239,In_132,In_251);
nor U240 (N_240,In_738,In_559);
or U241 (N_241,In_705,In_334);
nand U242 (N_242,In_666,In_349);
nand U243 (N_243,In_121,In_11);
xnor U244 (N_244,In_210,In_119);
nand U245 (N_245,In_639,In_41);
nand U246 (N_246,In_54,In_264);
or U247 (N_247,In_536,In_360);
nand U248 (N_248,In_660,In_619);
nor U249 (N_249,In_1,In_193);
xor U250 (N_250,In_698,In_473);
nand U251 (N_251,In_282,In_476);
nor U252 (N_252,In_292,In_391);
and U253 (N_253,In_655,In_654);
nor U254 (N_254,In_663,In_342);
nor U255 (N_255,In_153,In_726);
or U256 (N_256,In_8,In_340);
nand U257 (N_257,In_138,In_327);
or U258 (N_258,In_118,In_321);
nand U259 (N_259,In_357,In_117);
nor U260 (N_260,In_189,In_688);
nor U261 (N_261,In_20,In_278);
nand U262 (N_262,In_316,In_82);
nor U263 (N_263,In_640,In_495);
nor U264 (N_264,In_291,In_561);
or U265 (N_265,In_36,In_584);
nor U266 (N_266,In_592,In_274);
xnor U267 (N_267,In_328,In_529);
or U268 (N_268,In_162,In_387);
xnor U269 (N_269,In_378,In_505);
nand U270 (N_270,In_217,In_232);
and U271 (N_271,In_723,In_724);
nor U272 (N_272,In_486,In_369);
nor U273 (N_273,In_15,In_419);
or U274 (N_274,In_736,In_707);
nor U275 (N_275,In_225,In_456);
or U276 (N_276,In_625,In_370);
or U277 (N_277,In_371,In_386);
nor U278 (N_278,In_503,In_92);
nor U279 (N_279,In_556,In_307);
nor U280 (N_280,In_40,In_509);
nand U281 (N_281,In_455,In_519);
nand U282 (N_282,In_535,In_368);
nand U283 (N_283,In_527,In_730);
and U284 (N_284,In_243,In_333);
and U285 (N_285,In_26,In_365);
xnor U286 (N_286,In_299,In_725);
or U287 (N_287,In_113,In_337);
nand U288 (N_288,In_465,In_171);
nand U289 (N_289,In_245,In_533);
or U290 (N_290,In_422,In_552);
nor U291 (N_291,In_466,In_662);
xnor U292 (N_292,In_173,In_175);
nor U293 (N_293,In_223,In_679);
xnor U294 (N_294,In_701,In_123);
or U295 (N_295,In_539,In_548);
and U296 (N_296,In_613,In_5);
or U297 (N_297,In_421,In_283);
and U298 (N_298,In_413,In_406);
nor U299 (N_299,In_55,In_176);
xnor U300 (N_300,In_296,In_735);
nand U301 (N_301,In_485,In_414);
nor U302 (N_302,In_601,In_167);
and U303 (N_303,In_269,In_13);
nand U304 (N_304,In_32,In_348);
nor U305 (N_305,In_435,In_154);
xor U306 (N_306,In_50,In_256);
nand U307 (N_307,In_122,In_75);
nor U308 (N_308,In_630,In_507);
xor U309 (N_309,In_470,In_446);
xor U310 (N_310,In_145,In_259);
nor U311 (N_311,In_129,In_134);
nor U312 (N_312,In_241,In_732);
nand U313 (N_313,In_314,In_281);
nand U314 (N_314,In_257,In_266);
xor U315 (N_315,In_70,In_549);
or U316 (N_316,In_677,In_164);
xor U317 (N_317,In_265,In_3);
xnor U318 (N_318,In_445,In_377);
xnor U319 (N_319,In_332,In_608);
nor U320 (N_320,In_746,In_66);
and U321 (N_321,In_574,In_77);
nor U322 (N_322,In_498,In_647);
and U323 (N_323,In_528,In_394);
xnor U324 (N_324,In_45,In_722);
nand U325 (N_325,In_303,In_590);
or U326 (N_326,In_90,In_308);
and U327 (N_327,In_614,In_233);
or U328 (N_328,In_336,In_474);
or U329 (N_329,In_181,In_131);
xor U330 (N_330,In_300,In_744);
nor U331 (N_331,In_504,In_646);
or U332 (N_332,In_379,In_560);
and U333 (N_333,In_81,In_191);
or U334 (N_334,In_635,In_228);
nor U335 (N_335,In_242,In_396);
and U336 (N_336,In_491,In_564);
xnor U337 (N_337,In_637,In_506);
nand U338 (N_338,In_76,In_384);
xnor U339 (N_339,In_658,In_353);
and U340 (N_340,In_616,In_127);
and U341 (N_341,In_78,In_224);
nand U342 (N_342,In_652,In_56);
nand U343 (N_343,In_656,In_748);
xor U344 (N_344,In_464,In_235);
and U345 (N_345,In_302,In_531);
and U346 (N_346,In_511,In_568);
or U347 (N_347,In_240,In_526);
nor U348 (N_348,In_695,In_372);
nand U349 (N_349,In_188,In_170);
nor U350 (N_350,In_161,In_234);
nand U351 (N_351,In_543,In_718);
xor U352 (N_352,In_468,In_399);
xor U353 (N_353,In_581,In_31);
and U354 (N_354,In_177,In_367);
or U355 (N_355,In_33,In_325);
or U356 (N_356,In_516,In_633);
xor U357 (N_357,In_411,In_452);
or U358 (N_358,In_605,In_267);
xor U359 (N_359,In_159,In_522);
or U360 (N_360,In_313,In_629);
or U361 (N_361,In_589,In_621);
or U362 (N_362,In_697,In_339);
nor U363 (N_363,In_246,In_6);
or U364 (N_364,In_672,In_375);
xnor U365 (N_365,In_423,In_444);
nor U366 (N_366,In_218,In_68);
nand U367 (N_367,In_201,In_277);
nand U368 (N_368,In_407,In_612);
nand U369 (N_369,In_547,In_681);
xor U370 (N_370,In_312,In_230);
xnor U371 (N_371,In_98,In_636);
nor U372 (N_372,In_494,In_659);
nor U373 (N_373,In_609,In_211);
nand U374 (N_374,In_376,In_335);
xor U375 (N_375,In_69,In_116);
and U376 (N_376,In_107,In_375);
nand U377 (N_377,In_108,In_496);
or U378 (N_378,In_313,In_256);
and U379 (N_379,In_101,In_17);
nor U380 (N_380,In_171,In_325);
xnor U381 (N_381,In_244,In_265);
and U382 (N_382,In_719,In_527);
nand U383 (N_383,In_651,In_27);
nor U384 (N_384,In_189,In_464);
xor U385 (N_385,In_115,In_12);
nor U386 (N_386,In_195,In_186);
nand U387 (N_387,In_300,In_711);
xnor U388 (N_388,In_115,In_616);
xor U389 (N_389,In_323,In_135);
or U390 (N_390,In_431,In_385);
nor U391 (N_391,In_253,In_303);
nand U392 (N_392,In_14,In_378);
or U393 (N_393,In_290,In_38);
xnor U394 (N_394,In_491,In_554);
or U395 (N_395,In_392,In_298);
or U396 (N_396,In_439,In_202);
and U397 (N_397,In_158,In_338);
xor U398 (N_398,In_450,In_372);
and U399 (N_399,In_586,In_21);
xnor U400 (N_400,In_376,In_104);
and U401 (N_401,In_373,In_570);
xor U402 (N_402,In_316,In_65);
xor U403 (N_403,In_118,In_636);
nand U404 (N_404,In_101,In_633);
nor U405 (N_405,In_715,In_655);
nand U406 (N_406,In_154,In_30);
and U407 (N_407,In_670,In_735);
or U408 (N_408,In_110,In_175);
or U409 (N_409,In_712,In_471);
or U410 (N_410,In_479,In_440);
or U411 (N_411,In_398,In_594);
xnor U412 (N_412,In_312,In_454);
or U413 (N_413,In_623,In_55);
and U414 (N_414,In_145,In_541);
xnor U415 (N_415,In_486,In_392);
and U416 (N_416,In_298,In_658);
nor U417 (N_417,In_418,In_604);
nor U418 (N_418,In_333,In_636);
or U419 (N_419,In_164,In_736);
and U420 (N_420,In_610,In_49);
and U421 (N_421,In_88,In_205);
and U422 (N_422,In_383,In_435);
nor U423 (N_423,In_546,In_488);
nand U424 (N_424,In_245,In_334);
or U425 (N_425,In_498,In_243);
or U426 (N_426,In_437,In_552);
nand U427 (N_427,In_101,In_690);
nand U428 (N_428,In_97,In_625);
nor U429 (N_429,In_532,In_481);
xor U430 (N_430,In_442,In_232);
xor U431 (N_431,In_560,In_183);
nor U432 (N_432,In_277,In_31);
and U433 (N_433,In_544,In_593);
and U434 (N_434,In_295,In_270);
or U435 (N_435,In_621,In_622);
xnor U436 (N_436,In_726,In_40);
xnor U437 (N_437,In_574,In_745);
nor U438 (N_438,In_666,In_425);
nor U439 (N_439,In_118,In_492);
and U440 (N_440,In_199,In_423);
xnor U441 (N_441,In_744,In_87);
or U442 (N_442,In_687,In_484);
xnor U443 (N_443,In_651,In_638);
and U444 (N_444,In_409,In_536);
or U445 (N_445,In_395,In_304);
nor U446 (N_446,In_572,In_499);
and U447 (N_447,In_60,In_628);
and U448 (N_448,In_684,In_359);
xnor U449 (N_449,In_314,In_203);
nand U450 (N_450,In_116,In_686);
and U451 (N_451,In_558,In_8);
nand U452 (N_452,In_664,In_85);
or U453 (N_453,In_648,In_688);
or U454 (N_454,In_208,In_35);
nor U455 (N_455,In_456,In_122);
nand U456 (N_456,In_66,In_670);
xor U457 (N_457,In_534,In_375);
nor U458 (N_458,In_116,In_363);
xor U459 (N_459,In_151,In_68);
or U460 (N_460,In_497,In_17);
and U461 (N_461,In_574,In_100);
nand U462 (N_462,In_428,In_638);
nand U463 (N_463,In_587,In_492);
xor U464 (N_464,In_62,In_561);
xor U465 (N_465,In_149,In_184);
nand U466 (N_466,In_285,In_56);
and U467 (N_467,In_565,In_628);
and U468 (N_468,In_600,In_127);
and U469 (N_469,In_88,In_234);
and U470 (N_470,In_140,In_575);
nor U471 (N_471,In_400,In_419);
nor U472 (N_472,In_69,In_450);
xor U473 (N_473,In_135,In_582);
nand U474 (N_474,In_204,In_272);
or U475 (N_475,In_542,In_46);
nor U476 (N_476,In_592,In_642);
nor U477 (N_477,In_708,In_246);
nor U478 (N_478,In_147,In_665);
or U479 (N_479,In_630,In_408);
or U480 (N_480,In_420,In_362);
nor U481 (N_481,In_393,In_171);
and U482 (N_482,In_219,In_352);
nand U483 (N_483,In_395,In_447);
and U484 (N_484,In_735,In_632);
xnor U485 (N_485,In_311,In_701);
and U486 (N_486,In_320,In_537);
nand U487 (N_487,In_650,In_200);
nand U488 (N_488,In_10,In_57);
and U489 (N_489,In_32,In_340);
nand U490 (N_490,In_576,In_477);
nor U491 (N_491,In_321,In_345);
xnor U492 (N_492,In_268,In_241);
xnor U493 (N_493,In_113,In_164);
or U494 (N_494,In_611,In_617);
nor U495 (N_495,In_64,In_449);
nand U496 (N_496,In_95,In_513);
and U497 (N_497,In_433,In_631);
or U498 (N_498,In_338,In_112);
nand U499 (N_499,In_3,In_407);
and U500 (N_500,In_461,In_247);
xnor U501 (N_501,In_472,In_685);
xor U502 (N_502,In_668,In_142);
and U503 (N_503,In_388,In_288);
and U504 (N_504,In_461,In_64);
xnor U505 (N_505,In_270,In_339);
xor U506 (N_506,In_112,In_145);
xor U507 (N_507,In_269,In_372);
and U508 (N_508,In_348,In_271);
or U509 (N_509,In_503,In_229);
xor U510 (N_510,In_179,In_743);
nor U511 (N_511,In_457,In_351);
nand U512 (N_512,In_663,In_1);
xnor U513 (N_513,In_229,In_391);
or U514 (N_514,In_342,In_217);
nand U515 (N_515,In_616,In_173);
and U516 (N_516,In_427,In_79);
nor U517 (N_517,In_31,In_626);
and U518 (N_518,In_37,In_577);
nand U519 (N_519,In_91,In_472);
nand U520 (N_520,In_214,In_386);
xnor U521 (N_521,In_424,In_713);
nor U522 (N_522,In_5,In_585);
or U523 (N_523,In_126,In_588);
and U524 (N_524,In_614,In_570);
nand U525 (N_525,In_430,In_278);
and U526 (N_526,In_551,In_519);
or U527 (N_527,In_679,In_672);
nand U528 (N_528,In_57,In_560);
xnor U529 (N_529,In_717,In_340);
and U530 (N_530,In_331,In_704);
or U531 (N_531,In_45,In_209);
xnor U532 (N_532,In_136,In_705);
nor U533 (N_533,In_186,In_639);
xnor U534 (N_534,In_174,In_307);
nand U535 (N_535,In_576,In_590);
xor U536 (N_536,In_119,In_230);
or U537 (N_537,In_191,In_375);
nand U538 (N_538,In_556,In_421);
or U539 (N_539,In_727,In_141);
nand U540 (N_540,In_344,In_280);
nand U541 (N_541,In_507,In_46);
or U542 (N_542,In_695,In_347);
and U543 (N_543,In_81,In_702);
or U544 (N_544,In_365,In_544);
nand U545 (N_545,In_605,In_9);
or U546 (N_546,In_697,In_660);
nand U547 (N_547,In_157,In_693);
or U548 (N_548,In_251,In_486);
and U549 (N_549,In_374,In_28);
nand U550 (N_550,In_716,In_191);
nor U551 (N_551,In_420,In_599);
and U552 (N_552,In_235,In_741);
or U553 (N_553,In_685,In_513);
nor U554 (N_554,In_491,In_660);
nor U555 (N_555,In_14,In_120);
nand U556 (N_556,In_503,In_38);
nand U557 (N_557,In_547,In_709);
xor U558 (N_558,In_661,In_529);
and U559 (N_559,In_212,In_234);
and U560 (N_560,In_723,In_112);
xor U561 (N_561,In_14,In_712);
nand U562 (N_562,In_349,In_385);
nand U563 (N_563,In_409,In_163);
xnor U564 (N_564,In_652,In_744);
or U565 (N_565,In_601,In_701);
and U566 (N_566,In_655,In_458);
nand U567 (N_567,In_47,In_265);
or U568 (N_568,In_608,In_578);
xor U569 (N_569,In_495,In_401);
or U570 (N_570,In_495,In_232);
or U571 (N_571,In_214,In_14);
or U572 (N_572,In_415,In_632);
and U573 (N_573,In_342,In_581);
nand U574 (N_574,In_264,In_661);
nand U575 (N_575,In_501,In_282);
nand U576 (N_576,In_107,In_638);
or U577 (N_577,In_305,In_418);
nand U578 (N_578,In_185,In_502);
and U579 (N_579,In_350,In_110);
or U580 (N_580,In_545,In_508);
nor U581 (N_581,In_494,In_596);
and U582 (N_582,In_374,In_532);
xor U583 (N_583,In_112,In_439);
nand U584 (N_584,In_323,In_738);
nand U585 (N_585,In_725,In_723);
or U586 (N_586,In_235,In_416);
or U587 (N_587,In_42,In_71);
or U588 (N_588,In_493,In_511);
nand U589 (N_589,In_645,In_197);
xnor U590 (N_590,In_577,In_278);
or U591 (N_591,In_577,In_365);
or U592 (N_592,In_124,In_492);
and U593 (N_593,In_58,In_623);
or U594 (N_594,In_397,In_282);
nor U595 (N_595,In_81,In_510);
and U596 (N_596,In_189,In_400);
and U597 (N_597,In_646,In_651);
or U598 (N_598,In_459,In_92);
nor U599 (N_599,In_663,In_370);
nand U600 (N_600,In_527,In_397);
or U601 (N_601,In_80,In_733);
and U602 (N_602,In_684,In_8);
nor U603 (N_603,In_731,In_685);
nor U604 (N_604,In_299,In_686);
or U605 (N_605,In_607,In_237);
nor U606 (N_606,In_139,In_357);
nor U607 (N_607,In_83,In_277);
xor U608 (N_608,In_494,In_50);
and U609 (N_609,In_466,In_639);
or U610 (N_610,In_509,In_522);
or U611 (N_611,In_185,In_27);
nor U612 (N_612,In_169,In_123);
or U613 (N_613,In_430,In_254);
and U614 (N_614,In_56,In_15);
nand U615 (N_615,In_612,In_110);
nand U616 (N_616,In_80,In_683);
and U617 (N_617,In_632,In_680);
and U618 (N_618,In_721,In_233);
or U619 (N_619,In_560,In_648);
xor U620 (N_620,In_13,In_308);
or U621 (N_621,In_35,In_217);
nor U622 (N_622,In_213,In_13);
and U623 (N_623,In_715,In_13);
nand U624 (N_624,In_686,In_121);
xor U625 (N_625,In_63,In_215);
xor U626 (N_626,In_662,In_53);
and U627 (N_627,In_88,In_4);
nand U628 (N_628,In_352,In_429);
nor U629 (N_629,In_636,In_313);
xor U630 (N_630,In_21,In_153);
nand U631 (N_631,In_634,In_666);
or U632 (N_632,In_144,In_57);
nor U633 (N_633,In_667,In_312);
and U634 (N_634,In_332,In_662);
and U635 (N_635,In_559,In_234);
or U636 (N_636,In_363,In_61);
or U637 (N_637,In_288,In_520);
nand U638 (N_638,In_576,In_749);
nor U639 (N_639,In_350,In_637);
and U640 (N_640,In_558,In_418);
nor U641 (N_641,In_241,In_353);
nor U642 (N_642,In_582,In_485);
nand U643 (N_643,In_627,In_740);
or U644 (N_644,In_110,In_663);
xnor U645 (N_645,In_356,In_330);
xnor U646 (N_646,In_319,In_426);
xor U647 (N_647,In_267,In_565);
nand U648 (N_648,In_158,In_3);
and U649 (N_649,In_115,In_624);
or U650 (N_650,In_615,In_629);
nand U651 (N_651,In_380,In_382);
or U652 (N_652,In_108,In_740);
xnor U653 (N_653,In_444,In_344);
or U654 (N_654,In_274,In_57);
or U655 (N_655,In_369,In_749);
or U656 (N_656,In_649,In_269);
or U657 (N_657,In_327,In_664);
nor U658 (N_658,In_240,In_519);
nor U659 (N_659,In_264,In_524);
and U660 (N_660,In_106,In_551);
xor U661 (N_661,In_749,In_270);
xor U662 (N_662,In_103,In_233);
or U663 (N_663,In_730,In_674);
nor U664 (N_664,In_27,In_340);
or U665 (N_665,In_52,In_81);
and U666 (N_666,In_80,In_546);
nand U667 (N_667,In_196,In_154);
xnor U668 (N_668,In_2,In_285);
xor U669 (N_669,In_38,In_137);
xor U670 (N_670,In_520,In_64);
and U671 (N_671,In_455,In_79);
xor U672 (N_672,In_465,In_249);
and U673 (N_673,In_36,In_535);
or U674 (N_674,In_328,In_77);
or U675 (N_675,In_427,In_337);
and U676 (N_676,In_593,In_615);
and U677 (N_677,In_72,In_28);
nor U678 (N_678,In_610,In_147);
or U679 (N_679,In_688,In_465);
or U680 (N_680,In_93,In_640);
and U681 (N_681,In_590,In_243);
xor U682 (N_682,In_144,In_237);
or U683 (N_683,In_459,In_739);
xor U684 (N_684,In_36,In_652);
or U685 (N_685,In_327,In_620);
nand U686 (N_686,In_285,In_180);
nand U687 (N_687,In_12,In_494);
nor U688 (N_688,In_9,In_179);
or U689 (N_689,In_33,In_231);
nand U690 (N_690,In_197,In_554);
xnor U691 (N_691,In_168,In_151);
and U692 (N_692,In_79,In_506);
xnor U693 (N_693,In_60,In_247);
nand U694 (N_694,In_298,In_249);
nor U695 (N_695,In_454,In_128);
or U696 (N_696,In_173,In_538);
nor U697 (N_697,In_156,In_720);
xor U698 (N_698,In_101,In_597);
nand U699 (N_699,In_538,In_355);
nand U700 (N_700,In_274,In_118);
xor U701 (N_701,In_325,In_603);
nor U702 (N_702,In_748,In_749);
or U703 (N_703,In_675,In_552);
and U704 (N_704,In_258,In_229);
or U705 (N_705,In_555,In_539);
nor U706 (N_706,In_489,In_352);
nand U707 (N_707,In_567,In_22);
and U708 (N_708,In_175,In_39);
or U709 (N_709,In_564,In_725);
nand U710 (N_710,In_28,In_93);
or U711 (N_711,In_28,In_531);
nor U712 (N_712,In_145,In_717);
or U713 (N_713,In_227,In_148);
nand U714 (N_714,In_272,In_102);
nor U715 (N_715,In_245,In_301);
nor U716 (N_716,In_504,In_46);
nor U717 (N_717,In_439,In_433);
and U718 (N_718,In_67,In_3);
nor U719 (N_719,In_636,In_538);
and U720 (N_720,In_10,In_144);
nand U721 (N_721,In_187,In_679);
xor U722 (N_722,In_62,In_694);
or U723 (N_723,In_20,In_360);
nand U724 (N_724,In_114,In_581);
xor U725 (N_725,In_410,In_19);
nor U726 (N_726,In_229,In_745);
nor U727 (N_727,In_138,In_492);
nand U728 (N_728,In_23,In_679);
and U729 (N_729,In_521,In_687);
nand U730 (N_730,In_668,In_249);
xnor U731 (N_731,In_725,In_342);
and U732 (N_732,In_118,In_512);
and U733 (N_733,In_246,In_107);
nor U734 (N_734,In_597,In_0);
and U735 (N_735,In_749,In_355);
nor U736 (N_736,In_173,In_653);
or U737 (N_737,In_667,In_10);
xnor U738 (N_738,In_264,In_277);
nand U739 (N_739,In_563,In_287);
xor U740 (N_740,In_81,In_32);
or U741 (N_741,In_156,In_341);
nor U742 (N_742,In_595,In_690);
nand U743 (N_743,In_134,In_139);
or U744 (N_744,In_265,In_397);
xor U745 (N_745,In_177,In_369);
nor U746 (N_746,In_164,In_204);
or U747 (N_747,In_694,In_530);
or U748 (N_748,In_146,In_314);
nand U749 (N_749,In_599,In_126);
and U750 (N_750,In_229,In_730);
or U751 (N_751,In_593,In_395);
xor U752 (N_752,In_598,In_124);
nand U753 (N_753,In_146,In_353);
xnor U754 (N_754,In_524,In_378);
nand U755 (N_755,In_258,In_372);
nor U756 (N_756,In_656,In_671);
nor U757 (N_757,In_324,In_398);
or U758 (N_758,In_517,In_369);
nand U759 (N_759,In_693,In_185);
or U760 (N_760,In_350,In_270);
and U761 (N_761,In_144,In_460);
nor U762 (N_762,In_664,In_259);
or U763 (N_763,In_744,In_573);
nor U764 (N_764,In_10,In_99);
nand U765 (N_765,In_351,In_343);
and U766 (N_766,In_569,In_563);
or U767 (N_767,In_364,In_325);
nand U768 (N_768,In_104,In_385);
xnor U769 (N_769,In_491,In_180);
nand U770 (N_770,In_510,In_742);
nand U771 (N_771,In_476,In_260);
and U772 (N_772,In_488,In_706);
nand U773 (N_773,In_574,In_385);
nand U774 (N_774,In_462,In_637);
nand U775 (N_775,In_209,In_11);
xor U776 (N_776,In_362,In_193);
nor U777 (N_777,In_493,In_54);
and U778 (N_778,In_489,In_477);
and U779 (N_779,In_652,In_690);
xor U780 (N_780,In_395,In_375);
nor U781 (N_781,In_213,In_456);
and U782 (N_782,In_625,In_675);
nor U783 (N_783,In_656,In_60);
xor U784 (N_784,In_526,In_397);
and U785 (N_785,In_361,In_160);
or U786 (N_786,In_662,In_546);
nor U787 (N_787,In_609,In_543);
nor U788 (N_788,In_147,In_501);
nor U789 (N_789,In_286,In_320);
nor U790 (N_790,In_39,In_517);
xnor U791 (N_791,In_162,In_608);
nand U792 (N_792,In_272,In_320);
and U793 (N_793,In_93,In_668);
nor U794 (N_794,In_99,In_117);
and U795 (N_795,In_216,In_218);
and U796 (N_796,In_479,In_304);
xor U797 (N_797,In_725,In_560);
xnor U798 (N_798,In_255,In_89);
xor U799 (N_799,In_139,In_610);
nand U800 (N_800,In_447,In_164);
nor U801 (N_801,In_622,In_385);
nor U802 (N_802,In_710,In_230);
or U803 (N_803,In_473,In_26);
and U804 (N_804,In_363,In_569);
xor U805 (N_805,In_683,In_444);
and U806 (N_806,In_679,In_748);
or U807 (N_807,In_360,In_569);
or U808 (N_808,In_378,In_658);
or U809 (N_809,In_381,In_18);
and U810 (N_810,In_594,In_609);
xor U811 (N_811,In_184,In_528);
nor U812 (N_812,In_221,In_685);
nand U813 (N_813,In_168,In_407);
xnor U814 (N_814,In_183,In_205);
or U815 (N_815,In_182,In_277);
or U816 (N_816,In_191,In_11);
xnor U817 (N_817,In_674,In_503);
nand U818 (N_818,In_466,In_697);
xnor U819 (N_819,In_573,In_593);
or U820 (N_820,In_581,In_627);
nand U821 (N_821,In_671,In_648);
xnor U822 (N_822,In_197,In_747);
xnor U823 (N_823,In_15,In_310);
or U824 (N_824,In_512,In_188);
nor U825 (N_825,In_737,In_308);
nand U826 (N_826,In_539,In_684);
and U827 (N_827,In_327,In_308);
nor U828 (N_828,In_385,In_430);
xor U829 (N_829,In_569,In_118);
nor U830 (N_830,In_690,In_467);
or U831 (N_831,In_166,In_723);
nand U832 (N_832,In_350,In_742);
and U833 (N_833,In_737,In_454);
nor U834 (N_834,In_505,In_300);
and U835 (N_835,In_676,In_173);
or U836 (N_836,In_132,In_596);
or U837 (N_837,In_430,In_248);
nand U838 (N_838,In_24,In_154);
nor U839 (N_839,In_94,In_145);
xnor U840 (N_840,In_380,In_448);
nor U841 (N_841,In_59,In_423);
or U842 (N_842,In_505,In_440);
or U843 (N_843,In_497,In_638);
nand U844 (N_844,In_66,In_25);
nor U845 (N_845,In_349,In_116);
nand U846 (N_846,In_0,In_370);
and U847 (N_847,In_194,In_223);
nand U848 (N_848,In_137,In_562);
nand U849 (N_849,In_184,In_115);
or U850 (N_850,In_80,In_93);
xor U851 (N_851,In_747,In_677);
xor U852 (N_852,In_745,In_127);
nand U853 (N_853,In_434,In_222);
or U854 (N_854,In_214,In_51);
or U855 (N_855,In_392,In_526);
nor U856 (N_856,In_126,In_403);
nand U857 (N_857,In_647,In_539);
nand U858 (N_858,In_341,In_131);
nand U859 (N_859,In_376,In_47);
nand U860 (N_860,In_527,In_619);
nand U861 (N_861,In_564,In_293);
and U862 (N_862,In_153,In_119);
xor U863 (N_863,In_127,In_125);
nor U864 (N_864,In_180,In_88);
xnor U865 (N_865,In_703,In_431);
and U866 (N_866,In_308,In_319);
and U867 (N_867,In_193,In_695);
nor U868 (N_868,In_294,In_137);
nor U869 (N_869,In_34,In_242);
or U870 (N_870,In_735,In_118);
xnor U871 (N_871,In_635,In_428);
nand U872 (N_872,In_405,In_218);
nand U873 (N_873,In_608,In_265);
nand U874 (N_874,In_357,In_214);
or U875 (N_875,In_200,In_728);
xnor U876 (N_876,In_651,In_398);
or U877 (N_877,In_580,In_433);
and U878 (N_878,In_704,In_381);
nor U879 (N_879,In_675,In_317);
nand U880 (N_880,In_492,In_713);
or U881 (N_881,In_709,In_147);
xor U882 (N_882,In_145,In_357);
xor U883 (N_883,In_529,In_261);
xnor U884 (N_884,In_437,In_343);
or U885 (N_885,In_557,In_280);
nor U886 (N_886,In_720,In_393);
nor U887 (N_887,In_559,In_732);
xor U888 (N_888,In_443,In_1);
xnor U889 (N_889,In_495,In_686);
or U890 (N_890,In_506,In_89);
nor U891 (N_891,In_275,In_228);
xnor U892 (N_892,In_734,In_45);
or U893 (N_893,In_575,In_320);
or U894 (N_894,In_147,In_130);
nand U895 (N_895,In_621,In_450);
or U896 (N_896,In_745,In_429);
xor U897 (N_897,In_126,In_428);
or U898 (N_898,In_215,In_519);
and U899 (N_899,In_69,In_93);
or U900 (N_900,In_253,In_217);
xnor U901 (N_901,In_586,In_516);
or U902 (N_902,In_711,In_1);
and U903 (N_903,In_359,In_530);
and U904 (N_904,In_591,In_539);
or U905 (N_905,In_231,In_180);
nand U906 (N_906,In_192,In_474);
nor U907 (N_907,In_645,In_111);
nand U908 (N_908,In_615,In_470);
and U909 (N_909,In_188,In_681);
nor U910 (N_910,In_104,In_643);
nand U911 (N_911,In_681,In_693);
nor U912 (N_912,In_630,In_99);
xor U913 (N_913,In_673,In_369);
and U914 (N_914,In_441,In_560);
nand U915 (N_915,In_308,In_254);
xnor U916 (N_916,In_77,In_153);
nor U917 (N_917,In_437,In_517);
xor U918 (N_918,In_631,In_497);
nand U919 (N_919,In_468,In_231);
nor U920 (N_920,In_246,In_468);
nor U921 (N_921,In_532,In_540);
and U922 (N_922,In_75,In_546);
nand U923 (N_923,In_182,In_687);
or U924 (N_924,In_462,In_234);
or U925 (N_925,In_107,In_411);
nor U926 (N_926,In_75,In_511);
nand U927 (N_927,In_669,In_203);
or U928 (N_928,In_622,In_217);
and U929 (N_929,In_564,In_708);
xor U930 (N_930,In_86,In_95);
xnor U931 (N_931,In_381,In_393);
or U932 (N_932,In_642,In_672);
nand U933 (N_933,In_290,In_186);
and U934 (N_934,In_740,In_24);
or U935 (N_935,In_158,In_167);
and U936 (N_936,In_708,In_670);
nor U937 (N_937,In_667,In_692);
nand U938 (N_938,In_49,In_190);
nor U939 (N_939,In_191,In_39);
and U940 (N_940,In_233,In_570);
xor U941 (N_941,In_179,In_379);
or U942 (N_942,In_188,In_743);
nor U943 (N_943,In_298,In_326);
nor U944 (N_944,In_111,In_206);
nand U945 (N_945,In_701,In_357);
and U946 (N_946,In_39,In_6);
nor U947 (N_947,In_52,In_385);
xnor U948 (N_948,In_219,In_71);
nor U949 (N_949,In_264,In_465);
or U950 (N_950,In_134,In_513);
xor U951 (N_951,In_335,In_282);
and U952 (N_952,In_697,In_548);
nand U953 (N_953,In_440,In_301);
and U954 (N_954,In_14,In_498);
or U955 (N_955,In_241,In_131);
and U956 (N_956,In_237,In_105);
nor U957 (N_957,In_417,In_544);
nor U958 (N_958,In_500,In_292);
nor U959 (N_959,In_429,In_89);
xnor U960 (N_960,In_401,In_427);
xor U961 (N_961,In_123,In_513);
xor U962 (N_962,In_328,In_582);
or U963 (N_963,In_508,In_633);
nor U964 (N_964,In_65,In_2);
nor U965 (N_965,In_613,In_20);
nor U966 (N_966,In_432,In_220);
xnor U967 (N_967,In_643,In_717);
nand U968 (N_968,In_686,In_87);
or U969 (N_969,In_121,In_640);
nor U970 (N_970,In_453,In_42);
or U971 (N_971,In_434,In_216);
nand U972 (N_972,In_637,In_705);
nor U973 (N_973,In_231,In_444);
nor U974 (N_974,In_21,In_417);
and U975 (N_975,In_230,In_426);
nor U976 (N_976,In_451,In_680);
and U977 (N_977,In_724,In_483);
and U978 (N_978,In_391,In_87);
nor U979 (N_979,In_77,In_29);
nand U980 (N_980,In_621,In_171);
and U981 (N_981,In_29,In_358);
nor U982 (N_982,In_547,In_15);
nor U983 (N_983,In_537,In_11);
nor U984 (N_984,In_725,In_335);
xor U985 (N_985,In_466,In_56);
or U986 (N_986,In_58,In_120);
nand U987 (N_987,In_61,In_63);
xor U988 (N_988,In_432,In_41);
or U989 (N_989,In_310,In_86);
or U990 (N_990,In_150,In_174);
or U991 (N_991,In_163,In_184);
and U992 (N_992,In_729,In_348);
nand U993 (N_993,In_492,In_328);
xor U994 (N_994,In_509,In_612);
xnor U995 (N_995,In_498,In_299);
nor U996 (N_996,In_435,In_38);
xor U997 (N_997,In_200,In_125);
and U998 (N_998,In_360,In_496);
nor U999 (N_999,In_420,In_740);
and U1000 (N_1000,N_801,N_361);
nor U1001 (N_1001,N_668,N_536);
nand U1002 (N_1002,N_627,N_466);
and U1003 (N_1003,N_686,N_243);
nor U1004 (N_1004,N_57,N_484);
nand U1005 (N_1005,N_750,N_184);
nor U1006 (N_1006,N_73,N_939);
nor U1007 (N_1007,N_395,N_103);
and U1008 (N_1008,N_274,N_837);
nand U1009 (N_1009,N_676,N_33);
nor U1010 (N_1010,N_611,N_502);
nor U1011 (N_1011,N_157,N_195);
nand U1012 (N_1012,N_222,N_400);
or U1013 (N_1013,N_964,N_945);
or U1014 (N_1014,N_598,N_424);
nor U1015 (N_1015,N_820,N_476);
nor U1016 (N_1016,N_538,N_467);
xnor U1017 (N_1017,N_75,N_171);
xor U1018 (N_1018,N_997,N_50);
or U1019 (N_1019,N_143,N_416);
and U1020 (N_1020,N_347,N_90);
nor U1021 (N_1021,N_960,N_373);
xnor U1022 (N_1022,N_398,N_998);
and U1023 (N_1023,N_43,N_612);
xor U1024 (N_1024,N_636,N_615);
nor U1025 (N_1025,N_3,N_7);
and U1026 (N_1026,N_827,N_712);
nand U1027 (N_1027,N_115,N_851);
nand U1028 (N_1028,N_664,N_803);
nor U1029 (N_1029,N_950,N_591);
or U1030 (N_1030,N_432,N_463);
xnor U1031 (N_1031,N_849,N_113);
or U1032 (N_1032,N_863,N_443);
nor U1033 (N_1033,N_220,N_64);
and U1034 (N_1034,N_568,N_899);
xnor U1035 (N_1035,N_815,N_540);
nor U1036 (N_1036,N_300,N_177);
and U1037 (N_1037,N_437,N_341);
or U1038 (N_1038,N_384,N_768);
nor U1039 (N_1039,N_358,N_897);
nand U1040 (N_1040,N_67,N_826);
or U1041 (N_1041,N_532,N_715);
or U1042 (N_1042,N_814,N_747);
nor U1043 (N_1043,N_218,N_892);
nand U1044 (N_1044,N_819,N_645);
and U1045 (N_1045,N_138,N_282);
xor U1046 (N_1046,N_527,N_778);
and U1047 (N_1047,N_971,N_531);
nor U1048 (N_1048,N_264,N_24);
nor U1049 (N_1049,N_936,N_185);
nand U1050 (N_1050,N_306,N_574);
xor U1051 (N_1051,N_528,N_418);
nor U1052 (N_1052,N_952,N_112);
xnor U1053 (N_1053,N_757,N_925);
or U1054 (N_1054,N_411,N_391);
nor U1055 (N_1055,N_514,N_326);
or U1056 (N_1056,N_900,N_507);
or U1057 (N_1057,N_60,N_500);
or U1058 (N_1058,N_216,N_412);
and U1059 (N_1059,N_436,N_253);
and U1060 (N_1060,N_131,N_82);
xor U1061 (N_1061,N_992,N_891);
nand U1062 (N_1062,N_367,N_335);
nand U1063 (N_1063,N_553,N_984);
or U1064 (N_1064,N_250,N_859);
nand U1065 (N_1065,N_640,N_551);
nand U1066 (N_1066,N_135,N_555);
or U1067 (N_1067,N_771,N_908);
and U1068 (N_1068,N_816,N_456);
or U1069 (N_1069,N_840,N_213);
or U1070 (N_1070,N_45,N_372);
nor U1071 (N_1071,N_15,N_333);
and U1072 (N_1072,N_864,N_359);
xnor U1073 (N_1073,N_343,N_419);
or U1074 (N_1074,N_988,N_728);
xnor U1075 (N_1075,N_6,N_935);
or U1076 (N_1076,N_161,N_839);
xnor U1077 (N_1077,N_30,N_902);
nor U1078 (N_1078,N_922,N_348);
or U1079 (N_1079,N_46,N_989);
or U1080 (N_1080,N_807,N_552);
xnor U1081 (N_1081,N_37,N_408);
and U1082 (N_1082,N_59,N_522);
nand U1083 (N_1083,N_353,N_210);
and U1084 (N_1084,N_190,N_606);
and U1085 (N_1085,N_774,N_928);
xnor U1086 (N_1086,N_308,N_413);
and U1087 (N_1087,N_594,N_967);
xor U1088 (N_1088,N_550,N_77);
xnor U1089 (N_1089,N_219,N_236);
nor U1090 (N_1090,N_89,N_449);
and U1091 (N_1091,N_503,N_862);
nand U1092 (N_1092,N_71,N_610);
nor U1093 (N_1093,N_614,N_366);
xnor U1094 (N_1094,N_402,N_569);
xor U1095 (N_1095,N_710,N_619);
or U1096 (N_1096,N_524,N_795);
nand U1097 (N_1097,N_489,N_340);
or U1098 (N_1098,N_764,N_926);
or U1099 (N_1099,N_963,N_211);
nand U1100 (N_1100,N_872,N_84);
xnor U1101 (N_1101,N_278,N_773);
nand U1102 (N_1102,N_187,N_180);
nand U1103 (N_1103,N_453,N_338);
or U1104 (N_1104,N_110,N_323);
nand U1105 (N_1105,N_311,N_42);
nor U1106 (N_1106,N_792,N_812);
and U1107 (N_1107,N_356,N_968);
xnor U1108 (N_1108,N_566,N_172);
and U1109 (N_1109,N_633,N_106);
nand U1110 (N_1110,N_442,N_590);
nor U1111 (N_1111,N_973,N_886);
and U1112 (N_1112,N_593,N_705);
or U1113 (N_1113,N_128,N_123);
nor U1114 (N_1114,N_934,N_842);
xor U1115 (N_1115,N_208,N_10);
or U1116 (N_1116,N_369,N_345);
nand U1117 (N_1117,N_260,N_966);
or U1118 (N_1118,N_870,N_677);
or U1119 (N_1119,N_699,N_317);
nor U1120 (N_1120,N_144,N_125);
nand U1121 (N_1121,N_752,N_105);
or U1122 (N_1122,N_846,N_544);
xnor U1123 (N_1123,N_319,N_787);
or U1124 (N_1124,N_630,N_32);
nand U1125 (N_1125,N_255,N_702);
nor U1126 (N_1126,N_200,N_990);
or U1127 (N_1127,N_580,N_396);
xor U1128 (N_1128,N_501,N_206);
nand U1129 (N_1129,N_478,N_887);
nand U1130 (N_1130,N_469,N_920);
xnor U1131 (N_1131,N_533,N_941);
nor U1132 (N_1132,N_652,N_822);
nor U1133 (N_1133,N_513,N_257);
or U1134 (N_1134,N_35,N_25);
xor U1135 (N_1135,N_599,N_487);
or U1136 (N_1136,N_94,N_164);
xor U1137 (N_1137,N_87,N_504);
nor U1138 (N_1138,N_687,N_543);
or U1139 (N_1139,N_850,N_431);
and U1140 (N_1140,N_318,N_517);
and U1141 (N_1141,N_570,N_913);
xnor U1142 (N_1142,N_96,N_389);
or U1143 (N_1143,N_270,N_423);
nand U1144 (N_1144,N_944,N_604);
xor U1145 (N_1145,N_811,N_322);
nor U1146 (N_1146,N_102,N_21);
and U1147 (N_1147,N_706,N_777);
nor U1148 (N_1148,N_780,N_22);
nand U1149 (N_1149,N_393,N_735);
nand U1150 (N_1150,N_13,N_68);
xnor U1151 (N_1151,N_62,N_587);
or U1152 (N_1152,N_882,N_472);
nor U1153 (N_1153,N_394,N_556);
or U1154 (N_1154,N_756,N_344);
and U1155 (N_1155,N_267,N_695);
nor U1156 (N_1156,N_422,N_781);
and U1157 (N_1157,N_197,N_554);
nor U1158 (N_1158,N_404,N_738);
nand U1159 (N_1159,N_266,N_921);
nand U1160 (N_1160,N_249,N_217);
nor U1161 (N_1161,N_154,N_374);
nand U1162 (N_1162,N_49,N_616);
or U1163 (N_1163,N_224,N_12);
and U1164 (N_1164,N_831,N_938);
and U1165 (N_1165,N_262,N_54);
and U1166 (N_1166,N_387,N_621);
xor U1167 (N_1167,N_401,N_292);
nor U1168 (N_1168,N_644,N_1);
nand U1169 (N_1169,N_450,N_804);
xnor U1170 (N_1170,N_429,N_525);
xor U1171 (N_1171,N_198,N_709);
or U1172 (N_1172,N_101,N_956);
xnor U1173 (N_1173,N_798,N_910);
and U1174 (N_1174,N_537,N_203);
and U1175 (N_1175,N_579,N_914);
and U1176 (N_1176,N_916,N_231);
nand U1177 (N_1177,N_523,N_17);
or U1178 (N_1178,N_475,N_588);
nor U1179 (N_1179,N_854,N_767);
xor U1180 (N_1180,N_119,N_368);
xnor U1181 (N_1181,N_390,N_188);
xnor U1182 (N_1182,N_689,N_337);
nand U1183 (N_1183,N_701,N_104);
nand U1184 (N_1184,N_302,N_427);
xnor U1185 (N_1185,N_417,N_558);
and U1186 (N_1186,N_294,N_488);
nand U1187 (N_1187,N_946,N_824);
and U1188 (N_1188,N_797,N_508);
and U1189 (N_1189,N_58,N_518);
xor U1190 (N_1190,N_958,N_482);
and U1191 (N_1191,N_703,N_832);
nand U1192 (N_1192,N_40,N_468);
nor U1193 (N_1193,N_847,N_228);
xnor U1194 (N_1194,N_675,N_760);
and U1195 (N_1195,N_166,N_376);
and U1196 (N_1196,N_70,N_321);
nor U1197 (N_1197,N_785,N_625);
nor U1198 (N_1198,N_483,N_107);
and U1199 (N_1199,N_279,N_957);
nor U1200 (N_1200,N_861,N_269);
nor U1201 (N_1201,N_829,N_929);
nand U1202 (N_1202,N_806,N_191);
xor U1203 (N_1203,N_520,N_986);
xnor U1204 (N_1204,N_919,N_951);
xnor U1205 (N_1205,N_268,N_906);
nand U1206 (N_1206,N_438,N_491);
nand U1207 (N_1207,N_983,N_371);
nand U1208 (N_1208,N_617,N_201);
nand U1209 (N_1209,N_660,N_284);
and U1210 (N_1210,N_982,N_624);
xor U1211 (N_1211,N_461,N_698);
or U1212 (N_1212,N_170,N_717);
nand U1213 (N_1213,N_405,N_932);
nor U1214 (N_1214,N_307,N_133);
nand U1215 (N_1215,N_26,N_940);
nor U1216 (N_1216,N_79,N_707);
nand U1217 (N_1217,N_140,N_221);
nand U1218 (N_1218,N_691,N_460);
and U1219 (N_1219,N_34,N_127);
and U1220 (N_1220,N_793,N_354);
nand U1221 (N_1221,N_98,N_214);
and U1222 (N_1222,N_742,N_975);
xnor U1223 (N_1223,N_970,N_66);
nor U1224 (N_1224,N_288,N_152);
or U1225 (N_1225,N_679,N_600);
nand U1226 (N_1226,N_490,N_202);
or U1227 (N_1227,N_603,N_877);
nand U1228 (N_1228,N_830,N_565);
or U1229 (N_1229,N_305,N_521);
nor U1230 (N_1230,N_923,N_749);
nand U1231 (N_1231,N_205,N_790);
nand U1232 (N_1232,N_454,N_770);
nand U1233 (N_1233,N_397,N_651);
or U1234 (N_1234,N_539,N_626);
nand U1235 (N_1235,N_734,N_193);
nand U1236 (N_1236,N_407,N_758);
xor U1237 (N_1237,N_999,N_917);
xor U1238 (N_1238,N_56,N_572);
nand U1239 (N_1239,N_233,N_263);
nor U1240 (N_1240,N_159,N_741);
xor U1241 (N_1241,N_927,N_315);
xnor U1242 (N_1242,N_385,N_296);
and U1243 (N_1243,N_497,N_959);
or U1244 (N_1244,N_823,N_678);
nor U1245 (N_1245,N_716,N_731);
or U1246 (N_1246,N_696,N_100);
and U1247 (N_1247,N_894,N_808);
nor U1248 (N_1248,N_969,N_352);
or U1249 (N_1249,N_176,N_242);
or U1250 (N_1250,N_441,N_976);
nand U1251 (N_1251,N_471,N_560);
and U1252 (N_1252,N_481,N_167);
nor U1253 (N_1253,N_465,N_324);
and U1254 (N_1254,N_435,N_196);
and U1255 (N_1255,N_893,N_141);
xnor U1256 (N_1256,N_226,N_247);
xnor U1257 (N_1257,N_459,N_666);
or U1258 (N_1258,N_667,N_646);
nand U1259 (N_1259,N_800,N_755);
nor U1260 (N_1260,N_753,N_496);
xor U1261 (N_1261,N_541,N_884);
and U1262 (N_1262,N_479,N_700);
nand U1263 (N_1263,N_207,N_301);
nor U1264 (N_1264,N_866,N_360);
xnor U1265 (N_1265,N_445,N_534);
and U1266 (N_1266,N_199,N_406);
nand U1267 (N_1267,N_911,N_457);
nor U1268 (N_1268,N_662,N_194);
xor U1269 (N_1269,N_31,N_163);
nand U1270 (N_1270,N_18,N_669);
nand U1271 (N_1271,N_589,N_791);
and U1272 (N_1272,N_72,N_95);
nand U1273 (N_1273,N_277,N_156);
nand U1274 (N_1274,N_304,N_312);
or U1275 (N_1275,N_276,N_325);
or U1276 (N_1276,N_93,N_52);
xor U1277 (N_1277,N_410,N_868);
and U1278 (N_1278,N_448,N_142);
and U1279 (N_1279,N_557,N_381);
and U1280 (N_1280,N_836,N_150);
nor U1281 (N_1281,N_786,N_844);
and U1282 (N_1282,N_470,N_809);
nand U1283 (N_1283,N_44,N_509);
nand U1284 (N_1284,N_299,N_281);
or U1285 (N_1285,N_949,N_293);
xor U1286 (N_1286,N_158,N_122);
nor U1287 (N_1287,N_357,N_178);
nor U1288 (N_1288,N_751,N_746);
nand U1289 (N_1289,N_561,N_799);
nor U1290 (N_1290,N_271,N_629);
nor U1291 (N_1291,N_545,N_869);
nor U1292 (N_1292,N_272,N_813);
nand U1293 (N_1293,N_209,N_974);
or U1294 (N_1294,N_942,N_334);
nor U1295 (N_1295,N_597,N_151);
or U1296 (N_1296,N_953,N_915);
xor U1297 (N_1297,N_637,N_828);
xnor U1298 (N_1298,N_673,N_92);
and U1299 (N_1299,N_174,N_765);
and U1300 (N_1300,N_613,N_519);
xnor U1301 (N_1301,N_720,N_36);
nand U1302 (N_1302,N_74,N_879);
xnor U1303 (N_1303,N_848,N_769);
and U1304 (N_1304,N_160,N_860);
nor U1305 (N_1305,N_559,N_108);
or U1306 (N_1306,N_895,N_888);
or U1307 (N_1307,N_297,N_147);
xnor U1308 (N_1308,N_355,N_346);
nor U1309 (N_1309,N_648,N_562);
nor U1310 (N_1310,N_120,N_530);
xnor U1311 (N_1311,N_954,N_240);
nor U1312 (N_1312,N_499,N_745);
and U1313 (N_1313,N_825,N_409);
nor U1314 (N_1314,N_261,N_230);
nand U1315 (N_1315,N_386,N_632);
or U1316 (N_1316,N_251,N_28);
xnor U1317 (N_1317,N_280,N_99);
nand U1318 (N_1318,N_414,N_721);
and U1319 (N_1319,N_474,N_19);
xor U1320 (N_1320,N_320,N_486);
xnor U1321 (N_1321,N_779,N_295);
and U1322 (N_1322,N_314,N_229);
or U1323 (N_1323,N_153,N_912);
or U1324 (N_1324,N_252,N_783);
xor U1325 (N_1325,N_41,N_955);
or U1326 (N_1326,N_241,N_232);
and U1327 (N_1327,N_439,N_192);
nor U1328 (N_1328,N_4,N_546);
and U1329 (N_1329,N_548,N_607);
xnor U1330 (N_1330,N_817,N_980);
nand U1331 (N_1331,N_370,N_571);
xor U1332 (N_1332,N_789,N_286);
or U1333 (N_1333,N_165,N_724);
nand U1334 (N_1334,N_665,N_582);
and U1335 (N_1335,N_458,N_697);
xor U1336 (N_1336,N_447,N_117);
nand U1337 (N_1337,N_529,N_515);
or U1338 (N_1338,N_111,N_874);
or U1339 (N_1339,N_256,N_55);
nor U1340 (N_1340,N_480,N_933);
xnor U1341 (N_1341,N_585,N_740);
nand U1342 (N_1342,N_116,N_993);
and U1343 (N_1343,N_681,N_48);
nand U1344 (N_1344,N_985,N_215);
or U1345 (N_1345,N_265,N_609);
or U1346 (N_1346,N_618,N_841);
or U1347 (N_1347,N_592,N_455);
nand U1348 (N_1348,N_237,N_692);
nor U1349 (N_1349,N_670,N_189);
nor U1350 (N_1350,N_183,N_506);
xor U1351 (N_1351,N_858,N_563);
xnor U1352 (N_1352,N_909,N_602);
or U1353 (N_1353,N_623,N_867);
nor U1354 (N_1354,N_29,N_245);
and U1355 (N_1355,N_362,N_329);
or U1356 (N_1356,N_155,N_303);
nor U1357 (N_1357,N_462,N_642);
and U1358 (N_1358,N_118,N_730);
or U1359 (N_1359,N_725,N_399);
nand U1360 (N_1360,N_688,N_547);
xnor U1361 (N_1361,N_885,N_595);
nor U1362 (N_1362,N_759,N_126);
nor U1363 (N_1363,N_577,N_363);
or U1364 (N_1364,N_901,N_332);
and U1365 (N_1365,N_8,N_244);
and U1366 (N_1366,N_873,N_327);
nand U1367 (N_1367,N_145,N_981);
or U1368 (N_1368,N_88,N_235);
xor U1369 (N_1369,N_737,N_246);
xor U1370 (N_1370,N_336,N_169);
and U1371 (N_1371,N_39,N_857);
nand U1372 (N_1372,N_78,N_9);
nand U1373 (N_1373,N_146,N_683);
and U1374 (N_1374,N_69,N_259);
or U1375 (N_1375,N_994,N_498);
nor U1376 (N_1376,N_754,N_181);
and U1377 (N_1377,N_114,N_130);
or U1378 (N_1378,N_810,N_289);
nand U1379 (N_1379,N_583,N_930);
nor U1380 (N_1380,N_918,N_896);
nor U1381 (N_1381,N_661,N_446);
and U1382 (N_1382,N_380,N_473);
nand U1383 (N_1383,N_80,N_682);
and U1384 (N_1384,N_654,N_238);
or U1385 (N_1385,N_744,N_309);
or U1386 (N_1386,N_641,N_464);
and U1387 (N_1387,N_516,N_248);
or U1388 (N_1388,N_148,N_382);
nor U1389 (N_1389,N_485,N_659);
nand U1390 (N_1390,N_907,N_671);
xor U1391 (N_1391,N_225,N_510);
nand U1392 (N_1392,N_784,N_726);
nor U1393 (N_1393,N_420,N_132);
nand U1394 (N_1394,N_378,N_511);
nand U1395 (N_1395,N_898,N_0);
nor U1396 (N_1396,N_647,N_880);
or U1397 (N_1397,N_173,N_643);
nor U1398 (N_1398,N_136,N_351);
nor U1399 (N_1399,N_285,N_904);
nand U1400 (N_1400,N_83,N_889);
and U1401 (N_1401,N_856,N_727);
and U1402 (N_1402,N_972,N_776);
and U1403 (N_1403,N_878,N_5);
and U1404 (N_1404,N_492,N_124);
nand U1405 (N_1405,N_121,N_65);
nor U1406 (N_1406,N_403,N_835);
nor U1407 (N_1407,N_137,N_38);
or U1408 (N_1408,N_328,N_622);
nor U1409 (N_1409,N_549,N_796);
xnor U1410 (N_1410,N_805,N_379);
nor U1411 (N_1411,N_578,N_743);
or U1412 (N_1412,N_494,N_634);
and U1413 (N_1413,N_273,N_51);
xnor U1414 (N_1414,N_505,N_290);
nand U1415 (N_1415,N_876,N_81);
or U1416 (N_1416,N_162,N_179);
and U1417 (N_1417,N_575,N_631);
xnor U1418 (N_1418,N_16,N_584);
nor U1419 (N_1419,N_63,N_535);
nor U1420 (N_1420,N_937,N_310);
nor U1421 (N_1421,N_714,N_766);
xnor U1422 (N_1422,N_86,N_495);
nand U1423 (N_1423,N_608,N_477);
nand U1424 (N_1424,N_794,N_694);
or U1425 (N_1425,N_576,N_821);
nand U1426 (N_1426,N_452,N_961);
nand U1427 (N_1427,N_865,N_134);
xor U1428 (N_1428,N_739,N_526);
or U1429 (N_1429,N_685,N_392);
or U1430 (N_1430,N_962,N_875);
xor U1431 (N_1431,N_168,N_905);
nor U1432 (N_1432,N_987,N_881);
xnor U1433 (N_1433,N_947,N_722);
or U1434 (N_1434,N_61,N_2);
nand U1435 (N_1435,N_680,N_313);
nor U1436 (N_1436,N_129,N_658);
nand U1437 (N_1437,N_415,N_655);
nor U1438 (N_1438,N_175,N_713);
nand U1439 (N_1439,N_931,N_85);
nor U1440 (N_1440,N_542,N_212);
and U1441 (N_1441,N_635,N_639);
or U1442 (N_1442,N_339,N_364);
or U1443 (N_1443,N_802,N_512);
nor U1444 (N_1444,N_283,N_53);
nor U1445 (N_1445,N_342,N_239);
nand U1446 (N_1446,N_991,N_977);
nand U1447 (N_1447,N_596,N_444);
or U1448 (N_1448,N_833,N_650);
nand U1449 (N_1449,N_223,N_564);
and U1450 (N_1450,N_428,N_782);
nor U1451 (N_1451,N_425,N_903);
nand U1452 (N_1452,N_204,N_91);
xnor U1453 (N_1453,N_736,N_139);
nand U1454 (N_1454,N_924,N_349);
and U1455 (N_1455,N_14,N_788);
nand U1456 (N_1456,N_451,N_995);
or U1457 (N_1457,N_965,N_275);
or U1458 (N_1458,N_27,N_430);
nor U1459 (N_1459,N_871,N_434);
nand U1460 (N_1460,N_834,N_843);
nor U1461 (N_1461,N_663,N_657);
and U1462 (N_1462,N_287,N_601);
nor U1463 (N_1463,N_883,N_331);
xnor U1464 (N_1464,N_649,N_638);
and U1465 (N_1465,N_818,N_772);
or U1466 (N_1466,N_708,N_733);
and U1467 (N_1467,N_704,N_711);
xnor U1468 (N_1468,N_388,N_763);
and U1469 (N_1469,N_978,N_656);
nand U1470 (N_1470,N_762,N_761);
nand U1471 (N_1471,N_690,N_732);
nand U1472 (N_1472,N_440,N_365);
xnor U1473 (N_1473,N_838,N_729);
or U1474 (N_1474,N_421,N_298);
or U1475 (N_1475,N_47,N_97);
xnor U1476 (N_1476,N_186,N_620);
nand U1477 (N_1477,N_493,N_109);
xor U1478 (N_1478,N_996,N_375);
and U1479 (N_1479,N_433,N_350);
xor U1480 (N_1480,N_684,N_672);
nand U1481 (N_1481,N_948,N_845);
nand U1482 (N_1482,N_674,N_254);
nor U1483 (N_1483,N_330,N_979);
and U1484 (N_1484,N_718,N_853);
xor U1485 (N_1485,N_23,N_149);
and U1486 (N_1486,N_76,N_890);
or U1487 (N_1487,N_426,N_855);
xor U1488 (N_1488,N_258,N_227);
nand U1489 (N_1489,N_775,N_567);
and U1490 (N_1490,N_693,N_573);
and U1491 (N_1491,N_291,N_605);
or U1492 (N_1492,N_748,N_852);
and U1493 (N_1493,N_628,N_581);
xor U1494 (N_1494,N_586,N_943);
xnor U1495 (N_1495,N_182,N_723);
nand U1496 (N_1496,N_234,N_383);
and U1497 (N_1497,N_20,N_316);
nor U1498 (N_1498,N_719,N_377);
or U1499 (N_1499,N_653,N_11);
or U1500 (N_1500,N_614,N_17);
and U1501 (N_1501,N_22,N_540);
nor U1502 (N_1502,N_59,N_71);
nor U1503 (N_1503,N_696,N_205);
xnor U1504 (N_1504,N_569,N_124);
nor U1505 (N_1505,N_673,N_773);
nand U1506 (N_1506,N_341,N_230);
nand U1507 (N_1507,N_700,N_671);
nand U1508 (N_1508,N_305,N_515);
or U1509 (N_1509,N_863,N_907);
or U1510 (N_1510,N_964,N_470);
nor U1511 (N_1511,N_58,N_996);
or U1512 (N_1512,N_15,N_382);
and U1513 (N_1513,N_175,N_344);
nand U1514 (N_1514,N_25,N_730);
or U1515 (N_1515,N_181,N_901);
and U1516 (N_1516,N_749,N_98);
nor U1517 (N_1517,N_705,N_562);
xnor U1518 (N_1518,N_415,N_361);
and U1519 (N_1519,N_34,N_362);
and U1520 (N_1520,N_866,N_746);
xnor U1521 (N_1521,N_74,N_36);
nand U1522 (N_1522,N_328,N_206);
xnor U1523 (N_1523,N_562,N_311);
or U1524 (N_1524,N_724,N_577);
nor U1525 (N_1525,N_769,N_148);
and U1526 (N_1526,N_413,N_179);
and U1527 (N_1527,N_979,N_803);
xnor U1528 (N_1528,N_576,N_248);
nor U1529 (N_1529,N_594,N_619);
xnor U1530 (N_1530,N_502,N_420);
and U1531 (N_1531,N_702,N_30);
and U1532 (N_1532,N_928,N_351);
xnor U1533 (N_1533,N_543,N_479);
nand U1534 (N_1534,N_572,N_81);
nand U1535 (N_1535,N_940,N_927);
or U1536 (N_1536,N_618,N_184);
nand U1537 (N_1537,N_903,N_923);
xnor U1538 (N_1538,N_614,N_442);
and U1539 (N_1539,N_375,N_575);
nor U1540 (N_1540,N_847,N_195);
or U1541 (N_1541,N_195,N_730);
nor U1542 (N_1542,N_413,N_266);
or U1543 (N_1543,N_757,N_97);
nor U1544 (N_1544,N_664,N_953);
or U1545 (N_1545,N_454,N_345);
and U1546 (N_1546,N_327,N_335);
and U1547 (N_1547,N_951,N_717);
or U1548 (N_1548,N_749,N_813);
nor U1549 (N_1549,N_972,N_583);
or U1550 (N_1550,N_156,N_522);
xor U1551 (N_1551,N_260,N_788);
xnor U1552 (N_1552,N_196,N_391);
nand U1553 (N_1553,N_746,N_823);
and U1554 (N_1554,N_701,N_187);
nor U1555 (N_1555,N_842,N_563);
or U1556 (N_1556,N_540,N_741);
xnor U1557 (N_1557,N_243,N_294);
nand U1558 (N_1558,N_749,N_470);
nand U1559 (N_1559,N_105,N_530);
nand U1560 (N_1560,N_26,N_312);
nor U1561 (N_1561,N_467,N_448);
nand U1562 (N_1562,N_444,N_202);
nand U1563 (N_1563,N_764,N_181);
and U1564 (N_1564,N_256,N_692);
xor U1565 (N_1565,N_596,N_506);
nor U1566 (N_1566,N_872,N_359);
and U1567 (N_1567,N_774,N_935);
nor U1568 (N_1568,N_653,N_479);
nand U1569 (N_1569,N_121,N_589);
nand U1570 (N_1570,N_424,N_37);
nand U1571 (N_1571,N_737,N_40);
nand U1572 (N_1572,N_280,N_446);
nor U1573 (N_1573,N_176,N_707);
and U1574 (N_1574,N_462,N_434);
nand U1575 (N_1575,N_50,N_226);
nor U1576 (N_1576,N_622,N_569);
and U1577 (N_1577,N_687,N_383);
or U1578 (N_1578,N_448,N_426);
or U1579 (N_1579,N_418,N_680);
and U1580 (N_1580,N_407,N_213);
and U1581 (N_1581,N_849,N_325);
and U1582 (N_1582,N_111,N_225);
nor U1583 (N_1583,N_908,N_106);
or U1584 (N_1584,N_891,N_89);
nand U1585 (N_1585,N_478,N_935);
nand U1586 (N_1586,N_446,N_637);
and U1587 (N_1587,N_70,N_900);
xor U1588 (N_1588,N_493,N_236);
xnor U1589 (N_1589,N_860,N_466);
xor U1590 (N_1590,N_855,N_519);
nor U1591 (N_1591,N_12,N_838);
and U1592 (N_1592,N_561,N_202);
and U1593 (N_1593,N_235,N_933);
and U1594 (N_1594,N_241,N_136);
and U1595 (N_1595,N_572,N_90);
xor U1596 (N_1596,N_198,N_854);
and U1597 (N_1597,N_231,N_280);
or U1598 (N_1598,N_951,N_784);
or U1599 (N_1599,N_119,N_678);
xnor U1600 (N_1600,N_692,N_975);
nand U1601 (N_1601,N_25,N_685);
and U1602 (N_1602,N_758,N_955);
nor U1603 (N_1603,N_778,N_21);
nor U1604 (N_1604,N_348,N_356);
xor U1605 (N_1605,N_628,N_497);
xnor U1606 (N_1606,N_236,N_337);
or U1607 (N_1607,N_255,N_239);
nor U1608 (N_1608,N_815,N_835);
nor U1609 (N_1609,N_596,N_335);
nor U1610 (N_1610,N_723,N_509);
nand U1611 (N_1611,N_940,N_382);
xnor U1612 (N_1612,N_340,N_872);
xnor U1613 (N_1613,N_791,N_194);
xnor U1614 (N_1614,N_953,N_248);
xnor U1615 (N_1615,N_970,N_435);
xor U1616 (N_1616,N_495,N_813);
or U1617 (N_1617,N_399,N_840);
and U1618 (N_1618,N_4,N_437);
and U1619 (N_1619,N_234,N_224);
or U1620 (N_1620,N_714,N_877);
nand U1621 (N_1621,N_111,N_832);
xnor U1622 (N_1622,N_573,N_571);
nor U1623 (N_1623,N_688,N_689);
xor U1624 (N_1624,N_438,N_735);
or U1625 (N_1625,N_655,N_673);
nor U1626 (N_1626,N_960,N_372);
and U1627 (N_1627,N_379,N_744);
and U1628 (N_1628,N_557,N_637);
nor U1629 (N_1629,N_333,N_443);
and U1630 (N_1630,N_311,N_903);
or U1631 (N_1631,N_614,N_597);
xnor U1632 (N_1632,N_749,N_652);
and U1633 (N_1633,N_810,N_949);
nor U1634 (N_1634,N_458,N_679);
or U1635 (N_1635,N_441,N_162);
nor U1636 (N_1636,N_520,N_219);
nor U1637 (N_1637,N_98,N_74);
nor U1638 (N_1638,N_131,N_512);
nor U1639 (N_1639,N_777,N_330);
or U1640 (N_1640,N_182,N_869);
and U1641 (N_1641,N_937,N_439);
xnor U1642 (N_1642,N_264,N_953);
and U1643 (N_1643,N_374,N_233);
and U1644 (N_1644,N_265,N_780);
nor U1645 (N_1645,N_307,N_739);
nor U1646 (N_1646,N_598,N_486);
or U1647 (N_1647,N_81,N_353);
nand U1648 (N_1648,N_216,N_564);
or U1649 (N_1649,N_653,N_503);
or U1650 (N_1650,N_922,N_6);
or U1651 (N_1651,N_441,N_227);
and U1652 (N_1652,N_127,N_994);
or U1653 (N_1653,N_213,N_169);
nor U1654 (N_1654,N_218,N_605);
nand U1655 (N_1655,N_163,N_437);
or U1656 (N_1656,N_269,N_547);
xor U1657 (N_1657,N_491,N_970);
nand U1658 (N_1658,N_10,N_408);
xor U1659 (N_1659,N_206,N_825);
and U1660 (N_1660,N_473,N_177);
nor U1661 (N_1661,N_509,N_796);
xnor U1662 (N_1662,N_40,N_519);
nor U1663 (N_1663,N_424,N_528);
nor U1664 (N_1664,N_741,N_110);
nor U1665 (N_1665,N_162,N_858);
or U1666 (N_1666,N_60,N_978);
and U1667 (N_1667,N_195,N_193);
nor U1668 (N_1668,N_447,N_692);
and U1669 (N_1669,N_876,N_641);
nor U1670 (N_1670,N_445,N_477);
and U1671 (N_1671,N_636,N_136);
nor U1672 (N_1672,N_392,N_843);
xnor U1673 (N_1673,N_35,N_465);
nand U1674 (N_1674,N_907,N_815);
nand U1675 (N_1675,N_767,N_864);
or U1676 (N_1676,N_883,N_54);
nand U1677 (N_1677,N_603,N_604);
xor U1678 (N_1678,N_842,N_622);
nand U1679 (N_1679,N_179,N_866);
and U1680 (N_1680,N_267,N_922);
xor U1681 (N_1681,N_506,N_980);
nor U1682 (N_1682,N_625,N_918);
and U1683 (N_1683,N_94,N_956);
or U1684 (N_1684,N_542,N_96);
nand U1685 (N_1685,N_419,N_987);
xor U1686 (N_1686,N_542,N_862);
nand U1687 (N_1687,N_7,N_279);
xnor U1688 (N_1688,N_50,N_72);
nand U1689 (N_1689,N_674,N_34);
and U1690 (N_1690,N_270,N_14);
and U1691 (N_1691,N_535,N_234);
xnor U1692 (N_1692,N_540,N_257);
and U1693 (N_1693,N_880,N_78);
or U1694 (N_1694,N_783,N_566);
and U1695 (N_1695,N_717,N_894);
or U1696 (N_1696,N_879,N_532);
or U1697 (N_1697,N_588,N_915);
nor U1698 (N_1698,N_179,N_851);
nand U1699 (N_1699,N_238,N_910);
xor U1700 (N_1700,N_711,N_394);
or U1701 (N_1701,N_517,N_868);
and U1702 (N_1702,N_432,N_340);
nor U1703 (N_1703,N_402,N_562);
nand U1704 (N_1704,N_805,N_415);
or U1705 (N_1705,N_885,N_854);
nor U1706 (N_1706,N_478,N_840);
nand U1707 (N_1707,N_513,N_29);
nor U1708 (N_1708,N_601,N_424);
nand U1709 (N_1709,N_416,N_10);
nor U1710 (N_1710,N_564,N_527);
or U1711 (N_1711,N_778,N_532);
and U1712 (N_1712,N_598,N_288);
nor U1713 (N_1713,N_184,N_993);
xor U1714 (N_1714,N_564,N_569);
nand U1715 (N_1715,N_790,N_340);
or U1716 (N_1716,N_694,N_602);
xnor U1717 (N_1717,N_742,N_330);
nand U1718 (N_1718,N_310,N_700);
nor U1719 (N_1719,N_557,N_32);
or U1720 (N_1720,N_137,N_293);
nor U1721 (N_1721,N_683,N_577);
and U1722 (N_1722,N_620,N_490);
nor U1723 (N_1723,N_428,N_499);
xor U1724 (N_1724,N_519,N_383);
and U1725 (N_1725,N_99,N_138);
xor U1726 (N_1726,N_631,N_684);
and U1727 (N_1727,N_505,N_186);
or U1728 (N_1728,N_950,N_586);
xor U1729 (N_1729,N_171,N_15);
nand U1730 (N_1730,N_833,N_620);
xor U1731 (N_1731,N_756,N_151);
xor U1732 (N_1732,N_397,N_55);
or U1733 (N_1733,N_731,N_423);
nand U1734 (N_1734,N_642,N_539);
or U1735 (N_1735,N_144,N_492);
nor U1736 (N_1736,N_494,N_394);
nor U1737 (N_1737,N_203,N_395);
xor U1738 (N_1738,N_434,N_600);
or U1739 (N_1739,N_411,N_459);
and U1740 (N_1740,N_231,N_72);
xnor U1741 (N_1741,N_244,N_433);
and U1742 (N_1742,N_329,N_840);
or U1743 (N_1743,N_167,N_512);
xor U1744 (N_1744,N_600,N_545);
nor U1745 (N_1745,N_34,N_835);
xnor U1746 (N_1746,N_76,N_0);
or U1747 (N_1747,N_377,N_80);
and U1748 (N_1748,N_76,N_344);
nor U1749 (N_1749,N_614,N_114);
nand U1750 (N_1750,N_984,N_771);
and U1751 (N_1751,N_854,N_981);
nand U1752 (N_1752,N_140,N_250);
and U1753 (N_1753,N_115,N_836);
xnor U1754 (N_1754,N_94,N_493);
nor U1755 (N_1755,N_763,N_997);
or U1756 (N_1756,N_90,N_970);
nor U1757 (N_1757,N_847,N_879);
nor U1758 (N_1758,N_707,N_178);
nor U1759 (N_1759,N_587,N_71);
nand U1760 (N_1760,N_263,N_826);
nor U1761 (N_1761,N_103,N_55);
nand U1762 (N_1762,N_386,N_315);
xor U1763 (N_1763,N_600,N_206);
and U1764 (N_1764,N_294,N_423);
nand U1765 (N_1765,N_445,N_876);
xor U1766 (N_1766,N_25,N_153);
and U1767 (N_1767,N_627,N_863);
or U1768 (N_1768,N_903,N_509);
or U1769 (N_1769,N_693,N_646);
nor U1770 (N_1770,N_935,N_279);
nand U1771 (N_1771,N_771,N_505);
xnor U1772 (N_1772,N_814,N_464);
nor U1773 (N_1773,N_955,N_844);
xor U1774 (N_1774,N_295,N_789);
xor U1775 (N_1775,N_846,N_712);
xnor U1776 (N_1776,N_346,N_402);
or U1777 (N_1777,N_661,N_384);
or U1778 (N_1778,N_16,N_150);
xor U1779 (N_1779,N_136,N_791);
nor U1780 (N_1780,N_114,N_122);
or U1781 (N_1781,N_588,N_147);
and U1782 (N_1782,N_133,N_79);
and U1783 (N_1783,N_72,N_112);
or U1784 (N_1784,N_893,N_258);
and U1785 (N_1785,N_860,N_600);
or U1786 (N_1786,N_356,N_366);
xor U1787 (N_1787,N_879,N_326);
and U1788 (N_1788,N_178,N_526);
nor U1789 (N_1789,N_341,N_316);
nand U1790 (N_1790,N_406,N_547);
nand U1791 (N_1791,N_430,N_777);
xnor U1792 (N_1792,N_538,N_427);
and U1793 (N_1793,N_469,N_317);
nand U1794 (N_1794,N_477,N_259);
xnor U1795 (N_1795,N_712,N_456);
or U1796 (N_1796,N_861,N_920);
or U1797 (N_1797,N_248,N_336);
nand U1798 (N_1798,N_772,N_431);
xnor U1799 (N_1799,N_289,N_398);
nand U1800 (N_1800,N_894,N_771);
xor U1801 (N_1801,N_677,N_604);
or U1802 (N_1802,N_378,N_959);
and U1803 (N_1803,N_35,N_227);
nor U1804 (N_1804,N_856,N_597);
xnor U1805 (N_1805,N_42,N_244);
and U1806 (N_1806,N_141,N_754);
xnor U1807 (N_1807,N_668,N_361);
or U1808 (N_1808,N_918,N_388);
xor U1809 (N_1809,N_375,N_370);
nor U1810 (N_1810,N_305,N_653);
nand U1811 (N_1811,N_25,N_12);
nand U1812 (N_1812,N_896,N_408);
nor U1813 (N_1813,N_588,N_167);
nor U1814 (N_1814,N_242,N_897);
xnor U1815 (N_1815,N_405,N_99);
xor U1816 (N_1816,N_969,N_329);
or U1817 (N_1817,N_906,N_972);
nand U1818 (N_1818,N_479,N_688);
and U1819 (N_1819,N_380,N_431);
nand U1820 (N_1820,N_175,N_867);
nand U1821 (N_1821,N_529,N_266);
and U1822 (N_1822,N_45,N_518);
nor U1823 (N_1823,N_332,N_441);
or U1824 (N_1824,N_176,N_920);
and U1825 (N_1825,N_424,N_109);
xnor U1826 (N_1826,N_634,N_3);
xnor U1827 (N_1827,N_20,N_808);
or U1828 (N_1828,N_679,N_803);
xor U1829 (N_1829,N_628,N_616);
nand U1830 (N_1830,N_132,N_19);
nand U1831 (N_1831,N_975,N_482);
nand U1832 (N_1832,N_519,N_520);
and U1833 (N_1833,N_246,N_987);
xor U1834 (N_1834,N_529,N_597);
nor U1835 (N_1835,N_14,N_948);
nand U1836 (N_1836,N_955,N_748);
or U1837 (N_1837,N_33,N_136);
and U1838 (N_1838,N_483,N_498);
nand U1839 (N_1839,N_358,N_392);
xor U1840 (N_1840,N_108,N_255);
and U1841 (N_1841,N_813,N_589);
xnor U1842 (N_1842,N_986,N_680);
or U1843 (N_1843,N_318,N_85);
and U1844 (N_1844,N_756,N_204);
xor U1845 (N_1845,N_456,N_407);
xor U1846 (N_1846,N_594,N_75);
nand U1847 (N_1847,N_992,N_545);
xnor U1848 (N_1848,N_770,N_917);
nor U1849 (N_1849,N_565,N_430);
nand U1850 (N_1850,N_308,N_389);
nand U1851 (N_1851,N_3,N_169);
nand U1852 (N_1852,N_920,N_530);
nor U1853 (N_1853,N_345,N_271);
nand U1854 (N_1854,N_245,N_799);
or U1855 (N_1855,N_339,N_389);
or U1856 (N_1856,N_253,N_355);
or U1857 (N_1857,N_691,N_604);
or U1858 (N_1858,N_484,N_997);
or U1859 (N_1859,N_363,N_552);
nand U1860 (N_1860,N_383,N_832);
or U1861 (N_1861,N_894,N_19);
xnor U1862 (N_1862,N_765,N_669);
nand U1863 (N_1863,N_460,N_684);
and U1864 (N_1864,N_5,N_952);
nor U1865 (N_1865,N_781,N_341);
or U1866 (N_1866,N_57,N_866);
xor U1867 (N_1867,N_642,N_782);
and U1868 (N_1868,N_311,N_735);
xnor U1869 (N_1869,N_280,N_613);
and U1870 (N_1870,N_139,N_463);
xor U1871 (N_1871,N_602,N_141);
nor U1872 (N_1872,N_542,N_275);
and U1873 (N_1873,N_832,N_914);
xor U1874 (N_1874,N_91,N_944);
or U1875 (N_1875,N_684,N_630);
xor U1876 (N_1876,N_646,N_786);
nor U1877 (N_1877,N_589,N_320);
nand U1878 (N_1878,N_687,N_241);
and U1879 (N_1879,N_911,N_463);
or U1880 (N_1880,N_920,N_914);
or U1881 (N_1881,N_242,N_283);
nand U1882 (N_1882,N_848,N_291);
nand U1883 (N_1883,N_507,N_380);
or U1884 (N_1884,N_570,N_35);
and U1885 (N_1885,N_505,N_246);
nand U1886 (N_1886,N_369,N_869);
nand U1887 (N_1887,N_600,N_927);
or U1888 (N_1888,N_19,N_765);
xnor U1889 (N_1889,N_775,N_299);
nand U1890 (N_1890,N_88,N_313);
and U1891 (N_1891,N_444,N_938);
nand U1892 (N_1892,N_760,N_43);
xnor U1893 (N_1893,N_173,N_849);
and U1894 (N_1894,N_772,N_394);
nor U1895 (N_1895,N_289,N_685);
or U1896 (N_1896,N_260,N_544);
nor U1897 (N_1897,N_444,N_412);
and U1898 (N_1898,N_490,N_501);
nor U1899 (N_1899,N_418,N_262);
nand U1900 (N_1900,N_819,N_647);
or U1901 (N_1901,N_376,N_760);
nand U1902 (N_1902,N_107,N_933);
or U1903 (N_1903,N_941,N_359);
nand U1904 (N_1904,N_800,N_184);
or U1905 (N_1905,N_649,N_480);
nand U1906 (N_1906,N_892,N_390);
and U1907 (N_1907,N_829,N_54);
nand U1908 (N_1908,N_616,N_617);
and U1909 (N_1909,N_524,N_402);
nor U1910 (N_1910,N_158,N_982);
and U1911 (N_1911,N_220,N_108);
nor U1912 (N_1912,N_605,N_679);
nor U1913 (N_1913,N_806,N_236);
xnor U1914 (N_1914,N_200,N_715);
nand U1915 (N_1915,N_482,N_591);
or U1916 (N_1916,N_44,N_388);
and U1917 (N_1917,N_510,N_639);
xor U1918 (N_1918,N_75,N_414);
and U1919 (N_1919,N_728,N_110);
nand U1920 (N_1920,N_388,N_785);
nor U1921 (N_1921,N_184,N_903);
nand U1922 (N_1922,N_451,N_739);
and U1923 (N_1923,N_75,N_86);
and U1924 (N_1924,N_564,N_195);
xor U1925 (N_1925,N_565,N_239);
or U1926 (N_1926,N_99,N_31);
nand U1927 (N_1927,N_993,N_891);
and U1928 (N_1928,N_666,N_365);
nand U1929 (N_1929,N_19,N_997);
or U1930 (N_1930,N_591,N_334);
nor U1931 (N_1931,N_558,N_221);
xor U1932 (N_1932,N_10,N_977);
or U1933 (N_1933,N_955,N_848);
nand U1934 (N_1934,N_48,N_22);
or U1935 (N_1935,N_148,N_653);
and U1936 (N_1936,N_202,N_379);
and U1937 (N_1937,N_283,N_700);
or U1938 (N_1938,N_354,N_463);
nand U1939 (N_1939,N_278,N_916);
nor U1940 (N_1940,N_176,N_605);
nor U1941 (N_1941,N_961,N_823);
nor U1942 (N_1942,N_79,N_306);
nor U1943 (N_1943,N_790,N_828);
nor U1944 (N_1944,N_562,N_581);
or U1945 (N_1945,N_60,N_466);
and U1946 (N_1946,N_170,N_431);
or U1947 (N_1947,N_329,N_100);
xnor U1948 (N_1948,N_97,N_487);
xnor U1949 (N_1949,N_617,N_991);
xnor U1950 (N_1950,N_766,N_259);
nor U1951 (N_1951,N_290,N_937);
or U1952 (N_1952,N_488,N_287);
xnor U1953 (N_1953,N_155,N_602);
and U1954 (N_1954,N_808,N_348);
nand U1955 (N_1955,N_459,N_481);
or U1956 (N_1956,N_572,N_250);
nor U1957 (N_1957,N_415,N_875);
nor U1958 (N_1958,N_939,N_82);
and U1959 (N_1959,N_906,N_195);
or U1960 (N_1960,N_855,N_823);
nor U1961 (N_1961,N_776,N_997);
xor U1962 (N_1962,N_63,N_811);
and U1963 (N_1963,N_796,N_249);
or U1964 (N_1964,N_35,N_3);
or U1965 (N_1965,N_521,N_97);
xnor U1966 (N_1966,N_441,N_286);
and U1967 (N_1967,N_566,N_956);
and U1968 (N_1968,N_109,N_895);
or U1969 (N_1969,N_733,N_664);
and U1970 (N_1970,N_144,N_217);
nor U1971 (N_1971,N_506,N_311);
and U1972 (N_1972,N_866,N_600);
xor U1973 (N_1973,N_247,N_745);
or U1974 (N_1974,N_869,N_526);
xnor U1975 (N_1975,N_898,N_507);
and U1976 (N_1976,N_142,N_306);
or U1977 (N_1977,N_283,N_307);
nand U1978 (N_1978,N_268,N_511);
and U1979 (N_1979,N_59,N_913);
nor U1980 (N_1980,N_352,N_889);
xnor U1981 (N_1981,N_26,N_689);
nor U1982 (N_1982,N_877,N_821);
or U1983 (N_1983,N_230,N_431);
or U1984 (N_1984,N_924,N_899);
or U1985 (N_1985,N_855,N_605);
or U1986 (N_1986,N_289,N_435);
nand U1987 (N_1987,N_741,N_845);
and U1988 (N_1988,N_993,N_438);
nand U1989 (N_1989,N_180,N_928);
and U1990 (N_1990,N_321,N_999);
nand U1991 (N_1991,N_979,N_925);
nor U1992 (N_1992,N_482,N_903);
or U1993 (N_1993,N_758,N_603);
xnor U1994 (N_1994,N_322,N_15);
nand U1995 (N_1995,N_325,N_967);
nand U1996 (N_1996,N_374,N_894);
and U1997 (N_1997,N_782,N_870);
or U1998 (N_1998,N_718,N_30);
xnor U1999 (N_1999,N_57,N_614);
xor U2000 (N_2000,N_1499,N_1278);
xor U2001 (N_2001,N_1395,N_1429);
nand U2002 (N_2002,N_1461,N_1952);
xor U2003 (N_2003,N_1249,N_1557);
nand U2004 (N_2004,N_1166,N_1611);
or U2005 (N_2005,N_1162,N_1860);
or U2006 (N_2006,N_1801,N_1511);
nand U2007 (N_2007,N_1772,N_1531);
nand U2008 (N_2008,N_1583,N_1233);
xnor U2009 (N_2009,N_1354,N_1389);
and U2010 (N_2010,N_1115,N_1375);
and U2011 (N_2011,N_1972,N_1175);
nand U2012 (N_2012,N_1623,N_1417);
or U2013 (N_2013,N_1776,N_1255);
and U2014 (N_2014,N_1290,N_1157);
nor U2015 (N_2015,N_1271,N_1446);
xnor U2016 (N_2016,N_1096,N_1041);
nor U2017 (N_2017,N_1247,N_1535);
nand U2018 (N_2018,N_1288,N_1027);
or U2019 (N_2019,N_1785,N_1879);
nand U2020 (N_2020,N_1664,N_1077);
xor U2021 (N_2021,N_1450,N_1010);
or U2022 (N_2022,N_1198,N_1242);
and U2023 (N_2023,N_1858,N_1745);
xor U2024 (N_2024,N_1241,N_1159);
nor U2025 (N_2025,N_1413,N_1128);
xor U2026 (N_2026,N_1209,N_1831);
and U2027 (N_2027,N_1964,N_1773);
and U2028 (N_2028,N_1980,N_1550);
or U2029 (N_2029,N_1385,N_1713);
nand U2030 (N_2030,N_1055,N_1030);
nor U2031 (N_2031,N_1747,N_1421);
or U2032 (N_2032,N_1236,N_1903);
and U2033 (N_2033,N_1709,N_1377);
xnor U2034 (N_2034,N_1830,N_1070);
and U2035 (N_2035,N_1280,N_1599);
and U2036 (N_2036,N_1138,N_1983);
xnor U2037 (N_2037,N_1533,N_1305);
xor U2038 (N_2038,N_1558,N_1348);
nor U2039 (N_2039,N_1434,N_1496);
nand U2040 (N_2040,N_1107,N_1135);
nand U2041 (N_2041,N_1390,N_1338);
nor U2042 (N_2042,N_1037,N_1799);
nand U2043 (N_2043,N_1451,N_1267);
nor U2044 (N_2044,N_1941,N_1444);
nand U2045 (N_2045,N_1582,N_1396);
and U2046 (N_2046,N_1838,N_1775);
xor U2047 (N_2047,N_1925,N_1362);
or U2048 (N_2048,N_1105,N_1475);
or U2049 (N_2049,N_1503,N_1594);
and U2050 (N_2050,N_1464,N_1373);
nand U2051 (N_2051,N_1784,N_1516);
and U2052 (N_2052,N_1662,N_1192);
xnor U2053 (N_2053,N_1562,N_1724);
nor U2054 (N_2054,N_1978,N_1920);
xor U2055 (N_2055,N_1976,N_1645);
nand U2056 (N_2056,N_1191,N_1315);
nand U2057 (N_2057,N_1102,N_1302);
and U2058 (N_2058,N_1552,N_1600);
nor U2059 (N_2059,N_1842,N_1203);
xor U2060 (N_2060,N_1639,N_1561);
or U2061 (N_2061,N_1497,N_1462);
xnor U2062 (N_2062,N_1569,N_1722);
and U2063 (N_2063,N_1670,N_1289);
nor U2064 (N_2064,N_1851,N_1335);
nor U2065 (N_2065,N_1098,N_1194);
xor U2066 (N_2066,N_1666,N_1769);
xnor U2067 (N_2067,N_1577,N_1548);
and U2068 (N_2068,N_1627,N_1796);
nor U2069 (N_2069,N_1628,N_1788);
xnor U2070 (N_2070,N_1509,N_1843);
or U2071 (N_2071,N_1877,N_1384);
or U2072 (N_2072,N_1572,N_1766);
nand U2073 (N_2073,N_1119,N_1146);
and U2074 (N_2074,N_1728,N_1261);
xor U2075 (N_2075,N_1597,N_1716);
nand U2076 (N_2076,N_1401,N_1609);
xnor U2077 (N_2077,N_1833,N_1500);
and U2078 (N_2078,N_1221,N_1381);
and U2079 (N_2079,N_1235,N_1519);
xnor U2080 (N_2080,N_1132,N_1306);
xor U2081 (N_2081,N_1379,N_1588);
nand U2082 (N_2082,N_1074,N_1479);
or U2083 (N_2083,N_1440,N_1590);
nor U2084 (N_2084,N_1602,N_1770);
or U2085 (N_2085,N_1215,N_1977);
nor U2086 (N_2086,N_1647,N_1488);
nor U2087 (N_2087,N_1303,N_1892);
nand U2088 (N_2088,N_1011,N_1510);
and U2089 (N_2089,N_1369,N_1167);
nand U2090 (N_2090,N_1739,N_1878);
nand U2091 (N_2091,N_1922,N_1699);
and U2092 (N_2092,N_1176,N_1953);
or U2093 (N_2093,N_1126,N_1622);
and U2094 (N_2094,N_1603,N_1678);
xor U2095 (N_2095,N_1629,N_1934);
xnor U2096 (N_2096,N_1484,N_1002);
xor U2097 (N_2097,N_1090,N_1383);
or U2098 (N_2098,N_1145,N_1353);
nand U2099 (N_2099,N_1813,N_1436);
or U2100 (N_2100,N_1542,N_1994);
nor U2101 (N_2101,N_1341,N_1615);
and U2102 (N_2102,N_1553,N_1610);
nor U2103 (N_2103,N_1168,N_1259);
or U2104 (N_2104,N_1575,N_1836);
xor U2105 (N_2105,N_1131,N_1940);
xor U2106 (N_2106,N_1642,N_1887);
xnor U2107 (N_2107,N_1640,N_1874);
and U2108 (N_2108,N_1149,N_1756);
or U2109 (N_2109,N_1201,N_1616);
and U2110 (N_2110,N_1698,N_1026);
and U2111 (N_2111,N_1673,N_1021);
or U2112 (N_2112,N_1815,N_1680);
or U2113 (N_2113,N_1153,N_1792);
nor U2114 (N_2114,N_1189,N_1706);
and U2115 (N_2115,N_1365,N_1826);
and U2116 (N_2116,N_1525,N_1586);
nand U2117 (N_2117,N_1942,N_1276);
and U2118 (N_2118,N_1015,N_1309);
nor U2119 (N_2119,N_1791,N_1214);
xnor U2120 (N_2120,N_1950,N_1998);
xnor U2121 (N_2121,N_1927,N_1202);
xor U2122 (N_2122,N_1867,N_1483);
and U2123 (N_2123,N_1472,N_1322);
and U2124 (N_2124,N_1493,N_1841);
and U2125 (N_2125,N_1546,N_1900);
xnor U2126 (N_2126,N_1974,N_1334);
nand U2127 (N_2127,N_1891,N_1559);
or U2128 (N_2128,N_1489,N_1237);
and U2129 (N_2129,N_1823,N_1344);
xnor U2130 (N_2130,N_1258,N_1697);
xor U2131 (N_2131,N_1343,N_1094);
nor U2132 (N_2132,N_1283,N_1832);
nand U2133 (N_2133,N_1857,N_1393);
or U2134 (N_2134,N_1106,N_1693);
and U2135 (N_2135,N_1257,N_1056);
and U2136 (N_2136,N_1243,N_1150);
or U2137 (N_2137,N_1431,N_1391);
or U2138 (N_2138,N_1337,N_1207);
and U2139 (N_2139,N_1671,N_1733);
nor U2140 (N_2140,N_1862,N_1284);
xnor U2141 (N_2141,N_1545,N_1859);
nor U2142 (N_2142,N_1076,N_1804);
and U2143 (N_2143,N_1232,N_1460);
or U2144 (N_2144,N_1151,N_1211);
and U2145 (N_2145,N_1287,N_1342);
and U2146 (N_2146,N_1144,N_1817);
and U2147 (N_2147,N_1574,N_1311);
nor U2148 (N_2148,N_1755,N_1449);
nor U2149 (N_2149,N_1441,N_1178);
nand U2150 (N_2150,N_1522,N_1478);
and U2151 (N_2151,N_1031,N_1795);
and U2152 (N_2152,N_1184,N_1154);
or U2153 (N_2153,N_1644,N_1665);
nor U2154 (N_2154,N_1125,N_1789);
xnor U2155 (N_2155,N_1040,N_1187);
and U2156 (N_2156,N_1883,N_1465);
and U2157 (N_2157,N_1683,N_1660);
xnor U2158 (N_2158,N_1081,N_1814);
nor U2159 (N_2159,N_1414,N_1181);
xor U2160 (N_2160,N_1643,N_1825);
nor U2161 (N_2161,N_1452,N_1293);
or U2162 (N_2162,N_1244,N_1212);
and U2163 (N_2163,N_1620,N_1116);
or U2164 (N_2164,N_1428,N_1112);
and U2165 (N_2165,N_1649,N_1996);
nand U2166 (N_2166,N_1477,N_1560);
nand U2167 (N_2167,N_1505,N_1346);
and U2168 (N_2168,N_1173,N_1058);
xnor U2169 (N_2169,N_1955,N_1938);
or U2170 (N_2170,N_1073,N_1871);
or U2171 (N_2171,N_1592,N_1371);
nand U2172 (N_2172,N_1818,N_1845);
xnor U2173 (N_2173,N_1480,N_1459);
xnor U2174 (N_2174,N_1069,N_1193);
or U2175 (N_2175,N_1219,N_1973);
nor U2176 (N_2176,N_1866,N_1689);
xor U2177 (N_2177,N_1811,N_1494);
or U2178 (N_2178,N_1091,N_1439);
xor U2179 (N_2179,N_1888,N_1238);
xnor U2180 (N_2180,N_1536,N_1279);
nor U2181 (N_2181,N_1540,N_1367);
nand U2182 (N_2182,N_1884,N_1918);
xnor U2183 (N_2183,N_1024,N_1797);
xnor U2184 (N_2184,N_1712,N_1741);
nand U2185 (N_2185,N_1708,N_1963);
nor U2186 (N_2186,N_1266,N_1448);
nand U2187 (N_2187,N_1675,N_1876);
xnor U2188 (N_2188,N_1677,N_1003);
nor U2189 (N_2189,N_1001,N_1298);
or U2190 (N_2190,N_1299,N_1374);
nor U2191 (N_2191,N_1382,N_1913);
xnor U2192 (N_2192,N_1812,N_1632);
xor U2193 (N_2193,N_1358,N_1029);
and U2194 (N_2194,N_1598,N_1607);
nor U2195 (N_2195,N_1435,N_1250);
and U2196 (N_2196,N_1409,N_1226);
or U2197 (N_2197,N_1171,N_1679);
or U2198 (N_2198,N_1196,N_1174);
nor U2199 (N_2199,N_1840,N_1805);
nor U2200 (N_2200,N_1028,N_1372);
and U2201 (N_2201,N_1111,N_1412);
xnor U2202 (N_2202,N_1667,N_1966);
or U2203 (N_2203,N_1361,N_1835);
xor U2204 (N_2204,N_1433,N_1160);
nor U2205 (N_2205,N_1053,N_1947);
nor U2206 (N_2206,N_1430,N_1397);
nor U2207 (N_2207,N_1803,N_1039);
and U2208 (N_2208,N_1437,N_1084);
nand U2209 (N_2209,N_1406,N_1944);
or U2210 (N_2210,N_1317,N_1723);
xor U2211 (N_2211,N_1177,N_1291);
or U2212 (N_2212,N_1961,N_1861);
nand U2213 (N_2213,N_1188,N_1839);
and U2214 (N_2214,N_1061,N_1099);
nand U2215 (N_2215,N_1340,N_1764);
nand U2216 (N_2216,N_1227,N_1929);
or U2217 (N_2217,N_1988,N_1721);
or U2218 (N_2218,N_1333,N_1601);
nand U2219 (N_2219,N_1345,N_1968);
nor U2220 (N_2220,N_1200,N_1727);
nand U2221 (N_2221,N_1245,N_1685);
nor U2222 (N_2222,N_1323,N_1325);
and U2223 (N_2223,N_1914,N_1587);
nand U2224 (N_2224,N_1515,N_1272);
xnor U2225 (N_2225,N_1148,N_1425);
or U2226 (N_2226,N_1718,N_1674);
nand U2227 (N_2227,N_1619,N_1652);
xor U2228 (N_2228,N_1204,N_1329);
nor U2229 (N_2229,N_1183,N_1682);
xor U2230 (N_2230,N_1130,N_1658);
nand U2231 (N_2231,N_1103,N_1777);
xor U2232 (N_2232,N_1447,N_1498);
nand U2233 (N_2233,N_1270,N_1370);
or U2234 (N_2234,N_1705,N_1532);
nand U2235 (N_2235,N_1294,N_1239);
nand U2236 (N_2236,N_1692,N_1765);
xnor U2237 (N_2237,N_1962,N_1100);
or U2238 (N_2238,N_1012,N_1471);
nor U2239 (N_2239,N_1045,N_1134);
or U2240 (N_2240,N_1411,N_1710);
xor U2241 (N_2241,N_1514,N_1386);
and U2242 (N_2242,N_1538,N_1418);
xnor U2243 (N_2243,N_1419,N_1916);
nor U2244 (N_2244,N_1736,N_1093);
nor U2245 (N_2245,N_1400,N_1919);
nor U2246 (N_2246,N_1806,N_1704);
xor U2247 (N_2247,N_1956,N_1407);
nor U2248 (N_2248,N_1800,N_1019);
nor U2249 (N_2249,N_1984,N_1265);
xor U2250 (N_2250,N_1101,N_1108);
and U2251 (N_2251,N_1332,N_1368);
xnor U2252 (N_2252,N_1117,N_1256);
or U2253 (N_2253,N_1468,N_1218);
or U2254 (N_2254,N_1864,N_1886);
nor U2255 (N_2255,N_1199,N_1473);
or U2256 (N_2256,N_1481,N_1376);
or U2257 (N_2257,N_1424,N_1197);
or U2258 (N_2258,N_1732,N_1633);
and U2259 (N_2259,N_1565,N_1681);
xor U2260 (N_2260,N_1992,N_1097);
nor U2261 (N_2261,N_1408,N_1520);
xor U2262 (N_2262,N_1646,N_1895);
and U2263 (N_2263,N_1771,N_1206);
or U2264 (N_2264,N_1230,N_1926);
or U2265 (N_2265,N_1458,N_1120);
or U2266 (N_2266,N_1985,N_1141);
nor U2267 (N_2267,N_1047,N_1513);
and U2268 (N_2268,N_1790,N_1224);
and U2269 (N_2269,N_1834,N_1454);
or U2270 (N_2270,N_1273,N_1139);
and U2271 (N_2271,N_1474,N_1222);
nor U2272 (N_2272,N_1737,N_1210);
and U2273 (N_2273,N_1630,N_1025);
and U2274 (N_2274,N_1281,N_1443);
nor U2275 (N_2275,N_1626,N_1634);
nand U2276 (N_2276,N_1808,N_1277);
or U2277 (N_2277,N_1608,N_1856);
and U2278 (N_2278,N_1528,N_1969);
nand U2279 (N_2279,N_1750,N_1264);
and U2280 (N_2280,N_1008,N_1006);
xnor U2281 (N_2281,N_1051,N_1023);
nand U2282 (N_2282,N_1742,N_1182);
nand U2283 (N_2283,N_1578,N_1110);
xnor U2284 (N_2284,N_1912,N_1999);
or U2285 (N_2285,N_1663,N_1223);
xor U2286 (N_2286,N_1286,N_1898);
xnor U2287 (N_2287,N_1085,N_1229);
nor U2288 (N_2288,N_1216,N_1981);
or U2289 (N_2289,N_1180,N_1989);
xor U2290 (N_2290,N_1780,N_1951);
nand U2291 (N_2291,N_1863,N_1032);
and U2292 (N_2292,N_1476,N_1970);
nand U2293 (N_2293,N_1924,N_1336);
xor U2294 (N_2294,N_1915,N_1676);
or U2295 (N_2295,N_1104,N_1517);
or U2296 (N_2296,N_1339,N_1547);
nand U2297 (N_2297,N_1521,N_1868);
nor U2298 (N_2298,N_1364,N_1827);
nand U2299 (N_2299,N_1469,N_1059);
or U2300 (N_2300,N_1136,N_1072);
and U2301 (N_2301,N_1979,N_1802);
xor U2302 (N_2302,N_1725,N_1591);
or U2303 (N_2303,N_1958,N_1275);
nand U2304 (N_2304,N_1568,N_1930);
nand U2305 (N_2305,N_1759,N_1809);
and U2306 (N_2306,N_1967,N_1416);
nand U2307 (N_2307,N_1388,N_1088);
nand U2308 (N_2308,N_1965,N_1762);
nor U2309 (N_2309,N_1000,N_1993);
or U2310 (N_2310,N_1301,N_1080);
xnor U2311 (N_2311,N_1621,N_1684);
xnor U2312 (N_2312,N_1618,N_1847);
nor U2313 (N_2313,N_1351,N_1043);
and U2314 (N_2314,N_1405,N_1314);
xor U2315 (N_2315,N_1086,N_1313);
xor U2316 (N_2316,N_1321,N_1075);
xor U2317 (N_2317,N_1359,N_1512);
and U2318 (N_2318,N_1318,N_1566);
or U2319 (N_2319,N_1089,N_1829);
nor U2320 (N_2320,N_1767,N_1567);
and U2321 (N_2321,N_1997,N_1579);
and U2322 (N_2322,N_1638,N_1885);
and U2323 (N_2323,N_1046,N_1004);
or U2324 (N_2324,N_1897,N_1822);
xnor U2325 (N_2325,N_1923,N_1902);
nor U2326 (N_2326,N_1690,N_1543);
nor U2327 (N_2327,N_1324,N_1357);
or U2328 (N_2328,N_1606,N_1544);
nand U2329 (N_2329,N_1508,N_1873);
nor U2330 (N_2330,N_1456,N_1534);
nor U2331 (N_2331,N_1016,N_1754);
or U2332 (N_2332,N_1636,N_1155);
nor U2333 (N_2333,N_1524,N_1482);
nand U2334 (N_2334,N_1415,N_1635);
nor U2335 (N_2335,N_1890,N_1501);
nand U2336 (N_2336,N_1641,N_1172);
nand U2337 (N_2337,N_1399,N_1231);
or U2338 (N_2338,N_1703,N_1758);
nor U2339 (N_2339,N_1893,N_1328);
nand U2340 (N_2340,N_1975,N_1783);
or U2341 (N_2341,N_1297,N_1463);
xor U2342 (N_2342,N_1453,N_1714);
nor U2343 (N_2343,N_1398,N_1848);
and U2344 (N_2344,N_1687,N_1855);
nand U2345 (N_2345,N_1786,N_1854);
and U2346 (N_2346,N_1604,N_1052);
and U2347 (N_2347,N_1778,N_1147);
or U2348 (N_2348,N_1048,N_1467);
and U2349 (N_2349,N_1164,N_1905);
xnor U2350 (N_2350,N_1695,N_1217);
and U2351 (N_2351,N_1816,N_1190);
nand U2352 (N_2352,N_1349,N_1220);
nor U2353 (N_2353,N_1571,N_1949);
nand U2354 (N_2354,N_1140,N_1865);
nor U2355 (N_2355,N_1360,N_1248);
or U2356 (N_2356,N_1828,N_1083);
nor U2357 (N_2357,N_1113,N_1987);
xor U2358 (N_2358,N_1121,N_1960);
nor U2359 (N_2359,N_1054,N_1819);
xnor U2360 (N_2360,N_1022,N_1761);
or U2361 (N_2361,N_1637,N_1700);
and U2362 (N_2362,N_1504,N_1327);
nand U2363 (N_2363,N_1347,N_1779);
nand U2364 (N_2364,N_1928,N_1551);
and U2365 (N_2365,N_1143,N_1404);
nand U2366 (N_2366,N_1352,N_1161);
and U2367 (N_2367,N_1486,N_1487);
nor U2368 (N_2368,N_1751,N_1654);
xor U2369 (N_2369,N_1844,N_1793);
nor U2370 (N_2370,N_1529,N_1485);
xnor U2371 (N_2371,N_1807,N_1720);
or U2372 (N_2372,N_1445,N_1837);
xor U2373 (N_2373,N_1881,N_1526);
or U2374 (N_2374,N_1044,N_1875);
and U2375 (N_2375,N_1007,N_1730);
or U2376 (N_2376,N_1078,N_1282);
and U2377 (N_2377,N_1020,N_1087);
xor U2378 (N_2378,N_1186,N_1423);
nand U2379 (N_2379,N_1537,N_1296);
xnor U2380 (N_2380,N_1991,N_1506);
nand U2381 (N_2381,N_1648,N_1995);
and U2382 (N_2382,N_1410,N_1071);
nand U2383 (N_2383,N_1403,N_1959);
and U2384 (N_2384,N_1906,N_1554);
or U2385 (N_2385,N_1907,N_1331);
nor U2386 (N_2386,N_1208,N_1035);
nor U2387 (N_2387,N_1909,N_1749);
nand U2388 (N_2388,N_1669,N_1285);
nand U2389 (N_2389,N_1225,N_1179);
nor U2390 (N_2390,N_1185,N_1904);
or U2391 (N_2391,N_1355,N_1853);
or U2392 (N_2392,N_1326,N_1613);
nor U2393 (N_2393,N_1810,N_1631);
nand U2394 (N_2394,N_1300,N_1165);
or U2395 (N_2395,N_1363,N_1316);
nor U2396 (N_2396,N_1492,N_1917);
nor U2397 (N_2397,N_1240,N_1570);
xnor U2398 (N_2398,N_1158,N_1872);
nor U2399 (N_2399,N_1065,N_1009);
nand U2400 (N_2400,N_1014,N_1308);
and U2401 (N_2401,N_1757,N_1005);
xor U2402 (N_2402,N_1114,N_1580);
nor U2403 (N_2403,N_1653,N_1251);
nor U2404 (N_2404,N_1614,N_1049);
nand U2405 (N_2405,N_1262,N_1067);
nand U2406 (N_2406,N_1549,N_1668);
and U2407 (N_2407,N_1123,N_1911);
or U2408 (N_2408,N_1584,N_1596);
xor U2409 (N_2409,N_1254,N_1118);
or U2410 (N_2410,N_1034,N_1731);
nand U2411 (N_2411,N_1882,N_1782);
nand U2412 (N_2412,N_1387,N_1711);
nand U2413 (N_2413,N_1932,N_1744);
nand U2414 (N_2414,N_1899,N_1939);
or U2415 (N_2415,N_1013,N_1696);
xnor U2416 (N_2416,N_1846,N_1470);
and U2417 (N_2417,N_1948,N_1438);
nor U2418 (N_2418,N_1901,N_1760);
or U2419 (N_2419,N_1931,N_1060);
xor U2420 (N_2420,N_1142,N_1295);
or U2421 (N_2421,N_1908,N_1707);
or U2422 (N_2422,N_1933,N_1936);
or U2423 (N_2423,N_1523,N_1935);
nor U2424 (N_2424,N_1982,N_1057);
nand U2425 (N_2425,N_1869,N_1394);
nand U2426 (N_2426,N_1079,N_1957);
xnor U2427 (N_2427,N_1442,N_1420);
nor U2428 (N_2428,N_1320,N_1378);
or U2429 (N_2429,N_1743,N_1686);
nor U2430 (N_2430,N_1539,N_1850);
and U2431 (N_2431,N_1870,N_1124);
nand U2432 (N_2432,N_1849,N_1457);
xor U2433 (N_2433,N_1205,N_1556);
nand U2434 (N_2434,N_1986,N_1921);
nor U2435 (N_2435,N_1246,N_1292);
and U2436 (N_2436,N_1050,N_1495);
xnor U2437 (N_2437,N_1426,N_1127);
nand U2438 (N_2438,N_1129,N_1954);
and U2439 (N_2439,N_1527,N_1319);
nor U2440 (N_2440,N_1530,N_1774);
and U2441 (N_2441,N_1234,N_1109);
and U2442 (N_2442,N_1787,N_1068);
or U2443 (N_2443,N_1133,N_1502);
xnor U2444 (N_2444,N_1170,N_1794);
or U2445 (N_2445,N_1651,N_1573);
and U2446 (N_2446,N_1702,N_1064);
or U2447 (N_2447,N_1672,N_1253);
and U2448 (N_2448,N_1274,N_1466);
and U2449 (N_2449,N_1563,N_1455);
xor U2450 (N_2450,N_1095,N_1945);
or U2451 (N_2451,N_1585,N_1392);
nor U2452 (N_2452,N_1852,N_1748);
or U2453 (N_2453,N_1092,N_1330);
or U2454 (N_2454,N_1661,N_1726);
nor U2455 (N_2455,N_1033,N_1380);
or U2456 (N_2456,N_1688,N_1307);
nor U2457 (N_2457,N_1659,N_1541);
or U2458 (N_2458,N_1402,N_1937);
or U2459 (N_2459,N_1729,N_1213);
nand U2460 (N_2460,N_1719,N_1593);
or U2461 (N_2461,N_1734,N_1304);
nand U2462 (N_2462,N_1889,N_1946);
and U2463 (N_2463,N_1657,N_1971);
and U2464 (N_2464,N_1625,N_1612);
xnor U2465 (N_2465,N_1312,N_1605);
and U2466 (N_2466,N_1763,N_1735);
or U2467 (N_2467,N_1507,N_1701);
nor U2468 (N_2468,N_1310,N_1356);
and U2469 (N_2469,N_1894,N_1752);
xnor U2470 (N_2470,N_1062,N_1715);
nor U2471 (N_2471,N_1263,N_1195);
xor U2472 (N_2472,N_1581,N_1268);
nor U2473 (N_2473,N_1821,N_1066);
nor U2474 (N_2474,N_1156,N_1163);
nand U2475 (N_2475,N_1617,N_1017);
and U2476 (N_2476,N_1595,N_1824);
nor U2477 (N_2477,N_1422,N_1650);
nor U2478 (N_2478,N_1820,N_1152);
and U2479 (N_2479,N_1082,N_1880);
and U2480 (N_2480,N_1655,N_1691);
nor U2481 (N_2481,N_1491,N_1228);
and U2482 (N_2482,N_1555,N_1350);
xor U2483 (N_2483,N_1122,N_1260);
nand U2484 (N_2484,N_1589,N_1943);
or U2485 (N_2485,N_1564,N_1717);
or U2486 (N_2486,N_1694,N_1740);
nand U2487 (N_2487,N_1518,N_1896);
and U2488 (N_2488,N_1366,N_1432);
nand U2489 (N_2489,N_1624,N_1018);
nor U2490 (N_2490,N_1738,N_1576);
nand U2491 (N_2491,N_1063,N_1746);
and U2492 (N_2492,N_1910,N_1252);
and U2493 (N_2493,N_1038,N_1990);
nor U2494 (N_2494,N_1753,N_1781);
nand U2495 (N_2495,N_1169,N_1490);
nor U2496 (N_2496,N_1656,N_1768);
or U2497 (N_2497,N_1427,N_1042);
nand U2498 (N_2498,N_1798,N_1269);
and U2499 (N_2499,N_1137,N_1036);
nand U2500 (N_2500,N_1812,N_1005);
nor U2501 (N_2501,N_1535,N_1081);
or U2502 (N_2502,N_1691,N_1248);
nor U2503 (N_2503,N_1467,N_1739);
xnor U2504 (N_2504,N_1976,N_1826);
xnor U2505 (N_2505,N_1226,N_1768);
and U2506 (N_2506,N_1081,N_1095);
and U2507 (N_2507,N_1365,N_1395);
and U2508 (N_2508,N_1077,N_1224);
nand U2509 (N_2509,N_1886,N_1990);
and U2510 (N_2510,N_1606,N_1133);
or U2511 (N_2511,N_1848,N_1101);
xor U2512 (N_2512,N_1267,N_1562);
nor U2513 (N_2513,N_1897,N_1798);
xnor U2514 (N_2514,N_1506,N_1004);
or U2515 (N_2515,N_1949,N_1133);
and U2516 (N_2516,N_1249,N_1562);
nor U2517 (N_2517,N_1962,N_1982);
nand U2518 (N_2518,N_1432,N_1695);
nand U2519 (N_2519,N_1870,N_1612);
and U2520 (N_2520,N_1141,N_1432);
xor U2521 (N_2521,N_1825,N_1100);
or U2522 (N_2522,N_1565,N_1279);
xnor U2523 (N_2523,N_1437,N_1803);
xor U2524 (N_2524,N_1048,N_1738);
or U2525 (N_2525,N_1675,N_1307);
and U2526 (N_2526,N_1293,N_1673);
nor U2527 (N_2527,N_1459,N_1240);
nor U2528 (N_2528,N_1140,N_1721);
nor U2529 (N_2529,N_1264,N_1065);
nor U2530 (N_2530,N_1196,N_1428);
nand U2531 (N_2531,N_1851,N_1119);
or U2532 (N_2532,N_1386,N_1104);
or U2533 (N_2533,N_1982,N_1223);
and U2534 (N_2534,N_1652,N_1426);
or U2535 (N_2535,N_1681,N_1745);
or U2536 (N_2536,N_1588,N_1820);
nor U2537 (N_2537,N_1494,N_1250);
nor U2538 (N_2538,N_1865,N_1196);
nand U2539 (N_2539,N_1342,N_1794);
and U2540 (N_2540,N_1238,N_1160);
nand U2541 (N_2541,N_1981,N_1927);
nand U2542 (N_2542,N_1729,N_1554);
nor U2543 (N_2543,N_1030,N_1650);
nand U2544 (N_2544,N_1150,N_1546);
or U2545 (N_2545,N_1381,N_1395);
nand U2546 (N_2546,N_1787,N_1386);
nand U2547 (N_2547,N_1836,N_1386);
nand U2548 (N_2548,N_1903,N_1460);
and U2549 (N_2549,N_1595,N_1845);
and U2550 (N_2550,N_1938,N_1768);
nor U2551 (N_2551,N_1660,N_1956);
xnor U2552 (N_2552,N_1128,N_1308);
xor U2553 (N_2553,N_1897,N_1337);
xor U2554 (N_2554,N_1023,N_1762);
nor U2555 (N_2555,N_1581,N_1767);
nand U2556 (N_2556,N_1174,N_1606);
xnor U2557 (N_2557,N_1026,N_1318);
nand U2558 (N_2558,N_1843,N_1344);
or U2559 (N_2559,N_1572,N_1544);
and U2560 (N_2560,N_1002,N_1560);
or U2561 (N_2561,N_1150,N_1043);
nand U2562 (N_2562,N_1204,N_1855);
and U2563 (N_2563,N_1642,N_1760);
nor U2564 (N_2564,N_1729,N_1891);
nand U2565 (N_2565,N_1652,N_1608);
and U2566 (N_2566,N_1028,N_1324);
xnor U2567 (N_2567,N_1144,N_1800);
nor U2568 (N_2568,N_1310,N_1841);
or U2569 (N_2569,N_1718,N_1796);
xnor U2570 (N_2570,N_1292,N_1778);
and U2571 (N_2571,N_1377,N_1653);
xor U2572 (N_2572,N_1983,N_1100);
or U2573 (N_2573,N_1886,N_1705);
and U2574 (N_2574,N_1446,N_1473);
nand U2575 (N_2575,N_1256,N_1495);
nand U2576 (N_2576,N_1317,N_1500);
or U2577 (N_2577,N_1922,N_1746);
xor U2578 (N_2578,N_1257,N_1782);
xnor U2579 (N_2579,N_1646,N_1429);
nand U2580 (N_2580,N_1195,N_1836);
nor U2581 (N_2581,N_1747,N_1171);
and U2582 (N_2582,N_1042,N_1680);
or U2583 (N_2583,N_1664,N_1158);
nor U2584 (N_2584,N_1755,N_1705);
xnor U2585 (N_2585,N_1817,N_1616);
xnor U2586 (N_2586,N_1014,N_1376);
nand U2587 (N_2587,N_1435,N_1209);
nor U2588 (N_2588,N_1164,N_1894);
nor U2589 (N_2589,N_1994,N_1565);
nor U2590 (N_2590,N_1115,N_1121);
and U2591 (N_2591,N_1179,N_1981);
and U2592 (N_2592,N_1985,N_1363);
xor U2593 (N_2593,N_1596,N_1251);
or U2594 (N_2594,N_1876,N_1912);
nor U2595 (N_2595,N_1598,N_1074);
nor U2596 (N_2596,N_1784,N_1511);
and U2597 (N_2597,N_1293,N_1026);
nor U2598 (N_2598,N_1527,N_1720);
or U2599 (N_2599,N_1230,N_1973);
nor U2600 (N_2600,N_1222,N_1650);
xnor U2601 (N_2601,N_1165,N_1237);
nand U2602 (N_2602,N_1834,N_1869);
nor U2603 (N_2603,N_1035,N_1878);
or U2604 (N_2604,N_1170,N_1805);
nand U2605 (N_2605,N_1436,N_1311);
and U2606 (N_2606,N_1406,N_1317);
xor U2607 (N_2607,N_1484,N_1512);
xor U2608 (N_2608,N_1604,N_1789);
nand U2609 (N_2609,N_1951,N_1552);
and U2610 (N_2610,N_1008,N_1512);
xor U2611 (N_2611,N_1344,N_1266);
xor U2612 (N_2612,N_1480,N_1270);
or U2613 (N_2613,N_1160,N_1147);
or U2614 (N_2614,N_1705,N_1353);
or U2615 (N_2615,N_1597,N_1325);
or U2616 (N_2616,N_1475,N_1487);
nor U2617 (N_2617,N_1994,N_1926);
and U2618 (N_2618,N_1992,N_1421);
and U2619 (N_2619,N_1117,N_1132);
nor U2620 (N_2620,N_1684,N_1505);
nand U2621 (N_2621,N_1430,N_1624);
nor U2622 (N_2622,N_1558,N_1611);
nor U2623 (N_2623,N_1966,N_1753);
nor U2624 (N_2624,N_1471,N_1431);
nor U2625 (N_2625,N_1604,N_1911);
or U2626 (N_2626,N_1129,N_1390);
nand U2627 (N_2627,N_1217,N_1073);
nor U2628 (N_2628,N_1924,N_1656);
or U2629 (N_2629,N_1204,N_1822);
nand U2630 (N_2630,N_1486,N_1762);
and U2631 (N_2631,N_1371,N_1423);
or U2632 (N_2632,N_1954,N_1121);
nand U2633 (N_2633,N_1017,N_1320);
nor U2634 (N_2634,N_1271,N_1310);
nor U2635 (N_2635,N_1850,N_1021);
and U2636 (N_2636,N_1470,N_1829);
or U2637 (N_2637,N_1042,N_1726);
or U2638 (N_2638,N_1315,N_1194);
and U2639 (N_2639,N_1582,N_1238);
nand U2640 (N_2640,N_1268,N_1007);
nand U2641 (N_2641,N_1148,N_1466);
nand U2642 (N_2642,N_1776,N_1234);
nor U2643 (N_2643,N_1919,N_1311);
and U2644 (N_2644,N_1086,N_1059);
and U2645 (N_2645,N_1535,N_1064);
or U2646 (N_2646,N_1994,N_1899);
or U2647 (N_2647,N_1039,N_1868);
xnor U2648 (N_2648,N_1935,N_1701);
nand U2649 (N_2649,N_1303,N_1265);
nor U2650 (N_2650,N_1700,N_1847);
nand U2651 (N_2651,N_1942,N_1301);
and U2652 (N_2652,N_1382,N_1686);
or U2653 (N_2653,N_1236,N_1442);
or U2654 (N_2654,N_1409,N_1541);
xnor U2655 (N_2655,N_1272,N_1780);
or U2656 (N_2656,N_1324,N_1902);
nand U2657 (N_2657,N_1479,N_1064);
and U2658 (N_2658,N_1774,N_1708);
nand U2659 (N_2659,N_1805,N_1898);
xor U2660 (N_2660,N_1696,N_1402);
and U2661 (N_2661,N_1329,N_1283);
xor U2662 (N_2662,N_1819,N_1198);
nor U2663 (N_2663,N_1310,N_1560);
and U2664 (N_2664,N_1189,N_1937);
xnor U2665 (N_2665,N_1917,N_1529);
or U2666 (N_2666,N_1011,N_1260);
and U2667 (N_2667,N_1327,N_1891);
nor U2668 (N_2668,N_1643,N_1794);
and U2669 (N_2669,N_1269,N_1954);
nand U2670 (N_2670,N_1054,N_1603);
nand U2671 (N_2671,N_1869,N_1821);
and U2672 (N_2672,N_1203,N_1251);
xor U2673 (N_2673,N_1400,N_1457);
nor U2674 (N_2674,N_1614,N_1134);
nor U2675 (N_2675,N_1910,N_1548);
nor U2676 (N_2676,N_1986,N_1922);
xnor U2677 (N_2677,N_1626,N_1197);
nor U2678 (N_2678,N_1051,N_1374);
nor U2679 (N_2679,N_1770,N_1592);
and U2680 (N_2680,N_1095,N_1323);
nor U2681 (N_2681,N_1752,N_1822);
nor U2682 (N_2682,N_1960,N_1519);
nand U2683 (N_2683,N_1867,N_1634);
nor U2684 (N_2684,N_1017,N_1793);
and U2685 (N_2685,N_1532,N_1736);
nor U2686 (N_2686,N_1858,N_1853);
and U2687 (N_2687,N_1217,N_1904);
nand U2688 (N_2688,N_1478,N_1939);
nor U2689 (N_2689,N_1073,N_1117);
nor U2690 (N_2690,N_1817,N_1234);
xor U2691 (N_2691,N_1417,N_1290);
nand U2692 (N_2692,N_1930,N_1817);
or U2693 (N_2693,N_1084,N_1960);
xnor U2694 (N_2694,N_1817,N_1575);
nand U2695 (N_2695,N_1812,N_1551);
or U2696 (N_2696,N_1229,N_1876);
or U2697 (N_2697,N_1318,N_1867);
or U2698 (N_2698,N_1772,N_1037);
xnor U2699 (N_2699,N_1468,N_1383);
and U2700 (N_2700,N_1445,N_1885);
nand U2701 (N_2701,N_1676,N_1846);
xnor U2702 (N_2702,N_1014,N_1411);
nand U2703 (N_2703,N_1595,N_1483);
nand U2704 (N_2704,N_1903,N_1064);
xor U2705 (N_2705,N_1437,N_1245);
xnor U2706 (N_2706,N_1286,N_1237);
and U2707 (N_2707,N_1825,N_1801);
xor U2708 (N_2708,N_1743,N_1126);
and U2709 (N_2709,N_1746,N_1920);
nand U2710 (N_2710,N_1755,N_1937);
or U2711 (N_2711,N_1538,N_1317);
xnor U2712 (N_2712,N_1799,N_1451);
and U2713 (N_2713,N_1083,N_1643);
nand U2714 (N_2714,N_1742,N_1856);
xor U2715 (N_2715,N_1807,N_1916);
and U2716 (N_2716,N_1602,N_1581);
nor U2717 (N_2717,N_1723,N_1809);
nor U2718 (N_2718,N_1443,N_1537);
xor U2719 (N_2719,N_1562,N_1787);
xor U2720 (N_2720,N_1107,N_1653);
and U2721 (N_2721,N_1421,N_1904);
xnor U2722 (N_2722,N_1254,N_1435);
nand U2723 (N_2723,N_1883,N_1834);
and U2724 (N_2724,N_1074,N_1798);
xor U2725 (N_2725,N_1981,N_1205);
or U2726 (N_2726,N_1369,N_1937);
xor U2727 (N_2727,N_1757,N_1430);
xor U2728 (N_2728,N_1163,N_1064);
or U2729 (N_2729,N_1333,N_1886);
xnor U2730 (N_2730,N_1294,N_1945);
nor U2731 (N_2731,N_1691,N_1308);
or U2732 (N_2732,N_1529,N_1442);
nor U2733 (N_2733,N_1796,N_1352);
nand U2734 (N_2734,N_1624,N_1609);
or U2735 (N_2735,N_1825,N_1030);
and U2736 (N_2736,N_1425,N_1487);
and U2737 (N_2737,N_1733,N_1448);
nand U2738 (N_2738,N_1506,N_1954);
nand U2739 (N_2739,N_1888,N_1330);
and U2740 (N_2740,N_1293,N_1346);
and U2741 (N_2741,N_1655,N_1699);
and U2742 (N_2742,N_1967,N_1420);
nand U2743 (N_2743,N_1373,N_1499);
and U2744 (N_2744,N_1871,N_1750);
nand U2745 (N_2745,N_1139,N_1081);
xor U2746 (N_2746,N_1645,N_1048);
and U2747 (N_2747,N_1641,N_1821);
or U2748 (N_2748,N_1969,N_1953);
nand U2749 (N_2749,N_1982,N_1726);
nand U2750 (N_2750,N_1350,N_1556);
or U2751 (N_2751,N_1207,N_1726);
nand U2752 (N_2752,N_1958,N_1108);
and U2753 (N_2753,N_1541,N_1586);
nand U2754 (N_2754,N_1139,N_1895);
or U2755 (N_2755,N_1958,N_1307);
nor U2756 (N_2756,N_1850,N_1674);
nor U2757 (N_2757,N_1333,N_1017);
or U2758 (N_2758,N_1000,N_1111);
or U2759 (N_2759,N_1273,N_1644);
nand U2760 (N_2760,N_1453,N_1534);
nand U2761 (N_2761,N_1888,N_1535);
nor U2762 (N_2762,N_1052,N_1960);
xor U2763 (N_2763,N_1277,N_1913);
xnor U2764 (N_2764,N_1616,N_1918);
xnor U2765 (N_2765,N_1683,N_1351);
nand U2766 (N_2766,N_1652,N_1486);
nor U2767 (N_2767,N_1065,N_1477);
nand U2768 (N_2768,N_1809,N_1578);
nand U2769 (N_2769,N_1587,N_1620);
or U2770 (N_2770,N_1191,N_1941);
or U2771 (N_2771,N_1612,N_1766);
nor U2772 (N_2772,N_1556,N_1094);
nand U2773 (N_2773,N_1473,N_1855);
nand U2774 (N_2774,N_1091,N_1530);
or U2775 (N_2775,N_1975,N_1717);
nor U2776 (N_2776,N_1179,N_1857);
and U2777 (N_2777,N_1125,N_1255);
or U2778 (N_2778,N_1729,N_1005);
or U2779 (N_2779,N_1599,N_1551);
nand U2780 (N_2780,N_1521,N_1062);
xor U2781 (N_2781,N_1003,N_1634);
nand U2782 (N_2782,N_1749,N_1440);
or U2783 (N_2783,N_1770,N_1502);
or U2784 (N_2784,N_1239,N_1331);
xnor U2785 (N_2785,N_1549,N_1223);
nor U2786 (N_2786,N_1059,N_1319);
and U2787 (N_2787,N_1240,N_1136);
xor U2788 (N_2788,N_1959,N_1124);
xnor U2789 (N_2789,N_1782,N_1998);
xnor U2790 (N_2790,N_1364,N_1119);
nand U2791 (N_2791,N_1020,N_1539);
xor U2792 (N_2792,N_1680,N_1829);
nand U2793 (N_2793,N_1705,N_1359);
and U2794 (N_2794,N_1165,N_1870);
nand U2795 (N_2795,N_1854,N_1695);
or U2796 (N_2796,N_1860,N_1619);
and U2797 (N_2797,N_1866,N_1704);
and U2798 (N_2798,N_1770,N_1831);
nand U2799 (N_2799,N_1273,N_1325);
and U2800 (N_2800,N_1096,N_1134);
nor U2801 (N_2801,N_1692,N_1070);
nand U2802 (N_2802,N_1011,N_1085);
nand U2803 (N_2803,N_1698,N_1562);
nand U2804 (N_2804,N_1072,N_1394);
nor U2805 (N_2805,N_1536,N_1210);
xnor U2806 (N_2806,N_1525,N_1466);
nand U2807 (N_2807,N_1548,N_1545);
and U2808 (N_2808,N_1237,N_1563);
or U2809 (N_2809,N_1202,N_1486);
or U2810 (N_2810,N_1590,N_1725);
or U2811 (N_2811,N_1670,N_1843);
and U2812 (N_2812,N_1654,N_1220);
xnor U2813 (N_2813,N_1761,N_1997);
nand U2814 (N_2814,N_1622,N_1157);
or U2815 (N_2815,N_1578,N_1714);
nand U2816 (N_2816,N_1990,N_1207);
nor U2817 (N_2817,N_1344,N_1783);
and U2818 (N_2818,N_1527,N_1633);
nand U2819 (N_2819,N_1338,N_1750);
nor U2820 (N_2820,N_1798,N_1414);
and U2821 (N_2821,N_1690,N_1761);
xor U2822 (N_2822,N_1059,N_1530);
xnor U2823 (N_2823,N_1124,N_1308);
nand U2824 (N_2824,N_1606,N_1131);
nor U2825 (N_2825,N_1472,N_1829);
or U2826 (N_2826,N_1599,N_1361);
nor U2827 (N_2827,N_1108,N_1665);
nand U2828 (N_2828,N_1603,N_1498);
xor U2829 (N_2829,N_1807,N_1268);
and U2830 (N_2830,N_1980,N_1442);
or U2831 (N_2831,N_1358,N_1353);
or U2832 (N_2832,N_1656,N_1860);
or U2833 (N_2833,N_1789,N_1099);
xnor U2834 (N_2834,N_1718,N_1159);
nand U2835 (N_2835,N_1068,N_1348);
xnor U2836 (N_2836,N_1501,N_1801);
and U2837 (N_2837,N_1172,N_1870);
xor U2838 (N_2838,N_1779,N_1306);
and U2839 (N_2839,N_1560,N_1932);
and U2840 (N_2840,N_1007,N_1619);
or U2841 (N_2841,N_1940,N_1003);
or U2842 (N_2842,N_1292,N_1075);
or U2843 (N_2843,N_1700,N_1737);
nor U2844 (N_2844,N_1043,N_1854);
xnor U2845 (N_2845,N_1804,N_1188);
nand U2846 (N_2846,N_1665,N_1480);
nand U2847 (N_2847,N_1236,N_1054);
nand U2848 (N_2848,N_1407,N_1516);
and U2849 (N_2849,N_1090,N_1770);
nor U2850 (N_2850,N_1745,N_1255);
nand U2851 (N_2851,N_1641,N_1591);
nand U2852 (N_2852,N_1752,N_1131);
xor U2853 (N_2853,N_1331,N_1176);
and U2854 (N_2854,N_1292,N_1188);
nor U2855 (N_2855,N_1369,N_1578);
or U2856 (N_2856,N_1978,N_1381);
or U2857 (N_2857,N_1666,N_1997);
nor U2858 (N_2858,N_1368,N_1841);
or U2859 (N_2859,N_1991,N_1961);
or U2860 (N_2860,N_1564,N_1361);
xor U2861 (N_2861,N_1992,N_1278);
xnor U2862 (N_2862,N_1645,N_1146);
nor U2863 (N_2863,N_1693,N_1493);
xnor U2864 (N_2864,N_1590,N_1972);
or U2865 (N_2865,N_1157,N_1613);
xor U2866 (N_2866,N_1268,N_1578);
nand U2867 (N_2867,N_1529,N_1264);
or U2868 (N_2868,N_1263,N_1056);
or U2869 (N_2869,N_1353,N_1090);
or U2870 (N_2870,N_1740,N_1867);
xor U2871 (N_2871,N_1505,N_1430);
nand U2872 (N_2872,N_1771,N_1591);
nor U2873 (N_2873,N_1503,N_1163);
nand U2874 (N_2874,N_1466,N_1465);
xor U2875 (N_2875,N_1400,N_1140);
nand U2876 (N_2876,N_1430,N_1098);
nand U2877 (N_2877,N_1134,N_1236);
nand U2878 (N_2878,N_1798,N_1971);
xnor U2879 (N_2879,N_1626,N_1958);
and U2880 (N_2880,N_1981,N_1869);
and U2881 (N_2881,N_1824,N_1593);
or U2882 (N_2882,N_1169,N_1177);
nand U2883 (N_2883,N_1177,N_1830);
or U2884 (N_2884,N_1742,N_1625);
nand U2885 (N_2885,N_1922,N_1356);
xnor U2886 (N_2886,N_1494,N_1115);
or U2887 (N_2887,N_1035,N_1274);
or U2888 (N_2888,N_1774,N_1374);
nand U2889 (N_2889,N_1813,N_1282);
nand U2890 (N_2890,N_1722,N_1051);
and U2891 (N_2891,N_1413,N_1658);
xor U2892 (N_2892,N_1748,N_1610);
and U2893 (N_2893,N_1347,N_1255);
nand U2894 (N_2894,N_1396,N_1767);
and U2895 (N_2895,N_1199,N_1198);
nor U2896 (N_2896,N_1506,N_1120);
and U2897 (N_2897,N_1478,N_1115);
nor U2898 (N_2898,N_1308,N_1550);
or U2899 (N_2899,N_1000,N_1907);
xor U2900 (N_2900,N_1547,N_1577);
xor U2901 (N_2901,N_1240,N_1327);
xnor U2902 (N_2902,N_1124,N_1115);
and U2903 (N_2903,N_1777,N_1869);
and U2904 (N_2904,N_1881,N_1491);
or U2905 (N_2905,N_1257,N_1958);
and U2906 (N_2906,N_1148,N_1855);
or U2907 (N_2907,N_1316,N_1248);
and U2908 (N_2908,N_1813,N_1806);
and U2909 (N_2909,N_1228,N_1533);
nor U2910 (N_2910,N_1975,N_1465);
nor U2911 (N_2911,N_1249,N_1219);
nand U2912 (N_2912,N_1738,N_1637);
or U2913 (N_2913,N_1436,N_1561);
xor U2914 (N_2914,N_1355,N_1527);
nor U2915 (N_2915,N_1833,N_1402);
and U2916 (N_2916,N_1814,N_1487);
or U2917 (N_2917,N_1858,N_1669);
or U2918 (N_2918,N_1242,N_1603);
and U2919 (N_2919,N_1168,N_1042);
nand U2920 (N_2920,N_1140,N_1635);
nor U2921 (N_2921,N_1812,N_1068);
and U2922 (N_2922,N_1800,N_1520);
and U2923 (N_2923,N_1497,N_1603);
or U2924 (N_2924,N_1139,N_1149);
and U2925 (N_2925,N_1810,N_1476);
and U2926 (N_2926,N_1286,N_1001);
or U2927 (N_2927,N_1752,N_1763);
xor U2928 (N_2928,N_1700,N_1265);
or U2929 (N_2929,N_1141,N_1140);
nand U2930 (N_2930,N_1228,N_1999);
and U2931 (N_2931,N_1891,N_1204);
xnor U2932 (N_2932,N_1235,N_1388);
and U2933 (N_2933,N_1708,N_1640);
and U2934 (N_2934,N_1549,N_1149);
or U2935 (N_2935,N_1380,N_1006);
or U2936 (N_2936,N_1460,N_1920);
and U2937 (N_2937,N_1212,N_1419);
and U2938 (N_2938,N_1465,N_1408);
nor U2939 (N_2939,N_1241,N_1328);
and U2940 (N_2940,N_1104,N_1742);
xor U2941 (N_2941,N_1501,N_1281);
nor U2942 (N_2942,N_1294,N_1818);
or U2943 (N_2943,N_1391,N_1553);
or U2944 (N_2944,N_1279,N_1568);
nor U2945 (N_2945,N_1909,N_1795);
or U2946 (N_2946,N_1401,N_1767);
nand U2947 (N_2947,N_1926,N_1020);
and U2948 (N_2948,N_1900,N_1568);
or U2949 (N_2949,N_1828,N_1119);
xor U2950 (N_2950,N_1829,N_1198);
nor U2951 (N_2951,N_1933,N_1734);
nand U2952 (N_2952,N_1472,N_1899);
xnor U2953 (N_2953,N_1211,N_1668);
nand U2954 (N_2954,N_1980,N_1428);
nand U2955 (N_2955,N_1203,N_1925);
nor U2956 (N_2956,N_1065,N_1159);
nand U2957 (N_2957,N_1750,N_1642);
and U2958 (N_2958,N_1926,N_1687);
or U2959 (N_2959,N_1806,N_1639);
and U2960 (N_2960,N_1378,N_1415);
nand U2961 (N_2961,N_1931,N_1301);
and U2962 (N_2962,N_1911,N_1642);
or U2963 (N_2963,N_1360,N_1981);
and U2964 (N_2964,N_1409,N_1049);
and U2965 (N_2965,N_1464,N_1147);
and U2966 (N_2966,N_1493,N_1142);
nand U2967 (N_2967,N_1417,N_1169);
nor U2968 (N_2968,N_1579,N_1220);
or U2969 (N_2969,N_1459,N_1742);
xor U2970 (N_2970,N_1133,N_1365);
or U2971 (N_2971,N_1131,N_1779);
or U2972 (N_2972,N_1373,N_1222);
and U2973 (N_2973,N_1076,N_1459);
nor U2974 (N_2974,N_1820,N_1620);
or U2975 (N_2975,N_1328,N_1465);
nand U2976 (N_2976,N_1646,N_1947);
nor U2977 (N_2977,N_1948,N_1579);
or U2978 (N_2978,N_1374,N_1823);
or U2979 (N_2979,N_1231,N_1258);
or U2980 (N_2980,N_1606,N_1332);
xnor U2981 (N_2981,N_1219,N_1705);
and U2982 (N_2982,N_1370,N_1380);
nand U2983 (N_2983,N_1863,N_1342);
or U2984 (N_2984,N_1479,N_1845);
or U2985 (N_2985,N_1818,N_1262);
and U2986 (N_2986,N_1325,N_1580);
nand U2987 (N_2987,N_1711,N_1943);
nand U2988 (N_2988,N_1492,N_1247);
and U2989 (N_2989,N_1724,N_1817);
and U2990 (N_2990,N_1032,N_1329);
nand U2991 (N_2991,N_1259,N_1569);
nor U2992 (N_2992,N_1088,N_1384);
xnor U2993 (N_2993,N_1199,N_1541);
nand U2994 (N_2994,N_1611,N_1019);
nor U2995 (N_2995,N_1645,N_1087);
or U2996 (N_2996,N_1743,N_1382);
nor U2997 (N_2997,N_1347,N_1847);
xor U2998 (N_2998,N_1872,N_1320);
or U2999 (N_2999,N_1778,N_1353);
nor U3000 (N_3000,N_2076,N_2032);
nand U3001 (N_3001,N_2951,N_2701);
xnor U3002 (N_3002,N_2341,N_2140);
nand U3003 (N_3003,N_2323,N_2769);
nor U3004 (N_3004,N_2711,N_2114);
and U3005 (N_3005,N_2549,N_2641);
nand U3006 (N_3006,N_2239,N_2523);
nand U3007 (N_3007,N_2040,N_2288);
nand U3008 (N_3008,N_2011,N_2995);
and U3009 (N_3009,N_2803,N_2459);
or U3010 (N_3010,N_2061,N_2853);
nand U3011 (N_3011,N_2103,N_2563);
or U3012 (N_3012,N_2683,N_2691);
nand U3013 (N_3013,N_2539,N_2737);
xnor U3014 (N_3014,N_2677,N_2287);
nor U3015 (N_3015,N_2172,N_2765);
nand U3016 (N_3016,N_2504,N_2059);
or U3017 (N_3017,N_2966,N_2414);
and U3018 (N_3018,N_2536,N_2983);
or U3019 (N_3019,N_2912,N_2532);
nand U3020 (N_3020,N_2715,N_2687);
nand U3021 (N_3021,N_2098,N_2581);
or U3022 (N_3022,N_2418,N_2731);
nor U3023 (N_3023,N_2436,N_2285);
nand U3024 (N_3024,N_2351,N_2516);
or U3025 (N_3025,N_2298,N_2369);
xor U3026 (N_3026,N_2102,N_2545);
nand U3027 (N_3027,N_2343,N_2176);
nor U3028 (N_3028,N_2625,N_2283);
nor U3029 (N_3029,N_2049,N_2222);
nand U3030 (N_3030,N_2502,N_2530);
xnor U3031 (N_3031,N_2881,N_2120);
or U3032 (N_3032,N_2566,N_2484);
xnor U3033 (N_3033,N_2583,N_2847);
nor U3034 (N_3034,N_2774,N_2992);
xnor U3035 (N_3035,N_2470,N_2599);
nor U3036 (N_3036,N_2827,N_2648);
nor U3037 (N_3037,N_2277,N_2713);
and U3038 (N_3038,N_2171,N_2953);
or U3039 (N_3039,N_2888,N_2156);
xnor U3040 (N_3040,N_2155,N_2101);
nor U3041 (N_3041,N_2704,N_2255);
xor U3042 (N_3042,N_2350,N_2699);
or U3043 (N_3043,N_2107,N_2857);
nor U3044 (N_3044,N_2968,N_2196);
or U3045 (N_3045,N_2832,N_2038);
nand U3046 (N_3046,N_2707,N_2919);
nor U3047 (N_3047,N_2430,N_2085);
xor U3048 (N_3048,N_2670,N_2396);
nand U3049 (N_3049,N_2985,N_2634);
nor U3050 (N_3050,N_2465,N_2525);
and U3051 (N_3051,N_2817,N_2117);
and U3052 (N_3052,N_2052,N_2513);
and U3053 (N_3053,N_2237,N_2307);
or U3054 (N_3054,N_2265,N_2392);
or U3055 (N_3055,N_2997,N_2965);
nor U3056 (N_3056,N_2375,N_2408);
or U3057 (N_3057,N_2901,N_2553);
or U3058 (N_3058,N_2791,N_2591);
or U3059 (N_3059,N_2128,N_2201);
nor U3060 (N_3060,N_2570,N_2945);
and U3061 (N_3061,N_2730,N_2001);
nand U3062 (N_3062,N_2329,N_2863);
xnor U3063 (N_3063,N_2007,N_2585);
or U3064 (N_3064,N_2686,N_2131);
nand U3065 (N_3065,N_2862,N_2509);
and U3066 (N_3066,N_2238,N_2145);
nand U3067 (N_3067,N_2931,N_2230);
xnor U3068 (N_3068,N_2478,N_2274);
xnor U3069 (N_3069,N_2104,N_2397);
and U3070 (N_3070,N_2417,N_2772);
xor U3071 (N_3071,N_2554,N_2015);
or U3072 (N_3072,N_2856,N_2506);
xnor U3073 (N_3073,N_2276,N_2666);
and U3074 (N_3074,N_2651,N_2622);
nor U3075 (N_3075,N_2705,N_2439);
and U3076 (N_3076,N_2378,N_2607);
nand U3077 (N_3077,N_2148,N_2796);
xnor U3078 (N_3078,N_2173,N_2998);
and U3079 (N_3079,N_2499,N_2886);
and U3080 (N_3080,N_2161,N_2434);
or U3081 (N_3081,N_2234,N_2629);
or U3082 (N_3082,N_2324,N_2095);
and U3083 (N_3083,N_2046,N_2891);
and U3084 (N_3084,N_2223,N_2093);
or U3085 (N_3085,N_2790,N_2619);
or U3086 (N_3086,N_2267,N_2740);
nand U3087 (N_3087,N_2376,N_2835);
or U3088 (N_3088,N_2170,N_2137);
and U3089 (N_3089,N_2944,N_2003);
and U3090 (N_3090,N_2824,N_2218);
nor U3091 (N_3091,N_2754,N_2957);
xnor U3092 (N_3092,N_2312,N_2169);
nand U3093 (N_3093,N_2349,N_2981);
nor U3094 (N_3094,N_2537,N_2658);
or U3095 (N_3095,N_2527,N_2577);
or U3096 (N_3096,N_2209,N_2647);
xnor U3097 (N_3097,N_2511,N_2895);
or U3098 (N_3098,N_2216,N_2108);
nor U3099 (N_3099,N_2936,N_2004);
and U3100 (N_3100,N_2280,N_2593);
and U3101 (N_3101,N_2240,N_2183);
and U3102 (N_3102,N_2066,N_2159);
nand U3103 (N_3103,N_2531,N_2733);
or U3104 (N_3104,N_2720,N_2675);
nor U3105 (N_3105,N_2541,N_2884);
xnor U3106 (N_3106,N_2958,N_2785);
or U3107 (N_3107,N_2975,N_2952);
and U3108 (N_3108,N_2758,N_2005);
and U3109 (N_3109,N_2556,N_2270);
and U3110 (N_3110,N_2809,N_2567);
nor U3111 (N_3111,N_2197,N_2892);
or U3112 (N_3112,N_2473,N_2828);
nor U3113 (N_3113,N_2249,N_2810);
nor U3114 (N_3114,N_2174,N_2401);
or U3115 (N_3115,N_2657,N_2075);
nor U3116 (N_3116,N_2391,N_2819);
nor U3117 (N_3117,N_2424,N_2048);
xnor U3118 (N_3118,N_2446,N_2843);
and U3119 (N_3119,N_2212,N_2461);
nand U3120 (N_3120,N_2661,N_2008);
xnor U3121 (N_3121,N_2248,N_2193);
or U3122 (N_3122,N_2384,N_2875);
and U3123 (N_3123,N_2800,N_2388);
nand U3124 (N_3124,N_2515,N_2632);
nand U3125 (N_3125,N_2741,N_2512);
or U3126 (N_3126,N_2668,N_2157);
and U3127 (N_3127,N_2637,N_2564);
or U3128 (N_3128,N_2057,N_2825);
nor U3129 (N_3129,N_2425,N_2943);
nor U3130 (N_3130,N_2910,N_2115);
xor U3131 (N_3131,N_2578,N_2894);
nor U3132 (N_3132,N_2551,N_2605);
xnor U3133 (N_3133,N_2986,N_2961);
nand U3134 (N_3134,N_2721,N_2010);
nor U3135 (N_3135,N_2175,N_2487);
or U3136 (N_3136,N_2042,N_2002);
nand U3137 (N_3137,N_2533,N_2921);
xor U3138 (N_3138,N_2153,N_2822);
xnor U3139 (N_3139,N_2595,N_2929);
xnor U3140 (N_3140,N_2660,N_2452);
nor U3141 (N_3141,N_2873,N_2678);
or U3142 (N_3142,N_2177,N_2023);
nand U3143 (N_3143,N_2263,N_2165);
nor U3144 (N_3144,N_2896,N_2882);
and U3145 (N_3145,N_2597,N_2256);
or U3146 (N_3146,N_2543,N_2821);
xor U3147 (N_3147,N_2696,N_2044);
or U3148 (N_3148,N_2594,N_2067);
xnor U3149 (N_3149,N_2991,N_2264);
or U3150 (N_3150,N_2590,N_2962);
nand U3151 (N_3151,N_2782,N_2574);
nand U3152 (N_3152,N_2664,N_2694);
nand U3153 (N_3153,N_2762,N_2372);
and U3154 (N_3154,N_2259,N_2618);
or U3155 (N_3155,N_2208,N_2739);
xnor U3156 (N_3156,N_2804,N_2289);
or U3157 (N_3157,N_2146,N_2292);
or U3158 (N_3158,N_2420,N_2878);
xnor U3159 (N_3159,N_2189,N_2584);
or U3160 (N_3160,N_2559,N_2144);
and U3161 (N_3161,N_2738,N_2013);
and U3162 (N_3162,N_2517,N_2744);
nor U3163 (N_3163,N_2521,N_2451);
or U3164 (N_3164,N_2950,N_2606);
or U3165 (N_3165,N_2770,N_2572);
or U3166 (N_3166,N_2164,N_2088);
nand U3167 (N_3167,N_2316,N_2195);
xnor U3168 (N_3168,N_2411,N_2490);
or U3169 (N_3169,N_2639,N_2295);
nor U3170 (N_3170,N_2609,N_2415);
or U3171 (N_3171,N_2009,N_2464);
nand U3172 (N_3172,N_2442,N_2946);
nand U3173 (N_3173,N_2226,N_2074);
nand U3174 (N_3174,N_2163,N_2868);
xnor U3175 (N_3175,N_2020,N_2444);
xor U3176 (N_3176,N_2488,N_2520);
nand U3177 (N_3177,N_2072,N_2681);
nand U3178 (N_3178,N_2272,N_2054);
and U3179 (N_3179,N_2718,N_2555);
and U3180 (N_3180,N_2132,N_2058);
nor U3181 (N_3181,N_2064,N_2854);
or U3182 (N_3182,N_2271,N_2359);
nor U3183 (N_3183,N_2846,N_2213);
and U3184 (N_3184,N_2304,N_2848);
xnor U3185 (N_3185,N_2775,N_2763);
nor U3186 (N_3186,N_2296,N_2081);
xnor U3187 (N_3187,N_2188,N_2507);
nand U3188 (N_3188,N_2018,N_2231);
xnor U3189 (N_3189,N_2210,N_2709);
nor U3190 (N_3190,N_2253,N_2217);
or U3191 (N_3191,N_2906,N_2037);
nand U3192 (N_3192,N_2385,N_2897);
nand U3193 (N_3193,N_2680,N_2347);
xnor U3194 (N_3194,N_2671,N_2708);
xnor U3195 (N_3195,N_2849,N_2180);
and U3196 (N_3196,N_2982,N_2776);
and U3197 (N_3197,N_2663,N_2766);
xnor U3198 (N_3198,N_2834,N_2063);
or U3199 (N_3199,N_2764,N_2435);
or U3200 (N_3200,N_2938,N_2753);
nand U3201 (N_3201,N_2600,N_2345);
xnor U3202 (N_3202,N_2544,N_2250);
nand U3203 (N_3203,N_2045,N_2105);
nor U3204 (N_3204,N_2876,N_2505);
nor U3205 (N_3205,N_2035,N_2712);
or U3206 (N_3206,N_2149,N_2976);
nor U3207 (N_3207,N_2870,N_2562);
nand U3208 (N_3208,N_2460,N_2529);
and U3209 (N_3209,N_2717,N_2221);
nand U3210 (N_3210,N_2855,N_2016);
or U3211 (N_3211,N_2869,N_2565);
or U3212 (N_3212,N_2603,N_2746);
xnor U3213 (N_3213,N_2330,N_2080);
and U3214 (N_3214,N_2542,N_2322);
nor U3215 (N_3215,N_2728,N_2269);
nand U3216 (N_3216,N_2698,N_2142);
and U3217 (N_3217,N_2202,N_2643);
and U3218 (N_3218,N_2327,N_2242);
and U3219 (N_3219,N_2797,N_2458);
nand U3220 (N_3220,N_2495,N_2914);
nor U3221 (N_3221,N_2727,N_2403);
and U3222 (N_3222,N_2337,N_2662);
xnor U3223 (N_3223,N_2432,N_2191);
or U3224 (N_3224,N_2996,N_2429);
or U3225 (N_3225,N_2281,N_2443);
nand U3226 (N_3226,N_2973,N_2902);
nor U3227 (N_3227,N_2911,N_2909);
xor U3228 (N_3228,N_2192,N_2794);
and U3229 (N_3229,N_2476,N_2748);
xnor U3230 (N_3230,N_2812,N_2722);
nand U3231 (N_3231,N_2336,N_2447);
xor U3232 (N_3232,N_2123,N_2325);
nor U3233 (N_3233,N_2871,N_2926);
xnor U3234 (N_3234,N_2353,N_2649);
or U3235 (N_3235,N_2482,N_2211);
xnor U3236 (N_3236,N_2227,N_2829);
or U3237 (N_3237,N_2154,N_2094);
or U3238 (N_3238,N_2528,N_2302);
or U3239 (N_3239,N_2273,N_2342);
nor U3240 (N_3240,N_2837,N_2127);
and U3241 (N_3241,N_2060,N_2383);
xor U3242 (N_3242,N_2437,N_2241);
or U3243 (N_3243,N_2413,N_2806);
and U3244 (N_3244,N_2700,N_2959);
nor U3245 (N_3245,N_2994,N_2286);
nor U3246 (N_3246,N_2228,N_2284);
and U3247 (N_3247,N_2781,N_2334);
nor U3248 (N_3248,N_2260,N_2510);
nand U3249 (N_3249,N_2308,N_2029);
nand U3250 (N_3250,N_2395,N_2314);
and U3251 (N_3251,N_2409,N_2317);
or U3252 (N_3252,N_2313,N_2017);
nand U3253 (N_3253,N_2031,N_2203);
and U3254 (N_3254,N_2579,N_2757);
and U3255 (N_3255,N_2646,N_2377);
nand U3256 (N_3256,N_2360,N_2747);
nor U3257 (N_3257,N_2078,N_2940);
nor U3258 (N_3258,N_2736,N_2311);
xnor U3259 (N_3259,N_2110,N_2485);
xnor U3260 (N_3260,N_2423,N_2729);
or U3261 (N_3261,N_2224,N_2610);
xor U3262 (N_3262,N_2598,N_2640);
and U3263 (N_3263,N_2568,N_2365);
xor U3264 (N_3264,N_2993,N_2503);
xnor U3265 (N_3265,N_2225,N_2960);
xnor U3266 (N_3266,N_2974,N_2546);
nand U3267 (N_3267,N_2582,N_2596);
or U3268 (N_3268,N_2449,N_2977);
or U3269 (N_3269,N_2462,N_2550);
xor U3270 (N_3270,N_2805,N_2771);
xnor U3271 (N_3271,N_2129,N_2331);
nand U3272 (N_3272,N_2245,N_2162);
xor U3273 (N_3273,N_2320,N_2811);
and U3274 (N_3274,N_2306,N_2310);
nor U3275 (N_3275,N_2780,N_2421);
and U3276 (N_3276,N_2293,N_2150);
nand U3277 (N_3277,N_2971,N_2494);
or U3278 (N_3278,N_2963,N_2084);
xnor U3279 (N_3279,N_2158,N_2022);
nand U3280 (N_3280,N_2820,N_2055);
xor U3281 (N_3281,N_2692,N_2319);
or U3282 (N_3282,N_2328,N_2168);
xor U3283 (N_3283,N_2915,N_2258);
xor U3284 (N_3284,N_2885,N_2669);
xor U3285 (N_3285,N_2589,N_2676);
xor U3286 (N_3286,N_2455,N_2100);
xnor U3287 (N_3287,N_2761,N_2166);
or U3288 (N_3288,N_2339,N_2592);
nor U3289 (N_3289,N_2755,N_2370);
xor U3290 (N_3290,N_2920,N_2742);
and U3291 (N_3291,N_2852,N_2734);
xnor U3292 (N_3292,N_2905,N_2890);
xor U3293 (N_3293,N_2041,N_2089);
and U3294 (N_3294,N_2814,N_2326);
or U3295 (N_3295,N_2925,N_2611);
nor U3296 (N_3296,N_2864,N_2642);
nor U3297 (N_3297,N_2367,N_2466);
nand U3298 (N_3298,N_2299,N_2400);
nand U3299 (N_3299,N_2893,N_2534);
or U3300 (N_3300,N_2399,N_2665);
xnor U3301 (N_3301,N_2069,N_2338);
and U3302 (N_3302,N_2724,N_2489);
nand U3303 (N_3303,N_2404,N_2768);
nand U3304 (N_3304,N_2673,N_2179);
nor U3305 (N_3305,N_2725,N_2019);
nor U3306 (N_3306,N_2082,N_2346);
nand U3307 (N_3307,N_2918,N_2062);
nor U3308 (N_3308,N_2964,N_2500);
nand U3309 (N_3309,N_2538,N_2119);
nand U3310 (N_3310,N_2125,N_2999);
and U3311 (N_3311,N_2109,N_2616);
and U3312 (N_3312,N_2980,N_2898);
xnor U3313 (N_3313,N_2949,N_2695);
nand U3314 (N_3314,N_2118,N_2454);
xor U3315 (N_3315,N_2519,N_2380);
nor U3316 (N_3316,N_2947,N_2087);
xnor U3317 (N_3317,N_2294,N_2624);
nand U3318 (N_3318,N_2627,N_2321);
xnor U3319 (N_3319,N_2071,N_2988);
or U3320 (N_3320,N_2841,N_2937);
or U3321 (N_3321,N_2867,N_2205);
xor U3322 (N_3322,N_2232,N_2047);
xor U3323 (N_3323,N_2039,N_2386);
nor U3324 (N_3324,N_2838,N_2941);
xnor U3325 (N_3325,N_2547,N_2548);
and U3326 (N_3326,N_2877,N_2970);
xor U3327 (N_3327,N_2978,N_2361);
or U3328 (N_3328,N_2097,N_2799);
and U3329 (N_3329,N_2352,N_2151);
nand U3330 (N_3330,N_2623,N_2024);
nor U3331 (N_3331,N_2540,N_2186);
nand U3332 (N_3332,N_2143,N_2410);
or U3333 (N_3333,N_2026,N_2795);
nand U3334 (N_3334,N_2121,N_2552);
xnor U3335 (N_3335,N_2501,N_2786);
or U3336 (N_3336,N_2588,N_2030);
nand U3337 (N_3337,N_2972,N_2381);
or U3338 (N_3338,N_2613,N_2368);
or U3339 (N_3339,N_2823,N_2621);
or U3340 (N_3340,N_2934,N_2469);
or U3341 (N_3341,N_2922,N_2575);
nand U3342 (N_3342,N_2935,N_2928);
or U3343 (N_3343,N_2778,N_2141);
or U3344 (N_3344,N_2363,N_2422);
nand U3345 (N_3345,N_2291,N_2573);
nor U3346 (N_3346,N_2924,N_2569);
and U3347 (N_3347,N_2880,N_2526);
nand U3348 (N_3348,N_2942,N_2684);
or U3349 (N_3349,N_2122,N_2441);
or U3350 (N_3350,N_2077,N_2068);
nand U3351 (N_3351,N_2254,N_2364);
nor U3352 (N_3352,N_2056,N_2850);
xor U3353 (N_3353,N_2356,N_2251);
xor U3354 (N_3354,N_2086,N_2830);
xor U3355 (N_3355,N_2514,N_2990);
nand U3356 (N_3356,N_2252,N_2792);
or U3357 (N_3357,N_2969,N_2620);
and U3358 (N_3358,N_2178,N_2220);
xor U3359 (N_3359,N_2198,N_2858);
or U3360 (N_3360,N_2344,N_2138);
xor U3361 (N_3361,N_2036,N_2126);
nor U3362 (N_3362,N_2112,N_2362);
nor U3363 (N_3363,N_2006,N_2468);
and U3364 (N_3364,N_2644,N_2608);
and U3365 (N_3365,N_2070,N_2842);
nand U3366 (N_3366,N_2628,N_2714);
and U3367 (N_3367,N_2340,N_2073);
nor U3368 (N_3368,N_2358,N_2474);
nand U3369 (N_3369,N_2779,N_2558);
xor U3370 (N_3370,N_2652,N_2366);
and U3371 (N_3371,N_2818,N_2690);
xor U3372 (N_3372,N_2576,N_2246);
xor U3373 (N_3373,N_2518,N_2389);
nor U3374 (N_3374,N_2726,N_2079);
nor U3375 (N_3375,N_2000,N_2426);
nand U3376 (N_3376,N_2839,N_2014);
nor U3377 (N_3377,N_2907,N_2402);
nand U3378 (N_3378,N_2206,N_2913);
xor U3379 (N_3379,N_2152,N_2348);
and U3380 (N_3380,N_2354,N_2735);
or U3381 (N_3381,N_2654,N_2865);
xnor U3382 (N_3382,N_2844,N_2498);
nor U3383 (N_3383,N_2134,N_2394);
and U3384 (N_3384,N_2243,N_2840);
or U3385 (N_3385,N_2390,N_2393);
or U3386 (N_3386,N_2587,N_2851);
xnor U3387 (N_3387,N_2773,N_2745);
xnor U3388 (N_3388,N_2416,N_2214);
xnor U3389 (N_3389,N_2428,N_2453);
or U3390 (N_3390,N_2719,N_2244);
nor U3391 (N_3391,N_2257,N_2147);
nand U3392 (N_3392,N_2908,N_2167);
or U3393 (N_3393,N_2374,N_2379);
and U3394 (N_3394,N_2387,N_2967);
nand U3395 (N_3395,N_2685,N_2065);
nand U3396 (N_3396,N_2229,N_2989);
nor U3397 (N_3397,N_2887,N_2626);
xor U3398 (N_3398,N_2879,N_2382);
xnor U3399 (N_3399,N_2332,N_2614);
nand U3400 (N_3400,N_2560,N_2412);
nor U3401 (N_3401,N_2612,N_2866);
nor U3402 (N_3402,N_2113,N_2752);
nor U3403 (N_3403,N_2638,N_2903);
nand U3404 (N_3404,N_2034,N_2028);
and U3405 (N_3405,N_2784,N_2092);
nor U3406 (N_3406,N_2586,N_2497);
xnor U3407 (N_3407,N_2440,N_2448);
or U3408 (N_3408,N_2053,N_2833);
nor U3409 (N_3409,N_2290,N_2043);
nor U3410 (N_3410,N_2012,N_2266);
nor U3411 (N_3411,N_2801,N_2679);
xnor U3412 (N_3412,N_2027,N_2215);
nor U3413 (N_3413,N_2522,N_2483);
or U3414 (N_3414,N_2406,N_2682);
nor U3415 (N_3415,N_2333,N_2481);
nor U3416 (N_3416,N_2813,N_2508);
and U3417 (N_3417,N_2636,N_2710);
or U3418 (N_3418,N_2802,N_2933);
and U3419 (N_3419,N_2743,N_2207);
xor U3420 (N_3420,N_2979,N_2674);
nand U3421 (N_3421,N_2492,N_2561);
nand U3422 (N_3422,N_2789,N_2956);
xor U3423 (N_3423,N_2486,N_2659);
nand U3424 (N_3424,N_2859,N_2580);
nor U3425 (N_3425,N_2667,N_2635);
xor U3426 (N_3426,N_2706,N_2111);
or U3427 (N_3427,N_2405,N_2315);
xor U3428 (N_3428,N_2091,N_2524);
nor U3429 (N_3429,N_2831,N_2932);
nand U3430 (N_3430,N_2419,N_2874);
and U3431 (N_3431,N_2653,N_2457);
and U3432 (N_3432,N_2645,N_2672);
nor U3433 (N_3433,N_2693,N_2948);
or U3434 (N_3434,N_2357,N_2096);
nor U3435 (N_3435,N_2278,N_2954);
nor U3436 (N_3436,N_2557,N_2025);
and U3437 (N_3437,N_2135,N_2601);
and U3438 (N_3438,N_2496,N_2106);
or U3439 (N_3439,N_2194,N_2181);
or U3440 (N_3440,N_2472,N_2984);
or U3441 (N_3441,N_2261,N_2815);
xor U3442 (N_3442,N_2355,N_2927);
and U3443 (N_3443,N_2631,N_2475);
xor U3444 (N_3444,N_2450,N_2247);
nand U3445 (N_3445,N_2783,N_2427);
xor U3446 (N_3446,N_2275,N_2467);
xor U3447 (N_3447,N_2433,N_2463);
and U3448 (N_3448,N_2493,N_2571);
or U3449 (N_3449,N_2160,N_2445);
xor U3450 (N_3450,N_2872,N_2688);
and U3451 (N_3451,N_2756,N_2916);
xnor U3452 (N_3452,N_2335,N_2305);
nor U3453 (N_3453,N_2050,N_2407);
nand U3454 (N_3454,N_2656,N_2816);
xnor U3455 (N_3455,N_2187,N_2617);
or U3456 (N_3456,N_2438,N_2900);
or U3457 (N_3457,N_2703,N_2182);
nand U3458 (N_3458,N_2301,N_2861);
nand U3459 (N_3459,N_2297,N_2860);
xnor U3460 (N_3460,N_2279,N_2124);
xor U3461 (N_3461,N_2917,N_2139);
or U3462 (N_3462,N_2955,N_2689);
and U3463 (N_3463,N_2808,N_2751);
nor U3464 (N_3464,N_2051,N_2491);
nor U3465 (N_3465,N_2116,N_2759);
and U3466 (N_3466,N_2480,N_2090);
and U3467 (N_3467,N_2750,N_2262);
and U3468 (N_3468,N_2615,N_2889);
nor U3469 (N_3469,N_2236,N_2199);
nor U3470 (N_3470,N_2185,N_2836);
or U3471 (N_3471,N_2723,N_2268);
and U3472 (N_3472,N_2807,N_2471);
and U3473 (N_3473,N_2767,N_2987);
and U3474 (N_3474,N_2303,N_2904);
and U3475 (N_3475,N_2398,N_2697);
xnor U3476 (N_3476,N_2749,N_2130);
nand U3477 (N_3477,N_2235,N_2373);
and U3478 (N_3478,N_2535,N_2371);
and U3479 (N_3479,N_2318,N_2099);
nand U3480 (N_3480,N_2939,N_2477);
nand U3481 (N_3481,N_2788,N_2923);
xor U3482 (N_3482,N_2777,N_2431);
nand U3483 (N_3483,N_2309,N_2760);
xnor U3484 (N_3484,N_2300,N_2204);
and U3485 (N_3485,N_2633,N_2650);
xnor U3486 (N_3486,N_2655,N_2899);
or U3487 (N_3487,N_2282,N_2930);
and U3488 (N_3488,N_2033,N_2826);
or U3489 (N_3489,N_2200,N_2479);
or U3490 (N_3490,N_2798,N_2630);
nand U3491 (N_3491,N_2787,N_2456);
or U3492 (N_3492,N_2083,N_2219);
nand U3493 (N_3493,N_2136,N_2702);
nand U3494 (N_3494,N_2190,N_2133);
nand U3495 (N_3495,N_2716,N_2845);
or U3496 (N_3496,N_2602,N_2021);
and U3497 (N_3497,N_2793,N_2184);
or U3498 (N_3498,N_2604,N_2732);
xor U3499 (N_3499,N_2883,N_2233);
xor U3500 (N_3500,N_2654,N_2361);
xor U3501 (N_3501,N_2796,N_2911);
or U3502 (N_3502,N_2271,N_2186);
xnor U3503 (N_3503,N_2646,N_2359);
or U3504 (N_3504,N_2453,N_2058);
nand U3505 (N_3505,N_2199,N_2109);
nor U3506 (N_3506,N_2349,N_2312);
nor U3507 (N_3507,N_2165,N_2195);
or U3508 (N_3508,N_2570,N_2020);
and U3509 (N_3509,N_2386,N_2896);
nor U3510 (N_3510,N_2765,N_2053);
and U3511 (N_3511,N_2016,N_2160);
nor U3512 (N_3512,N_2912,N_2459);
and U3513 (N_3513,N_2419,N_2493);
and U3514 (N_3514,N_2229,N_2917);
nand U3515 (N_3515,N_2545,N_2958);
xnor U3516 (N_3516,N_2468,N_2639);
or U3517 (N_3517,N_2615,N_2628);
and U3518 (N_3518,N_2912,N_2754);
nor U3519 (N_3519,N_2430,N_2345);
and U3520 (N_3520,N_2215,N_2623);
xor U3521 (N_3521,N_2927,N_2488);
xor U3522 (N_3522,N_2971,N_2657);
and U3523 (N_3523,N_2158,N_2572);
xor U3524 (N_3524,N_2948,N_2827);
or U3525 (N_3525,N_2283,N_2552);
and U3526 (N_3526,N_2706,N_2655);
or U3527 (N_3527,N_2149,N_2307);
xor U3528 (N_3528,N_2616,N_2904);
nor U3529 (N_3529,N_2295,N_2605);
and U3530 (N_3530,N_2574,N_2958);
and U3531 (N_3531,N_2794,N_2109);
xor U3532 (N_3532,N_2568,N_2076);
or U3533 (N_3533,N_2783,N_2563);
or U3534 (N_3534,N_2847,N_2744);
nor U3535 (N_3535,N_2544,N_2595);
nor U3536 (N_3536,N_2997,N_2802);
or U3537 (N_3537,N_2770,N_2277);
or U3538 (N_3538,N_2900,N_2022);
nor U3539 (N_3539,N_2216,N_2092);
nand U3540 (N_3540,N_2328,N_2364);
and U3541 (N_3541,N_2500,N_2476);
nand U3542 (N_3542,N_2191,N_2591);
and U3543 (N_3543,N_2573,N_2093);
nand U3544 (N_3544,N_2358,N_2402);
or U3545 (N_3545,N_2985,N_2763);
and U3546 (N_3546,N_2669,N_2719);
nor U3547 (N_3547,N_2405,N_2685);
or U3548 (N_3548,N_2505,N_2499);
or U3549 (N_3549,N_2189,N_2280);
and U3550 (N_3550,N_2617,N_2041);
xnor U3551 (N_3551,N_2064,N_2143);
and U3552 (N_3552,N_2894,N_2969);
or U3553 (N_3553,N_2199,N_2981);
xnor U3554 (N_3554,N_2952,N_2651);
nand U3555 (N_3555,N_2678,N_2569);
or U3556 (N_3556,N_2044,N_2035);
or U3557 (N_3557,N_2822,N_2693);
and U3558 (N_3558,N_2499,N_2293);
nand U3559 (N_3559,N_2570,N_2673);
xor U3560 (N_3560,N_2025,N_2273);
nand U3561 (N_3561,N_2651,N_2596);
or U3562 (N_3562,N_2020,N_2263);
or U3563 (N_3563,N_2894,N_2973);
xnor U3564 (N_3564,N_2039,N_2704);
xnor U3565 (N_3565,N_2900,N_2837);
nor U3566 (N_3566,N_2337,N_2441);
xor U3567 (N_3567,N_2256,N_2671);
xor U3568 (N_3568,N_2614,N_2378);
and U3569 (N_3569,N_2182,N_2597);
or U3570 (N_3570,N_2932,N_2824);
nor U3571 (N_3571,N_2086,N_2702);
xnor U3572 (N_3572,N_2931,N_2005);
or U3573 (N_3573,N_2413,N_2363);
nor U3574 (N_3574,N_2270,N_2589);
or U3575 (N_3575,N_2279,N_2363);
or U3576 (N_3576,N_2312,N_2452);
and U3577 (N_3577,N_2969,N_2723);
nand U3578 (N_3578,N_2796,N_2658);
and U3579 (N_3579,N_2732,N_2979);
or U3580 (N_3580,N_2705,N_2595);
nand U3581 (N_3581,N_2550,N_2090);
and U3582 (N_3582,N_2869,N_2487);
nor U3583 (N_3583,N_2336,N_2850);
and U3584 (N_3584,N_2805,N_2654);
and U3585 (N_3585,N_2566,N_2075);
or U3586 (N_3586,N_2928,N_2479);
or U3587 (N_3587,N_2159,N_2533);
or U3588 (N_3588,N_2089,N_2210);
and U3589 (N_3589,N_2360,N_2562);
xnor U3590 (N_3590,N_2865,N_2332);
nand U3591 (N_3591,N_2753,N_2414);
nor U3592 (N_3592,N_2339,N_2283);
and U3593 (N_3593,N_2508,N_2271);
nor U3594 (N_3594,N_2799,N_2620);
xnor U3595 (N_3595,N_2737,N_2990);
or U3596 (N_3596,N_2257,N_2206);
or U3597 (N_3597,N_2897,N_2399);
and U3598 (N_3598,N_2666,N_2880);
and U3599 (N_3599,N_2247,N_2237);
and U3600 (N_3600,N_2358,N_2675);
and U3601 (N_3601,N_2004,N_2002);
xnor U3602 (N_3602,N_2326,N_2771);
and U3603 (N_3603,N_2464,N_2861);
and U3604 (N_3604,N_2589,N_2141);
and U3605 (N_3605,N_2816,N_2043);
or U3606 (N_3606,N_2741,N_2951);
xnor U3607 (N_3607,N_2157,N_2111);
xor U3608 (N_3608,N_2163,N_2739);
nand U3609 (N_3609,N_2245,N_2644);
xnor U3610 (N_3610,N_2764,N_2150);
or U3611 (N_3611,N_2996,N_2926);
nand U3612 (N_3612,N_2412,N_2700);
nor U3613 (N_3613,N_2867,N_2528);
or U3614 (N_3614,N_2266,N_2857);
nor U3615 (N_3615,N_2136,N_2726);
xor U3616 (N_3616,N_2022,N_2440);
or U3617 (N_3617,N_2963,N_2704);
nand U3618 (N_3618,N_2447,N_2696);
and U3619 (N_3619,N_2559,N_2956);
nor U3620 (N_3620,N_2401,N_2022);
nand U3621 (N_3621,N_2995,N_2737);
nor U3622 (N_3622,N_2400,N_2171);
nand U3623 (N_3623,N_2431,N_2922);
and U3624 (N_3624,N_2382,N_2362);
xor U3625 (N_3625,N_2010,N_2708);
or U3626 (N_3626,N_2518,N_2865);
and U3627 (N_3627,N_2848,N_2249);
nand U3628 (N_3628,N_2753,N_2600);
or U3629 (N_3629,N_2595,N_2715);
xnor U3630 (N_3630,N_2006,N_2730);
nor U3631 (N_3631,N_2479,N_2145);
or U3632 (N_3632,N_2728,N_2295);
xnor U3633 (N_3633,N_2898,N_2821);
nand U3634 (N_3634,N_2815,N_2648);
or U3635 (N_3635,N_2418,N_2411);
or U3636 (N_3636,N_2165,N_2473);
nand U3637 (N_3637,N_2160,N_2758);
and U3638 (N_3638,N_2641,N_2237);
and U3639 (N_3639,N_2058,N_2996);
nor U3640 (N_3640,N_2748,N_2757);
xor U3641 (N_3641,N_2466,N_2122);
or U3642 (N_3642,N_2662,N_2967);
or U3643 (N_3643,N_2588,N_2545);
xnor U3644 (N_3644,N_2624,N_2262);
or U3645 (N_3645,N_2705,N_2816);
nand U3646 (N_3646,N_2382,N_2080);
xor U3647 (N_3647,N_2912,N_2815);
nand U3648 (N_3648,N_2890,N_2689);
or U3649 (N_3649,N_2653,N_2650);
and U3650 (N_3650,N_2139,N_2081);
and U3651 (N_3651,N_2025,N_2435);
nand U3652 (N_3652,N_2243,N_2473);
nand U3653 (N_3653,N_2227,N_2052);
nor U3654 (N_3654,N_2224,N_2973);
and U3655 (N_3655,N_2369,N_2524);
or U3656 (N_3656,N_2380,N_2574);
xor U3657 (N_3657,N_2133,N_2502);
xor U3658 (N_3658,N_2425,N_2824);
or U3659 (N_3659,N_2493,N_2175);
nor U3660 (N_3660,N_2645,N_2143);
or U3661 (N_3661,N_2970,N_2823);
nor U3662 (N_3662,N_2575,N_2319);
or U3663 (N_3663,N_2202,N_2980);
nor U3664 (N_3664,N_2971,N_2259);
and U3665 (N_3665,N_2057,N_2389);
nor U3666 (N_3666,N_2145,N_2543);
xnor U3667 (N_3667,N_2006,N_2289);
nor U3668 (N_3668,N_2312,N_2197);
or U3669 (N_3669,N_2560,N_2872);
nor U3670 (N_3670,N_2319,N_2141);
or U3671 (N_3671,N_2392,N_2617);
xor U3672 (N_3672,N_2022,N_2009);
and U3673 (N_3673,N_2377,N_2169);
and U3674 (N_3674,N_2251,N_2478);
nand U3675 (N_3675,N_2642,N_2465);
or U3676 (N_3676,N_2780,N_2194);
and U3677 (N_3677,N_2073,N_2377);
and U3678 (N_3678,N_2877,N_2680);
or U3679 (N_3679,N_2991,N_2927);
nor U3680 (N_3680,N_2469,N_2703);
nor U3681 (N_3681,N_2531,N_2645);
xnor U3682 (N_3682,N_2917,N_2884);
nand U3683 (N_3683,N_2967,N_2601);
and U3684 (N_3684,N_2883,N_2139);
nand U3685 (N_3685,N_2221,N_2613);
and U3686 (N_3686,N_2220,N_2166);
xor U3687 (N_3687,N_2124,N_2519);
xnor U3688 (N_3688,N_2360,N_2760);
or U3689 (N_3689,N_2542,N_2361);
nor U3690 (N_3690,N_2492,N_2160);
xor U3691 (N_3691,N_2365,N_2815);
nand U3692 (N_3692,N_2956,N_2107);
and U3693 (N_3693,N_2704,N_2650);
xnor U3694 (N_3694,N_2362,N_2477);
and U3695 (N_3695,N_2558,N_2321);
nor U3696 (N_3696,N_2094,N_2443);
and U3697 (N_3697,N_2308,N_2362);
and U3698 (N_3698,N_2708,N_2301);
or U3699 (N_3699,N_2542,N_2355);
nor U3700 (N_3700,N_2029,N_2213);
nand U3701 (N_3701,N_2144,N_2153);
and U3702 (N_3702,N_2165,N_2215);
xnor U3703 (N_3703,N_2405,N_2050);
nor U3704 (N_3704,N_2944,N_2210);
nand U3705 (N_3705,N_2250,N_2625);
or U3706 (N_3706,N_2624,N_2981);
xor U3707 (N_3707,N_2590,N_2307);
and U3708 (N_3708,N_2754,N_2584);
and U3709 (N_3709,N_2754,N_2558);
or U3710 (N_3710,N_2389,N_2307);
xnor U3711 (N_3711,N_2145,N_2615);
xor U3712 (N_3712,N_2296,N_2927);
xnor U3713 (N_3713,N_2224,N_2388);
xnor U3714 (N_3714,N_2666,N_2748);
nand U3715 (N_3715,N_2478,N_2482);
xor U3716 (N_3716,N_2160,N_2911);
xnor U3717 (N_3717,N_2928,N_2844);
and U3718 (N_3718,N_2647,N_2931);
and U3719 (N_3719,N_2359,N_2469);
nor U3720 (N_3720,N_2074,N_2067);
nor U3721 (N_3721,N_2707,N_2965);
and U3722 (N_3722,N_2081,N_2457);
nand U3723 (N_3723,N_2052,N_2886);
or U3724 (N_3724,N_2836,N_2802);
nor U3725 (N_3725,N_2562,N_2642);
nand U3726 (N_3726,N_2087,N_2713);
and U3727 (N_3727,N_2407,N_2388);
xnor U3728 (N_3728,N_2424,N_2464);
or U3729 (N_3729,N_2569,N_2710);
nor U3730 (N_3730,N_2380,N_2338);
nor U3731 (N_3731,N_2334,N_2582);
xnor U3732 (N_3732,N_2418,N_2873);
xor U3733 (N_3733,N_2289,N_2282);
or U3734 (N_3734,N_2905,N_2538);
and U3735 (N_3735,N_2897,N_2568);
nand U3736 (N_3736,N_2435,N_2730);
and U3737 (N_3737,N_2100,N_2019);
and U3738 (N_3738,N_2659,N_2164);
nand U3739 (N_3739,N_2202,N_2115);
xnor U3740 (N_3740,N_2701,N_2761);
nor U3741 (N_3741,N_2847,N_2654);
nor U3742 (N_3742,N_2970,N_2557);
or U3743 (N_3743,N_2885,N_2862);
nand U3744 (N_3744,N_2141,N_2947);
and U3745 (N_3745,N_2647,N_2702);
nand U3746 (N_3746,N_2221,N_2515);
nand U3747 (N_3747,N_2689,N_2423);
nor U3748 (N_3748,N_2694,N_2006);
or U3749 (N_3749,N_2071,N_2594);
and U3750 (N_3750,N_2669,N_2408);
xnor U3751 (N_3751,N_2628,N_2958);
xor U3752 (N_3752,N_2975,N_2761);
nor U3753 (N_3753,N_2184,N_2468);
or U3754 (N_3754,N_2981,N_2073);
nor U3755 (N_3755,N_2096,N_2473);
nand U3756 (N_3756,N_2672,N_2709);
nand U3757 (N_3757,N_2268,N_2234);
nand U3758 (N_3758,N_2551,N_2614);
and U3759 (N_3759,N_2867,N_2666);
nand U3760 (N_3760,N_2204,N_2747);
nor U3761 (N_3761,N_2193,N_2224);
nor U3762 (N_3762,N_2293,N_2802);
nor U3763 (N_3763,N_2132,N_2254);
nand U3764 (N_3764,N_2020,N_2270);
nand U3765 (N_3765,N_2102,N_2490);
nor U3766 (N_3766,N_2070,N_2039);
xor U3767 (N_3767,N_2231,N_2332);
nor U3768 (N_3768,N_2215,N_2236);
nor U3769 (N_3769,N_2099,N_2003);
and U3770 (N_3770,N_2392,N_2467);
xor U3771 (N_3771,N_2454,N_2318);
nand U3772 (N_3772,N_2100,N_2888);
or U3773 (N_3773,N_2178,N_2009);
or U3774 (N_3774,N_2252,N_2802);
xnor U3775 (N_3775,N_2774,N_2974);
xor U3776 (N_3776,N_2593,N_2097);
and U3777 (N_3777,N_2239,N_2799);
nand U3778 (N_3778,N_2790,N_2039);
and U3779 (N_3779,N_2467,N_2044);
nand U3780 (N_3780,N_2094,N_2836);
and U3781 (N_3781,N_2117,N_2276);
nand U3782 (N_3782,N_2104,N_2531);
nor U3783 (N_3783,N_2750,N_2039);
or U3784 (N_3784,N_2021,N_2664);
or U3785 (N_3785,N_2743,N_2523);
or U3786 (N_3786,N_2699,N_2911);
and U3787 (N_3787,N_2521,N_2714);
xnor U3788 (N_3788,N_2215,N_2039);
xor U3789 (N_3789,N_2447,N_2161);
nor U3790 (N_3790,N_2159,N_2880);
xnor U3791 (N_3791,N_2174,N_2520);
and U3792 (N_3792,N_2571,N_2637);
and U3793 (N_3793,N_2459,N_2412);
nor U3794 (N_3794,N_2779,N_2538);
and U3795 (N_3795,N_2910,N_2854);
nor U3796 (N_3796,N_2232,N_2638);
nor U3797 (N_3797,N_2742,N_2495);
xor U3798 (N_3798,N_2336,N_2865);
or U3799 (N_3799,N_2790,N_2680);
nand U3800 (N_3800,N_2689,N_2541);
nand U3801 (N_3801,N_2582,N_2218);
or U3802 (N_3802,N_2372,N_2964);
and U3803 (N_3803,N_2202,N_2777);
or U3804 (N_3804,N_2448,N_2040);
and U3805 (N_3805,N_2773,N_2088);
and U3806 (N_3806,N_2251,N_2310);
xnor U3807 (N_3807,N_2246,N_2161);
nor U3808 (N_3808,N_2715,N_2341);
or U3809 (N_3809,N_2967,N_2575);
or U3810 (N_3810,N_2915,N_2462);
xnor U3811 (N_3811,N_2874,N_2105);
or U3812 (N_3812,N_2573,N_2090);
nor U3813 (N_3813,N_2108,N_2410);
nand U3814 (N_3814,N_2886,N_2842);
nand U3815 (N_3815,N_2474,N_2289);
or U3816 (N_3816,N_2801,N_2678);
nand U3817 (N_3817,N_2776,N_2118);
or U3818 (N_3818,N_2288,N_2060);
nor U3819 (N_3819,N_2190,N_2545);
or U3820 (N_3820,N_2826,N_2872);
and U3821 (N_3821,N_2567,N_2258);
nor U3822 (N_3822,N_2074,N_2772);
nor U3823 (N_3823,N_2197,N_2266);
or U3824 (N_3824,N_2257,N_2215);
and U3825 (N_3825,N_2427,N_2923);
or U3826 (N_3826,N_2400,N_2500);
or U3827 (N_3827,N_2511,N_2350);
and U3828 (N_3828,N_2976,N_2435);
nor U3829 (N_3829,N_2759,N_2147);
or U3830 (N_3830,N_2237,N_2057);
nand U3831 (N_3831,N_2203,N_2551);
and U3832 (N_3832,N_2845,N_2893);
and U3833 (N_3833,N_2434,N_2774);
nand U3834 (N_3834,N_2219,N_2970);
or U3835 (N_3835,N_2493,N_2355);
nand U3836 (N_3836,N_2875,N_2420);
xnor U3837 (N_3837,N_2099,N_2606);
and U3838 (N_3838,N_2832,N_2301);
and U3839 (N_3839,N_2212,N_2077);
xor U3840 (N_3840,N_2691,N_2763);
or U3841 (N_3841,N_2519,N_2813);
nand U3842 (N_3842,N_2851,N_2345);
and U3843 (N_3843,N_2345,N_2076);
nor U3844 (N_3844,N_2234,N_2646);
nor U3845 (N_3845,N_2057,N_2691);
xor U3846 (N_3846,N_2368,N_2455);
xor U3847 (N_3847,N_2671,N_2849);
and U3848 (N_3848,N_2135,N_2766);
or U3849 (N_3849,N_2896,N_2884);
nand U3850 (N_3850,N_2422,N_2620);
xor U3851 (N_3851,N_2544,N_2599);
xor U3852 (N_3852,N_2978,N_2128);
nor U3853 (N_3853,N_2913,N_2369);
nor U3854 (N_3854,N_2305,N_2883);
or U3855 (N_3855,N_2260,N_2556);
xnor U3856 (N_3856,N_2220,N_2836);
nand U3857 (N_3857,N_2956,N_2543);
nor U3858 (N_3858,N_2044,N_2366);
nand U3859 (N_3859,N_2863,N_2321);
nand U3860 (N_3860,N_2037,N_2796);
and U3861 (N_3861,N_2009,N_2438);
nor U3862 (N_3862,N_2805,N_2963);
xnor U3863 (N_3863,N_2313,N_2943);
or U3864 (N_3864,N_2467,N_2154);
xor U3865 (N_3865,N_2863,N_2137);
or U3866 (N_3866,N_2586,N_2126);
xnor U3867 (N_3867,N_2249,N_2606);
or U3868 (N_3868,N_2704,N_2485);
or U3869 (N_3869,N_2443,N_2129);
nand U3870 (N_3870,N_2263,N_2395);
or U3871 (N_3871,N_2116,N_2141);
or U3872 (N_3872,N_2377,N_2728);
or U3873 (N_3873,N_2791,N_2289);
nor U3874 (N_3874,N_2635,N_2934);
and U3875 (N_3875,N_2380,N_2046);
nand U3876 (N_3876,N_2515,N_2716);
nand U3877 (N_3877,N_2947,N_2206);
nor U3878 (N_3878,N_2547,N_2569);
nand U3879 (N_3879,N_2102,N_2958);
or U3880 (N_3880,N_2271,N_2949);
xnor U3881 (N_3881,N_2819,N_2034);
nor U3882 (N_3882,N_2501,N_2484);
xor U3883 (N_3883,N_2651,N_2452);
nor U3884 (N_3884,N_2754,N_2283);
xor U3885 (N_3885,N_2566,N_2651);
and U3886 (N_3886,N_2293,N_2122);
or U3887 (N_3887,N_2632,N_2742);
and U3888 (N_3888,N_2411,N_2349);
or U3889 (N_3889,N_2850,N_2275);
nand U3890 (N_3890,N_2393,N_2538);
nor U3891 (N_3891,N_2730,N_2082);
nor U3892 (N_3892,N_2944,N_2206);
xnor U3893 (N_3893,N_2617,N_2519);
and U3894 (N_3894,N_2717,N_2746);
nand U3895 (N_3895,N_2049,N_2227);
nor U3896 (N_3896,N_2764,N_2349);
nor U3897 (N_3897,N_2810,N_2595);
xor U3898 (N_3898,N_2160,N_2899);
xor U3899 (N_3899,N_2240,N_2763);
or U3900 (N_3900,N_2465,N_2811);
nor U3901 (N_3901,N_2242,N_2351);
and U3902 (N_3902,N_2916,N_2236);
nand U3903 (N_3903,N_2014,N_2771);
and U3904 (N_3904,N_2304,N_2909);
or U3905 (N_3905,N_2538,N_2428);
nor U3906 (N_3906,N_2142,N_2085);
nor U3907 (N_3907,N_2939,N_2850);
nand U3908 (N_3908,N_2013,N_2339);
or U3909 (N_3909,N_2602,N_2092);
or U3910 (N_3910,N_2592,N_2139);
nor U3911 (N_3911,N_2363,N_2491);
and U3912 (N_3912,N_2001,N_2994);
xor U3913 (N_3913,N_2718,N_2162);
and U3914 (N_3914,N_2609,N_2386);
nand U3915 (N_3915,N_2062,N_2006);
or U3916 (N_3916,N_2697,N_2986);
nor U3917 (N_3917,N_2465,N_2591);
nand U3918 (N_3918,N_2228,N_2520);
nand U3919 (N_3919,N_2324,N_2125);
nand U3920 (N_3920,N_2696,N_2324);
xor U3921 (N_3921,N_2725,N_2955);
nand U3922 (N_3922,N_2903,N_2952);
nor U3923 (N_3923,N_2129,N_2986);
xnor U3924 (N_3924,N_2255,N_2932);
or U3925 (N_3925,N_2390,N_2663);
or U3926 (N_3926,N_2392,N_2131);
nand U3927 (N_3927,N_2081,N_2586);
nand U3928 (N_3928,N_2083,N_2275);
nor U3929 (N_3929,N_2418,N_2315);
xnor U3930 (N_3930,N_2066,N_2333);
xnor U3931 (N_3931,N_2675,N_2817);
and U3932 (N_3932,N_2306,N_2055);
xor U3933 (N_3933,N_2990,N_2008);
xor U3934 (N_3934,N_2113,N_2138);
nand U3935 (N_3935,N_2344,N_2311);
or U3936 (N_3936,N_2783,N_2823);
or U3937 (N_3937,N_2482,N_2362);
nand U3938 (N_3938,N_2785,N_2062);
or U3939 (N_3939,N_2257,N_2799);
nand U3940 (N_3940,N_2785,N_2993);
or U3941 (N_3941,N_2114,N_2914);
or U3942 (N_3942,N_2586,N_2362);
nand U3943 (N_3943,N_2659,N_2781);
and U3944 (N_3944,N_2204,N_2809);
nor U3945 (N_3945,N_2064,N_2862);
nand U3946 (N_3946,N_2531,N_2498);
nand U3947 (N_3947,N_2476,N_2911);
or U3948 (N_3948,N_2053,N_2658);
xor U3949 (N_3949,N_2278,N_2317);
and U3950 (N_3950,N_2982,N_2576);
xor U3951 (N_3951,N_2405,N_2294);
nor U3952 (N_3952,N_2227,N_2304);
xnor U3953 (N_3953,N_2790,N_2995);
or U3954 (N_3954,N_2283,N_2202);
or U3955 (N_3955,N_2278,N_2284);
or U3956 (N_3956,N_2768,N_2006);
xor U3957 (N_3957,N_2346,N_2469);
nand U3958 (N_3958,N_2411,N_2544);
and U3959 (N_3959,N_2531,N_2461);
and U3960 (N_3960,N_2306,N_2796);
and U3961 (N_3961,N_2162,N_2061);
xnor U3962 (N_3962,N_2855,N_2644);
nand U3963 (N_3963,N_2675,N_2464);
nand U3964 (N_3964,N_2635,N_2296);
nand U3965 (N_3965,N_2705,N_2791);
and U3966 (N_3966,N_2084,N_2381);
and U3967 (N_3967,N_2891,N_2014);
nor U3968 (N_3968,N_2610,N_2329);
and U3969 (N_3969,N_2081,N_2806);
and U3970 (N_3970,N_2958,N_2618);
xnor U3971 (N_3971,N_2239,N_2054);
or U3972 (N_3972,N_2204,N_2093);
nand U3973 (N_3973,N_2711,N_2254);
nor U3974 (N_3974,N_2459,N_2537);
nor U3975 (N_3975,N_2829,N_2448);
or U3976 (N_3976,N_2374,N_2333);
nand U3977 (N_3977,N_2332,N_2472);
and U3978 (N_3978,N_2763,N_2480);
or U3979 (N_3979,N_2118,N_2556);
and U3980 (N_3980,N_2440,N_2043);
xnor U3981 (N_3981,N_2201,N_2189);
or U3982 (N_3982,N_2294,N_2107);
nand U3983 (N_3983,N_2499,N_2598);
nand U3984 (N_3984,N_2863,N_2755);
xnor U3985 (N_3985,N_2682,N_2998);
xnor U3986 (N_3986,N_2647,N_2537);
or U3987 (N_3987,N_2487,N_2968);
and U3988 (N_3988,N_2119,N_2918);
nand U3989 (N_3989,N_2258,N_2341);
or U3990 (N_3990,N_2533,N_2262);
xnor U3991 (N_3991,N_2754,N_2994);
nor U3992 (N_3992,N_2513,N_2986);
and U3993 (N_3993,N_2212,N_2876);
or U3994 (N_3994,N_2248,N_2276);
or U3995 (N_3995,N_2645,N_2421);
nand U3996 (N_3996,N_2475,N_2540);
and U3997 (N_3997,N_2699,N_2040);
xnor U3998 (N_3998,N_2475,N_2782);
nand U3999 (N_3999,N_2864,N_2210);
nor U4000 (N_4000,N_3288,N_3217);
nand U4001 (N_4001,N_3073,N_3204);
xnor U4002 (N_4002,N_3958,N_3406);
and U4003 (N_4003,N_3690,N_3069);
nor U4004 (N_4004,N_3911,N_3870);
xnor U4005 (N_4005,N_3248,N_3014);
and U4006 (N_4006,N_3591,N_3006);
or U4007 (N_4007,N_3494,N_3655);
nor U4008 (N_4008,N_3200,N_3873);
or U4009 (N_4009,N_3330,N_3303);
xnor U4010 (N_4010,N_3684,N_3077);
or U4011 (N_4011,N_3434,N_3806);
nand U4012 (N_4012,N_3084,N_3218);
xnor U4013 (N_4013,N_3948,N_3427);
or U4014 (N_4014,N_3514,N_3548);
nor U4015 (N_4015,N_3665,N_3866);
and U4016 (N_4016,N_3348,N_3926);
nor U4017 (N_4017,N_3029,N_3479);
nor U4018 (N_4018,N_3286,N_3225);
xor U4019 (N_4019,N_3780,N_3475);
nor U4020 (N_4020,N_3630,N_3659);
nor U4021 (N_4021,N_3071,N_3679);
nor U4022 (N_4022,N_3867,N_3956);
and U4023 (N_4023,N_3423,N_3589);
and U4024 (N_4024,N_3291,N_3784);
and U4025 (N_4025,N_3505,N_3112);
nand U4026 (N_4026,N_3544,N_3275);
or U4027 (N_4027,N_3818,N_3497);
nor U4028 (N_4028,N_3448,N_3632);
nor U4029 (N_4029,N_3499,N_3741);
or U4030 (N_4030,N_3724,N_3740);
nor U4031 (N_4031,N_3546,N_3436);
nand U4032 (N_4032,N_3731,N_3637);
nand U4033 (N_4033,N_3509,N_3524);
nand U4034 (N_4034,N_3835,N_3369);
and U4035 (N_4035,N_3641,N_3270);
or U4036 (N_4036,N_3067,N_3660);
nor U4037 (N_4037,N_3263,N_3652);
xor U4038 (N_4038,N_3207,N_3120);
and U4039 (N_4039,N_3094,N_3629);
or U4040 (N_4040,N_3139,N_3278);
nor U4041 (N_4041,N_3689,N_3875);
nor U4042 (N_4042,N_3441,N_3726);
and U4043 (N_4043,N_3848,N_3242);
xnor U4044 (N_4044,N_3306,N_3613);
and U4045 (N_4045,N_3919,N_3929);
or U4046 (N_4046,N_3047,N_3667);
nor U4047 (N_4047,N_3876,N_3028);
xnor U4048 (N_4048,N_3066,N_3776);
nor U4049 (N_4049,N_3636,N_3164);
nor U4050 (N_4050,N_3482,N_3778);
and U4051 (N_4051,N_3093,N_3577);
nor U4052 (N_4052,N_3119,N_3393);
xor U4053 (N_4053,N_3705,N_3447);
xnor U4054 (N_4054,N_3566,N_3522);
xor U4055 (N_4055,N_3663,N_3717);
and U4056 (N_4056,N_3944,N_3742);
and U4057 (N_4057,N_3032,N_3203);
or U4058 (N_4058,N_3010,N_3311);
or U4059 (N_4059,N_3481,N_3575);
nor U4060 (N_4060,N_3335,N_3015);
nand U4061 (N_4061,N_3592,N_3949);
and U4062 (N_4062,N_3904,N_3332);
nor U4063 (N_4063,N_3349,N_3520);
xor U4064 (N_4064,N_3430,N_3553);
or U4065 (N_4065,N_3772,N_3621);
nand U4066 (N_4066,N_3765,N_3243);
nor U4067 (N_4067,N_3386,N_3402);
nand U4068 (N_4068,N_3187,N_3221);
nor U4069 (N_4069,N_3860,N_3413);
and U4070 (N_4070,N_3083,N_3209);
nand U4071 (N_4071,N_3343,N_3905);
or U4072 (N_4072,N_3082,N_3839);
nand U4073 (N_4073,N_3519,N_3955);
xor U4074 (N_4074,N_3930,N_3301);
or U4075 (N_4075,N_3820,N_3634);
nand U4076 (N_4076,N_3049,N_3896);
xnor U4077 (N_4077,N_3931,N_3991);
nand U4078 (N_4078,N_3739,N_3357);
and U4079 (N_4079,N_3709,N_3421);
nand U4080 (N_4080,N_3523,N_3838);
nor U4081 (N_4081,N_3967,N_3939);
nand U4082 (N_4082,N_3317,N_3147);
nand U4083 (N_4083,N_3893,N_3650);
nand U4084 (N_4084,N_3972,N_3236);
nor U4085 (N_4085,N_3194,N_3000);
nor U4086 (N_4086,N_3272,N_3247);
nor U4087 (N_4087,N_3053,N_3359);
xnor U4088 (N_4088,N_3233,N_3950);
nand U4089 (N_4089,N_3574,N_3572);
nor U4090 (N_4090,N_3175,N_3170);
nor U4091 (N_4091,N_3785,N_3358);
xor U4092 (N_4092,N_3859,N_3401);
nor U4093 (N_4093,N_3114,N_3858);
xor U4094 (N_4094,N_3294,N_3622);
or U4095 (N_4095,N_3816,N_3452);
and U4096 (N_4096,N_3669,N_3962);
xor U4097 (N_4097,N_3188,N_3189);
or U4098 (N_4098,N_3850,N_3855);
and U4099 (N_4099,N_3989,N_3582);
or U4100 (N_4100,N_3791,N_3122);
and U4101 (N_4101,N_3789,N_3018);
xnor U4102 (N_4102,N_3283,N_3970);
or U4103 (N_4103,N_3150,N_3975);
or U4104 (N_4104,N_3923,N_3543);
xnor U4105 (N_4105,N_3292,N_3124);
xnor U4106 (N_4106,N_3063,N_3033);
nand U4107 (N_4107,N_3353,N_3998);
or U4108 (N_4108,N_3722,N_3107);
or U4109 (N_4109,N_3298,N_3536);
nor U4110 (N_4110,N_3415,N_3422);
nor U4111 (N_4111,N_3597,N_3994);
nor U4112 (N_4112,N_3437,N_3815);
xnor U4113 (N_4113,N_3959,N_3134);
nand U4114 (N_4114,N_3163,N_3885);
nor U4115 (N_4115,N_3501,N_3091);
nand U4116 (N_4116,N_3503,N_3912);
nand U4117 (N_4117,N_3617,N_3891);
and U4118 (N_4118,N_3079,N_3644);
nand U4119 (N_4119,N_3414,N_3165);
nand U4120 (N_4120,N_3156,N_3313);
or U4121 (N_4121,N_3356,N_3823);
or U4122 (N_4122,N_3732,N_3770);
or U4123 (N_4123,N_3057,N_3439);
xnor U4124 (N_4124,N_3444,N_3065);
nand U4125 (N_4125,N_3915,N_3048);
xnor U4126 (N_4126,N_3039,N_3372);
xnor U4127 (N_4127,N_3109,N_3232);
and U4128 (N_4128,N_3058,N_3419);
nor U4129 (N_4129,N_3877,N_3390);
nand U4130 (N_4130,N_3932,N_3586);
or U4131 (N_4131,N_3351,N_3800);
or U4132 (N_4132,N_3516,N_3830);
xor U4133 (N_4133,N_3723,N_3310);
nor U4134 (N_4134,N_3677,N_3141);
xor U4135 (N_4135,N_3092,N_3697);
xor U4136 (N_4136,N_3545,N_3469);
nor U4137 (N_4137,N_3746,N_3003);
nand U4138 (N_4138,N_3990,N_3149);
or U4139 (N_4139,N_3625,N_3542);
or U4140 (N_4140,N_3155,N_3551);
nor U4141 (N_4141,N_3133,N_3676);
and U4142 (N_4142,N_3786,N_3809);
nor U4143 (N_4143,N_3927,N_3244);
nor U4144 (N_4144,N_3396,N_3797);
nor U4145 (N_4145,N_3276,N_3355);
xnor U4146 (N_4146,N_3052,N_3813);
xnor U4147 (N_4147,N_3704,N_3824);
nor U4148 (N_4148,N_3730,N_3296);
nor U4149 (N_4149,N_3579,N_3309);
xnor U4150 (N_4150,N_3515,N_3999);
and U4151 (N_4151,N_3417,N_3320);
nor U4152 (N_4152,N_3836,N_3727);
and U4153 (N_4153,N_3087,N_3090);
or U4154 (N_4154,N_3025,N_3454);
or U4155 (N_4155,N_3115,N_3059);
nor U4156 (N_4156,N_3535,N_3375);
xor U4157 (N_4157,N_3701,N_3455);
xnor U4158 (N_4158,N_3504,N_3779);
nand U4159 (N_4159,N_3965,N_3817);
xnor U4160 (N_4160,N_3861,N_3166);
xor U4161 (N_4161,N_3183,N_3947);
and U4162 (N_4162,N_3054,N_3795);
or U4163 (N_4163,N_3321,N_3235);
xor U4164 (N_4164,N_3849,N_3841);
or U4165 (N_4165,N_3097,N_3078);
nor U4166 (N_4166,N_3653,N_3131);
nor U4167 (N_4167,N_3633,N_3814);
and U4168 (N_4168,N_3022,N_3997);
and U4169 (N_4169,N_3521,N_3675);
nand U4170 (N_4170,N_3555,N_3719);
or U4171 (N_4171,N_3237,N_3347);
and U4172 (N_4172,N_3981,N_3012);
nor U4173 (N_4173,N_3416,N_3318);
nor U4174 (N_4174,N_3500,N_3853);
nand U4175 (N_4175,N_3095,N_3027);
nor U4176 (N_4176,N_3196,N_3651);
nand U4177 (N_4177,N_3408,N_3388);
nand U4178 (N_4178,N_3743,N_3716);
nor U4179 (N_4179,N_3464,N_3395);
nor U4180 (N_4180,N_3510,N_3277);
xnor U4181 (N_4181,N_3623,N_3532);
nor U4182 (N_4182,N_3987,N_3710);
xor U4183 (N_4183,N_3174,N_3692);
nor U4184 (N_4184,N_3736,N_3898);
xor U4185 (N_4185,N_3599,N_3255);
nand U4186 (N_4186,N_3993,N_3037);
nor U4187 (N_4187,N_3755,N_3411);
or U4188 (N_4188,N_3483,N_3996);
and U4189 (N_4189,N_3338,N_3334);
or U4190 (N_4190,N_3002,N_3089);
or U4191 (N_4191,N_3009,N_3127);
or U4192 (N_4192,N_3230,N_3365);
nor U4193 (N_4193,N_3664,N_3280);
nand U4194 (N_4194,N_3790,N_3878);
xor U4195 (N_4195,N_3506,N_3160);
xnor U4196 (N_4196,N_3403,N_3412);
nor U4197 (N_4197,N_3714,N_3474);
nand U4198 (N_4198,N_3034,N_3088);
xnor U4199 (N_4199,N_3863,N_3668);
and U4200 (N_4200,N_3370,N_3264);
nor U4201 (N_4201,N_3945,N_3256);
nor U4202 (N_4202,N_3587,N_3565);
or U4203 (N_4203,N_3612,N_3289);
nor U4204 (N_4204,N_3980,N_3645);
nor U4205 (N_4205,N_3748,N_3902);
and U4206 (N_4206,N_3178,N_3627);
or U4207 (N_4207,N_3397,N_3104);
and U4208 (N_4208,N_3450,N_3721);
and U4209 (N_4209,N_3713,N_3061);
nand U4210 (N_4210,N_3894,N_3470);
xor U4211 (N_4211,N_3908,N_3268);
nand U4212 (N_4212,N_3459,N_3352);
nor U4213 (N_4213,N_3857,N_3041);
and U4214 (N_4214,N_3478,N_3021);
xor U4215 (N_4215,N_3030,N_3661);
nor U4216 (N_4216,N_3773,N_3140);
xnor U4217 (N_4217,N_3974,N_3238);
xnor U4218 (N_4218,N_3538,N_3252);
nand U4219 (N_4219,N_3763,N_3529);
or U4220 (N_4220,N_3314,N_3143);
and U4221 (N_4221,N_3312,N_3512);
nor U4222 (N_4222,N_3821,N_3913);
and U4223 (N_4223,N_3620,N_3971);
and U4224 (N_4224,N_3890,N_3060);
nor U4225 (N_4225,N_3451,N_3747);
or U4226 (N_4226,N_3605,N_3328);
nor U4227 (N_4227,N_3865,N_3552);
nor U4228 (N_4228,N_3608,N_3327);
nand U4229 (N_4229,N_3805,N_3757);
nand U4230 (N_4230,N_3812,N_3261);
nand U4231 (N_4231,N_3775,N_3564);
and U4232 (N_4232,N_3363,N_3480);
nor U4233 (N_4233,N_3085,N_3583);
or U4234 (N_4234,N_3936,N_3300);
nor U4235 (N_4235,N_3837,N_3562);
xnor U4236 (N_4236,N_3429,N_3585);
xnor U4237 (N_4237,N_3639,N_3273);
nor U4238 (N_4238,N_3703,N_3628);
or U4239 (N_4239,N_3984,N_3978);
and U4240 (N_4240,N_3219,N_3135);
xor U4241 (N_4241,N_3842,N_3517);
and U4242 (N_4242,N_3560,N_3561);
and U4243 (N_4243,N_3550,N_3304);
nor U4244 (N_4244,N_3154,N_3316);
or U4245 (N_4245,N_3121,N_3466);
or U4246 (N_4246,N_3642,N_3745);
nand U4247 (N_4247,N_3619,N_3195);
xor U4248 (N_4248,N_3662,N_3986);
nor U4249 (N_4249,N_3654,N_3610);
nor U4250 (N_4250,N_3920,N_3371);
and U4251 (N_4251,N_3964,N_3138);
xnor U4252 (N_4252,N_3125,N_3700);
nand U4253 (N_4253,N_3907,N_3428);
nand U4254 (N_4254,N_3151,N_3738);
and U4255 (N_4255,N_3148,N_3274);
nand U4256 (N_4256,N_3126,N_3308);
nor U4257 (N_4257,N_3110,N_3979);
nor U4258 (N_4258,N_3854,N_3381);
xnor U4259 (N_4259,N_3040,N_3366);
or U4260 (N_4260,N_3952,N_3391);
nor U4261 (N_4261,N_3011,N_3081);
or U4262 (N_4262,N_3262,N_3957);
nand U4263 (N_4263,N_3693,N_3305);
and U4264 (N_4264,N_3489,N_3803);
nor U4265 (N_4265,N_3377,N_3581);
nand U4266 (N_4266,N_3631,N_3250);
nor U4267 (N_4267,N_3493,N_3603);
or U4268 (N_4268,N_3744,N_3229);
nand U4269 (N_4269,N_3333,N_3976);
or U4270 (N_4270,N_3531,N_3206);
nor U4271 (N_4271,N_3568,N_3337);
or U4272 (N_4272,N_3265,N_3339);
xor U4273 (N_4273,N_3076,N_3137);
nor U4274 (N_4274,N_3389,N_3442);
and U4275 (N_4275,N_3511,N_3008);
or U4276 (N_4276,N_3508,N_3281);
nor U4277 (N_4277,N_3426,N_3168);
nor U4278 (N_4278,N_3758,N_3768);
or U4279 (N_4279,N_3573,N_3559);
and U4280 (N_4280,N_3656,N_3344);
nor U4281 (N_4281,N_3394,N_3099);
xor U4282 (N_4282,N_3346,N_3044);
xor U4283 (N_4283,N_3862,N_3977);
xnor U4284 (N_4284,N_3802,N_3883);
xor U4285 (N_4285,N_3068,N_3223);
and U4286 (N_4286,N_3686,N_3062);
nor U4287 (N_4287,N_3173,N_3198);
xor U4288 (N_4288,N_3539,N_3671);
nand U4289 (N_4289,N_3036,N_3525);
nand U4290 (N_4290,N_3602,N_3874);
nand U4291 (N_4291,N_3934,N_3215);
or U4292 (N_4292,N_3982,N_3694);
nor U4293 (N_4293,N_3285,N_3191);
nor U4294 (N_4294,N_3762,N_3540);
and U4295 (N_4295,N_3941,N_3491);
nor U4296 (N_4296,N_3624,N_3100);
nor U4297 (N_4297,N_3105,N_3513);
nand U4298 (N_4298,N_3829,N_3162);
nor U4299 (N_4299,N_3496,N_3373);
or U4300 (N_4300,N_3647,N_3903);
nor U4301 (N_4301,N_3329,N_3208);
nand U4302 (N_4302,N_3781,N_3595);
and U4303 (N_4303,N_3340,N_3869);
or U4304 (N_4304,N_3611,N_3899);
and U4305 (N_4305,N_3988,N_3350);
or U4306 (N_4306,N_3074,N_3407);
and U4307 (N_4307,N_3995,N_3326);
or U4308 (N_4308,N_3213,N_3845);
nor U4309 (N_4309,N_3533,N_3492);
nand U4310 (N_4310,N_3844,N_3942);
nor U4311 (N_4311,N_3658,N_3753);
and U4312 (N_4312,N_3128,N_3596);
nor U4313 (N_4313,N_3578,N_3354);
or U4314 (N_4314,N_3488,N_3751);
nand U4315 (N_4315,N_3678,N_3794);
xnor U4316 (N_4316,N_3360,N_3635);
nand U4317 (N_4317,N_3224,N_3146);
xor U4318 (N_4318,N_3212,N_3144);
and U4319 (N_4319,N_3897,N_3901);
or U4320 (N_4320,N_3681,N_3868);
nor U4321 (N_4321,N_3457,N_3240);
or U4322 (N_4322,N_3969,N_3881);
nor U4323 (N_4323,N_3670,N_3171);
nand U4324 (N_4324,N_3072,N_3588);
xnor U4325 (N_4325,N_3331,N_3928);
or U4326 (N_4326,N_3017,N_3192);
nand U4327 (N_4327,N_3123,N_3013);
xnor U4328 (N_4328,N_3176,N_3271);
xor U4329 (N_4329,N_3290,N_3961);
and U4330 (N_4330,N_3056,N_3259);
or U4331 (N_4331,N_3810,N_3387);
nand U4332 (N_4332,N_3819,N_3117);
nand U4333 (N_4333,N_3251,N_3020);
nor U4334 (N_4334,N_3832,N_3563);
xnor U4335 (N_4335,N_3777,N_3879);
xor U4336 (N_4336,N_3638,N_3383);
or U4337 (N_4337,N_3438,N_3473);
or U4338 (N_4338,N_3759,N_3487);
xor U4339 (N_4339,N_3895,N_3769);
nand U4340 (N_4340,N_3534,N_3657);
nand U4341 (N_4341,N_3080,N_3527);
nand U4342 (N_4342,N_3900,N_3297);
or U4343 (N_4343,N_3910,N_3729);
xor U4344 (N_4344,N_3458,N_3502);
nor U4345 (N_4345,N_3606,N_3718);
xnor U4346 (N_4346,N_3465,N_3463);
xnor U4347 (N_4347,N_3699,N_3197);
and U4348 (N_4348,N_3646,N_3205);
or U4349 (N_4349,N_3179,N_3707);
and U4350 (N_4350,N_3851,N_3616);
or U4351 (N_4351,N_3211,N_3345);
nand U4352 (N_4352,N_3886,N_3210);
nor U4353 (N_4353,N_3129,N_3571);
nand U4354 (N_4354,N_3698,N_3440);
and U4355 (N_4355,N_3136,N_3456);
or U4356 (N_4356,N_3973,N_3376);
nand U4357 (N_4357,N_3185,N_3600);
and U4358 (N_4358,N_3557,N_3547);
nor U4359 (N_4359,N_3096,N_3368);
xor U4360 (N_4360,N_3361,N_3295);
and U4361 (N_4361,N_3051,N_3254);
nor U4362 (N_4362,N_3822,N_3498);
and U4363 (N_4363,N_3055,N_3946);
nor U4364 (N_4364,N_3688,N_3378);
or U4365 (N_4365,N_3601,N_3342);
and U4366 (N_4366,N_3598,N_3951);
xnor U4367 (N_4367,N_3766,N_3756);
or U4368 (N_4368,N_3834,N_3398);
nor U4369 (N_4369,N_3968,N_3827);
nor U4370 (N_4370,N_3324,N_3453);
or U4371 (N_4371,N_3798,N_3880);
nand U4372 (N_4372,N_3385,N_3943);
xnor U4373 (N_4373,N_3788,N_3249);
nor U4374 (N_4374,N_3924,N_3992);
or U4375 (N_4375,N_3169,N_3098);
and U4376 (N_4376,N_3963,N_3284);
nor U4377 (N_4377,N_3490,N_3476);
or U4378 (N_4378,N_3222,N_3594);
and U4379 (N_4379,N_3177,N_3446);
nand U4380 (N_4380,N_3399,N_3761);
nor U4381 (N_4381,N_3673,N_3672);
or U4382 (N_4382,N_3214,N_3925);
nor U4383 (N_4383,N_3228,N_3269);
nand U4384 (N_4384,N_3220,N_3685);
or U4385 (N_4385,N_3840,N_3026);
and U4386 (N_4386,N_3202,N_3193);
or U4387 (N_4387,N_3158,N_3728);
xnor U4388 (N_4388,N_3917,N_3260);
nor U4389 (N_4389,N_3167,N_3691);
and U4390 (N_4390,N_3760,N_3216);
or U4391 (N_4391,N_3906,N_3528);
nor U4392 (N_4392,N_3038,N_3180);
xor U4393 (N_4393,N_3468,N_3793);
nor U4394 (N_4394,N_3570,N_3425);
and U4395 (N_4395,N_3418,N_3367);
xnor U4396 (N_4396,N_3674,N_3828);
or U4397 (N_4397,N_3181,N_3884);
and U4398 (N_4398,N_3299,N_3796);
nand U4399 (N_4399,N_3246,N_3231);
or U4400 (N_4400,N_3695,N_3764);
nor U4401 (N_4401,N_3102,N_3045);
nand U4402 (N_4402,N_3683,N_3737);
and U4403 (N_4403,N_3954,N_3584);
nor U4404 (N_4404,N_3118,N_3435);
or U4405 (N_4405,N_3257,N_3364);
and U4406 (N_4406,N_3130,N_3856);
nor U4407 (N_4407,N_3725,N_3307);
xor U4408 (N_4408,N_3576,N_3031);
and U4409 (N_4409,N_3420,N_3293);
nor U4410 (N_4410,N_3172,N_3733);
nor U4411 (N_4411,N_3882,N_3101);
or U4412 (N_4412,N_3405,N_3922);
and U4413 (N_4413,N_3558,N_3404);
xor U4414 (N_4414,N_3801,N_3921);
nand U4415 (N_4415,N_3752,N_3266);
nor U4416 (N_4416,N_3282,N_3462);
xor U4417 (N_4417,N_3864,N_3161);
and U4418 (N_4418,N_3241,N_3019);
nor U4419 (N_4419,N_3537,N_3384);
nor U4420 (N_4420,N_3409,N_3715);
nand U4421 (N_4421,N_3182,N_3593);
and U4422 (N_4422,N_3050,N_3199);
nor U4423 (N_4423,N_3774,N_3070);
nor U4424 (N_4424,N_3771,N_3042);
and U4425 (N_4425,N_3892,N_3935);
or U4426 (N_4426,N_3916,N_3460);
or U4427 (N_4427,N_3825,N_3495);
or U4428 (N_4428,N_3315,N_3024);
or U4429 (N_4429,N_3735,N_3445);
and U4430 (N_4430,N_3750,N_3507);
xor U4431 (N_4431,N_3549,N_3734);
or U4432 (N_4432,N_3322,N_3145);
nand U4433 (N_4433,N_3159,N_3467);
and U4434 (N_4434,N_3833,N_3471);
xor U4435 (N_4435,N_3258,N_3245);
or U4436 (N_4436,N_3323,N_3847);
or U4437 (N_4437,N_3708,N_3615);
nor U4438 (N_4438,N_3607,N_3909);
or U4439 (N_4439,N_3108,N_3767);
nand U4440 (N_4440,N_3554,N_3227);
nand U4441 (N_4441,N_3190,N_3424);
xor U4442 (N_4442,N_3604,N_3103);
xnor U4443 (N_4443,N_3783,N_3712);
or U4444 (N_4444,N_3754,N_3807);
or U4445 (N_4445,N_3287,N_3648);
nand U4446 (N_4446,N_3449,N_3113);
nand U4447 (N_4447,N_3541,N_3400);
and U4448 (N_4448,N_3319,N_3702);
nand U4449 (N_4449,N_3852,N_3279);
or U4450 (N_4450,N_3485,N_3914);
and U4451 (N_4451,N_3614,N_3787);
nand U4452 (N_4452,N_3302,N_3918);
nand U4453 (N_4453,N_3804,N_3808);
nand U4454 (N_4454,N_3938,N_3267);
nor U4455 (N_4455,N_3443,N_3872);
nand U4456 (N_4456,N_3016,N_3720);
nand U4457 (N_4457,N_3142,N_3530);
nor U4458 (N_4458,N_3239,N_3116);
and U4459 (N_4459,N_3831,N_3043);
and U4460 (N_4460,N_3687,N_3846);
or U4461 (N_4461,N_3086,N_3472);
nor U4462 (N_4462,N_3392,N_3518);
nand U4463 (N_4463,N_3001,N_3484);
nand U4464 (N_4464,N_3432,N_3640);
xnor U4465 (N_4465,N_3792,N_3711);
xnor U4466 (N_4466,N_3749,N_3580);
or U4467 (N_4467,N_3526,N_3410);
xnor U4468 (N_4468,N_3609,N_3843);
nand U4469 (N_4469,N_3153,N_3132);
and U4470 (N_4470,N_3706,N_3888);
nand U4471 (N_4471,N_3960,N_3682);
or U4472 (N_4472,N_3618,N_3184);
and U4473 (N_4473,N_3666,N_3226);
xnor U4474 (N_4474,N_3007,N_3782);
nor U4475 (N_4475,N_3643,N_3871);
and U4476 (N_4476,N_3887,N_3374);
or U4477 (N_4477,N_3889,N_3023);
or U4478 (N_4478,N_3380,N_3937);
or U4479 (N_4479,N_3433,N_3075);
xor U4480 (N_4480,N_3811,N_3336);
xnor U4481 (N_4481,N_3004,N_3035);
nand U4482 (N_4482,N_3953,N_3696);
and U4483 (N_4483,N_3201,N_3005);
or U4484 (N_4484,N_3983,N_3157);
or U4485 (N_4485,N_3111,N_3431);
xor U4486 (N_4486,N_3461,N_3649);
or U4487 (N_4487,N_3106,N_3826);
or U4488 (N_4488,N_3985,N_3152);
nor U4489 (N_4489,N_3362,N_3569);
or U4490 (N_4490,N_3234,N_3379);
or U4491 (N_4491,N_3186,N_3325);
and U4492 (N_4492,N_3486,N_3933);
and U4493 (N_4493,N_3626,N_3253);
nand U4494 (N_4494,N_3341,N_3046);
nor U4495 (N_4495,N_3966,N_3799);
nor U4496 (N_4496,N_3590,N_3680);
nor U4497 (N_4497,N_3567,N_3382);
and U4498 (N_4498,N_3556,N_3940);
or U4499 (N_4499,N_3064,N_3477);
and U4500 (N_4500,N_3345,N_3068);
and U4501 (N_4501,N_3671,N_3918);
nor U4502 (N_4502,N_3542,N_3581);
nand U4503 (N_4503,N_3776,N_3094);
or U4504 (N_4504,N_3312,N_3687);
xnor U4505 (N_4505,N_3615,N_3024);
and U4506 (N_4506,N_3213,N_3850);
nand U4507 (N_4507,N_3746,N_3551);
nor U4508 (N_4508,N_3204,N_3395);
xor U4509 (N_4509,N_3900,N_3382);
nand U4510 (N_4510,N_3137,N_3784);
nor U4511 (N_4511,N_3368,N_3486);
or U4512 (N_4512,N_3349,N_3255);
and U4513 (N_4513,N_3056,N_3605);
or U4514 (N_4514,N_3460,N_3827);
nand U4515 (N_4515,N_3636,N_3733);
xnor U4516 (N_4516,N_3831,N_3183);
or U4517 (N_4517,N_3458,N_3284);
and U4518 (N_4518,N_3275,N_3480);
or U4519 (N_4519,N_3616,N_3870);
nand U4520 (N_4520,N_3402,N_3074);
xnor U4521 (N_4521,N_3911,N_3675);
and U4522 (N_4522,N_3679,N_3865);
xnor U4523 (N_4523,N_3199,N_3305);
nand U4524 (N_4524,N_3005,N_3261);
xnor U4525 (N_4525,N_3054,N_3576);
and U4526 (N_4526,N_3542,N_3668);
or U4527 (N_4527,N_3677,N_3242);
or U4528 (N_4528,N_3918,N_3004);
nand U4529 (N_4529,N_3365,N_3749);
or U4530 (N_4530,N_3990,N_3268);
and U4531 (N_4531,N_3868,N_3228);
nand U4532 (N_4532,N_3538,N_3008);
or U4533 (N_4533,N_3608,N_3478);
nand U4534 (N_4534,N_3564,N_3873);
nand U4535 (N_4535,N_3068,N_3901);
or U4536 (N_4536,N_3635,N_3654);
nand U4537 (N_4537,N_3798,N_3789);
or U4538 (N_4538,N_3433,N_3989);
and U4539 (N_4539,N_3978,N_3121);
or U4540 (N_4540,N_3282,N_3717);
or U4541 (N_4541,N_3114,N_3979);
xor U4542 (N_4542,N_3809,N_3946);
xor U4543 (N_4543,N_3926,N_3850);
xnor U4544 (N_4544,N_3935,N_3615);
nand U4545 (N_4545,N_3203,N_3424);
and U4546 (N_4546,N_3130,N_3592);
or U4547 (N_4547,N_3631,N_3235);
and U4548 (N_4548,N_3645,N_3262);
and U4549 (N_4549,N_3474,N_3412);
nand U4550 (N_4550,N_3437,N_3750);
nor U4551 (N_4551,N_3384,N_3998);
xor U4552 (N_4552,N_3347,N_3673);
xnor U4553 (N_4553,N_3178,N_3137);
nor U4554 (N_4554,N_3203,N_3772);
nand U4555 (N_4555,N_3421,N_3973);
nor U4556 (N_4556,N_3875,N_3083);
nand U4557 (N_4557,N_3170,N_3252);
nor U4558 (N_4558,N_3585,N_3257);
nor U4559 (N_4559,N_3670,N_3463);
and U4560 (N_4560,N_3790,N_3533);
xnor U4561 (N_4561,N_3883,N_3221);
nor U4562 (N_4562,N_3993,N_3897);
and U4563 (N_4563,N_3130,N_3974);
nand U4564 (N_4564,N_3807,N_3925);
nor U4565 (N_4565,N_3317,N_3161);
and U4566 (N_4566,N_3149,N_3230);
or U4567 (N_4567,N_3538,N_3247);
nand U4568 (N_4568,N_3113,N_3305);
xor U4569 (N_4569,N_3652,N_3817);
xnor U4570 (N_4570,N_3253,N_3616);
or U4571 (N_4571,N_3595,N_3952);
nand U4572 (N_4572,N_3391,N_3721);
nand U4573 (N_4573,N_3910,N_3930);
and U4574 (N_4574,N_3233,N_3895);
nand U4575 (N_4575,N_3553,N_3727);
nand U4576 (N_4576,N_3400,N_3833);
and U4577 (N_4577,N_3545,N_3268);
nor U4578 (N_4578,N_3412,N_3385);
nand U4579 (N_4579,N_3107,N_3251);
nand U4580 (N_4580,N_3381,N_3938);
nor U4581 (N_4581,N_3151,N_3836);
nor U4582 (N_4582,N_3728,N_3650);
or U4583 (N_4583,N_3303,N_3644);
and U4584 (N_4584,N_3971,N_3185);
nor U4585 (N_4585,N_3233,N_3181);
and U4586 (N_4586,N_3829,N_3535);
and U4587 (N_4587,N_3888,N_3605);
xnor U4588 (N_4588,N_3178,N_3621);
or U4589 (N_4589,N_3762,N_3201);
and U4590 (N_4590,N_3196,N_3176);
nor U4591 (N_4591,N_3944,N_3243);
nand U4592 (N_4592,N_3210,N_3909);
and U4593 (N_4593,N_3078,N_3096);
and U4594 (N_4594,N_3884,N_3518);
nand U4595 (N_4595,N_3676,N_3618);
nand U4596 (N_4596,N_3428,N_3196);
nor U4597 (N_4597,N_3184,N_3423);
xor U4598 (N_4598,N_3491,N_3333);
nor U4599 (N_4599,N_3473,N_3106);
xor U4600 (N_4600,N_3041,N_3505);
and U4601 (N_4601,N_3893,N_3377);
nand U4602 (N_4602,N_3806,N_3533);
and U4603 (N_4603,N_3294,N_3955);
or U4604 (N_4604,N_3938,N_3556);
xnor U4605 (N_4605,N_3228,N_3163);
or U4606 (N_4606,N_3606,N_3032);
nand U4607 (N_4607,N_3343,N_3278);
nand U4608 (N_4608,N_3018,N_3605);
or U4609 (N_4609,N_3313,N_3344);
xnor U4610 (N_4610,N_3677,N_3205);
nand U4611 (N_4611,N_3439,N_3394);
xor U4612 (N_4612,N_3812,N_3853);
nor U4613 (N_4613,N_3606,N_3180);
or U4614 (N_4614,N_3280,N_3698);
nor U4615 (N_4615,N_3650,N_3875);
nor U4616 (N_4616,N_3394,N_3244);
and U4617 (N_4617,N_3676,N_3139);
nand U4618 (N_4618,N_3598,N_3937);
xnor U4619 (N_4619,N_3532,N_3484);
nand U4620 (N_4620,N_3919,N_3882);
xor U4621 (N_4621,N_3212,N_3436);
xnor U4622 (N_4622,N_3907,N_3810);
xnor U4623 (N_4623,N_3409,N_3608);
nor U4624 (N_4624,N_3168,N_3804);
xor U4625 (N_4625,N_3372,N_3443);
and U4626 (N_4626,N_3021,N_3961);
nand U4627 (N_4627,N_3513,N_3519);
or U4628 (N_4628,N_3443,N_3505);
nor U4629 (N_4629,N_3326,N_3976);
nand U4630 (N_4630,N_3110,N_3708);
xor U4631 (N_4631,N_3199,N_3047);
or U4632 (N_4632,N_3139,N_3586);
nor U4633 (N_4633,N_3403,N_3427);
xor U4634 (N_4634,N_3575,N_3644);
or U4635 (N_4635,N_3253,N_3697);
nor U4636 (N_4636,N_3329,N_3823);
nand U4637 (N_4637,N_3726,N_3091);
or U4638 (N_4638,N_3882,N_3060);
or U4639 (N_4639,N_3797,N_3021);
and U4640 (N_4640,N_3225,N_3151);
or U4641 (N_4641,N_3155,N_3412);
nor U4642 (N_4642,N_3423,N_3079);
or U4643 (N_4643,N_3737,N_3348);
nor U4644 (N_4644,N_3983,N_3067);
nor U4645 (N_4645,N_3932,N_3087);
nor U4646 (N_4646,N_3326,N_3807);
or U4647 (N_4647,N_3984,N_3866);
xor U4648 (N_4648,N_3016,N_3539);
xnor U4649 (N_4649,N_3800,N_3666);
and U4650 (N_4650,N_3167,N_3661);
nor U4651 (N_4651,N_3555,N_3685);
and U4652 (N_4652,N_3819,N_3913);
nor U4653 (N_4653,N_3118,N_3813);
nor U4654 (N_4654,N_3892,N_3053);
xnor U4655 (N_4655,N_3883,N_3576);
and U4656 (N_4656,N_3710,N_3525);
or U4657 (N_4657,N_3927,N_3536);
nor U4658 (N_4658,N_3527,N_3567);
or U4659 (N_4659,N_3510,N_3015);
xnor U4660 (N_4660,N_3329,N_3197);
nor U4661 (N_4661,N_3544,N_3636);
and U4662 (N_4662,N_3075,N_3686);
and U4663 (N_4663,N_3786,N_3026);
xnor U4664 (N_4664,N_3687,N_3426);
or U4665 (N_4665,N_3008,N_3449);
nand U4666 (N_4666,N_3655,N_3610);
or U4667 (N_4667,N_3816,N_3921);
xor U4668 (N_4668,N_3640,N_3731);
and U4669 (N_4669,N_3473,N_3650);
nand U4670 (N_4670,N_3151,N_3570);
nand U4671 (N_4671,N_3094,N_3367);
xnor U4672 (N_4672,N_3800,N_3335);
xor U4673 (N_4673,N_3227,N_3653);
nand U4674 (N_4674,N_3110,N_3206);
nor U4675 (N_4675,N_3472,N_3944);
and U4676 (N_4676,N_3487,N_3441);
nand U4677 (N_4677,N_3638,N_3109);
nor U4678 (N_4678,N_3105,N_3209);
and U4679 (N_4679,N_3300,N_3670);
and U4680 (N_4680,N_3145,N_3886);
nand U4681 (N_4681,N_3103,N_3966);
nor U4682 (N_4682,N_3167,N_3816);
and U4683 (N_4683,N_3580,N_3016);
xor U4684 (N_4684,N_3664,N_3169);
nand U4685 (N_4685,N_3931,N_3054);
nand U4686 (N_4686,N_3148,N_3077);
nand U4687 (N_4687,N_3961,N_3967);
xor U4688 (N_4688,N_3167,N_3409);
nand U4689 (N_4689,N_3547,N_3036);
and U4690 (N_4690,N_3441,N_3439);
or U4691 (N_4691,N_3657,N_3109);
or U4692 (N_4692,N_3362,N_3087);
xor U4693 (N_4693,N_3232,N_3330);
and U4694 (N_4694,N_3868,N_3637);
nand U4695 (N_4695,N_3516,N_3562);
xor U4696 (N_4696,N_3716,N_3314);
nand U4697 (N_4697,N_3091,N_3911);
nand U4698 (N_4698,N_3413,N_3700);
or U4699 (N_4699,N_3036,N_3054);
or U4700 (N_4700,N_3161,N_3002);
nor U4701 (N_4701,N_3907,N_3148);
nand U4702 (N_4702,N_3421,N_3339);
or U4703 (N_4703,N_3322,N_3152);
xor U4704 (N_4704,N_3849,N_3327);
nor U4705 (N_4705,N_3311,N_3974);
xor U4706 (N_4706,N_3956,N_3263);
and U4707 (N_4707,N_3566,N_3183);
or U4708 (N_4708,N_3939,N_3569);
nor U4709 (N_4709,N_3893,N_3474);
nand U4710 (N_4710,N_3866,N_3525);
nor U4711 (N_4711,N_3210,N_3689);
xor U4712 (N_4712,N_3674,N_3974);
nor U4713 (N_4713,N_3985,N_3558);
nand U4714 (N_4714,N_3066,N_3085);
and U4715 (N_4715,N_3089,N_3012);
nand U4716 (N_4716,N_3551,N_3780);
nor U4717 (N_4717,N_3394,N_3353);
or U4718 (N_4718,N_3224,N_3708);
xnor U4719 (N_4719,N_3044,N_3521);
or U4720 (N_4720,N_3916,N_3177);
nor U4721 (N_4721,N_3318,N_3881);
and U4722 (N_4722,N_3957,N_3187);
nor U4723 (N_4723,N_3508,N_3396);
and U4724 (N_4724,N_3715,N_3752);
and U4725 (N_4725,N_3735,N_3118);
and U4726 (N_4726,N_3598,N_3031);
nor U4727 (N_4727,N_3623,N_3973);
xnor U4728 (N_4728,N_3340,N_3836);
nand U4729 (N_4729,N_3719,N_3940);
nor U4730 (N_4730,N_3290,N_3597);
nand U4731 (N_4731,N_3416,N_3156);
or U4732 (N_4732,N_3738,N_3755);
xor U4733 (N_4733,N_3421,N_3488);
and U4734 (N_4734,N_3976,N_3742);
nand U4735 (N_4735,N_3001,N_3376);
xor U4736 (N_4736,N_3751,N_3805);
nand U4737 (N_4737,N_3342,N_3521);
nand U4738 (N_4738,N_3625,N_3912);
nand U4739 (N_4739,N_3149,N_3625);
nor U4740 (N_4740,N_3468,N_3657);
xor U4741 (N_4741,N_3709,N_3303);
nor U4742 (N_4742,N_3933,N_3869);
and U4743 (N_4743,N_3548,N_3116);
nor U4744 (N_4744,N_3501,N_3167);
nand U4745 (N_4745,N_3151,N_3611);
and U4746 (N_4746,N_3274,N_3164);
and U4747 (N_4747,N_3380,N_3711);
nor U4748 (N_4748,N_3948,N_3667);
or U4749 (N_4749,N_3975,N_3265);
and U4750 (N_4750,N_3142,N_3065);
nor U4751 (N_4751,N_3780,N_3579);
nor U4752 (N_4752,N_3942,N_3302);
or U4753 (N_4753,N_3264,N_3230);
and U4754 (N_4754,N_3615,N_3965);
or U4755 (N_4755,N_3792,N_3875);
nor U4756 (N_4756,N_3847,N_3015);
or U4757 (N_4757,N_3234,N_3657);
and U4758 (N_4758,N_3391,N_3473);
or U4759 (N_4759,N_3835,N_3946);
nand U4760 (N_4760,N_3688,N_3564);
nand U4761 (N_4761,N_3467,N_3145);
and U4762 (N_4762,N_3952,N_3169);
xnor U4763 (N_4763,N_3896,N_3736);
nor U4764 (N_4764,N_3129,N_3476);
and U4765 (N_4765,N_3987,N_3981);
nor U4766 (N_4766,N_3608,N_3267);
nor U4767 (N_4767,N_3613,N_3480);
xor U4768 (N_4768,N_3199,N_3736);
nor U4769 (N_4769,N_3706,N_3841);
xnor U4770 (N_4770,N_3622,N_3077);
and U4771 (N_4771,N_3359,N_3572);
or U4772 (N_4772,N_3340,N_3079);
nor U4773 (N_4773,N_3441,N_3399);
and U4774 (N_4774,N_3198,N_3983);
and U4775 (N_4775,N_3363,N_3672);
or U4776 (N_4776,N_3519,N_3046);
nand U4777 (N_4777,N_3683,N_3129);
and U4778 (N_4778,N_3275,N_3496);
nand U4779 (N_4779,N_3901,N_3067);
and U4780 (N_4780,N_3085,N_3207);
or U4781 (N_4781,N_3900,N_3870);
nor U4782 (N_4782,N_3931,N_3874);
nor U4783 (N_4783,N_3937,N_3469);
xor U4784 (N_4784,N_3964,N_3089);
and U4785 (N_4785,N_3698,N_3339);
and U4786 (N_4786,N_3250,N_3513);
and U4787 (N_4787,N_3141,N_3154);
nand U4788 (N_4788,N_3005,N_3817);
nor U4789 (N_4789,N_3287,N_3832);
or U4790 (N_4790,N_3088,N_3894);
and U4791 (N_4791,N_3338,N_3341);
xnor U4792 (N_4792,N_3333,N_3263);
xnor U4793 (N_4793,N_3671,N_3057);
xor U4794 (N_4794,N_3217,N_3347);
and U4795 (N_4795,N_3593,N_3541);
xnor U4796 (N_4796,N_3909,N_3375);
or U4797 (N_4797,N_3861,N_3739);
xor U4798 (N_4798,N_3662,N_3212);
xnor U4799 (N_4799,N_3013,N_3897);
xor U4800 (N_4800,N_3135,N_3149);
and U4801 (N_4801,N_3485,N_3722);
and U4802 (N_4802,N_3763,N_3512);
and U4803 (N_4803,N_3943,N_3378);
or U4804 (N_4804,N_3867,N_3942);
or U4805 (N_4805,N_3617,N_3688);
xor U4806 (N_4806,N_3909,N_3125);
or U4807 (N_4807,N_3987,N_3630);
and U4808 (N_4808,N_3625,N_3410);
or U4809 (N_4809,N_3441,N_3602);
nor U4810 (N_4810,N_3927,N_3731);
nand U4811 (N_4811,N_3606,N_3588);
nand U4812 (N_4812,N_3698,N_3012);
and U4813 (N_4813,N_3477,N_3260);
nor U4814 (N_4814,N_3280,N_3600);
and U4815 (N_4815,N_3461,N_3239);
nor U4816 (N_4816,N_3005,N_3048);
or U4817 (N_4817,N_3082,N_3306);
nand U4818 (N_4818,N_3541,N_3407);
xnor U4819 (N_4819,N_3484,N_3920);
or U4820 (N_4820,N_3595,N_3616);
nor U4821 (N_4821,N_3327,N_3125);
and U4822 (N_4822,N_3968,N_3195);
xor U4823 (N_4823,N_3482,N_3765);
xnor U4824 (N_4824,N_3030,N_3640);
xor U4825 (N_4825,N_3043,N_3314);
nor U4826 (N_4826,N_3298,N_3603);
xor U4827 (N_4827,N_3919,N_3868);
and U4828 (N_4828,N_3040,N_3759);
xnor U4829 (N_4829,N_3773,N_3322);
or U4830 (N_4830,N_3741,N_3272);
xnor U4831 (N_4831,N_3121,N_3212);
nor U4832 (N_4832,N_3515,N_3061);
and U4833 (N_4833,N_3100,N_3129);
nor U4834 (N_4834,N_3870,N_3562);
xnor U4835 (N_4835,N_3027,N_3034);
nor U4836 (N_4836,N_3330,N_3607);
xor U4837 (N_4837,N_3105,N_3424);
and U4838 (N_4838,N_3604,N_3651);
xnor U4839 (N_4839,N_3521,N_3587);
xnor U4840 (N_4840,N_3674,N_3670);
nand U4841 (N_4841,N_3684,N_3694);
nor U4842 (N_4842,N_3297,N_3167);
xnor U4843 (N_4843,N_3114,N_3028);
or U4844 (N_4844,N_3967,N_3557);
xnor U4845 (N_4845,N_3142,N_3909);
or U4846 (N_4846,N_3817,N_3188);
nor U4847 (N_4847,N_3155,N_3505);
or U4848 (N_4848,N_3081,N_3831);
xnor U4849 (N_4849,N_3899,N_3698);
xor U4850 (N_4850,N_3114,N_3810);
and U4851 (N_4851,N_3559,N_3306);
and U4852 (N_4852,N_3619,N_3503);
xnor U4853 (N_4853,N_3573,N_3625);
xnor U4854 (N_4854,N_3854,N_3566);
nand U4855 (N_4855,N_3447,N_3066);
xnor U4856 (N_4856,N_3609,N_3478);
and U4857 (N_4857,N_3423,N_3805);
xnor U4858 (N_4858,N_3492,N_3017);
and U4859 (N_4859,N_3734,N_3559);
or U4860 (N_4860,N_3509,N_3884);
nor U4861 (N_4861,N_3394,N_3535);
nor U4862 (N_4862,N_3489,N_3449);
xor U4863 (N_4863,N_3573,N_3990);
xnor U4864 (N_4864,N_3451,N_3949);
nor U4865 (N_4865,N_3260,N_3643);
nor U4866 (N_4866,N_3482,N_3440);
and U4867 (N_4867,N_3606,N_3789);
nand U4868 (N_4868,N_3262,N_3391);
or U4869 (N_4869,N_3893,N_3090);
or U4870 (N_4870,N_3930,N_3715);
and U4871 (N_4871,N_3489,N_3119);
nor U4872 (N_4872,N_3350,N_3415);
nor U4873 (N_4873,N_3915,N_3413);
or U4874 (N_4874,N_3082,N_3135);
nor U4875 (N_4875,N_3579,N_3039);
and U4876 (N_4876,N_3894,N_3701);
xor U4877 (N_4877,N_3696,N_3932);
nand U4878 (N_4878,N_3639,N_3740);
nor U4879 (N_4879,N_3075,N_3477);
nand U4880 (N_4880,N_3994,N_3873);
xnor U4881 (N_4881,N_3623,N_3287);
xnor U4882 (N_4882,N_3621,N_3345);
nor U4883 (N_4883,N_3980,N_3431);
or U4884 (N_4884,N_3712,N_3771);
nor U4885 (N_4885,N_3894,N_3473);
and U4886 (N_4886,N_3997,N_3734);
nor U4887 (N_4887,N_3198,N_3120);
nand U4888 (N_4888,N_3799,N_3318);
nand U4889 (N_4889,N_3984,N_3512);
and U4890 (N_4890,N_3666,N_3822);
nor U4891 (N_4891,N_3094,N_3721);
and U4892 (N_4892,N_3595,N_3234);
or U4893 (N_4893,N_3304,N_3221);
nand U4894 (N_4894,N_3705,N_3988);
nand U4895 (N_4895,N_3191,N_3907);
nor U4896 (N_4896,N_3364,N_3244);
and U4897 (N_4897,N_3277,N_3365);
nor U4898 (N_4898,N_3018,N_3432);
nand U4899 (N_4899,N_3970,N_3171);
and U4900 (N_4900,N_3300,N_3854);
nand U4901 (N_4901,N_3311,N_3212);
or U4902 (N_4902,N_3880,N_3290);
nand U4903 (N_4903,N_3897,N_3717);
xor U4904 (N_4904,N_3817,N_3722);
xnor U4905 (N_4905,N_3397,N_3520);
nand U4906 (N_4906,N_3909,N_3746);
or U4907 (N_4907,N_3488,N_3289);
nor U4908 (N_4908,N_3434,N_3732);
nand U4909 (N_4909,N_3065,N_3022);
nand U4910 (N_4910,N_3503,N_3894);
xnor U4911 (N_4911,N_3032,N_3592);
nor U4912 (N_4912,N_3790,N_3427);
and U4913 (N_4913,N_3062,N_3236);
nor U4914 (N_4914,N_3414,N_3847);
nor U4915 (N_4915,N_3068,N_3660);
nor U4916 (N_4916,N_3512,N_3378);
xor U4917 (N_4917,N_3594,N_3071);
or U4918 (N_4918,N_3096,N_3154);
and U4919 (N_4919,N_3736,N_3829);
or U4920 (N_4920,N_3796,N_3776);
nand U4921 (N_4921,N_3126,N_3056);
xnor U4922 (N_4922,N_3152,N_3126);
nand U4923 (N_4923,N_3087,N_3509);
xor U4924 (N_4924,N_3371,N_3498);
nor U4925 (N_4925,N_3411,N_3591);
xor U4926 (N_4926,N_3168,N_3246);
xor U4927 (N_4927,N_3639,N_3302);
nor U4928 (N_4928,N_3242,N_3600);
xnor U4929 (N_4929,N_3998,N_3718);
or U4930 (N_4930,N_3702,N_3554);
and U4931 (N_4931,N_3296,N_3977);
nand U4932 (N_4932,N_3205,N_3471);
nand U4933 (N_4933,N_3788,N_3196);
or U4934 (N_4934,N_3099,N_3603);
or U4935 (N_4935,N_3115,N_3084);
nor U4936 (N_4936,N_3658,N_3130);
xnor U4937 (N_4937,N_3029,N_3360);
or U4938 (N_4938,N_3186,N_3797);
or U4939 (N_4939,N_3767,N_3421);
and U4940 (N_4940,N_3268,N_3707);
or U4941 (N_4941,N_3415,N_3596);
nand U4942 (N_4942,N_3291,N_3970);
nand U4943 (N_4943,N_3214,N_3392);
xnor U4944 (N_4944,N_3464,N_3938);
or U4945 (N_4945,N_3729,N_3480);
nand U4946 (N_4946,N_3502,N_3026);
nand U4947 (N_4947,N_3947,N_3667);
and U4948 (N_4948,N_3597,N_3427);
or U4949 (N_4949,N_3176,N_3575);
nand U4950 (N_4950,N_3133,N_3693);
nor U4951 (N_4951,N_3056,N_3386);
xnor U4952 (N_4952,N_3518,N_3633);
nor U4953 (N_4953,N_3833,N_3141);
nor U4954 (N_4954,N_3391,N_3632);
xnor U4955 (N_4955,N_3441,N_3419);
nand U4956 (N_4956,N_3425,N_3784);
or U4957 (N_4957,N_3245,N_3433);
and U4958 (N_4958,N_3809,N_3523);
or U4959 (N_4959,N_3600,N_3612);
nand U4960 (N_4960,N_3382,N_3711);
nor U4961 (N_4961,N_3526,N_3035);
nor U4962 (N_4962,N_3830,N_3235);
nor U4963 (N_4963,N_3297,N_3035);
nor U4964 (N_4964,N_3033,N_3218);
nor U4965 (N_4965,N_3743,N_3250);
xor U4966 (N_4966,N_3573,N_3715);
and U4967 (N_4967,N_3644,N_3770);
nand U4968 (N_4968,N_3897,N_3899);
nor U4969 (N_4969,N_3282,N_3112);
nand U4970 (N_4970,N_3612,N_3324);
and U4971 (N_4971,N_3060,N_3966);
or U4972 (N_4972,N_3603,N_3477);
xor U4973 (N_4973,N_3014,N_3104);
nor U4974 (N_4974,N_3369,N_3093);
xnor U4975 (N_4975,N_3474,N_3037);
or U4976 (N_4976,N_3468,N_3652);
nor U4977 (N_4977,N_3856,N_3330);
nor U4978 (N_4978,N_3089,N_3271);
xnor U4979 (N_4979,N_3485,N_3740);
xor U4980 (N_4980,N_3251,N_3699);
nand U4981 (N_4981,N_3965,N_3196);
xnor U4982 (N_4982,N_3696,N_3927);
nor U4983 (N_4983,N_3557,N_3488);
and U4984 (N_4984,N_3068,N_3034);
nand U4985 (N_4985,N_3639,N_3891);
nand U4986 (N_4986,N_3446,N_3073);
nand U4987 (N_4987,N_3028,N_3229);
and U4988 (N_4988,N_3840,N_3223);
xnor U4989 (N_4989,N_3031,N_3888);
or U4990 (N_4990,N_3581,N_3428);
xnor U4991 (N_4991,N_3176,N_3472);
nor U4992 (N_4992,N_3200,N_3543);
and U4993 (N_4993,N_3500,N_3760);
or U4994 (N_4994,N_3174,N_3920);
nand U4995 (N_4995,N_3885,N_3056);
or U4996 (N_4996,N_3689,N_3379);
and U4997 (N_4997,N_3880,N_3626);
xor U4998 (N_4998,N_3560,N_3230);
nand U4999 (N_4999,N_3195,N_3283);
or UO_0 (O_0,N_4493,N_4017);
xor UO_1 (O_1,N_4437,N_4343);
and UO_2 (O_2,N_4953,N_4451);
or UO_3 (O_3,N_4967,N_4519);
nand UO_4 (O_4,N_4187,N_4290);
nor UO_5 (O_5,N_4701,N_4047);
nand UO_6 (O_6,N_4293,N_4863);
nor UO_7 (O_7,N_4101,N_4284);
or UO_8 (O_8,N_4150,N_4462);
nand UO_9 (O_9,N_4163,N_4487);
nor UO_10 (O_10,N_4814,N_4763);
nand UO_11 (O_11,N_4535,N_4956);
nand UO_12 (O_12,N_4422,N_4465);
or UO_13 (O_13,N_4344,N_4223);
nor UO_14 (O_14,N_4200,N_4933);
or UO_15 (O_15,N_4044,N_4970);
nor UO_16 (O_16,N_4033,N_4474);
nand UO_17 (O_17,N_4983,N_4229);
and UO_18 (O_18,N_4892,N_4592);
xnor UO_19 (O_19,N_4038,N_4713);
nor UO_20 (O_20,N_4475,N_4809);
or UO_21 (O_21,N_4553,N_4283);
and UO_22 (O_22,N_4010,N_4723);
xnor UO_23 (O_23,N_4346,N_4472);
nor UO_24 (O_24,N_4049,N_4749);
nor UO_25 (O_25,N_4595,N_4756);
xor UO_26 (O_26,N_4784,N_4115);
and UO_27 (O_27,N_4483,N_4160);
or UO_28 (O_28,N_4051,N_4254);
and UO_29 (O_29,N_4895,N_4311);
or UO_30 (O_30,N_4159,N_4875);
nand UO_31 (O_31,N_4380,N_4637);
nand UO_32 (O_32,N_4707,N_4816);
xor UO_33 (O_33,N_4011,N_4968);
or UO_34 (O_34,N_4419,N_4665);
and UO_35 (O_35,N_4906,N_4166);
nor UO_36 (O_36,N_4316,N_4812);
or UO_37 (O_37,N_4641,N_4040);
nand UO_38 (O_38,N_4204,N_4025);
and UO_39 (O_39,N_4324,N_4164);
and UO_40 (O_40,N_4512,N_4239);
nand UO_41 (O_41,N_4542,N_4277);
nand UO_42 (O_42,N_4417,N_4959);
nor UO_43 (O_43,N_4338,N_4209);
or UO_44 (O_44,N_4735,N_4696);
and UO_45 (O_45,N_4249,N_4389);
nor UO_46 (O_46,N_4711,N_4184);
nor UO_47 (O_47,N_4515,N_4503);
nand UO_48 (O_48,N_4445,N_4818);
nor UO_49 (O_49,N_4598,N_4815);
xor UO_50 (O_50,N_4618,N_4785);
or UO_51 (O_51,N_4583,N_4729);
xor UO_52 (O_52,N_4568,N_4761);
nor UO_53 (O_53,N_4514,N_4823);
xnor UO_54 (O_54,N_4772,N_4167);
and UO_55 (O_55,N_4221,N_4003);
nor UO_56 (O_56,N_4386,N_4926);
xor UO_57 (O_57,N_4181,N_4786);
xnor UO_58 (O_58,N_4335,N_4725);
nand UO_59 (O_59,N_4456,N_4990);
or UO_60 (O_60,N_4601,N_4098);
nor UO_61 (O_61,N_4278,N_4227);
nand UO_62 (O_62,N_4196,N_4775);
nor UO_63 (O_63,N_4144,N_4234);
and UO_64 (O_64,N_4804,N_4864);
or UO_65 (O_65,N_4647,N_4691);
or UO_66 (O_66,N_4908,N_4332);
nand UO_67 (O_67,N_4082,N_4076);
and UO_68 (O_68,N_4297,N_4479);
and UO_69 (O_69,N_4602,N_4243);
nand UO_70 (O_70,N_4370,N_4416);
and UO_71 (O_71,N_4631,N_4039);
or UO_72 (O_72,N_4799,N_4868);
or UO_73 (O_73,N_4937,N_4915);
nand UO_74 (O_74,N_4710,N_4807);
xor UO_75 (O_75,N_4048,N_4853);
and UO_76 (O_76,N_4174,N_4927);
xnor UO_77 (O_77,N_4310,N_4750);
nand UO_78 (O_78,N_4790,N_4432);
nor UO_79 (O_79,N_4273,N_4436);
and UO_80 (O_80,N_4947,N_4575);
nor UO_81 (O_81,N_4907,N_4973);
or UO_82 (O_82,N_4458,N_4858);
nand UO_83 (O_83,N_4328,N_4849);
and UO_84 (O_84,N_4476,N_4366);
xor UO_85 (O_85,N_4484,N_4766);
nor UO_86 (O_86,N_4700,N_4274);
and UO_87 (O_87,N_4615,N_4492);
or UO_88 (O_88,N_4646,N_4850);
xnor UO_89 (O_89,N_4517,N_4971);
xnor UO_90 (O_90,N_4188,N_4609);
or UO_91 (O_91,N_4326,N_4014);
or UO_92 (O_92,N_4401,N_4097);
and UO_93 (O_93,N_4758,N_4655);
xnor UO_94 (O_94,N_4393,N_4533);
and UO_95 (O_95,N_4275,N_4670);
xnor UO_96 (O_96,N_4315,N_4018);
nand UO_97 (O_97,N_4288,N_4240);
nand UO_98 (O_98,N_4330,N_4720);
nand UO_99 (O_99,N_4726,N_4762);
nand UO_100 (O_100,N_4903,N_4912);
nor UO_101 (O_101,N_4616,N_4803);
xor UO_102 (O_102,N_4950,N_4439);
and UO_103 (O_103,N_4702,N_4813);
and UO_104 (O_104,N_4091,N_4737);
or UO_105 (O_105,N_4360,N_4295);
nor UO_106 (O_106,N_4218,N_4265);
nand UO_107 (O_107,N_4377,N_4177);
and UO_108 (O_108,N_4825,N_4224);
nor UO_109 (O_109,N_4689,N_4337);
nand UO_110 (O_110,N_4651,N_4065);
xnor UO_111 (O_111,N_4543,N_4367);
xnor UO_112 (O_112,N_4427,N_4331);
or UO_113 (O_113,N_4500,N_4420);
xor UO_114 (O_114,N_4605,N_4957);
nand UO_115 (O_115,N_4482,N_4312);
xnor UO_116 (O_116,N_4653,N_4120);
xor UO_117 (O_117,N_4067,N_4920);
nor UO_118 (O_118,N_4534,N_4211);
xnor UO_119 (O_119,N_4153,N_4410);
or UO_120 (O_120,N_4627,N_4658);
nor UO_121 (O_121,N_4888,N_4934);
nand UO_122 (O_122,N_4123,N_4571);
xor UO_123 (O_123,N_4574,N_4373);
and UO_124 (O_124,N_4644,N_4528);
and UO_125 (O_125,N_4020,N_4552);
xor UO_126 (O_126,N_4806,N_4567);
nor UO_127 (O_127,N_4524,N_4536);
nor UO_128 (O_128,N_4576,N_4449);
nand UO_129 (O_129,N_4395,N_4341);
xor UO_130 (O_130,N_4501,N_4801);
xor UO_131 (O_131,N_4760,N_4418);
xnor UO_132 (O_132,N_4506,N_4012);
or UO_133 (O_133,N_4199,N_4885);
nand UO_134 (O_134,N_4245,N_4488);
or UO_135 (O_135,N_4925,N_4064);
nor UO_136 (O_136,N_4250,N_4382);
nor UO_137 (O_137,N_4596,N_4185);
or UO_138 (O_138,N_4860,N_4997);
and UO_139 (O_139,N_4149,N_4485);
nand UO_140 (O_140,N_4917,N_4563);
nand UO_141 (O_141,N_4736,N_4024);
xor UO_142 (O_142,N_4588,N_4727);
xnor UO_143 (O_143,N_4198,N_4015);
xor UO_144 (O_144,N_4448,N_4403);
xnor UO_145 (O_145,N_4113,N_4960);
nor UO_146 (O_146,N_4043,N_4969);
nor UO_147 (O_147,N_4954,N_4028);
nor UO_148 (O_148,N_4792,N_4699);
and UO_149 (O_149,N_4182,N_4765);
and UO_150 (O_150,N_4509,N_4179);
or UO_151 (O_151,N_4016,N_4292);
and UO_152 (O_152,N_4294,N_4610);
or UO_153 (O_153,N_4408,N_4964);
or UO_154 (O_154,N_4491,N_4347);
and UO_155 (O_155,N_4352,N_4554);
xnor UO_156 (O_156,N_4397,N_4222);
or UO_157 (O_157,N_4638,N_4137);
xor UO_158 (O_158,N_4489,N_4220);
nand UO_159 (O_159,N_4780,N_4027);
xor UO_160 (O_160,N_4837,N_4267);
xnor UO_161 (O_161,N_4752,N_4683);
nand UO_162 (O_162,N_4572,N_4923);
or UO_163 (O_163,N_4963,N_4624);
nand UO_164 (O_164,N_4998,N_4833);
xnor UO_165 (O_165,N_4186,N_4276);
nand UO_166 (O_166,N_4755,N_4890);
or UO_167 (O_167,N_4384,N_4302);
xnor UO_168 (O_168,N_4077,N_4207);
nand UO_169 (O_169,N_4935,N_4244);
and UO_170 (O_170,N_4272,N_4680);
and UO_171 (O_171,N_4090,N_4452);
nor UO_172 (O_172,N_4074,N_4949);
nor UO_173 (O_173,N_4879,N_4363);
nand UO_174 (O_174,N_4891,N_4687);
or UO_175 (O_175,N_4991,N_4241);
and UO_176 (O_176,N_4431,N_4168);
xor UO_177 (O_177,N_4883,N_4495);
nor UO_178 (O_178,N_4505,N_4928);
nand UO_179 (O_179,N_4771,N_4866);
and UO_180 (O_180,N_4381,N_4261);
nand UO_181 (O_181,N_4037,N_4733);
or UO_182 (O_182,N_4424,N_4371);
nor UO_183 (O_183,N_4652,N_4108);
nor UO_184 (O_184,N_4429,N_4642);
and UO_185 (O_185,N_4414,N_4197);
or UO_186 (O_186,N_4394,N_4544);
nor UO_187 (O_187,N_4939,N_4719);
and UO_188 (O_188,N_4682,N_4820);
nand UO_189 (O_189,N_4805,N_4550);
or UO_190 (O_190,N_4876,N_4821);
or UO_191 (O_191,N_4231,N_4769);
xor UO_192 (O_192,N_4320,N_4791);
xnor UO_193 (O_193,N_4390,N_4190);
xor UO_194 (O_194,N_4004,N_4191);
or UO_195 (O_195,N_4260,N_4158);
nor UO_196 (O_196,N_4387,N_4477);
nor UO_197 (O_197,N_4654,N_4802);
or UO_198 (O_198,N_4661,N_4839);
or UO_199 (O_199,N_4532,N_4841);
nor UO_200 (O_200,N_4604,N_4035);
nor UO_201 (O_201,N_4425,N_4659);
nor UO_202 (O_202,N_4777,N_4561);
nand UO_203 (O_203,N_4455,N_4834);
xnor UO_204 (O_204,N_4731,N_4444);
nand UO_205 (O_205,N_4754,N_4021);
or UO_206 (O_206,N_4882,N_4832);
nand UO_207 (O_207,N_4175,N_4753);
and UO_208 (O_208,N_4636,N_4135);
xor UO_209 (O_209,N_4856,N_4600);
or UO_210 (O_210,N_4225,N_4523);
and UO_211 (O_211,N_4840,N_4046);
nor UO_212 (O_212,N_4442,N_4447);
xor UO_213 (O_213,N_4413,N_4466);
nand UO_214 (O_214,N_4092,N_4900);
or UO_215 (O_215,N_4263,N_4541);
xor UO_216 (O_216,N_4518,N_4857);
nor UO_217 (O_217,N_4759,N_4287);
and UO_218 (O_218,N_4103,N_4111);
nand UO_219 (O_219,N_4171,N_4694);
nor UO_220 (O_220,N_4649,N_4635);
nor UO_221 (O_221,N_4264,N_4214);
nor UO_222 (O_222,N_4105,N_4606);
or UO_223 (O_223,N_4728,N_4936);
and UO_224 (O_224,N_4996,N_4955);
nand UO_225 (O_225,N_4121,N_4388);
or UO_226 (O_226,N_4742,N_4904);
nor UO_227 (O_227,N_4846,N_4952);
xnor UO_228 (O_228,N_4268,N_4102);
nand UO_229 (O_229,N_4613,N_4918);
or UO_230 (O_230,N_4675,N_4704);
and UO_231 (O_231,N_4869,N_4593);
xnor UO_232 (O_232,N_4086,N_4855);
nor UO_233 (O_233,N_4392,N_4862);
xnor UO_234 (O_234,N_4141,N_4994);
and UO_235 (O_235,N_4146,N_4938);
or UO_236 (O_236,N_4083,N_4705);
and UO_237 (O_237,N_4189,N_4573);
or UO_238 (O_238,N_4826,N_4851);
nand UO_239 (O_239,N_4607,N_4006);
nand UO_240 (O_240,N_4339,N_4486);
and UO_241 (O_241,N_4995,N_4434);
or UO_242 (O_242,N_4348,N_4162);
and UO_243 (O_243,N_4002,N_4376);
nor UO_244 (O_244,N_4819,N_4664);
nor UO_245 (O_245,N_4831,N_4537);
nor UO_246 (O_246,N_4139,N_4504);
nand UO_247 (O_247,N_4365,N_4143);
nor UO_248 (O_248,N_4560,N_4527);
and UO_249 (O_249,N_4865,N_4581);
xnor UO_250 (O_250,N_4611,N_4496);
nand UO_251 (O_251,N_4421,N_4075);
nand UO_252 (O_252,N_4256,N_4824);
or UO_253 (O_253,N_4842,N_4800);
xor UO_254 (O_254,N_4570,N_4467);
xnor UO_255 (O_255,N_4859,N_4986);
or UO_256 (O_256,N_4230,N_4678);
or UO_257 (O_257,N_4697,N_4122);
nor UO_258 (O_258,N_4612,N_4404);
xor UO_259 (O_259,N_4258,N_4867);
nor UO_260 (O_260,N_4650,N_4280);
xor UO_261 (O_261,N_4585,N_4169);
xor UO_262 (O_262,N_4525,N_4172);
and UO_263 (O_263,N_4718,N_4242);
nand UO_264 (O_264,N_4978,N_4872);
nor UO_265 (O_265,N_4481,N_4236);
nand UO_266 (O_266,N_4099,N_4126);
or UO_267 (O_267,N_4531,N_4657);
nand UO_268 (O_268,N_4291,N_4402);
nand UO_269 (O_269,N_4253,N_4133);
nor UO_270 (O_270,N_4690,N_4835);
nor UO_271 (O_271,N_4453,N_4714);
xnor UO_272 (O_272,N_4881,N_4929);
or UO_273 (O_273,N_4019,N_4999);
and UO_274 (O_274,N_4548,N_4454);
and UO_275 (O_275,N_4559,N_4178);
or UO_276 (O_276,N_4134,N_4982);
or UO_277 (O_277,N_4180,N_4473);
or UO_278 (O_278,N_4345,N_4887);
nor UO_279 (O_279,N_4944,N_4406);
nor UO_280 (O_280,N_4237,N_4539);
nor UO_281 (O_281,N_4490,N_4361);
nand UO_282 (O_282,N_4112,N_4958);
or UO_283 (O_283,N_4088,N_4993);
xnor UO_284 (O_284,N_4461,N_4157);
nor UO_285 (O_285,N_4068,N_4564);
nand UO_286 (O_286,N_4358,N_4587);
xnor UO_287 (O_287,N_4464,N_4679);
and UO_288 (O_288,N_4746,N_4087);
or UO_289 (O_289,N_4838,N_4125);
xnor UO_290 (O_290,N_4216,N_4693);
nand UO_291 (O_291,N_4362,N_4235);
nand UO_292 (O_292,N_4364,N_4206);
nand UO_293 (O_293,N_4708,N_4577);
xnor UO_294 (O_294,N_4247,N_4201);
nand UO_295 (O_295,N_4943,N_4961);
nor UO_296 (O_296,N_4545,N_4562);
and UO_297 (O_297,N_4692,N_4329);
or UO_298 (O_298,N_4219,N_4036);
or UO_299 (O_299,N_4407,N_4089);
nor UO_300 (O_300,N_4972,N_4079);
nor UO_301 (O_301,N_4323,N_4811);
or UO_302 (O_302,N_4194,N_4730);
nand UO_303 (O_303,N_4632,N_4673);
nand UO_304 (O_304,N_4050,N_4980);
or UO_305 (O_305,N_4138,N_4305);
and UO_306 (O_306,N_4547,N_4057);
and UO_307 (O_307,N_4989,N_4794);
nor UO_308 (O_308,N_4584,N_4822);
nand UO_309 (O_309,N_4405,N_4001);
nor UO_310 (O_310,N_4617,N_4142);
or UO_311 (O_311,N_4176,N_4210);
nand UO_312 (O_312,N_4000,N_4745);
or UO_313 (O_313,N_4529,N_4671);
nor UO_314 (O_314,N_4639,N_4266);
or UO_315 (O_315,N_4469,N_4976);
nand UO_316 (O_316,N_4896,N_4007);
nor UO_317 (O_317,N_4498,N_4586);
or UO_318 (O_318,N_4228,N_4217);
nor UO_319 (O_319,N_4783,N_4965);
or UO_320 (O_320,N_4070,N_4880);
or UO_321 (O_321,N_4289,N_4154);
nand UO_322 (O_322,N_4286,N_4147);
or UO_323 (O_323,N_4748,N_4977);
or UO_324 (O_324,N_4032,N_4298);
xor UO_325 (O_325,N_4318,N_4941);
and UO_326 (O_326,N_4359,N_4597);
and UO_327 (O_327,N_4252,N_4852);
nor UO_328 (O_328,N_4457,N_4913);
nand UO_329 (O_329,N_4668,N_4546);
and UO_330 (O_330,N_4396,N_4279);
nand UO_331 (O_331,N_4340,N_4828);
and UO_332 (O_332,N_4282,N_4281);
xnor UO_333 (O_333,N_4676,N_4556);
xnor UO_334 (O_334,N_4321,N_4423);
and UO_335 (O_335,N_4688,N_4441);
nand UO_336 (O_336,N_4170,N_4470);
or UO_337 (O_337,N_4910,N_4357);
nand UO_338 (O_338,N_4059,N_4619);
xnor UO_339 (O_339,N_4966,N_4873);
and UO_340 (O_340,N_4349,N_4871);
and UO_341 (O_341,N_4368,N_4764);
or UO_342 (O_342,N_4334,N_4902);
and UO_343 (O_343,N_4152,N_4757);
nand UO_344 (O_344,N_4056,N_4930);
xor UO_345 (O_345,N_4681,N_4626);
nor UO_346 (O_346,N_4921,N_4127);
and UO_347 (O_347,N_4041,N_4981);
and UO_348 (O_348,N_4732,N_4080);
nand UO_349 (O_349,N_4580,N_4478);
nand UO_350 (O_350,N_4129,N_4148);
xnor UO_351 (O_351,N_4540,N_4155);
or UO_352 (O_352,N_4594,N_4031);
nor UO_353 (O_353,N_4795,N_4717);
or UO_354 (O_354,N_4914,N_4005);
and UO_355 (O_355,N_4307,N_4435);
xnor UO_356 (O_356,N_4712,N_4569);
nand UO_357 (O_357,N_4459,N_4614);
nor UO_358 (O_358,N_4052,N_4590);
xor UO_359 (O_359,N_4262,N_4428);
or UO_360 (O_360,N_4911,N_4055);
nand UO_361 (O_361,N_4270,N_4847);
nand UO_362 (O_362,N_4640,N_4513);
nor UO_363 (O_363,N_4589,N_4106);
or UO_364 (O_364,N_4124,N_4034);
nand UO_365 (O_365,N_4116,N_4591);
nor UO_366 (O_366,N_4660,N_4674);
nand UO_367 (O_367,N_4743,N_4356);
and UO_368 (O_368,N_4029,N_4095);
nor UO_369 (O_369,N_4212,N_4426);
nand UO_370 (O_370,N_4383,N_4248);
and UO_371 (O_371,N_4085,N_4299);
nand UO_372 (O_372,N_4603,N_4629);
nor UO_373 (O_373,N_4656,N_4238);
xnor UO_374 (O_374,N_4399,N_4100);
and UO_375 (O_375,N_4739,N_4450);
or UO_376 (O_376,N_4740,N_4355);
and UO_377 (O_377,N_4433,N_4202);
nand UO_378 (O_378,N_4317,N_4817);
nand UO_379 (O_379,N_4333,N_4770);
nor UO_380 (O_380,N_4165,N_4026);
xor UO_381 (O_381,N_4919,N_4372);
nor UO_382 (O_382,N_4984,N_4130);
nand UO_383 (O_383,N_4829,N_4716);
nand UO_384 (O_384,N_4107,N_4257);
or UO_385 (O_385,N_4945,N_4599);
nor UO_386 (O_386,N_4565,N_4136);
nor UO_387 (O_387,N_4053,N_4412);
nand UO_388 (O_388,N_4350,N_4843);
nor UO_389 (O_389,N_4667,N_4669);
or UO_390 (O_390,N_4507,N_4030);
nor UO_391 (O_391,N_4259,N_4686);
xnor UO_392 (O_392,N_4663,N_4620);
nor UO_393 (O_393,N_4411,N_4854);
and UO_394 (O_394,N_4797,N_4430);
xnor UO_395 (O_395,N_4516,N_4768);
nand UO_396 (O_396,N_4008,N_4830);
nor UO_397 (O_397,N_4520,N_4798);
nand UO_398 (O_398,N_4375,N_4508);
xnor UO_399 (O_399,N_4415,N_4905);
or UO_400 (O_400,N_4861,N_4269);
or UO_401 (O_401,N_4063,N_4314);
or UO_402 (O_402,N_4023,N_4071);
nand UO_403 (O_403,N_4974,N_4118);
xor UO_404 (O_404,N_4932,N_4521);
and UO_405 (O_405,N_4140,N_4979);
or UO_406 (O_406,N_4931,N_4622);
nor UO_407 (O_407,N_4848,N_4555);
and UO_408 (O_408,N_4893,N_4870);
xnor UO_409 (O_409,N_4566,N_4400);
and UO_410 (O_410,N_4899,N_4884);
xnor UO_411 (O_411,N_4379,N_4303);
nor UO_412 (O_412,N_4625,N_4827);
nor UO_413 (O_413,N_4579,N_4354);
and UO_414 (O_414,N_4721,N_4342);
xnor UO_415 (O_415,N_4096,N_4510);
nand UO_416 (O_416,N_4192,N_4378);
xor UO_417 (O_417,N_4538,N_4463);
or UO_418 (O_418,N_4987,N_4131);
xnor UO_419 (O_419,N_4962,N_4215);
xor UO_420 (O_420,N_4066,N_4183);
nand UO_421 (O_421,N_4774,N_4151);
xor UO_422 (O_422,N_4145,N_4351);
nand UO_423 (O_423,N_4013,N_4988);
xor UO_424 (O_424,N_4722,N_4078);
xnor UO_425 (O_425,N_4119,N_4336);
and UO_426 (O_426,N_4073,N_4877);
nand UO_427 (O_427,N_4084,N_4940);
xnor UO_428 (O_428,N_4810,N_4634);
nor UO_429 (O_429,N_4643,N_4985);
xor UO_430 (O_430,N_4409,N_4738);
or UO_431 (O_431,N_4787,N_4385);
xor UO_432 (O_432,N_4781,N_4499);
and UO_433 (O_433,N_4203,N_4301);
xnor UO_434 (O_434,N_4042,N_4789);
or UO_435 (O_435,N_4782,N_4114);
nor UO_436 (O_436,N_4557,N_4916);
or UO_437 (O_437,N_4069,N_4703);
and UO_438 (O_438,N_4440,N_4698);
nand UO_439 (O_439,N_4666,N_4578);
nor UO_440 (O_440,N_4951,N_4391);
nor UO_441 (O_441,N_4468,N_4497);
or UO_442 (O_442,N_4208,N_4744);
and UO_443 (O_443,N_4117,N_4886);
xor UO_444 (O_444,N_4773,N_4246);
nor UO_445 (O_445,N_4161,N_4975);
nor UO_446 (O_446,N_4844,N_4793);
nand UO_447 (O_447,N_4551,N_4709);
nor UO_448 (O_448,N_4608,N_4889);
or UO_449 (O_449,N_4309,N_4924);
nand UO_450 (O_450,N_4226,N_4128);
xor UO_451 (O_451,N_4327,N_4110);
nand UO_452 (O_452,N_4271,N_4621);
xnor UO_453 (O_453,N_4526,N_4480);
and UO_454 (O_454,N_4094,N_4062);
and UO_455 (O_455,N_4648,N_4845);
or UO_456 (O_456,N_4522,N_4104);
or UO_457 (O_457,N_4662,N_4779);
or UO_458 (O_458,N_4874,N_4623);
and UO_459 (O_459,N_4285,N_4374);
nand UO_460 (O_460,N_4878,N_4685);
nand UO_461 (O_461,N_4061,N_4894);
nand UO_462 (O_462,N_4081,N_4897);
or UO_463 (O_463,N_4695,N_4741);
nor UO_464 (O_464,N_4306,N_4942);
or UO_465 (O_465,N_4582,N_4058);
nand UO_466 (O_466,N_4778,N_4558);
or UO_467 (O_467,N_4398,N_4808);
nor UO_468 (O_468,N_4132,N_4313);
or UO_469 (O_469,N_4296,N_4369);
nor UO_470 (O_470,N_4630,N_4322);
and UO_471 (O_471,N_4308,N_4093);
or UO_472 (O_472,N_4645,N_4045);
nand UO_473 (O_473,N_4909,N_4195);
nand UO_474 (O_474,N_4251,N_4460);
nand UO_475 (O_475,N_4549,N_4747);
and UO_476 (O_476,N_4511,N_4232);
and UO_477 (O_477,N_4193,N_4767);
nor UO_478 (O_478,N_4724,N_4672);
or UO_479 (O_479,N_4922,N_4233);
nor UO_480 (O_480,N_4054,N_4901);
xnor UO_481 (O_481,N_4446,N_4706);
xor UO_482 (O_482,N_4633,N_4734);
and UO_483 (O_483,N_4898,N_4751);
xnor UO_484 (O_484,N_4205,N_4471);
and UO_485 (O_485,N_4325,N_4060);
or UO_486 (O_486,N_4109,N_4530);
or UO_487 (O_487,N_4255,N_4300);
or UO_488 (O_488,N_4443,N_4156);
nor UO_489 (O_489,N_4946,N_4796);
and UO_490 (O_490,N_4628,N_4304);
nor UO_491 (O_491,N_4213,N_4438);
and UO_492 (O_492,N_4319,N_4072);
nand UO_493 (O_493,N_4677,N_4715);
nor UO_494 (O_494,N_4948,N_4502);
nor UO_495 (O_495,N_4173,N_4022);
or UO_496 (O_496,N_4836,N_4788);
and UO_497 (O_497,N_4494,N_4353);
nand UO_498 (O_498,N_4684,N_4776);
nand UO_499 (O_499,N_4992,N_4009);
or UO_500 (O_500,N_4313,N_4037);
or UO_501 (O_501,N_4774,N_4939);
xor UO_502 (O_502,N_4908,N_4285);
or UO_503 (O_503,N_4157,N_4752);
nor UO_504 (O_504,N_4949,N_4775);
or UO_505 (O_505,N_4876,N_4597);
nor UO_506 (O_506,N_4908,N_4675);
or UO_507 (O_507,N_4536,N_4773);
nor UO_508 (O_508,N_4081,N_4303);
xnor UO_509 (O_509,N_4403,N_4309);
and UO_510 (O_510,N_4814,N_4355);
and UO_511 (O_511,N_4200,N_4983);
xor UO_512 (O_512,N_4303,N_4572);
nand UO_513 (O_513,N_4102,N_4149);
nand UO_514 (O_514,N_4691,N_4604);
nor UO_515 (O_515,N_4142,N_4174);
nor UO_516 (O_516,N_4674,N_4796);
nand UO_517 (O_517,N_4295,N_4069);
or UO_518 (O_518,N_4083,N_4103);
xor UO_519 (O_519,N_4901,N_4178);
or UO_520 (O_520,N_4364,N_4887);
or UO_521 (O_521,N_4702,N_4751);
nand UO_522 (O_522,N_4309,N_4698);
nor UO_523 (O_523,N_4829,N_4288);
and UO_524 (O_524,N_4962,N_4577);
and UO_525 (O_525,N_4634,N_4100);
or UO_526 (O_526,N_4303,N_4789);
and UO_527 (O_527,N_4578,N_4702);
and UO_528 (O_528,N_4690,N_4949);
nor UO_529 (O_529,N_4309,N_4591);
or UO_530 (O_530,N_4787,N_4950);
nand UO_531 (O_531,N_4128,N_4612);
or UO_532 (O_532,N_4411,N_4439);
or UO_533 (O_533,N_4097,N_4996);
or UO_534 (O_534,N_4518,N_4236);
nand UO_535 (O_535,N_4571,N_4839);
nor UO_536 (O_536,N_4250,N_4530);
nand UO_537 (O_537,N_4269,N_4420);
xor UO_538 (O_538,N_4008,N_4218);
or UO_539 (O_539,N_4584,N_4266);
or UO_540 (O_540,N_4463,N_4433);
xor UO_541 (O_541,N_4950,N_4877);
nand UO_542 (O_542,N_4343,N_4134);
xnor UO_543 (O_543,N_4214,N_4881);
nand UO_544 (O_544,N_4605,N_4117);
nor UO_545 (O_545,N_4452,N_4119);
xnor UO_546 (O_546,N_4516,N_4263);
and UO_547 (O_547,N_4056,N_4326);
nand UO_548 (O_548,N_4578,N_4807);
nor UO_549 (O_549,N_4189,N_4896);
or UO_550 (O_550,N_4652,N_4323);
and UO_551 (O_551,N_4062,N_4082);
nor UO_552 (O_552,N_4067,N_4629);
and UO_553 (O_553,N_4287,N_4101);
nand UO_554 (O_554,N_4782,N_4195);
or UO_555 (O_555,N_4681,N_4283);
or UO_556 (O_556,N_4252,N_4487);
nand UO_557 (O_557,N_4139,N_4686);
and UO_558 (O_558,N_4187,N_4840);
nor UO_559 (O_559,N_4172,N_4529);
and UO_560 (O_560,N_4427,N_4831);
xor UO_561 (O_561,N_4029,N_4438);
nor UO_562 (O_562,N_4397,N_4381);
or UO_563 (O_563,N_4818,N_4299);
and UO_564 (O_564,N_4981,N_4442);
and UO_565 (O_565,N_4445,N_4449);
nand UO_566 (O_566,N_4098,N_4921);
or UO_567 (O_567,N_4507,N_4518);
xnor UO_568 (O_568,N_4801,N_4440);
xor UO_569 (O_569,N_4272,N_4790);
or UO_570 (O_570,N_4558,N_4324);
nor UO_571 (O_571,N_4545,N_4121);
or UO_572 (O_572,N_4314,N_4774);
nand UO_573 (O_573,N_4178,N_4286);
nand UO_574 (O_574,N_4750,N_4249);
nor UO_575 (O_575,N_4584,N_4369);
xnor UO_576 (O_576,N_4962,N_4388);
nor UO_577 (O_577,N_4737,N_4495);
xor UO_578 (O_578,N_4629,N_4695);
nand UO_579 (O_579,N_4816,N_4549);
xnor UO_580 (O_580,N_4521,N_4785);
nand UO_581 (O_581,N_4938,N_4814);
and UO_582 (O_582,N_4777,N_4789);
and UO_583 (O_583,N_4089,N_4387);
nor UO_584 (O_584,N_4443,N_4105);
nand UO_585 (O_585,N_4779,N_4814);
nand UO_586 (O_586,N_4817,N_4587);
and UO_587 (O_587,N_4343,N_4863);
nand UO_588 (O_588,N_4465,N_4074);
nand UO_589 (O_589,N_4888,N_4413);
xnor UO_590 (O_590,N_4508,N_4822);
or UO_591 (O_591,N_4772,N_4513);
xor UO_592 (O_592,N_4103,N_4433);
nand UO_593 (O_593,N_4248,N_4075);
or UO_594 (O_594,N_4773,N_4718);
nand UO_595 (O_595,N_4219,N_4090);
nor UO_596 (O_596,N_4276,N_4809);
or UO_597 (O_597,N_4654,N_4121);
and UO_598 (O_598,N_4971,N_4231);
nor UO_599 (O_599,N_4214,N_4955);
nand UO_600 (O_600,N_4626,N_4062);
nand UO_601 (O_601,N_4020,N_4219);
nor UO_602 (O_602,N_4659,N_4523);
nor UO_603 (O_603,N_4003,N_4608);
nor UO_604 (O_604,N_4717,N_4980);
nor UO_605 (O_605,N_4842,N_4398);
nor UO_606 (O_606,N_4704,N_4797);
xnor UO_607 (O_607,N_4741,N_4781);
nor UO_608 (O_608,N_4455,N_4435);
xor UO_609 (O_609,N_4177,N_4116);
and UO_610 (O_610,N_4988,N_4910);
xor UO_611 (O_611,N_4419,N_4440);
nor UO_612 (O_612,N_4260,N_4021);
and UO_613 (O_613,N_4413,N_4217);
nor UO_614 (O_614,N_4254,N_4549);
nor UO_615 (O_615,N_4786,N_4277);
and UO_616 (O_616,N_4347,N_4544);
and UO_617 (O_617,N_4142,N_4555);
or UO_618 (O_618,N_4105,N_4514);
nor UO_619 (O_619,N_4851,N_4264);
nor UO_620 (O_620,N_4478,N_4681);
xnor UO_621 (O_621,N_4221,N_4611);
or UO_622 (O_622,N_4592,N_4991);
or UO_623 (O_623,N_4554,N_4607);
and UO_624 (O_624,N_4485,N_4722);
nor UO_625 (O_625,N_4715,N_4714);
or UO_626 (O_626,N_4600,N_4563);
and UO_627 (O_627,N_4166,N_4410);
and UO_628 (O_628,N_4104,N_4570);
nor UO_629 (O_629,N_4171,N_4504);
nor UO_630 (O_630,N_4298,N_4439);
and UO_631 (O_631,N_4463,N_4142);
nor UO_632 (O_632,N_4219,N_4335);
nand UO_633 (O_633,N_4298,N_4161);
nor UO_634 (O_634,N_4637,N_4562);
nand UO_635 (O_635,N_4615,N_4658);
or UO_636 (O_636,N_4427,N_4745);
nand UO_637 (O_637,N_4814,N_4669);
and UO_638 (O_638,N_4536,N_4243);
nor UO_639 (O_639,N_4330,N_4723);
nand UO_640 (O_640,N_4470,N_4831);
nand UO_641 (O_641,N_4036,N_4519);
and UO_642 (O_642,N_4153,N_4074);
and UO_643 (O_643,N_4972,N_4213);
or UO_644 (O_644,N_4111,N_4194);
and UO_645 (O_645,N_4720,N_4834);
and UO_646 (O_646,N_4508,N_4836);
and UO_647 (O_647,N_4832,N_4867);
and UO_648 (O_648,N_4063,N_4624);
nor UO_649 (O_649,N_4526,N_4709);
or UO_650 (O_650,N_4197,N_4250);
xnor UO_651 (O_651,N_4757,N_4066);
nor UO_652 (O_652,N_4267,N_4790);
or UO_653 (O_653,N_4189,N_4601);
or UO_654 (O_654,N_4713,N_4559);
nand UO_655 (O_655,N_4190,N_4623);
xnor UO_656 (O_656,N_4582,N_4335);
nand UO_657 (O_657,N_4891,N_4820);
and UO_658 (O_658,N_4008,N_4303);
nand UO_659 (O_659,N_4704,N_4985);
nand UO_660 (O_660,N_4296,N_4400);
nor UO_661 (O_661,N_4337,N_4339);
nand UO_662 (O_662,N_4355,N_4016);
nand UO_663 (O_663,N_4614,N_4892);
and UO_664 (O_664,N_4579,N_4192);
nor UO_665 (O_665,N_4504,N_4967);
or UO_666 (O_666,N_4850,N_4505);
nor UO_667 (O_667,N_4294,N_4307);
and UO_668 (O_668,N_4526,N_4242);
and UO_669 (O_669,N_4508,N_4166);
and UO_670 (O_670,N_4709,N_4193);
xnor UO_671 (O_671,N_4544,N_4060);
nor UO_672 (O_672,N_4847,N_4839);
and UO_673 (O_673,N_4934,N_4287);
nor UO_674 (O_674,N_4300,N_4095);
or UO_675 (O_675,N_4542,N_4991);
xnor UO_676 (O_676,N_4388,N_4481);
nand UO_677 (O_677,N_4015,N_4549);
xnor UO_678 (O_678,N_4466,N_4338);
xor UO_679 (O_679,N_4374,N_4385);
xor UO_680 (O_680,N_4920,N_4440);
xor UO_681 (O_681,N_4813,N_4295);
or UO_682 (O_682,N_4006,N_4917);
nor UO_683 (O_683,N_4360,N_4202);
nand UO_684 (O_684,N_4608,N_4052);
and UO_685 (O_685,N_4222,N_4826);
and UO_686 (O_686,N_4839,N_4173);
xor UO_687 (O_687,N_4085,N_4122);
xnor UO_688 (O_688,N_4577,N_4423);
xnor UO_689 (O_689,N_4112,N_4298);
or UO_690 (O_690,N_4774,N_4660);
or UO_691 (O_691,N_4397,N_4042);
nor UO_692 (O_692,N_4683,N_4550);
nor UO_693 (O_693,N_4916,N_4626);
nand UO_694 (O_694,N_4522,N_4907);
or UO_695 (O_695,N_4115,N_4761);
xnor UO_696 (O_696,N_4493,N_4139);
and UO_697 (O_697,N_4925,N_4400);
or UO_698 (O_698,N_4531,N_4277);
or UO_699 (O_699,N_4247,N_4297);
or UO_700 (O_700,N_4742,N_4602);
or UO_701 (O_701,N_4800,N_4487);
or UO_702 (O_702,N_4742,N_4032);
xor UO_703 (O_703,N_4931,N_4025);
or UO_704 (O_704,N_4419,N_4313);
xnor UO_705 (O_705,N_4869,N_4473);
or UO_706 (O_706,N_4386,N_4283);
xnor UO_707 (O_707,N_4658,N_4580);
and UO_708 (O_708,N_4754,N_4234);
or UO_709 (O_709,N_4130,N_4041);
and UO_710 (O_710,N_4783,N_4493);
or UO_711 (O_711,N_4911,N_4615);
nor UO_712 (O_712,N_4529,N_4200);
nor UO_713 (O_713,N_4524,N_4364);
nand UO_714 (O_714,N_4881,N_4986);
nor UO_715 (O_715,N_4539,N_4649);
xor UO_716 (O_716,N_4978,N_4239);
nor UO_717 (O_717,N_4061,N_4528);
nor UO_718 (O_718,N_4599,N_4743);
or UO_719 (O_719,N_4331,N_4210);
nand UO_720 (O_720,N_4884,N_4461);
xor UO_721 (O_721,N_4083,N_4730);
nor UO_722 (O_722,N_4001,N_4846);
xnor UO_723 (O_723,N_4474,N_4404);
and UO_724 (O_724,N_4792,N_4905);
or UO_725 (O_725,N_4341,N_4706);
or UO_726 (O_726,N_4304,N_4940);
xor UO_727 (O_727,N_4958,N_4975);
nand UO_728 (O_728,N_4068,N_4495);
nand UO_729 (O_729,N_4896,N_4158);
nor UO_730 (O_730,N_4002,N_4895);
nand UO_731 (O_731,N_4939,N_4280);
nand UO_732 (O_732,N_4215,N_4816);
nor UO_733 (O_733,N_4986,N_4588);
or UO_734 (O_734,N_4677,N_4834);
nand UO_735 (O_735,N_4836,N_4642);
nand UO_736 (O_736,N_4092,N_4761);
nand UO_737 (O_737,N_4470,N_4370);
nor UO_738 (O_738,N_4179,N_4706);
or UO_739 (O_739,N_4185,N_4898);
xnor UO_740 (O_740,N_4176,N_4864);
xnor UO_741 (O_741,N_4570,N_4973);
xnor UO_742 (O_742,N_4895,N_4249);
xnor UO_743 (O_743,N_4906,N_4536);
nand UO_744 (O_744,N_4779,N_4460);
xnor UO_745 (O_745,N_4703,N_4839);
and UO_746 (O_746,N_4559,N_4762);
or UO_747 (O_747,N_4465,N_4591);
or UO_748 (O_748,N_4857,N_4532);
or UO_749 (O_749,N_4421,N_4247);
xor UO_750 (O_750,N_4589,N_4810);
or UO_751 (O_751,N_4971,N_4198);
xnor UO_752 (O_752,N_4364,N_4049);
nand UO_753 (O_753,N_4539,N_4409);
and UO_754 (O_754,N_4198,N_4274);
or UO_755 (O_755,N_4182,N_4502);
and UO_756 (O_756,N_4085,N_4448);
nor UO_757 (O_757,N_4437,N_4518);
xnor UO_758 (O_758,N_4686,N_4547);
nand UO_759 (O_759,N_4094,N_4900);
or UO_760 (O_760,N_4454,N_4967);
and UO_761 (O_761,N_4372,N_4222);
or UO_762 (O_762,N_4319,N_4047);
nand UO_763 (O_763,N_4455,N_4290);
nor UO_764 (O_764,N_4640,N_4182);
or UO_765 (O_765,N_4527,N_4932);
nand UO_766 (O_766,N_4199,N_4044);
xor UO_767 (O_767,N_4331,N_4929);
xor UO_768 (O_768,N_4271,N_4423);
or UO_769 (O_769,N_4951,N_4139);
nand UO_770 (O_770,N_4474,N_4065);
xor UO_771 (O_771,N_4014,N_4663);
xor UO_772 (O_772,N_4354,N_4590);
nand UO_773 (O_773,N_4479,N_4336);
nand UO_774 (O_774,N_4910,N_4583);
nor UO_775 (O_775,N_4352,N_4943);
and UO_776 (O_776,N_4622,N_4918);
xor UO_777 (O_777,N_4761,N_4228);
nand UO_778 (O_778,N_4488,N_4093);
or UO_779 (O_779,N_4640,N_4273);
nor UO_780 (O_780,N_4081,N_4871);
nand UO_781 (O_781,N_4770,N_4755);
xor UO_782 (O_782,N_4266,N_4493);
nor UO_783 (O_783,N_4262,N_4869);
xnor UO_784 (O_784,N_4262,N_4903);
xor UO_785 (O_785,N_4149,N_4458);
nand UO_786 (O_786,N_4855,N_4704);
and UO_787 (O_787,N_4699,N_4568);
nor UO_788 (O_788,N_4523,N_4637);
nand UO_789 (O_789,N_4689,N_4460);
and UO_790 (O_790,N_4073,N_4353);
and UO_791 (O_791,N_4796,N_4537);
nor UO_792 (O_792,N_4661,N_4464);
xor UO_793 (O_793,N_4502,N_4000);
nor UO_794 (O_794,N_4631,N_4187);
and UO_795 (O_795,N_4670,N_4970);
and UO_796 (O_796,N_4595,N_4990);
and UO_797 (O_797,N_4258,N_4938);
xor UO_798 (O_798,N_4601,N_4996);
or UO_799 (O_799,N_4230,N_4451);
nand UO_800 (O_800,N_4438,N_4620);
nor UO_801 (O_801,N_4571,N_4562);
nand UO_802 (O_802,N_4524,N_4735);
nand UO_803 (O_803,N_4089,N_4032);
xor UO_804 (O_804,N_4892,N_4499);
or UO_805 (O_805,N_4085,N_4892);
nand UO_806 (O_806,N_4464,N_4264);
nand UO_807 (O_807,N_4396,N_4930);
xnor UO_808 (O_808,N_4574,N_4231);
xor UO_809 (O_809,N_4887,N_4758);
and UO_810 (O_810,N_4099,N_4220);
or UO_811 (O_811,N_4939,N_4604);
or UO_812 (O_812,N_4752,N_4090);
nand UO_813 (O_813,N_4183,N_4648);
or UO_814 (O_814,N_4212,N_4180);
nand UO_815 (O_815,N_4431,N_4779);
or UO_816 (O_816,N_4406,N_4703);
and UO_817 (O_817,N_4617,N_4957);
nand UO_818 (O_818,N_4908,N_4280);
and UO_819 (O_819,N_4094,N_4636);
nand UO_820 (O_820,N_4517,N_4015);
or UO_821 (O_821,N_4663,N_4878);
and UO_822 (O_822,N_4097,N_4462);
nand UO_823 (O_823,N_4703,N_4606);
nor UO_824 (O_824,N_4769,N_4911);
xor UO_825 (O_825,N_4119,N_4662);
nor UO_826 (O_826,N_4505,N_4036);
and UO_827 (O_827,N_4458,N_4659);
nand UO_828 (O_828,N_4872,N_4073);
nor UO_829 (O_829,N_4047,N_4005);
nor UO_830 (O_830,N_4368,N_4050);
nor UO_831 (O_831,N_4636,N_4459);
xnor UO_832 (O_832,N_4559,N_4486);
xor UO_833 (O_833,N_4580,N_4344);
xnor UO_834 (O_834,N_4002,N_4824);
nand UO_835 (O_835,N_4045,N_4851);
xnor UO_836 (O_836,N_4563,N_4433);
and UO_837 (O_837,N_4506,N_4030);
or UO_838 (O_838,N_4047,N_4119);
xnor UO_839 (O_839,N_4407,N_4980);
xnor UO_840 (O_840,N_4094,N_4607);
nand UO_841 (O_841,N_4386,N_4225);
xor UO_842 (O_842,N_4950,N_4260);
nand UO_843 (O_843,N_4834,N_4261);
xor UO_844 (O_844,N_4857,N_4208);
xnor UO_845 (O_845,N_4073,N_4204);
nand UO_846 (O_846,N_4658,N_4455);
nand UO_847 (O_847,N_4817,N_4466);
nand UO_848 (O_848,N_4218,N_4097);
and UO_849 (O_849,N_4319,N_4511);
xnor UO_850 (O_850,N_4875,N_4299);
xnor UO_851 (O_851,N_4509,N_4944);
nor UO_852 (O_852,N_4264,N_4181);
and UO_853 (O_853,N_4462,N_4640);
xor UO_854 (O_854,N_4619,N_4451);
nand UO_855 (O_855,N_4176,N_4313);
xor UO_856 (O_856,N_4260,N_4028);
nand UO_857 (O_857,N_4393,N_4439);
or UO_858 (O_858,N_4097,N_4852);
nor UO_859 (O_859,N_4794,N_4609);
nand UO_860 (O_860,N_4312,N_4201);
or UO_861 (O_861,N_4906,N_4132);
nor UO_862 (O_862,N_4408,N_4272);
xnor UO_863 (O_863,N_4435,N_4845);
or UO_864 (O_864,N_4988,N_4162);
nor UO_865 (O_865,N_4896,N_4733);
xnor UO_866 (O_866,N_4928,N_4197);
or UO_867 (O_867,N_4882,N_4430);
nand UO_868 (O_868,N_4499,N_4091);
xnor UO_869 (O_869,N_4202,N_4251);
nor UO_870 (O_870,N_4275,N_4063);
and UO_871 (O_871,N_4596,N_4662);
xor UO_872 (O_872,N_4490,N_4705);
or UO_873 (O_873,N_4427,N_4611);
or UO_874 (O_874,N_4256,N_4408);
xor UO_875 (O_875,N_4466,N_4908);
nand UO_876 (O_876,N_4370,N_4924);
nand UO_877 (O_877,N_4381,N_4096);
and UO_878 (O_878,N_4119,N_4648);
xor UO_879 (O_879,N_4367,N_4943);
or UO_880 (O_880,N_4945,N_4505);
nand UO_881 (O_881,N_4251,N_4633);
nand UO_882 (O_882,N_4204,N_4712);
and UO_883 (O_883,N_4407,N_4189);
nand UO_884 (O_884,N_4056,N_4750);
xor UO_885 (O_885,N_4412,N_4416);
xor UO_886 (O_886,N_4465,N_4767);
xnor UO_887 (O_887,N_4437,N_4740);
or UO_888 (O_888,N_4435,N_4220);
nand UO_889 (O_889,N_4893,N_4136);
or UO_890 (O_890,N_4822,N_4665);
nand UO_891 (O_891,N_4304,N_4702);
or UO_892 (O_892,N_4455,N_4847);
nand UO_893 (O_893,N_4958,N_4376);
nand UO_894 (O_894,N_4014,N_4396);
nor UO_895 (O_895,N_4727,N_4715);
and UO_896 (O_896,N_4515,N_4343);
and UO_897 (O_897,N_4281,N_4365);
or UO_898 (O_898,N_4193,N_4637);
and UO_899 (O_899,N_4697,N_4660);
nand UO_900 (O_900,N_4139,N_4006);
nor UO_901 (O_901,N_4976,N_4286);
and UO_902 (O_902,N_4548,N_4272);
nand UO_903 (O_903,N_4911,N_4109);
and UO_904 (O_904,N_4826,N_4882);
xor UO_905 (O_905,N_4028,N_4492);
or UO_906 (O_906,N_4687,N_4675);
nand UO_907 (O_907,N_4031,N_4285);
xor UO_908 (O_908,N_4338,N_4127);
or UO_909 (O_909,N_4079,N_4853);
or UO_910 (O_910,N_4604,N_4569);
nand UO_911 (O_911,N_4631,N_4472);
xor UO_912 (O_912,N_4645,N_4882);
nor UO_913 (O_913,N_4383,N_4428);
xnor UO_914 (O_914,N_4396,N_4756);
nand UO_915 (O_915,N_4731,N_4294);
nor UO_916 (O_916,N_4614,N_4117);
nand UO_917 (O_917,N_4958,N_4146);
xor UO_918 (O_918,N_4082,N_4919);
or UO_919 (O_919,N_4215,N_4413);
nor UO_920 (O_920,N_4596,N_4324);
nand UO_921 (O_921,N_4332,N_4569);
xnor UO_922 (O_922,N_4548,N_4660);
nor UO_923 (O_923,N_4328,N_4712);
and UO_924 (O_924,N_4367,N_4278);
xnor UO_925 (O_925,N_4430,N_4582);
nand UO_926 (O_926,N_4442,N_4793);
nand UO_927 (O_927,N_4196,N_4647);
xnor UO_928 (O_928,N_4498,N_4375);
xor UO_929 (O_929,N_4399,N_4452);
nand UO_930 (O_930,N_4058,N_4978);
and UO_931 (O_931,N_4143,N_4292);
and UO_932 (O_932,N_4133,N_4534);
or UO_933 (O_933,N_4677,N_4553);
and UO_934 (O_934,N_4307,N_4652);
and UO_935 (O_935,N_4465,N_4880);
or UO_936 (O_936,N_4645,N_4972);
xnor UO_937 (O_937,N_4224,N_4109);
and UO_938 (O_938,N_4813,N_4211);
nor UO_939 (O_939,N_4210,N_4222);
xnor UO_940 (O_940,N_4467,N_4744);
and UO_941 (O_941,N_4532,N_4394);
or UO_942 (O_942,N_4714,N_4395);
or UO_943 (O_943,N_4611,N_4326);
or UO_944 (O_944,N_4850,N_4587);
or UO_945 (O_945,N_4911,N_4428);
xor UO_946 (O_946,N_4102,N_4208);
nand UO_947 (O_947,N_4324,N_4106);
or UO_948 (O_948,N_4240,N_4313);
nand UO_949 (O_949,N_4211,N_4283);
nor UO_950 (O_950,N_4379,N_4263);
and UO_951 (O_951,N_4210,N_4028);
xnor UO_952 (O_952,N_4256,N_4442);
or UO_953 (O_953,N_4790,N_4029);
or UO_954 (O_954,N_4782,N_4395);
xnor UO_955 (O_955,N_4367,N_4011);
xnor UO_956 (O_956,N_4467,N_4970);
nand UO_957 (O_957,N_4685,N_4922);
or UO_958 (O_958,N_4098,N_4988);
nand UO_959 (O_959,N_4818,N_4961);
nor UO_960 (O_960,N_4231,N_4138);
and UO_961 (O_961,N_4809,N_4535);
and UO_962 (O_962,N_4612,N_4547);
nor UO_963 (O_963,N_4784,N_4633);
xnor UO_964 (O_964,N_4736,N_4578);
xnor UO_965 (O_965,N_4558,N_4112);
nor UO_966 (O_966,N_4354,N_4999);
nor UO_967 (O_967,N_4496,N_4459);
nor UO_968 (O_968,N_4572,N_4192);
nor UO_969 (O_969,N_4278,N_4088);
nand UO_970 (O_970,N_4193,N_4926);
or UO_971 (O_971,N_4025,N_4982);
or UO_972 (O_972,N_4929,N_4422);
nand UO_973 (O_973,N_4189,N_4477);
or UO_974 (O_974,N_4484,N_4013);
and UO_975 (O_975,N_4178,N_4232);
xor UO_976 (O_976,N_4009,N_4075);
and UO_977 (O_977,N_4651,N_4323);
and UO_978 (O_978,N_4855,N_4491);
nor UO_979 (O_979,N_4017,N_4838);
and UO_980 (O_980,N_4012,N_4577);
and UO_981 (O_981,N_4462,N_4972);
and UO_982 (O_982,N_4396,N_4440);
or UO_983 (O_983,N_4604,N_4995);
or UO_984 (O_984,N_4994,N_4080);
xnor UO_985 (O_985,N_4219,N_4243);
or UO_986 (O_986,N_4698,N_4373);
nand UO_987 (O_987,N_4245,N_4837);
nand UO_988 (O_988,N_4987,N_4675);
nand UO_989 (O_989,N_4662,N_4098);
xnor UO_990 (O_990,N_4249,N_4482);
nor UO_991 (O_991,N_4968,N_4246);
or UO_992 (O_992,N_4987,N_4620);
or UO_993 (O_993,N_4700,N_4794);
nor UO_994 (O_994,N_4154,N_4384);
or UO_995 (O_995,N_4126,N_4163);
and UO_996 (O_996,N_4993,N_4248);
xor UO_997 (O_997,N_4219,N_4217);
nand UO_998 (O_998,N_4126,N_4709);
nor UO_999 (O_999,N_4048,N_4216);
endmodule