module basic_1500_15000_2000_3_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10001,N_10002,N_10003,N_10004,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10016,N_10017,N_10018,N_10019,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10038,N_10040,N_10041,N_10044,N_10045,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10054,N_10055,N_10056,N_10057,N_10059,N_10060,N_10062,N_10063,N_10064,N_10065,N_10067,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10079,N_10081,N_10082,N_10083,N_10084,N_10086,N_10087,N_10088,N_10091,N_10092,N_10093,N_10094,N_10095,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10104,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10117,N_10118,N_10120,N_10121,N_10122,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10184,N_10185,N_10186,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10196,N_10197,N_10198,N_10199,N_10200,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10215,N_10216,N_10217,N_10218,N_10219,N_10221,N_10223,N_10224,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10235,N_10236,N_10237,N_10238,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10249,N_10250,N_10252,N_10255,N_10256,N_10258,N_10259,N_10261,N_10262,N_10264,N_10265,N_10270,N_10272,N_10273,N_10275,N_10277,N_10278,N_10279,N_10281,N_10283,N_10284,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10296,N_10297,N_10299,N_10300,N_10301,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10332,N_10333,N_10337,N_10339,N_10340,N_10341,N_10344,N_10345,N_10347,N_10348,N_10350,N_10351,N_10352,N_10354,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10403,N_10404,N_10405,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10414,N_10415,N_10416,N_10417,N_10419,N_10420,N_10421,N_10424,N_10426,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10445,N_10446,N_10448,N_10449,N_10451,N_10452,N_10454,N_10455,N_10456,N_10457,N_10458,N_10460,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10476,N_10477,N_10479,N_10480,N_10481,N_10482,N_10484,N_10487,N_10488,N_10489,N_10490,N_10492,N_10494,N_10495,N_10496,N_10499,N_10500,N_10503,N_10505,N_10507,N_10508,N_10509,N_10510,N_10511,N_10515,N_10516,N_10517,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10526,N_10528,N_10529,N_10530,N_10531,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10545,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10561,N_10562,N_10563,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10573,N_10574,N_10577,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10594,N_10596,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10606,N_10607,N_10608,N_10609,N_10610,N_10612,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10628,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10659,N_10660,N_10661,N_10662,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10680,N_10681,N_10683,N_10684,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10703,N_10704,N_10705,N_10706,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10728,N_10730,N_10731,N_10733,N_10735,N_10738,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10749,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10771,N_10772,N_10773,N_10775,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10792,N_10793,N_10795,N_10796,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10840,N_10841,N_10842,N_10843,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10860,N_10861,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10882,N_10883,N_10884,N_10886,N_10887,N_10888,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10916,N_10917,N_10918,N_10920,N_10921,N_10923,N_10924,N_10925,N_10926,N_10929,N_10930,N_10931,N_10932,N_10933,N_10936,N_10938,N_10939,N_10941,N_10943,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10964,N_10965,N_10968,N_10969,N_10971,N_10972,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10981,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11009,N_11011,N_11012,N_11013,N_11015,N_11016,N_11017,N_11018,N_11019,N_11021,N_11022,N_11024,N_11025,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11045,N_11046,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11079,N_11081,N_11082,N_11083,N_11084,N_11086,N_11087,N_11088,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11130,N_11131,N_11132,N_11134,N_11135,N_11136,N_11137,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11158,N_11159,N_11160,N_11162,N_11164,N_11166,N_11167,N_11168,N_11171,N_11172,N_11174,N_11175,N_11178,N_11179,N_11180,N_11181,N_11183,N_11186,N_11187,N_11188,N_11189,N_11191,N_11192,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11202,N_11203,N_11204,N_11205,N_11207,N_11208,N_11209,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11241,N_11242,N_11243,N_11244,N_11247,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11259,N_11260,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11292,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11310,N_11311,N_11312,N_11313,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11324,N_11325,N_11326,N_11327,N_11328,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11338,N_11339,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11353,N_11354,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11375,N_11377,N_11381,N_11383,N_11384,N_11385,N_11387,N_11388,N_11389,N_11390,N_11391,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11401,N_11402,N_11403,N_11404,N_11405,N_11407,N_11409,N_11410,N_11411,N_11412,N_11414,N_11415,N_11416,N_11417,N_11419,N_11420,N_11421,N_11422,N_11424,N_11425,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11438,N_11439,N_11440,N_11441,N_11445,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11466,N_11468,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11482,N_11483,N_11484,N_11486,N_11487,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11522,N_11523,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11544,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11556,N_11557,N_11558,N_11559,N_11561,N_11562,N_11564,N_11565,N_11566,N_11568,N_11570,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11592,N_11594,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11616,N_11617,N_11618,N_11619,N_11621,N_11622,N_11624,N_11625,N_11626,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11676,N_11677,N_11678,N_11679,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11714,N_11715,N_11716,N_11717,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11758,N_11759,N_11760,N_11761,N_11766,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11778,N_11780,N_11781,N_11782,N_11783,N_11785,N_11788,N_11790,N_11791,N_11792,N_11793,N_11794,N_11796,N_11797,N_11798,N_11799,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11811,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11842,N_11843,N_11844,N_11845,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11858,N_11859,N_11860,N_11861,N_11863,N_11864,N_11865,N_11866,N_11867,N_11869,N_11870,N_11872,N_11873,N_11874,N_11875,N_11879,N_11880,N_11881,N_11883,N_11885,N_11886,N_11887,N_11888,N_11890,N_11891,N_11893,N_11894,N_11895,N_11896,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11905,N_11907,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11916,N_11917,N_11919,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11941,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11954,N_11955,N_11956,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11967,N_11968,N_11969,N_11970,N_11971,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11980,N_11981,N_11982,N_11984,N_11985,N_11986,N_11987,N_11989,N_11990,N_11991,N_11992,N_11994,N_11995,N_11996,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12013,N_12015,N_12016,N_12017,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12035,N_12036,N_12037,N_12039,N_12041,N_12042,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12083,N_12084,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12101,N_12102,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12131,N_12132,N_12133,N_12134,N_12136,N_12137,N_12138,N_12139,N_12141,N_12142,N_12143,N_12144,N_12146,N_12147,N_12149,N_12150,N_12151,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12161,N_12162,N_12164,N_12166,N_12167,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12178,N_12179,N_12180,N_12181,N_12182,N_12184,N_12185,N_12186,N_12188,N_12191,N_12192,N_12193,N_12194,N_12195,N_12197,N_12198,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12208,N_12209,N_12211,N_12212,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12236,N_12237,N_12238,N_12239,N_12240,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12254,N_12255,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12288,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12305,N_12307,N_12308,N_12309,N_12310,N_12311,N_12314,N_12316,N_12318,N_12320,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12333,N_12334,N_12335,N_12336,N_12337,N_12339,N_12341,N_12342,N_12343,N_12345,N_12348,N_12349,N_12351,N_12352,N_12353,N_12355,N_12356,N_12357,N_12358,N_12359,N_12361,N_12362,N_12365,N_12366,N_12367,N_12369,N_12370,N_12371,N_12373,N_12374,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12386,N_12387,N_12389,N_12390,N_12392,N_12393,N_12394,N_12395,N_12399,N_12400,N_12402,N_12403,N_12404,N_12405,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12428,N_12429,N_12430,N_12431,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12444,N_12445,N_12449,N_12450,N_12452,N_12453,N_12454,N_12457,N_12458,N_12459,N_12460,N_12461,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12481,N_12482,N_12483,N_12484,N_12486,N_12487,N_12488,N_12489,N_12490,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12513,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12546,N_12547,N_12548,N_12549,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12562,N_12563,N_12564,N_12565,N_12568,N_12569,N_12571,N_12572,N_12573,N_12574,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12583,N_12584,N_12585,N_12586,N_12587,N_12589,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12609,N_12610,N_12611,N_12612,N_12613,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12638,N_12639,N_12640,N_12641,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12664,N_12665,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12684,N_12686,N_12687,N_12688,N_12689,N_12690,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12700,N_12701,N_12702,N_12703,N_12705,N_12706,N_12708,N_12709,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12737,N_12738,N_12739,N_12741,N_12742,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12764,N_12765,N_12767,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12782,N_12783,N_12784,N_12785,N_12786,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12804,N_12805,N_12806,N_12807,N_12808,N_12810,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12823,N_12825,N_12826,N_12827,N_12828,N_12829,N_12831,N_12832,N_12834,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12847,N_12848,N_12849,N_12850,N_12852,N_12853,N_12855,N_12856,N_12857,N_12858,N_12860,N_12862,N_12863,N_12864,N_12867,N_12869,N_12872,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12882,N_12883,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12909,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12920,N_12921,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12971,N_12973,N_12974,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12983,N_12984,N_12987,N_12988,N_12991,N_12992,N_12993,N_12994,N_12996,N_12997,N_12999,N_13001,N_13002,N_13003,N_13005,N_13007,N_13008,N_13009,N_13010,N_13011,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13022,N_13023,N_13024,N_13025,N_13026,N_13029,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13041,N_13042,N_13044,N_13046,N_13047,N_13048,N_13049,N_13050,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13061,N_13062,N_13063,N_13064,N_13068,N_13069,N_13070,N_13071,N_13073,N_13074,N_13075,N_13077,N_13079,N_13080,N_13081,N_13082,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13107,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13118,N_13119,N_13120,N_13121,N_13122,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13134,N_13135,N_13136,N_13138,N_13139,N_13140,N_13141,N_13143,N_13144,N_13145,N_13147,N_13148,N_13149,N_13150,N_13152,N_13153,N_13155,N_13156,N_13158,N_13159,N_13160,N_13161,N_13164,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13187,N_13190,N_13191,N_13192,N_13195,N_13197,N_13199,N_13200,N_13202,N_13203,N_13204,N_13205,N_13208,N_13209,N_13210,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13229,N_13230,N_13231,N_13232,N_13233,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13265,N_13266,N_13267,N_13268,N_13269,N_13271,N_13273,N_13274,N_13275,N_13278,N_13279,N_13280,N_13282,N_13283,N_13284,N_13285,N_13286,N_13288,N_13289,N_13290,N_13292,N_13294,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13307,N_13308,N_13309,N_13311,N_13312,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13323,N_13324,N_13325,N_13326,N_13328,N_13329,N_13330,N_13331,N_13332,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13360,N_13361,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13375,N_13376,N_13378,N_13379,N_13381,N_13382,N_13383,N_13385,N_13386,N_13387,N_13388,N_13389,N_13392,N_13393,N_13394,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13431,N_13432,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13467,N_13468,N_13469,N_13473,N_13474,N_13475,N_13476,N_13478,N_13479,N_13480,N_13482,N_13483,N_13484,N_13485,N_13487,N_13488,N_13489,N_13490,N_13493,N_13494,N_13495,N_13496,N_13499,N_13501,N_13503,N_13504,N_13506,N_13507,N_13508,N_13509,N_13510,N_13512,N_13513,N_13516,N_13517,N_13518,N_13519,N_13520,N_13523,N_13524,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13548,N_13549,N_13550,N_13551,N_13552,N_13554,N_13555,N_13557,N_13559,N_13560,N_13562,N_13563,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13573,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13604,N_13605,N_13606,N_13607,N_13608,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13620,N_13621,N_13624,N_13625,N_13626,N_13627,N_13628,N_13630,N_13631,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13648,N_13649,N_13650,N_13651,N_13652,N_13657,N_13659,N_13661,N_13662,N_13663,N_13664,N_13666,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13678,N_13679,N_13680,N_13681,N_13682,N_13684,N_13686,N_13687,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13696,N_13697,N_13698,N_13699,N_13700,N_13703,N_13704,N_13705,N_13706,N_13708,N_13709,N_13710,N_13711,N_13713,N_13715,N_13716,N_13717,N_13718,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13735,N_13736,N_13738,N_13739,N_13741,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13754,N_13755,N_13756,N_13759,N_13761,N_13762,N_13763,N_13765,N_13766,N_13767,N_13769,N_13771,N_13772,N_13773,N_13775,N_13776,N_13777,N_13778,N_13780,N_13781,N_13782,N_13783,N_13784,N_13786,N_13787,N_13788,N_13789,N_13791,N_13792,N_13794,N_13795,N_13796,N_13797,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13812,N_13813,N_13815,N_13816,N_13817,N_13819,N_13820,N_13821,N_13822,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13835,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13863,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13872,N_13873,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13885,N_13886,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13897,N_13898,N_13901,N_13902,N_13905,N_13906,N_13907,N_13908,N_13909,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13925,N_13926,N_13927,N_13929,N_13930,N_13931,N_13933,N_13935,N_13936,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13952,N_13953,N_13955,N_13956,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13965,N_13966,N_13967,N_13968,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14017,N_14019,N_14020,N_14022,N_14023,N_14024,N_14025,N_14029,N_14031,N_14033,N_14034,N_14036,N_14038,N_14039,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14051,N_14052,N_14053,N_14054,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14066,N_14068,N_14069,N_14070,N_14071,N_14072,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14084,N_14085,N_14086,N_14089,N_14090,N_14091,N_14092,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14109,N_14110,N_14111,N_14112,N_14113,N_14115,N_14116,N_14117,N_14119,N_14120,N_14121,N_14122,N_14124,N_14125,N_14126,N_14127,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14143,N_14144,N_14145,N_14146,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14169,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14178,N_14179,N_14181,N_14182,N_14184,N_14185,N_14186,N_14187,N_14188,N_14190,N_14192,N_14193,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14211,N_14212,N_14213,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14246,N_14247,N_14248,N_14249,N_14250,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14262,N_14264,N_14266,N_14267,N_14268,N_14270,N_14271,N_14272,N_14273,N_14275,N_14276,N_14277,N_14278,N_14279,N_14281,N_14282,N_14283,N_14284,N_14285,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14326,N_14328,N_14330,N_14331,N_14332,N_14334,N_14336,N_14338,N_14339,N_14340,N_14342,N_14346,N_14347,N_14348,N_14349,N_14351,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14362,N_14363,N_14364,N_14365,N_14366,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14377,N_14378,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14399,N_14400,N_14401,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14423,N_14424,N_14425,N_14426,N_14430,N_14431,N_14432,N_14433,N_14434,N_14436,N_14438,N_14439,N_14440,N_14441,N_14443,N_14444,N_14445,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14492,N_14493,N_14494,N_14495,N_14497,N_14499,N_14500,N_14503,N_14504,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14538,N_14539,N_14540,N_14542,N_14545,N_14546,N_14547,N_14548,N_14550,N_14551,N_14552,N_14553,N_14555,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14577,N_14578,N_14579,N_14580,N_14581,N_14583,N_14584,N_14589,N_14590,N_14591,N_14592,N_14595,N_14596,N_14599,N_14601,N_14602,N_14603,N_14605,N_14606,N_14607,N_14608,N_14609,N_14612,N_14613,N_14614,N_14615,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14636,N_14640,N_14641,N_14643,N_14644,N_14645,N_14646,N_14647,N_14649,N_14650,N_14654,N_14655,N_14656,N_14658,N_14660,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14670,N_14672,N_14673,N_14674,N_14675,N_14676,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14689,N_14690,N_14691,N_14692,N_14694,N_14695,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14709,N_14711,N_14712,N_14713,N_14714,N_14715,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14731,N_14732,N_14733,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14743,N_14744,N_14745,N_14746,N_14748,N_14749,N_14750,N_14752,N_14754,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14764,N_14765,N_14767,N_14768,N_14769,N_14770,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14780,N_14781,N_14782,N_14783,N_14785,N_14786,N_14787,N_14789,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14805,N_14806,N_14808,N_14810,N_14813,N_14817,N_14818,N_14819,N_14821,N_14822,N_14824,N_14825,N_14826,N_14827,N_14830,N_14831,N_14832,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14844,N_14846,N_14847,N_14851,N_14852,N_14853,N_14854,N_14855,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14874,N_14876,N_14877,N_14879,N_14880,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14911,N_14912,N_14913,N_14914,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14928,N_14929,N_14930,N_14932,N_14934,N_14935,N_14936,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14954,N_14955,N_14956,N_14957,N_14959,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14972,N_14973,N_14974,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14986,N_14987,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_222,In_400);
nand U1 (N_1,In_174,In_424);
or U2 (N_2,In_270,In_1034);
xnor U3 (N_3,In_601,In_1070);
nand U4 (N_4,In_187,In_412);
or U5 (N_5,In_1350,In_846);
or U6 (N_6,In_479,In_120);
xnor U7 (N_7,In_1454,In_926);
nor U8 (N_8,In_1038,In_1299);
or U9 (N_9,In_1440,In_506);
or U10 (N_10,In_943,In_93);
nor U11 (N_11,In_1474,In_1475);
and U12 (N_12,In_1412,In_733);
or U13 (N_13,In_746,In_1426);
nor U14 (N_14,In_1497,In_491);
xnor U15 (N_15,In_1394,In_442);
or U16 (N_16,In_96,In_142);
xor U17 (N_17,In_1053,In_299);
nor U18 (N_18,In_903,In_518);
xnor U19 (N_19,In_1376,In_1175);
xor U20 (N_20,In_257,In_841);
or U21 (N_21,In_282,In_769);
nand U22 (N_22,In_27,In_304);
nor U23 (N_23,In_526,In_1035);
nand U24 (N_24,In_835,In_1476);
xnor U25 (N_25,In_188,In_156);
nand U26 (N_26,In_105,In_229);
or U27 (N_27,In_962,In_267);
nand U28 (N_28,In_625,In_923);
nor U29 (N_29,In_1495,In_1110);
nand U30 (N_30,In_492,In_496);
nor U31 (N_31,In_1095,In_1319);
nor U32 (N_32,In_1007,In_931);
nand U33 (N_33,In_171,In_1107);
nor U34 (N_34,In_1121,In_1159);
and U35 (N_35,In_677,In_644);
nand U36 (N_36,In_1245,In_1073);
nand U37 (N_37,In_1260,In_87);
or U38 (N_38,In_398,In_629);
nor U39 (N_39,In_432,In_390);
nor U40 (N_40,In_1209,In_408);
and U41 (N_41,In_568,In_210);
xnor U42 (N_42,In_1400,In_366);
and U43 (N_43,In_322,In_704);
nand U44 (N_44,In_1261,In_839);
nor U45 (N_45,In_633,In_1193);
nand U46 (N_46,In_612,In_1407);
or U47 (N_47,In_60,In_944);
or U48 (N_48,In_183,In_384);
and U49 (N_49,In_1360,In_805);
or U50 (N_50,In_972,In_732);
nand U51 (N_51,In_1258,In_1353);
and U52 (N_52,In_72,In_696);
and U53 (N_53,In_1304,In_974);
and U54 (N_54,In_1392,In_28);
nor U55 (N_55,In_129,In_859);
or U56 (N_56,In_177,In_193);
or U57 (N_57,In_1137,In_1220);
nor U58 (N_58,In_75,In_1082);
nand U59 (N_59,In_471,In_488);
xnor U60 (N_60,In_434,In_1344);
xor U61 (N_61,In_61,In_1165);
or U62 (N_62,In_1181,In_619);
nand U63 (N_63,In_416,In_305);
nor U64 (N_64,In_636,In_428);
or U65 (N_65,In_138,In_1133);
and U66 (N_66,In_1281,In_1373);
xor U67 (N_67,In_1347,In_350);
or U68 (N_68,In_191,In_295);
and U69 (N_69,In_49,In_701);
or U70 (N_70,In_1183,In_111);
nor U71 (N_71,In_1225,In_1036);
nor U72 (N_72,In_346,In_64);
or U73 (N_73,In_809,In_969);
xnor U74 (N_74,In_1105,In_914);
and U75 (N_75,In_976,In_220);
and U76 (N_76,In_1386,In_531);
nor U77 (N_77,In_600,In_461);
and U78 (N_78,In_648,In_760);
nor U79 (N_79,In_1291,In_803);
xnor U80 (N_80,In_1419,In_453);
xnor U81 (N_81,In_1187,In_388);
and U82 (N_82,In_1072,In_891);
and U83 (N_83,In_6,In_235);
and U84 (N_84,In_1442,In_659);
nor U85 (N_85,In_166,In_475);
nand U86 (N_86,In_317,In_233);
and U87 (N_87,In_54,In_377);
nor U88 (N_88,In_345,In_418);
or U89 (N_89,In_1453,In_1152);
and U90 (N_90,In_785,In_389);
nor U91 (N_91,In_1354,In_1459);
nor U92 (N_92,In_1264,In_1008);
nand U93 (N_93,In_1092,In_318);
xnor U94 (N_94,In_213,In_737);
nand U95 (N_95,In_1224,In_36);
and U96 (N_96,In_1162,In_770);
nand U97 (N_97,In_1172,In_1303);
nor U98 (N_98,In_1102,In_620);
or U99 (N_99,In_922,In_279);
xor U100 (N_100,In_975,In_478);
xnor U101 (N_101,In_1109,In_1000);
or U102 (N_102,In_731,In_1012);
xnor U103 (N_103,In_1408,In_796);
and U104 (N_104,In_827,In_735);
nor U105 (N_105,In_106,In_1307);
nor U106 (N_106,In_519,In_118);
xor U107 (N_107,In_186,In_31);
and U108 (N_108,In_965,In_830);
xor U109 (N_109,In_550,In_1276);
or U110 (N_110,In_817,In_1483);
xnor U111 (N_111,In_481,In_507);
and U112 (N_112,In_705,In_140);
or U113 (N_113,In_1460,In_1315);
xnor U114 (N_114,In_407,In_379);
or U115 (N_115,In_1246,In_865);
xor U116 (N_116,In_843,In_949);
and U117 (N_117,In_1485,In_530);
or U118 (N_118,In_825,In_929);
nand U119 (N_119,In_406,In_1016);
or U120 (N_120,In_1463,In_589);
nand U121 (N_121,In_800,In_444);
xor U122 (N_122,In_1179,In_1215);
or U123 (N_123,In_273,In_940);
xor U124 (N_124,In_595,In_62);
xor U125 (N_125,In_1122,In_1287);
and U126 (N_126,In_1279,In_660);
nor U127 (N_127,In_413,In_1479);
xnor U128 (N_128,In_980,In_41);
xnor U129 (N_129,In_1283,In_1021);
and U130 (N_130,In_992,In_1249);
and U131 (N_131,In_1481,In_924);
or U132 (N_132,In_1135,In_288);
nand U133 (N_133,In_730,In_276);
xnor U134 (N_134,In_338,In_1241);
nor U135 (N_135,In_269,In_1156);
xnor U136 (N_136,In_1418,In_837);
nand U137 (N_137,In_1484,In_694);
or U138 (N_138,In_672,In_290);
nand U139 (N_139,In_1368,In_647);
nand U140 (N_140,In_561,In_1268);
nand U141 (N_141,In_393,In_352);
and U142 (N_142,In_375,In_1234);
nand U143 (N_143,In_543,In_570);
nand U144 (N_144,In_856,In_109);
and U145 (N_145,In_981,In_246);
and U146 (N_146,In_313,In_307);
or U147 (N_147,In_954,In_30);
nor U148 (N_148,In_1409,In_1056);
and U149 (N_149,In_199,In_1118);
nand U150 (N_150,In_15,In_314);
and U151 (N_151,In_627,In_897);
or U152 (N_152,In_948,In_172);
and U153 (N_153,In_368,In_414);
and U154 (N_154,In_429,In_242);
xor U155 (N_155,In_592,In_831);
and U156 (N_156,In_1158,In_1085);
and U157 (N_157,In_968,In_882);
and U158 (N_158,In_904,In_1112);
or U159 (N_159,In_1089,In_632);
or U160 (N_160,In_484,In_997);
and U161 (N_161,In_739,In_1232);
xor U162 (N_162,In_925,In_33);
or U163 (N_163,In_17,In_994);
xor U164 (N_164,In_1065,In_333);
nor U165 (N_165,In_1169,In_1014);
and U166 (N_166,In_819,In_510);
nor U167 (N_167,In_117,In_744);
or U168 (N_168,In_115,In_983);
and U169 (N_169,In_999,In_802);
nand U170 (N_170,In_901,In_48);
nor U171 (N_171,In_624,In_1123);
nor U172 (N_172,In_749,In_359);
or U173 (N_173,In_579,In_670);
nor U174 (N_174,In_702,In_1028);
nor U175 (N_175,In_1151,In_437);
xnor U176 (N_176,In_291,In_970);
nand U177 (N_177,In_467,In_417);
xor U178 (N_178,In_371,In_150);
or U179 (N_179,In_854,In_1136);
or U180 (N_180,In_480,In_750);
nand U181 (N_181,In_263,In_516);
and U182 (N_182,In_1163,In_144);
xor U183 (N_183,In_939,In_1450);
and U184 (N_184,In_1239,In_391);
xnor U185 (N_185,In_798,In_1348);
nor U186 (N_186,In_905,In_214);
or U187 (N_187,In_205,In_661);
nand U188 (N_188,In_1037,In_883);
and U189 (N_189,In_973,In_907);
nand U190 (N_190,In_208,In_1295);
and U191 (N_191,In_761,In_112);
nor U192 (N_192,In_1214,In_961);
and U193 (N_193,In_1486,In_327);
nor U194 (N_194,In_896,In_887);
xnor U195 (N_195,In_296,In_792);
or U196 (N_196,In_861,In_362);
nor U197 (N_197,In_50,In_137);
and U198 (N_198,In_1157,In_1425);
xnor U199 (N_199,In_43,In_1010);
xor U200 (N_200,In_94,In_122);
nand U201 (N_201,In_126,In_281);
xor U202 (N_202,In_1115,In_185);
or U203 (N_203,In_868,In_173);
xor U204 (N_204,In_203,In_522);
nor U205 (N_205,In_811,In_202);
and U206 (N_206,In_682,In_131);
nor U207 (N_207,In_878,In_86);
xor U208 (N_208,In_228,In_1243);
nand U209 (N_209,In_1043,In_476);
xnor U210 (N_210,In_495,In_740);
xnor U211 (N_211,In_1445,In_283);
and U212 (N_212,In_993,In_168);
nor U213 (N_213,In_1168,In_351);
and U214 (N_214,In_574,In_247);
nor U215 (N_215,In_1274,In_1084);
nand U216 (N_216,In_1222,In_571);
xor U217 (N_217,In_306,In_19);
nand U218 (N_218,In_1026,In_1447);
nor U219 (N_219,In_1393,In_829);
and U220 (N_220,In_1269,In_1013);
and U221 (N_221,In_603,In_13);
nand U222 (N_222,In_845,In_666);
or U223 (N_223,In_842,In_53);
or U224 (N_224,In_312,In_330);
or U225 (N_225,In_628,In_280);
nand U226 (N_226,In_1430,In_919);
xor U227 (N_227,In_630,In_1480);
xor U228 (N_228,In_611,In_1321);
or U229 (N_229,In_626,In_42);
xnor U230 (N_230,In_1042,In_609);
xor U231 (N_231,In_723,In_1332);
and U232 (N_232,In_405,In_675);
nand U233 (N_233,In_423,In_1455);
nand U234 (N_234,In_245,In_365);
or U235 (N_235,In_1100,In_409);
nand U236 (N_236,In_98,In_427);
nor U237 (N_237,In_466,In_308);
nand U238 (N_238,In_286,In_1417);
and U239 (N_239,In_727,In_271);
or U240 (N_240,In_380,In_1211);
nand U241 (N_241,In_0,In_930);
nand U242 (N_242,In_1490,In_547);
xor U243 (N_243,In_1044,In_1491);
xor U244 (N_244,In_1174,In_420);
xnor U245 (N_245,In_680,In_1231);
and U246 (N_246,In_794,In_1171);
nor U247 (N_247,In_544,In_256);
and U248 (N_248,In_219,In_1247);
nand U249 (N_249,In_78,In_458);
nand U250 (N_250,In_797,In_344);
nor U251 (N_251,In_1032,In_1147);
xor U252 (N_252,In_1326,In_606);
nor U253 (N_253,In_1004,In_321);
nor U254 (N_254,In_332,In_277);
or U255 (N_255,In_248,In_1015);
nor U256 (N_256,In_482,In_646);
xnor U257 (N_257,In_751,In_1433);
or U258 (N_258,In_1219,In_1421);
nand U259 (N_259,In_1254,In_1296);
nand U260 (N_260,In_1054,In_575);
nor U261 (N_261,In_806,In_422);
nor U262 (N_262,In_664,In_1025);
and U263 (N_263,In_1297,In_446);
or U264 (N_264,In_1443,In_381);
or U265 (N_265,In_1049,In_58);
or U266 (N_266,In_1461,In_1127);
and U267 (N_267,In_1478,In_642);
xnor U268 (N_268,In_272,In_1359);
xnor U269 (N_269,In_537,In_1005);
or U270 (N_270,In_951,In_486);
nand U271 (N_271,In_40,In_1235);
or U272 (N_272,In_370,In_1040);
or U273 (N_273,In_1079,In_70);
xnor U274 (N_274,In_523,In_671);
and U275 (N_275,In_20,In_847);
nor U276 (N_276,In_711,In_353);
nand U277 (N_277,In_278,In_726);
and U278 (N_278,In_1464,In_713);
and U279 (N_279,In_781,In_734);
nand U280 (N_280,In_1385,In_443);
xnor U281 (N_281,In_436,In_967);
nand U282 (N_282,In_977,In_237);
xnor U283 (N_283,In_1126,In_425);
nand U284 (N_284,In_1275,In_114);
xor U285 (N_285,In_1208,In_617);
nand U286 (N_286,In_251,In_56);
or U287 (N_287,In_1190,In_989);
and U288 (N_288,In_789,In_767);
xor U289 (N_289,In_867,In_364);
xor U290 (N_290,In_16,In_1302);
nand U291 (N_291,In_116,In_473);
and U292 (N_292,In_752,In_127);
nor U293 (N_293,In_1128,In_1221);
nand U294 (N_294,In_1017,In_936);
and U295 (N_295,In_1227,In_293);
or U296 (N_296,In_971,In_988);
nand U297 (N_297,In_801,In_259);
nand U298 (N_298,In_884,In_950);
or U299 (N_299,In_435,In_196);
and U300 (N_300,In_1194,In_655);
or U301 (N_301,In_71,In_1041);
nor U302 (N_302,In_1131,In_906);
or U303 (N_303,In_1201,In_1370);
nor U304 (N_304,In_1191,In_598);
or U305 (N_305,In_464,In_615);
or U306 (N_306,In_768,In_665);
nor U307 (N_307,In_1244,In_310);
nor U308 (N_308,In_978,In_149);
xnor U309 (N_309,In_1378,In_37);
and U310 (N_310,In_838,In_650);
and U311 (N_311,In_132,In_152);
nor U312 (N_312,In_240,In_928);
nor U313 (N_313,In_1331,In_1120);
nor U314 (N_314,In_754,In_1024);
xnor U315 (N_315,In_74,In_1031);
nor U316 (N_316,In_1472,In_175);
xor U317 (N_317,In_758,In_101);
nor U318 (N_318,In_591,In_549);
xor U319 (N_319,In_532,In_1064);
nor U320 (N_320,In_542,In_700);
and U321 (N_321,In_1259,In_169);
or U322 (N_322,In_946,In_1387);
and U323 (N_323,In_404,In_1143);
xnor U324 (N_324,In_160,In_294);
and U325 (N_325,In_1027,In_95);
and U326 (N_326,In_1200,In_123);
nor U327 (N_327,In_1205,In_662);
nor U328 (N_328,In_657,In_490);
xnor U329 (N_329,In_764,In_315);
and U330 (N_330,In_1351,In_1406);
and U331 (N_331,In_703,In_691);
nand U332 (N_332,In_1184,In_864);
xnor U333 (N_333,In_1057,In_1199);
xor U334 (N_334,In_439,In_772);
and U335 (N_335,In_1177,In_4);
and U336 (N_336,In_415,In_1144);
and U337 (N_337,In_1423,In_584);
xnor U338 (N_338,In_1164,In_987);
or U339 (N_339,In_1062,In_546);
or U340 (N_340,In_722,In_690);
nand U341 (N_341,In_715,In_128);
nand U342 (N_342,In_335,In_525);
and U343 (N_343,In_1397,In_1306);
nor U344 (N_344,In_1388,In_1271);
nor U345 (N_345,In_728,In_824);
nand U346 (N_346,In_374,In_863);
nand U347 (N_347,In_658,In_1342);
or U348 (N_348,In_258,In_300);
or U349 (N_349,In_500,In_206);
nand U350 (N_350,In_182,In_1093);
or U351 (N_351,In_511,In_729);
or U352 (N_352,In_1142,In_1337);
xor U353 (N_353,In_1067,In_1290);
nor U354 (N_354,In_515,In_55);
xor U355 (N_355,In_339,In_419);
nor U356 (N_356,In_462,In_382);
nand U357 (N_357,In_483,In_1277);
and U358 (N_358,In_1237,In_355);
or U359 (N_359,In_1236,In_261);
nor U360 (N_360,In_1132,In_285);
xor U361 (N_361,In_504,In_757);
nor U362 (N_362,In_618,In_1233);
and U363 (N_363,In_1019,In_956);
and U364 (N_364,In_885,In_309);
and U365 (N_365,In_320,In_807);
nor U366 (N_366,In_871,In_472);
and U367 (N_367,In_763,In_814);
or U368 (N_368,In_201,In_44);
and U369 (N_369,In_836,In_1381);
xor U370 (N_370,In_164,In_1195);
and U371 (N_371,In_1002,In_230);
nand U372 (N_372,In_91,In_1161);
nor U373 (N_373,In_1153,In_1316);
nand U374 (N_374,In_1011,In_902);
nand U375 (N_375,In_681,In_585);
and U376 (N_376,In_1372,In_254);
or U377 (N_377,In_890,In_387);
xor U378 (N_378,In_262,In_759);
nor U379 (N_379,In_813,In_1140);
and U380 (N_380,In_1061,In_832);
xnor U381 (N_381,In_941,In_1116);
or U382 (N_382,In_1050,In_996);
nor U383 (N_383,In_431,In_583);
xor U384 (N_384,In_82,In_474);
nand U385 (N_385,In_323,In_343);
or U386 (N_386,In_146,In_621);
xnor U387 (N_387,In_912,In_1009);
and U388 (N_388,In_1023,In_1148);
nor U389 (N_389,In_687,In_298);
or U390 (N_390,In_100,In_1402);
and U391 (N_391,In_909,In_1470);
nand U392 (N_392,In_1248,In_102);
xnor U393 (N_393,In_1203,In_1436);
and U394 (N_394,In_1001,In_1059);
or U395 (N_395,In_512,In_1060);
and U396 (N_396,In_1288,In_910);
and U397 (N_397,In_157,In_198);
xnor U398 (N_398,In_1074,In_778);
xnor U399 (N_399,In_745,In_1322);
nand U400 (N_400,In_217,In_1047);
nor U401 (N_401,In_623,In_348);
nand U402 (N_402,In_945,In_594);
nand U403 (N_403,In_556,In_1086);
nand U404 (N_404,In_1366,In_1451);
nand U405 (N_405,In_640,In_99);
and U406 (N_406,In_421,In_1180);
nor U407 (N_407,In_238,In_51);
nor U408 (N_408,In_777,In_107);
nor U409 (N_409,In_1379,In_849);
nor U410 (N_410,In_1160,In_287);
or U411 (N_411,In_678,In_334);
xnor U412 (N_412,In_1380,In_869);
and U413 (N_413,In_1091,In_1336);
xnor U414 (N_414,In_855,In_979);
nor U415 (N_415,In_1437,In_14);
and U416 (N_416,In_1401,In_3);
and U417 (N_417,In_1146,In_1081);
and U418 (N_418,In_493,In_139);
xnor U419 (N_419,In_1098,In_65);
xor U420 (N_420,In_587,In_1045);
nor U421 (N_421,In_643,In_73);
nor U422 (N_422,In_1301,In_656);
nand U423 (N_423,In_1155,In_524);
xnor U424 (N_424,In_337,In_1108);
or U425 (N_425,In_888,In_674);
nand U426 (N_426,In_148,In_1489);
xor U427 (N_427,In_477,In_81);
xor U428 (N_428,In_953,In_514);
nor U429 (N_429,In_1345,In_1446);
nor U430 (N_430,In_1206,In_1106);
xnor U431 (N_431,In_508,In_1312);
and U432 (N_432,In_818,In_376);
nand U433 (N_433,In_358,In_685);
xnor U434 (N_434,In_1189,In_249);
and U435 (N_435,In_121,In_1469);
nand U436 (N_436,In_1328,In_103);
nor U437 (N_437,In_1363,In_1075);
nand U438 (N_438,In_1333,In_1265);
and U439 (N_439,In_639,In_1251);
and U440 (N_440,In_1444,In_899);
and U441 (N_441,In_637,In_141);
xor U442 (N_442,In_79,In_717);
nor U443 (N_443,In_39,In_373);
and U444 (N_444,In_812,In_59);
and U445 (N_445,In_1051,In_34);
nor U446 (N_446,In_569,In_255);
or U447 (N_447,In_253,In_113);
xnor U448 (N_448,In_718,In_534);
nor U449 (N_449,In_565,In_178);
or U450 (N_450,In_808,In_1327);
xnor U451 (N_451,In_21,In_212);
and U452 (N_452,In_1192,In_553);
or U453 (N_453,In_1167,In_485);
nand U454 (N_454,In_1,In_1055);
or U455 (N_455,In_452,In_505);
nand U456 (N_456,In_342,In_225);
xor U457 (N_457,In_135,In_908);
and U458 (N_458,In_635,In_1358);
nand U459 (N_459,In_1252,In_1267);
xor U460 (N_460,In_959,In_83);
nand U461 (N_461,In_935,In_1101);
nand U462 (N_462,In_1488,In_1431);
nand U463 (N_463,In_533,In_1130);
nand U464 (N_464,In_154,In_1256);
xor U465 (N_465,In_52,In_881);
nor U466 (N_466,In_143,In_1238);
xor U467 (N_467,In_145,In_274);
nand U468 (N_468,In_1077,In_302);
xor U469 (N_469,In_89,In_12);
and U470 (N_470,In_1405,In_554);
nor U471 (N_471,In_634,In_1399);
or U472 (N_472,In_155,In_38);
nor U473 (N_473,In_1066,In_762);
nand U474 (N_474,In_189,In_698);
and U475 (N_475,In_470,In_775);
nor U476 (N_476,In_557,In_572);
xnor U477 (N_477,In_581,In_821);
and U478 (N_478,In_1294,In_963);
nand U479 (N_479,In_450,In_984);
or U480 (N_480,In_264,In_638);
nand U481 (N_481,In_877,In_1340);
nor U482 (N_482,In_870,In_576);
or U483 (N_483,In_297,In_456);
or U484 (N_484,In_67,In_879);
xnor U485 (N_485,In_652,In_403);
and U486 (N_486,In_354,In_231);
or U487 (N_487,In_826,In_325);
or U488 (N_488,In_1398,In_218);
or U489 (N_489,In_1438,In_957);
or U490 (N_490,In_784,In_834);
nor U491 (N_491,In_289,In_560);
nand U492 (N_492,In_426,In_517);
or U493 (N_493,In_853,In_1103);
nor U494 (N_494,In_689,In_934);
xor U495 (N_495,In_190,In_918);
xnor U496 (N_496,In_1414,In_23);
or U497 (N_497,In_577,In_1210);
nand U498 (N_498,In_361,In_663);
nor U499 (N_499,In_1117,In_130);
nor U500 (N_500,In_669,In_159);
or U501 (N_501,In_607,In_236);
nor U502 (N_502,In_326,In_783);
or U503 (N_503,In_593,In_782);
xor U504 (N_504,In_378,In_1145);
nor U505 (N_505,In_736,In_136);
xor U506 (N_506,In_340,In_455);
nand U507 (N_507,In_933,In_699);
xor U508 (N_508,In_367,In_932);
and U509 (N_509,In_68,In_184);
xnor U510 (N_510,In_1069,In_1305);
xor U511 (N_511,In_1223,In_1341);
or U512 (N_512,In_873,In_163);
and U513 (N_513,In_747,In_688);
xor U514 (N_514,In_104,In_1330);
xor U515 (N_515,In_937,In_108);
nand U516 (N_516,In_920,In_349);
and U517 (N_517,In_395,In_766);
and U518 (N_518,In_958,In_324);
nand U519 (N_519,In_24,In_386);
or U520 (N_520,In_1111,In_331);
xnor U521 (N_521,In_1389,In_982);
nand U522 (N_522,In_588,In_90);
or U523 (N_523,In_162,In_1289);
and U524 (N_524,In_528,In_1125);
nand U525 (N_525,In_551,In_1226);
or U526 (N_526,In_35,In_328);
nor U527 (N_527,In_1329,In_582);
nor U528 (N_528,In_1313,In_580);
xor U529 (N_529,In_604,In_596);
nor U530 (N_530,In_707,In_1466);
nor U531 (N_531,In_529,In_753);
xnor U532 (N_532,In_709,In_97);
nand U533 (N_533,In_1395,In_469);
nor U534 (N_534,In_1173,In_250);
nand U535 (N_535,In_1449,In_179);
or U536 (N_536,In_147,In_161);
nand U537 (N_537,In_1204,In_1424);
nor U538 (N_538,In_714,In_497);
nand U539 (N_539,In_2,In_402);
and U540 (N_540,In_1046,In_501);
nor U541 (N_541,In_1196,In_360);
and U542 (N_542,In_776,In_852);
or U543 (N_543,In_1188,In_917);
xnor U544 (N_544,In_911,In_445);
and U545 (N_545,In_536,In_57);
nor U546 (N_546,In_1018,In_697);
nor U547 (N_547,In_1094,In_1422);
or U548 (N_548,In_29,In_921);
and U549 (N_549,In_1403,In_874);
xnor U550 (N_550,In_11,In_1090);
nor U551 (N_551,In_399,In_742);
xnor U552 (N_552,In_1361,In_851);
xor U553 (N_553,In_433,In_1456);
nand U554 (N_554,In_1349,In_26);
nand U555 (N_555,In_1139,In_1355);
nor U556 (N_556,In_559,In_894);
nand U557 (N_557,In_1242,In_683);
nand U558 (N_558,In_1310,In_708);
xnor U559 (N_559,In_676,In_645);
xnor U560 (N_560,In_1429,In_562);
nand U561 (N_561,In_741,In_447);
nor U562 (N_562,In_1052,In_724);
xor U563 (N_563,In_494,In_88);
or U564 (N_564,In_215,In_1314);
or U565 (N_565,In_1377,In_1030);
and U566 (N_566,In_810,In_430);
xnor U567 (N_567,In_211,In_372);
nand U568 (N_568,In_875,In_25);
or U569 (N_569,In_578,In_1352);
and U570 (N_570,In_686,In_153);
or U571 (N_571,In_341,In_301);
xnor U572 (N_572,In_952,In_92);
nand U573 (N_573,In_706,In_124);
nand U574 (N_574,In_1207,In_947);
nor U575 (N_575,In_1104,In_986);
or U576 (N_576,In_942,In_1150);
nor U577 (N_577,In_862,In_1096);
xnor U578 (N_578,In_181,In_719);
and U579 (N_579,In_964,In_1427);
nor U580 (N_580,In_828,In_209);
and U581 (N_581,In_76,In_872);
and U582 (N_582,In_1334,In_85);
or U583 (N_583,In_1298,In_487);
xor U584 (N_584,In_1230,In_1202);
nor U585 (N_585,In_241,In_716);
and U586 (N_586,In_833,In_895);
and U587 (N_587,In_1468,In_1383);
or U588 (N_588,In_649,In_848);
or U589 (N_589,In_1166,In_1217);
xor U590 (N_590,In_468,In_397);
nand U591 (N_591,In_1457,In_653);
or U592 (N_592,In_779,In_1229);
nand U593 (N_593,In_564,In_448);
nand U594 (N_594,In_1250,In_990);
xor U595 (N_595,In_1266,In_319);
xnor U596 (N_596,In_538,In_773);
nand U597 (N_597,In_170,In_548);
and U598 (N_598,In_651,In_622);
xor U599 (N_599,In_1218,In_1113);
or U600 (N_600,In_252,In_955);
nor U601 (N_601,In_226,In_77);
xor U602 (N_602,In_521,In_7);
xor U603 (N_603,In_527,In_613);
and U604 (N_604,In_204,In_110);
nand U605 (N_605,In_900,In_1253);
and U606 (N_606,In_1467,In_1346);
and U607 (N_607,In_260,In_499);
or U608 (N_608,In_1415,In_1362);
or U609 (N_609,In_1058,In_1308);
nand U610 (N_610,In_311,In_465);
nand U611 (N_611,In_1138,In_1323);
and U612 (N_612,In_1124,In_563);
nor U613 (N_613,In_725,In_771);
nand U614 (N_614,In_1416,In_1324);
xnor U615 (N_615,In_1318,In_292);
nor U616 (N_616,In_610,In_133);
or U617 (N_617,In_1441,In_216);
xnor U618 (N_618,In_134,In_755);
nor U619 (N_619,In_440,In_938);
nand U620 (N_620,In_539,In_679);
xnor U621 (N_621,In_857,In_1029);
xor U622 (N_622,In_1339,In_513);
or U623 (N_623,In_275,In_1033);
or U624 (N_624,In_1212,In_1325);
and U625 (N_625,In_915,In_791);
xor U626 (N_626,In_1228,In_66);
nor U627 (N_627,In_991,In_1410);
and U628 (N_628,In_151,In_599);
nor U629 (N_629,In_1338,In_1097);
xnor U630 (N_630,In_765,In_927);
nor U631 (N_631,In_995,In_892);
or U632 (N_632,In_1404,In_357);
nand U633 (N_633,In_602,In_840);
nand U634 (N_634,In_266,In_780);
or U635 (N_635,In_1471,In_1465);
xnor U636 (N_636,In_459,In_449);
nand U637 (N_637,In_5,In_1048);
or U638 (N_638,In_743,In_265);
and U639 (N_639,In_268,In_232);
xor U640 (N_640,In_1343,In_463);
or U641 (N_641,In_1255,In_1335);
and U642 (N_642,In_1278,In_1068);
nand U643 (N_643,In_1240,In_916);
nor U644 (N_644,In_1320,In_535);
nand U645 (N_645,In_509,In_1458);
and U646 (N_646,In_654,In_1292);
nor U647 (N_647,In_860,In_1076);
xor U648 (N_648,In_356,In_1197);
nand U649 (N_649,In_605,In_392);
nor U650 (N_650,In_552,In_1272);
nor U651 (N_651,In_1487,In_804);
nand U652 (N_652,In_1494,In_748);
nand U653 (N_653,In_1432,In_47);
xnor U654 (N_654,In_195,In_738);
nand U655 (N_655,In_790,In_32);
nand U656 (N_656,In_913,In_438);
nor U657 (N_657,In_1129,In_1493);
nor U658 (N_658,In_1375,In_411);
or U659 (N_659,In_1428,In_641);
or U660 (N_660,In_1462,In_84);
xor U661 (N_661,In_799,In_45);
xnor U662 (N_662,In_1411,In_197);
and U663 (N_663,In_502,In_558);
xor U664 (N_664,In_347,In_316);
nor U665 (N_665,In_385,In_369);
or U666 (N_666,In_823,In_489);
nand U667 (N_667,In_586,In_1216);
xor U668 (N_668,In_567,In_396);
and U669 (N_669,In_1178,In_693);
nand U670 (N_670,In_787,In_401);
or U671 (N_671,In_880,In_631);
nand U672 (N_672,In_889,In_960);
xnor U673 (N_673,In_793,In_224);
xor U674 (N_674,In_69,In_668);
and U675 (N_675,In_1367,In_1391);
and U676 (N_676,In_207,In_1477);
nor U677 (N_677,In_720,In_1039);
xor U678 (N_678,In_8,In_673);
nor U679 (N_679,In_1365,In_1285);
nor U680 (N_680,In_234,In_80);
and U681 (N_681,In_1390,In_1182);
xnor U682 (N_682,In_966,In_200);
nand U683 (N_683,In_721,In_1176);
or U684 (N_684,In_893,In_460);
xnor U685 (N_685,In_158,In_1071);
nor U686 (N_686,In_1280,In_1022);
or U687 (N_687,In_1356,In_1452);
nand U688 (N_688,In_597,In_1020);
or U689 (N_689,In_774,In_1198);
and U690 (N_690,In_1099,In_1083);
and U691 (N_691,In_1311,In_1498);
nor U692 (N_692,In_1263,In_1114);
or U693 (N_693,In_608,In_383);
xor U694 (N_694,In_1087,In_573);
nand U695 (N_695,In_284,In_540);
xnor U696 (N_696,In_555,In_303);
xnor U697 (N_697,In_441,In_545);
and U698 (N_698,In_410,In_1300);
and U699 (N_699,In_898,In_1213);
nor U700 (N_700,In_1270,In_1309);
and U701 (N_701,In_167,In_165);
or U702 (N_702,In_10,In_1496);
nand U703 (N_703,In_1006,In_1088);
or U704 (N_704,In_712,In_866);
nor U705 (N_705,In_692,In_454);
nor U706 (N_706,In_1413,In_457);
and U707 (N_707,In_1170,In_520);
nor U708 (N_708,In_498,In_1434);
xnor U709 (N_709,In_1284,In_844);
and U710 (N_710,In_1482,In_590);
or U711 (N_711,In_1257,In_1384);
nor U712 (N_712,In_1141,In_566);
and U713 (N_713,In_451,In_1420);
nand U714 (N_714,In_1364,In_239);
or U715 (N_715,In_1396,In_1262);
nand U716 (N_716,In_756,In_125);
or U717 (N_717,In_18,In_363);
nand U718 (N_718,In_998,In_1369);
xor U719 (N_719,In_667,In_1473);
and U720 (N_720,In_788,In_876);
xor U721 (N_721,In_1078,In_1134);
nor U722 (N_722,In_1439,In_850);
or U723 (N_723,In_1374,In_194);
and U724 (N_724,In_816,In_1293);
or U725 (N_725,In_176,In_1149);
nor U726 (N_726,In_221,In_614);
or U727 (N_727,In_684,In_815);
xor U728 (N_728,In_1080,In_1185);
nor U729 (N_729,In_985,In_119);
xor U730 (N_730,In_394,In_192);
or U731 (N_731,In_786,In_1282);
nor U732 (N_732,In_243,In_1273);
and U733 (N_733,In_22,In_1448);
or U734 (N_734,In_1186,In_46);
or U735 (N_735,In_1382,In_503);
nand U736 (N_736,In_795,In_329);
and U737 (N_737,In_616,In_1492);
nor U738 (N_738,In_541,In_1286);
or U739 (N_739,In_1371,In_223);
and U740 (N_740,In_180,In_244);
nand U741 (N_741,In_710,In_1357);
nand U742 (N_742,In_1063,In_858);
nand U743 (N_743,In_1499,In_695);
xor U744 (N_744,In_1003,In_822);
or U745 (N_745,In_1154,In_1119);
xor U746 (N_746,In_63,In_1317);
and U747 (N_747,In_1435,In_336);
xnor U748 (N_748,In_820,In_9);
or U749 (N_749,In_886,In_227);
and U750 (N_750,In_837,In_794);
nor U751 (N_751,In_801,In_883);
nand U752 (N_752,In_1214,In_454);
or U753 (N_753,In_863,In_508);
xor U754 (N_754,In_827,In_1464);
xnor U755 (N_755,In_1308,In_23);
or U756 (N_756,In_955,In_904);
xnor U757 (N_757,In_735,In_623);
or U758 (N_758,In_555,In_791);
xnor U759 (N_759,In_621,In_1368);
or U760 (N_760,In_569,In_1341);
or U761 (N_761,In_1272,In_512);
nand U762 (N_762,In_975,In_157);
and U763 (N_763,In_299,In_799);
nor U764 (N_764,In_1102,In_1091);
nor U765 (N_765,In_570,In_409);
or U766 (N_766,In_660,In_663);
xnor U767 (N_767,In_1222,In_864);
or U768 (N_768,In_827,In_363);
xor U769 (N_769,In_1276,In_182);
or U770 (N_770,In_189,In_264);
nor U771 (N_771,In_1286,In_266);
nor U772 (N_772,In_720,In_1290);
and U773 (N_773,In_1054,In_51);
nor U774 (N_774,In_442,In_1121);
nor U775 (N_775,In_574,In_581);
nand U776 (N_776,In_1022,In_797);
and U777 (N_777,In_761,In_663);
or U778 (N_778,In_287,In_791);
nor U779 (N_779,In_1200,In_597);
nand U780 (N_780,In_282,In_902);
nor U781 (N_781,In_157,In_1114);
or U782 (N_782,In_157,In_630);
or U783 (N_783,In_1280,In_396);
nand U784 (N_784,In_1300,In_1030);
and U785 (N_785,In_1329,In_205);
nor U786 (N_786,In_514,In_525);
nor U787 (N_787,In_378,In_751);
nor U788 (N_788,In_613,In_1316);
or U789 (N_789,In_601,In_955);
xor U790 (N_790,In_402,In_758);
or U791 (N_791,In_552,In_1345);
nand U792 (N_792,In_287,In_606);
nand U793 (N_793,In_1017,In_260);
nor U794 (N_794,In_261,In_270);
nor U795 (N_795,In_858,In_185);
nand U796 (N_796,In_151,In_1334);
or U797 (N_797,In_480,In_1000);
and U798 (N_798,In_522,In_1397);
nand U799 (N_799,In_519,In_891);
nand U800 (N_800,In_36,In_625);
nand U801 (N_801,In_689,In_488);
xor U802 (N_802,In_409,In_1093);
and U803 (N_803,In_717,In_1089);
xor U804 (N_804,In_1279,In_371);
and U805 (N_805,In_1199,In_756);
xor U806 (N_806,In_387,In_424);
nor U807 (N_807,In_492,In_770);
nor U808 (N_808,In_1400,In_651);
nand U809 (N_809,In_1272,In_594);
or U810 (N_810,In_778,In_1291);
and U811 (N_811,In_1185,In_1123);
nand U812 (N_812,In_1409,In_52);
or U813 (N_813,In_1469,In_402);
xnor U814 (N_814,In_687,In_156);
and U815 (N_815,In_310,In_1364);
nor U816 (N_816,In_615,In_1108);
nor U817 (N_817,In_1057,In_980);
nand U818 (N_818,In_752,In_1199);
nor U819 (N_819,In_1412,In_948);
nor U820 (N_820,In_623,In_1495);
nand U821 (N_821,In_343,In_1013);
xnor U822 (N_822,In_814,In_707);
nand U823 (N_823,In_418,In_252);
xnor U824 (N_824,In_1230,In_761);
or U825 (N_825,In_77,In_448);
or U826 (N_826,In_1459,In_547);
or U827 (N_827,In_25,In_1288);
and U828 (N_828,In_1212,In_1);
or U829 (N_829,In_1458,In_1006);
nor U830 (N_830,In_457,In_1294);
xor U831 (N_831,In_828,In_1440);
nand U832 (N_832,In_1413,In_3);
or U833 (N_833,In_945,In_1248);
nand U834 (N_834,In_95,In_255);
xnor U835 (N_835,In_1058,In_829);
and U836 (N_836,In_777,In_1399);
and U837 (N_837,In_291,In_684);
and U838 (N_838,In_1405,In_628);
xnor U839 (N_839,In_1253,In_392);
nor U840 (N_840,In_700,In_95);
nor U841 (N_841,In_858,In_789);
nand U842 (N_842,In_1297,In_485);
nand U843 (N_843,In_1298,In_450);
nor U844 (N_844,In_1093,In_668);
or U845 (N_845,In_1024,In_962);
nand U846 (N_846,In_210,In_197);
nor U847 (N_847,In_1099,In_64);
nand U848 (N_848,In_73,In_1478);
nor U849 (N_849,In_274,In_518);
xnor U850 (N_850,In_469,In_1140);
xor U851 (N_851,In_850,In_1363);
nor U852 (N_852,In_137,In_476);
xnor U853 (N_853,In_788,In_1283);
nor U854 (N_854,In_1279,In_1483);
nand U855 (N_855,In_319,In_960);
nand U856 (N_856,In_1485,In_1104);
nor U857 (N_857,In_153,In_1102);
nor U858 (N_858,In_786,In_1496);
and U859 (N_859,In_458,In_1414);
nand U860 (N_860,In_1220,In_1258);
and U861 (N_861,In_412,In_697);
nand U862 (N_862,In_764,In_1268);
or U863 (N_863,In_504,In_1044);
nand U864 (N_864,In_524,In_155);
nor U865 (N_865,In_628,In_691);
or U866 (N_866,In_1284,In_832);
nand U867 (N_867,In_170,In_727);
and U868 (N_868,In_59,In_1418);
and U869 (N_869,In_1279,In_1160);
nand U870 (N_870,In_174,In_403);
nand U871 (N_871,In_505,In_566);
nor U872 (N_872,In_947,In_795);
and U873 (N_873,In_436,In_1085);
nand U874 (N_874,In_937,In_556);
and U875 (N_875,In_813,In_207);
and U876 (N_876,In_877,In_911);
and U877 (N_877,In_337,In_1353);
nand U878 (N_878,In_669,In_25);
nor U879 (N_879,In_398,In_354);
nand U880 (N_880,In_875,In_1173);
or U881 (N_881,In_583,In_99);
nand U882 (N_882,In_201,In_658);
and U883 (N_883,In_776,In_826);
or U884 (N_884,In_376,In_1122);
and U885 (N_885,In_1235,In_1308);
nor U886 (N_886,In_825,In_476);
and U887 (N_887,In_439,In_885);
or U888 (N_888,In_1331,In_379);
xnor U889 (N_889,In_1357,In_103);
and U890 (N_890,In_414,In_37);
nor U891 (N_891,In_746,In_284);
nor U892 (N_892,In_22,In_961);
nand U893 (N_893,In_185,In_303);
nor U894 (N_894,In_1012,In_151);
and U895 (N_895,In_549,In_502);
xnor U896 (N_896,In_224,In_558);
nor U897 (N_897,In_806,In_333);
and U898 (N_898,In_464,In_304);
and U899 (N_899,In_1362,In_256);
nand U900 (N_900,In_1018,In_1292);
nor U901 (N_901,In_406,In_159);
nor U902 (N_902,In_989,In_687);
nor U903 (N_903,In_1335,In_60);
and U904 (N_904,In_974,In_388);
nor U905 (N_905,In_406,In_602);
nand U906 (N_906,In_549,In_1252);
or U907 (N_907,In_1343,In_1039);
or U908 (N_908,In_1420,In_896);
xor U909 (N_909,In_998,In_1425);
xor U910 (N_910,In_969,In_673);
and U911 (N_911,In_1240,In_205);
nand U912 (N_912,In_380,In_54);
xor U913 (N_913,In_1480,In_1055);
nand U914 (N_914,In_737,In_691);
and U915 (N_915,In_722,In_1129);
nand U916 (N_916,In_1110,In_660);
and U917 (N_917,In_132,In_1062);
nand U918 (N_918,In_1186,In_1488);
and U919 (N_919,In_1002,In_1347);
xnor U920 (N_920,In_1215,In_407);
xnor U921 (N_921,In_928,In_364);
and U922 (N_922,In_387,In_1165);
nand U923 (N_923,In_1346,In_1192);
xor U924 (N_924,In_474,In_490);
nand U925 (N_925,In_801,In_1313);
nand U926 (N_926,In_715,In_209);
nand U927 (N_927,In_2,In_1056);
nor U928 (N_928,In_568,In_1393);
nand U929 (N_929,In_862,In_532);
and U930 (N_930,In_969,In_270);
or U931 (N_931,In_485,In_799);
nor U932 (N_932,In_20,In_695);
xnor U933 (N_933,In_317,In_902);
xor U934 (N_934,In_775,In_187);
nor U935 (N_935,In_635,In_70);
or U936 (N_936,In_1317,In_386);
and U937 (N_937,In_1015,In_70);
xor U938 (N_938,In_138,In_886);
or U939 (N_939,In_230,In_366);
nor U940 (N_940,In_1246,In_414);
and U941 (N_941,In_744,In_963);
nor U942 (N_942,In_1433,In_181);
and U943 (N_943,In_231,In_488);
xor U944 (N_944,In_561,In_153);
and U945 (N_945,In_1399,In_374);
nand U946 (N_946,In_64,In_459);
nand U947 (N_947,In_1325,In_1375);
or U948 (N_948,In_918,In_902);
nand U949 (N_949,In_343,In_1078);
nor U950 (N_950,In_612,In_944);
nand U951 (N_951,In_1237,In_136);
xnor U952 (N_952,In_1346,In_1468);
or U953 (N_953,In_782,In_781);
xor U954 (N_954,In_1095,In_634);
nand U955 (N_955,In_52,In_435);
and U956 (N_956,In_1329,In_879);
xnor U957 (N_957,In_829,In_847);
or U958 (N_958,In_202,In_291);
or U959 (N_959,In_1422,In_1196);
or U960 (N_960,In_1086,In_196);
nor U961 (N_961,In_1331,In_196);
or U962 (N_962,In_864,In_1153);
xnor U963 (N_963,In_165,In_259);
nor U964 (N_964,In_369,In_430);
nand U965 (N_965,In_1158,In_1132);
or U966 (N_966,In_650,In_144);
nand U967 (N_967,In_547,In_1181);
or U968 (N_968,In_1111,In_1205);
xor U969 (N_969,In_701,In_6);
and U970 (N_970,In_649,In_1419);
or U971 (N_971,In_875,In_345);
nor U972 (N_972,In_419,In_911);
or U973 (N_973,In_991,In_1174);
nand U974 (N_974,In_1273,In_137);
xor U975 (N_975,In_700,In_1346);
and U976 (N_976,In_1206,In_1122);
xor U977 (N_977,In_182,In_750);
xor U978 (N_978,In_803,In_523);
nor U979 (N_979,In_1240,In_214);
nor U980 (N_980,In_731,In_30);
nor U981 (N_981,In_1300,In_776);
or U982 (N_982,In_1353,In_982);
xnor U983 (N_983,In_1036,In_561);
or U984 (N_984,In_725,In_590);
and U985 (N_985,In_851,In_1277);
nand U986 (N_986,In_1405,In_22);
xor U987 (N_987,In_100,In_242);
and U988 (N_988,In_1201,In_356);
nand U989 (N_989,In_240,In_686);
nand U990 (N_990,In_467,In_21);
or U991 (N_991,In_678,In_856);
and U992 (N_992,In_56,In_62);
nand U993 (N_993,In_467,In_1391);
xnor U994 (N_994,In_562,In_1398);
nand U995 (N_995,In_272,In_591);
nor U996 (N_996,In_149,In_1028);
xor U997 (N_997,In_1259,In_233);
nor U998 (N_998,In_410,In_745);
or U999 (N_999,In_276,In_954);
xnor U1000 (N_1000,In_516,In_1273);
nand U1001 (N_1001,In_815,In_629);
and U1002 (N_1002,In_253,In_1225);
nand U1003 (N_1003,In_513,In_967);
xor U1004 (N_1004,In_873,In_852);
xor U1005 (N_1005,In_1384,In_10);
xor U1006 (N_1006,In_222,In_1003);
nor U1007 (N_1007,In_1283,In_1400);
xnor U1008 (N_1008,In_597,In_25);
and U1009 (N_1009,In_472,In_1168);
and U1010 (N_1010,In_509,In_760);
or U1011 (N_1011,In_84,In_928);
or U1012 (N_1012,In_244,In_428);
nand U1013 (N_1013,In_971,In_722);
nor U1014 (N_1014,In_1286,In_513);
nand U1015 (N_1015,In_439,In_214);
and U1016 (N_1016,In_1079,In_980);
or U1017 (N_1017,In_683,In_672);
or U1018 (N_1018,In_502,In_212);
nand U1019 (N_1019,In_976,In_1123);
nand U1020 (N_1020,In_1059,In_691);
nand U1021 (N_1021,In_869,In_56);
or U1022 (N_1022,In_898,In_530);
xnor U1023 (N_1023,In_1342,In_836);
nand U1024 (N_1024,In_1255,In_719);
nand U1025 (N_1025,In_1464,In_1234);
nor U1026 (N_1026,In_1014,In_659);
xnor U1027 (N_1027,In_723,In_205);
xor U1028 (N_1028,In_922,In_1268);
xor U1029 (N_1029,In_524,In_359);
and U1030 (N_1030,In_44,In_1323);
xnor U1031 (N_1031,In_136,In_822);
xnor U1032 (N_1032,In_21,In_294);
or U1033 (N_1033,In_305,In_1003);
or U1034 (N_1034,In_641,In_363);
xor U1035 (N_1035,In_696,In_1425);
or U1036 (N_1036,In_582,In_1110);
nand U1037 (N_1037,In_474,In_1087);
xor U1038 (N_1038,In_613,In_1312);
xnor U1039 (N_1039,In_637,In_57);
xor U1040 (N_1040,In_404,In_1130);
nor U1041 (N_1041,In_1261,In_451);
nand U1042 (N_1042,In_908,In_1182);
nand U1043 (N_1043,In_154,In_672);
nor U1044 (N_1044,In_936,In_552);
nor U1045 (N_1045,In_1446,In_712);
nor U1046 (N_1046,In_218,In_679);
or U1047 (N_1047,In_1429,In_1133);
nand U1048 (N_1048,In_1275,In_35);
and U1049 (N_1049,In_188,In_288);
nand U1050 (N_1050,In_559,In_211);
nand U1051 (N_1051,In_72,In_693);
xnor U1052 (N_1052,In_542,In_311);
or U1053 (N_1053,In_696,In_104);
and U1054 (N_1054,In_197,In_1486);
nor U1055 (N_1055,In_564,In_62);
and U1056 (N_1056,In_873,In_15);
and U1057 (N_1057,In_104,In_633);
nor U1058 (N_1058,In_536,In_678);
xor U1059 (N_1059,In_730,In_1324);
nor U1060 (N_1060,In_593,In_1116);
nand U1061 (N_1061,In_480,In_1254);
nand U1062 (N_1062,In_394,In_189);
nor U1063 (N_1063,In_961,In_941);
or U1064 (N_1064,In_1153,In_1287);
and U1065 (N_1065,In_1182,In_1323);
nand U1066 (N_1066,In_1215,In_1110);
and U1067 (N_1067,In_734,In_857);
nor U1068 (N_1068,In_1212,In_1227);
xor U1069 (N_1069,In_74,In_981);
xnor U1070 (N_1070,In_1400,In_473);
or U1071 (N_1071,In_1028,In_914);
and U1072 (N_1072,In_183,In_1261);
nand U1073 (N_1073,In_798,In_777);
or U1074 (N_1074,In_1165,In_1263);
nor U1075 (N_1075,In_277,In_1181);
xor U1076 (N_1076,In_121,In_294);
nand U1077 (N_1077,In_1111,In_355);
nor U1078 (N_1078,In_1265,In_674);
nor U1079 (N_1079,In_1168,In_1472);
nand U1080 (N_1080,In_1409,In_436);
nor U1081 (N_1081,In_1487,In_481);
or U1082 (N_1082,In_1262,In_837);
nor U1083 (N_1083,In_880,In_210);
or U1084 (N_1084,In_730,In_1091);
and U1085 (N_1085,In_90,In_1127);
and U1086 (N_1086,In_765,In_526);
nand U1087 (N_1087,In_452,In_858);
nand U1088 (N_1088,In_389,In_944);
nand U1089 (N_1089,In_258,In_689);
and U1090 (N_1090,In_1113,In_1475);
nand U1091 (N_1091,In_572,In_122);
and U1092 (N_1092,In_1099,In_1052);
or U1093 (N_1093,In_1320,In_313);
nor U1094 (N_1094,In_641,In_1007);
xor U1095 (N_1095,In_950,In_448);
nand U1096 (N_1096,In_464,In_692);
xor U1097 (N_1097,In_1135,In_380);
xor U1098 (N_1098,In_1017,In_156);
or U1099 (N_1099,In_1338,In_1269);
xor U1100 (N_1100,In_1492,In_1292);
or U1101 (N_1101,In_87,In_1430);
or U1102 (N_1102,In_323,In_1323);
nand U1103 (N_1103,In_307,In_128);
and U1104 (N_1104,In_176,In_1167);
nand U1105 (N_1105,In_1112,In_1345);
and U1106 (N_1106,In_441,In_782);
xor U1107 (N_1107,In_320,In_966);
nand U1108 (N_1108,In_400,In_992);
nand U1109 (N_1109,In_192,In_1342);
xnor U1110 (N_1110,In_377,In_1480);
or U1111 (N_1111,In_1057,In_36);
and U1112 (N_1112,In_393,In_135);
or U1113 (N_1113,In_32,In_37);
xnor U1114 (N_1114,In_1087,In_292);
xor U1115 (N_1115,In_152,In_1439);
nand U1116 (N_1116,In_784,In_1025);
xnor U1117 (N_1117,In_620,In_451);
and U1118 (N_1118,In_321,In_1331);
xnor U1119 (N_1119,In_1415,In_86);
nand U1120 (N_1120,In_195,In_1145);
and U1121 (N_1121,In_385,In_115);
nand U1122 (N_1122,In_168,In_1395);
nand U1123 (N_1123,In_409,In_399);
nor U1124 (N_1124,In_329,In_365);
nand U1125 (N_1125,In_1289,In_1391);
nor U1126 (N_1126,In_1322,In_726);
and U1127 (N_1127,In_688,In_207);
nor U1128 (N_1128,In_350,In_282);
and U1129 (N_1129,In_811,In_1119);
nor U1130 (N_1130,In_1448,In_819);
xnor U1131 (N_1131,In_1159,In_841);
and U1132 (N_1132,In_846,In_8);
nand U1133 (N_1133,In_211,In_948);
nand U1134 (N_1134,In_659,In_906);
xor U1135 (N_1135,In_824,In_128);
nand U1136 (N_1136,In_1402,In_563);
xnor U1137 (N_1137,In_1475,In_845);
or U1138 (N_1138,In_165,In_1367);
and U1139 (N_1139,In_794,In_51);
and U1140 (N_1140,In_225,In_37);
xnor U1141 (N_1141,In_315,In_1328);
or U1142 (N_1142,In_523,In_338);
xor U1143 (N_1143,In_233,In_1079);
nand U1144 (N_1144,In_311,In_1179);
or U1145 (N_1145,In_510,In_222);
nor U1146 (N_1146,In_682,In_297);
nor U1147 (N_1147,In_61,In_1168);
and U1148 (N_1148,In_97,In_1027);
xnor U1149 (N_1149,In_836,In_978);
xnor U1150 (N_1150,In_848,In_643);
or U1151 (N_1151,In_414,In_652);
nor U1152 (N_1152,In_568,In_750);
xnor U1153 (N_1153,In_495,In_1360);
nand U1154 (N_1154,In_564,In_618);
nand U1155 (N_1155,In_80,In_1471);
or U1156 (N_1156,In_144,In_203);
and U1157 (N_1157,In_1331,In_1421);
nand U1158 (N_1158,In_521,In_1482);
and U1159 (N_1159,In_797,In_1436);
nor U1160 (N_1160,In_1115,In_1354);
nor U1161 (N_1161,In_663,In_467);
nor U1162 (N_1162,In_234,In_790);
nor U1163 (N_1163,In_1290,In_562);
xor U1164 (N_1164,In_272,In_1468);
or U1165 (N_1165,In_239,In_323);
nand U1166 (N_1166,In_1173,In_1396);
nand U1167 (N_1167,In_378,In_58);
or U1168 (N_1168,In_1391,In_179);
or U1169 (N_1169,In_839,In_912);
nand U1170 (N_1170,In_593,In_201);
xnor U1171 (N_1171,In_1305,In_932);
and U1172 (N_1172,In_126,In_328);
nand U1173 (N_1173,In_1330,In_749);
nor U1174 (N_1174,In_316,In_1195);
nor U1175 (N_1175,In_774,In_99);
or U1176 (N_1176,In_119,In_260);
or U1177 (N_1177,In_807,In_916);
and U1178 (N_1178,In_855,In_1070);
or U1179 (N_1179,In_1283,In_850);
nand U1180 (N_1180,In_40,In_893);
nor U1181 (N_1181,In_1014,In_882);
xnor U1182 (N_1182,In_1315,In_69);
or U1183 (N_1183,In_527,In_1361);
and U1184 (N_1184,In_1490,In_623);
xor U1185 (N_1185,In_217,In_1473);
and U1186 (N_1186,In_296,In_1091);
xor U1187 (N_1187,In_1492,In_435);
nor U1188 (N_1188,In_1471,In_1062);
xor U1189 (N_1189,In_76,In_1424);
and U1190 (N_1190,In_89,In_1009);
xor U1191 (N_1191,In_1495,In_1452);
and U1192 (N_1192,In_276,In_862);
or U1193 (N_1193,In_488,In_1328);
or U1194 (N_1194,In_643,In_309);
nand U1195 (N_1195,In_565,In_576);
and U1196 (N_1196,In_760,In_1479);
or U1197 (N_1197,In_139,In_1139);
or U1198 (N_1198,In_1234,In_622);
nand U1199 (N_1199,In_607,In_428);
xor U1200 (N_1200,In_1240,In_674);
nor U1201 (N_1201,In_876,In_296);
nor U1202 (N_1202,In_854,In_1168);
and U1203 (N_1203,In_651,In_552);
xnor U1204 (N_1204,In_33,In_978);
xnor U1205 (N_1205,In_1,In_1088);
xnor U1206 (N_1206,In_918,In_416);
nand U1207 (N_1207,In_575,In_303);
or U1208 (N_1208,In_715,In_1491);
nor U1209 (N_1209,In_333,In_378);
and U1210 (N_1210,In_1294,In_332);
and U1211 (N_1211,In_47,In_630);
nor U1212 (N_1212,In_236,In_941);
nand U1213 (N_1213,In_229,In_837);
xnor U1214 (N_1214,In_1133,In_229);
nand U1215 (N_1215,In_724,In_621);
nor U1216 (N_1216,In_633,In_1333);
nand U1217 (N_1217,In_1394,In_38);
and U1218 (N_1218,In_825,In_951);
nand U1219 (N_1219,In_332,In_884);
nor U1220 (N_1220,In_136,In_394);
nand U1221 (N_1221,In_57,In_384);
or U1222 (N_1222,In_470,In_771);
xor U1223 (N_1223,In_803,In_532);
xnor U1224 (N_1224,In_1290,In_435);
or U1225 (N_1225,In_354,In_711);
xor U1226 (N_1226,In_311,In_120);
nand U1227 (N_1227,In_560,In_18);
nor U1228 (N_1228,In_765,In_1489);
and U1229 (N_1229,In_387,In_392);
xor U1230 (N_1230,In_501,In_238);
or U1231 (N_1231,In_698,In_1447);
nor U1232 (N_1232,In_1398,In_1152);
or U1233 (N_1233,In_897,In_67);
nor U1234 (N_1234,In_918,In_456);
nand U1235 (N_1235,In_1394,In_1379);
nand U1236 (N_1236,In_85,In_1180);
and U1237 (N_1237,In_1443,In_802);
nand U1238 (N_1238,In_120,In_1151);
and U1239 (N_1239,In_204,In_1058);
nand U1240 (N_1240,In_855,In_1090);
or U1241 (N_1241,In_697,In_721);
xnor U1242 (N_1242,In_1409,In_16);
and U1243 (N_1243,In_1159,In_1470);
and U1244 (N_1244,In_812,In_1218);
nor U1245 (N_1245,In_624,In_1443);
or U1246 (N_1246,In_818,In_270);
and U1247 (N_1247,In_288,In_178);
xnor U1248 (N_1248,In_847,In_680);
and U1249 (N_1249,In_437,In_755);
or U1250 (N_1250,In_487,In_1343);
or U1251 (N_1251,In_891,In_12);
or U1252 (N_1252,In_711,In_1287);
xor U1253 (N_1253,In_939,In_47);
and U1254 (N_1254,In_443,In_252);
nand U1255 (N_1255,In_1225,In_332);
and U1256 (N_1256,In_188,In_1270);
xnor U1257 (N_1257,In_163,In_702);
and U1258 (N_1258,In_192,In_1480);
nand U1259 (N_1259,In_77,In_1433);
xor U1260 (N_1260,In_526,In_86);
or U1261 (N_1261,In_279,In_815);
or U1262 (N_1262,In_877,In_988);
nand U1263 (N_1263,In_773,In_652);
or U1264 (N_1264,In_239,In_341);
or U1265 (N_1265,In_823,In_745);
xor U1266 (N_1266,In_983,In_127);
nand U1267 (N_1267,In_399,In_1008);
nand U1268 (N_1268,In_305,In_1490);
nand U1269 (N_1269,In_1167,In_787);
or U1270 (N_1270,In_1213,In_341);
nand U1271 (N_1271,In_835,In_1434);
or U1272 (N_1272,In_627,In_1372);
or U1273 (N_1273,In_582,In_734);
nand U1274 (N_1274,In_764,In_572);
and U1275 (N_1275,In_918,In_923);
and U1276 (N_1276,In_285,In_52);
nor U1277 (N_1277,In_269,In_1003);
xor U1278 (N_1278,In_960,In_664);
nor U1279 (N_1279,In_986,In_227);
xnor U1280 (N_1280,In_1220,In_1343);
and U1281 (N_1281,In_395,In_399);
and U1282 (N_1282,In_506,In_1369);
or U1283 (N_1283,In_218,In_641);
nand U1284 (N_1284,In_496,In_278);
nor U1285 (N_1285,In_593,In_595);
and U1286 (N_1286,In_1266,In_227);
nand U1287 (N_1287,In_1039,In_1209);
nand U1288 (N_1288,In_122,In_1164);
and U1289 (N_1289,In_522,In_1298);
nor U1290 (N_1290,In_225,In_920);
nand U1291 (N_1291,In_1330,In_468);
or U1292 (N_1292,In_227,In_1068);
xnor U1293 (N_1293,In_991,In_416);
nand U1294 (N_1294,In_248,In_786);
nand U1295 (N_1295,In_643,In_1162);
nand U1296 (N_1296,In_956,In_392);
nand U1297 (N_1297,In_724,In_660);
xnor U1298 (N_1298,In_1230,In_1312);
and U1299 (N_1299,In_1328,In_1382);
nand U1300 (N_1300,In_295,In_1162);
nand U1301 (N_1301,In_505,In_463);
nor U1302 (N_1302,In_1250,In_1015);
or U1303 (N_1303,In_1422,In_401);
or U1304 (N_1304,In_134,In_992);
nor U1305 (N_1305,In_999,In_477);
or U1306 (N_1306,In_176,In_1463);
nand U1307 (N_1307,In_900,In_432);
nand U1308 (N_1308,In_305,In_1203);
or U1309 (N_1309,In_604,In_1233);
nand U1310 (N_1310,In_1448,In_1492);
xnor U1311 (N_1311,In_234,In_1124);
nor U1312 (N_1312,In_50,In_1202);
nand U1313 (N_1313,In_682,In_1185);
and U1314 (N_1314,In_1079,In_833);
and U1315 (N_1315,In_813,In_864);
or U1316 (N_1316,In_1366,In_381);
or U1317 (N_1317,In_288,In_461);
or U1318 (N_1318,In_963,In_95);
nor U1319 (N_1319,In_816,In_1099);
nand U1320 (N_1320,In_1149,In_524);
or U1321 (N_1321,In_767,In_1342);
or U1322 (N_1322,In_566,In_1213);
xor U1323 (N_1323,In_1284,In_671);
and U1324 (N_1324,In_378,In_1476);
nor U1325 (N_1325,In_1026,In_1414);
xnor U1326 (N_1326,In_396,In_331);
and U1327 (N_1327,In_877,In_1452);
xor U1328 (N_1328,In_485,In_396);
and U1329 (N_1329,In_241,In_780);
or U1330 (N_1330,In_1063,In_1235);
nor U1331 (N_1331,In_114,In_1243);
or U1332 (N_1332,In_761,In_707);
xor U1333 (N_1333,In_1308,In_187);
or U1334 (N_1334,In_525,In_74);
or U1335 (N_1335,In_95,In_134);
or U1336 (N_1336,In_670,In_26);
nor U1337 (N_1337,In_50,In_159);
or U1338 (N_1338,In_766,In_391);
and U1339 (N_1339,In_893,In_876);
or U1340 (N_1340,In_1093,In_977);
or U1341 (N_1341,In_167,In_694);
xor U1342 (N_1342,In_1489,In_1104);
or U1343 (N_1343,In_387,In_577);
nor U1344 (N_1344,In_468,In_8);
nand U1345 (N_1345,In_553,In_1302);
xor U1346 (N_1346,In_412,In_611);
nor U1347 (N_1347,In_913,In_728);
nand U1348 (N_1348,In_7,In_423);
xor U1349 (N_1349,In_1218,In_1467);
and U1350 (N_1350,In_723,In_1377);
nor U1351 (N_1351,In_233,In_880);
nand U1352 (N_1352,In_84,In_1111);
xor U1353 (N_1353,In_660,In_1401);
xor U1354 (N_1354,In_806,In_667);
nor U1355 (N_1355,In_588,In_1054);
or U1356 (N_1356,In_1337,In_323);
and U1357 (N_1357,In_581,In_76);
nor U1358 (N_1358,In_448,In_57);
and U1359 (N_1359,In_838,In_1367);
or U1360 (N_1360,In_1110,In_1152);
xor U1361 (N_1361,In_1484,In_422);
or U1362 (N_1362,In_266,In_74);
xor U1363 (N_1363,In_1449,In_490);
xor U1364 (N_1364,In_125,In_1189);
nor U1365 (N_1365,In_1086,In_854);
and U1366 (N_1366,In_921,In_991);
nor U1367 (N_1367,In_1038,In_1291);
nand U1368 (N_1368,In_254,In_1045);
or U1369 (N_1369,In_351,In_6);
nand U1370 (N_1370,In_1013,In_284);
xnor U1371 (N_1371,In_46,In_1461);
and U1372 (N_1372,In_392,In_1278);
xor U1373 (N_1373,In_810,In_258);
or U1374 (N_1374,In_146,In_1047);
or U1375 (N_1375,In_89,In_285);
and U1376 (N_1376,In_102,In_217);
nand U1377 (N_1377,In_302,In_1302);
nor U1378 (N_1378,In_1286,In_934);
nand U1379 (N_1379,In_1400,In_764);
or U1380 (N_1380,In_779,In_483);
xnor U1381 (N_1381,In_470,In_772);
xor U1382 (N_1382,In_531,In_1001);
and U1383 (N_1383,In_272,In_1370);
xnor U1384 (N_1384,In_219,In_17);
and U1385 (N_1385,In_1055,In_226);
nor U1386 (N_1386,In_1297,In_914);
and U1387 (N_1387,In_1222,In_1068);
or U1388 (N_1388,In_1337,In_655);
nand U1389 (N_1389,In_493,In_1483);
nand U1390 (N_1390,In_99,In_905);
and U1391 (N_1391,In_249,In_1312);
nand U1392 (N_1392,In_961,In_1055);
nand U1393 (N_1393,In_67,In_1319);
xnor U1394 (N_1394,In_111,In_357);
nor U1395 (N_1395,In_137,In_412);
xor U1396 (N_1396,In_996,In_872);
nor U1397 (N_1397,In_785,In_76);
or U1398 (N_1398,In_95,In_374);
and U1399 (N_1399,In_375,In_996);
or U1400 (N_1400,In_1157,In_194);
and U1401 (N_1401,In_727,In_1471);
and U1402 (N_1402,In_126,In_814);
nor U1403 (N_1403,In_1471,In_431);
xnor U1404 (N_1404,In_495,In_273);
and U1405 (N_1405,In_1211,In_920);
or U1406 (N_1406,In_1271,In_1219);
nand U1407 (N_1407,In_1088,In_471);
nand U1408 (N_1408,In_589,In_227);
nor U1409 (N_1409,In_379,In_55);
nor U1410 (N_1410,In_299,In_1423);
and U1411 (N_1411,In_986,In_1188);
nor U1412 (N_1412,In_749,In_99);
or U1413 (N_1413,In_1361,In_1377);
xor U1414 (N_1414,In_184,In_260);
or U1415 (N_1415,In_687,In_244);
or U1416 (N_1416,In_1204,In_1318);
xor U1417 (N_1417,In_614,In_1082);
and U1418 (N_1418,In_716,In_1180);
or U1419 (N_1419,In_1397,In_943);
or U1420 (N_1420,In_1059,In_1422);
nor U1421 (N_1421,In_997,In_1436);
and U1422 (N_1422,In_593,In_76);
nand U1423 (N_1423,In_360,In_999);
xor U1424 (N_1424,In_700,In_937);
xor U1425 (N_1425,In_1035,In_528);
xnor U1426 (N_1426,In_1266,In_1145);
xnor U1427 (N_1427,In_498,In_546);
nor U1428 (N_1428,In_839,In_526);
and U1429 (N_1429,In_1252,In_625);
and U1430 (N_1430,In_1361,In_857);
or U1431 (N_1431,In_1289,In_1075);
and U1432 (N_1432,In_1301,In_1055);
nor U1433 (N_1433,In_1248,In_662);
nand U1434 (N_1434,In_275,In_641);
nor U1435 (N_1435,In_233,In_6);
nor U1436 (N_1436,In_718,In_457);
xor U1437 (N_1437,In_664,In_529);
nand U1438 (N_1438,In_20,In_838);
xor U1439 (N_1439,In_776,In_1098);
nor U1440 (N_1440,In_113,In_986);
or U1441 (N_1441,In_634,In_883);
and U1442 (N_1442,In_16,In_582);
nor U1443 (N_1443,In_187,In_345);
xor U1444 (N_1444,In_1375,In_1213);
nor U1445 (N_1445,In_950,In_763);
and U1446 (N_1446,In_341,In_813);
nand U1447 (N_1447,In_384,In_770);
xor U1448 (N_1448,In_1167,In_282);
xor U1449 (N_1449,In_339,In_924);
nor U1450 (N_1450,In_729,In_999);
and U1451 (N_1451,In_363,In_389);
nand U1452 (N_1452,In_1318,In_695);
nand U1453 (N_1453,In_1466,In_1088);
or U1454 (N_1454,In_11,In_403);
or U1455 (N_1455,In_712,In_1348);
xnor U1456 (N_1456,In_822,In_542);
nor U1457 (N_1457,In_404,In_955);
or U1458 (N_1458,In_950,In_936);
nor U1459 (N_1459,In_779,In_790);
nor U1460 (N_1460,In_698,In_990);
nand U1461 (N_1461,In_724,In_89);
or U1462 (N_1462,In_1357,In_1321);
nand U1463 (N_1463,In_255,In_231);
or U1464 (N_1464,In_316,In_1025);
xor U1465 (N_1465,In_576,In_1319);
xor U1466 (N_1466,In_575,In_944);
xor U1467 (N_1467,In_844,In_1064);
and U1468 (N_1468,In_70,In_851);
and U1469 (N_1469,In_366,In_74);
and U1470 (N_1470,In_560,In_1484);
or U1471 (N_1471,In_527,In_484);
nand U1472 (N_1472,In_552,In_1121);
nand U1473 (N_1473,In_306,In_80);
xnor U1474 (N_1474,In_1208,In_43);
or U1475 (N_1475,In_57,In_1144);
and U1476 (N_1476,In_826,In_1143);
and U1477 (N_1477,In_1219,In_496);
and U1478 (N_1478,In_1152,In_235);
and U1479 (N_1479,In_397,In_903);
xnor U1480 (N_1480,In_382,In_1454);
nor U1481 (N_1481,In_532,In_740);
nand U1482 (N_1482,In_431,In_1349);
xnor U1483 (N_1483,In_1053,In_536);
and U1484 (N_1484,In_272,In_839);
and U1485 (N_1485,In_1123,In_293);
xor U1486 (N_1486,In_40,In_413);
or U1487 (N_1487,In_152,In_1076);
xor U1488 (N_1488,In_1223,In_1484);
or U1489 (N_1489,In_821,In_1080);
and U1490 (N_1490,In_1313,In_769);
and U1491 (N_1491,In_645,In_1205);
and U1492 (N_1492,In_447,In_1493);
nand U1493 (N_1493,In_521,In_378);
nand U1494 (N_1494,In_611,In_353);
nand U1495 (N_1495,In_678,In_486);
nand U1496 (N_1496,In_216,In_766);
nand U1497 (N_1497,In_688,In_962);
and U1498 (N_1498,In_539,In_988);
nand U1499 (N_1499,In_1469,In_1043);
xnor U1500 (N_1500,In_1399,In_1058);
nand U1501 (N_1501,In_801,In_1110);
nand U1502 (N_1502,In_169,In_25);
and U1503 (N_1503,In_22,In_178);
nand U1504 (N_1504,In_956,In_656);
nand U1505 (N_1505,In_591,In_187);
and U1506 (N_1506,In_1192,In_360);
nand U1507 (N_1507,In_1465,In_617);
or U1508 (N_1508,In_749,In_211);
nand U1509 (N_1509,In_387,In_1249);
and U1510 (N_1510,In_1113,In_828);
nand U1511 (N_1511,In_1150,In_1388);
nand U1512 (N_1512,In_17,In_1001);
or U1513 (N_1513,In_187,In_444);
nand U1514 (N_1514,In_663,In_219);
nand U1515 (N_1515,In_342,In_469);
xor U1516 (N_1516,In_675,In_303);
nor U1517 (N_1517,In_540,In_277);
nor U1518 (N_1518,In_613,In_856);
xnor U1519 (N_1519,In_1008,In_954);
nor U1520 (N_1520,In_140,In_765);
nand U1521 (N_1521,In_80,In_348);
nor U1522 (N_1522,In_1200,In_585);
and U1523 (N_1523,In_89,In_217);
xnor U1524 (N_1524,In_546,In_577);
or U1525 (N_1525,In_247,In_656);
or U1526 (N_1526,In_1336,In_46);
or U1527 (N_1527,In_774,In_817);
nor U1528 (N_1528,In_1076,In_786);
or U1529 (N_1529,In_379,In_113);
nand U1530 (N_1530,In_834,In_908);
nor U1531 (N_1531,In_1128,In_1419);
nand U1532 (N_1532,In_265,In_54);
or U1533 (N_1533,In_547,In_1088);
and U1534 (N_1534,In_723,In_1307);
nand U1535 (N_1535,In_277,In_1119);
nand U1536 (N_1536,In_1433,In_1193);
xnor U1537 (N_1537,In_43,In_425);
nand U1538 (N_1538,In_383,In_39);
xor U1539 (N_1539,In_1263,In_737);
or U1540 (N_1540,In_751,In_960);
nor U1541 (N_1541,In_360,In_182);
nor U1542 (N_1542,In_918,In_1281);
nand U1543 (N_1543,In_1117,In_1228);
and U1544 (N_1544,In_197,In_1372);
or U1545 (N_1545,In_378,In_1456);
xor U1546 (N_1546,In_1350,In_1030);
nor U1547 (N_1547,In_544,In_125);
nand U1548 (N_1548,In_301,In_961);
nor U1549 (N_1549,In_79,In_1328);
nor U1550 (N_1550,In_763,In_1087);
nand U1551 (N_1551,In_1306,In_737);
xnor U1552 (N_1552,In_1084,In_103);
and U1553 (N_1553,In_941,In_10);
and U1554 (N_1554,In_630,In_189);
and U1555 (N_1555,In_839,In_1198);
or U1556 (N_1556,In_1046,In_1349);
xnor U1557 (N_1557,In_1485,In_1266);
and U1558 (N_1558,In_1227,In_549);
xnor U1559 (N_1559,In_810,In_371);
nand U1560 (N_1560,In_1277,In_42);
or U1561 (N_1561,In_1162,In_1340);
or U1562 (N_1562,In_1267,In_1394);
and U1563 (N_1563,In_1197,In_92);
and U1564 (N_1564,In_162,In_981);
and U1565 (N_1565,In_1151,In_550);
xnor U1566 (N_1566,In_258,In_885);
xnor U1567 (N_1567,In_730,In_412);
nand U1568 (N_1568,In_180,In_1405);
and U1569 (N_1569,In_695,In_836);
nand U1570 (N_1570,In_143,In_676);
nor U1571 (N_1571,In_2,In_712);
xor U1572 (N_1572,In_908,In_858);
or U1573 (N_1573,In_966,In_905);
xor U1574 (N_1574,In_694,In_202);
or U1575 (N_1575,In_1157,In_479);
and U1576 (N_1576,In_1350,In_780);
xnor U1577 (N_1577,In_781,In_563);
xnor U1578 (N_1578,In_352,In_48);
and U1579 (N_1579,In_662,In_1391);
nor U1580 (N_1580,In_497,In_129);
nor U1581 (N_1581,In_1058,In_1449);
nor U1582 (N_1582,In_1011,In_1212);
and U1583 (N_1583,In_311,In_1005);
xor U1584 (N_1584,In_1029,In_1384);
or U1585 (N_1585,In_982,In_105);
and U1586 (N_1586,In_1264,In_470);
or U1587 (N_1587,In_1380,In_396);
nor U1588 (N_1588,In_587,In_1173);
and U1589 (N_1589,In_1163,In_589);
nor U1590 (N_1590,In_1413,In_1018);
or U1591 (N_1591,In_640,In_105);
nor U1592 (N_1592,In_1302,In_1237);
xor U1593 (N_1593,In_207,In_746);
and U1594 (N_1594,In_329,In_94);
or U1595 (N_1595,In_934,In_29);
or U1596 (N_1596,In_780,In_127);
nor U1597 (N_1597,In_877,In_929);
and U1598 (N_1598,In_1385,In_133);
and U1599 (N_1599,In_721,In_237);
and U1600 (N_1600,In_30,In_572);
xor U1601 (N_1601,In_756,In_1267);
or U1602 (N_1602,In_417,In_119);
nor U1603 (N_1603,In_244,In_671);
or U1604 (N_1604,In_313,In_665);
nand U1605 (N_1605,In_792,In_743);
nor U1606 (N_1606,In_705,In_892);
nor U1607 (N_1607,In_479,In_611);
nor U1608 (N_1608,In_675,In_832);
nor U1609 (N_1609,In_978,In_313);
and U1610 (N_1610,In_947,In_692);
xnor U1611 (N_1611,In_1474,In_583);
nand U1612 (N_1612,In_424,In_989);
or U1613 (N_1613,In_663,In_1278);
or U1614 (N_1614,In_1223,In_1342);
nand U1615 (N_1615,In_1080,In_564);
or U1616 (N_1616,In_1467,In_1243);
nor U1617 (N_1617,In_1495,In_849);
xnor U1618 (N_1618,In_1495,In_1089);
nor U1619 (N_1619,In_1000,In_144);
xor U1620 (N_1620,In_163,In_1449);
or U1621 (N_1621,In_8,In_72);
or U1622 (N_1622,In_311,In_498);
nand U1623 (N_1623,In_203,In_370);
nand U1624 (N_1624,In_1332,In_1024);
or U1625 (N_1625,In_1188,In_494);
or U1626 (N_1626,In_125,In_669);
and U1627 (N_1627,In_628,In_716);
and U1628 (N_1628,In_598,In_715);
or U1629 (N_1629,In_1281,In_56);
or U1630 (N_1630,In_1464,In_1012);
nor U1631 (N_1631,In_1399,In_1427);
xnor U1632 (N_1632,In_1039,In_634);
nand U1633 (N_1633,In_494,In_1140);
xor U1634 (N_1634,In_1359,In_359);
and U1635 (N_1635,In_1143,In_407);
xor U1636 (N_1636,In_1332,In_108);
xnor U1637 (N_1637,In_603,In_1285);
xor U1638 (N_1638,In_183,In_1432);
xor U1639 (N_1639,In_399,In_1428);
xnor U1640 (N_1640,In_1,In_426);
nand U1641 (N_1641,In_1412,In_1494);
nand U1642 (N_1642,In_1499,In_1385);
nand U1643 (N_1643,In_1214,In_874);
nor U1644 (N_1644,In_112,In_1002);
or U1645 (N_1645,In_1142,In_1089);
or U1646 (N_1646,In_950,In_777);
and U1647 (N_1647,In_676,In_1492);
nand U1648 (N_1648,In_1192,In_769);
and U1649 (N_1649,In_434,In_1317);
xor U1650 (N_1650,In_542,In_853);
nor U1651 (N_1651,In_394,In_1305);
nand U1652 (N_1652,In_851,In_1170);
and U1653 (N_1653,In_384,In_1375);
nor U1654 (N_1654,In_1489,In_151);
nor U1655 (N_1655,In_1289,In_1196);
nand U1656 (N_1656,In_1408,In_271);
xnor U1657 (N_1657,In_128,In_1122);
xor U1658 (N_1658,In_271,In_1466);
nand U1659 (N_1659,In_241,In_1065);
nand U1660 (N_1660,In_980,In_1421);
and U1661 (N_1661,In_62,In_305);
and U1662 (N_1662,In_931,In_752);
xor U1663 (N_1663,In_775,In_1351);
and U1664 (N_1664,In_1194,In_792);
or U1665 (N_1665,In_23,In_540);
nand U1666 (N_1666,In_399,In_1449);
nand U1667 (N_1667,In_83,In_399);
nor U1668 (N_1668,In_24,In_528);
nor U1669 (N_1669,In_1222,In_1270);
xor U1670 (N_1670,In_448,In_786);
or U1671 (N_1671,In_1433,In_389);
and U1672 (N_1672,In_735,In_794);
or U1673 (N_1673,In_1418,In_784);
and U1674 (N_1674,In_1293,In_1384);
nor U1675 (N_1675,In_661,In_135);
nor U1676 (N_1676,In_699,In_234);
nand U1677 (N_1677,In_1306,In_1457);
xor U1678 (N_1678,In_886,In_1483);
nor U1679 (N_1679,In_700,In_1277);
and U1680 (N_1680,In_846,In_1138);
and U1681 (N_1681,In_82,In_178);
or U1682 (N_1682,In_534,In_612);
nand U1683 (N_1683,In_346,In_76);
or U1684 (N_1684,In_111,In_1053);
xor U1685 (N_1685,In_546,In_313);
or U1686 (N_1686,In_906,In_49);
nor U1687 (N_1687,In_1371,In_634);
nor U1688 (N_1688,In_542,In_1315);
and U1689 (N_1689,In_404,In_701);
nor U1690 (N_1690,In_1391,In_1175);
or U1691 (N_1691,In_787,In_688);
xor U1692 (N_1692,In_790,In_1116);
or U1693 (N_1693,In_271,In_1236);
nor U1694 (N_1694,In_818,In_1214);
xnor U1695 (N_1695,In_982,In_1450);
xor U1696 (N_1696,In_842,In_447);
or U1697 (N_1697,In_1420,In_151);
xor U1698 (N_1698,In_687,In_497);
and U1699 (N_1699,In_906,In_792);
xnor U1700 (N_1700,In_341,In_1369);
xnor U1701 (N_1701,In_1108,In_1314);
nor U1702 (N_1702,In_41,In_578);
nand U1703 (N_1703,In_238,In_751);
nand U1704 (N_1704,In_148,In_249);
and U1705 (N_1705,In_949,In_1201);
xor U1706 (N_1706,In_1191,In_971);
xor U1707 (N_1707,In_886,In_562);
nand U1708 (N_1708,In_1261,In_643);
nand U1709 (N_1709,In_652,In_1191);
nand U1710 (N_1710,In_1345,In_50);
or U1711 (N_1711,In_115,In_527);
xor U1712 (N_1712,In_101,In_416);
or U1713 (N_1713,In_1402,In_838);
nor U1714 (N_1714,In_243,In_864);
nor U1715 (N_1715,In_338,In_146);
or U1716 (N_1716,In_688,In_95);
and U1717 (N_1717,In_118,In_657);
and U1718 (N_1718,In_1215,In_961);
nor U1719 (N_1719,In_411,In_1130);
nand U1720 (N_1720,In_959,In_1460);
and U1721 (N_1721,In_1334,In_1125);
nand U1722 (N_1722,In_678,In_669);
xor U1723 (N_1723,In_1364,In_562);
xnor U1724 (N_1724,In_1223,In_162);
nand U1725 (N_1725,In_63,In_113);
nand U1726 (N_1726,In_902,In_710);
nor U1727 (N_1727,In_1276,In_390);
and U1728 (N_1728,In_426,In_814);
xor U1729 (N_1729,In_1159,In_1293);
nor U1730 (N_1730,In_179,In_871);
and U1731 (N_1731,In_371,In_113);
or U1732 (N_1732,In_163,In_581);
xnor U1733 (N_1733,In_1272,In_511);
and U1734 (N_1734,In_1323,In_1253);
xnor U1735 (N_1735,In_797,In_407);
or U1736 (N_1736,In_712,In_454);
and U1737 (N_1737,In_466,In_1365);
nor U1738 (N_1738,In_1275,In_309);
and U1739 (N_1739,In_1090,In_470);
xnor U1740 (N_1740,In_969,In_497);
nand U1741 (N_1741,In_489,In_385);
nand U1742 (N_1742,In_709,In_728);
xor U1743 (N_1743,In_252,In_157);
and U1744 (N_1744,In_543,In_1483);
nand U1745 (N_1745,In_1153,In_468);
or U1746 (N_1746,In_196,In_1345);
and U1747 (N_1747,In_1153,In_1158);
or U1748 (N_1748,In_666,In_89);
nand U1749 (N_1749,In_1440,In_1012);
nand U1750 (N_1750,In_1497,In_177);
or U1751 (N_1751,In_1479,In_15);
and U1752 (N_1752,In_1330,In_1327);
nor U1753 (N_1753,In_134,In_298);
and U1754 (N_1754,In_554,In_472);
nor U1755 (N_1755,In_65,In_1413);
xnor U1756 (N_1756,In_952,In_415);
nor U1757 (N_1757,In_671,In_239);
nand U1758 (N_1758,In_690,In_695);
nor U1759 (N_1759,In_496,In_1420);
and U1760 (N_1760,In_476,In_656);
nand U1761 (N_1761,In_1478,In_1019);
and U1762 (N_1762,In_657,In_745);
and U1763 (N_1763,In_1399,In_1321);
and U1764 (N_1764,In_10,In_471);
xnor U1765 (N_1765,In_4,In_1388);
nor U1766 (N_1766,In_401,In_985);
xnor U1767 (N_1767,In_487,In_861);
xor U1768 (N_1768,In_1488,In_751);
or U1769 (N_1769,In_1112,In_1284);
and U1770 (N_1770,In_1483,In_994);
and U1771 (N_1771,In_319,In_1332);
xor U1772 (N_1772,In_994,In_289);
or U1773 (N_1773,In_1065,In_225);
and U1774 (N_1774,In_106,In_328);
xnor U1775 (N_1775,In_778,In_1422);
nand U1776 (N_1776,In_314,In_937);
xor U1777 (N_1777,In_1279,In_1408);
nand U1778 (N_1778,In_161,In_919);
or U1779 (N_1779,In_614,In_408);
or U1780 (N_1780,In_1458,In_691);
and U1781 (N_1781,In_739,In_1332);
nand U1782 (N_1782,In_57,In_1216);
or U1783 (N_1783,In_402,In_780);
nand U1784 (N_1784,In_1359,In_536);
nand U1785 (N_1785,In_514,In_751);
nand U1786 (N_1786,In_249,In_163);
nand U1787 (N_1787,In_692,In_822);
and U1788 (N_1788,In_1137,In_596);
nor U1789 (N_1789,In_962,In_158);
nor U1790 (N_1790,In_1340,In_778);
nand U1791 (N_1791,In_374,In_158);
nand U1792 (N_1792,In_684,In_206);
or U1793 (N_1793,In_461,In_973);
nor U1794 (N_1794,In_549,In_1416);
nor U1795 (N_1795,In_1409,In_982);
nand U1796 (N_1796,In_130,In_1166);
nor U1797 (N_1797,In_1352,In_379);
and U1798 (N_1798,In_911,In_1182);
xnor U1799 (N_1799,In_1319,In_1497);
xor U1800 (N_1800,In_1482,In_1388);
nand U1801 (N_1801,In_1067,In_1391);
nand U1802 (N_1802,In_484,In_1324);
and U1803 (N_1803,In_953,In_1462);
nand U1804 (N_1804,In_903,In_519);
nor U1805 (N_1805,In_1298,In_669);
and U1806 (N_1806,In_1196,In_1005);
nand U1807 (N_1807,In_36,In_225);
xor U1808 (N_1808,In_405,In_1220);
nor U1809 (N_1809,In_1313,In_11);
nor U1810 (N_1810,In_1479,In_955);
nand U1811 (N_1811,In_1237,In_1214);
xor U1812 (N_1812,In_28,In_56);
xnor U1813 (N_1813,In_1328,In_690);
xnor U1814 (N_1814,In_777,In_874);
or U1815 (N_1815,In_919,In_810);
and U1816 (N_1816,In_1163,In_1415);
nand U1817 (N_1817,In_1363,In_266);
nor U1818 (N_1818,In_1411,In_596);
nor U1819 (N_1819,In_14,In_620);
and U1820 (N_1820,In_1037,In_1197);
or U1821 (N_1821,In_466,In_780);
nor U1822 (N_1822,In_295,In_83);
nand U1823 (N_1823,In_1210,In_208);
nor U1824 (N_1824,In_777,In_875);
or U1825 (N_1825,In_339,In_1453);
nand U1826 (N_1826,In_231,In_1343);
nand U1827 (N_1827,In_1370,In_156);
and U1828 (N_1828,In_863,In_68);
or U1829 (N_1829,In_838,In_817);
or U1830 (N_1830,In_897,In_14);
or U1831 (N_1831,In_401,In_611);
xnor U1832 (N_1832,In_1299,In_692);
nor U1833 (N_1833,In_515,In_48);
nor U1834 (N_1834,In_325,In_912);
and U1835 (N_1835,In_438,In_329);
nor U1836 (N_1836,In_1352,In_1409);
and U1837 (N_1837,In_52,In_608);
and U1838 (N_1838,In_1032,In_37);
nand U1839 (N_1839,In_1221,In_976);
xnor U1840 (N_1840,In_570,In_1481);
nand U1841 (N_1841,In_1089,In_1051);
xor U1842 (N_1842,In_796,In_375);
and U1843 (N_1843,In_180,In_395);
nand U1844 (N_1844,In_705,In_290);
or U1845 (N_1845,In_396,In_473);
xnor U1846 (N_1846,In_649,In_856);
and U1847 (N_1847,In_138,In_611);
xnor U1848 (N_1848,In_431,In_188);
nor U1849 (N_1849,In_16,In_272);
or U1850 (N_1850,In_1239,In_455);
and U1851 (N_1851,In_502,In_579);
xor U1852 (N_1852,In_247,In_1020);
nand U1853 (N_1853,In_109,In_812);
or U1854 (N_1854,In_759,In_290);
or U1855 (N_1855,In_346,In_562);
nand U1856 (N_1856,In_459,In_1024);
nand U1857 (N_1857,In_1142,In_590);
nand U1858 (N_1858,In_374,In_1202);
nand U1859 (N_1859,In_672,In_378);
or U1860 (N_1860,In_71,In_763);
nor U1861 (N_1861,In_824,In_442);
or U1862 (N_1862,In_863,In_502);
xnor U1863 (N_1863,In_1114,In_948);
nand U1864 (N_1864,In_1433,In_320);
xor U1865 (N_1865,In_697,In_852);
or U1866 (N_1866,In_680,In_181);
or U1867 (N_1867,In_1026,In_1013);
nand U1868 (N_1868,In_355,In_636);
xnor U1869 (N_1869,In_162,In_345);
nand U1870 (N_1870,In_1136,In_37);
or U1871 (N_1871,In_591,In_48);
xnor U1872 (N_1872,In_566,In_148);
nor U1873 (N_1873,In_494,In_970);
or U1874 (N_1874,In_433,In_1094);
nand U1875 (N_1875,In_292,In_233);
nand U1876 (N_1876,In_349,In_118);
nand U1877 (N_1877,In_1148,In_165);
nor U1878 (N_1878,In_759,In_1445);
nand U1879 (N_1879,In_197,In_1092);
xnor U1880 (N_1880,In_1294,In_1217);
nand U1881 (N_1881,In_364,In_989);
xor U1882 (N_1882,In_1000,In_517);
xnor U1883 (N_1883,In_376,In_1496);
and U1884 (N_1884,In_242,In_743);
nor U1885 (N_1885,In_198,In_984);
nand U1886 (N_1886,In_1161,In_1154);
nor U1887 (N_1887,In_1455,In_1405);
and U1888 (N_1888,In_758,In_1358);
nand U1889 (N_1889,In_960,In_988);
nand U1890 (N_1890,In_1306,In_537);
nor U1891 (N_1891,In_101,In_1090);
or U1892 (N_1892,In_51,In_993);
nor U1893 (N_1893,In_359,In_1078);
or U1894 (N_1894,In_152,In_1408);
xnor U1895 (N_1895,In_357,In_824);
and U1896 (N_1896,In_302,In_1288);
nand U1897 (N_1897,In_1054,In_76);
or U1898 (N_1898,In_312,In_902);
nor U1899 (N_1899,In_1381,In_1395);
nor U1900 (N_1900,In_744,In_1379);
nand U1901 (N_1901,In_1113,In_436);
xnor U1902 (N_1902,In_225,In_338);
nand U1903 (N_1903,In_532,In_969);
or U1904 (N_1904,In_298,In_282);
nor U1905 (N_1905,In_382,In_521);
xnor U1906 (N_1906,In_1496,In_424);
nor U1907 (N_1907,In_1102,In_1334);
xor U1908 (N_1908,In_614,In_870);
nor U1909 (N_1909,In_917,In_16);
or U1910 (N_1910,In_1450,In_769);
or U1911 (N_1911,In_769,In_1079);
nor U1912 (N_1912,In_313,In_741);
xnor U1913 (N_1913,In_1042,In_1234);
or U1914 (N_1914,In_570,In_774);
nor U1915 (N_1915,In_1018,In_565);
nor U1916 (N_1916,In_292,In_1140);
and U1917 (N_1917,In_994,In_881);
and U1918 (N_1918,In_335,In_227);
xnor U1919 (N_1919,In_541,In_62);
nor U1920 (N_1920,In_359,In_516);
nor U1921 (N_1921,In_875,In_1175);
or U1922 (N_1922,In_1273,In_15);
xnor U1923 (N_1923,In_127,In_1062);
and U1924 (N_1924,In_85,In_382);
nand U1925 (N_1925,In_1121,In_837);
or U1926 (N_1926,In_174,In_423);
nor U1927 (N_1927,In_1122,In_64);
or U1928 (N_1928,In_253,In_1196);
and U1929 (N_1929,In_1497,In_1353);
xnor U1930 (N_1930,In_308,In_505);
xnor U1931 (N_1931,In_170,In_1127);
and U1932 (N_1932,In_886,In_1042);
nor U1933 (N_1933,In_25,In_617);
xnor U1934 (N_1934,In_667,In_1179);
or U1935 (N_1935,In_1103,In_169);
xor U1936 (N_1936,In_188,In_603);
or U1937 (N_1937,In_769,In_572);
or U1938 (N_1938,In_1432,In_1431);
nor U1939 (N_1939,In_9,In_36);
xor U1940 (N_1940,In_1369,In_770);
xor U1941 (N_1941,In_1464,In_1362);
nand U1942 (N_1942,In_33,In_1117);
xnor U1943 (N_1943,In_412,In_1371);
and U1944 (N_1944,In_536,In_297);
and U1945 (N_1945,In_847,In_824);
nand U1946 (N_1946,In_1248,In_310);
xnor U1947 (N_1947,In_1217,In_667);
nor U1948 (N_1948,In_43,In_541);
xnor U1949 (N_1949,In_902,In_1486);
and U1950 (N_1950,In_1008,In_1146);
xor U1951 (N_1951,In_1297,In_613);
nor U1952 (N_1952,In_53,In_1335);
nor U1953 (N_1953,In_302,In_690);
xor U1954 (N_1954,In_158,In_1400);
nand U1955 (N_1955,In_1057,In_728);
and U1956 (N_1956,In_1167,In_362);
and U1957 (N_1957,In_695,In_1284);
or U1958 (N_1958,In_1376,In_55);
and U1959 (N_1959,In_325,In_800);
or U1960 (N_1960,In_490,In_398);
or U1961 (N_1961,In_650,In_501);
nor U1962 (N_1962,In_566,In_1361);
and U1963 (N_1963,In_291,In_1257);
nand U1964 (N_1964,In_986,In_814);
nor U1965 (N_1965,In_1291,In_1009);
nand U1966 (N_1966,In_486,In_1448);
or U1967 (N_1967,In_122,In_373);
or U1968 (N_1968,In_1267,In_1372);
or U1969 (N_1969,In_119,In_1273);
and U1970 (N_1970,In_954,In_198);
or U1971 (N_1971,In_1201,In_1135);
nand U1972 (N_1972,In_1041,In_1105);
nor U1973 (N_1973,In_582,In_634);
nor U1974 (N_1974,In_932,In_1090);
nor U1975 (N_1975,In_308,In_1347);
nand U1976 (N_1976,In_10,In_1085);
and U1977 (N_1977,In_1006,In_96);
and U1978 (N_1978,In_1301,In_1438);
and U1979 (N_1979,In_159,In_1428);
nand U1980 (N_1980,In_33,In_1452);
nor U1981 (N_1981,In_1254,In_945);
and U1982 (N_1982,In_984,In_1236);
and U1983 (N_1983,In_1402,In_251);
and U1984 (N_1984,In_605,In_44);
nor U1985 (N_1985,In_612,In_1026);
and U1986 (N_1986,In_363,In_786);
and U1987 (N_1987,In_1023,In_58);
or U1988 (N_1988,In_1300,In_1365);
nand U1989 (N_1989,In_1149,In_711);
nor U1990 (N_1990,In_733,In_491);
xor U1991 (N_1991,In_1076,In_196);
or U1992 (N_1992,In_1094,In_581);
or U1993 (N_1993,In_1315,In_63);
nand U1994 (N_1994,In_599,In_195);
nand U1995 (N_1995,In_338,In_783);
nor U1996 (N_1996,In_646,In_240);
nor U1997 (N_1997,In_1322,In_649);
xnor U1998 (N_1998,In_1211,In_831);
and U1999 (N_1999,In_1013,In_1498);
and U2000 (N_2000,In_993,In_1302);
nor U2001 (N_2001,In_1173,In_1297);
nand U2002 (N_2002,In_1093,In_896);
xnor U2003 (N_2003,In_1099,In_1039);
nand U2004 (N_2004,In_1191,In_465);
and U2005 (N_2005,In_1014,In_654);
nand U2006 (N_2006,In_618,In_1474);
and U2007 (N_2007,In_991,In_706);
nor U2008 (N_2008,In_366,In_884);
xnor U2009 (N_2009,In_624,In_387);
nand U2010 (N_2010,In_353,In_941);
nor U2011 (N_2011,In_560,In_21);
or U2012 (N_2012,In_168,In_213);
and U2013 (N_2013,In_399,In_689);
xnor U2014 (N_2014,In_627,In_1167);
xor U2015 (N_2015,In_1351,In_33);
and U2016 (N_2016,In_1283,In_1002);
nand U2017 (N_2017,In_1437,In_351);
nand U2018 (N_2018,In_1242,In_1304);
or U2019 (N_2019,In_411,In_698);
or U2020 (N_2020,In_190,In_294);
nand U2021 (N_2021,In_909,In_837);
nand U2022 (N_2022,In_1422,In_888);
nand U2023 (N_2023,In_583,In_436);
and U2024 (N_2024,In_722,In_1323);
nand U2025 (N_2025,In_1192,In_1249);
nand U2026 (N_2026,In_371,In_328);
nand U2027 (N_2027,In_70,In_1223);
nor U2028 (N_2028,In_77,In_394);
nand U2029 (N_2029,In_493,In_247);
nor U2030 (N_2030,In_290,In_1171);
and U2031 (N_2031,In_15,In_240);
nor U2032 (N_2032,In_671,In_1400);
nor U2033 (N_2033,In_635,In_308);
xor U2034 (N_2034,In_947,In_37);
or U2035 (N_2035,In_114,In_1377);
nor U2036 (N_2036,In_1237,In_1439);
and U2037 (N_2037,In_1179,In_545);
nand U2038 (N_2038,In_535,In_1344);
nand U2039 (N_2039,In_1078,In_1026);
and U2040 (N_2040,In_241,In_1292);
xnor U2041 (N_2041,In_424,In_863);
xnor U2042 (N_2042,In_1383,In_996);
nor U2043 (N_2043,In_355,In_675);
nand U2044 (N_2044,In_884,In_640);
nand U2045 (N_2045,In_1180,In_1457);
and U2046 (N_2046,In_319,In_645);
nand U2047 (N_2047,In_1290,In_323);
and U2048 (N_2048,In_1250,In_154);
or U2049 (N_2049,In_1022,In_228);
xor U2050 (N_2050,In_971,In_1115);
and U2051 (N_2051,In_493,In_113);
and U2052 (N_2052,In_867,In_868);
nor U2053 (N_2053,In_1455,In_570);
and U2054 (N_2054,In_959,In_203);
or U2055 (N_2055,In_397,In_827);
nor U2056 (N_2056,In_415,In_695);
xor U2057 (N_2057,In_340,In_1458);
xor U2058 (N_2058,In_1304,In_1394);
nor U2059 (N_2059,In_1393,In_1370);
xor U2060 (N_2060,In_1493,In_268);
nor U2061 (N_2061,In_186,In_1174);
nand U2062 (N_2062,In_1181,In_1174);
nand U2063 (N_2063,In_311,In_1069);
and U2064 (N_2064,In_1273,In_675);
or U2065 (N_2065,In_161,In_1196);
and U2066 (N_2066,In_619,In_584);
xor U2067 (N_2067,In_886,In_1109);
and U2068 (N_2068,In_956,In_1404);
xnor U2069 (N_2069,In_70,In_488);
or U2070 (N_2070,In_1261,In_252);
nand U2071 (N_2071,In_1201,In_1104);
or U2072 (N_2072,In_295,In_633);
nand U2073 (N_2073,In_1039,In_317);
nor U2074 (N_2074,In_605,In_267);
nand U2075 (N_2075,In_331,In_1262);
nor U2076 (N_2076,In_1334,In_300);
and U2077 (N_2077,In_136,In_1239);
nor U2078 (N_2078,In_459,In_461);
nand U2079 (N_2079,In_1261,In_45);
or U2080 (N_2080,In_161,In_393);
nor U2081 (N_2081,In_825,In_357);
or U2082 (N_2082,In_1068,In_163);
or U2083 (N_2083,In_1284,In_1255);
or U2084 (N_2084,In_547,In_660);
or U2085 (N_2085,In_406,In_1372);
and U2086 (N_2086,In_97,In_1015);
xor U2087 (N_2087,In_1408,In_373);
xor U2088 (N_2088,In_666,In_196);
xor U2089 (N_2089,In_846,In_247);
nand U2090 (N_2090,In_326,In_444);
nand U2091 (N_2091,In_412,In_945);
xnor U2092 (N_2092,In_464,In_630);
or U2093 (N_2093,In_1428,In_1061);
nor U2094 (N_2094,In_1439,In_525);
or U2095 (N_2095,In_967,In_1186);
xnor U2096 (N_2096,In_371,In_623);
and U2097 (N_2097,In_240,In_1481);
nor U2098 (N_2098,In_832,In_1359);
nand U2099 (N_2099,In_653,In_639);
nor U2100 (N_2100,In_1353,In_210);
or U2101 (N_2101,In_412,In_1207);
nand U2102 (N_2102,In_878,In_322);
xor U2103 (N_2103,In_1200,In_903);
nor U2104 (N_2104,In_1349,In_410);
xnor U2105 (N_2105,In_442,In_78);
nand U2106 (N_2106,In_1147,In_1458);
xor U2107 (N_2107,In_908,In_427);
nor U2108 (N_2108,In_17,In_1082);
nand U2109 (N_2109,In_135,In_917);
nand U2110 (N_2110,In_871,In_463);
nor U2111 (N_2111,In_1002,In_873);
or U2112 (N_2112,In_324,In_1450);
nand U2113 (N_2113,In_584,In_829);
and U2114 (N_2114,In_915,In_51);
xnor U2115 (N_2115,In_315,In_411);
nand U2116 (N_2116,In_735,In_1040);
or U2117 (N_2117,In_848,In_557);
nand U2118 (N_2118,In_318,In_1065);
or U2119 (N_2119,In_163,In_239);
nor U2120 (N_2120,In_678,In_1328);
nand U2121 (N_2121,In_688,In_1095);
xnor U2122 (N_2122,In_432,In_960);
or U2123 (N_2123,In_362,In_253);
nand U2124 (N_2124,In_1145,In_873);
and U2125 (N_2125,In_810,In_893);
nand U2126 (N_2126,In_850,In_514);
nand U2127 (N_2127,In_49,In_384);
and U2128 (N_2128,In_963,In_287);
xor U2129 (N_2129,In_1427,In_1296);
nand U2130 (N_2130,In_419,In_639);
and U2131 (N_2131,In_608,In_285);
xor U2132 (N_2132,In_1390,In_61);
and U2133 (N_2133,In_11,In_458);
xnor U2134 (N_2134,In_133,In_875);
or U2135 (N_2135,In_1297,In_612);
or U2136 (N_2136,In_43,In_967);
and U2137 (N_2137,In_454,In_1159);
xor U2138 (N_2138,In_112,In_1077);
or U2139 (N_2139,In_408,In_613);
nand U2140 (N_2140,In_1016,In_434);
nand U2141 (N_2141,In_180,In_847);
nand U2142 (N_2142,In_1189,In_1236);
or U2143 (N_2143,In_195,In_60);
and U2144 (N_2144,In_381,In_823);
or U2145 (N_2145,In_163,In_445);
and U2146 (N_2146,In_541,In_745);
or U2147 (N_2147,In_1044,In_1158);
or U2148 (N_2148,In_1350,In_48);
nand U2149 (N_2149,In_319,In_1089);
xor U2150 (N_2150,In_197,In_786);
and U2151 (N_2151,In_1440,In_315);
or U2152 (N_2152,In_602,In_902);
or U2153 (N_2153,In_256,In_583);
nand U2154 (N_2154,In_323,In_1360);
or U2155 (N_2155,In_469,In_1468);
nor U2156 (N_2156,In_1467,In_1140);
nor U2157 (N_2157,In_1462,In_1355);
xor U2158 (N_2158,In_817,In_1154);
xor U2159 (N_2159,In_463,In_480);
or U2160 (N_2160,In_1170,In_102);
xnor U2161 (N_2161,In_1070,In_269);
and U2162 (N_2162,In_184,In_21);
and U2163 (N_2163,In_88,In_251);
and U2164 (N_2164,In_326,In_806);
xor U2165 (N_2165,In_1100,In_1460);
nand U2166 (N_2166,In_1267,In_515);
nand U2167 (N_2167,In_1207,In_853);
and U2168 (N_2168,In_1343,In_702);
nor U2169 (N_2169,In_1329,In_1327);
or U2170 (N_2170,In_110,In_802);
xor U2171 (N_2171,In_498,In_660);
nor U2172 (N_2172,In_600,In_326);
nor U2173 (N_2173,In_1139,In_588);
xnor U2174 (N_2174,In_1114,In_778);
nor U2175 (N_2175,In_1258,In_1006);
nand U2176 (N_2176,In_51,In_1198);
and U2177 (N_2177,In_963,In_497);
or U2178 (N_2178,In_113,In_746);
or U2179 (N_2179,In_857,In_599);
nand U2180 (N_2180,In_1134,In_1186);
nor U2181 (N_2181,In_287,In_1361);
or U2182 (N_2182,In_369,In_968);
nor U2183 (N_2183,In_770,In_1067);
xor U2184 (N_2184,In_746,In_698);
and U2185 (N_2185,In_266,In_1280);
xnor U2186 (N_2186,In_1308,In_181);
or U2187 (N_2187,In_884,In_1166);
or U2188 (N_2188,In_216,In_872);
xor U2189 (N_2189,In_279,In_484);
nor U2190 (N_2190,In_775,In_393);
nor U2191 (N_2191,In_267,In_1086);
nor U2192 (N_2192,In_642,In_1311);
and U2193 (N_2193,In_1039,In_1044);
xor U2194 (N_2194,In_1003,In_160);
nor U2195 (N_2195,In_1125,In_73);
xnor U2196 (N_2196,In_1329,In_401);
nand U2197 (N_2197,In_1000,In_379);
or U2198 (N_2198,In_1216,In_503);
and U2199 (N_2199,In_1492,In_317);
or U2200 (N_2200,In_913,In_1221);
nor U2201 (N_2201,In_919,In_85);
and U2202 (N_2202,In_798,In_993);
or U2203 (N_2203,In_776,In_579);
xnor U2204 (N_2204,In_506,In_1188);
or U2205 (N_2205,In_624,In_1404);
nor U2206 (N_2206,In_521,In_510);
nand U2207 (N_2207,In_452,In_1426);
nand U2208 (N_2208,In_729,In_1016);
nand U2209 (N_2209,In_647,In_696);
nand U2210 (N_2210,In_1117,In_549);
nand U2211 (N_2211,In_9,In_63);
nor U2212 (N_2212,In_345,In_1288);
nor U2213 (N_2213,In_930,In_143);
xnor U2214 (N_2214,In_1423,In_378);
nor U2215 (N_2215,In_433,In_1181);
xnor U2216 (N_2216,In_868,In_376);
and U2217 (N_2217,In_571,In_717);
xnor U2218 (N_2218,In_686,In_257);
and U2219 (N_2219,In_988,In_1012);
or U2220 (N_2220,In_128,In_576);
nor U2221 (N_2221,In_1496,In_601);
and U2222 (N_2222,In_819,In_966);
nand U2223 (N_2223,In_285,In_73);
nand U2224 (N_2224,In_1023,In_1275);
nor U2225 (N_2225,In_1238,In_1038);
and U2226 (N_2226,In_919,In_993);
or U2227 (N_2227,In_137,In_158);
nor U2228 (N_2228,In_251,In_990);
xor U2229 (N_2229,In_599,In_366);
xor U2230 (N_2230,In_247,In_1243);
nor U2231 (N_2231,In_546,In_1127);
and U2232 (N_2232,In_1262,In_1358);
nor U2233 (N_2233,In_510,In_989);
xnor U2234 (N_2234,In_566,In_722);
xnor U2235 (N_2235,In_852,In_441);
nor U2236 (N_2236,In_275,In_634);
nand U2237 (N_2237,In_1290,In_988);
or U2238 (N_2238,In_1359,In_685);
nand U2239 (N_2239,In_284,In_842);
xor U2240 (N_2240,In_1407,In_34);
and U2241 (N_2241,In_734,In_400);
nand U2242 (N_2242,In_249,In_362);
or U2243 (N_2243,In_893,In_364);
or U2244 (N_2244,In_254,In_613);
or U2245 (N_2245,In_854,In_798);
nor U2246 (N_2246,In_1250,In_722);
and U2247 (N_2247,In_600,In_101);
nor U2248 (N_2248,In_1365,In_799);
nor U2249 (N_2249,In_647,In_667);
or U2250 (N_2250,In_135,In_379);
xor U2251 (N_2251,In_703,In_993);
or U2252 (N_2252,In_408,In_1181);
nor U2253 (N_2253,In_204,In_1009);
nor U2254 (N_2254,In_706,In_11);
nor U2255 (N_2255,In_743,In_111);
nor U2256 (N_2256,In_96,In_602);
xnor U2257 (N_2257,In_1125,In_1059);
or U2258 (N_2258,In_1080,In_285);
xor U2259 (N_2259,In_1024,In_26);
and U2260 (N_2260,In_436,In_423);
and U2261 (N_2261,In_222,In_201);
nand U2262 (N_2262,In_815,In_837);
xor U2263 (N_2263,In_436,In_295);
nor U2264 (N_2264,In_755,In_421);
nand U2265 (N_2265,In_731,In_1288);
nand U2266 (N_2266,In_520,In_938);
and U2267 (N_2267,In_653,In_535);
nand U2268 (N_2268,In_1441,In_1407);
nand U2269 (N_2269,In_976,In_476);
and U2270 (N_2270,In_1004,In_1328);
or U2271 (N_2271,In_869,In_284);
nor U2272 (N_2272,In_450,In_760);
xor U2273 (N_2273,In_656,In_1490);
or U2274 (N_2274,In_800,In_9);
xnor U2275 (N_2275,In_1236,In_1204);
and U2276 (N_2276,In_472,In_1242);
and U2277 (N_2277,In_745,In_194);
or U2278 (N_2278,In_226,In_568);
or U2279 (N_2279,In_682,In_1005);
and U2280 (N_2280,In_631,In_1145);
nor U2281 (N_2281,In_1206,In_855);
nor U2282 (N_2282,In_40,In_970);
xnor U2283 (N_2283,In_18,In_1066);
or U2284 (N_2284,In_732,In_858);
or U2285 (N_2285,In_1406,In_61);
nor U2286 (N_2286,In_348,In_1142);
xnor U2287 (N_2287,In_1444,In_597);
nand U2288 (N_2288,In_251,In_867);
xor U2289 (N_2289,In_683,In_1258);
and U2290 (N_2290,In_930,In_689);
and U2291 (N_2291,In_987,In_1289);
nand U2292 (N_2292,In_1274,In_168);
xor U2293 (N_2293,In_544,In_364);
xnor U2294 (N_2294,In_1186,In_687);
and U2295 (N_2295,In_286,In_198);
nor U2296 (N_2296,In_655,In_560);
or U2297 (N_2297,In_1129,In_765);
and U2298 (N_2298,In_677,In_728);
nand U2299 (N_2299,In_1164,In_1067);
xnor U2300 (N_2300,In_885,In_144);
nor U2301 (N_2301,In_1102,In_451);
nor U2302 (N_2302,In_928,In_312);
or U2303 (N_2303,In_673,In_361);
xnor U2304 (N_2304,In_629,In_46);
and U2305 (N_2305,In_644,In_147);
and U2306 (N_2306,In_746,In_714);
or U2307 (N_2307,In_721,In_701);
nand U2308 (N_2308,In_851,In_1136);
or U2309 (N_2309,In_1389,In_1009);
or U2310 (N_2310,In_1332,In_559);
nor U2311 (N_2311,In_1081,In_1141);
and U2312 (N_2312,In_476,In_1342);
nand U2313 (N_2313,In_63,In_315);
or U2314 (N_2314,In_445,In_567);
nand U2315 (N_2315,In_115,In_670);
xor U2316 (N_2316,In_170,In_251);
nor U2317 (N_2317,In_94,In_370);
nor U2318 (N_2318,In_554,In_549);
xor U2319 (N_2319,In_1244,In_728);
or U2320 (N_2320,In_439,In_726);
xor U2321 (N_2321,In_670,In_13);
xor U2322 (N_2322,In_542,In_1108);
nand U2323 (N_2323,In_96,In_1264);
or U2324 (N_2324,In_1354,In_1051);
xnor U2325 (N_2325,In_1032,In_1043);
and U2326 (N_2326,In_1444,In_1248);
nor U2327 (N_2327,In_1141,In_541);
or U2328 (N_2328,In_1388,In_453);
or U2329 (N_2329,In_554,In_157);
and U2330 (N_2330,In_5,In_1253);
xor U2331 (N_2331,In_689,In_43);
nand U2332 (N_2332,In_1345,In_778);
nor U2333 (N_2333,In_1331,In_798);
nand U2334 (N_2334,In_302,In_733);
xor U2335 (N_2335,In_993,In_670);
xor U2336 (N_2336,In_792,In_870);
nor U2337 (N_2337,In_720,In_469);
nand U2338 (N_2338,In_85,In_321);
nand U2339 (N_2339,In_615,In_202);
or U2340 (N_2340,In_1417,In_494);
nor U2341 (N_2341,In_110,In_715);
and U2342 (N_2342,In_196,In_520);
xnor U2343 (N_2343,In_150,In_1435);
xnor U2344 (N_2344,In_728,In_770);
and U2345 (N_2345,In_1393,In_1499);
nor U2346 (N_2346,In_507,In_1179);
or U2347 (N_2347,In_41,In_180);
xnor U2348 (N_2348,In_910,In_352);
xor U2349 (N_2349,In_1244,In_973);
or U2350 (N_2350,In_1344,In_635);
or U2351 (N_2351,In_1145,In_922);
or U2352 (N_2352,In_641,In_68);
nor U2353 (N_2353,In_1358,In_446);
or U2354 (N_2354,In_382,In_464);
and U2355 (N_2355,In_1019,In_1080);
or U2356 (N_2356,In_882,In_845);
xnor U2357 (N_2357,In_1402,In_1033);
or U2358 (N_2358,In_1072,In_242);
and U2359 (N_2359,In_1199,In_1271);
or U2360 (N_2360,In_433,In_451);
and U2361 (N_2361,In_1234,In_1087);
nor U2362 (N_2362,In_1118,In_1153);
nand U2363 (N_2363,In_1499,In_1215);
or U2364 (N_2364,In_1283,In_974);
nor U2365 (N_2365,In_1402,In_1334);
nand U2366 (N_2366,In_265,In_501);
nor U2367 (N_2367,In_942,In_383);
and U2368 (N_2368,In_875,In_620);
nor U2369 (N_2369,In_679,In_93);
and U2370 (N_2370,In_395,In_449);
nor U2371 (N_2371,In_498,In_383);
or U2372 (N_2372,In_785,In_368);
or U2373 (N_2373,In_1202,In_803);
or U2374 (N_2374,In_409,In_1392);
or U2375 (N_2375,In_414,In_594);
xnor U2376 (N_2376,In_309,In_1032);
nor U2377 (N_2377,In_457,In_872);
and U2378 (N_2378,In_980,In_402);
or U2379 (N_2379,In_965,In_970);
or U2380 (N_2380,In_114,In_535);
or U2381 (N_2381,In_261,In_1240);
nand U2382 (N_2382,In_702,In_453);
nand U2383 (N_2383,In_1216,In_436);
nor U2384 (N_2384,In_2,In_958);
xor U2385 (N_2385,In_789,In_189);
nor U2386 (N_2386,In_1309,In_1223);
nor U2387 (N_2387,In_69,In_1000);
xor U2388 (N_2388,In_946,In_888);
nor U2389 (N_2389,In_957,In_403);
and U2390 (N_2390,In_1486,In_1002);
and U2391 (N_2391,In_1454,In_456);
or U2392 (N_2392,In_411,In_43);
xor U2393 (N_2393,In_910,In_399);
or U2394 (N_2394,In_629,In_317);
nand U2395 (N_2395,In_362,In_942);
nor U2396 (N_2396,In_760,In_36);
and U2397 (N_2397,In_985,In_726);
xor U2398 (N_2398,In_1290,In_258);
or U2399 (N_2399,In_1305,In_474);
or U2400 (N_2400,In_252,In_992);
xnor U2401 (N_2401,In_384,In_519);
nor U2402 (N_2402,In_1338,In_1204);
nand U2403 (N_2403,In_815,In_931);
nor U2404 (N_2404,In_1066,In_1167);
nor U2405 (N_2405,In_1410,In_308);
or U2406 (N_2406,In_1270,In_343);
and U2407 (N_2407,In_362,In_929);
xor U2408 (N_2408,In_502,In_643);
nor U2409 (N_2409,In_1050,In_1163);
nand U2410 (N_2410,In_386,In_93);
nor U2411 (N_2411,In_905,In_1193);
or U2412 (N_2412,In_1425,In_1043);
xor U2413 (N_2413,In_1414,In_1013);
and U2414 (N_2414,In_1344,In_307);
nand U2415 (N_2415,In_1335,In_1478);
nand U2416 (N_2416,In_1056,In_1088);
or U2417 (N_2417,In_1117,In_1011);
nand U2418 (N_2418,In_444,In_895);
nand U2419 (N_2419,In_256,In_1234);
or U2420 (N_2420,In_912,In_1081);
or U2421 (N_2421,In_566,In_384);
xnor U2422 (N_2422,In_958,In_545);
and U2423 (N_2423,In_824,In_1076);
nor U2424 (N_2424,In_1210,In_1457);
and U2425 (N_2425,In_1382,In_1039);
xnor U2426 (N_2426,In_414,In_761);
nor U2427 (N_2427,In_660,In_761);
nand U2428 (N_2428,In_844,In_851);
or U2429 (N_2429,In_234,In_1484);
nor U2430 (N_2430,In_968,In_1252);
nor U2431 (N_2431,In_1115,In_425);
nand U2432 (N_2432,In_1165,In_822);
and U2433 (N_2433,In_1182,In_585);
xnor U2434 (N_2434,In_696,In_1193);
and U2435 (N_2435,In_623,In_564);
xnor U2436 (N_2436,In_99,In_719);
nand U2437 (N_2437,In_180,In_19);
and U2438 (N_2438,In_890,In_206);
and U2439 (N_2439,In_1387,In_35);
and U2440 (N_2440,In_555,In_635);
nand U2441 (N_2441,In_608,In_778);
or U2442 (N_2442,In_1108,In_878);
nand U2443 (N_2443,In_354,In_952);
nor U2444 (N_2444,In_774,In_447);
nand U2445 (N_2445,In_888,In_1364);
or U2446 (N_2446,In_1334,In_1321);
nand U2447 (N_2447,In_1197,In_199);
xnor U2448 (N_2448,In_1443,In_287);
nor U2449 (N_2449,In_1259,In_562);
nand U2450 (N_2450,In_664,In_902);
or U2451 (N_2451,In_763,In_1133);
and U2452 (N_2452,In_1071,In_559);
nand U2453 (N_2453,In_137,In_369);
nand U2454 (N_2454,In_1273,In_783);
nor U2455 (N_2455,In_147,In_805);
xor U2456 (N_2456,In_226,In_706);
and U2457 (N_2457,In_499,In_1219);
xnor U2458 (N_2458,In_355,In_186);
xor U2459 (N_2459,In_438,In_1128);
or U2460 (N_2460,In_592,In_465);
and U2461 (N_2461,In_1158,In_632);
xor U2462 (N_2462,In_104,In_1498);
nor U2463 (N_2463,In_57,In_466);
or U2464 (N_2464,In_824,In_1221);
nor U2465 (N_2465,In_647,In_220);
or U2466 (N_2466,In_758,In_701);
xor U2467 (N_2467,In_14,In_759);
or U2468 (N_2468,In_1324,In_816);
or U2469 (N_2469,In_83,In_6);
nor U2470 (N_2470,In_148,In_989);
and U2471 (N_2471,In_502,In_441);
nand U2472 (N_2472,In_240,In_153);
and U2473 (N_2473,In_860,In_1155);
nor U2474 (N_2474,In_407,In_387);
nor U2475 (N_2475,In_641,In_1287);
xor U2476 (N_2476,In_1257,In_1445);
nor U2477 (N_2477,In_60,In_1276);
and U2478 (N_2478,In_1302,In_899);
nand U2479 (N_2479,In_360,In_821);
xnor U2480 (N_2480,In_1327,In_299);
nor U2481 (N_2481,In_356,In_1267);
nor U2482 (N_2482,In_1356,In_659);
or U2483 (N_2483,In_440,In_1433);
nand U2484 (N_2484,In_1199,In_893);
or U2485 (N_2485,In_676,In_475);
or U2486 (N_2486,In_1403,In_1434);
nor U2487 (N_2487,In_1161,In_620);
nand U2488 (N_2488,In_99,In_531);
or U2489 (N_2489,In_1045,In_909);
xnor U2490 (N_2490,In_1135,In_1217);
nor U2491 (N_2491,In_831,In_37);
and U2492 (N_2492,In_1060,In_222);
and U2493 (N_2493,In_548,In_1471);
nor U2494 (N_2494,In_55,In_638);
or U2495 (N_2495,In_207,In_973);
and U2496 (N_2496,In_1057,In_1200);
or U2497 (N_2497,In_1213,In_4);
or U2498 (N_2498,In_1366,In_741);
nor U2499 (N_2499,In_857,In_1367);
and U2500 (N_2500,In_224,In_1109);
nor U2501 (N_2501,In_1168,In_760);
and U2502 (N_2502,In_1468,In_1464);
nor U2503 (N_2503,In_777,In_851);
nand U2504 (N_2504,In_916,In_604);
and U2505 (N_2505,In_1244,In_1285);
and U2506 (N_2506,In_1122,In_547);
nand U2507 (N_2507,In_701,In_267);
and U2508 (N_2508,In_412,In_1341);
or U2509 (N_2509,In_1443,In_817);
nand U2510 (N_2510,In_962,In_1222);
nor U2511 (N_2511,In_1221,In_735);
and U2512 (N_2512,In_1111,In_8);
nor U2513 (N_2513,In_689,In_1081);
and U2514 (N_2514,In_618,In_334);
xnor U2515 (N_2515,In_250,In_612);
or U2516 (N_2516,In_986,In_854);
nand U2517 (N_2517,In_666,In_440);
xor U2518 (N_2518,In_312,In_1088);
nor U2519 (N_2519,In_415,In_60);
nand U2520 (N_2520,In_451,In_1000);
or U2521 (N_2521,In_906,In_34);
nand U2522 (N_2522,In_1038,In_1237);
and U2523 (N_2523,In_394,In_109);
and U2524 (N_2524,In_1157,In_980);
or U2525 (N_2525,In_330,In_24);
nand U2526 (N_2526,In_89,In_759);
or U2527 (N_2527,In_1310,In_1222);
xnor U2528 (N_2528,In_39,In_782);
or U2529 (N_2529,In_691,In_1258);
xor U2530 (N_2530,In_791,In_688);
nand U2531 (N_2531,In_233,In_418);
or U2532 (N_2532,In_577,In_1100);
and U2533 (N_2533,In_811,In_953);
and U2534 (N_2534,In_1107,In_1284);
or U2535 (N_2535,In_363,In_1446);
and U2536 (N_2536,In_623,In_502);
or U2537 (N_2537,In_410,In_1316);
xnor U2538 (N_2538,In_1017,In_253);
or U2539 (N_2539,In_1054,In_501);
and U2540 (N_2540,In_345,In_130);
xnor U2541 (N_2541,In_839,In_398);
nand U2542 (N_2542,In_1477,In_836);
and U2543 (N_2543,In_1002,In_1459);
and U2544 (N_2544,In_2,In_1059);
nand U2545 (N_2545,In_578,In_441);
nand U2546 (N_2546,In_648,In_607);
or U2547 (N_2547,In_127,In_1267);
and U2548 (N_2548,In_205,In_935);
xnor U2549 (N_2549,In_589,In_137);
or U2550 (N_2550,In_1393,In_772);
or U2551 (N_2551,In_1105,In_931);
nand U2552 (N_2552,In_945,In_360);
nor U2553 (N_2553,In_541,In_1445);
or U2554 (N_2554,In_520,In_1220);
nor U2555 (N_2555,In_1247,In_942);
nor U2556 (N_2556,In_1251,In_1408);
xnor U2557 (N_2557,In_1134,In_606);
nand U2558 (N_2558,In_510,In_54);
or U2559 (N_2559,In_288,In_1073);
nand U2560 (N_2560,In_331,In_1184);
nor U2561 (N_2561,In_869,In_1023);
nand U2562 (N_2562,In_1459,In_1466);
nor U2563 (N_2563,In_851,In_1000);
xor U2564 (N_2564,In_1332,In_417);
nor U2565 (N_2565,In_1111,In_966);
nor U2566 (N_2566,In_200,In_1108);
nand U2567 (N_2567,In_266,In_1357);
and U2568 (N_2568,In_310,In_1269);
nor U2569 (N_2569,In_1337,In_564);
nor U2570 (N_2570,In_1302,In_1296);
or U2571 (N_2571,In_349,In_822);
nand U2572 (N_2572,In_278,In_919);
xor U2573 (N_2573,In_341,In_582);
or U2574 (N_2574,In_1358,In_1421);
xnor U2575 (N_2575,In_1379,In_506);
xor U2576 (N_2576,In_886,In_721);
and U2577 (N_2577,In_872,In_671);
nand U2578 (N_2578,In_188,In_1424);
and U2579 (N_2579,In_315,In_952);
nor U2580 (N_2580,In_1142,In_93);
nor U2581 (N_2581,In_405,In_684);
nor U2582 (N_2582,In_757,In_1112);
xnor U2583 (N_2583,In_1362,In_1118);
or U2584 (N_2584,In_0,In_179);
or U2585 (N_2585,In_1113,In_631);
xnor U2586 (N_2586,In_1100,In_1428);
or U2587 (N_2587,In_1011,In_128);
and U2588 (N_2588,In_1191,In_1397);
nor U2589 (N_2589,In_563,In_1169);
or U2590 (N_2590,In_299,In_343);
and U2591 (N_2591,In_26,In_320);
nor U2592 (N_2592,In_815,In_952);
nand U2593 (N_2593,In_860,In_776);
and U2594 (N_2594,In_1446,In_1227);
nor U2595 (N_2595,In_609,In_1400);
nand U2596 (N_2596,In_1055,In_915);
nor U2597 (N_2597,In_760,In_1106);
nand U2598 (N_2598,In_1116,In_552);
nand U2599 (N_2599,In_266,In_380);
and U2600 (N_2600,In_780,In_1130);
nand U2601 (N_2601,In_360,In_1246);
nor U2602 (N_2602,In_386,In_367);
and U2603 (N_2603,In_67,In_443);
and U2604 (N_2604,In_267,In_388);
and U2605 (N_2605,In_1003,In_1017);
nand U2606 (N_2606,In_797,In_1098);
xnor U2607 (N_2607,In_746,In_125);
or U2608 (N_2608,In_576,In_634);
nand U2609 (N_2609,In_1408,In_1249);
nor U2610 (N_2610,In_1174,In_850);
nand U2611 (N_2611,In_717,In_1282);
or U2612 (N_2612,In_412,In_1073);
or U2613 (N_2613,In_579,In_1348);
and U2614 (N_2614,In_728,In_278);
nor U2615 (N_2615,In_227,In_1373);
and U2616 (N_2616,In_867,In_6);
and U2617 (N_2617,In_675,In_723);
nand U2618 (N_2618,In_493,In_1334);
nand U2619 (N_2619,In_803,In_1225);
nand U2620 (N_2620,In_1314,In_710);
xor U2621 (N_2621,In_7,In_294);
or U2622 (N_2622,In_1359,In_534);
xnor U2623 (N_2623,In_1472,In_47);
xnor U2624 (N_2624,In_1454,In_978);
xor U2625 (N_2625,In_930,In_1079);
or U2626 (N_2626,In_1364,In_1322);
nor U2627 (N_2627,In_77,In_864);
nor U2628 (N_2628,In_230,In_1336);
xor U2629 (N_2629,In_1427,In_1449);
or U2630 (N_2630,In_157,In_1122);
or U2631 (N_2631,In_202,In_21);
or U2632 (N_2632,In_1467,In_1386);
xnor U2633 (N_2633,In_1377,In_432);
xor U2634 (N_2634,In_1187,In_674);
xnor U2635 (N_2635,In_402,In_240);
and U2636 (N_2636,In_533,In_1415);
nor U2637 (N_2637,In_1092,In_813);
nor U2638 (N_2638,In_1345,In_792);
xor U2639 (N_2639,In_250,In_191);
or U2640 (N_2640,In_115,In_476);
nor U2641 (N_2641,In_390,In_113);
and U2642 (N_2642,In_177,In_1108);
nor U2643 (N_2643,In_156,In_1254);
or U2644 (N_2644,In_1318,In_1169);
xor U2645 (N_2645,In_807,In_915);
xnor U2646 (N_2646,In_252,In_1220);
nor U2647 (N_2647,In_112,In_265);
nor U2648 (N_2648,In_634,In_1434);
or U2649 (N_2649,In_402,In_65);
nand U2650 (N_2650,In_329,In_823);
nor U2651 (N_2651,In_773,In_1075);
xor U2652 (N_2652,In_395,In_1155);
or U2653 (N_2653,In_1227,In_758);
or U2654 (N_2654,In_1073,In_321);
and U2655 (N_2655,In_1116,In_7);
nor U2656 (N_2656,In_459,In_1251);
xor U2657 (N_2657,In_970,In_1237);
nand U2658 (N_2658,In_1013,In_17);
and U2659 (N_2659,In_548,In_1468);
nand U2660 (N_2660,In_858,In_925);
or U2661 (N_2661,In_190,In_908);
and U2662 (N_2662,In_1012,In_127);
xnor U2663 (N_2663,In_162,In_1180);
or U2664 (N_2664,In_412,In_892);
nor U2665 (N_2665,In_911,In_236);
xor U2666 (N_2666,In_796,In_389);
nor U2667 (N_2667,In_846,In_765);
or U2668 (N_2668,In_1176,In_46);
nor U2669 (N_2669,In_657,In_1479);
or U2670 (N_2670,In_1232,In_156);
xor U2671 (N_2671,In_938,In_1213);
and U2672 (N_2672,In_359,In_331);
nand U2673 (N_2673,In_962,In_494);
or U2674 (N_2674,In_1196,In_1446);
xnor U2675 (N_2675,In_1350,In_28);
and U2676 (N_2676,In_1061,In_684);
or U2677 (N_2677,In_1095,In_22);
nor U2678 (N_2678,In_838,In_1135);
nand U2679 (N_2679,In_1331,In_511);
or U2680 (N_2680,In_142,In_240);
nor U2681 (N_2681,In_403,In_1113);
and U2682 (N_2682,In_803,In_166);
and U2683 (N_2683,In_613,In_407);
or U2684 (N_2684,In_458,In_896);
and U2685 (N_2685,In_789,In_1413);
nand U2686 (N_2686,In_1304,In_1349);
nor U2687 (N_2687,In_394,In_680);
nor U2688 (N_2688,In_1254,In_451);
nor U2689 (N_2689,In_1128,In_1024);
and U2690 (N_2690,In_1370,In_1020);
xnor U2691 (N_2691,In_603,In_542);
or U2692 (N_2692,In_1334,In_645);
xor U2693 (N_2693,In_1020,In_503);
xnor U2694 (N_2694,In_631,In_1345);
and U2695 (N_2695,In_745,In_1031);
xnor U2696 (N_2696,In_1050,In_77);
nor U2697 (N_2697,In_351,In_556);
nand U2698 (N_2698,In_824,In_249);
nor U2699 (N_2699,In_702,In_1115);
and U2700 (N_2700,In_1474,In_617);
xor U2701 (N_2701,In_1327,In_1227);
nand U2702 (N_2702,In_854,In_992);
or U2703 (N_2703,In_1444,In_565);
nor U2704 (N_2704,In_425,In_513);
nand U2705 (N_2705,In_1023,In_471);
or U2706 (N_2706,In_63,In_717);
nand U2707 (N_2707,In_614,In_589);
xnor U2708 (N_2708,In_1279,In_698);
and U2709 (N_2709,In_278,In_1196);
xor U2710 (N_2710,In_21,In_470);
and U2711 (N_2711,In_749,In_449);
or U2712 (N_2712,In_1309,In_68);
xnor U2713 (N_2713,In_745,In_920);
nor U2714 (N_2714,In_990,In_1009);
nor U2715 (N_2715,In_1109,In_1469);
xor U2716 (N_2716,In_1351,In_209);
and U2717 (N_2717,In_130,In_402);
nor U2718 (N_2718,In_858,In_414);
nor U2719 (N_2719,In_1002,In_1278);
or U2720 (N_2720,In_878,In_606);
or U2721 (N_2721,In_84,In_1038);
or U2722 (N_2722,In_1435,In_468);
xnor U2723 (N_2723,In_483,In_1423);
and U2724 (N_2724,In_656,In_216);
nand U2725 (N_2725,In_1052,In_978);
and U2726 (N_2726,In_194,In_688);
or U2727 (N_2727,In_1180,In_1047);
or U2728 (N_2728,In_1041,In_1315);
or U2729 (N_2729,In_584,In_1024);
or U2730 (N_2730,In_959,In_312);
nand U2731 (N_2731,In_779,In_231);
xor U2732 (N_2732,In_779,In_1498);
or U2733 (N_2733,In_483,In_1272);
nand U2734 (N_2734,In_889,In_393);
nor U2735 (N_2735,In_579,In_798);
or U2736 (N_2736,In_1245,In_595);
nor U2737 (N_2737,In_1273,In_1238);
nand U2738 (N_2738,In_633,In_1473);
or U2739 (N_2739,In_372,In_656);
xor U2740 (N_2740,In_1149,In_1070);
or U2741 (N_2741,In_1053,In_857);
and U2742 (N_2742,In_908,In_555);
nand U2743 (N_2743,In_225,In_1189);
nand U2744 (N_2744,In_954,In_188);
or U2745 (N_2745,In_689,In_131);
and U2746 (N_2746,In_623,In_929);
nand U2747 (N_2747,In_1370,In_1367);
or U2748 (N_2748,In_1034,In_1220);
nand U2749 (N_2749,In_1034,In_1094);
and U2750 (N_2750,In_89,In_294);
xor U2751 (N_2751,In_821,In_909);
and U2752 (N_2752,In_1068,In_936);
and U2753 (N_2753,In_1306,In_496);
nor U2754 (N_2754,In_577,In_853);
nor U2755 (N_2755,In_1293,In_899);
xor U2756 (N_2756,In_1053,In_1183);
or U2757 (N_2757,In_1456,In_1117);
nand U2758 (N_2758,In_259,In_316);
nand U2759 (N_2759,In_84,In_822);
nor U2760 (N_2760,In_871,In_786);
and U2761 (N_2761,In_753,In_784);
or U2762 (N_2762,In_72,In_423);
and U2763 (N_2763,In_868,In_244);
xnor U2764 (N_2764,In_802,In_584);
nand U2765 (N_2765,In_1434,In_1250);
xnor U2766 (N_2766,In_671,In_50);
or U2767 (N_2767,In_1061,In_1083);
or U2768 (N_2768,In_20,In_1192);
xnor U2769 (N_2769,In_124,In_1464);
or U2770 (N_2770,In_1124,In_1469);
or U2771 (N_2771,In_744,In_1427);
or U2772 (N_2772,In_617,In_959);
xnor U2773 (N_2773,In_400,In_264);
nor U2774 (N_2774,In_1180,In_1419);
and U2775 (N_2775,In_179,In_251);
and U2776 (N_2776,In_844,In_843);
xnor U2777 (N_2777,In_20,In_841);
xor U2778 (N_2778,In_284,In_192);
and U2779 (N_2779,In_358,In_652);
and U2780 (N_2780,In_133,In_667);
or U2781 (N_2781,In_1285,In_1446);
nand U2782 (N_2782,In_1180,In_239);
and U2783 (N_2783,In_119,In_633);
nand U2784 (N_2784,In_853,In_536);
or U2785 (N_2785,In_1277,In_848);
nand U2786 (N_2786,In_1204,In_1484);
and U2787 (N_2787,In_1309,In_983);
or U2788 (N_2788,In_379,In_367);
xnor U2789 (N_2789,In_1123,In_608);
nor U2790 (N_2790,In_1372,In_510);
xor U2791 (N_2791,In_985,In_62);
nor U2792 (N_2792,In_115,In_636);
and U2793 (N_2793,In_179,In_1262);
nand U2794 (N_2794,In_1349,In_625);
or U2795 (N_2795,In_203,In_629);
xor U2796 (N_2796,In_962,In_2);
nand U2797 (N_2797,In_169,In_1424);
nand U2798 (N_2798,In_541,In_259);
nor U2799 (N_2799,In_1173,In_932);
or U2800 (N_2800,In_739,In_111);
or U2801 (N_2801,In_790,In_1134);
or U2802 (N_2802,In_255,In_549);
nand U2803 (N_2803,In_699,In_93);
xnor U2804 (N_2804,In_702,In_781);
nand U2805 (N_2805,In_288,In_417);
or U2806 (N_2806,In_48,In_594);
nor U2807 (N_2807,In_352,In_856);
xnor U2808 (N_2808,In_146,In_1423);
and U2809 (N_2809,In_1375,In_371);
xor U2810 (N_2810,In_1470,In_225);
or U2811 (N_2811,In_335,In_37);
or U2812 (N_2812,In_694,In_1201);
nor U2813 (N_2813,In_488,In_1259);
and U2814 (N_2814,In_152,In_1139);
or U2815 (N_2815,In_930,In_629);
xor U2816 (N_2816,In_946,In_940);
nand U2817 (N_2817,In_716,In_575);
nor U2818 (N_2818,In_829,In_395);
nand U2819 (N_2819,In_344,In_1058);
nand U2820 (N_2820,In_1108,In_619);
and U2821 (N_2821,In_565,In_760);
nand U2822 (N_2822,In_1029,In_578);
or U2823 (N_2823,In_1348,In_1246);
nor U2824 (N_2824,In_940,In_630);
nor U2825 (N_2825,In_142,In_1109);
nor U2826 (N_2826,In_796,In_396);
nor U2827 (N_2827,In_1175,In_272);
and U2828 (N_2828,In_1429,In_420);
xnor U2829 (N_2829,In_361,In_8);
and U2830 (N_2830,In_208,In_966);
xnor U2831 (N_2831,In_1088,In_365);
nand U2832 (N_2832,In_950,In_630);
and U2833 (N_2833,In_133,In_780);
and U2834 (N_2834,In_93,In_111);
xor U2835 (N_2835,In_12,In_251);
xnor U2836 (N_2836,In_1375,In_1295);
or U2837 (N_2837,In_48,In_758);
or U2838 (N_2838,In_931,In_142);
nand U2839 (N_2839,In_726,In_1204);
and U2840 (N_2840,In_244,In_1254);
or U2841 (N_2841,In_1157,In_103);
and U2842 (N_2842,In_596,In_85);
nor U2843 (N_2843,In_165,In_1430);
xor U2844 (N_2844,In_879,In_351);
xor U2845 (N_2845,In_663,In_1246);
xnor U2846 (N_2846,In_127,In_1155);
nor U2847 (N_2847,In_879,In_1029);
and U2848 (N_2848,In_1081,In_833);
nand U2849 (N_2849,In_1321,In_737);
or U2850 (N_2850,In_810,In_169);
xor U2851 (N_2851,In_836,In_169);
nor U2852 (N_2852,In_807,In_561);
or U2853 (N_2853,In_25,In_2);
nand U2854 (N_2854,In_909,In_1124);
nor U2855 (N_2855,In_1203,In_493);
or U2856 (N_2856,In_1053,In_1112);
nand U2857 (N_2857,In_51,In_1487);
nand U2858 (N_2858,In_238,In_1315);
nand U2859 (N_2859,In_839,In_1197);
and U2860 (N_2860,In_868,In_1145);
or U2861 (N_2861,In_159,In_1318);
or U2862 (N_2862,In_996,In_219);
xnor U2863 (N_2863,In_965,In_1300);
nand U2864 (N_2864,In_852,In_61);
and U2865 (N_2865,In_1423,In_626);
xnor U2866 (N_2866,In_1093,In_16);
and U2867 (N_2867,In_1010,In_1489);
or U2868 (N_2868,In_1155,In_1214);
nor U2869 (N_2869,In_1433,In_1467);
nand U2870 (N_2870,In_257,In_373);
or U2871 (N_2871,In_1102,In_355);
nand U2872 (N_2872,In_214,In_888);
and U2873 (N_2873,In_799,In_1087);
and U2874 (N_2874,In_847,In_1425);
nand U2875 (N_2875,In_259,In_637);
nor U2876 (N_2876,In_1249,In_1287);
nor U2877 (N_2877,In_1065,In_971);
nor U2878 (N_2878,In_683,In_1447);
or U2879 (N_2879,In_24,In_1308);
nand U2880 (N_2880,In_1211,In_659);
or U2881 (N_2881,In_427,In_566);
and U2882 (N_2882,In_1071,In_850);
nand U2883 (N_2883,In_1405,In_1464);
nor U2884 (N_2884,In_1101,In_642);
xnor U2885 (N_2885,In_689,In_38);
and U2886 (N_2886,In_573,In_703);
xor U2887 (N_2887,In_374,In_808);
nand U2888 (N_2888,In_331,In_1003);
and U2889 (N_2889,In_476,In_269);
nand U2890 (N_2890,In_920,In_90);
nor U2891 (N_2891,In_1444,In_1358);
and U2892 (N_2892,In_377,In_1214);
and U2893 (N_2893,In_289,In_1043);
nand U2894 (N_2894,In_1440,In_1430);
nand U2895 (N_2895,In_586,In_296);
and U2896 (N_2896,In_679,In_1033);
xor U2897 (N_2897,In_639,In_938);
nand U2898 (N_2898,In_901,In_214);
xor U2899 (N_2899,In_734,In_349);
nand U2900 (N_2900,In_979,In_140);
or U2901 (N_2901,In_573,In_579);
nor U2902 (N_2902,In_250,In_1474);
or U2903 (N_2903,In_936,In_415);
or U2904 (N_2904,In_1401,In_1022);
nand U2905 (N_2905,In_1372,In_1459);
xnor U2906 (N_2906,In_1307,In_1013);
and U2907 (N_2907,In_1498,In_372);
nor U2908 (N_2908,In_293,In_312);
nand U2909 (N_2909,In_608,In_551);
nor U2910 (N_2910,In_1014,In_1222);
or U2911 (N_2911,In_269,In_749);
and U2912 (N_2912,In_29,In_540);
or U2913 (N_2913,In_1246,In_1306);
and U2914 (N_2914,In_354,In_976);
nor U2915 (N_2915,In_1004,In_247);
or U2916 (N_2916,In_317,In_1273);
or U2917 (N_2917,In_551,In_641);
nand U2918 (N_2918,In_1321,In_1427);
nor U2919 (N_2919,In_689,In_1044);
nand U2920 (N_2920,In_41,In_1310);
xnor U2921 (N_2921,In_292,In_1272);
nand U2922 (N_2922,In_507,In_1264);
xnor U2923 (N_2923,In_678,In_403);
or U2924 (N_2924,In_253,In_1438);
nand U2925 (N_2925,In_734,In_298);
nor U2926 (N_2926,In_712,In_151);
or U2927 (N_2927,In_53,In_562);
or U2928 (N_2928,In_1129,In_113);
nor U2929 (N_2929,In_889,In_719);
nor U2930 (N_2930,In_1381,In_775);
xnor U2931 (N_2931,In_1086,In_29);
nor U2932 (N_2932,In_1455,In_280);
or U2933 (N_2933,In_621,In_210);
nor U2934 (N_2934,In_160,In_1462);
nand U2935 (N_2935,In_1072,In_885);
and U2936 (N_2936,In_771,In_723);
nor U2937 (N_2937,In_764,In_325);
xnor U2938 (N_2938,In_237,In_204);
or U2939 (N_2939,In_336,In_244);
nor U2940 (N_2940,In_1133,In_452);
or U2941 (N_2941,In_683,In_1472);
nand U2942 (N_2942,In_796,In_945);
and U2943 (N_2943,In_921,In_76);
or U2944 (N_2944,In_8,In_166);
or U2945 (N_2945,In_286,In_994);
and U2946 (N_2946,In_16,In_1042);
xnor U2947 (N_2947,In_41,In_865);
nor U2948 (N_2948,In_1014,In_916);
xor U2949 (N_2949,In_885,In_1097);
or U2950 (N_2950,In_1104,In_1097);
xor U2951 (N_2951,In_780,In_1298);
xor U2952 (N_2952,In_397,In_147);
and U2953 (N_2953,In_1449,In_1166);
and U2954 (N_2954,In_1042,In_730);
nand U2955 (N_2955,In_96,In_1198);
nor U2956 (N_2956,In_1361,In_1285);
and U2957 (N_2957,In_1277,In_595);
nand U2958 (N_2958,In_118,In_224);
nand U2959 (N_2959,In_867,In_944);
nand U2960 (N_2960,In_1282,In_709);
nor U2961 (N_2961,In_1499,In_1022);
or U2962 (N_2962,In_54,In_635);
nand U2963 (N_2963,In_1354,In_1291);
xnor U2964 (N_2964,In_1424,In_1309);
xor U2965 (N_2965,In_1110,In_1279);
and U2966 (N_2966,In_1317,In_484);
nor U2967 (N_2967,In_587,In_220);
nor U2968 (N_2968,In_435,In_1322);
and U2969 (N_2969,In_377,In_33);
xor U2970 (N_2970,In_759,In_8);
and U2971 (N_2971,In_1377,In_1249);
nand U2972 (N_2972,In_158,In_1350);
nor U2973 (N_2973,In_1373,In_1461);
xor U2974 (N_2974,In_859,In_894);
and U2975 (N_2975,In_213,In_4);
nand U2976 (N_2976,In_1182,In_1061);
xnor U2977 (N_2977,In_126,In_652);
xnor U2978 (N_2978,In_125,In_504);
nor U2979 (N_2979,In_782,In_1187);
xor U2980 (N_2980,In_97,In_1233);
nor U2981 (N_2981,In_1474,In_1268);
or U2982 (N_2982,In_1167,In_1307);
or U2983 (N_2983,In_713,In_1332);
xnor U2984 (N_2984,In_697,In_390);
or U2985 (N_2985,In_1290,In_772);
xor U2986 (N_2986,In_153,In_301);
and U2987 (N_2987,In_1170,In_1342);
or U2988 (N_2988,In_766,In_805);
nor U2989 (N_2989,In_1018,In_278);
nor U2990 (N_2990,In_213,In_526);
nor U2991 (N_2991,In_463,In_1136);
or U2992 (N_2992,In_530,In_220);
and U2993 (N_2993,In_335,In_659);
and U2994 (N_2994,In_1253,In_939);
or U2995 (N_2995,In_1252,In_754);
nand U2996 (N_2996,In_1264,In_917);
xnor U2997 (N_2997,In_187,In_1237);
xnor U2998 (N_2998,In_901,In_116);
or U2999 (N_2999,In_553,In_825);
nor U3000 (N_3000,In_368,In_500);
and U3001 (N_3001,In_840,In_1149);
xnor U3002 (N_3002,In_974,In_799);
nand U3003 (N_3003,In_431,In_1313);
xnor U3004 (N_3004,In_645,In_510);
and U3005 (N_3005,In_43,In_1163);
and U3006 (N_3006,In_745,In_664);
or U3007 (N_3007,In_1487,In_665);
nor U3008 (N_3008,In_72,In_687);
nor U3009 (N_3009,In_513,In_1450);
nor U3010 (N_3010,In_607,In_273);
or U3011 (N_3011,In_527,In_980);
nor U3012 (N_3012,In_770,In_1313);
nor U3013 (N_3013,In_626,In_1096);
nor U3014 (N_3014,In_352,In_1271);
nor U3015 (N_3015,In_984,In_1028);
and U3016 (N_3016,In_1183,In_1133);
and U3017 (N_3017,In_1197,In_1060);
nand U3018 (N_3018,In_406,In_38);
xor U3019 (N_3019,In_169,In_271);
xnor U3020 (N_3020,In_1345,In_839);
nand U3021 (N_3021,In_609,In_671);
nor U3022 (N_3022,In_135,In_1169);
xnor U3023 (N_3023,In_784,In_445);
or U3024 (N_3024,In_1282,In_474);
nor U3025 (N_3025,In_1407,In_748);
or U3026 (N_3026,In_1370,In_958);
and U3027 (N_3027,In_423,In_1210);
or U3028 (N_3028,In_282,In_34);
xor U3029 (N_3029,In_576,In_1090);
or U3030 (N_3030,In_58,In_457);
or U3031 (N_3031,In_909,In_1269);
xnor U3032 (N_3032,In_1213,In_77);
xnor U3033 (N_3033,In_926,In_1275);
xor U3034 (N_3034,In_729,In_47);
nand U3035 (N_3035,In_1290,In_178);
or U3036 (N_3036,In_1209,In_577);
xor U3037 (N_3037,In_289,In_1210);
xor U3038 (N_3038,In_1262,In_1278);
or U3039 (N_3039,In_1402,In_1118);
or U3040 (N_3040,In_1133,In_1446);
nand U3041 (N_3041,In_691,In_1194);
nor U3042 (N_3042,In_291,In_1158);
nor U3043 (N_3043,In_594,In_844);
nand U3044 (N_3044,In_621,In_1061);
xnor U3045 (N_3045,In_911,In_20);
nand U3046 (N_3046,In_126,In_131);
nand U3047 (N_3047,In_1338,In_39);
and U3048 (N_3048,In_1100,In_404);
nor U3049 (N_3049,In_1006,In_576);
xor U3050 (N_3050,In_240,In_608);
xnor U3051 (N_3051,In_1047,In_1365);
nand U3052 (N_3052,In_644,In_831);
and U3053 (N_3053,In_1071,In_263);
nand U3054 (N_3054,In_1288,In_516);
nor U3055 (N_3055,In_1175,In_1346);
nor U3056 (N_3056,In_785,In_1220);
nor U3057 (N_3057,In_152,In_1431);
and U3058 (N_3058,In_731,In_1105);
nor U3059 (N_3059,In_235,In_492);
and U3060 (N_3060,In_1069,In_1419);
and U3061 (N_3061,In_379,In_884);
nand U3062 (N_3062,In_1265,In_404);
xnor U3063 (N_3063,In_189,In_1202);
xnor U3064 (N_3064,In_604,In_1330);
nor U3065 (N_3065,In_1262,In_797);
nor U3066 (N_3066,In_561,In_1410);
nor U3067 (N_3067,In_2,In_697);
xor U3068 (N_3068,In_902,In_946);
nor U3069 (N_3069,In_728,In_898);
or U3070 (N_3070,In_392,In_936);
xnor U3071 (N_3071,In_973,In_452);
and U3072 (N_3072,In_1140,In_1000);
xnor U3073 (N_3073,In_1456,In_295);
or U3074 (N_3074,In_945,In_1028);
and U3075 (N_3075,In_1478,In_973);
nand U3076 (N_3076,In_488,In_284);
xor U3077 (N_3077,In_995,In_974);
and U3078 (N_3078,In_1341,In_347);
nor U3079 (N_3079,In_107,In_519);
or U3080 (N_3080,In_834,In_879);
xnor U3081 (N_3081,In_1407,In_556);
nor U3082 (N_3082,In_90,In_535);
and U3083 (N_3083,In_1253,In_886);
nor U3084 (N_3084,In_940,In_290);
nor U3085 (N_3085,In_1272,In_1260);
xor U3086 (N_3086,In_11,In_162);
and U3087 (N_3087,In_217,In_369);
nand U3088 (N_3088,In_1451,In_1410);
nand U3089 (N_3089,In_1050,In_482);
or U3090 (N_3090,In_298,In_787);
nand U3091 (N_3091,In_1090,In_94);
nand U3092 (N_3092,In_65,In_814);
or U3093 (N_3093,In_622,In_1497);
or U3094 (N_3094,In_418,In_1463);
and U3095 (N_3095,In_1040,In_77);
or U3096 (N_3096,In_362,In_188);
and U3097 (N_3097,In_396,In_1303);
xor U3098 (N_3098,In_1220,In_1441);
and U3099 (N_3099,In_615,In_1291);
xnor U3100 (N_3100,In_1069,In_635);
nand U3101 (N_3101,In_230,In_17);
or U3102 (N_3102,In_806,In_1100);
and U3103 (N_3103,In_163,In_2);
or U3104 (N_3104,In_868,In_104);
nand U3105 (N_3105,In_153,In_614);
nor U3106 (N_3106,In_350,In_284);
xnor U3107 (N_3107,In_809,In_78);
xor U3108 (N_3108,In_835,In_1293);
nor U3109 (N_3109,In_401,In_1133);
and U3110 (N_3110,In_537,In_41);
or U3111 (N_3111,In_198,In_1052);
or U3112 (N_3112,In_630,In_236);
xor U3113 (N_3113,In_678,In_723);
or U3114 (N_3114,In_142,In_1302);
nand U3115 (N_3115,In_1120,In_915);
or U3116 (N_3116,In_1403,In_207);
xnor U3117 (N_3117,In_1148,In_16);
nor U3118 (N_3118,In_596,In_164);
and U3119 (N_3119,In_1164,In_918);
xor U3120 (N_3120,In_668,In_1064);
or U3121 (N_3121,In_1295,In_1115);
or U3122 (N_3122,In_879,In_121);
nand U3123 (N_3123,In_216,In_844);
nand U3124 (N_3124,In_322,In_1290);
xnor U3125 (N_3125,In_19,In_1159);
or U3126 (N_3126,In_1490,In_209);
or U3127 (N_3127,In_1061,In_498);
and U3128 (N_3128,In_42,In_538);
nand U3129 (N_3129,In_1128,In_1146);
xnor U3130 (N_3130,In_732,In_1361);
xor U3131 (N_3131,In_383,In_497);
nand U3132 (N_3132,In_101,In_970);
nor U3133 (N_3133,In_1012,In_1173);
xnor U3134 (N_3134,In_1293,In_1071);
nand U3135 (N_3135,In_877,In_44);
nor U3136 (N_3136,In_1172,In_742);
nor U3137 (N_3137,In_918,In_1374);
xor U3138 (N_3138,In_16,In_2);
xnor U3139 (N_3139,In_1341,In_111);
xnor U3140 (N_3140,In_709,In_1456);
nand U3141 (N_3141,In_962,In_771);
and U3142 (N_3142,In_1253,In_1255);
and U3143 (N_3143,In_181,In_688);
or U3144 (N_3144,In_1089,In_755);
nor U3145 (N_3145,In_1004,In_446);
xnor U3146 (N_3146,In_1170,In_344);
and U3147 (N_3147,In_763,In_664);
or U3148 (N_3148,In_744,In_1173);
xor U3149 (N_3149,In_807,In_751);
nand U3150 (N_3150,In_1448,In_736);
nand U3151 (N_3151,In_1435,In_341);
nor U3152 (N_3152,In_265,In_1432);
xor U3153 (N_3153,In_119,In_647);
nand U3154 (N_3154,In_547,In_460);
nand U3155 (N_3155,In_1488,In_758);
or U3156 (N_3156,In_1134,In_1155);
and U3157 (N_3157,In_212,In_507);
and U3158 (N_3158,In_669,In_20);
nand U3159 (N_3159,In_336,In_1347);
or U3160 (N_3160,In_723,In_273);
nand U3161 (N_3161,In_1103,In_488);
xnor U3162 (N_3162,In_842,In_1397);
or U3163 (N_3163,In_1215,In_1297);
or U3164 (N_3164,In_938,In_777);
xnor U3165 (N_3165,In_1225,In_116);
nor U3166 (N_3166,In_1011,In_1040);
nor U3167 (N_3167,In_242,In_208);
and U3168 (N_3168,In_1274,In_1484);
or U3169 (N_3169,In_72,In_680);
and U3170 (N_3170,In_357,In_603);
nand U3171 (N_3171,In_32,In_1006);
nand U3172 (N_3172,In_123,In_1321);
and U3173 (N_3173,In_802,In_707);
and U3174 (N_3174,In_562,In_348);
or U3175 (N_3175,In_547,In_388);
or U3176 (N_3176,In_809,In_1301);
or U3177 (N_3177,In_697,In_1154);
and U3178 (N_3178,In_641,In_1491);
or U3179 (N_3179,In_997,In_1009);
nor U3180 (N_3180,In_157,In_991);
nand U3181 (N_3181,In_746,In_869);
nand U3182 (N_3182,In_1483,In_465);
xor U3183 (N_3183,In_41,In_826);
xnor U3184 (N_3184,In_1246,In_122);
or U3185 (N_3185,In_56,In_448);
xor U3186 (N_3186,In_337,In_1066);
or U3187 (N_3187,In_1126,In_963);
nand U3188 (N_3188,In_1049,In_1255);
nand U3189 (N_3189,In_2,In_892);
and U3190 (N_3190,In_295,In_787);
nand U3191 (N_3191,In_718,In_1385);
nor U3192 (N_3192,In_58,In_285);
xor U3193 (N_3193,In_1383,In_679);
or U3194 (N_3194,In_277,In_1206);
nand U3195 (N_3195,In_531,In_990);
nand U3196 (N_3196,In_876,In_539);
nand U3197 (N_3197,In_1011,In_301);
xnor U3198 (N_3198,In_1221,In_338);
xor U3199 (N_3199,In_487,In_72);
xor U3200 (N_3200,In_389,In_802);
nand U3201 (N_3201,In_175,In_570);
or U3202 (N_3202,In_1241,In_1212);
xnor U3203 (N_3203,In_182,In_210);
and U3204 (N_3204,In_1369,In_920);
and U3205 (N_3205,In_548,In_779);
xnor U3206 (N_3206,In_1173,In_726);
or U3207 (N_3207,In_584,In_13);
and U3208 (N_3208,In_331,In_996);
nor U3209 (N_3209,In_1246,In_211);
nand U3210 (N_3210,In_465,In_978);
xor U3211 (N_3211,In_1164,In_1461);
or U3212 (N_3212,In_653,In_343);
and U3213 (N_3213,In_155,In_365);
nor U3214 (N_3214,In_82,In_1098);
nand U3215 (N_3215,In_198,In_1463);
nor U3216 (N_3216,In_1095,In_594);
nor U3217 (N_3217,In_1381,In_1011);
xnor U3218 (N_3218,In_1254,In_1066);
xor U3219 (N_3219,In_352,In_1472);
nor U3220 (N_3220,In_1138,In_546);
xnor U3221 (N_3221,In_658,In_58);
or U3222 (N_3222,In_298,In_308);
xnor U3223 (N_3223,In_1404,In_731);
or U3224 (N_3224,In_887,In_362);
nor U3225 (N_3225,In_453,In_957);
nor U3226 (N_3226,In_1332,In_735);
nor U3227 (N_3227,In_219,In_1003);
xnor U3228 (N_3228,In_1287,In_1375);
nor U3229 (N_3229,In_761,In_357);
xnor U3230 (N_3230,In_1427,In_999);
nand U3231 (N_3231,In_767,In_1401);
nand U3232 (N_3232,In_302,In_807);
or U3233 (N_3233,In_1305,In_1258);
or U3234 (N_3234,In_1202,In_753);
or U3235 (N_3235,In_746,In_237);
xnor U3236 (N_3236,In_106,In_189);
nand U3237 (N_3237,In_1473,In_1478);
or U3238 (N_3238,In_612,In_1365);
nand U3239 (N_3239,In_604,In_29);
and U3240 (N_3240,In_118,In_1405);
or U3241 (N_3241,In_1325,In_473);
nand U3242 (N_3242,In_547,In_971);
nand U3243 (N_3243,In_630,In_995);
or U3244 (N_3244,In_879,In_230);
nand U3245 (N_3245,In_622,In_719);
nor U3246 (N_3246,In_689,In_263);
nand U3247 (N_3247,In_671,In_292);
nand U3248 (N_3248,In_659,In_681);
or U3249 (N_3249,In_1067,In_473);
xor U3250 (N_3250,In_1116,In_999);
nor U3251 (N_3251,In_682,In_1099);
nand U3252 (N_3252,In_605,In_1028);
or U3253 (N_3253,In_1257,In_656);
and U3254 (N_3254,In_1349,In_1059);
nand U3255 (N_3255,In_545,In_479);
nand U3256 (N_3256,In_504,In_734);
nand U3257 (N_3257,In_252,In_960);
nand U3258 (N_3258,In_552,In_788);
and U3259 (N_3259,In_123,In_390);
nand U3260 (N_3260,In_220,In_173);
or U3261 (N_3261,In_736,In_394);
and U3262 (N_3262,In_1193,In_1341);
nand U3263 (N_3263,In_1463,In_211);
or U3264 (N_3264,In_1438,In_1440);
nor U3265 (N_3265,In_1444,In_306);
nor U3266 (N_3266,In_274,In_747);
nand U3267 (N_3267,In_1105,In_179);
nand U3268 (N_3268,In_676,In_1370);
nor U3269 (N_3269,In_1240,In_303);
nand U3270 (N_3270,In_1347,In_515);
and U3271 (N_3271,In_1108,In_1465);
and U3272 (N_3272,In_572,In_676);
nand U3273 (N_3273,In_128,In_11);
nor U3274 (N_3274,In_401,In_1111);
or U3275 (N_3275,In_1061,In_77);
or U3276 (N_3276,In_93,In_210);
or U3277 (N_3277,In_692,In_838);
or U3278 (N_3278,In_280,In_740);
nor U3279 (N_3279,In_167,In_1114);
and U3280 (N_3280,In_568,In_412);
or U3281 (N_3281,In_1061,In_990);
xor U3282 (N_3282,In_424,In_140);
nor U3283 (N_3283,In_929,In_1041);
nor U3284 (N_3284,In_620,In_476);
and U3285 (N_3285,In_18,In_340);
and U3286 (N_3286,In_388,In_293);
nand U3287 (N_3287,In_1284,In_522);
or U3288 (N_3288,In_1001,In_1124);
or U3289 (N_3289,In_447,In_284);
nor U3290 (N_3290,In_1078,In_785);
nand U3291 (N_3291,In_1288,In_649);
nor U3292 (N_3292,In_147,In_1438);
nor U3293 (N_3293,In_795,In_203);
xnor U3294 (N_3294,In_880,In_483);
and U3295 (N_3295,In_842,In_1248);
and U3296 (N_3296,In_1242,In_488);
nand U3297 (N_3297,In_1301,In_988);
xnor U3298 (N_3298,In_979,In_1200);
or U3299 (N_3299,In_224,In_673);
or U3300 (N_3300,In_549,In_200);
or U3301 (N_3301,In_345,In_566);
and U3302 (N_3302,In_1389,In_932);
xnor U3303 (N_3303,In_272,In_1274);
and U3304 (N_3304,In_250,In_239);
xnor U3305 (N_3305,In_158,In_424);
and U3306 (N_3306,In_127,In_717);
and U3307 (N_3307,In_1011,In_1130);
nor U3308 (N_3308,In_309,In_658);
and U3309 (N_3309,In_736,In_1154);
nor U3310 (N_3310,In_1211,In_1202);
and U3311 (N_3311,In_279,In_630);
or U3312 (N_3312,In_842,In_604);
xor U3313 (N_3313,In_1397,In_469);
xnor U3314 (N_3314,In_368,In_131);
nor U3315 (N_3315,In_437,In_592);
and U3316 (N_3316,In_61,In_510);
or U3317 (N_3317,In_478,In_1267);
nand U3318 (N_3318,In_1403,In_583);
nor U3319 (N_3319,In_48,In_235);
or U3320 (N_3320,In_1253,In_113);
nand U3321 (N_3321,In_235,In_880);
or U3322 (N_3322,In_1289,In_243);
nor U3323 (N_3323,In_1164,In_1446);
nor U3324 (N_3324,In_1262,In_1426);
xnor U3325 (N_3325,In_1394,In_477);
nor U3326 (N_3326,In_993,In_174);
nand U3327 (N_3327,In_463,In_1432);
xor U3328 (N_3328,In_828,In_579);
and U3329 (N_3329,In_804,In_515);
and U3330 (N_3330,In_1208,In_643);
and U3331 (N_3331,In_292,In_97);
or U3332 (N_3332,In_595,In_636);
xnor U3333 (N_3333,In_406,In_1300);
and U3334 (N_3334,In_1412,In_400);
and U3335 (N_3335,In_910,In_1169);
and U3336 (N_3336,In_1115,In_473);
nand U3337 (N_3337,In_587,In_439);
xnor U3338 (N_3338,In_1411,In_214);
or U3339 (N_3339,In_814,In_620);
nor U3340 (N_3340,In_664,In_1397);
nor U3341 (N_3341,In_1484,In_279);
and U3342 (N_3342,In_1093,In_474);
xnor U3343 (N_3343,In_1235,In_541);
xor U3344 (N_3344,In_261,In_485);
nor U3345 (N_3345,In_709,In_75);
nor U3346 (N_3346,In_15,In_302);
nor U3347 (N_3347,In_936,In_183);
xor U3348 (N_3348,In_264,In_101);
or U3349 (N_3349,In_968,In_748);
nor U3350 (N_3350,In_1273,In_610);
xnor U3351 (N_3351,In_592,In_672);
nor U3352 (N_3352,In_779,In_468);
xnor U3353 (N_3353,In_199,In_916);
nor U3354 (N_3354,In_1435,In_1364);
nor U3355 (N_3355,In_126,In_501);
or U3356 (N_3356,In_789,In_559);
nand U3357 (N_3357,In_141,In_680);
or U3358 (N_3358,In_557,In_1349);
and U3359 (N_3359,In_1168,In_800);
xor U3360 (N_3360,In_867,In_489);
nand U3361 (N_3361,In_456,In_1224);
nand U3362 (N_3362,In_548,In_687);
or U3363 (N_3363,In_141,In_776);
or U3364 (N_3364,In_261,In_1277);
and U3365 (N_3365,In_1037,In_1395);
or U3366 (N_3366,In_91,In_1094);
or U3367 (N_3367,In_1352,In_312);
nor U3368 (N_3368,In_1093,In_1440);
nor U3369 (N_3369,In_1087,In_1143);
nor U3370 (N_3370,In_1368,In_248);
nand U3371 (N_3371,In_1266,In_946);
or U3372 (N_3372,In_355,In_706);
nand U3373 (N_3373,In_958,In_956);
or U3374 (N_3374,In_606,In_801);
nand U3375 (N_3375,In_395,In_857);
or U3376 (N_3376,In_984,In_917);
xnor U3377 (N_3377,In_1336,In_130);
nand U3378 (N_3378,In_1114,In_722);
nor U3379 (N_3379,In_542,In_1317);
nand U3380 (N_3380,In_1466,In_620);
and U3381 (N_3381,In_755,In_470);
and U3382 (N_3382,In_375,In_597);
xnor U3383 (N_3383,In_120,In_135);
and U3384 (N_3384,In_1223,In_536);
xor U3385 (N_3385,In_991,In_50);
nand U3386 (N_3386,In_550,In_477);
xnor U3387 (N_3387,In_238,In_642);
or U3388 (N_3388,In_319,In_1282);
and U3389 (N_3389,In_848,In_726);
and U3390 (N_3390,In_4,In_1377);
xor U3391 (N_3391,In_1060,In_971);
xnor U3392 (N_3392,In_1294,In_644);
and U3393 (N_3393,In_1203,In_425);
nand U3394 (N_3394,In_525,In_428);
and U3395 (N_3395,In_144,In_1155);
nor U3396 (N_3396,In_1004,In_1020);
nand U3397 (N_3397,In_726,In_881);
and U3398 (N_3398,In_1034,In_812);
xnor U3399 (N_3399,In_576,In_910);
and U3400 (N_3400,In_478,In_281);
and U3401 (N_3401,In_1287,In_1051);
nor U3402 (N_3402,In_311,In_166);
nor U3403 (N_3403,In_1077,In_66);
xnor U3404 (N_3404,In_115,In_1499);
nand U3405 (N_3405,In_195,In_143);
xor U3406 (N_3406,In_588,In_415);
xor U3407 (N_3407,In_665,In_464);
or U3408 (N_3408,In_188,In_265);
nand U3409 (N_3409,In_1317,In_65);
or U3410 (N_3410,In_649,In_817);
nor U3411 (N_3411,In_1236,In_632);
nor U3412 (N_3412,In_665,In_1444);
nor U3413 (N_3413,In_1491,In_95);
nor U3414 (N_3414,In_472,In_1213);
and U3415 (N_3415,In_1293,In_1093);
nor U3416 (N_3416,In_1178,In_864);
nor U3417 (N_3417,In_1303,In_140);
xnor U3418 (N_3418,In_891,In_439);
and U3419 (N_3419,In_665,In_630);
nor U3420 (N_3420,In_1227,In_837);
xnor U3421 (N_3421,In_1359,In_406);
xnor U3422 (N_3422,In_765,In_47);
nand U3423 (N_3423,In_439,In_164);
or U3424 (N_3424,In_629,In_784);
nor U3425 (N_3425,In_292,In_1254);
and U3426 (N_3426,In_1030,In_986);
and U3427 (N_3427,In_106,In_147);
and U3428 (N_3428,In_908,In_460);
nand U3429 (N_3429,In_164,In_1149);
xnor U3430 (N_3430,In_842,In_1035);
or U3431 (N_3431,In_4,In_355);
nand U3432 (N_3432,In_1220,In_1447);
and U3433 (N_3433,In_1185,In_1477);
or U3434 (N_3434,In_543,In_1094);
and U3435 (N_3435,In_780,In_130);
xor U3436 (N_3436,In_1253,In_619);
xnor U3437 (N_3437,In_121,In_454);
and U3438 (N_3438,In_389,In_477);
nand U3439 (N_3439,In_1061,In_1475);
or U3440 (N_3440,In_378,In_1474);
or U3441 (N_3441,In_157,In_425);
xor U3442 (N_3442,In_602,In_466);
nand U3443 (N_3443,In_1108,In_1118);
nor U3444 (N_3444,In_546,In_1474);
or U3445 (N_3445,In_58,In_1235);
and U3446 (N_3446,In_704,In_209);
xor U3447 (N_3447,In_631,In_816);
xnor U3448 (N_3448,In_308,In_225);
xor U3449 (N_3449,In_883,In_1126);
xor U3450 (N_3450,In_892,In_152);
nand U3451 (N_3451,In_1333,In_231);
nor U3452 (N_3452,In_1178,In_1224);
and U3453 (N_3453,In_1232,In_1101);
xor U3454 (N_3454,In_964,In_894);
nand U3455 (N_3455,In_167,In_1243);
xnor U3456 (N_3456,In_1415,In_1061);
nand U3457 (N_3457,In_966,In_1183);
nor U3458 (N_3458,In_1459,In_13);
nor U3459 (N_3459,In_1286,In_1361);
and U3460 (N_3460,In_826,In_1140);
or U3461 (N_3461,In_52,In_1302);
or U3462 (N_3462,In_1190,In_504);
xnor U3463 (N_3463,In_1224,In_1471);
nand U3464 (N_3464,In_817,In_1030);
or U3465 (N_3465,In_663,In_877);
or U3466 (N_3466,In_749,In_1132);
nand U3467 (N_3467,In_782,In_1406);
nand U3468 (N_3468,In_66,In_641);
and U3469 (N_3469,In_615,In_723);
nand U3470 (N_3470,In_1141,In_1239);
xnor U3471 (N_3471,In_1273,In_250);
nand U3472 (N_3472,In_959,In_526);
or U3473 (N_3473,In_826,In_1164);
nor U3474 (N_3474,In_122,In_17);
and U3475 (N_3475,In_539,In_1214);
nand U3476 (N_3476,In_556,In_128);
and U3477 (N_3477,In_1339,In_237);
or U3478 (N_3478,In_1102,In_368);
nand U3479 (N_3479,In_1119,In_229);
nand U3480 (N_3480,In_1015,In_160);
and U3481 (N_3481,In_207,In_430);
nand U3482 (N_3482,In_610,In_108);
xnor U3483 (N_3483,In_1013,In_683);
nand U3484 (N_3484,In_1409,In_1233);
and U3485 (N_3485,In_595,In_1369);
or U3486 (N_3486,In_1453,In_1007);
and U3487 (N_3487,In_1159,In_288);
or U3488 (N_3488,In_1357,In_838);
nor U3489 (N_3489,In_406,In_186);
nand U3490 (N_3490,In_548,In_307);
nor U3491 (N_3491,In_278,In_164);
xnor U3492 (N_3492,In_791,In_298);
nand U3493 (N_3493,In_1124,In_1436);
nor U3494 (N_3494,In_1464,In_649);
nand U3495 (N_3495,In_282,In_1090);
and U3496 (N_3496,In_943,In_8);
and U3497 (N_3497,In_998,In_229);
xor U3498 (N_3498,In_1395,In_1375);
nand U3499 (N_3499,In_1473,In_304);
nor U3500 (N_3500,In_1057,In_392);
xnor U3501 (N_3501,In_151,In_425);
and U3502 (N_3502,In_806,In_611);
nand U3503 (N_3503,In_900,In_727);
nand U3504 (N_3504,In_645,In_558);
nand U3505 (N_3505,In_961,In_1095);
nand U3506 (N_3506,In_242,In_1173);
and U3507 (N_3507,In_368,In_1140);
xnor U3508 (N_3508,In_614,In_1023);
nor U3509 (N_3509,In_1325,In_1328);
or U3510 (N_3510,In_234,In_194);
nor U3511 (N_3511,In_161,In_1474);
or U3512 (N_3512,In_1497,In_303);
xnor U3513 (N_3513,In_138,In_1242);
xnor U3514 (N_3514,In_57,In_800);
or U3515 (N_3515,In_156,In_973);
nand U3516 (N_3516,In_1228,In_561);
xor U3517 (N_3517,In_1375,In_1263);
nand U3518 (N_3518,In_896,In_1208);
nor U3519 (N_3519,In_14,In_1416);
xnor U3520 (N_3520,In_1451,In_762);
or U3521 (N_3521,In_770,In_1223);
nand U3522 (N_3522,In_575,In_501);
xnor U3523 (N_3523,In_332,In_654);
and U3524 (N_3524,In_1377,In_250);
and U3525 (N_3525,In_1028,In_1152);
nor U3526 (N_3526,In_900,In_259);
or U3527 (N_3527,In_1381,In_1326);
or U3528 (N_3528,In_650,In_609);
nand U3529 (N_3529,In_1284,In_164);
and U3530 (N_3530,In_802,In_535);
nand U3531 (N_3531,In_299,In_273);
nand U3532 (N_3532,In_120,In_548);
nand U3533 (N_3533,In_884,In_1178);
or U3534 (N_3534,In_1472,In_310);
or U3535 (N_3535,In_34,In_114);
nor U3536 (N_3536,In_46,In_1414);
nor U3537 (N_3537,In_271,In_1342);
or U3538 (N_3538,In_1094,In_935);
xor U3539 (N_3539,In_1353,In_1423);
or U3540 (N_3540,In_980,In_567);
nand U3541 (N_3541,In_1357,In_527);
or U3542 (N_3542,In_1237,In_863);
or U3543 (N_3543,In_990,In_424);
nor U3544 (N_3544,In_863,In_1077);
nand U3545 (N_3545,In_453,In_500);
nor U3546 (N_3546,In_1305,In_704);
or U3547 (N_3547,In_1456,In_304);
nor U3548 (N_3548,In_1026,In_302);
or U3549 (N_3549,In_753,In_34);
xor U3550 (N_3550,In_1124,In_1122);
or U3551 (N_3551,In_724,In_1260);
or U3552 (N_3552,In_438,In_49);
xor U3553 (N_3553,In_1157,In_869);
or U3554 (N_3554,In_233,In_946);
nor U3555 (N_3555,In_543,In_392);
xor U3556 (N_3556,In_285,In_1435);
or U3557 (N_3557,In_1045,In_108);
nand U3558 (N_3558,In_505,In_288);
and U3559 (N_3559,In_476,In_926);
xor U3560 (N_3560,In_75,In_616);
or U3561 (N_3561,In_3,In_1096);
nand U3562 (N_3562,In_294,In_806);
or U3563 (N_3563,In_196,In_581);
nor U3564 (N_3564,In_849,In_1368);
nor U3565 (N_3565,In_942,In_350);
or U3566 (N_3566,In_699,In_99);
nor U3567 (N_3567,In_312,In_1064);
or U3568 (N_3568,In_714,In_1207);
nand U3569 (N_3569,In_392,In_329);
and U3570 (N_3570,In_1238,In_1190);
nor U3571 (N_3571,In_770,In_1395);
xnor U3572 (N_3572,In_1255,In_761);
nand U3573 (N_3573,In_287,In_238);
and U3574 (N_3574,In_271,In_642);
nor U3575 (N_3575,In_394,In_1289);
nand U3576 (N_3576,In_382,In_642);
or U3577 (N_3577,In_443,In_1124);
or U3578 (N_3578,In_743,In_1203);
nor U3579 (N_3579,In_1057,In_623);
xor U3580 (N_3580,In_589,In_1244);
and U3581 (N_3581,In_1054,In_435);
and U3582 (N_3582,In_698,In_669);
xnor U3583 (N_3583,In_428,In_1081);
or U3584 (N_3584,In_1285,In_1248);
nor U3585 (N_3585,In_90,In_1119);
or U3586 (N_3586,In_193,In_1458);
xnor U3587 (N_3587,In_839,In_300);
nand U3588 (N_3588,In_254,In_238);
xor U3589 (N_3589,In_368,In_560);
nand U3590 (N_3590,In_187,In_1002);
xnor U3591 (N_3591,In_1486,In_1127);
nand U3592 (N_3592,In_1214,In_372);
or U3593 (N_3593,In_503,In_490);
nand U3594 (N_3594,In_831,In_674);
and U3595 (N_3595,In_266,In_503);
or U3596 (N_3596,In_1073,In_525);
or U3597 (N_3597,In_704,In_1497);
nor U3598 (N_3598,In_1147,In_1067);
and U3599 (N_3599,In_765,In_1376);
and U3600 (N_3600,In_15,In_975);
nand U3601 (N_3601,In_508,In_796);
xnor U3602 (N_3602,In_967,In_559);
nand U3603 (N_3603,In_780,In_1203);
nand U3604 (N_3604,In_215,In_153);
xor U3605 (N_3605,In_1233,In_125);
and U3606 (N_3606,In_1031,In_736);
xor U3607 (N_3607,In_771,In_274);
or U3608 (N_3608,In_844,In_308);
xnor U3609 (N_3609,In_1270,In_256);
nor U3610 (N_3610,In_942,In_1429);
nor U3611 (N_3611,In_1470,In_863);
nand U3612 (N_3612,In_846,In_35);
xnor U3613 (N_3613,In_389,In_631);
or U3614 (N_3614,In_1308,In_1376);
nor U3615 (N_3615,In_1224,In_910);
or U3616 (N_3616,In_1391,In_1354);
nand U3617 (N_3617,In_39,In_1032);
nand U3618 (N_3618,In_28,In_672);
xor U3619 (N_3619,In_883,In_714);
or U3620 (N_3620,In_426,In_1021);
nor U3621 (N_3621,In_1212,In_927);
nand U3622 (N_3622,In_1477,In_1439);
or U3623 (N_3623,In_1129,In_32);
nor U3624 (N_3624,In_454,In_584);
xnor U3625 (N_3625,In_972,In_1054);
and U3626 (N_3626,In_1439,In_536);
nand U3627 (N_3627,In_35,In_609);
or U3628 (N_3628,In_269,In_765);
or U3629 (N_3629,In_681,In_122);
nor U3630 (N_3630,In_1377,In_323);
xor U3631 (N_3631,In_1048,In_607);
nor U3632 (N_3632,In_147,In_347);
nor U3633 (N_3633,In_1011,In_600);
nand U3634 (N_3634,In_487,In_577);
nor U3635 (N_3635,In_1063,In_459);
xor U3636 (N_3636,In_444,In_974);
or U3637 (N_3637,In_605,In_38);
nor U3638 (N_3638,In_676,In_1215);
nand U3639 (N_3639,In_1144,In_14);
xnor U3640 (N_3640,In_252,In_1100);
or U3641 (N_3641,In_1471,In_1280);
nor U3642 (N_3642,In_116,In_1065);
or U3643 (N_3643,In_877,In_1332);
nor U3644 (N_3644,In_1128,In_554);
or U3645 (N_3645,In_1215,In_1265);
xor U3646 (N_3646,In_888,In_958);
xor U3647 (N_3647,In_857,In_479);
or U3648 (N_3648,In_486,In_782);
nor U3649 (N_3649,In_1031,In_1424);
xnor U3650 (N_3650,In_123,In_476);
nor U3651 (N_3651,In_902,In_1200);
nand U3652 (N_3652,In_383,In_1026);
xor U3653 (N_3653,In_780,In_420);
xnor U3654 (N_3654,In_370,In_604);
nand U3655 (N_3655,In_727,In_958);
or U3656 (N_3656,In_1469,In_1300);
nor U3657 (N_3657,In_1251,In_1346);
and U3658 (N_3658,In_1250,In_1406);
and U3659 (N_3659,In_1423,In_281);
nand U3660 (N_3660,In_1309,In_1037);
xnor U3661 (N_3661,In_936,In_233);
nor U3662 (N_3662,In_1050,In_1085);
xor U3663 (N_3663,In_711,In_704);
and U3664 (N_3664,In_70,In_1233);
xor U3665 (N_3665,In_1196,In_17);
xnor U3666 (N_3666,In_397,In_1103);
nor U3667 (N_3667,In_875,In_1353);
xor U3668 (N_3668,In_980,In_1183);
nand U3669 (N_3669,In_144,In_302);
nand U3670 (N_3670,In_242,In_404);
or U3671 (N_3671,In_1312,In_389);
and U3672 (N_3672,In_236,In_1295);
nor U3673 (N_3673,In_326,In_142);
or U3674 (N_3674,In_1142,In_1111);
nand U3675 (N_3675,In_627,In_767);
or U3676 (N_3676,In_1241,In_528);
and U3677 (N_3677,In_158,In_1213);
nor U3678 (N_3678,In_1031,In_817);
or U3679 (N_3679,In_272,In_488);
and U3680 (N_3680,In_322,In_316);
nand U3681 (N_3681,In_342,In_762);
or U3682 (N_3682,In_252,In_1491);
or U3683 (N_3683,In_1105,In_720);
and U3684 (N_3684,In_1206,In_673);
or U3685 (N_3685,In_105,In_1304);
nand U3686 (N_3686,In_847,In_1430);
nor U3687 (N_3687,In_1479,In_459);
nand U3688 (N_3688,In_820,In_689);
or U3689 (N_3689,In_667,In_40);
or U3690 (N_3690,In_1210,In_1165);
or U3691 (N_3691,In_1497,In_1355);
and U3692 (N_3692,In_1045,In_1434);
and U3693 (N_3693,In_993,In_74);
nand U3694 (N_3694,In_827,In_161);
nand U3695 (N_3695,In_1134,In_939);
or U3696 (N_3696,In_612,In_1020);
or U3697 (N_3697,In_1465,In_1245);
nor U3698 (N_3698,In_1470,In_418);
nor U3699 (N_3699,In_1097,In_656);
nor U3700 (N_3700,In_996,In_190);
nor U3701 (N_3701,In_958,In_815);
and U3702 (N_3702,In_776,In_690);
and U3703 (N_3703,In_915,In_385);
xnor U3704 (N_3704,In_301,In_1425);
nor U3705 (N_3705,In_229,In_98);
nand U3706 (N_3706,In_711,In_457);
nor U3707 (N_3707,In_1345,In_176);
nor U3708 (N_3708,In_672,In_1034);
or U3709 (N_3709,In_911,In_415);
xnor U3710 (N_3710,In_1064,In_1482);
nand U3711 (N_3711,In_830,In_662);
nor U3712 (N_3712,In_1199,In_377);
or U3713 (N_3713,In_174,In_1304);
or U3714 (N_3714,In_1116,In_1487);
or U3715 (N_3715,In_1472,In_642);
nand U3716 (N_3716,In_778,In_20);
nor U3717 (N_3717,In_874,In_471);
nor U3718 (N_3718,In_890,In_1459);
and U3719 (N_3719,In_1222,In_693);
or U3720 (N_3720,In_719,In_928);
xnor U3721 (N_3721,In_941,In_223);
and U3722 (N_3722,In_156,In_1361);
or U3723 (N_3723,In_686,In_333);
or U3724 (N_3724,In_580,In_758);
xnor U3725 (N_3725,In_527,In_62);
and U3726 (N_3726,In_1039,In_600);
nand U3727 (N_3727,In_814,In_411);
and U3728 (N_3728,In_764,In_973);
xnor U3729 (N_3729,In_1365,In_3);
xor U3730 (N_3730,In_1187,In_1181);
or U3731 (N_3731,In_594,In_744);
nor U3732 (N_3732,In_548,In_186);
nor U3733 (N_3733,In_323,In_846);
and U3734 (N_3734,In_1355,In_661);
or U3735 (N_3735,In_1437,In_747);
nor U3736 (N_3736,In_738,In_419);
and U3737 (N_3737,In_903,In_390);
xor U3738 (N_3738,In_125,In_83);
xnor U3739 (N_3739,In_576,In_1173);
nor U3740 (N_3740,In_196,In_1358);
or U3741 (N_3741,In_328,In_909);
xnor U3742 (N_3742,In_937,In_670);
and U3743 (N_3743,In_619,In_344);
or U3744 (N_3744,In_774,In_952);
xor U3745 (N_3745,In_792,In_257);
or U3746 (N_3746,In_467,In_993);
xnor U3747 (N_3747,In_43,In_1479);
xor U3748 (N_3748,In_12,In_983);
nor U3749 (N_3749,In_769,In_280);
xnor U3750 (N_3750,In_1041,In_631);
and U3751 (N_3751,In_1123,In_1239);
xnor U3752 (N_3752,In_1060,In_805);
or U3753 (N_3753,In_434,In_377);
nor U3754 (N_3754,In_415,In_423);
xor U3755 (N_3755,In_1426,In_640);
nor U3756 (N_3756,In_834,In_510);
and U3757 (N_3757,In_485,In_141);
and U3758 (N_3758,In_464,In_1287);
or U3759 (N_3759,In_640,In_564);
xnor U3760 (N_3760,In_1261,In_1026);
or U3761 (N_3761,In_1254,In_24);
or U3762 (N_3762,In_1010,In_317);
and U3763 (N_3763,In_782,In_267);
nor U3764 (N_3764,In_474,In_141);
nor U3765 (N_3765,In_405,In_424);
and U3766 (N_3766,In_448,In_1384);
or U3767 (N_3767,In_1253,In_892);
nor U3768 (N_3768,In_582,In_476);
nand U3769 (N_3769,In_7,In_896);
and U3770 (N_3770,In_751,In_1225);
nor U3771 (N_3771,In_439,In_1370);
nor U3772 (N_3772,In_1444,In_1390);
nand U3773 (N_3773,In_128,In_1298);
and U3774 (N_3774,In_127,In_84);
nand U3775 (N_3775,In_941,In_269);
or U3776 (N_3776,In_664,In_207);
nor U3777 (N_3777,In_691,In_57);
nand U3778 (N_3778,In_253,In_473);
and U3779 (N_3779,In_778,In_467);
nor U3780 (N_3780,In_1271,In_870);
nand U3781 (N_3781,In_1415,In_1006);
nor U3782 (N_3782,In_321,In_731);
nand U3783 (N_3783,In_84,In_1330);
nor U3784 (N_3784,In_694,In_730);
nor U3785 (N_3785,In_1266,In_1058);
or U3786 (N_3786,In_1429,In_249);
nand U3787 (N_3787,In_431,In_984);
xor U3788 (N_3788,In_591,In_915);
and U3789 (N_3789,In_198,In_406);
or U3790 (N_3790,In_369,In_884);
nand U3791 (N_3791,In_861,In_1072);
xor U3792 (N_3792,In_861,In_583);
xnor U3793 (N_3793,In_1166,In_1072);
or U3794 (N_3794,In_93,In_1096);
or U3795 (N_3795,In_1368,In_887);
nor U3796 (N_3796,In_87,In_707);
or U3797 (N_3797,In_138,In_1491);
nor U3798 (N_3798,In_976,In_755);
nor U3799 (N_3799,In_473,In_633);
nand U3800 (N_3800,In_1148,In_816);
xor U3801 (N_3801,In_1086,In_371);
nand U3802 (N_3802,In_463,In_740);
nor U3803 (N_3803,In_352,In_254);
xor U3804 (N_3804,In_774,In_541);
xnor U3805 (N_3805,In_1370,In_1483);
or U3806 (N_3806,In_1266,In_682);
xor U3807 (N_3807,In_516,In_366);
nand U3808 (N_3808,In_35,In_455);
xor U3809 (N_3809,In_367,In_475);
nor U3810 (N_3810,In_1026,In_751);
nor U3811 (N_3811,In_1412,In_162);
or U3812 (N_3812,In_170,In_107);
and U3813 (N_3813,In_1164,In_509);
and U3814 (N_3814,In_628,In_543);
or U3815 (N_3815,In_1285,In_1457);
nor U3816 (N_3816,In_452,In_707);
nor U3817 (N_3817,In_1100,In_582);
nand U3818 (N_3818,In_53,In_479);
nor U3819 (N_3819,In_1051,In_24);
or U3820 (N_3820,In_722,In_1213);
or U3821 (N_3821,In_814,In_420);
or U3822 (N_3822,In_680,In_1390);
or U3823 (N_3823,In_402,In_1407);
nor U3824 (N_3824,In_260,In_1305);
and U3825 (N_3825,In_869,In_539);
and U3826 (N_3826,In_787,In_843);
nor U3827 (N_3827,In_374,In_319);
or U3828 (N_3828,In_1006,In_72);
and U3829 (N_3829,In_1381,In_1128);
nand U3830 (N_3830,In_1426,In_134);
and U3831 (N_3831,In_188,In_1337);
nand U3832 (N_3832,In_1093,In_1024);
and U3833 (N_3833,In_401,In_332);
nand U3834 (N_3834,In_19,In_252);
xnor U3835 (N_3835,In_400,In_756);
nand U3836 (N_3836,In_614,In_1274);
xnor U3837 (N_3837,In_951,In_1203);
nor U3838 (N_3838,In_109,In_1475);
or U3839 (N_3839,In_625,In_1027);
nor U3840 (N_3840,In_31,In_97);
xnor U3841 (N_3841,In_1188,In_197);
xor U3842 (N_3842,In_945,In_787);
nor U3843 (N_3843,In_1019,In_62);
xnor U3844 (N_3844,In_1238,In_1292);
or U3845 (N_3845,In_883,In_1069);
nor U3846 (N_3846,In_1276,In_790);
and U3847 (N_3847,In_830,In_164);
and U3848 (N_3848,In_1338,In_483);
nand U3849 (N_3849,In_769,In_1426);
or U3850 (N_3850,In_565,In_990);
nor U3851 (N_3851,In_831,In_587);
and U3852 (N_3852,In_1311,In_471);
and U3853 (N_3853,In_640,In_764);
or U3854 (N_3854,In_1233,In_955);
and U3855 (N_3855,In_338,In_1150);
or U3856 (N_3856,In_14,In_553);
nor U3857 (N_3857,In_105,In_48);
nand U3858 (N_3858,In_714,In_1380);
nand U3859 (N_3859,In_1005,In_1483);
or U3860 (N_3860,In_1425,In_316);
or U3861 (N_3861,In_429,In_1002);
nor U3862 (N_3862,In_315,In_45);
or U3863 (N_3863,In_1325,In_1347);
xor U3864 (N_3864,In_668,In_77);
or U3865 (N_3865,In_1382,In_1449);
nor U3866 (N_3866,In_745,In_785);
nand U3867 (N_3867,In_267,In_648);
nor U3868 (N_3868,In_1097,In_210);
nand U3869 (N_3869,In_1041,In_692);
and U3870 (N_3870,In_1281,In_435);
or U3871 (N_3871,In_536,In_1293);
nor U3872 (N_3872,In_663,In_1340);
xor U3873 (N_3873,In_1089,In_747);
or U3874 (N_3874,In_912,In_48);
nand U3875 (N_3875,In_919,In_483);
xnor U3876 (N_3876,In_1014,In_637);
or U3877 (N_3877,In_25,In_302);
nor U3878 (N_3878,In_602,In_845);
and U3879 (N_3879,In_95,In_417);
nor U3880 (N_3880,In_413,In_905);
nor U3881 (N_3881,In_901,In_394);
and U3882 (N_3882,In_513,In_925);
nand U3883 (N_3883,In_843,In_551);
or U3884 (N_3884,In_1404,In_381);
nand U3885 (N_3885,In_1257,In_285);
nand U3886 (N_3886,In_1495,In_322);
nor U3887 (N_3887,In_1301,In_1234);
nor U3888 (N_3888,In_1407,In_108);
nand U3889 (N_3889,In_1165,In_756);
or U3890 (N_3890,In_970,In_771);
nor U3891 (N_3891,In_150,In_113);
nor U3892 (N_3892,In_87,In_1075);
nor U3893 (N_3893,In_507,In_1353);
xor U3894 (N_3894,In_1063,In_339);
nand U3895 (N_3895,In_380,In_73);
nand U3896 (N_3896,In_497,In_756);
and U3897 (N_3897,In_292,In_217);
and U3898 (N_3898,In_1005,In_1094);
or U3899 (N_3899,In_1185,In_726);
and U3900 (N_3900,In_45,In_972);
nor U3901 (N_3901,In_708,In_1146);
xor U3902 (N_3902,In_1099,In_1449);
and U3903 (N_3903,In_1051,In_1079);
and U3904 (N_3904,In_47,In_1033);
and U3905 (N_3905,In_1412,In_638);
nand U3906 (N_3906,In_1307,In_655);
or U3907 (N_3907,In_315,In_610);
nand U3908 (N_3908,In_196,In_282);
or U3909 (N_3909,In_1096,In_1336);
nor U3910 (N_3910,In_97,In_1465);
nand U3911 (N_3911,In_902,In_1195);
xnor U3912 (N_3912,In_185,In_366);
nand U3913 (N_3913,In_894,In_222);
xor U3914 (N_3914,In_1064,In_965);
nand U3915 (N_3915,In_586,In_48);
nand U3916 (N_3916,In_65,In_1060);
or U3917 (N_3917,In_584,In_749);
xnor U3918 (N_3918,In_547,In_637);
or U3919 (N_3919,In_1290,In_1302);
and U3920 (N_3920,In_1422,In_255);
nor U3921 (N_3921,In_1161,In_521);
nor U3922 (N_3922,In_1369,In_609);
nand U3923 (N_3923,In_1310,In_13);
or U3924 (N_3924,In_359,In_1170);
xnor U3925 (N_3925,In_171,In_538);
nor U3926 (N_3926,In_35,In_838);
or U3927 (N_3927,In_791,In_588);
nand U3928 (N_3928,In_423,In_226);
or U3929 (N_3929,In_22,In_1392);
or U3930 (N_3930,In_917,In_739);
and U3931 (N_3931,In_1128,In_1186);
nor U3932 (N_3932,In_1287,In_327);
nor U3933 (N_3933,In_986,In_210);
or U3934 (N_3934,In_1110,In_229);
nand U3935 (N_3935,In_621,In_448);
xor U3936 (N_3936,In_1102,In_424);
nand U3937 (N_3937,In_4,In_702);
nand U3938 (N_3938,In_1495,In_693);
or U3939 (N_3939,In_1483,In_345);
xnor U3940 (N_3940,In_44,In_1070);
and U3941 (N_3941,In_1057,In_1308);
nand U3942 (N_3942,In_130,In_972);
and U3943 (N_3943,In_1143,In_773);
nor U3944 (N_3944,In_744,In_1422);
xor U3945 (N_3945,In_617,In_742);
nand U3946 (N_3946,In_107,In_1043);
and U3947 (N_3947,In_1038,In_678);
or U3948 (N_3948,In_1304,In_1361);
and U3949 (N_3949,In_877,In_56);
nor U3950 (N_3950,In_1240,In_464);
and U3951 (N_3951,In_282,In_420);
or U3952 (N_3952,In_7,In_10);
xnor U3953 (N_3953,In_1196,In_894);
and U3954 (N_3954,In_119,In_664);
xnor U3955 (N_3955,In_538,In_1119);
xnor U3956 (N_3956,In_1435,In_1168);
or U3957 (N_3957,In_1175,In_1499);
and U3958 (N_3958,In_1017,In_674);
xnor U3959 (N_3959,In_878,In_508);
or U3960 (N_3960,In_830,In_345);
xnor U3961 (N_3961,In_77,In_1312);
nor U3962 (N_3962,In_482,In_26);
xnor U3963 (N_3963,In_735,In_229);
xor U3964 (N_3964,In_1332,In_178);
and U3965 (N_3965,In_235,In_113);
and U3966 (N_3966,In_436,In_1101);
nor U3967 (N_3967,In_208,In_1280);
and U3968 (N_3968,In_648,In_598);
xnor U3969 (N_3969,In_1143,In_977);
xnor U3970 (N_3970,In_215,In_1061);
or U3971 (N_3971,In_354,In_836);
nor U3972 (N_3972,In_539,In_778);
nor U3973 (N_3973,In_130,In_1238);
and U3974 (N_3974,In_377,In_1223);
and U3975 (N_3975,In_782,In_123);
nand U3976 (N_3976,In_424,In_834);
nand U3977 (N_3977,In_1494,In_891);
nor U3978 (N_3978,In_1020,In_162);
nand U3979 (N_3979,In_524,In_1299);
xor U3980 (N_3980,In_38,In_845);
nand U3981 (N_3981,In_594,In_1370);
xnor U3982 (N_3982,In_986,In_793);
xor U3983 (N_3983,In_844,In_1089);
nand U3984 (N_3984,In_1103,In_1226);
nor U3985 (N_3985,In_928,In_781);
nand U3986 (N_3986,In_254,In_39);
nor U3987 (N_3987,In_712,In_135);
nand U3988 (N_3988,In_1041,In_17);
or U3989 (N_3989,In_1240,In_71);
and U3990 (N_3990,In_509,In_702);
or U3991 (N_3991,In_802,In_814);
or U3992 (N_3992,In_280,In_337);
nor U3993 (N_3993,In_1459,In_1406);
nand U3994 (N_3994,In_1000,In_305);
and U3995 (N_3995,In_629,In_1290);
xor U3996 (N_3996,In_151,In_386);
nor U3997 (N_3997,In_1103,In_1232);
and U3998 (N_3998,In_341,In_707);
xnor U3999 (N_3999,In_322,In_37);
nand U4000 (N_4000,In_417,In_454);
and U4001 (N_4001,In_499,In_530);
nor U4002 (N_4002,In_726,In_117);
nand U4003 (N_4003,In_213,In_995);
xnor U4004 (N_4004,In_294,In_374);
nor U4005 (N_4005,In_1184,In_1398);
nand U4006 (N_4006,In_405,In_810);
nand U4007 (N_4007,In_626,In_1314);
nor U4008 (N_4008,In_824,In_1352);
nor U4009 (N_4009,In_1450,In_741);
xor U4010 (N_4010,In_97,In_723);
xnor U4011 (N_4011,In_1079,In_1098);
or U4012 (N_4012,In_300,In_1364);
and U4013 (N_4013,In_1216,In_439);
nor U4014 (N_4014,In_1387,In_444);
or U4015 (N_4015,In_1499,In_284);
and U4016 (N_4016,In_770,In_732);
xnor U4017 (N_4017,In_357,In_684);
or U4018 (N_4018,In_1225,In_1437);
nor U4019 (N_4019,In_87,In_357);
nor U4020 (N_4020,In_834,In_176);
nand U4021 (N_4021,In_869,In_533);
nand U4022 (N_4022,In_451,In_630);
nand U4023 (N_4023,In_1163,In_949);
xor U4024 (N_4024,In_97,In_333);
nor U4025 (N_4025,In_366,In_186);
nor U4026 (N_4026,In_791,In_1313);
and U4027 (N_4027,In_1030,In_774);
xnor U4028 (N_4028,In_1359,In_1367);
or U4029 (N_4029,In_708,In_811);
or U4030 (N_4030,In_1414,In_132);
nor U4031 (N_4031,In_799,In_819);
and U4032 (N_4032,In_311,In_1165);
nor U4033 (N_4033,In_1270,In_904);
or U4034 (N_4034,In_765,In_289);
nand U4035 (N_4035,In_578,In_710);
xnor U4036 (N_4036,In_1258,In_1033);
or U4037 (N_4037,In_1293,In_1010);
nor U4038 (N_4038,In_912,In_215);
or U4039 (N_4039,In_1018,In_1256);
nor U4040 (N_4040,In_240,In_1254);
nand U4041 (N_4041,In_1437,In_809);
nor U4042 (N_4042,In_206,In_483);
nand U4043 (N_4043,In_39,In_241);
or U4044 (N_4044,In_1424,In_1311);
xor U4045 (N_4045,In_79,In_826);
nand U4046 (N_4046,In_944,In_1488);
or U4047 (N_4047,In_664,In_633);
and U4048 (N_4048,In_596,In_390);
nand U4049 (N_4049,In_130,In_349);
or U4050 (N_4050,In_1015,In_1107);
or U4051 (N_4051,In_1427,In_439);
and U4052 (N_4052,In_250,In_552);
nor U4053 (N_4053,In_1456,In_223);
nor U4054 (N_4054,In_1267,In_778);
xor U4055 (N_4055,In_231,In_223);
nor U4056 (N_4056,In_1319,In_970);
xnor U4057 (N_4057,In_1347,In_753);
nand U4058 (N_4058,In_795,In_1078);
xor U4059 (N_4059,In_1404,In_207);
nor U4060 (N_4060,In_724,In_367);
nand U4061 (N_4061,In_1433,In_403);
nor U4062 (N_4062,In_996,In_558);
xnor U4063 (N_4063,In_833,In_900);
xor U4064 (N_4064,In_439,In_1261);
nor U4065 (N_4065,In_6,In_133);
nor U4066 (N_4066,In_1101,In_1458);
and U4067 (N_4067,In_1279,In_274);
or U4068 (N_4068,In_571,In_1189);
or U4069 (N_4069,In_1036,In_724);
nand U4070 (N_4070,In_1126,In_1094);
nand U4071 (N_4071,In_1415,In_508);
nor U4072 (N_4072,In_517,In_859);
or U4073 (N_4073,In_1453,In_1253);
nor U4074 (N_4074,In_248,In_14);
nor U4075 (N_4075,In_162,In_324);
or U4076 (N_4076,In_876,In_267);
nor U4077 (N_4077,In_422,In_1346);
or U4078 (N_4078,In_685,In_1276);
nor U4079 (N_4079,In_845,In_730);
nor U4080 (N_4080,In_368,In_1252);
nand U4081 (N_4081,In_1335,In_135);
nand U4082 (N_4082,In_636,In_276);
nor U4083 (N_4083,In_372,In_648);
nand U4084 (N_4084,In_39,In_893);
xnor U4085 (N_4085,In_666,In_44);
xor U4086 (N_4086,In_181,In_1455);
xor U4087 (N_4087,In_935,In_1085);
xnor U4088 (N_4088,In_1106,In_1467);
nor U4089 (N_4089,In_684,In_1482);
nor U4090 (N_4090,In_1156,In_770);
nor U4091 (N_4091,In_482,In_448);
nor U4092 (N_4092,In_252,In_85);
nand U4093 (N_4093,In_1316,In_583);
and U4094 (N_4094,In_66,In_1361);
nor U4095 (N_4095,In_84,In_1460);
or U4096 (N_4096,In_35,In_373);
and U4097 (N_4097,In_108,In_1314);
and U4098 (N_4098,In_1371,In_1373);
nor U4099 (N_4099,In_673,In_1441);
nor U4100 (N_4100,In_1191,In_1155);
nand U4101 (N_4101,In_818,In_1187);
xnor U4102 (N_4102,In_1171,In_451);
or U4103 (N_4103,In_234,In_193);
or U4104 (N_4104,In_278,In_376);
xnor U4105 (N_4105,In_1157,In_878);
nor U4106 (N_4106,In_101,In_223);
nand U4107 (N_4107,In_1001,In_405);
or U4108 (N_4108,In_809,In_766);
nand U4109 (N_4109,In_497,In_1224);
or U4110 (N_4110,In_830,In_236);
or U4111 (N_4111,In_1377,In_319);
or U4112 (N_4112,In_1144,In_1234);
or U4113 (N_4113,In_700,In_1343);
xnor U4114 (N_4114,In_675,In_475);
nor U4115 (N_4115,In_1386,In_770);
xor U4116 (N_4116,In_311,In_59);
or U4117 (N_4117,In_169,In_864);
xor U4118 (N_4118,In_679,In_495);
nand U4119 (N_4119,In_349,In_751);
nand U4120 (N_4120,In_583,In_1115);
nor U4121 (N_4121,In_730,In_761);
xnor U4122 (N_4122,In_268,In_67);
nand U4123 (N_4123,In_1421,In_666);
nand U4124 (N_4124,In_591,In_351);
nor U4125 (N_4125,In_573,In_1212);
and U4126 (N_4126,In_928,In_1066);
nand U4127 (N_4127,In_1175,In_124);
xor U4128 (N_4128,In_1429,In_6);
or U4129 (N_4129,In_1498,In_532);
and U4130 (N_4130,In_625,In_1056);
xor U4131 (N_4131,In_1328,In_945);
and U4132 (N_4132,In_943,In_1260);
nor U4133 (N_4133,In_1029,In_1436);
nand U4134 (N_4134,In_1457,In_1250);
and U4135 (N_4135,In_1394,In_79);
nor U4136 (N_4136,In_1191,In_87);
or U4137 (N_4137,In_1327,In_223);
nand U4138 (N_4138,In_619,In_173);
xnor U4139 (N_4139,In_184,In_49);
xnor U4140 (N_4140,In_728,In_1288);
xnor U4141 (N_4141,In_1407,In_787);
and U4142 (N_4142,In_609,In_581);
xnor U4143 (N_4143,In_76,In_1025);
and U4144 (N_4144,In_277,In_542);
or U4145 (N_4145,In_23,In_1236);
nand U4146 (N_4146,In_805,In_1441);
or U4147 (N_4147,In_623,In_758);
nand U4148 (N_4148,In_949,In_1330);
nor U4149 (N_4149,In_656,In_432);
and U4150 (N_4150,In_690,In_1058);
and U4151 (N_4151,In_1415,In_1374);
nand U4152 (N_4152,In_52,In_31);
xnor U4153 (N_4153,In_178,In_106);
nor U4154 (N_4154,In_311,In_12);
nor U4155 (N_4155,In_634,In_346);
nand U4156 (N_4156,In_708,In_1431);
nor U4157 (N_4157,In_165,In_540);
and U4158 (N_4158,In_548,In_223);
and U4159 (N_4159,In_1039,In_1189);
and U4160 (N_4160,In_1385,In_1171);
nand U4161 (N_4161,In_3,In_105);
nor U4162 (N_4162,In_1361,In_455);
nor U4163 (N_4163,In_354,In_454);
and U4164 (N_4164,In_909,In_878);
or U4165 (N_4165,In_292,In_552);
nor U4166 (N_4166,In_646,In_813);
nor U4167 (N_4167,In_1397,In_390);
nor U4168 (N_4168,In_820,In_101);
or U4169 (N_4169,In_330,In_733);
xnor U4170 (N_4170,In_954,In_1390);
xor U4171 (N_4171,In_1406,In_554);
or U4172 (N_4172,In_1315,In_827);
nor U4173 (N_4173,In_928,In_1346);
xor U4174 (N_4174,In_996,In_670);
xor U4175 (N_4175,In_786,In_490);
or U4176 (N_4176,In_638,In_167);
and U4177 (N_4177,In_1279,In_1011);
nor U4178 (N_4178,In_1472,In_86);
nand U4179 (N_4179,In_387,In_914);
nor U4180 (N_4180,In_843,In_124);
and U4181 (N_4181,In_1006,In_318);
nand U4182 (N_4182,In_491,In_767);
nand U4183 (N_4183,In_494,In_709);
or U4184 (N_4184,In_1174,In_514);
nor U4185 (N_4185,In_1054,In_36);
and U4186 (N_4186,In_300,In_227);
nand U4187 (N_4187,In_1458,In_1287);
or U4188 (N_4188,In_1420,In_1137);
and U4189 (N_4189,In_596,In_292);
nand U4190 (N_4190,In_494,In_696);
nor U4191 (N_4191,In_1064,In_1338);
xnor U4192 (N_4192,In_995,In_430);
nand U4193 (N_4193,In_305,In_301);
nand U4194 (N_4194,In_707,In_1370);
nor U4195 (N_4195,In_739,In_1249);
nor U4196 (N_4196,In_1339,In_1093);
or U4197 (N_4197,In_509,In_129);
nor U4198 (N_4198,In_567,In_63);
nand U4199 (N_4199,In_998,In_678);
nand U4200 (N_4200,In_994,In_1100);
or U4201 (N_4201,In_112,In_556);
or U4202 (N_4202,In_1365,In_1484);
and U4203 (N_4203,In_1444,In_121);
or U4204 (N_4204,In_764,In_282);
nand U4205 (N_4205,In_339,In_77);
nand U4206 (N_4206,In_708,In_1104);
or U4207 (N_4207,In_1417,In_237);
nand U4208 (N_4208,In_659,In_667);
or U4209 (N_4209,In_377,In_996);
nor U4210 (N_4210,In_623,In_359);
nor U4211 (N_4211,In_461,In_1157);
and U4212 (N_4212,In_1494,In_787);
xnor U4213 (N_4213,In_1085,In_1211);
nor U4214 (N_4214,In_460,In_1310);
nand U4215 (N_4215,In_1159,In_337);
nand U4216 (N_4216,In_1091,In_435);
or U4217 (N_4217,In_811,In_346);
nand U4218 (N_4218,In_1492,In_593);
and U4219 (N_4219,In_924,In_637);
and U4220 (N_4220,In_1267,In_508);
nor U4221 (N_4221,In_324,In_108);
or U4222 (N_4222,In_406,In_1031);
nand U4223 (N_4223,In_203,In_1006);
and U4224 (N_4224,In_83,In_1334);
xnor U4225 (N_4225,In_1300,In_417);
nand U4226 (N_4226,In_1336,In_3);
and U4227 (N_4227,In_330,In_494);
and U4228 (N_4228,In_22,In_788);
or U4229 (N_4229,In_1114,In_281);
nor U4230 (N_4230,In_1059,In_827);
and U4231 (N_4231,In_1376,In_1172);
xor U4232 (N_4232,In_1317,In_12);
and U4233 (N_4233,In_481,In_276);
xnor U4234 (N_4234,In_1377,In_32);
xnor U4235 (N_4235,In_1144,In_1487);
xnor U4236 (N_4236,In_1157,In_43);
xnor U4237 (N_4237,In_1467,In_269);
nor U4238 (N_4238,In_1419,In_9);
or U4239 (N_4239,In_1279,In_608);
or U4240 (N_4240,In_280,In_903);
nor U4241 (N_4241,In_336,In_404);
and U4242 (N_4242,In_372,In_1159);
or U4243 (N_4243,In_1219,In_375);
xnor U4244 (N_4244,In_529,In_1053);
xnor U4245 (N_4245,In_340,In_437);
nor U4246 (N_4246,In_855,In_86);
and U4247 (N_4247,In_186,In_1157);
or U4248 (N_4248,In_46,In_472);
nor U4249 (N_4249,In_129,In_1071);
xnor U4250 (N_4250,In_1276,In_1448);
xor U4251 (N_4251,In_721,In_421);
or U4252 (N_4252,In_997,In_828);
nor U4253 (N_4253,In_961,In_1108);
nor U4254 (N_4254,In_280,In_1292);
or U4255 (N_4255,In_203,In_1202);
nor U4256 (N_4256,In_931,In_812);
or U4257 (N_4257,In_916,In_0);
xnor U4258 (N_4258,In_1298,In_705);
and U4259 (N_4259,In_568,In_48);
and U4260 (N_4260,In_16,In_1235);
xnor U4261 (N_4261,In_1425,In_868);
xor U4262 (N_4262,In_118,In_1445);
and U4263 (N_4263,In_945,In_1052);
nor U4264 (N_4264,In_1173,In_1419);
xnor U4265 (N_4265,In_959,In_65);
xnor U4266 (N_4266,In_638,In_80);
and U4267 (N_4267,In_870,In_537);
nand U4268 (N_4268,In_1120,In_891);
xor U4269 (N_4269,In_1437,In_490);
nand U4270 (N_4270,In_920,In_223);
nand U4271 (N_4271,In_220,In_1134);
nor U4272 (N_4272,In_352,In_299);
nand U4273 (N_4273,In_735,In_505);
nand U4274 (N_4274,In_692,In_892);
or U4275 (N_4275,In_165,In_652);
xnor U4276 (N_4276,In_1272,In_875);
and U4277 (N_4277,In_1158,In_1366);
xnor U4278 (N_4278,In_393,In_185);
nand U4279 (N_4279,In_978,In_937);
nand U4280 (N_4280,In_955,In_450);
nor U4281 (N_4281,In_61,In_146);
xnor U4282 (N_4282,In_1212,In_1062);
nor U4283 (N_4283,In_97,In_68);
or U4284 (N_4284,In_538,In_138);
xor U4285 (N_4285,In_1249,In_939);
nor U4286 (N_4286,In_1402,In_1179);
or U4287 (N_4287,In_825,In_1140);
xor U4288 (N_4288,In_108,In_50);
or U4289 (N_4289,In_216,In_1301);
or U4290 (N_4290,In_415,In_169);
xnor U4291 (N_4291,In_1138,In_454);
xnor U4292 (N_4292,In_1393,In_1061);
nand U4293 (N_4293,In_1152,In_342);
nand U4294 (N_4294,In_195,In_1111);
and U4295 (N_4295,In_648,In_276);
nor U4296 (N_4296,In_218,In_342);
nand U4297 (N_4297,In_320,In_655);
and U4298 (N_4298,In_446,In_306);
or U4299 (N_4299,In_1165,In_167);
nand U4300 (N_4300,In_849,In_458);
nand U4301 (N_4301,In_332,In_1123);
or U4302 (N_4302,In_160,In_682);
and U4303 (N_4303,In_1001,In_533);
nand U4304 (N_4304,In_187,In_150);
or U4305 (N_4305,In_662,In_585);
or U4306 (N_4306,In_101,In_1330);
nor U4307 (N_4307,In_654,In_82);
xnor U4308 (N_4308,In_827,In_183);
or U4309 (N_4309,In_667,In_843);
xnor U4310 (N_4310,In_836,In_890);
and U4311 (N_4311,In_621,In_1328);
nand U4312 (N_4312,In_1403,In_999);
xnor U4313 (N_4313,In_644,In_1208);
or U4314 (N_4314,In_1216,In_1438);
nand U4315 (N_4315,In_529,In_714);
or U4316 (N_4316,In_170,In_1251);
or U4317 (N_4317,In_1153,In_1370);
or U4318 (N_4318,In_1435,In_580);
and U4319 (N_4319,In_1071,In_41);
and U4320 (N_4320,In_1068,In_219);
nand U4321 (N_4321,In_1365,In_1094);
and U4322 (N_4322,In_360,In_1098);
or U4323 (N_4323,In_686,In_499);
and U4324 (N_4324,In_255,In_1276);
nand U4325 (N_4325,In_115,In_234);
and U4326 (N_4326,In_1038,In_860);
nor U4327 (N_4327,In_1382,In_378);
nor U4328 (N_4328,In_531,In_187);
and U4329 (N_4329,In_1336,In_228);
xnor U4330 (N_4330,In_477,In_488);
or U4331 (N_4331,In_79,In_529);
nor U4332 (N_4332,In_856,In_1126);
nand U4333 (N_4333,In_422,In_265);
and U4334 (N_4334,In_71,In_378);
xor U4335 (N_4335,In_763,In_455);
or U4336 (N_4336,In_786,In_11);
nand U4337 (N_4337,In_32,In_68);
nor U4338 (N_4338,In_522,In_489);
nor U4339 (N_4339,In_1017,In_991);
xnor U4340 (N_4340,In_491,In_326);
or U4341 (N_4341,In_976,In_812);
and U4342 (N_4342,In_410,In_335);
nand U4343 (N_4343,In_170,In_601);
and U4344 (N_4344,In_734,In_88);
and U4345 (N_4345,In_289,In_1462);
nor U4346 (N_4346,In_1323,In_327);
and U4347 (N_4347,In_975,In_1243);
and U4348 (N_4348,In_370,In_440);
nand U4349 (N_4349,In_850,In_755);
nor U4350 (N_4350,In_713,In_366);
nor U4351 (N_4351,In_49,In_778);
nor U4352 (N_4352,In_1014,In_670);
and U4353 (N_4353,In_1015,In_186);
nand U4354 (N_4354,In_325,In_1065);
xor U4355 (N_4355,In_637,In_123);
xnor U4356 (N_4356,In_647,In_1360);
or U4357 (N_4357,In_442,In_1401);
xnor U4358 (N_4358,In_206,In_418);
and U4359 (N_4359,In_1148,In_64);
nand U4360 (N_4360,In_855,In_442);
nand U4361 (N_4361,In_106,In_1221);
and U4362 (N_4362,In_1005,In_1240);
or U4363 (N_4363,In_318,In_61);
or U4364 (N_4364,In_230,In_1313);
or U4365 (N_4365,In_1164,In_430);
and U4366 (N_4366,In_667,In_1386);
xnor U4367 (N_4367,In_852,In_1025);
or U4368 (N_4368,In_791,In_960);
nand U4369 (N_4369,In_1008,In_767);
nor U4370 (N_4370,In_704,In_818);
nor U4371 (N_4371,In_969,In_255);
and U4372 (N_4372,In_911,In_11);
or U4373 (N_4373,In_38,In_1466);
xnor U4374 (N_4374,In_1466,In_261);
nand U4375 (N_4375,In_257,In_1357);
nor U4376 (N_4376,In_1021,In_150);
nor U4377 (N_4377,In_1375,In_918);
and U4378 (N_4378,In_563,In_1163);
nand U4379 (N_4379,In_231,In_1185);
xor U4380 (N_4380,In_22,In_62);
or U4381 (N_4381,In_842,In_1301);
or U4382 (N_4382,In_241,In_173);
xnor U4383 (N_4383,In_1422,In_1332);
nand U4384 (N_4384,In_1378,In_101);
nor U4385 (N_4385,In_1223,In_1182);
nand U4386 (N_4386,In_367,In_828);
and U4387 (N_4387,In_175,In_380);
or U4388 (N_4388,In_1395,In_999);
or U4389 (N_4389,In_1492,In_830);
nor U4390 (N_4390,In_938,In_1461);
and U4391 (N_4391,In_1392,In_1393);
nor U4392 (N_4392,In_175,In_452);
xnor U4393 (N_4393,In_152,In_1443);
xnor U4394 (N_4394,In_758,In_659);
or U4395 (N_4395,In_862,In_344);
or U4396 (N_4396,In_1261,In_158);
or U4397 (N_4397,In_891,In_480);
xor U4398 (N_4398,In_328,In_1386);
nor U4399 (N_4399,In_1266,In_697);
nor U4400 (N_4400,In_195,In_44);
xnor U4401 (N_4401,In_588,In_905);
xor U4402 (N_4402,In_1401,In_200);
and U4403 (N_4403,In_1024,In_805);
or U4404 (N_4404,In_137,In_335);
or U4405 (N_4405,In_776,In_1434);
and U4406 (N_4406,In_913,In_567);
and U4407 (N_4407,In_1019,In_1002);
and U4408 (N_4408,In_1064,In_165);
xor U4409 (N_4409,In_839,In_1183);
or U4410 (N_4410,In_667,In_717);
or U4411 (N_4411,In_943,In_1432);
xnor U4412 (N_4412,In_1056,In_478);
and U4413 (N_4413,In_1406,In_635);
nand U4414 (N_4414,In_374,In_1227);
xor U4415 (N_4415,In_670,In_176);
nand U4416 (N_4416,In_767,In_634);
xnor U4417 (N_4417,In_721,In_209);
and U4418 (N_4418,In_1355,In_291);
or U4419 (N_4419,In_873,In_1344);
nand U4420 (N_4420,In_643,In_1392);
or U4421 (N_4421,In_868,In_303);
or U4422 (N_4422,In_912,In_520);
nor U4423 (N_4423,In_38,In_409);
nor U4424 (N_4424,In_1056,In_502);
nor U4425 (N_4425,In_703,In_2);
xnor U4426 (N_4426,In_559,In_118);
and U4427 (N_4427,In_198,In_89);
xnor U4428 (N_4428,In_666,In_278);
nor U4429 (N_4429,In_1263,In_384);
nand U4430 (N_4430,In_1368,In_262);
and U4431 (N_4431,In_854,In_1162);
nor U4432 (N_4432,In_125,In_873);
nand U4433 (N_4433,In_801,In_1378);
and U4434 (N_4434,In_808,In_126);
and U4435 (N_4435,In_832,In_1229);
and U4436 (N_4436,In_285,In_1292);
xnor U4437 (N_4437,In_562,In_337);
nand U4438 (N_4438,In_935,In_881);
and U4439 (N_4439,In_1400,In_73);
nor U4440 (N_4440,In_831,In_237);
nand U4441 (N_4441,In_674,In_192);
nand U4442 (N_4442,In_714,In_1004);
and U4443 (N_4443,In_1236,In_914);
nand U4444 (N_4444,In_309,In_929);
or U4445 (N_4445,In_1423,In_1207);
xnor U4446 (N_4446,In_1315,In_897);
or U4447 (N_4447,In_364,In_390);
nor U4448 (N_4448,In_737,In_11);
or U4449 (N_4449,In_356,In_538);
and U4450 (N_4450,In_81,In_727);
nand U4451 (N_4451,In_392,In_182);
nor U4452 (N_4452,In_549,In_1209);
xor U4453 (N_4453,In_872,In_789);
and U4454 (N_4454,In_55,In_582);
xnor U4455 (N_4455,In_536,In_399);
xnor U4456 (N_4456,In_891,In_1047);
nor U4457 (N_4457,In_866,In_409);
nor U4458 (N_4458,In_432,In_107);
and U4459 (N_4459,In_12,In_607);
or U4460 (N_4460,In_88,In_220);
and U4461 (N_4461,In_586,In_1058);
or U4462 (N_4462,In_288,In_615);
xor U4463 (N_4463,In_515,In_603);
xor U4464 (N_4464,In_415,In_352);
and U4465 (N_4465,In_894,In_29);
and U4466 (N_4466,In_217,In_255);
or U4467 (N_4467,In_1140,In_1301);
nand U4468 (N_4468,In_1163,In_331);
nand U4469 (N_4469,In_1352,In_1391);
nand U4470 (N_4470,In_1298,In_349);
or U4471 (N_4471,In_1047,In_132);
and U4472 (N_4472,In_63,In_691);
xnor U4473 (N_4473,In_641,In_1227);
or U4474 (N_4474,In_468,In_29);
xor U4475 (N_4475,In_1346,In_1422);
and U4476 (N_4476,In_507,In_592);
and U4477 (N_4477,In_1348,In_223);
and U4478 (N_4478,In_1225,In_412);
xnor U4479 (N_4479,In_608,In_396);
or U4480 (N_4480,In_828,In_1432);
and U4481 (N_4481,In_761,In_643);
and U4482 (N_4482,In_258,In_757);
nand U4483 (N_4483,In_819,In_387);
and U4484 (N_4484,In_673,In_852);
nand U4485 (N_4485,In_998,In_1119);
or U4486 (N_4486,In_158,In_1370);
nor U4487 (N_4487,In_129,In_505);
nor U4488 (N_4488,In_1068,In_1012);
nor U4489 (N_4489,In_245,In_551);
nor U4490 (N_4490,In_976,In_1020);
nand U4491 (N_4491,In_393,In_321);
xor U4492 (N_4492,In_1174,In_369);
xor U4493 (N_4493,In_524,In_805);
and U4494 (N_4494,In_190,In_1261);
nand U4495 (N_4495,In_689,In_1220);
and U4496 (N_4496,In_650,In_862);
or U4497 (N_4497,In_488,In_713);
xor U4498 (N_4498,In_886,In_1308);
nor U4499 (N_4499,In_761,In_905);
nor U4500 (N_4500,In_1067,In_18);
nor U4501 (N_4501,In_695,In_87);
xnor U4502 (N_4502,In_772,In_1406);
or U4503 (N_4503,In_623,In_501);
or U4504 (N_4504,In_1385,In_511);
nand U4505 (N_4505,In_1192,In_1011);
nand U4506 (N_4506,In_195,In_263);
nand U4507 (N_4507,In_1013,In_765);
nor U4508 (N_4508,In_162,In_1176);
or U4509 (N_4509,In_473,In_598);
xor U4510 (N_4510,In_1069,In_1164);
nand U4511 (N_4511,In_1350,In_684);
nor U4512 (N_4512,In_1158,In_520);
or U4513 (N_4513,In_155,In_141);
or U4514 (N_4514,In_1182,In_771);
nor U4515 (N_4515,In_671,In_642);
xnor U4516 (N_4516,In_20,In_332);
or U4517 (N_4517,In_509,In_549);
xnor U4518 (N_4518,In_654,In_325);
and U4519 (N_4519,In_78,In_1217);
nor U4520 (N_4520,In_922,In_1491);
and U4521 (N_4521,In_427,In_996);
xnor U4522 (N_4522,In_814,In_1113);
nor U4523 (N_4523,In_856,In_946);
nor U4524 (N_4524,In_290,In_299);
or U4525 (N_4525,In_100,In_884);
and U4526 (N_4526,In_449,In_959);
xor U4527 (N_4527,In_1093,In_894);
nor U4528 (N_4528,In_884,In_799);
xor U4529 (N_4529,In_1402,In_778);
nor U4530 (N_4530,In_1167,In_838);
nand U4531 (N_4531,In_243,In_907);
nand U4532 (N_4532,In_897,In_684);
nor U4533 (N_4533,In_396,In_471);
and U4534 (N_4534,In_1402,In_1213);
and U4535 (N_4535,In_947,In_1317);
xor U4536 (N_4536,In_1224,In_348);
nor U4537 (N_4537,In_293,In_731);
or U4538 (N_4538,In_75,In_114);
xor U4539 (N_4539,In_1248,In_851);
and U4540 (N_4540,In_876,In_371);
nor U4541 (N_4541,In_975,In_765);
or U4542 (N_4542,In_843,In_346);
or U4543 (N_4543,In_1272,In_650);
and U4544 (N_4544,In_193,In_258);
or U4545 (N_4545,In_1050,In_6);
nand U4546 (N_4546,In_238,In_1104);
or U4547 (N_4547,In_603,In_802);
and U4548 (N_4548,In_473,In_604);
xor U4549 (N_4549,In_63,In_1373);
or U4550 (N_4550,In_782,In_89);
nand U4551 (N_4551,In_66,In_832);
nor U4552 (N_4552,In_1362,In_391);
nor U4553 (N_4553,In_1382,In_808);
nand U4554 (N_4554,In_362,In_683);
xnor U4555 (N_4555,In_1238,In_1202);
and U4556 (N_4556,In_314,In_560);
xnor U4557 (N_4557,In_608,In_18);
nor U4558 (N_4558,In_448,In_164);
nor U4559 (N_4559,In_668,In_792);
nor U4560 (N_4560,In_695,In_171);
and U4561 (N_4561,In_578,In_191);
xor U4562 (N_4562,In_61,In_260);
nand U4563 (N_4563,In_435,In_1361);
and U4564 (N_4564,In_1205,In_145);
or U4565 (N_4565,In_982,In_701);
xor U4566 (N_4566,In_1164,In_721);
and U4567 (N_4567,In_1372,In_715);
xor U4568 (N_4568,In_879,In_47);
and U4569 (N_4569,In_45,In_1221);
and U4570 (N_4570,In_744,In_698);
and U4571 (N_4571,In_1294,In_272);
or U4572 (N_4572,In_1467,In_975);
and U4573 (N_4573,In_605,In_1241);
nor U4574 (N_4574,In_500,In_177);
nand U4575 (N_4575,In_1392,In_18);
nand U4576 (N_4576,In_299,In_553);
or U4577 (N_4577,In_89,In_530);
or U4578 (N_4578,In_1126,In_156);
xnor U4579 (N_4579,In_821,In_1231);
and U4580 (N_4580,In_1454,In_1140);
nor U4581 (N_4581,In_684,In_1421);
or U4582 (N_4582,In_401,In_503);
and U4583 (N_4583,In_1298,In_462);
and U4584 (N_4584,In_1386,In_716);
nand U4585 (N_4585,In_230,In_1423);
nand U4586 (N_4586,In_1166,In_991);
nor U4587 (N_4587,In_1004,In_852);
and U4588 (N_4588,In_1009,In_1296);
xnor U4589 (N_4589,In_1125,In_709);
nor U4590 (N_4590,In_1248,In_144);
xnor U4591 (N_4591,In_39,In_986);
xor U4592 (N_4592,In_1248,In_560);
xnor U4593 (N_4593,In_1014,In_577);
nand U4594 (N_4594,In_1070,In_1107);
nand U4595 (N_4595,In_610,In_1431);
and U4596 (N_4596,In_799,In_713);
and U4597 (N_4597,In_133,In_865);
or U4598 (N_4598,In_1262,In_550);
and U4599 (N_4599,In_1349,In_924);
or U4600 (N_4600,In_801,In_262);
nor U4601 (N_4601,In_264,In_411);
nor U4602 (N_4602,In_146,In_1376);
nand U4603 (N_4603,In_215,In_866);
and U4604 (N_4604,In_100,In_342);
nor U4605 (N_4605,In_1246,In_374);
and U4606 (N_4606,In_1037,In_146);
nor U4607 (N_4607,In_1459,In_1119);
nor U4608 (N_4608,In_21,In_189);
xnor U4609 (N_4609,In_525,In_1169);
nand U4610 (N_4610,In_1314,In_606);
and U4611 (N_4611,In_529,In_291);
and U4612 (N_4612,In_98,In_763);
nand U4613 (N_4613,In_1195,In_447);
nand U4614 (N_4614,In_1343,In_92);
or U4615 (N_4615,In_1281,In_1188);
nand U4616 (N_4616,In_1464,In_354);
or U4617 (N_4617,In_1256,In_759);
or U4618 (N_4618,In_1052,In_464);
nand U4619 (N_4619,In_1196,In_1017);
or U4620 (N_4620,In_621,In_900);
and U4621 (N_4621,In_171,In_485);
and U4622 (N_4622,In_678,In_741);
or U4623 (N_4623,In_175,In_1311);
nand U4624 (N_4624,In_348,In_1028);
and U4625 (N_4625,In_327,In_964);
or U4626 (N_4626,In_871,In_270);
nand U4627 (N_4627,In_838,In_830);
and U4628 (N_4628,In_1033,In_163);
or U4629 (N_4629,In_1369,In_958);
and U4630 (N_4630,In_535,In_569);
xor U4631 (N_4631,In_556,In_1332);
nor U4632 (N_4632,In_737,In_910);
or U4633 (N_4633,In_1265,In_224);
nand U4634 (N_4634,In_1337,In_30);
xor U4635 (N_4635,In_293,In_1087);
and U4636 (N_4636,In_1416,In_1200);
xor U4637 (N_4637,In_1397,In_790);
nor U4638 (N_4638,In_1036,In_1215);
nor U4639 (N_4639,In_52,In_689);
nand U4640 (N_4640,In_1450,In_514);
nand U4641 (N_4641,In_762,In_229);
nand U4642 (N_4642,In_795,In_1246);
nand U4643 (N_4643,In_1159,In_609);
and U4644 (N_4644,In_88,In_70);
xnor U4645 (N_4645,In_99,In_1332);
and U4646 (N_4646,In_290,In_953);
xor U4647 (N_4647,In_1194,In_986);
xnor U4648 (N_4648,In_430,In_189);
nor U4649 (N_4649,In_282,In_824);
or U4650 (N_4650,In_799,In_985);
and U4651 (N_4651,In_1263,In_1333);
or U4652 (N_4652,In_612,In_1338);
and U4653 (N_4653,In_413,In_974);
xor U4654 (N_4654,In_233,In_593);
and U4655 (N_4655,In_1392,In_846);
nor U4656 (N_4656,In_428,In_56);
nand U4657 (N_4657,In_1012,In_227);
or U4658 (N_4658,In_7,In_1432);
nand U4659 (N_4659,In_295,In_130);
or U4660 (N_4660,In_1216,In_84);
and U4661 (N_4661,In_1257,In_369);
and U4662 (N_4662,In_1439,In_491);
nor U4663 (N_4663,In_354,In_962);
xnor U4664 (N_4664,In_1362,In_222);
nand U4665 (N_4665,In_1367,In_796);
nor U4666 (N_4666,In_805,In_1382);
and U4667 (N_4667,In_1260,In_989);
and U4668 (N_4668,In_865,In_1340);
nand U4669 (N_4669,In_1194,In_763);
nand U4670 (N_4670,In_142,In_1144);
or U4671 (N_4671,In_1245,In_1344);
xor U4672 (N_4672,In_986,In_1327);
nor U4673 (N_4673,In_1427,In_567);
xnor U4674 (N_4674,In_792,In_437);
or U4675 (N_4675,In_31,In_1320);
xor U4676 (N_4676,In_487,In_27);
nand U4677 (N_4677,In_748,In_20);
or U4678 (N_4678,In_419,In_970);
nor U4679 (N_4679,In_857,In_166);
nor U4680 (N_4680,In_36,In_376);
xnor U4681 (N_4681,In_1265,In_1428);
and U4682 (N_4682,In_28,In_891);
or U4683 (N_4683,In_239,In_401);
and U4684 (N_4684,In_1321,In_380);
xor U4685 (N_4685,In_475,In_749);
and U4686 (N_4686,In_1324,In_1101);
xor U4687 (N_4687,In_183,In_806);
or U4688 (N_4688,In_828,In_832);
and U4689 (N_4689,In_447,In_160);
nand U4690 (N_4690,In_1331,In_163);
nor U4691 (N_4691,In_631,In_1201);
or U4692 (N_4692,In_1437,In_244);
and U4693 (N_4693,In_1445,In_338);
nor U4694 (N_4694,In_424,In_400);
or U4695 (N_4695,In_821,In_985);
nor U4696 (N_4696,In_1441,In_498);
xor U4697 (N_4697,In_249,In_54);
nor U4698 (N_4698,In_498,In_770);
and U4699 (N_4699,In_510,In_301);
nor U4700 (N_4700,In_1081,In_1205);
nand U4701 (N_4701,In_787,In_988);
nand U4702 (N_4702,In_191,In_675);
nor U4703 (N_4703,In_1131,In_16);
nor U4704 (N_4704,In_600,In_563);
nor U4705 (N_4705,In_237,In_807);
or U4706 (N_4706,In_963,In_1093);
and U4707 (N_4707,In_1441,In_1447);
or U4708 (N_4708,In_1043,In_392);
and U4709 (N_4709,In_520,In_528);
nor U4710 (N_4710,In_743,In_94);
or U4711 (N_4711,In_546,In_1210);
nand U4712 (N_4712,In_263,In_273);
or U4713 (N_4713,In_363,In_686);
or U4714 (N_4714,In_164,In_251);
nand U4715 (N_4715,In_346,In_847);
nor U4716 (N_4716,In_725,In_1380);
xor U4717 (N_4717,In_110,In_761);
or U4718 (N_4718,In_749,In_59);
and U4719 (N_4719,In_1008,In_1381);
xor U4720 (N_4720,In_888,In_119);
nand U4721 (N_4721,In_582,In_799);
or U4722 (N_4722,In_138,In_65);
nor U4723 (N_4723,In_1329,In_949);
xnor U4724 (N_4724,In_860,In_366);
and U4725 (N_4725,In_637,In_988);
xnor U4726 (N_4726,In_149,In_1497);
nor U4727 (N_4727,In_1000,In_82);
or U4728 (N_4728,In_1105,In_1145);
nor U4729 (N_4729,In_817,In_1349);
nor U4730 (N_4730,In_1255,In_1198);
or U4731 (N_4731,In_1355,In_755);
and U4732 (N_4732,In_1459,In_532);
or U4733 (N_4733,In_1387,In_888);
nor U4734 (N_4734,In_1194,In_13);
nor U4735 (N_4735,In_975,In_1248);
nand U4736 (N_4736,In_170,In_913);
xor U4737 (N_4737,In_834,In_663);
nand U4738 (N_4738,In_1035,In_74);
nor U4739 (N_4739,In_1332,In_847);
or U4740 (N_4740,In_1471,In_746);
or U4741 (N_4741,In_1250,In_164);
and U4742 (N_4742,In_84,In_794);
xor U4743 (N_4743,In_1204,In_818);
or U4744 (N_4744,In_897,In_1048);
xnor U4745 (N_4745,In_944,In_420);
nor U4746 (N_4746,In_1086,In_836);
xor U4747 (N_4747,In_415,In_1185);
xnor U4748 (N_4748,In_1118,In_1440);
nand U4749 (N_4749,In_604,In_598);
or U4750 (N_4750,In_54,In_1199);
nand U4751 (N_4751,In_427,In_1347);
or U4752 (N_4752,In_655,In_713);
nand U4753 (N_4753,In_1060,In_225);
nor U4754 (N_4754,In_1458,In_617);
xor U4755 (N_4755,In_1495,In_557);
nor U4756 (N_4756,In_1,In_1239);
nor U4757 (N_4757,In_436,In_1039);
nand U4758 (N_4758,In_361,In_896);
nor U4759 (N_4759,In_1050,In_82);
nand U4760 (N_4760,In_300,In_102);
nor U4761 (N_4761,In_442,In_1351);
or U4762 (N_4762,In_1465,In_58);
nor U4763 (N_4763,In_1011,In_680);
and U4764 (N_4764,In_71,In_721);
or U4765 (N_4765,In_1063,In_841);
and U4766 (N_4766,In_1019,In_329);
nor U4767 (N_4767,In_972,In_765);
xor U4768 (N_4768,In_777,In_64);
or U4769 (N_4769,In_1107,In_1330);
xnor U4770 (N_4770,In_54,In_67);
nor U4771 (N_4771,In_300,In_538);
xor U4772 (N_4772,In_292,In_803);
and U4773 (N_4773,In_524,In_683);
or U4774 (N_4774,In_797,In_744);
nor U4775 (N_4775,In_955,In_41);
nand U4776 (N_4776,In_987,In_27);
nand U4777 (N_4777,In_473,In_905);
xor U4778 (N_4778,In_536,In_1215);
or U4779 (N_4779,In_863,In_1386);
xor U4780 (N_4780,In_1101,In_924);
nand U4781 (N_4781,In_1301,In_306);
xor U4782 (N_4782,In_85,In_797);
or U4783 (N_4783,In_755,In_1079);
and U4784 (N_4784,In_24,In_1219);
nor U4785 (N_4785,In_325,In_747);
and U4786 (N_4786,In_46,In_791);
xnor U4787 (N_4787,In_504,In_1439);
nor U4788 (N_4788,In_231,In_473);
xor U4789 (N_4789,In_697,In_1440);
or U4790 (N_4790,In_788,In_531);
nand U4791 (N_4791,In_190,In_876);
nor U4792 (N_4792,In_989,In_1253);
nand U4793 (N_4793,In_1349,In_1454);
xnor U4794 (N_4794,In_475,In_376);
xnor U4795 (N_4795,In_1090,In_645);
nand U4796 (N_4796,In_1482,In_200);
nand U4797 (N_4797,In_369,In_33);
xnor U4798 (N_4798,In_1291,In_461);
nor U4799 (N_4799,In_1455,In_536);
nor U4800 (N_4800,In_1417,In_1251);
or U4801 (N_4801,In_1124,In_98);
nor U4802 (N_4802,In_71,In_982);
nand U4803 (N_4803,In_253,In_1195);
xnor U4804 (N_4804,In_1021,In_999);
xor U4805 (N_4805,In_271,In_1180);
or U4806 (N_4806,In_639,In_1055);
nand U4807 (N_4807,In_719,In_1023);
nand U4808 (N_4808,In_1372,In_355);
xnor U4809 (N_4809,In_1335,In_250);
nor U4810 (N_4810,In_142,In_1445);
and U4811 (N_4811,In_1198,In_332);
nor U4812 (N_4812,In_1231,In_337);
or U4813 (N_4813,In_1309,In_812);
and U4814 (N_4814,In_475,In_465);
nor U4815 (N_4815,In_54,In_1353);
and U4816 (N_4816,In_1370,In_1076);
nand U4817 (N_4817,In_158,In_485);
or U4818 (N_4818,In_944,In_178);
nor U4819 (N_4819,In_769,In_128);
xor U4820 (N_4820,In_1440,In_18);
nor U4821 (N_4821,In_435,In_296);
or U4822 (N_4822,In_1011,In_247);
xnor U4823 (N_4823,In_1191,In_758);
or U4824 (N_4824,In_1368,In_209);
nor U4825 (N_4825,In_1322,In_1166);
nor U4826 (N_4826,In_896,In_195);
and U4827 (N_4827,In_72,In_1295);
xnor U4828 (N_4828,In_1232,In_257);
or U4829 (N_4829,In_950,In_289);
and U4830 (N_4830,In_944,In_766);
xnor U4831 (N_4831,In_551,In_717);
and U4832 (N_4832,In_295,In_12);
and U4833 (N_4833,In_1051,In_284);
nand U4834 (N_4834,In_970,In_700);
nor U4835 (N_4835,In_1130,In_88);
nand U4836 (N_4836,In_139,In_435);
nor U4837 (N_4837,In_684,In_122);
or U4838 (N_4838,In_1077,In_979);
and U4839 (N_4839,In_571,In_1444);
xnor U4840 (N_4840,In_903,In_1074);
xor U4841 (N_4841,In_1036,In_1496);
nor U4842 (N_4842,In_639,In_976);
and U4843 (N_4843,In_1292,In_1362);
and U4844 (N_4844,In_936,In_1314);
xor U4845 (N_4845,In_1327,In_383);
or U4846 (N_4846,In_66,In_330);
nand U4847 (N_4847,In_701,In_549);
nor U4848 (N_4848,In_913,In_1053);
nand U4849 (N_4849,In_560,In_958);
or U4850 (N_4850,In_235,In_434);
and U4851 (N_4851,In_153,In_1482);
or U4852 (N_4852,In_294,In_1100);
or U4853 (N_4853,In_993,In_1309);
or U4854 (N_4854,In_1042,In_206);
and U4855 (N_4855,In_32,In_1335);
nor U4856 (N_4856,In_1189,In_1394);
or U4857 (N_4857,In_711,In_308);
and U4858 (N_4858,In_1415,In_428);
or U4859 (N_4859,In_1143,In_402);
or U4860 (N_4860,In_926,In_1001);
nand U4861 (N_4861,In_144,In_53);
or U4862 (N_4862,In_1404,In_1459);
nand U4863 (N_4863,In_365,In_851);
and U4864 (N_4864,In_402,In_922);
or U4865 (N_4865,In_1044,In_1369);
xnor U4866 (N_4866,In_1130,In_578);
xor U4867 (N_4867,In_307,In_1024);
and U4868 (N_4868,In_118,In_1112);
or U4869 (N_4869,In_678,In_181);
and U4870 (N_4870,In_151,In_1150);
and U4871 (N_4871,In_1254,In_396);
nor U4872 (N_4872,In_743,In_750);
nand U4873 (N_4873,In_748,In_539);
nand U4874 (N_4874,In_1085,In_392);
xnor U4875 (N_4875,In_49,In_543);
xor U4876 (N_4876,In_757,In_58);
xnor U4877 (N_4877,In_518,In_1284);
nand U4878 (N_4878,In_693,In_1404);
and U4879 (N_4879,In_690,In_359);
xnor U4880 (N_4880,In_1448,In_1413);
and U4881 (N_4881,In_843,In_960);
nor U4882 (N_4882,In_945,In_655);
nor U4883 (N_4883,In_1432,In_701);
xor U4884 (N_4884,In_975,In_679);
and U4885 (N_4885,In_648,In_1086);
nor U4886 (N_4886,In_667,In_981);
or U4887 (N_4887,In_425,In_18);
nor U4888 (N_4888,In_519,In_304);
or U4889 (N_4889,In_1192,In_671);
xor U4890 (N_4890,In_603,In_1069);
nor U4891 (N_4891,In_445,In_1100);
nand U4892 (N_4892,In_1132,In_459);
xor U4893 (N_4893,In_509,In_23);
nor U4894 (N_4894,In_1410,In_255);
nand U4895 (N_4895,In_42,In_319);
nand U4896 (N_4896,In_1185,In_236);
or U4897 (N_4897,In_16,In_927);
nand U4898 (N_4898,In_1099,In_65);
nor U4899 (N_4899,In_721,In_221);
xnor U4900 (N_4900,In_571,In_1426);
nand U4901 (N_4901,In_92,In_1288);
nor U4902 (N_4902,In_969,In_495);
xnor U4903 (N_4903,In_915,In_789);
and U4904 (N_4904,In_443,In_434);
or U4905 (N_4905,In_408,In_1115);
and U4906 (N_4906,In_1131,In_1035);
nand U4907 (N_4907,In_48,In_784);
xor U4908 (N_4908,In_1141,In_379);
and U4909 (N_4909,In_1107,In_1265);
and U4910 (N_4910,In_791,In_63);
nor U4911 (N_4911,In_808,In_1180);
nor U4912 (N_4912,In_875,In_1431);
nor U4913 (N_4913,In_1432,In_1396);
or U4914 (N_4914,In_1148,In_764);
xnor U4915 (N_4915,In_730,In_590);
and U4916 (N_4916,In_1238,In_547);
and U4917 (N_4917,In_1248,In_1113);
and U4918 (N_4918,In_1433,In_598);
and U4919 (N_4919,In_766,In_1353);
and U4920 (N_4920,In_506,In_173);
nor U4921 (N_4921,In_752,In_971);
nor U4922 (N_4922,In_563,In_472);
xor U4923 (N_4923,In_1153,In_914);
nand U4924 (N_4924,In_1238,In_1461);
nand U4925 (N_4925,In_855,In_980);
or U4926 (N_4926,In_162,In_826);
nor U4927 (N_4927,In_878,In_552);
and U4928 (N_4928,In_398,In_1278);
and U4929 (N_4929,In_1193,In_1248);
nand U4930 (N_4930,In_1452,In_727);
and U4931 (N_4931,In_1027,In_28);
nor U4932 (N_4932,In_1282,In_1174);
xnor U4933 (N_4933,In_544,In_765);
xnor U4934 (N_4934,In_1358,In_193);
and U4935 (N_4935,In_793,In_908);
or U4936 (N_4936,In_1480,In_465);
nand U4937 (N_4937,In_1110,In_322);
nand U4938 (N_4938,In_1185,In_263);
and U4939 (N_4939,In_1090,In_164);
nand U4940 (N_4940,In_990,In_1481);
and U4941 (N_4941,In_121,In_409);
nor U4942 (N_4942,In_911,In_187);
or U4943 (N_4943,In_268,In_1337);
xnor U4944 (N_4944,In_1047,In_1036);
or U4945 (N_4945,In_305,In_512);
and U4946 (N_4946,In_58,In_224);
or U4947 (N_4947,In_131,In_1059);
and U4948 (N_4948,In_1477,In_384);
nor U4949 (N_4949,In_658,In_361);
xnor U4950 (N_4950,In_407,In_799);
nand U4951 (N_4951,In_563,In_1346);
and U4952 (N_4952,In_1491,In_184);
nor U4953 (N_4953,In_168,In_464);
xor U4954 (N_4954,In_1166,In_845);
xnor U4955 (N_4955,In_947,In_545);
nand U4956 (N_4956,In_612,In_216);
nor U4957 (N_4957,In_1079,In_380);
nor U4958 (N_4958,In_858,In_749);
nand U4959 (N_4959,In_1011,In_171);
nor U4960 (N_4960,In_1451,In_536);
nand U4961 (N_4961,In_56,In_1291);
nand U4962 (N_4962,In_448,In_774);
xnor U4963 (N_4963,In_159,In_591);
or U4964 (N_4964,In_1434,In_1477);
xnor U4965 (N_4965,In_58,In_1275);
xnor U4966 (N_4966,In_1172,In_1498);
nor U4967 (N_4967,In_72,In_1493);
nand U4968 (N_4968,In_1447,In_1158);
and U4969 (N_4969,In_985,In_736);
nor U4970 (N_4970,In_934,In_204);
or U4971 (N_4971,In_1388,In_20);
or U4972 (N_4972,In_470,In_445);
or U4973 (N_4973,In_1365,In_463);
nand U4974 (N_4974,In_1180,In_1077);
or U4975 (N_4975,In_345,In_617);
and U4976 (N_4976,In_574,In_788);
or U4977 (N_4977,In_270,In_50);
nand U4978 (N_4978,In_151,In_334);
nand U4979 (N_4979,In_988,In_568);
nor U4980 (N_4980,In_506,In_471);
xor U4981 (N_4981,In_1290,In_1153);
or U4982 (N_4982,In_1253,In_145);
nand U4983 (N_4983,In_883,In_62);
or U4984 (N_4984,In_276,In_809);
or U4985 (N_4985,In_345,In_834);
or U4986 (N_4986,In_745,In_889);
nor U4987 (N_4987,In_1146,In_1030);
or U4988 (N_4988,In_491,In_421);
and U4989 (N_4989,In_1021,In_611);
nand U4990 (N_4990,In_689,In_1124);
or U4991 (N_4991,In_986,In_1448);
xnor U4992 (N_4992,In_1318,In_1227);
and U4993 (N_4993,In_735,In_1478);
and U4994 (N_4994,In_1364,In_886);
nor U4995 (N_4995,In_781,In_729);
xnor U4996 (N_4996,In_522,In_1044);
xor U4997 (N_4997,In_925,In_263);
and U4998 (N_4998,In_468,In_0);
or U4999 (N_4999,In_874,In_1204);
nor U5000 (N_5000,N_1610,N_1596);
and U5001 (N_5001,N_1771,N_621);
nor U5002 (N_5002,N_3694,N_343);
nand U5003 (N_5003,N_2275,N_3726);
nor U5004 (N_5004,N_2159,N_411);
nor U5005 (N_5005,N_540,N_1436);
or U5006 (N_5006,N_2993,N_3051);
nand U5007 (N_5007,N_492,N_4197);
xnor U5008 (N_5008,N_2301,N_280);
nor U5009 (N_5009,N_235,N_4971);
or U5010 (N_5010,N_1494,N_416);
or U5011 (N_5011,N_1674,N_4205);
or U5012 (N_5012,N_4858,N_4238);
and U5013 (N_5013,N_4829,N_1754);
nor U5014 (N_5014,N_2422,N_1570);
nor U5015 (N_5015,N_3551,N_3224);
nor U5016 (N_5016,N_2361,N_4187);
xor U5017 (N_5017,N_172,N_2151);
nor U5018 (N_5018,N_4619,N_582);
xnor U5019 (N_5019,N_3680,N_2714);
nor U5020 (N_5020,N_1045,N_1321);
nand U5021 (N_5021,N_41,N_1590);
xor U5022 (N_5022,N_2528,N_2152);
or U5023 (N_5023,N_4066,N_4873);
nor U5024 (N_5024,N_4748,N_3842);
and U5025 (N_5025,N_790,N_3632);
xor U5026 (N_5026,N_3939,N_1390);
or U5027 (N_5027,N_4114,N_3106);
and U5028 (N_5028,N_1,N_3588);
nand U5029 (N_5029,N_1351,N_533);
and U5030 (N_5030,N_2686,N_1244);
nand U5031 (N_5031,N_1406,N_722);
nand U5032 (N_5032,N_1174,N_4515);
xnor U5033 (N_5033,N_4417,N_3681);
and U5034 (N_5034,N_4223,N_186);
or U5035 (N_5035,N_4424,N_4574);
xor U5036 (N_5036,N_1496,N_3633);
xnor U5037 (N_5037,N_1548,N_1577);
xor U5038 (N_5038,N_3643,N_1209);
or U5039 (N_5039,N_2828,N_729);
nor U5040 (N_5040,N_3949,N_3866);
and U5041 (N_5041,N_2657,N_1755);
nand U5042 (N_5042,N_3017,N_652);
xnor U5043 (N_5043,N_3347,N_2386);
xnor U5044 (N_5044,N_3371,N_4906);
and U5045 (N_5045,N_3284,N_1629);
xnor U5046 (N_5046,N_1928,N_2757);
nor U5047 (N_5047,N_4561,N_1645);
and U5048 (N_5048,N_4026,N_2506);
and U5049 (N_5049,N_2273,N_4474);
xor U5050 (N_5050,N_3428,N_1361);
and U5051 (N_5051,N_1793,N_4013);
and U5052 (N_5052,N_2149,N_4936);
and U5053 (N_5053,N_4658,N_3293);
or U5054 (N_5054,N_4449,N_4563);
xnor U5055 (N_5055,N_846,N_4673);
xor U5056 (N_5056,N_4544,N_2392);
nor U5057 (N_5057,N_4554,N_2721);
nand U5058 (N_5058,N_701,N_1991);
nand U5059 (N_5059,N_2365,N_2784);
and U5060 (N_5060,N_3008,N_3395);
xnor U5061 (N_5061,N_2990,N_4470);
and U5062 (N_5062,N_4097,N_1862);
xor U5063 (N_5063,N_1118,N_4108);
nor U5064 (N_5064,N_30,N_1083);
xnor U5065 (N_5065,N_3087,N_4074);
and U5066 (N_5066,N_3171,N_919);
nand U5067 (N_5067,N_1753,N_1847);
xor U5068 (N_5068,N_1318,N_4568);
or U5069 (N_5069,N_2127,N_3070);
xor U5070 (N_5070,N_2296,N_2344);
nand U5071 (N_5071,N_261,N_4404);
nand U5072 (N_5072,N_2955,N_3707);
or U5073 (N_5073,N_631,N_3699);
nor U5074 (N_5074,N_1395,N_400);
and U5075 (N_5075,N_331,N_3378);
and U5076 (N_5076,N_578,N_3442);
or U5077 (N_5077,N_1331,N_3484);
nor U5078 (N_5078,N_2915,N_4476);
or U5079 (N_5079,N_4148,N_3568);
and U5080 (N_5080,N_3324,N_2023);
xor U5081 (N_5081,N_1587,N_544);
nand U5082 (N_5082,N_2705,N_4692);
nor U5083 (N_5083,N_2269,N_2608);
nor U5084 (N_5084,N_949,N_402);
nor U5085 (N_5085,N_1023,N_1861);
and U5086 (N_5086,N_1636,N_2450);
or U5087 (N_5087,N_1867,N_2548);
xor U5088 (N_5088,N_1574,N_315);
nor U5089 (N_5089,N_3461,N_75);
nor U5090 (N_5090,N_1280,N_1490);
xor U5091 (N_5091,N_1970,N_4096);
nand U5092 (N_5092,N_2055,N_2797);
xor U5093 (N_5093,N_3056,N_1612);
xor U5094 (N_5094,N_387,N_4229);
nand U5095 (N_5095,N_3407,N_1917);
nor U5096 (N_5096,N_951,N_1388);
xnor U5097 (N_5097,N_4932,N_1937);
xnor U5098 (N_5098,N_2138,N_3869);
xor U5099 (N_5099,N_926,N_2054);
nor U5100 (N_5100,N_3370,N_1507);
nand U5101 (N_5101,N_4968,N_433);
and U5102 (N_5102,N_4126,N_548);
or U5103 (N_5103,N_1263,N_589);
and U5104 (N_5104,N_2170,N_1890);
nor U5105 (N_5105,N_3006,N_1832);
or U5106 (N_5106,N_4282,N_3543);
nand U5107 (N_5107,N_1794,N_284);
nand U5108 (N_5108,N_1541,N_4200);
xor U5109 (N_5109,N_369,N_4764);
and U5110 (N_5110,N_2350,N_4448);
nand U5111 (N_5111,N_4718,N_1520);
and U5112 (N_5112,N_3848,N_4443);
nor U5113 (N_5113,N_2319,N_2626);
and U5114 (N_5114,N_160,N_368);
nand U5115 (N_5115,N_25,N_2562);
and U5116 (N_5116,N_2903,N_1271);
or U5117 (N_5117,N_4194,N_755);
or U5118 (N_5118,N_4738,N_3014);
nor U5119 (N_5119,N_3659,N_3291);
nor U5120 (N_5120,N_735,N_1257);
or U5121 (N_5121,N_1692,N_1880);
xnor U5122 (N_5122,N_3327,N_546);
and U5123 (N_5123,N_678,N_1342);
and U5124 (N_5124,N_4683,N_86);
nor U5125 (N_5125,N_18,N_4261);
and U5126 (N_5126,N_2413,N_691);
nor U5127 (N_5127,N_639,N_1500);
and U5128 (N_5128,N_1329,N_4918);
and U5129 (N_5129,N_458,N_214);
or U5130 (N_5130,N_4007,N_2015);
nand U5131 (N_5131,N_1821,N_989);
or U5132 (N_5132,N_2699,N_4796);
or U5133 (N_5133,N_3987,N_4479);
nand U5134 (N_5134,N_1872,N_2980);
nor U5135 (N_5135,N_1077,N_4857);
or U5136 (N_5136,N_1048,N_3228);
nor U5137 (N_5137,N_2096,N_3635);
xor U5138 (N_5138,N_2095,N_4178);
nand U5139 (N_5139,N_1094,N_3063);
nor U5140 (N_5140,N_2813,N_3487);
and U5141 (N_5141,N_4402,N_1243);
and U5142 (N_5142,N_62,N_1362);
nand U5143 (N_5143,N_1537,N_3620);
nand U5144 (N_5144,N_4629,N_1001);
xor U5145 (N_5145,N_4254,N_2433);
xor U5146 (N_5146,N_3522,N_1325);
nor U5147 (N_5147,N_1995,N_1979);
and U5148 (N_5148,N_3211,N_2162);
and U5149 (N_5149,N_1032,N_3970);
nand U5150 (N_5150,N_126,N_625);
and U5151 (N_5151,N_2382,N_675);
and U5152 (N_5152,N_3776,N_2524);
nor U5153 (N_5153,N_2728,N_3828);
nand U5154 (N_5154,N_3373,N_1037);
xnor U5155 (N_5155,N_4874,N_3737);
and U5156 (N_5156,N_2173,N_4961);
xnor U5157 (N_5157,N_291,N_2567);
and U5158 (N_5158,N_3241,N_2012);
and U5159 (N_5159,N_636,N_2338);
nor U5160 (N_5160,N_2930,N_915);
nor U5161 (N_5161,N_4980,N_3908);
nand U5162 (N_5162,N_689,N_3074);
nor U5163 (N_5163,N_3155,N_2855);
nand U5164 (N_5164,N_19,N_76);
nor U5165 (N_5165,N_2545,N_4422);
or U5166 (N_5166,N_4521,N_3937);
nor U5167 (N_5167,N_107,N_1007);
nand U5168 (N_5168,N_2617,N_728);
nor U5169 (N_5169,N_4868,N_3384);
nand U5170 (N_5170,N_993,N_571);
or U5171 (N_5171,N_3141,N_2972);
nand U5172 (N_5172,N_92,N_3863);
nand U5173 (N_5173,N_2364,N_1474);
nor U5174 (N_5174,N_1741,N_1260);
or U5175 (N_5175,N_2449,N_3901);
nor U5176 (N_5176,N_3001,N_3683);
xnor U5177 (N_5177,N_4856,N_2543);
nor U5178 (N_5178,N_1671,N_3798);
xnor U5179 (N_5179,N_435,N_1054);
and U5180 (N_5180,N_3372,N_462);
nand U5181 (N_5181,N_769,N_499);
xor U5182 (N_5182,N_3202,N_145);
xor U5183 (N_5183,N_3116,N_190);
or U5184 (N_5184,N_3296,N_773);
nand U5185 (N_5185,N_1141,N_590);
or U5186 (N_5186,N_897,N_2441);
and U5187 (N_5187,N_4080,N_1543);
nor U5188 (N_5188,N_1323,N_4728);
and U5189 (N_5189,N_2654,N_1288);
nor U5190 (N_5190,N_2230,N_2696);
or U5191 (N_5191,N_2878,N_1091);
or U5192 (N_5192,N_307,N_2651);
nand U5193 (N_5193,N_2925,N_136);
and U5194 (N_5194,N_1647,N_1497);
nor U5195 (N_5195,N_924,N_2363);
and U5196 (N_5196,N_4896,N_4835);
and U5197 (N_5197,N_4029,N_1585);
xnor U5198 (N_5198,N_1104,N_57);
nor U5199 (N_5199,N_4668,N_2438);
nand U5200 (N_5200,N_798,N_3130);
nor U5201 (N_5201,N_3611,N_2957);
and U5202 (N_5202,N_920,N_1643);
nor U5203 (N_5203,N_2034,N_2541);
and U5204 (N_5204,N_2675,N_4837);
xnor U5205 (N_5205,N_2819,N_2107);
nand U5206 (N_5206,N_3102,N_4297);
nand U5207 (N_5207,N_228,N_3058);
or U5208 (N_5208,N_4885,N_1020);
nand U5209 (N_5209,N_4504,N_1178);
xor U5210 (N_5210,N_2157,N_1655);
nand U5211 (N_5211,N_3689,N_4957);
and U5212 (N_5212,N_240,N_4712);
xnor U5213 (N_5213,N_3482,N_3899);
xnor U5214 (N_5214,N_3462,N_4503);
nor U5215 (N_5215,N_4320,N_4319);
xor U5216 (N_5216,N_2471,N_3005);
and U5217 (N_5217,N_3380,N_3921);
and U5218 (N_5218,N_3464,N_182);
nand U5219 (N_5219,N_109,N_4953);
and U5220 (N_5220,N_1787,N_1234);
xnor U5221 (N_5221,N_4087,N_1555);
or U5222 (N_5222,N_3121,N_3670);
nor U5223 (N_5223,N_4921,N_1146);
and U5224 (N_5224,N_3920,N_8);
or U5225 (N_5225,N_2971,N_3506);
or U5226 (N_5226,N_4484,N_204);
nor U5227 (N_5227,N_4999,N_4491);
xor U5228 (N_5228,N_2985,N_2777);
nand U5229 (N_5229,N_858,N_4979);
and U5230 (N_5230,N_4747,N_223);
nand U5231 (N_5231,N_1412,N_2292);
or U5232 (N_5232,N_2901,N_3069);
xor U5233 (N_5233,N_991,N_99);
or U5234 (N_5234,N_3795,N_4305);
nand U5235 (N_5235,N_114,N_1525);
and U5236 (N_5236,N_889,N_4162);
nor U5237 (N_5237,N_2771,N_4382);
nand U5238 (N_5238,N_1644,N_3529);
nand U5239 (N_5239,N_1954,N_2927);
nand U5240 (N_5240,N_3422,N_2519);
nand U5241 (N_5241,N_1857,N_4199);
and U5242 (N_5242,N_4407,N_2360);
or U5243 (N_5243,N_3287,N_560);
nor U5244 (N_5244,N_4710,N_3650);
xnor U5245 (N_5245,N_3587,N_1281);
nor U5246 (N_5246,N_3747,N_724);
or U5247 (N_5247,N_4102,N_1429);
nor U5248 (N_5248,N_1955,N_4165);
and U5249 (N_5249,N_4111,N_4793);
and U5250 (N_5250,N_189,N_2470);
nor U5251 (N_5251,N_699,N_4555);
and U5252 (N_5252,N_1557,N_3988);
xnor U5253 (N_5253,N_1877,N_2199);
nand U5254 (N_5254,N_1481,N_1873);
xnor U5255 (N_5255,N_1354,N_2482);
xnor U5256 (N_5256,N_4628,N_1560);
nor U5257 (N_5257,N_4944,N_2135);
xor U5258 (N_5258,N_2600,N_1367);
nand U5259 (N_5259,N_3193,N_4357);
and U5260 (N_5260,N_3825,N_1166);
nand U5261 (N_5261,N_4883,N_4630);
and U5262 (N_5262,N_3402,N_1634);
xor U5263 (N_5263,N_4091,N_1571);
nand U5264 (N_5264,N_1947,N_4751);
and U5265 (N_5265,N_4154,N_2517);
or U5266 (N_5266,N_570,N_3230);
xnor U5267 (N_5267,N_1062,N_4410);
or U5268 (N_5268,N_1295,N_285);
nor U5269 (N_5269,N_719,N_3311);
or U5270 (N_5270,N_312,N_3416);
or U5271 (N_5271,N_4132,N_4542);
nor U5272 (N_5272,N_1725,N_1215);
nor U5273 (N_5273,N_4020,N_1370);
and U5274 (N_5274,N_3978,N_2687);
nand U5275 (N_5275,N_3527,N_2209);
and U5276 (N_5276,N_1504,N_2581);
and U5277 (N_5277,N_3984,N_1138);
or U5278 (N_5278,N_2504,N_3082);
or U5279 (N_5279,N_992,N_3834);
xnor U5280 (N_5280,N_3467,N_4898);
nand U5281 (N_5281,N_3318,N_4733);
or U5282 (N_5282,N_3674,N_2277);
xor U5283 (N_5283,N_4820,N_826);
and U5284 (N_5284,N_2045,N_606);
or U5285 (N_5285,N_3278,N_3943);
or U5286 (N_5286,N_1828,N_562);
nor U5287 (N_5287,N_2025,N_4204);
nand U5288 (N_5288,N_3500,N_3596);
or U5289 (N_5289,N_2803,N_3275);
xnor U5290 (N_5290,N_2412,N_4144);
or U5291 (N_5291,N_1907,N_3267);
xor U5292 (N_5292,N_4564,N_3104);
xor U5293 (N_5293,N_4201,N_739);
xnor U5294 (N_5294,N_4441,N_1874);
or U5295 (N_5295,N_4966,N_4036);
nor U5296 (N_5296,N_2087,N_4175);
and U5297 (N_5297,N_687,N_3675);
xor U5298 (N_5298,N_592,N_3062);
xor U5299 (N_5299,N_3317,N_4250);
nand U5300 (N_5300,N_3796,N_2465);
and U5301 (N_5301,N_4602,N_923);
nor U5302 (N_5302,N_3367,N_267);
or U5303 (N_5303,N_2610,N_2492);
nor U5304 (N_5304,N_3332,N_1151);
and U5305 (N_5305,N_464,N_667);
and U5306 (N_5306,N_1391,N_2329);
nand U5307 (N_5307,N_3927,N_179);
and U5308 (N_5308,N_1355,N_4497);
xnor U5309 (N_5309,N_4789,N_1898);
nor U5310 (N_5310,N_4231,N_1482);
xor U5311 (N_5311,N_855,N_1373);
xnor U5312 (N_5312,N_2232,N_2720);
xor U5313 (N_5313,N_2516,N_3656);
nand U5314 (N_5314,N_273,N_850);
and U5315 (N_5315,N_513,N_3055);
or U5316 (N_5316,N_155,N_3786);
xnor U5317 (N_5317,N_1275,N_2487);
or U5318 (N_5318,N_3146,N_21);
or U5319 (N_5319,N_1074,N_1471);
nor U5320 (N_5320,N_3956,N_688);
nor U5321 (N_5321,N_1484,N_3710);
xnor U5322 (N_5322,N_1110,N_2768);
nor U5323 (N_5323,N_4069,N_2748);
nand U5324 (N_5324,N_1624,N_479);
xor U5325 (N_5325,N_2835,N_1819);
nand U5326 (N_5326,N_2084,N_586);
and U5327 (N_5327,N_3530,N_1971);
nor U5328 (N_5328,N_805,N_2461);
or U5329 (N_5329,N_4084,N_4765);
and U5330 (N_5330,N_1473,N_1221);
nand U5331 (N_5331,N_187,N_4622);
or U5332 (N_5332,N_2817,N_3509);
or U5333 (N_5333,N_1508,N_842);
nand U5334 (N_5334,N_975,N_2206);
xor U5335 (N_5335,N_1811,N_620);
nand U5336 (N_5336,N_1241,N_4060);
and U5337 (N_5337,N_1818,N_3405);
and U5338 (N_5338,N_4090,N_2463);
xnor U5339 (N_5339,N_1369,N_4294);
or U5340 (N_5340,N_4092,N_1068);
and U5341 (N_5341,N_4083,N_1478);
nand U5342 (N_5342,N_597,N_4444);
nand U5343 (N_5343,N_81,N_3281);
nand U5344 (N_5344,N_1977,N_3011);
xnor U5345 (N_5345,N_4335,N_1598);
nor U5346 (N_5346,N_3238,N_1777);
and U5347 (N_5347,N_1237,N_445);
nand U5348 (N_5348,N_1453,N_2333);
and U5349 (N_5349,N_2457,N_2962);
nor U5350 (N_5350,N_2847,N_4749);
or U5351 (N_5351,N_1393,N_736);
or U5352 (N_5352,N_4705,N_4725);
and U5353 (N_5353,N_686,N_1153);
nor U5354 (N_5354,N_3639,N_1733);
xor U5355 (N_5355,N_4587,N_4726);
nand U5356 (N_5356,N_221,N_4527);
nor U5357 (N_5357,N_1056,N_3678);
xnor U5358 (N_5358,N_340,N_1885);
and U5359 (N_5359,N_4578,N_1942);
xor U5360 (N_5360,N_2443,N_3410);
nand U5361 (N_5361,N_4744,N_591);
xor U5362 (N_5362,N_4797,N_1595);
nor U5363 (N_5363,N_1495,N_3358);
and U5364 (N_5364,N_1195,N_508);
nand U5365 (N_5365,N_3583,N_230);
or U5366 (N_5366,N_3301,N_281);
xor U5367 (N_5367,N_1035,N_3337);
or U5368 (N_5368,N_164,N_2538);
nor U5369 (N_5369,N_4420,N_1652);
and U5370 (N_5370,N_3837,N_3991);
xnor U5371 (N_5371,N_2631,N_1080);
nor U5372 (N_5372,N_2466,N_199);
and U5373 (N_5373,N_2369,N_1842);
nand U5374 (N_5374,N_4827,N_4845);
or U5375 (N_5375,N_4812,N_3456);
nand U5376 (N_5376,N_3375,N_4987);
nor U5377 (N_5377,N_595,N_3609);
and U5378 (N_5378,N_4485,N_1408);
or U5379 (N_5379,N_3905,N_1605);
or U5380 (N_5380,N_2073,N_2573);
and U5381 (N_5381,N_4643,N_4607);
or U5382 (N_5382,N_2359,N_2964);
or U5383 (N_5383,N_4455,N_4324);
and U5384 (N_5384,N_2348,N_4049);
xor U5385 (N_5385,N_1510,N_4522);
nand U5386 (N_5386,N_602,N_1681);
and U5387 (N_5387,N_242,N_4051);
or U5388 (N_5388,N_173,N_4805);
nand U5389 (N_5389,N_231,N_2841);
and U5390 (N_5390,N_3954,N_3858);
and U5391 (N_5391,N_741,N_3701);
nor U5392 (N_5392,N_1006,N_3239);
xor U5393 (N_5393,N_4945,N_4287);
nor U5394 (N_5394,N_52,N_2026);
or U5395 (N_5395,N_467,N_4477);
nand U5396 (N_5396,N_3963,N_598);
or U5397 (N_5397,N_1027,N_4890);
or U5398 (N_5398,N_4866,N_1722);
nor U5399 (N_5399,N_3974,N_506);
and U5400 (N_5400,N_1988,N_4262);
or U5401 (N_5401,N_1684,N_2346);
nand U5402 (N_5402,N_1588,N_2027);
xnor U5403 (N_5403,N_1090,N_2316);
and U5404 (N_5404,N_896,N_4513);
and U5405 (N_5405,N_1950,N_1366);
nand U5406 (N_5406,N_3919,N_1606);
nand U5407 (N_5407,N_2306,N_3809);
xnor U5408 (N_5408,N_626,N_4266);
xnor U5409 (N_5409,N_1107,N_2884);
xor U5410 (N_5410,N_717,N_2986);
or U5411 (N_5411,N_3857,N_4452);
nand U5412 (N_5412,N_2578,N_3816);
nor U5413 (N_5413,N_4021,N_3619);
xnor U5414 (N_5414,N_1120,N_295);
and U5415 (N_5415,N_780,N_1155);
nand U5416 (N_5416,N_4997,N_3401);
nor U5417 (N_5417,N_4716,N_2837);
nand U5418 (N_5418,N_2659,N_2263);
and U5419 (N_5419,N_2935,N_4881);
or U5420 (N_5420,N_2670,N_3714);
xor U5421 (N_5421,N_1274,N_4654);
nand U5422 (N_5422,N_821,N_3531);
nand U5423 (N_5423,N_1765,N_1929);
xor U5424 (N_5424,N_2838,N_2793);
nor U5425 (N_5425,N_3763,N_89);
nand U5426 (N_5426,N_3696,N_3010);
nor U5427 (N_5427,N_1173,N_1459);
and U5428 (N_5428,N_3466,N_49);
nand U5429 (N_5429,N_1308,N_927);
and U5430 (N_5430,N_2483,N_398);
xor U5431 (N_5431,N_2717,N_568);
or U5432 (N_5432,N_1921,N_2039);
or U5433 (N_5433,N_4946,N_913);
xnor U5434 (N_5434,N_4766,N_2940);
nor U5435 (N_5435,N_1569,N_1365);
nand U5436 (N_5436,N_3789,N_1403);
nand U5437 (N_5437,N_2900,N_4686);
or U5438 (N_5438,N_4572,N_4969);
and U5439 (N_5439,N_4865,N_3212);
nand U5440 (N_5440,N_4363,N_314);
or U5441 (N_5441,N_4028,N_4219);
nand U5442 (N_5442,N_262,N_1546);
xnor U5443 (N_5443,N_4188,N_429);
nand U5444 (N_5444,N_2380,N_2673);
nand U5445 (N_5445,N_4304,N_1302);
nor U5446 (N_5446,N_1043,N_3233);
or U5447 (N_5447,N_1619,N_2451);
nand U5448 (N_5448,N_2260,N_1310);
and U5449 (N_5449,N_372,N_731);
nor U5450 (N_5450,N_2020,N_4408);
nand U5451 (N_5451,N_672,N_515);
or U5452 (N_5452,N_3031,N_4112);
nand U5453 (N_5453,N_567,N_105);
or U5454 (N_5454,N_3071,N_654);
xor U5455 (N_5455,N_1661,N_500);
and U5456 (N_5456,N_194,N_3061);
or U5457 (N_5457,N_4173,N_1039);
nand U5458 (N_5458,N_3137,N_4939);
and U5459 (N_5459,N_4708,N_1581);
nor U5460 (N_5460,N_1816,N_1925);
nor U5461 (N_5461,N_3517,N_2899);
nor U5462 (N_5462,N_2709,N_4149);
or U5463 (N_5463,N_1224,N_191);
xor U5464 (N_5464,N_1071,N_3345);
and U5465 (N_5465,N_502,N_2692);
nor U5466 (N_5466,N_632,N_225);
or U5467 (N_5467,N_3120,N_348);
nor U5468 (N_5468,N_4350,N_3035);
or U5469 (N_5469,N_4687,N_2776);
nor U5470 (N_5470,N_704,N_4230);
and U5471 (N_5471,N_3854,N_3580);
nor U5472 (N_5472,N_1524,N_2355);
and U5473 (N_5473,N_1058,N_4806);
nand U5474 (N_5474,N_3925,N_565);
nor U5475 (N_5475,N_3297,N_1129);
nand U5476 (N_5476,N_3455,N_4481);
nor U5477 (N_5477,N_2833,N_4160);
xnor U5478 (N_5478,N_2808,N_1121);
nand U5479 (N_5479,N_3549,N_723);
xor U5480 (N_5480,N_745,N_520);
nand U5481 (N_5481,N_864,N_4253);
nand U5482 (N_5482,N_1079,N_345);
xnor U5483 (N_5483,N_824,N_3030);
xnor U5484 (N_5484,N_2535,N_3019);
or U5485 (N_5485,N_3057,N_335);
and U5486 (N_5486,N_3443,N_1330);
nand U5487 (N_5487,N_4798,N_1761);
nor U5488 (N_5488,N_4743,N_3762);
and U5489 (N_5489,N_3073,N_4581);
xor U5490 (N_5490,N_121,N_1812);
xnor U5491 (N_5491,N_3579,N_1868);
and U5492 (N_5492,N_4489,N_1608);
or U5493 (N_5493,N_4821,N_353);
and U5494 (N_5494,N_2307,N_2794);
nor U5495 (N_5495,N_2253,N_3232);
and U5496 (N_5496,N_1445,N_912);
nand U5497 (N_5497,N_48,N_1906);
or U5498 (N_5498,N_1517,N_2342);
or U5499 (N_5499,N_969,N_1164);
nor U5500 (N_5500,N_658,N_3430);
xor U5501 (N_5501,N_1716,N_3878);
or U5502 (N_5502,N_808,N_4398);
nor U5503 (N_5503,N_4843,N_4494);
or U5504 (N_5504,N_2224,N_1152);
or U5505 (N_5505,N_3237,N_1276);
xor U5506 (N_5506,N_4442,N_2791);
or U5507 (N_5507,N_2832,N_3495);
nor U5508 (N_5508,N_2630,N_985);
or U5509 (N_5509,N_2379,N_1827);
nand U5510 (N_5510,N_2700,N_967);
xnor U5511 (N_5511,N_1651,N_4888);
and U5512 (N_5512,N_4955,N_146);
xor U5513 (N_5513,N_4889,N_2210);
or U5514 (N_5514,N_661,N_176);
xor U5515 (N_5515,N_3493,N_2143);
and U5516 (N_5516,N_3460,N_1586);
nor U5517 (N_5517,N_3032,N_1087);
xnor U5518 (N_5518,N_1960,N_1347);
xnor U5519 (N_5519,N_2726,N_2373);
xnor U5520 (N_5520,N_2858,N_2689);
nand U5521 (N_5521,N_2007,N_1371);
or U5522 (N_5522,N_4973,N_157);
xnor U5523 (N_5523,N_981,N_3119);
or U5524 (N_5524,N_2425,N_493);
and U5525 (N_5525,N_4316,N_430);
nand U5526 (N_5526,N_702,N_2734);
and U5527 (N_5527,N_3218,N_3148);
or U5528 (N_5528,N_2521,N_59);
xnor U5529 (N_5529,N_3967,N_3615);
nand U5530 (N_5530,N_271,N_2091);
nor U5531 (N_5531,N_3458,N_3882);
nand U5532 (N_5532,N_3344,N_1172);
xor U5533 (N_5533,N_758,N_2399);
nand U5534 (N_5534,N_3894,N_2326);
and U5535 (N_5535,N_1358,N_2278);
or U5536 (N_5536,N_4169,N_3748);
or U5537 (N_5537,N_471,N_3865);
nor U5538 (N_5538,N_1536,N_3981);
nand U5539 (N_5539,N_2409,N_3750);
nand U5540 (N_5540,N_922,N_4326);
and U5541 (N_5541,N_2678,N_1304);
nor U5542 (N_5542,N_1600,N_4739);
and U5543 (N_5543,N_3135,N_3366);
nand U5544 (N_5544,N_1106,N_2737);
nand U5545 (N_5545,N_3195,N_3704);
nor U5546 (N_5546,N_1303,N_3829);
nand U5547 (N_5547,N_4085,N_1452);
and U5548 (N_5548,N_1593,N_1191);
and U5549 (N_5549,N_1024,N_998);
or U5550 (N_5550,N_4614,N_2762);
or U5551 (N_5551,N_787,N_3187);
or U5552 (N_5552,N_366,N_818);
xor U5553 (N_5553,N_666,N_814);
nor U5554 (N_5554,N_670,N_1749);
nand U5555 (N_5555,N_4537,N_272);
nand U5556 (N_5556,N_4756,N_2040);
and U5557 (N_5557,N_3013,N_2661);
nor U5558 (N_5558,N_1807,N_2396);
and U5559 (N_5559,N_2475,N_4236);
and U5560 (N_5560,N_3593,N_1213);
xor U5561 (N_5561,N_1943,N_4972);
and U5562 (N_5562,N_4068,N_970);
and U5563 (N_5563,N_1559,N_456);
nand U5564 (N_5564,N_2434,N_2501);
nand U5565 (N_5565,N_4719,N_2590);
nor U5566 (N_5566,N_3768,N_1618);
and U5567 (N_5567,N_3389,N_718);
nand U5568 (N_5568,N_1808,N_3185);
nor U5569 (N_5569,N_2973,N_2540);
nand U5570 (N_5570,N_4009,N_680);
nand U5571 (N_5571,N_2003,N_749);
or U5572 (N_5572,N_1205,N_1211);
xor U5573 (N_5573,N_2769,N_694);
or U5574 (N_5574,N_4958,N_637);
nand U5575 (N_5575,N_2367,N_4168);
nor U5576 (N_5576,N_3623,N_2178);
or U5577 (N_5577,N_3733,N_1568);
and U5578 (N_5578,N_4548,N_208);
nand U5579 (N_5579,N_2378,N_4644);
and U5580 (N_5580,N_3732,N_1981);
and U5581 (N_5581,N_539,N_3702);
xor U5582 (N_5582,N_3716,N_1134);
or U5583 (N_5583,N_630,N_2658);
xnor U5584 (N_5584,N_4433,N_4900);
nor U5585 (N_5585,N_3169,N_70);
and U5586 (N_5586,N_1112,N_3603);
and U5587 (N_5587,N_2556,N_2298);
nor U5588 (N_5588,N_645,N_1299);
xor U5589 (N_5589,N_1127,N_2056);
nand U5590 (N_5590,N_347,N_2052);
xnor U5591 (N_5591,N_1378,N_2375);
nor U5592 (N_5592,N_4251,N_1089);
nor U5593 (N_5593,N_2974,N_4355);
and U5594 (N_5594,N_2708,N_3891);
nor U5595 (N_5595,N_1964,N_2197);
or U5596 (N_5596,N_2607,N_4482);
and U5597 (N_5597,N_2041,N_298);
xor U5598 (N_5598,N_3952,N_4609);
nand U5599 (N_5599,N_2963,N_4315);
or U5600 (N_5600,N_1066,N_2534);
or U5601 (N_5601,N_2806,N_1298);
nor U5602 (N_5602,N_2145,N_1640);
nand U5603 (N_5603,N_2787,N_1806);
nand U5604 (N_5604,N_2752,N_3867);
and U5605 (N_5605,N_2530,N_2976);
xnor U5606 (N_5606,N_3946,N_1742);
or U5607 (N_5607,N_2381,N_4437);
and U5608 (N_5608,N_4904,N_2036);
nor U5609 (N_5609,N_1871,N_2010);
nor U5610 (N_5610,N_1855,N_1067);
nor U5611 (N_5611,N_373,N_2882);
or U5612 (N_5612,N_2848,N_916);
and U5613 (N_5613,N_4274,N_984);
or U5614 (N_5614,N_3631,N_3942);
nand U5615 (N_5615,N_193,N_1477);
or U5616 (N_5616,N_1025,N_768);
xor U5617 (N_5617,N_4788,N_3183);
or U5618 (N_5618,N_1597,N_3508);
nand U5619 (N_5619,N_143,N_389);
and U5620 (N_5620,N_4052,N_871);
xor U5621 (N_5621,N_3864,N_774);
or U5622 (N_5622,N_2515,N_3325);
xor U5623 (N_5623,N_3432,N_3663);
and U5624 (N_5624,N_894,N_2225);
nor U5625 (N_5625,N_3536,N_2906);
nor U5626 (N_5626,N_4483,N_881);
nand U5627 (N_5627,N_707,N_4425);
or U5628 (N_5628,N_3885,N_3602);
nor U5629 (N_5629,N_3640,N_4839);
or U5630 (N_5630,N_1105,N_3958);
and U5631 (N_5631,N_2554,N_1797);
or U5632 (N_5632,N_933,N_4996);
and U5633 (N_5633,N_614,N_1724);
xnor U5634 (N_5634,N_409,N_4191);
xor U5635 (N_5635,N_4283,N_4399);
or U5636 (N_5636,N_2710,N_4523);
nor U5637 (N_5637,N_381,N_4757);
and U5638 (N_5638,N_3986,N_2743);
xnor U5639 (N_5639,N_4895,N_3998);
or U5640 (N_5640,N_1439,N_3969);
xor U5641 (N_5641,N_2684,N_3161);
and U5642 (N_5642,N_2169,N_1814);
xnor U5643 (N_5643,N_2424,N_1059);
or U5644 (N_5644,N_1589,N_2886);
nand U5645 (N_5645,N_1572,N_2426);
or U5646 (N_5646,N_4682,N_3851);
nand U5647 (N_5647,N_4978,N_3447);
and U5648 (N_5648,N_149,N_1082);
nand U5649 (N_5649,N_1075,N_3727);
or U5650 (N_5650,N_779,N_3788);
nand U5651 (N_5651,N_2477,N_2038);
nor U5652 (N_5652,N_4190,N_3305);
nand U5653 (N_5653,N_465,N_3605);
and U5654 (N_5654,N_711,N_3453);
xnor U5655 (N_5655,N_2852,N_2931);
or U5656 (N_5656,N_1233,N_3273);
or U5657 (N_5657,N_1664,N_4511);
nor U5658 (N_5658,N_408,N_2706);
nor U5659 (N_5659,N_2401,N_1252);
or U5660 (N_5660,N_573,N_4288);
or U5661 (N_5661,N_3496,N_2814);
and U5662 (N_5662,N_738,N_1604);
nand U5663 (N_5663,N_1222,N_65);
nand U5664 (N_5664,N_1004,N_883);
or U5665 (N_5665,N_882,N_4549);
xor U5666 (N_5666,N_3944,N_2219);
or U5667 (N_5667,N_3491,N_2895);
nor U5668 (N_5668,N_4198,N_2198);
xor U5669 (N_5669,N_3566,N_660);
nor U5670 (N_5670,N_4956,N_3784);
or U5671 (N_5671,N_2207,N_2693);
and U5672 (N_5672,N_3098,N_3997);
or U5673 (N_5673,N_4634,N_4415);
nand U5674 (N_5674,N_1349,N_928);
xnor U5675 (N_5675,N_3236,N_2086);
nand U5676 (N_5676,N_1905,N_2097);
nor U5677 (N_5677,N_2954,N_3805);
and U5678 (N_5678,N_1846,N_2368);
nor U5679 (N_5679,N_2865,N_1864);
nand U5680 (N_5680,N_405,N_1642);
xor U5681 (N_5681,N_1277,N_817);
xor U5682 (N_5682,N_2377,N_1051);
and U5683 (N_5683,N_2476,N_3930);
and U5684 (N_5684,N_587,N_4340);
or U5685 (N_5685,N_2388,N_3652);
and U5686 (N_5686,N_357,N_29);
nor U5687 (N_5687,N_2137,N_3856);
xnor U5688 (N_5688,N_4700,N_2759);
nor U5689 (N_5689,N_4911,N_4930);
and U5690 (N_5690,N_2458,N_4438);
nor U5691 (N_5691,N_3923,N_2897);
nor U5692 (N_5692,N_1952,N_3697);
or U5693 (N_5693,N_893,N_1180);
nand U5694 (N_5694,N_3409,N_1161);
or U5695 (N_5695,N_3379,N_4291);
nand U5696 (N_5696,N_2989,N_4931);
nor U5697 (N_5697,N_2894,N_2764);
nor U5698 (N_5698,N_3552,N_2616);
xnor U5699 (N_5699,N_4280,N_3262);
and U5700 (N_5700,N_599,N_4531);
nor U5701 (N_5701,N_2741,N_2510);
xor U5702 (N_5702,N_3221,N_1799);
or U5703 (N_5703,N_1542,N_1663);
and U5704 (N_5704,N_4672,N_236);
nand U5705 (N_5705,N_1189,N_2332);
and U5706 (N_5706,N_2261,N_3875);
xnor U5707 (N_5707,N_1479,N_831);
and U5708 (N_5708,N_2440,N_4794);
nor U5709 (N_5709,N_1334,N_4412);
or U5710 (N_5710,N_1502,N_3249);
and U5711 (N_5711,N_941,N_380);
nor U5712 (N_5712,N_1665,N_607);
xnor U5713 (N_5713,N_4818,N_268);
nor U5714 (N_5714,N_2645,N_664);
and U5715 (N_5715,N_942,N_4395);
or U5716 (N_5716,N_3860,N_876);
xnor U5717 (N_5717,N_4892,N_4055);
and U5718 (N_5718,N_4934,N_791);
nor U5719 (N_5719,N_3444,N_28);
or U5720 (N_5720,N_2996,N_3368);
nand U5721 (N_5721,N_150,N_3922);
xnor U5722 (N_5722,N_651,N_2896);
nand U5723 (N_5723,N_3940,N_1719);
or U5724 (N_5724,N_4982,N_2498);
and U5725 (N_5725,N_4848,N_1448);
nor U5726 (N_5726,N_3159,N_1782);
or U5727 (N_5727,N_2415,N_3773);
or U5728 (N_5728,N_4400,N_3992);
nand U5729 (N_5729,N_337,N_1427);
xnor U5730 (N_5730,N_2189,N_2862);
and U5731 (N_5731,N_901,N_2648);
xnor U5732 (N_5732,N_1450,N_961);
or U5733 (N_5733,N_974,N_2289);
xor U5734 (N_5734,N_4880,N_3088);
nand U5735 (N_5735,N_3414,N_2448);
nand U5736 (N_5736,N_1433,N_4693);
nand U5737 (N_5737,N_1545,N_583);
or U5738 (N_5738,N_1009,N_1055);
nor U5739 (N_5739,N_2285,N_82);
or U5740 (N_5740,N_526,N_1860);
or U5741 (N_5741,N_1736,N_1583);
nand U5742 (N_5742,N_4121,N_793);
and U5743 (N_5743,N_2765,N_1046);
or U5744 (N_5744,N_1779,N_3009);
nor U5745 (N_5745,N_2282,N_1432);
and U5746 (N_5746,N_1328,N_584);
xnor U5747 (N_5747,N_3167,N_3523);
xnor U5748 (N_5748,N_4569,N_3154);
nand U5749 (N_5749,N_761,N_388);
nand U5750 (N_5750,N_1385,N_4171);
nor U5751 (N_5751,N_4975,N_1601);
or U5752 (N_5752,N_2998,N_1296);
or U5753 (N_5753,N_1904,N_4612);
and U5754 (N_5754,N_2725,N_796);
nand U5755 (N_5755,N_2662,N_2842);
or U5756 (N_5756,N_39,N_206);
or U5757 (N_5757,N_2995,N_2336);
and U5758 (N_5758,N_426,N_3556);
nor U5759 (N_5759,N_3077,N_46);
and U5760 (N_5760,N_2108,N_1204);
nand U5761 (N_5761,N_3572,N_638);
xnor U5762 (N_5762,N_2439,N_4127);
nand U5763 (N_5763,N_2732,N_1000);
xor U5764 (N_5764,N_853,N_2532);
nand U5765 (N_5765,N_3831,N_1987);
nand U5766 (N_5766,N_3538,N_211);
nor U5767 (N_5767,N_2923,N_4019);
or U5768 (N_5768,N_2861,N_1575);
xor U5769 (N_5769,N_3859,N_3897);
or U5770 (N_5770,N_3216,N_3686);
nor U5771 (N_5771,N_3331,N_4093);
and U5772 (N_5772,N_1423,N_3666);
xnor U5773 (N_5773,N_4870,N_7);
or U5774 (N_5774,N_4740,N_1040);
xnor U5775 (N_5775,N_1486,N_856);
nor U5776 (N_5776,N_4924,N_557);
or U5777 (N_5777,N_2605,N_3449);
nor U5778 (N_5778,N_4499,N_2627);
and U5779 (N_5779,N_1231,N_3067);
nor U5780 (N_5780,N_3836,N_4368);
or U5781 (N_5781,N_3473,N_1931);
and U5782 (N_5782,N_4983,N_2493);
nor U5783 (N_5783,N_2950,N_3793);
and U5784 (N_5784,N_3515,N_1143);
nand U5785 (N_5785,N_561,N_3382);
or U5786 (N_5786,N_2400,N_3242);
and U5787 (N_5787,N_2635,N_1212);
nor U5788 (N_5788,N_1435,N_2555);
or U5789 (N_5789,N_2877,N_4328);
and U5790 (N_5790,N_2221,N_2718);
and U5791 (N_5791,N_2825,N_1956);
nor U5792 (N_5792,N_350,N_4594);
and U5793 (N_5793,N_3896,N_2062);
and U5794 (N_5794,N_1830,N_1256);
nand U5795 (N_5795,N_3613,N_4046);
or U5796 (N_5796,N_238,N_175);
or U5797 (N_5797,N_3440,N_1676);
or U5798 (N_5798,N_2017,N_3739);
nand U5799 (N_5799,N_4057,N_1920);
nor U5800 (N_5800,N_437,N_971);
or U5801 (N_5801,N_1965,N_2561);
or U5802 (N_5802,N_809,N_1856);
nor U5803 (N_5803,N_4038,N_1790);
or U5804 (N_5804,N_3018,N_2566);
xnor U5805 (N_5805,N_4308,N_88);
xor U5806 (N_5806,N_2822,N_1875);
xnor U5807 (N_5807,N_1312,N_3279);
or U5808 (N_5808,N_753,N_279);
nand U5809 (N_5809,N_3386,N_2280);
and U5810 (N_5810,N_1554,N_2816);
nor U5811 (N_5811,N_360,N_1463);
and U5812 (N_5812,N_3096,N_2697);
nand U5813 (N_5813,N_1223,N_1049);
nand U5814 (N_5814,N_3192,N_4496);
and U5815 (N_5815,N_1228,N_4094);
nand U5816 (N_5816,N_3935,N_964);
nand U5817 (N_5817,N_2639,N_2688);
and U5818 (N_5818,N_3313,N_612);
or U5819 (N_5819,N_2851,N_1145);
xnor U5820 (N_5820,N_2559,N_2420);
nand U5821 (N_5821,N_1333,N_1192);
nand U5822 (N_5822,N_1932,N_3777);
nand U5823 (N_5823,N_1384,N_1485);
nor U5824 (N_5824,N_3612,N_2088);
and U5825 (N_5825,N_2912,N_1021);
nand U5826 (N_5826,N_4145,N_4141);
and U5827 (N_5827,N_203,N_4406);
nand U5828 (N_5828,N_2164,N_2274);
or U5829 (N_5829,N_2312,N_1467);
or U5830 (N_5830,N_2313,N_867);
nor U5831 (N_5831,N_1940,N_2512);
xor U5832 (N_5832,N_2455,N_1552);
xor U5833 (N_5833,N_1387,N_4015);
nor U5834 (N_5834,N_2499,N_441);
nand U5835 (N_5835,N_3348,N_256);
nand U5836 (N_5836,N_4699,N_656);
nand U5837 (N_5837,N_2460,N_903);
nand U5838 (N_5838,N_1284,N_929);
nand U5839 (N_5839,N_4808,N_4727);
nand U5840 (N_5840,N_3420,N_1966);
and U5841 (N_5841,N_3408,N_947);
xor U5842 (N_5842,N_501,N_148);
nor U5843 (N_5843,N_3092,N_851);
nand U5844 (N_5844,N_2325,N_2944);
xor U5845 (N_5845,N_47,N_269);
or U5846 (N_5846,N_3571,N_1011);
nor U5847 (N_5847,N_174,N_2634);
nor U5848 (N_5848,N_2114,N_2479);
nand U5849 (N_5849,N_3132,N_1489);
xnor U5850 (N_5850,N_1456,N_2866);
nand U5851 (N_5851,N_2002,N_2674);
xor U5852 (N_5852,N_2347,N_838);
or U5853 (N_5853,N_4863,N_2092);
or U5854 (N_5854,N_1246,N_3277);
nor U5855 (N_5855,N_1758,N_4354);
xor U5856 (N_5856,N_3962,N_2782);
xnor U5857 (N_5857,N_1627,N_3165);
or U5858 (N_5858,N_4942,N_3292);
and U5859 (N_5859,N_4348,N_2398);
nor U5860 (N_5860,N_3832,N_3059);
or U5861 (N_5861,N_865,N_4954);
and U5862 (N_5862,N_4995,N_1594);
nor U5863 (N_5863,N_3103,N_177);
nor U5864 (N_5864,N_2395,N_4761);
or U5865 (N_5865,N_489,N_2165);
or U5866 (N_5866,N_2323,N_2522);
nor U5867 (N_5867,N_4926,N_4279);
nor U5868 (N_5868,N_4018,N_2259);
xnor U5869 (N_5869,N_2549,N_2520);
nand U5870 (N_5870,N_2956,N_3111);
nand U5871 (N_5871,N_1657,N_3303);
or U5872 (N_5872,N_3871,N_2014);
nand U5873 (N_5873,N_3288,N_2234);
and U5874 (N_5874,N_344,N_2148);
or U5875 (N_5875,N_1983,N_4179);
or U5876 (N_5876,N_1731,N_4615);
or U5877 (N_5877,N_934,N_1128);
xnor U5878 (N_5878,N_43,N_3622);
and U5879 (N_5879,N_1573,N_3269);
nor U5880 (N_5880,N_757,N_1701);
or U5881 (N_5881,N_4210,N_4337);
or U5882 (N_5882,N_1673,N_2042);
xor U5883 (N_5883,N_4616,N_4676);
nor U5884 (N_5884,N_4217,N_532);
and U5885 (N_5885,N_1914,N_4176);
nor U5886 (N_5886,N_4631,N_748);
nor U5887 (N_5887,N_4541,N_1085);
nor U5888 (N_5888,N_3794,N_1934);
and U5889 (N_5889,N_4307,N_476);
nor U5890 (N_5890,N_3227,N_4030);
nand U5891 (N_5891,N_2072,N_715);
or U5892 (N_5892,N_3429,N_2778);
nor U5893 (N_5893,N_4016,N_2271);
and U5894 (N_5894,N_1449,N_4240);
or U5895 (N_5895,N_3849,N_4035);
and U5896 (N_5896,N_4401,N_4259);
nor U5897 (N_5897,N_3810,N_4461);
and U5898 (N_5898,N_3450,N_4303);
and U5899 (N_5899,N_3307,N_3948);
nand U5900 (N_5900,N_3047,N_4397);
or U5901 (N_5901,N_4369,N_3629);
xor U5902 (N_5902,N_2291,N_4840);
xnor U5903 (N_5903,N_3713,N_63);
xor U5904 (N_5904,N_444,N_1766);
or U5905 (N_5905,N_120,N_956);
xnor U5906 (N_5906,N_673,N_2711);
nor U5907 (N_5907,N_2831,N_1622);
nand U5908 (N_5908,N_963,N_2203);
or U5909 (N_5909,N_4648,N_4665);
and U5910 (N_5910,N_878,N_3608);
nor U5911 (N_5911,N_3668,N_4137);
xnor U5912 (N_5912,N_3156,N_1908);
nor U5913 (N_5913,N_795,N_79);
xnor U5914 (N_5914,N_917,N_1253);
nor U5915 (N_5915,N_2988,N_4707);
and U5916 (N_5916,N_4948,N_3099);
nor U5917 (N_5917,N_2507,N_255);
xnor U5918 (N_5918,N_264,N_2854);
or U5919 (N_5919,N_3692,N_1550);
or U5920 (N_5920,N_4908,N_668);
or U5921 (N_5921,N_2100,N_1053);
nand U5922 (N_5922,N_772,N_4161);
or U5923 (N_5923,N_542,N_771);
nor U5924 (N_5924,N_3511,N_3234);
or U5925 (N_5925,N_3830,N_875);
and U5926 (N_5926,N_994,N_2735);
nand U5927 (N_5927,N_2796,N_393);
xnor U5928 (N_5928,N_1527,N_1415);
nor U5929 (N_5929,N_3667,N_3147);
xnor U5930 (N_5930,N_4734,N_2830);
nand U5931 (N_5931,N_1052,N_628);
or U5932 (N_5932,N_525,N_3601);
and U5933 (N_5933,N_1123,N_2116);
and U5934 (N_5934,N_1897,N_1961);
nand U5935 (N_5935,N_4224,N_3342);
nor U5936 (N_5936,N_683,N_496);
or U5937 (N_5937,N_339,N_2564);
xnor U5938 (N_5938,N_3586,N_4006);
nand U5939 (N_5939,N_3539,N_1972);
nor U5940 (N_5940,N_2509,N_4559);
nor U5941 (N_5941,N_20,N_4894);
and U5942 (N_5942,N_4000,N_1465);
or U5943 (N_5943,N_2490,N_2286);
or U5944 (N_5944,N_1410,N_603);
nand U5945 (N_5945,N_2250,N_4059);
xnor U5946 (N_5946,N_623,N_2074);
and U5947 (N_5947,N_4591,N_1804);
and U5948 (N_5948,N_1301,N_3658);
nand U5949 (N_5949,N_712,N_1870);
nand U5950 (N_5950,N_1202,N_484);
xor U5951 (N_5951,N_104,N_3226);
nand U5952 (N_5952,N_3626,N_1710);
nand U5953 (N_5953,N_3814,N_2242);
nor U5954 (N_5954,N_2093,N_2124);
and U5955 (N_5955,N_469,N_1360);
nor U5956 (N_5956,N_4193,N_4010);
nor U5957 (N_5957,N_2755,N_4276);
nor U5958 (N_5958,N_4833,N_783);
and U5959 (N_5959,N_4935,N_2569);
or U5960 (N_5960,N_375,N_2552);
and U5961 (N_5961,N_531,N_1770);
and U5962 (N_5962,N_2867,N_2192);
or U5963 (N_5963,N_1472,N_278);
or U5964 (N_5964,N_3157,N_3996);
nand U5965 (N_5965,N_4753,N_3559);
and U5966 (N_5966,N_4031,N_3573);
xor U5967 (N_5967,N_2676,N_382);
nand U5968 (N_5968,N_3225,N_2550);
and U5969 (N_5969,N_3038,N_362);
nor U5970 (N_5970,N_2067,N_3915);
xnor U5971 (N_5971,N_803,N_3054);
xor U5972 (N_5972,N_220,N_2890);
or U5973 (N_5973,N_4964,N_4551);
nand U5974 (N_5974,N_4258,N_3528);
or U5975 (N_5975,N_1638,N_3945);
and U5976 (N_5976,N_644,N_4526);
nand U5977 (N_5977,N_2423,N_909);
xor U5978 (N_5978,N_3215,N_2918);
nor U5979 (N_5979,N_2656,N_4782);
nor U5980 (N_5980,N_2497,N_352);
xor U5981 (N_5981,N_3839,N_1498);
or U5982 (N_5982,N_2468,N_2913);
xnor U5983 (N_5983,N_3725,N_140);
nor U5984 (N_5984,N_2044,N_4689);
xor U5985 (N_5985,N_4110,N_820);
and U5986 (N_5986,N_3383,N_2139);
nand U5987 (N_5987,N_4860,N_4755);
nor U5988 (N_5988,N_486,N_3204);
nor U5989 (N_5989,N_3557,N_332);
nor U5990 (N_5990,N_4313,N_3044);
and U5991 (N_5991,N_1402,N_2763);
nand U5992 (N_5992,N_3387,N_3194);
xor U5993 (N_5993,N_4571,N_3434);
or U5994 (N_5994,N_3186,N_4177);
nand U5995 (N_5995,N_3843,N_4519);
nor U5996 (N_5996,N_407,N_3641);
xor U5997 (N_5997,N_4844,N_4427);
xnor U5998 (N_5998,N_3544,N_1030);
xnor U5999 (N_5999,N_3760,N_16);
and U6000 (N_6000,N_2167,N_1825);
or U6001 (N_6001,N_823,N_3209);
nor U6002 (N_6002,N_2144,N_2933);
or U6003 (N_6003,N_957,N_1963);
and U6004 (N_6004,N_420,N_2892);
xor U6005 (N_6005,N_1272,N_2582);
nand U6006 (N_6006,N_3647,N_1580);
nand U6007 (N_6007,N_1115,N_439);
and U6008 (N_6008,N_1278,N_2288);
xnor U6009 (N_6009,N_4823,N_785);
nor U6010 (N_6010,N_4039,N_3066);
and U6011 (N_6011,N_1014,N_3012);
nand U6012 (N_6012,N_2349,N_4436);
and U6013 (N_6013,N_3480,N_3672);
nor U6014 (N_6014,N_497,N_1029);
and U6015 (N_6015,N_152,N_3207);
nor U6016 (N_6016,N_210,N_1649);
nor U6017 (N_6017,N_310,N_655);
xnor U6018 (N_6018,N_3282,N_1938);
nor U6019 (N_6019,N_2739,N_1028);
nor U6020 (N_6020,N_4383,N_376);
nor U6021 (N_6021,N_227,N_1033);
or U6022 (N_6022,N_2187,N_2418);
xnor U6023 (N_6023,N_404,N_3910);
xor U6024 (N_6024,N_2871,N_1097);
or U6025 (N_6025,N_3616,N_4159);
nor U6026 (N_6026,N_4317,N_2331);
and U6027 (N_6027,N_1368,N_2857);
nor U6028 (N_6028,N_2473,N_370);
or U6029 (N_6029,N_2050,N_1293);
nor U6030 (N_6030,N_3801,N_2391);
or U6031 (N_6031,N_2428,N_4451);
xor U6032 (N_6032,N_473,N_4508);
and U6033 (N_6033,N_1137,N_4207);
xor U6034 (N_6034,N_2802,N_1343);
or U6035 (N_6035,N_2402,N_3016);
nor U6036 (N_6036,N_662,N_1564);
nand U6037 (N_6037,N_3909,N_3791);
nor U6038 (N_6038,N_4498,N_2961);
or U6039 (N_6039,N_2489,N_4241);
nor U6040 (N_6040,N_3705,N_4322);
nand U6041 (N_6041,N_447,N_3025);
nor U6042 (N_6042,N_4156,N_1767);
nor U6043 (N_6043,N_3804,N_3052);
nand U6044 (N_6044,N_3941,N_1464);
and U6045 (N_6045,N_351,N_4189);
xnor U6046 (N_6046,N_2864,N_5);
nand U6047 (N_6047,N_3687,N_2035);
and U6048 (N_6048,N_4901,N_98);
or U6049 (N_6049,N_3546,N_3289);
nand U6050 (N_6050,N_4070,N_1382);
nand U6051 (N_6051,N_122,N_3189);
and U6052 (N_6052,N_341,N_2220);
and U6053 (N_6053,N_1913,N_3197);
and U6054 (N_6054,N_3599,N_635);
xnor U6055 (N_6055,N_4893,N_819);
and U6056 (N_6056,N_3290,N_3600);
and U6057 (N_6057,N_2638,N_4147);
nor U6058 (N_6058,N_1357,N_2132);
nor U6059 (N_6059,N_1789,N_0);
xnor U6060 (N_6060,N_1584,N_4680);
nand U6061 (N_6061,N_3585,N_2115);
xnor U6062 (N_6062,N_579,N_215);
nor U6063 (N_6063,N_364,N_3792);
or U6064 (N_6064,N_3246,N_1116);
or U6065 (N_6065,N_2740,N_2760);
and U6066 (N_6066,N_22,N_84);
nor U6067 (N_6067,N_4103,N_1148);
or U6068 (N_6068,N_3499,N_2889);
xor U6069 (N_6069,N_4846,N_113);
nor U6070 (N_6070,N_4702,N_4390);
nand U6071 (N_6071,N_3114,N_421);
or U6072 (N_6072,N_2324,N_4758);
xor U6073 (N_6073,N_4220,N_4434);
or U6074 (N_6074,N_1454,N_3554);
and U6075 (N_6075,N_3028,N_4514);
and U6076 (N_6076,N_4237,N_1022);
or U6077 (N_6077,N_3299,N_2722);
nand U6078 (N_6078,N_3718,N_1413);
or U6079 (N_6079,N_249,N_1501);
nor U6080 (N_6080,N_4632,N_286);
nand U6081 (N_6081,N_288,N_619);
nor U6082 (N_6082,N_2780,N_323);
xnor U6083 (N_6083,N_4723,N_4285);
and U6084 (N_6084,N_2932,N_3532);
and U6085 (N_6085,N_1407,N_2410);
nor U6086 (N_6086,N_4976,N_2984);
and U6087 (N_6087,N_4075,N_1708);
and U6088 (N_6088,N_4041,N_2268);
or U6089 (N_6089,N_4824,N_4933);
xnor U6090 (N_6090,N_358,N_165);
or U6091 (N_6091,N_3570,N_999);
xnor U6092 (N_6092,N_101,N_333);
nand U6093 (N_6093,N_839,N_2751);
nor U6094 (N_6094,N_1683,N_383);
and U6095 (N_6095,N_1582,N_4618);
or U6096 (N_6096,N_4611,N_1084);
nor U6097 (N_6097,N_3563,N_3115);
and U6098 (N_6098,N_338,N_536);
or U6099 (N_6099,N_4656,N_4040);
nor U6100 (N_6100,N_3349,N_3966);
nor U6101 (N_6101,N_2081,N_4826);
nor U6102 (N_6102,N_3490,N_2076);
nand U6103 (N_6103,N_4558,N_908);
and U6104 (N_6104,N_3393,N_3244);
and U6105 (N_6105,N_1630,N_4597);
nor U6106 (N_6106,N_3168,N_3822);
or U6107 (N_6107,N_2715,N_2888);
nand U6108 (N_6108,N_2204,N_634);
xor U6109 (N_6109,N_1728,N_1980);
nor U6110 (N_6110,N_4486,N_4232);
nor U6111 (N_6111,N_450,N_2575);
nor U6112 (N_6112,N_3229,N_1532);
nor U6113 (N_6113,N_334,N_1678);
nand U6114 (N_6114,N_3448,N_425);
or U6115 (N_6115,N_4847,N_822);
and U6116 (N_6116,N_1930,N_1985);
or U6117 (N_6117,N_1801,N_4626);
nand U6118 (N_6118,N_3838,N_4260);
or U6119 (N_6119,N_4649,N_3844);
and U6120 (N_6120,N_3778,N_3085);
xnor U6121 (N_6121,N_744,N_4221);
and U6122 (N_6122,N_4142,N_2486);
or U6123 (N_6123,N_3740,N_4907);
or U6124 (N_6124,N_4048,N_943);
nand U6125 (N_6125,N_318,N_2459);
nor U6126 (N_6126,N_2354,N_1041);
nand U6127 (N_6127,N_682,N_2937);
or U6128 (N_6128,N_4822,N_4334);
nor U6129 (N_6129,N_2090,N_2756);
xnor U6130 (N_6130,N_4225,N_610);
xor U6131 (N_6131,N_2028,N_141);
nand U6132 (N_6132,N_259,N_3669);
xor U6133 (N_6133,N_3582,N_2049);
nor U6134 (N_6134,N_3706,N_2623);
and U6135 (N_6135,N_1114,N_2774);
xnor U6136 (N_6136,N_4807,N_1933);
and U6137 (N_6137,N_226,N_770);
or U6138 (N_6138,N_833,N_3661);
nand U6139 (N_6139,N_2366,N_3755);
or U6140 (N_6140,N_3889,N_877);
or U6141 (N_6141,N_4343,N_1455);
or U6142 (N_6142,N_1891,N_3698);
nor U6143 (N_6143,N_1883,N_1866);
or U6144 (N_6144,N_2959,N_2446);
xnor U6145 (N_6145,N_1973,N_4659);
or U6146 (N_6146,N_3469,N_2018);
xor U6147 (N_6147,N_4314,N_528);
nand U6148 (N_6148,N_3093,N_1540);
and U6149 (N_6149,N_45,N_3328);
xnor U6150 (N_6150,N_2632,N_692);
nand U6151 (N_6151,N_3971,N_3471);
nor U6152 (N_6152,N_3320,N_3502);
and U6153 (N_6153,N_955,N_1659);
or U6154 (N_6154,N_3723,N_2123);
or U6155 (N_6155,N_2953,N_2444);
and U6156 (N_6156,N_3808,N_1865);
and U6157 (N_6157,N_1648,N_1528);
and U6158 (N_6158,N_1699,N_3343);
nand U6159 (N_6159,N_2754,N_1924);
xnor U6160 (N_6160,N_1822,N_1493);
nand U6161 (N_6161,N_3604,N_4459);
nor U6162 (N_6162,N_3541,N_2106);
and U6163 (N_6163,N_1314,N_3027);
and U6164 (N_6164,N_1469,N_2233);
and U6165 (N_6165,N_475,N_2117);
nor U6166 (N_6166,N_3766,N_4745);
nor U6167 (N_6167,N_2683,N_2810);
nor U6168 (N_6168,N_2105,N_4181);
and U6169 (N_6169,N_1249,N_4529);
nand U6170 (N_6170,N_2749,N_4695);
nor U6171 (N_6171,N_1916,N_2599);
or U6172 (N_6172,N_2005,N_3591);
or U6173 (N_6173,N_2258,N_4938);
and U6174 (N_6174,N_1285,N_2805);
xor U6175 (N_6175,N_3757,N_2742);
nand U6176 (N_6176,N_1290,N_997);
xnor U6177 (N_6177,N_4388,N_2294);
nor U6178 (N_6178,N_1579,N_2695);
nor U6179 (N_6179,N_4076,N_2746);
or U6180 (N_6180,N_4435,N_2863);
nor U6181 (N_6181,N_44,N_3765);
or U6182 (N_6182,N_2929,N_2208);
nand U6183 (N_6183,N_4,N_488);
and U6184 (N_6184,N_830,N_3685);
nor U6185 (N_6185,N_866,N_2247);
nand U6186 (N_6186,N_2085,N_1687);
or U6187 (N_6187,N_3516,N_1746);
and U6188 (N_6188,N_1840,N_792);
nor U6189 (N_6189,N_4633,N_3526);
or U6190 (N_6190,N_2546,N_659);
nand U6191 (N_6191,N_2666,N_2214);
or U6192 (N_6192,N_2064,N_296);
or U6193 (N_6193,N_3451,N_3217);
xor U6194 (N_6194,N_3917,N_2531);
or U6195 (N_6195,N_4195,N_2077);
xnor U6196 (N_6196,N_3174,N_303);
and U6197 (N_6197,N_627,N_558);
xnor U6198 (N_6198,N_3679,N_1591);
and U6199 (N_6199,N_4671,N_657);
and U6200 (N_6200,N_2758,N_2790);
xnor U6201 (N_6201,N_4784,N_1944);
nor U6202 (N_6202,N_15,N_2542);
nor U6203 (N_6203,N_3664,N_3504);
nor U6204 (N_6204,N_4109,N_4851);
or U6205 (N_6205,N_494,N_4575);
xor U6206 (N_6206,N_4490,N_3351);
xor U6207 (N_6207,N_2059,N_3144);
nor U6208 (N_6208,N_2829,N_3152);
nor U6209 (N_6209,N_643,N_3547);
and U6210 (N_6210,N_3125,N_1951);
nand U6211 (N_6211,N_2704,N_3042);
and U6212 (N_6212,N_1734,N_1723);
xor U6213 (N_6213,N_3247,N_1823);
or U6214 (N_6214,N_1186,N_247);
nor U6215 (N_6215,N_918,N_4560);
and U6216 (N_6216,N_4516,N_4423);
or U6217 (N_6217,N_1763,N_4589);
nor U6218 (N_6218,N_3080,N_4704);
and U6219 (N_6219,N_2919,N_4405);
xnor U6220 (N_6220,N_1142,N_130);
xnor U6221 (N_6221,N_3369,N_1179);
and U6222 (N_6222,N_3437,N_200);
nand U6223 (N_6223,N_2526,N_4344);
xnor U6224 (N_6224,N_2818,N_3746);
xnor U6225 (N_6225,N_2029,N_794);
or U6226 (N_6226,N_4466,N_3590);
nor U6227 (N_6227,N_2249,N_4709);
and U6228 (N_6228,N_2175,N_2680);
nand U6229 (N_6229,N_1563,N_4750);
xnor U6230 (N_6230,N_2104,N_939);
nor U6231 (N_6231,N_4113,N_4735);
xor U6232 (N_6232,N_3191,N_3874);
xnor U6233 (N_6233,N_4086,N_4977);
xor U6234 (N_6234,N_4653,N_2120);
nor U6235 (N_6235,N_2201,N_85);
and U6236 (N_6236,N_1715,N_3627);
nand U6237 (N_6237,N_4877,N_4771);
and U6238 (N_6238,N_3086,N_1063);
or U6239 (N_6239,N_1529,N_385);
nand U6240 (N_6240,N_3800,N_2513);
nor U6241 (N_6241,N_1751,N_4082);
xnor U6242 (N_6242,N_4081,N_4411);
nor U6243 (N_6243,N_1886,N_50);
nand U6244 (N_6244,N_4791,N_2021);
or U6245 (N_6245,N_4003,N_4359);
and U6246 (N_6246,N_2134,N_2058);
or U6247 (N_6247,N_813,N_491);
and U6248 (N_6248,N_4301,N_477);
xor U6249 (N_6249,N_1088,N_3855);
xor U6250 (N_6250,N_446,N_594);
nor U6251 (N_6251,N_4585,N_2874);
nor U6252 (N_6252,N_112,N_3357);
nor U6253 (N_6253,N_3826,N_4802);
xor U6254 (N_6254,N_1017,N_2883);
or U6255 (N_6255,N_77,N_2727);
nor U6256 (N_6256,N_4785,N_551);
nand U6257 (N_6257,N_3388,N_3489);
nor U6258 (N_6258,N_3933,N_2156);
and U6259 (N_6259,N_1879,N_973);
nand U6260 (N_6260,N_3245,N_4737);
xor U6261 (N_6261,N_873,N_4621);
or U6262 (N_6262,N_1576,N_640);
and U6263 (N_6263,N_4500,N_4639);
and U6264 (N_6264,N_1470,N_2481);
or U6265 (N_6265,N_2583,N_811);
and U6266 (N_6266,N_514,N_2405);
nand U6267 (N_6267,N_2122,N_716);
and U6268 (N_6268,N_251,N_356);
xnor U6269 (N_6269,N_2154,N_3790);
or U6270 (N_6270,N_4077,N_4876);
nand U6271 (N_6271,N_3163,N_3876);
or U6272 (N_6272,N_3285,N_4339);
or U6273 (N_6273,N_3595,N_1187);
or U6274 (N_6274,N_2121,N_3982);
nor U6275 (N_6275,N_1611,N_3989);
and U6276 (N_6276,N_1072,N_2270);
xor U6277 (N_6277,N_1111,N_2174);
nor U6278 (N_6278,N_2495,N_1440);
xor U6279 (N_6279,N_4032,N_3110);
and U6280 (N_6280,N_2591,N_3719);
nor U6281 (N_6281,N_3465,N_158);
nor U6282 (N_6282,N_2303,N_4661);
xnor U6283 (N_6283,N_3254,N_3628);
nand U6284 (N_6284,N_3947,N_3598);
nand U6285 (N_6285,N_1405,N_1815);
nand U6286 (N_6286,N_3399,N_3363);
xor U6287 (N_6287,N_2352,N_1419);
or U6288 (N_6288,N_3079,N_4562);
nor U6289 (N_6289,N_569,N_3597);
xnor U6290 (N_6290,N_709,N_2502);
nor U6291 (N_6291,N_216,N_4582);
nor U6292 (N_6292,N_1505,N_2185);
nor U6293 (N_6293,N_244,N_4841);
or U6294 (N_6294,N_2795,N_898);
or U6295 (N_6295,N_4722,N_4512);
nor U6296 (N_6296,N_2975,N_2799);
or U6297 (N_6297,N_1010,N_3638);
or U6298 (N_6298,N_3049,N_4296);
nor U6299 (N_6299,N_413,N_2284);
nand U6300 (N_6300,N_4899,N_2057);
and U6301 (N_6301,N_3134,N_3175);
or U6302 (N_6302,N_4746,N_2437);
nor U6303 (N_6303,N_394,N_519);
nor U6304 (N_6304,N_2006,N_4678);
xor U6305 (N_6305,N_4100,N_2008);
xnor U6306 (N_6306,N_2603,N_3356);
and U6307 (N_6307,N_4509,N_1829);
and U6308 (N_6308,N_2999,N_153);
and U6309 (N_6309,N_1193,N_144);
and U6310 (N_6310,N_2411,N_1245);
nand U6311 (N_6311,N_4373,N_3753);
nor U6312 (N_6312,N_151,N_2474);
nor U6313 (N_6313,N_2511,N_836);
or U6314 (N_6314,N_2094,N_1688);
and U6315 (N_6315,N_4535,N_4460);
xnor U6316 (N_6316,N_1887,N_1992);
nor U6317 (N_6317,N_1417,N_4915);
nand U6318 (N_6318,N_4651,N_1628);
nor U6319 (N_6319,N_3514,N_642);
nand U6320 (N_6320,N_423,N_2048);
nand U6321 (N_6321,N_2619,N_900);
nor U6322 (N_6322,N_2445,N_4054);
and U6323 (N_6323,N_3398,N_4209);
nand U6324 (N_6324,N_2902,N_78);
xor U6325 (N_6325,N_2217,N_503);
or U6326 (N_6326,N_2246,N_4660);
xor U6327 (N_6327,N_4072,N_2281);
or U6328 (N_6328,N_844,N_3100);
nor U6329 (N_6329,N_1491,N_3634);
xnor U6330 (N_6330,N_4152,N_297);
nor U6331 (N_6331,N_3505,N_3729);
and U6332 (N_6332,N_4249,N_523);
and U6333 (N_6333,N_911,N_2587);
and U6334 (N_6334,N_3712,N_1654);
and U6335 (N_6335,N_4056,N_3250);
nand U6336 (N_6336,N_4329,N_4255);
or U6337 (N_6337,N_3993,N_1139);
nand U6338 (N_6338,N_4951,N_3263);
xnor U6339 (N_6339,N_1792,N_2452);
nor U6340 (N_6340,N_4391,N_1511);
and U6341 (N_6341,N_2724,N_3775);
and U6342 (N_6342,N_427,N_4859);
and U6343 (N_6343,N_4281,N_1957);
xnor U6344 (N_6344,N_3046,N_24);
and U6345 (N_6345,N_4362,N_4540);
nor U6346 (N_6346,N_1399,N_1745);
xnor U6347 (N_6347,N_2330,N_1784);
or U6348 (N_6348,N_2118,N_1392);
or U6349 (N_6349,N_4174,N_1292);
nor U6350 (N_6350,N_3743,N_1266);
xnor U6351 (N_6351,N_1076,N_746);
nor U6352 (N_6352,N_4380,N_4990);
nor U6353 (N_6353,N_4309,N_3138);
or U6354 (N_6354,N_3938,N_1609);
and U6355 (N_6355,N_4815,N_3439);
nor U6356 (N_6356,N_4849,N_1776);
and U6357 (N_6357,N_1533,N_2180);
or U6358 (N_6358,N_4732,N_2707);
or U6359 (N_6359,N_4440,N_765);
nand U6360 (N_6360,N_2978,N_843);
xnor U6361 (N_6361,N_1431,N_4421);
or U6362 (N_6362,N_2305,N_2300);
xnor U6363 (N_6363,N_1869,N_1826);
and U6364 (N_6364,N_4358,N_3494);
and U6365 (N_6365,N_4119,N_3730);
xor U6366 (N_6366,N_3653,N_4998);
xnor U6367 (N_6367,N_1768,N_3965);
nand U6368 (N_6368,N_538,N_3983);
or U6369 (N_6369,N_4520,N_2080);
and U6370 (N_6370,N_3654,N_543);
nor U6371 (N_6371,N_2943,N_2836);
or U6372 (N_6372,N_1889,N_4134);
and U6373 (N_6373,N_1876,N_4379);
nand U6374 (N_6374,N_4781,N_4349);
nand U6375 (N_6375,N_90,N_3180);
xnor U6376 (N_6376,N_4635,N_3976);
and U6377 (N_6377,N_2341,N_3396);
or U6378 (N_6378,N_1499,N_137);
nand U6379 (N_6379,N_4959,N_3994);
or U6380 (N_6380,N_3231,N_1780);
xnor U6381 (N_6381,N_4392,N_1713);
or U6382 (N_6382,N_3260,N_2611);
nor U6383 (N_6383,N_2394,N_4836);
xor U6384 (N_6384,N_3248,N_1837);
or U6385 (N_6385,N_2315,N_1158);
or U6386 (N_6386,N_1744,N_448);
xnor U6387 (N_6387,N_1984,N_3139);
nor U6388 (N_6388,N_2256,N_4608);
xnor U6389 (N_6389,N_4557,N_3574);
and U6390 (N_6390,N_3503,N_2942);
and U6391 (N_6391,N_921,N_2195);
nor U6392 (N_6392,N_461,N_4374);
and U6393 (N_6393,N_3459,N_212);
nor U6394 (N_6394,N_2885,N_2537);
or U6395 (N_6395,N_4023,N_859);
xnor U6396 (N_6396,N_4588,N_1602);
xor U6397 (N_6397,N_2417,N_3173);
and U6398 (N_6398,N_1795,N_4605);
or U6399 (N_6399,N_4960,N_2809);
and U6400 (N_6400,N_4952,N_2384);
nand U6401 (N_6401,N_1268,N_106);
nand U6402 (N_6402,N_3959,N_3964);
or U6403 (N_6403,N_3196,N_3149);
xor U6404 (N_6404,N_1424,N_618);
and U6405 (N_6405,N_4182,N_487);
or U6406 (N_6406,N_3893,N_2745);
nor U6407 (N_6407,N_3298,N_1339);
nor U6408 (N_6408,N_3581,N_54);
and U6409 (N_6409,N_3276,N_4741);
or U6410 (N_6410,N_3540,N_1140);
or U6411 (N_6411,N_4767,N_443);
nand U6412 (N_6412,N_2340,N_2030);
xor U6413 (N_6413,N_1124,N_1958);
and U6414 (N_6414,N_4278,N_725);
nand U6415 (N_6415,N_996,N_1073);
or U6416 (N_6416,N_3470,N_1468);
nor U6417 (N_6417,N_4151,N_1969);
nand U6418 (N_6418,N_3329,N_2098);
and U6419 (N_6419,N_67,N_706);
or U6420 (N_6420,N_3558,N_2514);
and U6421 (N_6421,N_510,N_4292);
or U6422 (N_6422,N_904,N_1131);
nand U6423 (N_6423,N_4211,N_3507);
nand U6424 (N_6424,N_2916,N_2155);
xor U6425 (N_6425,N_4300,N_1377);
and U6426 (N_6426,N_4879,N_982);
nand U6427 (N_6427,N_2589,N_4172);
nand U6428 (N_6428,N_161,N_2904);
nor U6429 (N_6429,N_35,N_2628);
and U6430 (N_6430,N_1551,N_1416);
nor U6431 (N_6431,N_2981,N_3662);
or U6432 (N_6432,N_378,N_3029);
xnor U6433 (N_6433,N_316,N_3105);
or U6434 (N_6434,N_3143,N_3758);
and U6435 (N_6435,N_2153,N_4623);
and U6436 (N_6436,N_2723,N_1332);
or U6437 (N_6437,N_3391,N_2505);
nor U6438 (N_6438,N_3340,N_3708);
xnor U6439 (N_6439,N_3764,N_845);
nor U6440 (N_6440,N_354,N_3835);
nor U6441 (N_6441,N_1986,N_1086);
nand U6442 (N_6442,N_3850,N_4290);
xnor U6443 (N_6443,N_2629,N_1521);
xor U6444 (N_6444,N_732,N_2614);
nor U6445 (N_6445,N_2240,N_4742);
and U6446 (N_6446,N_4034,N_2161);
nand U6447 (N_6447,N_852,N_1669);
nand U6448 (N_6448,N_2820,N_3824);
or U6449 (N_6449,N_4331,N_3642);
xor U6450 (N_6450,N_4792,N_4778);
nor U6451 (N_6451,N_3310,N_2702);
and U6452 (N_6452,N_4468,N_3695);
nand U6453 (N_6453,N_4720,N_633);
xnor U6454 (N_6454,N_3745,N_750);
nand U6455 (N_6455,N_395,N_4940);
xnor U6456 (N_6456,N_1998,N_1156);
and U6457 (N_6457,N_2147,N_192);
nand U6458 (N_6458,N_797,N_2202);
nor U6459 (N_6459,N_4202,N_577);
or U6460 (N_6460,N_2811,N_1662);
xnor U6461 (N_6461,N_4289,N_2733);
nand U6462 (N_6462,N_1703,N_4047);
nor U6463 (N_6463,N_4375,N_751);
nor U6464 (N_6464,N_4679,N_3026);
nand U6465 (N_6465,N_2527,N_217);
nand U6466 (N_6466,N_3636,N_1240);
or U6467 (N_6467,N_4855,N_1175);
nand U6468 (N_6468,N_4414,N_4409);
or U6469 (N_6469,N_4663,N_3312);
and U6470 (N_6470,N_4002,N_3205);
or U6471 (N_6471,N_3419,N_1042);
nor U6472 (N_6472,N_3252,N_3961);
and U6473 (N_6473,N_3400,N_3198);
and U6474 (N_6474,N_3339,N_3717);
xor U6475 (N_6475,N_3474,N_2644);
or U6476 (N_6476,N_449,N_857);
xnor U6477 (N_6477,N_2576,N_4637);
and U6478 (N_6478,N_3771,N_3118);
and U6479 (N_6479,N_1539,N_3272);
xor U6480 (N_6480,N_4123,N_4834);
and U6481 (N_6481,N_2839,N_4850);
xor U6482 (N_6482,N_3817,N_1096);
nand U6483 (N_6483,N_972,N_481);
xor U6484 (N_6484,N_2738,N_2397);
or U6485 (N_6485,N_3754,N_2158);
or U6486 (N_6486,N_1050,N_3525);
nand U6487 (N_6487,N_2222,N_3472);
and U6488 (N_6488,N_527,N_4454);
xnor U6489 (N_6489,N_1968,N_1422);
nor U6490 (N_6490,N_2669,N_277);
and U6491 (N_6491,N_3870,N_2053);
nor U6492 (N_6492,N_2881,N_1737);
nor U6493 (N_6493,N_4567,N_1900);
or U6494 (N_6494,N_60,N_1132);
nor U6495 (N_6495,N_4270,N_2523);
or U6496 (N_6496,N_752,N_2467);
and U6497 (N_6497,N_3562,N_766);
or U6498 (N_6498,N_1843,N_3177);
xnor U6499 (N_6499,N_3468,N_2000);
or U6500 (N_6500,N_304,N_3481);
nand U6501 (N_6501,N_776,N_2893);
nor U6502 (N_6502,N_1616,N_3353);
and U6503 (N_6503,N_233,N_4265);
nand U6504 (N_6504,N_812,N_1786);
nor U6505 (N_6505,N_69,N_4867);
nor U6506 (N_6506,N_2070,N_906);
xnor U6507 (N_6507,N_4909,N_2786);
xor U6508 (N_6508,N_549,N_371);
xnor U6509 (N_6509,N_3015,N_593);
nand U6510 (N_6510,N_1437,N_4384);
nand U6511 (N_6511,N_2252,N_4592);
nor U6512 (N_6512,N_265,N_3336);
or U6513 (N_6513,N_2873,N_2853);
nand U6514 (N_6514,N_979,N_1561);
nor U6515 (N_6515,N_3785,N_3206);
nor U6516 (N_6516,N_2712,N_2063);
or U6517 (N_6517,N_168,N_83);
and U6518 (N_6518,N_4580,N_397);
or U6519 (N_6519,N_2859,N_2267);
or U6520 (N_6520,N_827,N_309);
or U6521 (N_6521,N_4216,N_2168);
and U6522 (N_6522,N_4897,N_1306);
or U6523 (N_6523,N_3315,N_2539);
nand U6524 (N_6524,N_1639,N_258);
nand U6525 (N_6525,N_1418,N_2753);
nand U6526 (N_6526,N_27,N_2613);
and U6527 (N_6527,N_3884,N_1232);
or U6528 (N_6528,N_1149,N_890);
nand U6529 (N_6529,N_103,N_239);
nand U6530 (N_6530,N_4947,N_1759);
xor U6531 (N_6531,N_965,N_3091);
nand U6532 (N_6532,N_1679,N_3036);
xnor U6533 (N_6533,N_319,N_1711);
and U6534 (N_6534,N_4902,N_406);
nor U6535 (N_6535,N_2131,N_2529);
and U6536 (N_6536,N_438,N_1523);
xor U6537 (N_6537,N_4852,N_816);
or U6538 (N_6538,N_4768,N_1259);
xor U6539 (N_6539,N_4136,N_2664);
or U6540 (N_6540,N_2636,N_3319);
nor U6541 (N_6541,N_2690,N_863);
xor U6542 (N_6542,N_4312,N_3779);
xnor U6543 (N_6543,N_1363,N_1518);
xor U6544 (N_6544,N_3064,N_4729);
nand U6545 (N_6545,N_4667,N_3772);
xnor U6546 (N_6546,N_1781,N_4062);
xnor U6547 (N_6547,N_2066,N_807);
nand U6548 (N_6548,N_3452,N_432);
and U6549 (N_6549,N_4302,N_205);
xnor U6550 (N_6550,N_3621,N_884);
or U6551 (N_6551,N_209,N_111);
or U6552 (N_6552,N_36,N_196);
and U6553 (N_6553,N_2435,N_4553);
xnor U6554 (N_6554,N_1126,N_2211);
nor U6555 (N_6555,N_2150,N_4790);
nand U6556 (N_6556,N_2647,N_2844);
nand U6557 (N_6557,N_511,N_4800);
and U6558 (N_6558,N_2403,N_2798);
or U6559 (N_6559,N_1044,N_1936);
nand U6560 (N_6560,N_4239,N_698);
nor U6561 (N_6561,N_848,N_3645);
or U6562 (N_6562,N_322,N_4810);
nand U6563 (N_6563,N_535,N_97);
or U6564 (N_6564,N_1078,N_229);
xor U6565 (N_6565,N_2255,N_1167);
and U6566 (N_6566,N_1247,N_2357);
nor U6567 (N_6567,N_3140,N_1556);
and U6568 (N_6568,N_197,N_1389);
or U6569 (N_6569,N_3423,N_948);
or U6570 (N_6570,N_37,N_3034);
xnor U6571 (N_6571,N_451,N_615);
and U6572 (N_6572,N_4386,N_3179);
xnor U6573 (N_6573,N_4916,N_4385);
xor U6574 (N_6574,N_2130,N_861);
and U6575 (N_6575,N_4025,N_1948);
xnor U6576 (N_6576,N_2812,N_1839);
nand U6577 (N_6577,N_3199,N_3475);
or U6578 (N_6578,N_888,N_4487);
nor U6579 (N_6579,N_954,N_2299);
or U6580 (N_6580,N_74,N_2266);
nor U6581 (N_6581,N_3690,N_4603);
nor U6582 (N_6582,N_4949,N_4116);
or U6583 (N_6583,N_2840,N_1338);
or U6584 (N_6584,N_516,N_4596);
and U6585 (N_6585,N_524,N_1199);
nor U6586 (N_6586,N_4923,N_4345);
nand U6587 (N_6587,N_1446,N_541);
and U6588 (N_6588,N_4227,N_1005);
nand U6589 (N_6589,N_3050,N_2621);
and U6590 (N_6590,N_2374,N_472);
nand U6591 (N_6591,N_4604,N_775);
or U6592 (N_6592,N_325,N_4361);
xnor U6593 (N_6593,N_1177,N_390);
nor U6594 (N_6594,N_835,N_4212);
or U6595 (N_6595,N_23,N_1513);
and U6596 (N_6596,N_2133,N_1380);
and U6597 (N_6597,N_3251,N_2311);
xor U6598 (N_6598,N_1834,N_2068);
nor U6599 (N_6599,N_4817,N_1219);
or U6600 (N_6600,N_3255,N_2193);
or U6601 (N_6601,N_4576,N_1566);
or U6602 (N_6602,N_3477,N_125);
xor U6603 (N_6603,N_2602,N_4917);
xnor U6604 (N_6604,N_4657,N_1667);
nand U6605 (N_6605,N_938,N_2622);
nor U6606 (N_6606,N_1633,N_2646);
nand U6607 (N_6607,N_2671,N_1133);
xor U6608 (N_6608,N_2264,N_4257);
and U6609 (N_6609,N_4107,N_788);
nor U6610 (N_6610,N_1264,N_1682);
nor U6611 (N_6611,N_4646,N_3928);
and U6612 (N_6612,N_4170,N_3607);
nor U6613 (N_6613,N_436,N_275);
and U6614 (N_6614,N_2730,N_4360);
nor U6615 (N_6615,N_3361,N_2951);
nand U6616 (N_6616,N_3926,N_324);
and U6617 (N_6617,N_1730,N_3560);
or U6618 (N_6618,N_4590,N_810);
nor U6619 (N_6619,N_1397,N_142);
nand U6620 (N_6620,N_801,N_4140);
or U6621 (N_6621,N_3335,N_3200);
or U6622 (N_6622,N_554,N_4458);
nand U6623 (N_6623,N_1165,N_1113);
and U6624 (N_6624,N_4882,N_1756);
nand U6625 (N_6625,N_4053,N_3980);
or U6626 (N_6626,N_1670,N_219);
nand U6627 (N_6627,N_2113,N_4264);
xnor U6628 (N_6628,N_4992,N_1910);
and U6629 (N_6629,N_978,N_944);
nor U6630 (N_6630,N_1238,N_2921);
or U6631 (N_6631,N_4364,N_907);
or U6632 (N_6632,N_1401,N_2241);
and U6633 (N_6633,N_1748,N_3164);
or U6634 (N_6634,N_4323,N_1941);
nand U6635 (N_6635,N_1283,N_849);
xnor U6636 (N_6636,N_4215,N_1185);
and U6637 (N_6637,N_887,N_4752);
xnor U6638 (N_6638,N_2236,N_1512);
or U6639 (N_6639,N_509,N_359);
nand U6640 (N_6640,N_418,N_2869);
nand U6641 (N_6641,N_1309,N_4389);
nor U6642 (N_6642,N_550,N_902);
or U6643 (N_6643,N_3076,N_377);
and U6644 (N_6644,N_306,N_4625);
and U6645 (N_6645,N_3852,N_2321);
xor U6646 (N_6646,N_679,N_466);
or U6647 (N_6647,N_2290,N_4685);
nand U6648 (N_6648,N_4819,N_246);
or U6649 (N_6649,N_641,N_3403);
xor U6650 (N_6650,N_4118,N_2958);
nand U6651 (N_6651,N_3330,N_135);
and U6652 (N_6652,N_4432,N_3354);
and U6653 (N_6653,N_3213,N_3286);
xor U6654 (N_6654,N_3553,N_566);
or U6655 (N_6655,N_1660,N_4736);
nor U6656 (N_6656,N_3742,N_2652);
and U6657 (N_6657,N_2766,N_2389);
nor U6658 (N_6658,N_2334,N_53);
or U6659 (N_6659,N_2592,N_563);
or U6660 (N_6660,N_1760,N_1411);
nor U6661 (N_6661,N_4098,N_1813);
xor U6662 (N_6662,N_3131,N_3682);
or U6663 (N_6663,N_1783,N_767);
xnor U6664 (N_6664,N_1492,N_2160);
nand U6665 (N_6665,N_977,N_3820);
or U6666 (N_6666,N_100,N_2585);
nand U6667 (N_6667,N_976,N_2179);
and U6668 (N_6668,N_64,N_4674);
nand U6669 (N_6669,N_1320,N_1200);
xor U6670 (N_6670,N_201,N_1300);
xor U6671 (N_6671,N_2358,N_1108);
xor U6672 (N_6672,N_3735,N_3862);
and U6673 (N_6673,N_829,N_3425);
and U6674 (N_6674,N_2641,N_4416);
nand U6675 (N_6675,N_3985,N_2456);
xor U6676 (N_6676,N_2604,N_162);
xor U6677 (N_6677,N_2182,N_3724);
and U6678 (N_6678,N_2099,N_4681);
nand U6679 (N_6679,N_4532,N_169);
nor U6680 (N_6680,N_3136,N_3578);
nand U6681 (N_6681,N_4341,N_1428);
xor U6682 (N_6682,N_1982,N_3811);
or U6683 (N_6683,N_1425,N_117);
or U6684 (N_6684,N_2335,N_4507);
and U6685 (N_6685,N_4524,N_1340);
nand U6686 (N_6686,N_4690,N_457);
xnor U6687 (N_6687,N_410,N_3914);
or U6688 (N_6688,N_4298,N_3731);
and U6689 (N_6689,N_3569,N_3955);
nor U6690 (N_6690,N_950,N_293);
xnor U6691 (N_6691,N_3223,N_321);
and U6692 (N_6692,N_2977,N_552);
nand U6693 (N_6693,N_2694,N_2416);
xor U6694 (N_6694,N_248,N_1282);
nor U6695 (N_6695,N_282,N_4370);
nand U6696 (N_6696,N_468,N_953);
nand U6697 (N_6697,N_127,N_1122);
xnor U6698 (N_6698,N_3253,N_3756);
and U6699 (N_6699,N_4139,N_2860);
or U6700 (N_6700,N_3728,N_1188);
or U6701 (N_6701,N_3501,N_3736);
nand U6702 (N_6702,N_3898,N_3960);
or U6703 (N_6703,N_4017,N_3924);
nor U6704 (N_6704,N_4447,N_3438);
xnor U6705 (N_6705,N_2353,N_2390);
nor U6706 (N_6706,N_4311,N_1852);
or U6707 (N_6707,N_2815,N_3421);
and U6708 (N_6708,N_1379,N_4045);
nand U6709 (N_6709,N_2807,N_4670);
or U6710 (N_6710,N_1705,N_3270);
nand U6711 (N_6711,N_1270,N_2205);
and U6712 (N_6712,N_1514,N_504);
or U6713 (N_6713,N_1709,N_3833);
xor U6714 (N_6714,N_4577,N_305);
nand U6715 (N_6715,N_2547,N_1614);
or U6716 (N_6716,N_983,N_3333);
nor U6717 (N_6717,N_4786,N_128);
nand U6718 (N_6718,N_1962,N_2736);
or U6719 (N_6719,N_3610,N_4912);
and U6720 (N_6720,N_3433,N_4376);
nor U6721 (N_6721,N_778,N_1336);
or U6722 (N_6722,N_2031,N_1008);
nand U6723 (N_6723,N_1805,N_419);
nand U6724 (N_6724,N_3657,N_1810);
xnor U6725 (N_6725,N_937,N_3819);
nor U6726 (N_6726,N_3412,N_4593);
xnor U6727 (N_6727,N_2579,N_1394);
nand U6728 (N_6728,N_1348,N_4242);
nand U6729 (N_6729,N_2609,N_932);
xor U6730 (N_6730,N_1666,N_2494);
xnor U6731 (N_6731,N_123,N_4550);
and U6732 (N_6732,N_3182,N_4610);
xor U6733 (N_6733,N_1064,N_4636);
nor U6734 (N_6734,N_1562,N_2019);
and U6735 (N_6735,N_3485,N_2454);
xnor U6736 (N_6736,N_1098,N_4552);
and U6737 (N_6737,N_4620,N_4351);
or U6738 (N_6738,N_4937,N_4650);
or U6739 (N_6739,N_4666,N_2213);
nor U6740 (N_6740,N_3257,N_1136);
nor U6741 (N_6741,N_482,N_3881);
xor U6742 (N_6742,N_3002,N_4164);
nor U6743 (N_6743,N_1475,N_1239);
nand U6744 (N_6744,N_2351,N_483);
nand U6745 (N_6745,N_1526,N_1707);
and U6746 (N_6746,N_2119,N_1060);
nor U6747 (N_6747,N_1989,N_4528);
and U6748 (N_6748,N_3904,N_4277);
or U6749 (N_6749,N_4965,N_4131);
nand U6750 (N_6750,N_91,N_4510);
xnor U6751 (N_6751,N_885,N_1101);
nor U6752 (N_6752,N_721,N_1217);
nor U6753 (N_6753,N_178,N_2618);
nand U6754 (N_6754,N_1863,N_2022);
xor U6755 (N_6755,N_2229,N_4547);
xnor U6756 (N_6756,N_3280,N_4064);
or U6757 (N_6757,N_1409,N_4941);
nor U6758 (N_6758,N_1350,N_2215);
and U6759 (N_6759,N_1414,N_1878);
or U6760 (N_6760,N_2612,N_1796);
or U6761 (N_6761,N_2672,N_4192);
and U6762 (N_6762,N_3117,N_2560);
nand U6763 (N_6763,N_4974,N_4122);
xor U6764 (N_6764,N_2371,N_2834);
or U6765 (N_6765,N_4762,N_3160);
nand U6766 (N_6766,N_4234,N_3769);
or U6767 (N_6767,N_737,N_301);
nand U6768 (N_6768,N_1769,N_935);
nor U6769 (N_6769,N_3624,N_966);
or U6770 (N_6770,N_3671,N_4089);
xor U6771 (N_6771,N_4721,N_2876);
nor U6772 (N_6772,N_2924,N_730);
or U6773 (N_6773,N_2484,N_3907);
nand U6774 (N_6774,N_115,N_2643);
and U6775 (N_6775,N_93,N_4208);
nand U6776 (N_6776,N_2856,N_1953);
or U6777 (N_6777,N_1057,N_3065);
nand U6778 (N_6778,N_2129,N_960);
and U6779 (N_6779,N_243,N_2223);
xnor U6780 (N_6780,N_1198,N_3990);
and U6781 (N_6781,N_3693,N_3302);
nand U6782 (N_6782,N_2432,N_1615);
nor U6783 (N_6783,N_4332,N_4203);
nor U6784 (N_6784,N_4556,N_600);
nor U6785 (N_6785,N_4872,N_1599);
xnor U6786 (N_6786,N_4456,N_1015);
xor U6787 (N_6787,N_1269,N_3951);
nand U6788 (N_6788,N_1858,N_3537);
nor U6789 (N_6789,N_4801,N_3630);
nand U6790 (N_6790,N_3644,N_4166);
or U6791 (N_6791,N_2941,N_4677);
and U6792 (N_6792,N_3584,N_4058);
nor U6793 (N_6793,N_1637,N_1894);
xnor U6794 (N_6794,N_4518,N_4453);
nand U6795 (N_6795,N_1352,N_522);
xnor U6796 (N_6796,N_3806,N_2069);
and U6797 (N_6797,N_3314,N_4703);
and U6798 (N_6798,N_139,N_4104);
nor U6799 (N_6799,N_2407,N_1911);
nor U6800 (N_6800,N_959,N_129);
or U6801 (N_6801,N_2037,N_4462);
and U6802 (N_6802,N_4701,N_604);
nor U6803 (N_6803,N_17,N_2176);
nor U6804 (N_6804,N_3090,N_2920);
nand U6805 (N_6805,N_250,N_2872);
xnor U6806 (N_6806,N_2188,N_4828);
nor U6807 (N_6807,N_1324,N_4372);
and U6808 (N_6808,N_3665,N_4022);
nor U6809 (N_6809,N_3176,N_1458);
and U6810 (N_6810,N_1680,N_4985);
or U6811 (N_6811,N_1119,N_3781);
nor U6812 (N_6812,N_3306,N_3107);
nor U6813 (N_6813,N_3075,N_1668);
xor U6814 (N_6814,N_1381,N_1047);
nand U6815 (N_6815,N_1732,N_2681);
and U6816 (N_6816,N_1721,N_4675);
nor U6817 (N_6817,N_2967,N_452);
nand U6818 (N_6818,N_4099,N_2078);
xnor U6819 (N_6819,N_1718,N_700);
xor U6820 (N_6820,N_1689,N_762);
nand U6821 (N_6821,N_2279,N_2843);
xnor U6822 (N_6822,N_2485,N_1848);
nor U6823 (N_6823,N_391,N_1626);
or U6824 (N_6824,N_3818,N_2372);
nand U6825 (N_6825,N_4814,N_847);
nand U6826 (N_6826,N_1901,N_4155);
nor U6827 (N_6827,N_327,N_1785);
nand U6828 (N_6828,N_1476,N_3895);
or U6829 (N_6829,N_2004,N_4640);
nand U6830 (N_6830,N_1250,N_1218);
or U6831 (N_6831,N_4988,N_4691);
or U6832 (N_6832,N_4130,N_676);
xnor U6833 (N_6833,N_2243,N_1182);
xnor U6834 (N_6834,N_26,N_1841);
nor U6835 (N_6835,N_4226,N_4480);
xor U6836 (N_6836,N_4506,N_4989);
and U6837 (N_6837,N_4598,N_2488);
xor U6838 (N_6838,N_4472,N_1506);
or U6839 (N_6839,N_4760,N_1909);
xor U6840 (N_6840,N_799,N_58);
and U6841 (N_6841,N_2574,N_300);
nor U6842 (N_6842,N_649,N_1531);
or U6843 (N_6843,N_116,N_1170);
or U6844 (N_6844,N_257,N_224);
or U6845 (N_6845,N_2478,N_3902);
or U6846 (N_6846,N_1364,N_872);
nor U6847 (N_6847,N_56,N_4342);
xnor U6848 (N_6848,N_4246,N_3364);
and U6849 (N_6849,N_1650,N_237);
xor U6850 (N_6850,N_3261,N_4838);
nor U6851 (N_6851,N_3039,N_3124);
and U6852 (N_6852,N_3932,N_198);
nor U6853 (N_6853,N_986,N_3936);
or U6854 (N_6854,N_4271,N_1194);
or U6855 (N_6855,N_1788,N_4336);
xor U6856 (N_6856,N_3476,N_3457);
and U6857 (N_6857,N_498,N_1791);
nor U6858 (N_6858,N_3734,N_1623);
xnor U6859 (N_6859,N_1103,N_3890);
and U6860 (N_6860,N_1150,N_428);
nand U6861 (N_6861,N_470,N_260);
nor U6862 (N_6862,N_4993,N_1519);
nor U6863 (N_6863,N_2320,N_3355);
nand U6864 (N_6864,N_171,N_1578);
nor U6865 (N_6865,N_3846,N_3521);
and U6866 (N_6866,N_3492,N_4419);
and U6867 (N_6867,N_2827,N_3957);
or U6868 (N_6868,N_1747,N_1553);
and U6869 (N_6869,N_3823,N_3024);
nor U6870 (N_6870,N_4652,N_1447);
nand U6871 (N_6871,N_2948,N_4248);
nor U6872 (N_6872,N_1225,N_4129);
or U6873 (N_6873,N_1311,N_2393);
nor U6874 (N_6874,N_3023,N_685);
nor U6875 (N_6875,N_3845,N_3877);
and U6876 (N_6876,N_4133,N_1739);
and U6877 (N_6877,N_3222,N_4071);
or U6878 (N_6878,N_4150,N_32);
or U6879 (N_6879,N_2947,N_1923);
nor U6880 (N_6880,N_3170,N_55);
or U6881 (N_6881,N_674,N_94);
nor U6882 (N_6882,N_1307,N_1100);
or U6883 (N_6883,N_4891,N_1903);
and U6884 (N_6884,N_3931,N_4642);
nor U6885 (N_6885,N_365,N_4534);
or U6886 (N_6886,N_2287,N_1974);
and U6887 (N_6887,N_4803,N_2216);
or U6888 (N_6888,N_3128,N_2891);
xnor U6889 (N_6889,N_4467,N_3749);
or U6890 (N_6890,N_415,N_891);
xnor U6891 (N_6891,N_1461,N_3334);
nand U6892 (N_6892,N_1888,N_1850);
nand U6893 (N_6893,N_1327,N_1774);
and U6894 (N_6894,N_2345,N_1949);
nand U6895 (N_6895,N_3308,N_1694);
and U6896 (N_6896,N_1607,N_253);
nor U6897 (N_6897,N_2191,N_1695);
xnor U6898 (N_6898,N_3007,N_2184);
or U6899 (N_6899,N_743,N_202);
and U6900 (N_6900,N_4243,N_1881);
and U6901 (N_6901,N_2238,N_4641);
or U6902 (N_6902,N_4492,N_879);
nand U6903 (N_6903,N_2430,N_2668);
and U6904 (N_6904,N_3782,N_4431);
nor U6905 (N_6905,N_2,N_51);
or U6906 (N_6906,N_3565,N_3700);
nand U6907 (N_6907,N_2276,N_580);
nor U6908 (N_6908,N_832,N_4811);
and U6909 (N_6909,N_3021,N_3524);
xor U6910 (N_6910,N_1315,N_3780);
xor U6911 (N_6911,N_379,N_4495);
xor U6912 (N_6912,N_1229,N_1712);
nand U6913 (N_6913,N_3108,N_2262);
or U6914 (N_6914,N_3637,N_4338);
and U6915 (N_6915,N_1706,N_431);
xnor U6916 (N_6916,N_4042,N_3567);
or U6917 (N_6917,N_2655,N_2565);
and U6918 (N_6918,N_31,N_2141);
nand U6919 (N_6919,N_2804,N_1918);
xor U6920 (N_6920,N_1163,N_4831);
nand U6921 (N_6921,N_4862,N_4816);
and U6922 (N_6922,N_2642,N_3606);
nor U6923 (N_6923,N_4536,N_3265);
nand U6924 (N_6924,N_3346,N_3268);
xnor U6925 (N_6925,N_4214,N_2142);
and U6926 (N_6926,N_3188,N_4446);
or U6927 (N_6927,N_4011,N_2868);
and U6928 (N_6928,N_4970,N_3321);
and U6929 (N_6929,N_4365,N_355);
nand U6930 (N_6930,N_3445,N_2237);
nand U6931 (N_6931,N_4861,N_1726);
or U6932 (N_6932,N_4772,N_1743);
nand U6933 (N_6933,N_1635,N_1893);
nand U6934 (N_6934,N_1685,N_2408);
or U6935 (N_6935,N_3043,N_4439);
xor U6936 (N_6936,N_4488,N_3787);
nand U6937 (N_6937,N_3649,N_4124);
or U6938 (N_6938,N_4371,N_1845);
nand U6939 (N_6939,N_3812,N_4396);
nand U6940 (N_6940,N_13,N_2640);
or U6941 (N_6941,N_4600,N_2128);
and U6942 (N_6942,N_1922,N_2789);
and U6943 (N_6943,N_4299,N_1935);
xor U6944 (N_6944,N_703,N_605);
and U6945 (N_6945,N_4606,N_895);
xnor U6946 (N_6946,N_3813,N_1092);
nor U6947 (N_6947,N_274,N_3454);
nor U6948 (N_6948,N_3995,N_2032);
nand U6949 (N_6949,N_2339,N_4050);
xor U6950 (N_6950,N_1675,N_1441);
nor U6951 (N_6951,N_2761,N_1289);
or U6952 (N_6952,N_4913,N_665);
nor U6953 (N_6953,N_609,N_3162);
nor U6954 (N_6954,N_1844,N_2660);
and U6955 (N_6955,N_4001,N_342);
xor U6956 (N_6956,N_2496,N_2464);
nand U6957 (N_6957,N_207,N_308);
or U6958 (N_6958,N_2024,N_4012);
xor U6959 (N_6959,N_1999,N_118);
nor U6960 (N_6960,N_2462,N_4986);
xor U6961 (N_6961,N_2525,N_4730);
nor U6962 (N_6962,N_2337,N_3918);
and U6963 (N_6963,N_1400,N_95);
nand U6964 (N_6964,N_232,N_2043);
or U6965 (N_6965,N_328,N_2406);
and U6966 (N_6966,N_4775,N_4247);
and U6967 (N_6967,N_1515,N_1345);
or U6968 (N_6968,N_4573,N_3081);
xor U6969 (N_6969,N_1990,N_1882);
xnor U6970 (N_6970,N_4776,N_1690);
nand U6971 (N_6971,N_4008,N_61);
and U6972 (N_6972,N_2665,N_2716);
xor U6973 (N_6973,N_2667,N_3153);
and U6974 (N_6974,N_4403,N_4887);
and U6975 (N_6975,N_4043,N_802);
xor U6976 (N_6976,N_4984,N_2677);
or U6977 (N_6977,N_134,N_2272);
and U6978 (N_6978,N_3797,N_2109);
nand U6979 (N_6979,N_4377,N_727);
nor U6980 (N_6980,N_3783,N_2593);
xor U6981 (N_6981,N_4469,N_4770);
xnor U6982 (N_6982,N_3802,N_2553);
and U6983 (N_6983,N_2318,N_2879);
nor U6984 (N_6984,N_3722,N_990);
or U6985 (N_6985,N_2703,N_3376);
or U6986 (N_6986,N_3934,N_3322);
xor U6987 (N_6987,N_2744,N_2922);
and U6988 (N_6988,N_905,N_4275);
nor U6989 (N_6989,N_2783,N_3219);
xnor U6990 (N_6990,N_3853,N_530);
or U6991 (N_6991,N_3892,N_4769);
xor U6992 (N_6992,N_4910,N_1535);
or U6993 (N_6993,N_1646,N_4268);
or U6994 (N_6994,N_2615,N_1849);
and U6995 (N_6995,N_1538,N_453);
nor U6996 (N_6996,N_4967,N_4473);
or U6997 (N_6997,N_289,N_1258);
or U6998 (N_6998,N_3304,N_1102);
nand U6999 (N_6999,N_1184,N_3751);
and U7000 (N_7000,N_414,N_3214);
or U7001 (N_7001,N_2577,N_2327);
nor U7002 (N_7002,N_1693,N_695);
and U7003 (N_7003,N_1297,N_463);
and U7004 (N_7004,N_505,N_4809);
and U7005 (N_7005,N_759,N_3576);
and U7006 (N_7006,N_4570,N_786);
nand U7007 (N_7007,N_195,N_2685);
nor U7008 (N_7008,N_131,N_4799);
xnor U7009 (N_7009,N_3045,N_2551);
and U7010 (N_7010,N_156,N_4378);
nand U7011 (N_7011,N_4884,N_270);
nor U7012 (N_7012,N_4393,N_2239);
or U7013 (N_7013,N_2580,N_2328);
nand U7014 (N_7014,N_2051,N_4795);
xor U7015 (N_7015,N_4878,N_4381);
or U7016 (N_7016,N_4037,N_367);
or U7017 (N_7017,N_899,N_3166);
nor U7018 (N_7018,N_945,N_4566);
xor U7019 (N_7019,N_2429,N_1196);
and U7020 (N_7020,N_588,N_1207);
nor U7021 (N_7021,N_3264,N_412);
nor U7022 (N_7022,N_1341,N_1775);
nor U7023 (N_7023,N_3887,N_1656);
and U7024 (N_7024,N_3575,N_3415);
xor U7025 (N_7025,N_222,N_1625);
nand U7026 (N_7026,N_4586,N_1544);
nor U7027 (N_7027,N_2231,N_3208);
xnor U7028 (N_7028,N_4333,N_1034);
nand U7029 (N_7029,N_4465,N_14);
or U7030 (N_7030,N_2571,N_3190);
xor U7031 (N_7031,N_2945,N_784);
and U7032 (N_7032,N_2235,N_1549);
or U7033 (N_7033,N_474,N_3323);
nor U7034 (N_7034,N_2110,N_1316);
xor U7035 (N_7035,N_1824,N_2001);
and U7036 (N_7036,N_512,N_3392);
or U7037 (N_7037,N_4014,N_697);
nand U7038 (N_7038,N_1242,N_108);
nor U7039 (N_7039,N_3752,N_4777);
nor U7040 (N_7040,N_3184,N_3316);
nor U7041 (N_7041,N_1720,N_2898);
and U7042 (N_7042,N_4153,N_3542);
xor U7043 (N_7043,N_234,N_4669);
xor U7044 (N_7044,N_4428,N_3089);
nand U7045 (N_7045,N_4731,N_163);
or U7046 (N_7046,N_1038,N_4157);
nand U7047 (N_7047,N_3873,N_2649);
nor U7048 (N_7048,N_3709,N_4426);
nand U7049 (N_7049,N_3112,N_2966);
and U7050 (N_7050,N_4684,N_940);
nand U7051 (N_7051,N_2770,N_4950);
and U7052 (N_7052,N_2171,N_1460);
xnor U7053 (N_7053,N_1696,N_2908);
xnor U7054 (N_7054,N_3767,N_2781);
nand U7055 (N_7055,N_1248,N_4617);
or U7056 (N_7056,N_2826,N_2926);
nand U7057 (N_7057,N_1838,N_4306);
nand U7058 (N_7058,N_574,N_760);
xnor U7059 (N_7059,N_4638,N_2491);
or U7060 (N_7060,N_726,N_3181);
or U7061 (N_7061,N_4356,N_3377);
or U7062 (N_7062,N_3360,N_4662);
xnor U7063 (N_7063,N_485,N_860);
and U7064 (N_7064,N_3594,N_2983);
nand U7065 (N_7065,N_2071,N_714);
or U7066 (N_7066,N_1319,N_3427);
and U7067 (N_7067,N_3761,N_1031);
nand U7068 (N_7068,N_3078,N_1503);
xor U7069 (N_7069,N_349,N_2907);
xnor U7070 (N_7070,N_4871,N_3721);
or U7071 (N_7071,N_3020,N_1631);
xnor U7072 (N_7072,N_4413,N_1206);
nor U7073 (N_7073,N_1386,N_1026);
nand U7074 (N_7074,N_868,N_254);
nand U7075 (N_7075,N_1641,N_460);
and U7076 (N_7076,N_1592,N_1099);
nand U7077 (N_7077,N_3478,N_1326);
nand U7078 (N_7078,N_1836,N_2343);
nor U7079 (N_7079,N_2469,N_1613);
or U7080 (N_7080,N_1831,N_1125);
nand U7081 (N_7081,N_1798,N_2558);
xnor U7082 (N_7082,N_2472,N_1620);
xor U7083 (N_7083,N_4539,N_2533);
nand U7084 (N_7084,N_800,N_2075);
xor U7085 (N_7085,N_1353,N_671);
xor U7086 (N_7086,N_1421,N_2196);
xor U7087 (N_7087,N_1335,N_4830);
xor U7088 (N_7088,N_958,N_2245);
or U7089 (N_7089,N_4886,N_3040);
nor U7090 (N_7090,N_4222,N_4138);
and U7091 (N_7091,N_646,N_764);
nor U7092 (N_7092,N_4655,N_3625);
and U7093 (N_7093,N_1895,N_1603);
and U7094 (N_7094,N_1255,N_330);
or U7095 (N_7095,N_3053,N_2775);
and U7096 (N_7096,N_1750,N_1159);
xor U7097 (N_7097,N_3060,N_3133);
or U7098 (N_7098,N_1902,N_4095);
nor U7099 (N_7099,N_2404,N_4502);
xor U7100 (N_7100,N_575,N_4184);
or U7101 (N_7101,N_2218,N_4135);
or U7102 (N_7102,N_80,N_4180);
nand U7103 (N_7103,N_1919,N_213);
nor U7104 (N_7104,N_693,N_4263);
nand U7105 (N_7105,N_1176,N_3258);
or U7106 (N_7106,N_3703,N_4565);
nor U7107 (N_7107,N_3677,N_1567);
nor U7108 (N_7108,N_2713,N_1487);
nand U7109 (N_7109,N_2597,N_4697);
nand U7110 (N_7110,N_4033,N_1547);
xor U7111 (N_7111,N_1359,N_290);
nand U7112 (N_7112,N_3417,N_2011);
and U7113 (N_7113,N_3614,N_2140);
xor U7114 (N_7114,N_507,N_1617);
or U7115 (N_7115,N_4774,N_2870);
xor U7116 (N_7116,N_3720,N_1939);
nand U7117 (N_7117,N_3929,N_2588);
xnor U7118 (N_7118,N_87,N_2265);
or U7119 (N_7119,N_2186,N_708);
and U7120 (N_7120,N_1534,N_184);
nor U7121 (N_7121,N_601,N_781);
xnor U7122 (N_7122,N_874,N_4284);
nand U7123 (N_7123,N_2939,N_1565);
xnor U7124 (N_7124,N_2823,N_1530);
and U7125 (N_7125,N_529,N_66);
nor U7126 (N_7126,N_2650,N_2960);
or U7127 (N_7127,N_3271,N_1374);
nor U7128 (N_7128,N_886,N_3431);
or U7129 (N_7129,N_880,N_3240);
xnor U7130 (N_7130,N_3979,N_2779);
and U7131 (N_7131,N_4321,N_1273);
or U7132 (N_7132,N_3691,N_862);
xor U7133 (N_7133,N_1926,N_361);
nand U7134 (N_7134,N_617,N_4698);
nand U7135 (N_7135,N_1168,N_1800);
nand U7136 (N_7136,N_4724,N_1216);
xnor U7137 (N_7137,N_2568,N_2453);
and U7138 (N_7138,N_1896,N_4079);
nor U7139 (N_7139,N_3840,N_1109);
or U7140 (N_7140,N_1702,N_3827);
or U7141 (N_7141,N_454,N_756);
xor U7142 (N_7142,N_4272,N_2849);
or U7143 (N_7143,N_1488,N_3861);
or U7144 (N_7144,N_2046,N_2314);
and U7145 (N_7145,N_4780,N_1451);
and U7146 (N_7146,N_3651,N_2033);
nand U7147 (N_7147,N_1738,N_287);
nand U7148 (N_7148,N_837,N_2601);
xor U7149 (N_7149,N_2982,N_4120);
nand U7150 (N_7150,N_3488,N_3338);
xnor U7151 (N_7151,N_2427,N_1658);
or U7152 (N_7152,N_2772,N_2969);
or U7153 (N_7153,N_294,N_2994);
nor U7154 (N_7154,N_422,N_3033);
and U7155 (N_7155,N_3950,N_3326);
or U7156 (N_7156,N_1144,N_119);
xnor U7157 (N_7157,N_4706,N_311);
nor U7158 (N_7158,N_980,N_4927);
and U7159 (N_7159,N_2370,N_4327);
nand U7160 (N_7160,N_914,N_3122);
and U7161 (N_7161,N_3374,N_1466);
or U7162 (N_7162,N_1286,N_4919);
nor U7163 (N_7163,N_1967,N_3759);
and U7164 (N_7164,N_4325,N_4387);
and U7165 (N_7165,N_1522,N_2500);
and U7166 (N_7166,N_3618,N_608);
nand U7167 (N_7167,N_3973,N_4206);
nor U7168 (N_7168,N_4864,N_740);
nor U7169 (N_7169,N_3145,N_138);
xnor U7170 (N_7170,N_2606,N_1773);
xor U7171 (N_7171,N_4717,N_2792);
nor U7172 (N_7172,N_2965,N_1752);
or U7173 (N_7173,N_2997,N_3906);
nor U7174 (N_7174,N_3545,N_1686);
or U7175 (N_7175,N_4158,N_4318);
xnor U7176 (N_7176,N_2083,N_1251);
xnor U7177 (N_7177,N_4991,N_1226);
and U7178 (N_7178,N_3424,N_4125);
nand U7179 (N_7179,N_648,N_1197);
nand U7180 (N_7180,N_3872,N_3803);
nor U7181 (N_7181,N_4779,N_326);
nor U7182 (N_7182,N_931,N_4714);
and U7183 (N_7183,N_1480,N_1426);
nor U7184 (N_7184,N_3463,N_2952);
nand U7185 (N_7185,N_2181,N_6);
and U7186 (N_7186,N_1993,N_576);
nand U7187 (N_7187,N_1183,N_1442);
and U7188 (N_7188,N_3673,N_2013);
or U7189 (N_7189,N_3646,N_1069);
and U7190 (N_7190,N_1201,N_684);
xor U7191 (N_7191,N_4601,N_3004);
xnor U7192 (N_7192,N_1317,N_3352);
xnor U7193 (N_7193,N_952,N_266);
xnor U7194 (N_7194,N_166,N_96);
nor U7195 (N_7195,N_4295,N_2166);
nand U7196 (N_7196,N_3435,N_2190);
or U7197 (N_7197,N_854,N_3127);
and U7198 (N_7198,N_4711,N_2563);
xor U7199 (N_7199,N_2385,N_2419);
and U7200 (N_7200,N_1376,N_1287);
xnor U7201 (N_7201,N_3533,N_1236);
xnor U7202 (N_7202,N_3158,N_1398);
or U7203 (N_7203,N_1095,N_3520);
and U7204 (N_7204,N_4024,N_4273);
or U7205 (N_7205,N_1016,N_987);
or U7206 (N_7206,N_4163,N_870);
nand U7207 (N_7207,N_962,N_1714);
nor U7208 (N_7208,N_3365,N_2946);
nand U7209 (N_7209,N_3577,N_495);
nand U7210 (N_7210,N_3083,N_2850);
nand U7211 (N_7211,N_3441,N_9);
xnor U7212 (N_7212,N_696,N_2503);
xnor U7213 (N_7213,N_2663,N_2060);
nor U7214 (N_7214,N_68,N_2731);
xnor U7215 (N_7215,N_3676,N_3390);
nor U7216 (N_7216,N_1267,N_3341);
and U7217 (N_7217,N_363,N_4106);
xnor U7218 (N_7218,N_2125,N_3);
or U7219 (N_7219,N_3715,N_559);
or U7220 (N_7220,N_4196,N_2111);
xor U7221 (N_7221,N_73,N_1065);
nand U7222 (N_7222,N_1262,N_1356);
nand U7223 (N_7223,N_1945,N_2750);
xnor U7224 (N_7224,N_1443,N_1854);
and U7225 (N_7225,N_2518,N_1959);
nand U7226 (N_7226,N_2414,N_2065);
nand U7227 (N_7227,N_2914,N_1279);
and U7228 (N_7228,N_2244,N_4920);
and U7229 (N_7229,N_3483,N_3512);
nand U7230 (N_7230,N_2992,N_2101);
nor U7231 (N_7231,N_4267,N_2910);
and U7232 (N_7232,N_4352,N_3534);
or U7233 (N_7233,N_968,N_2293);
nand U7234 (N_7234,N_2309,N_1558);
or U7235 (N_7235,N_2679,N_2047);
nand U7236 (N_7236,N_995,N_124);
nor U7237 (N_7237,N_132,N_3883);
nand U7238 (N_7238,N_2936,N_2436);
and U7239 (N_7239,N_3660,N_147);
or U7240 (N_7240,N_2909,N_1203);
or U7241 (N_7241,N_384,N_777);
xor U7242 (N_7242,N_653,N_3178);
and U7243 (N_7243,N_2911,N_936);
nor U7244 (N_7244,N_1698,N_2383);
nand U7245 (N_7245,N_4546,N_3113);
and U7246 (N_7246,N_4842,N_2938);
xor U7247 (N_7247,N_681,N_3123);
nand U7248 (N_7248,N_1691,N_1994);
and U7249 (N_7249,N_3510,N_1160);
or U7250 (N_7250,N_1740,N_1444);
or U7251 (N_7251,N_2968,N_4061);
nand U7252 (N_7252,N_2544,N_4584);
nor U7253 (N_7253,N_2102,N_2653);
nor U7254 (N_7254,N_925,N_2586);
and U7255 (N_7255,N_1946,N_4533);
nand U7256 (N_7256,N_1430,N_1117);
or U7257 (N_7257,N_2257,N_1884);
and U7258 (N_7258,N_1434,N_4310);
or U7259 (N_7259,N_3220,N_3815);
xor U7260 (N_7260,N_3479,N_3513);
or U7261 (N_7261,N_3150,N_4233);
nand U7262 (N_7262,N_2970,N_4914);
and U7263 (N_7263,N_2821,N_650);
xnor U7264 (N_7264,N_1899,N_4595);
and U7265 (N_7265,N_4903,N_3436);
nor U7266 (N_7266,N_4394,N_4286);
nor U7267 (N_7267,N_2934,N_1912);
or U7268 (N_7268,N_2788,N_2227);
or U7269 (N_7269,N_263,N_4088);
and U7270 (N_7270,N_2987,N_442);
nand U7271 (N_7271,N_3413,N_4418);
nor U7272 (N_7272,N_2322,N_1019);
and U7273 (N_7273,N_2254,N_33);
or U7274 (N_7274,N_4143,N_3274);
or U7275 (N_7275,N_4256,N_910);
xor U7276 (N_7276,N_3519,N_1762);
xnor U7277 (N_7277,N_763,N_1012);
nor U7278 (N_7278,N_1291,N_3037);
or U7279 (N_7279,N_2594,N_1764);
nor U7280 (N_7280,N_1070,N_4475);
nor U7281 (N_7281,N_2767,N_1220);
nor U7282 (N_7282,N_2376,N_690);
or U7283 (N_7283,N_3295,N_4517);
nor U7284 (N_7284,N_547,N_1003);
nand U7285 (N_7285,N_545,N_417);
xor U7286 (N_7286,N_4501,N_1997);
xnor U7287 (N_7287,N_1018,N_1375);
nor U7288 (N_7288,N_3744,N_1337);
and U7289 (N_7289,N_2598,N_490);
xnor U7290 (N_7290,N_4905,N_1346);
or U7291 (N_7291,N_4783,N_1214);
and U7292 (N_7292,N_815,N_3774);
and U7293 (N_7293,N_4244,N_677);
and U7294 (N_7294,N_3548,N_3518);
and U7295 (N_7295,N_2431,N_3847);
nand U7296 (N_7296,N_3912,N_806);
nand U7297 (N_7297,N_2194,N_40);
or U7298 (N_7298,N_102,N_2701);
and U7299 (N_7299,N_2089,N_3072);
or U7300 (N_7300,N_4457,N_299);
or U7301 (N_7301,N_3589,N_4115);
xnor U7302 (N_7302,N_218,N_2949);
and U7303 (N_7303,N_1632,N_4464);
nand U7304 (N_7304,N_629,N_3868);
and U7305 (N_7305,N_1013,N_3022);
xnor U7306 (N_7306,N_2248,N_302);
or U7307 (N_7307,N_4101,N_4471);
nand U7308 (N_7308,N_2633,N_3350);
and U7309 (N_7309,N_2584,N_4543);
nand U7310 (N_7310,N_1230,N_2719);
and U7311 (N_7311,N_3201,N_4347);
and U7312 (N_7312,N_2387,N_2595);
xor U7313 (N_7313,N_521,N_2146);
or U7314 (N_7314,N_3097,N_3879);
nand U7315 (N_7315,N_2136,N_1677);
and U7316 (N_7316,N_434,N_1516);
xnor U7317 (N_7317,N_1978,N_1171);
nand U7318 (N_7318,N_346,N_4624);
or U7319 (N_7319,N_1344,N_71);
xnor U7320 (N_7320,N_537,N_4078);
nor U7321 (N_7321,N_3688,N_4117);
nor U7322 (N_7322,N_317,N_2283);
or U7323 (N_7323,N_2991,N_3094);
xnor U7324 (N_7324,N_1265,N_1210);
and U7325 (N_7325,N_4645,N_742);
nand U7326 (N_7326,N_2880,N_3911);
and U7327 (N_7327,N_3294,N_276);
nand U7328 (N_7328,N_2698,N_386);
nor U7329 (N_7329,N_4825,N_3256);
xnor U7330 (N_7330,N_622,N_1438);
xor U7331 (N_7331,N_185,N_4627);
and U7332 (N_7332,N_2016,N_3497);
xnor U7333 (N_7333,N_2103,N_2310);
nand U7334 (N_7334,N_4583,N_3535);
nor U7335 (N_7335,N_3084,N_245);
nand U7336 (N_7336,N_2846,N_1509);
nor U7337 (N_7337,N_283,N_4065);
nand U7338 (N_7338,N_1729,N_2442);
nand U7339 (N_7339,N_2061,N_1851);
nor U7340 (N_7340,N_1254,N_581);
nand U7341 (N_7341,N_1853,N_556);
or U7342 (N_7342,N_1915,N_1404);
nand U7343 (N_7343,N_1002,N_2729);
nor U7344 (N_7344,N_3109,N_1672);
nand U7345 (N_7345,N_4854,N_4925);
and U7346 (N_7346,N_34,N_3903);
or U7347 (N_7347,N_4773,N_1820);
or U7348 (N_7348,N_663,N_3426);
nand U7349 (N_7349,N_4929,N_2557);
nor U7350 (N_7350,N_841,N_2979);
or U7351 (N_7351,N_3068,N_3397);
and U7352 (N_7352,N_825,N_3913);
or U7353 (N_7353,N_2317,N_3418);
or U7354 (N_7354,N_4525,N_2226);
xnor U7355 (N_7355,N_3406,N_1833);
nor U7356 (N_7356,N_3880,N_2747);
xor U7357 (N_7357,N_1169,N_4367);
and U7358 (N_7358,N_2637,N_3821);
nor U7359 (N_7359,N_1181,N_3841);
nand U7360 (N_7360,N_720,N_518);
or U7361 (N_7361,N_4353,N_188);
and U7362 (N_7362,N_4713,N_2508);
and U7363 (N_7363,N_3711,N_4962);
nor U7364 (N_7364,N_4293,N_3770);
or U7365 (N_7365,N_2082,N_1081);
xnor U7366 (N_7366,N_2212,N_789);
and U7367 (N_7367,N_555,N_4067);
nor U7368 (N_7368,N_4269,N_3151);
nor U7369 (N_7369,N_710,N_1859);
nor U7370 (N_7370,N_3394,N_3684);
xor U7371 (N_7371,N_1772,N_4128);
or U7372 (N_7372,N_4445,N_3404);
nor U7373 (N_7373,N_1700,N_292);
nand U7374 (N_7374,N_4928,N_480);
and U7375 (N_7375,N_4218,N_320);
xor U7376 (N_7376,N_4005,N_4696);
xor U7377 (N_7377,N_4694,N_3235);
nand U7378 (N_7378,N_2845,N_4963);
xor U7379 (N_7379,N_2172,N_424);
or U7380 (N_7380,N_110,N_4530);
nand U7381 (N_7381,N_1383,N_2570);
nand U7382 (N_7382,N_840,N_2304);
xnor U7383 (N_7383,N_4430,N_1135);
and U7384 (N_7384,N_2691,N_2625);
and U7385 (N_7385,N_3203,N_4759);
and U7386 (N_7386,N_2362,N_3916);
xor U7387 (N_7387,N_4245,N_1061);
nand U7388 (N_7388,N_1036,N_4185);
or U7389 (N_7389,N_1093,N_1975);
nor U7390 (N_7390,N_669,N_1653);
xnor U7391 (N_7391,N_4346,N_534);
xnor U7392 (N_7392,N_1717,N_647);
or U7393 (N_7393,N_2421,N_2009);
xnor U7394 (N_7394,N_1261,N_3592);
and U7395 (N_7395,N_4146,N_3655);
xor U7396 (N_7396,N_4545,N_1157);
nand U7397 (N_7397,N_3309,N_2875);
nor U7398 (N_7398,N_3003,N_4688);
nand U7399 (N_7399,N_374,N_167);
or U7400 (N_7400,N_180,N_1976);
nor U7401 (N_7401,N_2163,N_988);
and U7402 (N_7402,N_3648,N_3041);
xnor U7403 (N_7403,N_4228,N_2302);
nand U7404 (N_7404,N_4105,N_4579);
nor U7405 (N_7405,N_4853,N_2824);
xor U7406 (N_7406,N_3738,N_4429);
or U7407 (N_7407,N_252,N_2887);
or U7408 (N_7408,N_1147,N_4715);
or U7409 (N_7409,N_4167,N_2773);
nand U7410 (N_7410,N_3243,N_705);
or U7411 (N_7411,N_3266,N_2295);
nor U7412 (N_7412,N_12,N_3385);
and U7413 (N_7413,N_1130,N_1396);
xnor U7414 (N_7414,N_4981,N_4044);
or U7415 (N_7415,N_782,N_38);
and U7416 (N_7416,N_4613,N_946);
nand U7417 (N_7417,N_1154,N_4505);
or U7418 (N_7418,N_4943,N_3172);
and U7419 (N_7419,N_11,N_613);
nand U7420 (N_7420,N_3486,N_3210);
nor U7421 (N_7421,N_1457,N_4450);
or U7422 (N_7422,N_834,N_1305);
nand U7423 (N_7423,N_241,N_3142);
and U7424 (N_7424,N_1735,N_159);
nor U7425 (N_7425,N_2928,N_133);
and U7426 (N_7426,N_154,N_2801);
and U7427 (N_7427,N_1697,N_733);
and U7428 (N_7428,N_4787,N_517);
nand U7429 (N_7429,N_4538,N_3799);
or U7430 (N_7430,N_596,N_4186);
nor U7431 (N_7431,N_2682,N_478);
nand U7432 (N_7432,N_3048,N_3101);
xnor U7433 (N_7433,N_4763,N_4813);
nor U7434 (N_7434,N_3411,N_2308);
nor U7435 (N_7435,N_2536,N_4599);
xnor U7436 (N_7436,N_3888,N_3886);
nor U7437 (N_7437,N_3000,N_2079);
or U7438 (N_7438,N_4463,N_1313);
and U7439 (N_7439,N_2624,N_1227);
nor U7440 (N_7440,N_624,N_329);
nor U7441 (N_7441,N_3555,N_2596);
and U7442 (N_7442,N_2800,N_1802);
or U7443 (N_7443,N_4922,N_2228);
xnor U7444 (N_7444,N_401,N_1835);
nand U7445 (N_7445,N_585,N_3362);
xnor U7446 (N_7446,N_2905,N_3741);
nor U7447 (N_7447,N_3259,N_4832);
and U7448 (N_7448,N_3095,N_828);
nand U7449 (N_7449,N_1190,N_1704);
or U7450 (N_7450,N_3953,N_4478);
and U7451 (N_7451,N_4004,N_336);
xor U7452 (N_7452,N_3999,N_3977);
nand U7453 (N_7453,N_804,N_1372);
nand U7454 (N_7454,N_2112,N_747);
nand U7455 (N_7455,N_4493,N_3126);
nor U7456 (N_7456,N_3359,N_1757);
xnor U7457 (N_7457,N_2297,N_4027);
xor U7458 (N_7458,N_3617,N_1809);
nand U7459 (N_7459,N_2785,N_1778);
or U7460 (N_7460,N_4869,N_3129);
or U7461 (N_7461,N_3900,N_4366);
and U7462 (N_7462,N_4994,N_611);
nor U7463 (N_7463,N_1817,N_1235);
and U7464 (N_7464,N_4213,N_572);
and U7465 (N_7465,N_2356,N_183);
xor U7466 (N_7466,N_4754,N_2251);
or U7467 (N_7467,N_616,N_2126);
and U7468 (N_7468,N_399,N_1208);
nand U7469 (N_7469,N_1803,N_1892);
xnor U7470 (N_7470,N_1420,N_396);
nand U7471 (N_7471,N_3381,N_2177);
nand U7472 (N_7472,N_3446,N_4063);
nor U7473 (N_7473,N_754,N_4647);
nand U7474 (N_7474,N_2572,N_1483);
or U7475 (N_7475,N_3968,N_72);
and U7476 (N_7476,N_3498,N_2480);
nand U7477 (N_7477,N_3972,N_4183);
and U7478 (N_7478,N_564,N_2200);
xnor U7479 (N_7479,N_1294,N_1462);
nor U7480 (N_7480,N_930,N_1322);
and U7481 (N_7481,N_3807,N_734);
xnor U7482 (N_7482,N_455,N_3283);
and U7483 (N_7483,N_4804,N_313);
nor U7484 (N_7484,N_2183,N_3550);
and U7485 (N_7485,N_170,N_869);
or U7486 (N_7486,N_4664,N_181);
or U7487 (N_7487,N_2620,N_10);
nand U7488 (N_7488,N_713,N_459);
nor U7489 (N_7489,N_553,N_2447);
nor U7490 (N_7490,N_3564,N_392);
nor U7491 (N_7491,N_892,N_4330);
and U7492 (N_7492,N_1996,N_4252);
nand U7493 (N_7493,N_3300,N_3561);
or U7494 (N_7494,N_42,N_1621);
xnor U7495 (N_7495,N_1162,N_440);
xnor U7496 (N_7496,N_1927,N_3975);
nand U7497 (N_7497,N_4073,N_403);
nor U7498 (N_7498,N_2917,N_4235);
xnor U7499 (N_7499,N_4875,N_1727);
nand U7500 (N_7500,N_3322,N_1074);
or U7501 (N_7501,N_4169,N_4076);
nand U7502 (N_7502,N_1442,N_1399);
xor U7503 (N_7503,N_3862,N_4550);
and U7504 (N_7504,N_463,N_4794);
xnor U7505 (N_7505,N_35,N_4046);
or U7506 (N_7506,N_222,N_3624);
or U7507 (N_7507,N_2489,N_685);
xor U7508 (N_7508,N_3676,N_2898);
nor U7509 (N_7509,N_2649,N_3643);
or U7510 (N_7510,N_4242,N_2929);
xnor U7511 (N_7511,N_422,N_3938);
nand U7512 (N_7512,N_3583,N_4789);
and U7513 (N_7513,N_3654,N_389);
nand U7514 (N_7514,N_3651,N_4253);
nand U7515 (N_7515,N_565,N_3047);
xor U7516 (N_7516,N_4669,N_3982);
nand U7517 (N_7517,N_51,N_4533);
nand U7518 (N_7518,N_3317,N_4065);
nand U7519 (N_7519,N_1222,N_2935);
xnor U7520 (N_7520,N_920,N_936);
and U7521 (N_7521,N_691,N_233);
nand U7522 (N_7522,N_4518,N_4342);
xnor U7523 (N_7523,N_3222,N_4506);
xnor U7524 (N_7524,N_1063,N_599);
nand U7525 (N_7525,N_4258,N_1206);
and U7526 (N_7526,N_4707,N_1655);
nand U7527 (N_7527,N_2796,N_7);
and U7528 (N_7528,N_877,N_2507);
and U7529 (N_7529,N_3752,N_4793);
nand U7530 (N_7530,N_2735,N_838);
nor U7531 (N_7531,N_4305,N_2255);
or U7532 (N_7532,N_3851,N_2385);
xnor U7533 (N_7533,N_2880,N_2695);
or U7534 (N_7534,N_784,N_624);
or U7535 (N_7535,N_4902,N_1785);
nor U7536 (N_7536,N_812,N_1496);
xor U7537 (N_7537,N_57,N_3524);
nand U7538 (N_7538,N_357,N_490);
or U7539 (N_7539,N_2151,N_3113);
or U7540 (N_7540,N_3919,N_999);
and U7541 (N_7541,N_1160,N_2402);
nand U7542 (N_7542,N_708,N_3583);
xnor U7543 (N_7543,N_1334,N_4448);
nor U7544 (N_7544,N_1062,N_419);
nand U7545 (N_7545,N_703,N_1937);
nor U7546 (N_7546,N_2660,N_778);
xor U7547 (N_7547,N_4104,N_1343);
and U7548 (N_7548,N_4751,N_4471);
xnor U7549 (N_7549,N_549,N_4155);
nor U7550 (N_7550,N_4160,N_594);
or U7551 (N_7551,N_1668,N_673);
xor U7552 (N_7552,N_686,N_926);
nand U7553 (N_7553,N_2094,N_2650);
xor U7554 (N_7554,N_2542,N_2809);
xor U7555 (N_7555,N_1709,N_3271);
and U7556 (N_7556,N_4950,N_1201);
and U7557 (N_7557,N_1561,N_2080);
xnor U7558 (N_7558,N_3511,N_4105);
xor U7559 (N_7559,N_502,N_3965);
nand U7560 (N_7560,N_4207,N_1670);
nand U7561 (N_7561,N_954,N_3078);
nor U7562 (N_7562,N_647,N_2034);
xnor U7563 (N_7563,N_2002,N_1820);
and U7564 (N_7564,N_4682,N_730);
xnor U7565 (N_7565,N_4650,N_4851);
or U7566 (N_7566,N_764,N_3068);
or U7567 (N_7567,N_2579,N_502);
or U7568 (N_7568,N_4557,N_3787);
nor U7569 (N_7569,N_468,N_959);
nor U7570 (N_7570,N_4246,N_1034);
and U7571 (N_7571,N_739,N_2311);
nor U7572 (N_7572,N_4290,N_1657);
xnor U7573 (N_7573,N_901,N_2035);
or U7574 (N_7574,N_3053,N_3551);
nor U7575 (N_7575,N_4478,N_2404);
or U7576 (N_7576,N_2410,N_4408);
or U7577 (N_7577,N_3061,N_4123);
and U7578 (N_7578,N_1588,N_207);
and U7579 (N_7579,N_1153,N_2229);
nand U7580 (N_7580,N_1831,N_4687);
nor U7581 (N_7581,N_1751,N_1664);
or U7582 (N_7582,N_1962,N_1018);
xor U7583 (N_7583,N_3486,N_1431);
and U7584 (N_7584,N_2161,N_4912);
nor U7585 (N_7585,N_3443,N_32);
nand U7586 (N_7586,N_4989,N_1413);
nand U7587 (N_7587,N_2236,N_2853);
xor U7588 (N_7588,N_145,N_3401);
or U7589 (N_7589,N_2558,N_2070);
or U7590 (N_7590,N_3157,N_1468);
nand U7591 (N_7591,N_2884,N_4457);
and U7592 (N_7592,N_77,N_4587);
nor U7593 (N_7593,N_1100,N_1317);
or U7594 (N_7594,N_3908,N_602);
xnor U7595 (N_7595,N_2758,N_2727);
and U7596 (N_7596,N_1929,N_253);
and U7597 (N_7597,N_2837,N_3151);
and U7598 (N_7598,N_3885,N_2929);
or U7599 (N_7599,N_1017,N_1413);
nand U7600 (N_7600,N_1781,N_3695);
xnor U7601 (N_7601,N_4191,N_286);
nor U7602 (N_7602,N_2913,N_4612);
or U7603 (N_7603,N_3704,N_4877);
nand U7604 (N_7604,N_4841,N_3099);
nand U7605 (N_7605,N_2498,N_1793);
and U7606 (N_7606,N_272,N_866);
nor U7607 (N_7607,N_1323,N_1778);
nor U7608 (N_7608,N_2556,N_279);
or U7609 (N_7609,N_4531,N_4279);
or U7610 (N_7610,N_3666,N_1021);
nand U7611 (N_7611,N_376,N_4922);
xor U7612 (N_7612,N_2966,N_4430);
or U7613 (N_7613,N_4069,N_4620);
nand U7614 (N_7614,N_3820,N_3188);
or U7615 (N_7615,N_645,N_1644);
xor U7616 (N_7616,N_1370,N_2339);
or U7617 (N_7617,N_1945,N_3143);
or U7618 (N_7618,N_2643,N_3344);
nor U7619 (N_7619,N_274,N_1526);
nand U7620 (N_7620,N_2225,N_678);
nor U7621 (N_7621,N_978,N_1057);
and U7622 (N_7622,N_1146,N_4955);
nor U7623 (N_7623,N_2858,N_4914);
or U7624 (N_7624,N_1408,N_2962);
and U7625 (N_7625,N_4596,N_1192);
and U7626 (N_7626,N_4251,N_1653);
xnor U7627 (N_7627,N_1928,N_1099);
xor U7628 (N_7628,N_2876,N_1710);
and U7629 (N_7629,N_3350,N_2698);
xor U7630 (N_7630,N_3004,N_1491);
nor U7631 (N_7631,N_1107,N_2704);
and U7632 (N_7632,N_2641,N_3781);
or U7633 (N_7633,N_4085,N_2663);
nor U7634 (N_7634,N_1286,N_2197);
nand U7635 (N_7635,N_4871,N_4328);
xor U7636 (N_7636,N_2283,N_2397);
or U7637 (N_7637,N_239,N_4324);
nand U7638 (N_7638,N_3217,N_2766);
xor U7639 (N_7639,N_2710,N_2206);
xnor U7640 (N_7640,N_3304,N_3942);
and U7641 (N_7641,N_3643,N_438);
xnor U7642 (N_7642,N_4404,N_3158);
or U7643 (N_7643,N_569,N_3001);
or U7644 (N_7644,N_3513,N_1537);
nand U7645 (N_7645,N_4021,N_3417);
nor U7646 (N_7646,N_1086,N_4969);
and U7647 (N_7647,N_304,N_3344);
nor U7648 (N_7648,N_3834,N_2016);
nor U7649 (N_7649,N_2140,N_4111);
xor U7650 (N_7650,N_860,N_3146);
nor U7651 (N_7651,N_4216,N_4024);
nor U7652 (N_7652,N_2177,N_534);
nor U7653 (N_7653,N_4610,N_3093);
nand U7654 (N_7654,N_3625,N_3882);
or U7655 (N_7655,N_4890,N_4145);
xor U7656 (N_7656,N_3534,N_1058);
xor U7657 (N_7657,N_3932,N_4098);
xnor U7658 (N_7658,N_3400,N_264);
and U7659 (N_7659,N_3843,N_1623);
nor U7660 (N_7660,N_3310,N_1967);
nand U7661 (N_7661,N_4917,N_3184);
nor U7662 (N_7662,N_3122,N_223);
nor U7663 (N_7663,N_1634,N_3225);
nand U7664 (N_7664,N_605,N_2051);
or U7665 (N_7665,N_4049,N_1162);
xor U7666 (N_7666,N_1178,N_2145);
nand U7667 (N_7667,N_750,N_3346);
and U7668 (N_7668,N_3514,N_4412);
xor U7669 (N_7669,N_2841,N_4414);
xor U7670 (N_7670,N_4639,N_4470);
or U7671 (N_7671,N_4552,N_3135);
xor U7672 (N_7672,N_3041,N_4227);
xnor U7673 (N_7673,N_4613,N_3701);
and U7674 (N_7674,N_4992,N_605);
and U7675 (N_7675,N_1104,N_2708);
nand U7676 (N_7676,N_969,N_83);
and U7677 (N_7677,N_2658,N_298);
nor U7678 (N_7678,N_2566,N_3992);
nand U7679 (N_7679,N_3794,N_2219);
nor U7680 (N_7680,N_2087,N_2779);
nor U7681 (N_7681,N_309,N_4908);
nand U7682 (N_7682,N_848,N_3729);
nand U7683 (N_7683,N_4453,N_3549);
nor U7684 (N_7684,N_3182,N_1050);
nor U7685 (N_7685,N_2915,N_4002);
nor U7686 (N_7686,N_4120,N_1114);
xnor U7687 (N_7687,N_3209,N_485);
xor U7688 (N_7688,N_547,N_1805);
nand U7689 (N_7689,N_4051,N_478);
and U7690 (N_7690,N_1573,N_827);
nand U7691 (N_7691,N_3319,N_1627);
and U7692 (N_7692,N_3764,N_1002);
nor U7693 (N_7693,N_3647,N_1777);
xnor U7694 (N_7694,N_4178,N_348);
and U7695 (N_7695,N_1388,N_4682);
xor U7696 (N_7696,N_1448,N_2303);
nor U7697 (N_7697,N_4221,N_244);
nand U7698 (N_7698,N_1609,N_2875);
and U7699 (N_7699,N_1560,N_4634);
nor U7700 (N_7700,N_4183,N_1382);
or U7701 (N_7701,N_4729,N_4938);
nor U7702 (N_7702,N_2287,N_1256);
nand U7703 (N_7703,N_3957,N_4104);
and U7704 (N_7704,N_1931,N_111);
nor U7705 (N_7705,N_3989,N_3825);
xnor U7706 (N_7706,N_4985,N_4612);
nand U7707 (N_7707,N_2714,N_2138);
nor U7708 (N_7708,N_3178,N_199);
or U7709 (N_7709,N_2126,N_4103);
or U7710 (N_7710,N_3795,N_880);
nand U7711 (N_7711,N_1299,N_2258);
and U7712 (N_7712,N_908,N_1488);
and U7713 (N_7713,N_3007,N_1324);
xnor U7714 (N_7714,N_3266,N_3572);
or U7715 (N_7715,N_3614,N_4676);
xnor U7716 (N_7716,N_501,N_1210);
nand U7717 (N_7717,N_1442,N_4295);
nand U7718 (N_7718,N_1390,N_1057);
or U7719 (N_7719,N_455,N_1555);
nand U7720 (N_7720,N_2354,N_3366);
nor U7721 (N_7721,N_2605,N_4138);
or U7722 (N_7722,N_4452,N_3052);
or U7723 (N_7723,N_2271,N_2552);
xor U7724 (N_7724,N_357,N_279);
or U7725 (N_7725,N_357,N_3039);
xor U7726 (N_7726,N_2753,N_651);
nor U7727 (N_7727,N_1184,N_1859);
nand U7728 (N_7728,N_2956,N_1910);
nor U7729 (N_7729,N_453,N_4256);
or U7730 (N_7730,N_4097,N_1495);
and U7731 (N_7731,N_1944,N_1788);
or U7732 (N_7732,N_1972,N_649);
and U7733 (N_7733,N_2453,N_4654);
xor U7734 (N_7734,N_1096,N_3442);
nor U7735 (N_7735,N_3985,N_1937);
and U7736 (N_7736,N_4899,N_3794);
xnor U7737 (N_7737,N_1341,N_1843);
or U7738 (N_7738,N_1373,N_3543);
nor U7739 (N_7739,N_2419,N_2628);
nand U7740 (N_7740,N_1300,N_1716);
nor U7741 (N_7741,N_393,N_1179);
nor U7742 (N_7742,N_2404,N_2384);
or U7743 (N_7743,N_3750,N_3337);
nand U7744 (N_7744,N_4623,N_497);
nor U7745 (N_7745,N_4551,N_2698);
nand U7746 (N_7746,N_4713,N_3088);
nand U7747 (N_7747,N_3783,N_1177);
and U7748 (N_7748,N_1202,N_2456);
nor U7749 (N_7749,N_1184,N_700);
and U7750 (N_7750,N_4100,N_4568);
or U7751 (N_7751,N_511,N_2352);
nand U7752 (N_7752,N_4626,N_3328);
and U7753 (N_7753,N_1289,N_918);
nor U7754 (N_7754,N_2463,N_4892);
xnor U7755 (N_7755,N_3463,N_3684);
or U7756 (N_7756,N_4306,N_1108);
nor U7757 (N_7757,N_3778,N_1131);
nand U7758 (N_7758,N_2665,N_4208);
xnor U7759 (N_7759,N_4460,N_194);
nor U7760 (N_7760,N_685,N_4260);
and U7761 (N_7761,N_3280,N_4123);
or U7762 (N_7762,N_3971,N_902);
nand U7763 (N_7763,N_2659,N_3335);
xnor U7764 (N_7764,N_3451,N_4575);
xor U7765 (N_7765,N_1331,N_7);
xnor U7766 (N_7766,N_4973,N_2511);
or U7767 (N_7767,N_685,N_2850);
nor U7768 (N_7768,N_29,N_1778);
nor U7769 (N_7769,N_4503,N_1244);
or U7770 (N_7770,N_2752,N_3069);
xnor U7771 (N_7771,N_3389,N_1498);
and U7772 (N_7772,N_3410,N_3616);
nand U7773 (N_7773,N_3789,N_2602);
or U7774 (N_7774,N_2455,N_2008);
nand U7775 (N_7775,N_2709,N_2546);
xor U7776 (N_7776,N_4350,N_2912);
or U7777 (N_7777,N_2087,N_635);
xor U7778 (N_7778,N_4032,N_3232);
or U7779 (N_7779,N_269,N_1155);
nor U7780 (N_7780,N_3768,N_3070);
or U7781 (N_7781,N_2034,N_1622);
nor U7782 (N_7782,N_1203,N_4276);
nand U7783 (N_7783,N_3107,N_468);
xnor U7784 (N_7784,N_833,N_4362);
nor U7785 (N_7785,N_3007,N_1984);
xor U7786 (N_7786,N_2869,N_4285);
or U7787 (N_7787,N_649,N_4025);
or U7788 (N_7788,N_881,N_1268);
nand U7789 (N_7789,N_293,N_3326);
or U7790 (N_7790,N_1731,N_1311);
xor U7791 (N_7791,N_2773,N_4342);
or U7792 (N_7792,N_4094,N_1264);
xnor U7793 (N_7793,N_3615,N_4193);
or U7794 (N_7794,N_3288,N_2357);
nor U7795 (N_7795,N_2108,N_1368);
xor U7796 (N_7796,N_3536,N_309);
or U7797 (N_7797,N_92,N_1873);
nor U7798 (N_7798,N_2243,N_4437);
or U7799 (N_7799,N_2212,N_2708);
nor U7800 (N_7800,N_62,N_2226);
nor U7801 (N_7801,N_3144,N_4357);
nand U7802 (N_7802,N_1295,N_3002);
or U7803 (N_7803,N_1535,N_3539);
xor U7804 (N_7804,N_572,N_2213);
nand U7805 (N_7805,N_4213,N_2421);
xor U7806 (N_7806,N_3579,N_1951);
and U7807 (N_7807,N_3917,N_3412);
nor U7808 (N_7808,N_3697,N_4798);
xor U7809 (N_7809,N_1548,N_852);
xnor U7810 (N_7810,N_3715,N_842);
nor U7811 (N_7811,N_62,N_622);
nor U7812 (N_7812,N_2540,N_2120);
or U7813 (N_7813,N_2363,N_4865);
and U7814 (N_7814,N_4896,N_3132);
or U7815 (N_7815,N_1729,N_693);
and U7816 (N_7816,N_4075,N_3065);
nand U7817 (N_7817,N_3385,N_3410);
xnor U7818 (N_7818,N_4211,N_4056);
nand U7819 (N_7819,N_189,N_1906);
and U7820 (N_7820,N_3323,N_3725);
or U7821 (N_7821,N_925,N_3373);
nor U7822 (N_7822,N_3260,N_3233);
nor U7823 (N_7823,N_4835,N_425);
or U7824 (N_7824,N_3418,N_2906);
or U7825 (N_7825,N_3471,N_2984);
or U7826 (N_7826,N_3548,N_4674);
or U7827 (N_7827,N_4490,N_3834);
or U7828 (N_7828,N_4692,N_4509);
nor U7829 (N_7829,N_652,N_2588);
xnor U7830 (N_7830,N_1003,N_3912);
xnor U7831 (N_7831,N_3492,N_488);
nor U7832 (N_7832,N_4307,N_4596);
or U7833 (N_7833,N_389,N_1815);
xnor U7834 (N_7834,N_790,N_2023);
nor U7835 (N_7835,N_37,N_2125);
nand U7836 (N_7836,N_1319,N_1502);
or U7837 (N_7837,N_2853,N_3861);
xor U7838 (N_7838,N_221,N_3810);
or U7839 (N_7839,N_421,N_3842);
and U7840 (N_7840,N_3490,N_2138);
and U7841 (N_7841,N_2024,N_4023);
or U7842 (N_7842,N_2258,N_1761);
or U7843 (N_7843,N_1464,N_1624);
xnor U7844 (N_7844,N_515,N_1139);
xor U7845 (N_7845,N_238,N_1152);
and U7846 (N_7846,N_3696,N_1252);
or U7847 (N_7847,N_396,N_1101);
nand U7848 (N_7848,N_775,N_2887);
xnor U7849 (N_7849,N_4343,N_4700);
nor U7850 (N_7850,N_979,N_391);
nor U7851 (N_7851,N_3701,N_923);
nor U7852 (N_7852,N_4633,N_1866);
and U7853 (N_7853,N_688,N_4294);
or U7854 (N_7854,N_3775,N_1480);
xnor U7855 (N_7855,N_3775,N_1531);
nand U7856 (N_7856,N_1141,N_3079);
xor U7857 (N_7857,N_477,N_723);
nand U7858 (N_7858,N_583,N_4227);
and U7859 (N_7859,N_3866,N_4290);
nor U7860 (N_7860,N_4440,N_1204);
or U7861 (N_7861,N_4780,N_86);
nor U7862 (N_7862,N_3901,N_3694);
nor U7863 (N_7863,N_502,N_327);
xor U7864 (N_7864,N_2025,N_3695);
xor U7865 (N_7865,N_370,N_4602);
and U7866 (N_7866,N_1405,N_3695);
nor U7867 (N_7867,N_3095,N_824);
or U7868 (N_7868,N_1292,N_4849);
and U7869 (N_7869,N_1410,N_1514);
nor U7870 (N_7870,N_2459,N_569);
nand U7871 (N_7871,N_2208,N_475);
nor U7872 (N_7872,N_3965,N_3789);
nand U7873 (N_7873,N_937,N_1917);
nand U7874 (N_7874,N_1460,N_2202);
nor U7875 (N_7875,N_4198,N_3404);
xnor U7876 (N_7876,N_970,N_1007);
or U7877 (N_7877,N_91,N_876);
and U7878 (N_7878,N_2055,N_3332);
nor U7879 (N_7879,N_1577,N_4156);
or U7880 (N_7880,N_995,N_1388);
nand U7881 (N_7881,N_4948,N_854);
nor U7882 (N_7882,N_2581,N_4790);
nor U7883 (N_7883,N_138,N_1141);
xor U7884 (N_7884,N_394,N_4444);
and U7885 (N_7885,N_241,N_2983);
xor U7886 (N_7886,N_2092,N_1523);
nand U7887 (N_7887,N_3464,N_4277);
nor U7888 (N_7888,N_233,N_2337);
or U7889 (N_7889,N_1659,N_459);
and U7890 (N_7890,N_3695,N_1980);
xor U7891 (N_7891,N_4803,N_4127);
or U7892 (N_7892,N_2021,N_3960);
and U7893 (N_7893,N_4418,N_3529);
and U7894 (N_7894,N_2351,N_3063);
nor U7895 (N_7895,N_215,N_392);
or U7896 (N_7896,N_2500,N_4876);
xor U7897 (N_7897,N_3362,N_3373);
or U7898 (N_7898,N_3685,N_4326);
or U7899 (N_7899,N_1778,N_1137);
and U7900 (N_7900,N_3300,N_582);
and U7901 (N_7901,N_2473,N_1534);
xnor U7902 (N_7902,N_2193,N_2481);
nor U7903 (N_7903,N_1696,N_1509);
or U7904 (N_7904,N_1726,N_1658);
xor U7905 (N_7905,N_3228,N_948);
nand U7906 (N_7906,N_1838,N_1846);
nor U7907 (N_7907,N_2001,N_4481);
nand U7908 (N_7908,N_1747,N_2704);
nand U7909 (N_7909,N_295,N_368);
or U7910 (N_7910,N_1552,N_430);
xor U7911 (N_7911,N_3566,N_2655);
or U7912 (N_7912,N_4374,N_2768);
nand U7913 (N_7913,N_3294,N_2117);
and U7914 (N_7914,N_1425,N_4704);
nor U7915 (N_7915,N_4966,N_4778);
nor U7916 (N_7916,N_2431,N_3460);
nand U7917 (N_7917,N_4262,N_70);
xnor U7918 (N_7918,N_3965,N_2582);
nand U7919 (N_7919,N_4524,N_294);
or U7920 (N_7920,N_4746,N_1259);
nand U7921 (N_7921,N_4550,N_3664);
and U7922 (N_7922,N_1559,N_64);
nand U7923 (N_7923,N_3269,N_441);
and U7924 (N_7924,N_2059,N_2641);
and U7925 (N_7925,N_1565,N_1995);
or U7926 (N_7926,N_246,N_610);
and U7927 (N_7927,N_4020,N_4652);
and U7928 (N_7928,N_518,N_2197);
xnor U7929 (N_7929,N_641,N_2717);
xnor U7930 (N_7930,N_2604,N_2305);
nor U7931 (N_7931,N_3971,N_4241);
and U7932 (N_7932,N_4673,N_2676);
nor U7933 (N_7933,N_2987,N_812);
and U7934 (N_7934,N_4678,N_3173);
nand U7935 (N_7935,N_3743,N_970);
and U7936 (N_7936,N_4488,N_4330);
and U7937 (N_7937,N_1502,N_196);
and U7938 (N_7938,N_3391,N_4055);
xnor U7939 (N_7939,N_2238,N_2433);
or U7940 (N_7940,N_2067,N_273);
nand U7941 (N_7941,N_406,N_3821);
and U7942 (N_7942,N_1073,N_2707);
xor U7943 (N_7943,N_4648,N_4485);
nor U7944 (N_7944,N_2094,N_1521);
or U7945 (N_7945,N_4765,N_532);
or U7946 (N_7946,N_990,N_4463);
nor U7947 (N_7947,N_3656,N_2658);
and U7948 (N_7948,N_182,N_141);
nand U7949 (N_7949,N_3324,N_1454);
xor U7950 (N_7950,N_3923,N_1479);
xor U7951 (N_7951,N_308,N_72);
xor U7952 (N_7952,N_3781,N_2927);
nor U7953 (N_7953,N_162,N_2878);
and U7954 (N_7954,N_1432,N_2864);
xor U7955 (N_7955,N_4079,N_4925);
nand U7956 (N_7956,N_2070,N_2423);
or U7957 (N_7957,N_875,N_1049);
and U7958 (N_7958,N_4983,N_3649);
nor U7959 (N_7959,N_1240,N_2763);
nor U7960 (N_7960,N_142,N_3547);
xnor U7961 (N_7961,N_4705,N_40);
nand U7962 (N_7962,N_1796,N_3080);
and U7963 (N_7963,N_2571,N_621);
or U7964 (N_7964,N_3152,N_2064);
and U7965 (N_7965,N_3861,N_3067);
xnor U7966 (N_7966,N_1531,N_261);
or U7967 (N_7967,N_4688,N_4047);
nor U7968 (N_7968,N_4461,N_4987);
and U7969 (N_7969,N_190,N_1308);
nand U7970 (N_7970,N_4248,N_1874);
or U7971 (N_7971,N_2524,N_3646);
nor U7972 (N_7972,N_4897,N_2868);
or U7973 (N_7973,N_3835,N_1704);
and U7974 (N_7974,N_3403,N_3558);
and U7975 (N_7975,N_1214,N_1376);
and U7976 (N_7976,N_1208,N_3142);
nand U7977 (N_7977,N_655,N_2427);
or U7978 (N_7978,N_761,N_3770);
nand U7979 (N_7979,N_30,N_1410);
xnor U7980 (N_7980,N_380,N_4684);
or U7981 (N_7981,N_4319,N_2302);
nand U7982 (N_7982,N_2045,N_4558);
or U7983 (N_7983,N_1402,N_813);
nand U7984 (N_7984,N_4425,N_4262);
nand U7985 (N_7985,N_3393,N_2632);
xnor U7986 (N_7986,N_2927,N_3524);
nor U7987 (N_7987,N_4428,N_4325);
or U7988 (N_7988,N_936,N_2188);
nand U7989 (N_7989,N_3137,N_3721);
and U7990 (N_7990,N_291,N_2632);
or U7991 (N_7991,N_712,N_2966);
or U7992 (N_7992,N_4569,N_766);
and U7993 (N_7993,N_4012,N_4958);
nor U7994 (N_7994,N_350,N_4136);
nor U7995 (N_7995,N_4723,N_741);
nor U7996 (N_7996,N_3420,N_572);
and U7997 (N_7997,N_4073,N_93);
nor U7998 (N_7998,N_338,N_2);
nor U7999 (N_7999,N_3276,N_209);
nor U8000 (N_8000,N_2914,N_357);
xor U8001 (N_8001,N_1405,N_3416);
or U8002 (N_8002,N_2860,N_4788);
nand U8003 (N_8003,N_4607,N_3814);
and U8004 (N_8004,N_4704,N_4314);
and U8005 (N_8005,N_1917,N_1280);
and U8006 (N_8006,N_3744,N_126);
nor U8007 (N_8007,N_2929,N_2971);
xnor U8008 (N_8008,N_234,N_4763);
nor U8009 (N_8009,N_3475,N_1297);
nand U8010 (N_8010,N_62,N_397);
nand U8011 (N_8011,N_4915,N_2900);
and U8012 (N_8012,N_1209,N_4110);
xor U8013 (N_8013,N_4964,N_4406);
nor U8014 (N_8014,N_2993,N_2777);
nand U8015 (N_8015,N_2749,N_285);
nand U8016 (N_8016,N_780,N_1856);
nand U8017 (N_8017,N_2657,N_4300);
nor U8018 (N_8018,N_586,N_662);
nand U8019 (N_8019,N_537,N_1089);
or U8020 (N_8020,N_4619,N_306);
nor U8021 (N_8021,N_2681,N_2083);
or U8022 (N_8022,N_4867,N_4590);
nand U8023 (N_8023,N_2905,N_4307);
or U8024 (N_8024,N_2880,N_18);
and U8025 (N_8025,N_3273,N_4657);
and U8026 (N_8026,N_1020,N_543);
nand U8027 (N_8027,N_1048,N_1204);
and U8028 (N_8028,N_4720,N_4630);
nand U8029 (N_8029,N_2140,N_3804);
or U8030 (N_8030,N_740,N_1540);
and U8031 (N_8031,N_4123,N_1561);
nor U8032 (N_8032,N_1159,N_1173);
nand U8033 (N_8033,N_4479,N_412);
and U8034 (N_8034,N_2860,N_4369);
nor U8035 (N_8035,N_4499,N_4975);
xor U8036 (N_8036,N_852,N_1599);
nand U8037 (N_8037,N_1135,N_1400);
and U8038 (N_8038,N_2283,N_1186);
nor U8039 (N_8039,N_1751,N_3792);
nand U8040 (N_8040,N_1000,N_4691);
nand U8041 (N_8041,N_706,N_2983);
nand U8042 (N_8042,N_609,N_4841);
and U8043 (N_8043,N_3636,N_3280);
nor U8044 (N_8044,N_206,N_179);
nand U8045 (N_8045,N_1074,N_1852);
nand U8046 (N_8046,N_4622,N_219);
and U8047 (N_8047,N_2717,N_685);
and U8048 (N_8048,N_3806,N_2210);
or U8049 (N_8049,N_1870,N_2573);
nor U8050 (N_8050,N_1659,N_1290);
xor U8051 (N_8051,N_1039,N_183);
nor U8052 (N_8052,N_2306,N_2931);
xnor U8053 (N_8053,N_3199,N_2998);
and U8054 (N_8054,N_2606,N_1592);
nand U8055 (N_8055,N_3190,N_4016);
xnor U8056 (N_8056,N_3649,N_2886);
xnor U8057 (N_8057,N_4542,N_334);
or U8058 (N_8058,N_3204,N_2140);
nor U8059 (N_8059,N_3778,N_3013);
xor U8060 (N_8060,N_4223,N_307);
xnor U8061 (N_8061,N_4412,N_51);
xor U8062 (N_8062,N_877,N_1888);
xor U8063 (N_8063,N_2784,N_1117);
and U8064 (N_8064,N_2987,N_660);
nor U8065 (N_8065,N_820,N_1907);
nor U8066 (N_8066,N_1514,N_2123);
and U8067 (N_8067,N_3955,N_4156);
nor U8068 (N_8068,N_4262,N_4036);
nand U8069 (N_8069,N_1752,N_1537);
nand U8070 (N_8070,N_561,N_352);
or U8071 (N_8071,N_4109,N_1181);
nand U8072 (N_8072,N_2470,N_4179);
nand U8073 (N_8073,N_4788,N_4856);
or U8074 (N_8074,N_4924,N_2481);
nor U8075 (N_8075,N_2451,N_175);
xor U8076 (N_8076,N_2498,N_2619);
or U8077 (N_8077,N_3565,N_4157);
nand U8078 (N_8078,N_1085,N_2729);
nand U8079 (N_8079,N_3318,N_295);
nor U8080 (N_8080,N_3330,N_1070);
nor U8081 (N_8081,N_3663,N_994);
and U8082 (N_8082,N_4603,N_236);
xor U8083 (N_8083,N_164,N_2113);
or U8084 (N_8084,N_3434,N_4050);
nand U8085 (N_8085,N_2888,N_3233);
nor U8086 (N_8086,N_4186,N_1007);
and U8087 (N_8087,N_281,N_4851);
nor U8088 (N_8088,N_654,N_2935);
and U8089 (N_8089,N_1822,N_2710);
xor U8090 (N_8090,N_1803,N_3798);
or U8091 (N_8091,N_3801,N_3696);
nand U8092 (N_8092,N_1692,N_1532);
and U8093 (N_8093,N_1384,N_2124);
xor U8094 (N_8094,N_3643,N_4316);
and U8095 (N_8095,N_4203,N_1058);
nand U8096 (N_8096,N_4876,N_2795);
and U8097 (N_8097,N_477,N_1530);
and U8098 (N_8098,N_1660,N_4376);
nand U8099 (N_8099,N_4724,N_1035);
nor U8100 (N_8100,N_3535,N_2392);
xor U8101 (N_8101,N_1240,N_392);
or U8102 (N_8102,N_3970,N_3363);
or U8103 (N_8103,N_1580,N_1538);
xor U8104 (N_8104,N_504,N_1654);
or U8105 (N_8105,N_3261,N_75);
xnor U8106 (N_8106,N_1112,N_3737);
xor U8107 (N_8107,N_1390,N_1134);
nand U8108 (N_8108,N_950,N_692);
xor U8109 (N_8109,N_1693,N_3030);
and U8110 (N_8110,N_268,N_2770);
and U8111 (N_8111,N_2167,N_872);
nor U8112 (N_8112,N_3521,N_38);
and U8113 (N_8113,N_2725,N_426);
and U8114 (N_8114,N_4752,N_4702);
xor U8115 (N_8115,N_1529,N_4836);
or U8116 (N_8116,N_4331,N_1794);
xor U8117 (N_8117,N_4787,N_3208);
nor U8118 (N_8118,N_2525,N_2251);
nor U8119 (N_8119,N_2876,N_3383);
nor U8120 (N_8120,N_44,N_741);
nand U8121 (N_8121,N_1341,N_2572);
or U8122 (N_8122,N_2312,N_3649);
and U8123 (N_8123,N_644,N_1889);
xnor U8124 (N_8124,N_406,N_1373);
or U8125 (N_8125,N_3956,N_1757);
and U8126 (N_8126,N_3770,N_1848);
nor U8127 (N_8127,N_855,N_3222);
xnor U8128 (N_8128,N_3455,N_4312);
xor U8129 (N_8129,N_3337,N_2145);
nand U8130 (N_8130,N_4444,N_4405);
xor U8131 (N_8131,N_3416,N_4790);
nand U8132 (N_8132,N_1280,N_3397);
nor U8133 (N_8133,N_654,N_2460);
nor U8134 (N_8134,N_3469,N_3694);
xor U8135 (N_8135,N_953,N_4577);
and U8136 (N_8136,N_58,N_1859);
and U8137 (N_8137,N_4863,N_388);
or U8138 (N_8138,N_540,N_4631);
or U8139 (N_8139,N_4242,N_3253);
and U8140 (N_8140,N_2150,N_4353);
or U8141 (N_8141,N_2317,N_1282);
nor U8142 (N_8142,N_2859,N_1785);
nand U8143 (N_8143,N_2268,N_1550);
or U8144 (N_8144,N_4995,N_4786);
and U8145 (N_8145,N_4320,N_1731);
nand U8146 (N_8146,N_1551,N_1920);
nor U8147 (N_8147,N_3833,N_3311);
nor U8148 (N_8148,N_2302,N_579);
xnor U8149 (N_8149,N_57,N_4680);
nand U8150 (N_8150,N_769,N_2483);
and U8151 (N_8151,N_4407,N_1013);
nor U8152 (N_8152,N_4958,N_3242);
and U8153 (N_8153,N_414,N_3873);
and U8154 (N_8154,N_2071,N_1677);
nand U8155 (N_8155,N_4457,N_1621);
xnor U8156 (N_8156,N_2628,N_1193);
and U8157 (N_8157,N_1457,N_3438);
nor U8158 (N_8158,N_4625,N_4292);
nand U8159 (N_8159,N_3345,N_3567);
nand U8160 (N_8160,N_385,N_2962);
nand U8161 (N_8161,N_770,N_3741);
nand U8162 (N_8162,N_106,N_1375);
nor U8163 (N_8163,N_2963,N_1522);
nand U8164 (N_8164,N_3335,N_4246);
xor U8165 (N_8165,N_4743,N_1545);
or U8166 (N_8166,N_1025,N_2574);
nand U8167 (N_8167,N_2337,N_3244);
and U8168 (N_8168,N_2620,N_42);
and U8169 (N_8169,N_4347,N_3971);
and U8170 (N_8170,N_3041,N_1482);
or U8171 (N_8171,N_110,N_3921);
nor U8172 (N_8172,N_1825,N_4385);
or U8173 (N_8173,N_3585,N_4968);
nand U8174 (N_8174,N_3017,N_3246);
nand U8175 (N_8175,N_2505,N_2329);
nand U8176 (N_8176,N_4590,N_3078);
or U8177 (N_8177,N_1583,N_4765);
nor U8178 (N_8178,N_780,N_2181);
and U8179 (N_8179,N_3260,N_1759);
or U8180 (N_8180,N_264,N_545);
nand U8181 (N_8181,N_3010,N_4545);
nor U8182 (N_8182,N_571,N_2808);
and U8183 (N_8183,N_1327,N_4252);
and U8184 (N_8184,N_4803,N_1364);
nand U8185 (N_8185,N_613,N_2834);
nand U8186 (N_8186,N_1205,N_2730);
xor U8187 (N_8187,N_3135,N_3385);
and U8188 (N_8188,N_4400,N_2643);
and U8189 (N_8189,N_3270,N_1256);
nand U8190 (N_8190,N_3376,N_4758);
nand U8191 (N_8191,N_1692,N_2257);
nor U8192 (N_8192,N_3354,N_589);
or U8193 (N_8193,N_3281,N_706);
or U8194 (N_8194,N_262,N_4398);
nand U8195 (N_8195,N_1013,N_843);
nand U8196 (N_8196,N_3855,N_3768);
xnor U8197 (N_8197,N_352,N_4270);
nor U8198 (N_8198,N_2202,N_2126);
xnor U8199 (N_8199,N_4145,N_4860);
or U8200 (N_8200,N_1030,N_1538);
and U8201 (N_8201,N_110,N_2007);
nand U8202 (N_8202,N_4840,N_1070);
or U8203 (N_8203,N_2229,N_4600);
nor U8204 (N_8204,N_2262,N_257);
nand U8205 (N_8205,N_2719,N_2067);
nand U8206 (N_8206,N_1074,N_2828);
nor U8207 (N_8207,N_1771,N_1308);
and U8208 (N_8208,N_1754,N_3743);
nand U8209 (N_8209,N_2512,N_4609);
and U8210 (N_8210,N_3351,N_4465);
or U8211 (N_8211,N_4267,N_2200);
or U8212 (N_8212,N_372,N_338);
nand U8213 (N_8213,N_2326,N_111);
nand U8214 (N_8214,N_2163,N_4063);
nand U8215 (N_8215,N_2943,N_1190);
and U8216 (N_8216,N_3894,N_569);
or U8217 (N_8217,N_3444,N_649);
nand U8218 (N_8218,N_3034,N_3617);
nand U8219 (N_8219,N_4416,N_2596);
nor U8220 (N_8220,N_516,N_905);
or U8221 (N_8221,N_2120,N_1776);
or U8222 (N_8222,N_855,N_4195);
xor U8223 (N_8223,N_3675,N_3246);
or U8224 (N_8224,N_1991,N_4130);
nor U8225 (N_8225,N_1215,N_1162);
or U8226 (N_8226,N_3472,N_3278);
xor U8227 (N_8227,N_1903,N_3900);
xor U8228 (N_8228,N_4148,N_4496);
nand U8229 (N_8229,N_1384,N_3996);
nor U8230 (N_8230,N_4101,N_2907);
and U8231 (N_8231,N_2548,N_1483);
nand U8232 (N_8232,N_1580,N_3783);
nor U8233 (N_8233,N_3715,N_3827);
or U8234 (N_8234,N_3052,N_1209);
or U8235 (N_8235,N_165,N_4658);
nor U8236 (N_8236,N_2573,N_906);
nor U8237 (N_8237,N_4641,N_2351);
nand U8238 (N_8238,N_971,N_872);
or U8239 (N_8239,N_1565,N_939);
or U8240 (N_8240,N_2096,N_2330);
xnor U8241 (N_8241,N_564,N_1652);
nand U8242 (N_8242,N_2926,N_2359);
nor U8243 (N_8243,N_4454,N_3523);
and U8244 (N_8244,N_3069,N_725);
nand U8245 (N_8245,N_3822,N_2588);
nand U8246 (N_8246,N_4080,N_4643);
xnor U8247 (N_8247,N_1134,N_823);
or U8248 (N_8248,N_1081,N_2254);
or U8249 (N_8249,N_1108,N_552);
and U8250 (N_8250,N_1141,N_3670);
and U8251 (N_8251,N_3358,N_1001);
or U8252 (N_8252,N_4865,N_3192);
nor U8253 (N_8253,N_2227,N_3497);
xor U8254 (N_8254,N_4723,N_3270);
nand U8255 (N_8255,N_1255,N_2553);
or U8256 (N_8256,N_989,N_1130);
or U8257 (N_8257,N_3635,N_2380);
or U8258 (N_8258,N_4945,N_582);
nand U8259 (N_8259,N_3391,N_4370);
and U8260 (N_8260,N_3717,N_1486);
xnor U8261 (N_8261,N_1969,N_142);
nor U8262 (N_8262,N_677,N_1101);
xnor U8263 (N_8263,N_603,N_1205);
and U8264 (N_8264,N_825,N_178);
nor U8265 (N_8265,N_4391,N_756);
xor U8266 (N_8266,N_446,N_2232);
nor U8267 (N_8267,N_3033,N_4000);
nand U8268 (N_8268,N_4354,N_1607);
and U8269 (N_8269,N_495,N_2914);
nor U8270 (N_8270,N_3153,N_2332);
and U8271 (N_8271,N_4341,N_1627);
or U8272 (N_8272,N_4122,N_1853);
xnor U8273 (N_8273,N_2029,N_3237);
or U8274 (N_8274,N_2058,N_4953);
and U8275 (N_8275,N_268,N_3334);
or U8276 (N_8276,N_2222,N_910);
or U8277 (N_8277,N_1238,N_4633);
or U8278 (N_8278,N_1227,N_758);
xnor U8279 (N_8279,N_3318,N_2233);
and U8280 (N_8280,N_494,N_1708);
xnor U8281 (N_8281,N_628,N_4458);
or U8282 (N_8282,N_2983,N_2854);
nand U8283 (N_8283,N_3317,N_4974);
nand U8284 (N_8284,N_683,N_1724);
xor U8285 (N_8285,N_3,N_3345);
nor U8286 (N_8286,N_1841,N_2461);
xnor U8287 (N_8287,N_1540,N_1755);
or U8288 (N_8288,N_1093,N_2785);
xnor U8289 (N_8289,N_1927,N_535);
or U8290 (N_8290,N_2378,N_2223);
nor U8291 (N_8291,N_1793,N_4872);
and U8292 (N_8292,N_3121,N_2322);
and U8293 (N_8293,N_4107,N_3426);
and U8294 (N_8294,N_3933,N_1284);
and U8295 (N_8295,N_4717,N_921);
or U8296 (N_8296,N_1680,N_3870);
nand U8297 (N_8297,N_3310,N_3422);
xnor U8298 (N_8298,N_4002,N_311);
xnor U8299 (N_8299,N_3219,N_4884);
and U8300 (N_8300,N_377,N_4226);
nor U8301 (N_8301,N_3149,N_1229);
and U8302 (N_8302,N_3017,N_3037);
nor U8303 (N_8303,N_3333,N_3852);
and U8304 (N_8304,N_3898,N_1539);
or U8305 (N_8305,N_2044,N_4283);
or U8306 (N_8306,N_437,N_363);
nor U8307 (N_8307,N_2505,N_2653);
nand U8308 (N_8308,N_2776,N_1170);
xnor U8309 (N_8309,N_1382,N_104);
nand U8310 (N_8310,N_2803,N_1831);
nand U8311 (N_8311,N_2191,N_1961);
nor U8312 (N_8312,N_4084,N_2703);
nor U8313 (N_8313,N_3950,N_2941);
or U8314 (N_8314,N_81,N_1475);
nor U8315 (N_8315,N_2782,N_1311);
nor U8316 (N_8316,N_2563,N_2614);
or U8317 (N_8317,N_3448,N_2752);
and U8318 (N_8318,N_4458,N_4306);
and U8319 (N_8319,N_2791,N_4336);
nand U8320 (N_8320,N_2298,N_1498);
nand U8321 (N_8321,N_2579,N_4432);
xnor U8322 (N_8322,N_1997,N_3249);
and U8323 (N_8323,N_838,N_1879);
and U8324 (N_8324,N_4416,N_753);
nand U8325 (N_8325,N_1023,N_1777);
nand U8326 (N_8326,N_3146,N_3268);
and U8327 (N_8327,N_1645,N_1610);
nand U8328 (N_8328,N_812,N_4978);
and U8329 (N_8329,N_2112,N_788);
xor U8330 (N_8330,N_1437,N_581);
and U8331 (N_8331,N_4875,N_4640);
xor U8332 (N_8332,N_2129,N_2514);
or U8333 (N_8333,N_108,N_794);
or U8334 (N_8334,N_2073,N_3685);
xnor U8335 (N_8335,N_3925,N_4320);
or U8336 (N_8336,N_1110,N_1748);
nand U8337 (N_8337,N_2390,N_3210);
nand U8338 (N_8338,N_3421,N_4882);
and U8339 (N_8339,N_0,N_1569);
xor U8340 (N_8340,N_1340,N_1188);
nor U8341 (N_8341,N_3275,N_1687);
nand U8342 (N_8342,N_460,N_3481);
or U8343 (N_8343,N_1939,N_4936);
or U8344 (N_8344,N_2971,N_618);
and U8345 (N_8345,N_1096,N_985);
nand U8346 (N_8346,N_2746,N_4531);
xnor U8347 (N_8347,N_2111,N_4269);
and U8348 (N_8348,N_93,N_4213);
nand U8349 (N_8349,N_591,N_4699);
nand U8350 (N_8350,N_2662,N_4052);
xor U8351 (N_8351,N_1922,N_1059);
and U8352 (N_8352,N_2934,N_1597);
or U8353 (N_8353,N_887,N_2594);
nor U8354 (N_8354,N_4781,N_830);
and U8355 (N_8355,N_2917,N_957);
nand U8356 (N_8356,N_1635,N_3577);
nor U8357 (N_8357,N_3100,N_618);
or U8358 (N_8358,N_3519,N_2313);
and U8359 (N_8359,N_218,N_967);
nand U8360 (N_8360,N_3319,N_3380);
nand U8361 (N_8361,N_801,N_2982);
nand U8362 (N_8362,N_2551,N_3365);
nor U8363 (N_8363,N_3374,N_2407);
or U8364 (N_8364,N_2444,N_3945);
nand U8365 (N_8365,N_689,N_4785);
or U8366 (N_8366,N_3682,N_1563);
nand U8367 (N_8367,N_2300,N_3865);
xor U8368 (N_8368,N_1952,N_4861);
nand U8369 (N_8369,N_4407,N_1501);
xnor U8370 (N_8370,N_4963,N_4138);
xor U8371 (N_8371,N_3542,N_1734);
nand U8372 (N_8372,N_547,N_3841);
xor U8373 (N_8373,N_2729,N_4746);
xnor U8374 (N_8374,N_4361,N_4);
nand U8375 (N_8375,N_51,N_2214);
xor U8376 (N_8376,N_3633,N_2666);
or U8377 (N_8377,N_4626,N_3539);
xnor U8378 (N_8378,N_2704,N_159);
nand U8379 (N_8379,N_847,N_2023);
xor U8380 (N_8380,N_105,N_3303);
xnor U8381 (N_8381,N_3472,N_1684);
and U8382 (N_8382,N_862,N_1828);
nor U8383 (N_8383,N_3829,N_3130);
nor U8384 (N_8384,N_3270,N_1675);
xnor U8385 (N_8385,N_4736,N_1232);
nor U8386 (N_8386,N_4616,N_1469);
or U8387 (N_8387,N_4950,N_1824);
and U8388 (N_8388,N_4020,N_1118);
or U8389 (N_8389,N_3090,N_3997);
or U8390 (N_8390,N_323,N_3853);
xor U8391 (N_8391,N_1883,N_3931);
xor U8392 (N_8392,N_2385,N_868);
xnor U8393 (N_8393,N_789,N_1931);
xnor U8394 (N_8394,N_1747,N_2072);
nor U8395 (N_8395,N_3634,N_2012);
xnor U8396 (N_8396,N_367,N_705);
nand U8397 (N_8397,N_3703,N_2920);
xnor U8398 (N_8398,N_3402,N_2317);
or U8399 (N_8399,N_1573,N_2933);
nor U8400 (N_8400,N_3704,N_1970);
and U8401 (N_8401,N_4657,N_2674);
xnor U8402 (N_8402,N_4744,N_4233);
nand U8403 (N_8403,N_3606,N_495);
nor U8404 (N_8404,N_4596,N_1169);
xor U8405 (N_8405,N_4792,N_3957);
and U8406 (N_8406,N_3077,N_4202);
nand U8407 (N_8407,N_572,N_21);
nor U8408 (N_8408,N_4975,N_2487);
xor U8409 (N_8409,N_1649,N_3311);
xor U8410 (N_8410,N_1672,N_2853);
nor U8411 (N_8411,N_2330,N_4143);
nor U8412 (N_8412,N_3431,N_4740);
or U8413 (N_8413,N_2640,N_4788);
nand U8414 (N_8414,N_690,N_2217);
nand U8415 (N_8415,N_1015,N_3941);
xnor U8416 (N_8416,N_2109,N_95);
or U8417 (N_8417,N_3726,N_2665);
nand U8418 (N_8418,N_1136,N_1288);
xnor U8419 (N_8419,N_1341,N_4551);
and U8420 (N_8420,N_2974,N_4972);
nand U8421 (N_8421,N_1465,N_4401);
or U8422 (N_8422,N_1900,N_3392);
and U8423 (N_8423,N_270,N_3513);
and U8424 (N_8424,N_2220,N_3197);
nand U8425 (N_8425,N_1883,N_68);
and U8426 (N_8426,N_1122,N_1860);
or U8427 (N_8427,N_452,N_3337);
or U8428 (N_8428,N_2360,N_2607);
nor U8429 (N_8429,N_3743,N_3716);
nand U8430 (N_8430,N_280,N_1434);
and U8431 (N_8431,N_3804,N_4509);
xnor U8432 (N_8432,N_2986,N_2579);
nor U8433 (N_8433,N_4888,N_565);
xnor U8434 (N_8434,N_646,N_3908);
or U8435 (N_8435,N_2702,N_3366);
or U8436 (N_8436,N_1605,N_1445);
nor U8437 (N_8437,N_2516,N_2210);
nand U8438 (N_8438,N_1126,N_749);
nand U8439 (N_8439,N_4392,N_1849);
and U8440 (N_8440,N_4152,N_1179);
and U8441 (N_8441,N_4291,N_4125);
xor U8442 (N_8442,N_4250,N_3002);
or U8443 (N_8443,N_406,N_172);
xnor U8444 (N_8444,N_3641,N_984);
and U8445 (N_8445,N_3263,N_233);
nor U8446 (N_8446,N_2028,N_2819);
nor U8447 (N_8447,N_1987,N_4799);
and U8448 (N_8448,N_4549,N_1484);
and U8449 (N_8449,N_4785,N_712);
xor U8450 (N_8450,N_4087,N_4071);
or U8451 (N_8451,N_2951,N_579);
and U8452 (N_8452,N_1603,N_3226);
nand U8453 (N_8453,N_273,N_3702);
and U8454 (N_8454,N_4519,N_3325);
xnor U8455 (N_8455,N_2062,N_3589);
nor U8456 (N_8456,N_2401,N_2456);
or U8457 (N_8457,N_2684,N_1236);
nand U8458 (N_8458,N_959,N_1549);
or U8459 (N_8459,N_1333,N_4312);
xor U8460 (N_8460,N_4124,N_3232);
or U8461 (N_8461,N_1836,N_2754);
and U8462 (N_8462,N_4859,N_3482);
xor U8463 (N_8463,N_3745,N_4007);
nor U8464 (N_8464,N_1497,N_4146);
nand U8465 (N_8465,N_2318,N_1036);
xor U8466 (N_8466,N_1488,N_1228);
and U8467 (N_8467,N_3793,N_1737);
and U8468 (N_8468,N_4855,N_4338);
nand U8469 (N_8469,N_2818,N_546);
xor U8470 (N_8470,N_3670,N_3888);
xor U8471 (N_8471,N_3332,N_4531);
xor U8472 (N_8472,N_4066,N_4859);
and U8473 (N_8473,N_1199,N_4929);
or U8474 (N_8474,N_3252,N_3384);
and U8475 (N_8475,N_812,N_3691);
and U8476 (N_8476,N_788,N_359);
and U8477 (N_8477,N_2001,N_4138);
nand U8478 (N_8478,N_681,N_3022);
nand U8479 (N_8479,N_2080,N_2060);
and U8480 (N_8480,N_4630,N_243);
xor U8481 (N_8481,N_4318,N_3256);
and U8482 (N_8482,N_4794,N_3434);
nand U8483 (N_8483,N_2472,N_1598);
nand U8484 (N_8484,N_2828,N_1660);
nand U8485 (N_8485,N_4781,N_4326);
xnor U8486 (N_8486,N_3907,N_4187);
or U8487 (N_8487,N_2373,N_4143);
nor U8488 (N_8488,N_1943,N_773);
or U8489 (N_8489,N_3593,N_1190);
nand U8490 (N_8490,N_1699,N_2903);
and U8491 (N_8491,N_1509,N_4805);
nand U8492 (N_8492,N_1981,N_3874);
xnor U8493 (N_8493,N_251,N_1439);
nand U8494 (N_8494,N_2712,N_2246);
and U8495 (N_8495,N_3556,N_3269);
nor U8496 (N_8496,N_1506,N_4787);
nand U8497 (N_8497,N_4845,N_4330);
and U8498 (N_8498,N_4972,N_3200);
xor U8499 (N_8499,N_3864,N_388);
nand U8500 (N_8500,N_3416,N_1135);
and U8501 (N_8501,N_2875,N_4941);
nor U8502 (N_8502,N_846,N_1606);
nor U8503 (N_8503,N_322,N_1948);
or U8504 (N_8504,N_1490,N_1166);
xnor U8505 (N_8505,N_2603,N_1018);
or U8506 (N_8506,N_4813,N_3518);
xnor U8507 (N_8507,N_1464,N_3824);
and U8508 (N_8508,N_4086,N_4310);
nor U8509 (N_8509,N_1480,N_1946);
and U8510 (N_8510,N_2366,N_2170);
and U8511 (N_8511,N_913,N_308);
nor U8512 (N_8512,N_4416,N_2853);
xnor U8513 (N_8513,N_877,N_3602);
and U8514 (N_8514,N_617,N_1836);
nor U8515 (N_8515,N_1130,N_3850);
or U8516 (N_8516,N_601,N_4255);
nor U8517 (N_8517,N_3858,N_4605);
nor U8518 (N_8518,N_2720,N_785);
xor U8519 (N_8519,N_263,N_1218);
nand U8520 (N_8520,N_3952,N_556);
nor U8521 (N_8521,N_1050,N_3559);
nand U8522 (N_8522,N_4440,N_3194);
and U8523 (N_8523,N_98,N_1915);
nor U8524 (N_8524,N_3431,N_3528);
nor U8525 (N_8525,N_4571,N_1169);
nand U8526 (N_8526,N_2107,N_4360);
nand U8527 (N_8527,N_556,N_2348);
or U8528 (N_8528,N_1018,N_1550);
or U8529 (N_8529,N_2392,N_67);
nand U8530 (N_8530,N_4809,N_4449);
nor U8531 (N_8531,N_4330,N_1125);
xor U8532 (N_8532,N_3477,N_2164);
and U8533 (N_8533,N_2827,N_3171);
nand U8534 (N_8534,N_2460,N_2905);
nand U8535 (N_8535,N_204,N_1413);
xnor U8536 (N_8536,N_3074,N_2528);
and U8537 (N_8537,N_4517,N_650);
or U8538 (N_8538,N_3976,N_2013);
and U8539 (N_8539,N_2418,N_2304);
nor U8540 (N_8540,N_1125,N_206);
and U8541 (N_8541,N_3884,N_2798);
or U8542 (N_8542,N_3281,N_4917);
xor U8543 (N_8543,N_1098,N_4545);
or U8544 (N_8544,N_2706,N_58);
and U8545 (N_8545,N_3995,N_295);
nor U8546 (N_8546,N_3612,N_213);
xnor U8547 (N_8547,N_743,N_51);
or U8548 (N_8548,N_2353,N_564);
and U8549 (N_8549,N_2729,N_2561);
nand U8550 (N_8550,N_4247,N_4370);
or U8551 (N_8551,N_1347,N_191);
or U8552 (N_8552,N_2930,N_1430);
or U8553 (N_8553,N_4254,N_158);
xor U8554 (N_8554,N_1721,N_4602);
or U8555 (N_8555,N_4545,N_2734);
xor U8556 (N_8556,N_1391,N_3556);
xor U8557 (N_8557,N_120,N_1234);
nor U8558 (N_8558,N_4554,N_54);
xor U8559 (N_8559,N_366,N_966);
nand U8560 (N_8560,N_22,N_1169);
xnor U8561 (N_8561,N_3914,N_4253);
or U8562 (N_8562,N_2721,N_3921);
nor U8563 (N_8563,N_2202,N_2879);
or U8564 (N_8564,N_955,N_1358);
and U8565 (N_8565,N_3685,N_4533);
and U8566 (N_8566,N_2029,N_3873);
and U8567 (N_8567,N_4508,N_3024);
xnor U8568 (N_8568,N_3694,N_1758);
or U8569 (N_8569,N_3876,N_839);
nand U8570 (N_8570,N_3664,N_2032);
or U8571 (N_8571,N_3487,N_2873);
nor U8572 (N_8572,N_3767,N_3921);
nor U8573 (N_8573,N_1988,N_1091);
and U8574 (N_8574,N_1010,N_1383);
and U8575 (N_8575,N_2828,N_4981);
xor U8576 (N_8576,N_3553,N_592);
or U8577 (N_8577,N_3948,N_1339);
and U8578 (N_8578,N_3723,N_106);
and U8579 (N_8579,N_2605,N_4684);
xnor U8580 (N_8580,N_4198,N_438);
and U8581 (N_8581,N_3964,N_4619);
nand U8582 (N_8582,N_4414,N_4379);
nor U8583 (N_8583,N_4325,N_3164);
and U8584 (N_8584,N_1300,N_3188);
nand U8585 (N_8585,N_2573,N_4645);
xor U8586 (N_8586,N_781,N_136);
and U8587 (N_8587,N_3084,N_4376);
or U8588 (N_8588,N_4967,N_4624);
or U8589 (N_8589,N_2932,N_3685);
nand U8590 (N_8590,N_2114,N_3331);
and U8591 (N_8591,N_1350,N_3331);
xor U8592 (N_8592,N_1051,N_4901);
nor U8593 (N_8593,N_2799,N_173);
nand U8594 (N_8594,N_4601,N_2004);
nand U8595 (N_8595,N_378,N_120);
and U8596 (N_8596,N_69,N_1926);
nor U8597 (N_8597,N_2381,N_4979);
and U8598 (N_8598,N_3328,N_190);
nand U8599 (N_8599,N_60,N_2347);
nor U8600 (N_8600,N_3899,N_2779);
nor U8601 (N_8601,N_3663,N_897);
xor U8602 (N_8602,N_1372,N_3040);
and U8603 (N_8603,N_3648,N_3150);
nor U8604 (N_8604,N_1305,N_3913);
nor U8605 (N_8605,N_4851,N_4224);
xor U8606 (N_8606,N_2669,N_857);
or U8607 (N_8607,N_3931,N_278);
and U8608 (N_8608,N_4250,N_1325);
nand U8609 (N_8609,N_574,N_791);
nor U8610 (N_8610,N_4692,N_983);
nand U8611 (N_8611,N_4844,N_2236);
or U8612 (N_8612,N_2682,N_3986);
xnor U8613 (N_8613,N_3642,N_2203);
nor U8614 (N_8614,N_2930,N_4264);
or U8615 (N_8615,N_1969,N_1105);
and U8616 (N_8616,N_2263,N_2255);
nor U8617 (N_8617,N_518,N_1817);
xor U8618 (N_8618,N_1414,N_4649);
nand U8619 (N_8619,N_3300,N_2454);
nor U8620 (N_8620,N_2463,N_3245);
and U8621 (N_8621,N_4500,N_2829);
and U8622 (N_8622,N_1079,N_3522);
xnor U8623 (N_8623,N_1734,N_1221);
xor U8624 (N_8624,N_161,N_3325);
xor U8625 (N_8625,N_1181,N_307);
xor U8626 (N_8626,N_4811,N_1236);
or U8627 (N_8627,N_4493,N_307);
xnor U8628 (N_8628,N_2867,N_2053);
and U8629 (N_8629,N_885,N_2503);
or U8630 (N_8630,N_336,N_4155);
nand U8631 (N_8631,N_874,N_543);
nand U8632 (N_8632,N_2014,N_3344);
xor U8633 (N_8633,N_1902,N_1665);
nand U8634 (N_8634,N_3420,N_2976);
xnor U8635 (N_8635,N_4892,N_517);
or U8636 (N_8636,N_2766,N_1537);
nor U8637 (N_8637,N_4828,N_4047);
xor U8638 (N_8638,N_1352,N_1134);
or U8639 (N_8639,N_3011,N_1620);
nand U8640 (N_8640,N_1395,N_1437);
and U8641 (N_8641,N_4341,N_3209);
and U8642 (N_8642,N_1622,N_4136);
xnor U8643 (N_8643,N_2059,N_3567);
or U8644 (N_8644,N_4341,N_1642);
nor U8645 (N_8645,N_1880,N_958);
and U8646 (N_8646,N_2549,N_3037);
xnor U8647 (N_8647,N_4084,N_3345);
nor U8648 (N_8648,N_3435,N_335);
xor U8649 (N_8649,N_4630,N_2569);
or U8650 (N_8650,N_2787,N_3235);
or U8651 (N_8651,N_4069,N_3750);
and U8652 (N_8652,N_2859,N_1119);
nand U8653 (N_8653,N_4167,N_4443);
or U8654 (N_8654,N_3731,N_4236);
nor U8655 (N_8655,N_1699,N_2792);
xnor U8656 (N_8656,N_1829,N_853);
nor U8657 (N_8657,N_1481,N_2999);
xor U8658 (N_8658,N_4022,N_4432);
nand U8659 (N_8659,N_666,N_331);
nor U8660 (N_8660,N_2237,N_2531);
and U8661 (N_8661,N_2693,N_1269);
and U8662 (N_8662,N_3655,N_1706);
nor U8663 (N_8663,N_4762,N_3919);
nand U8664 (N_8664,N_3925,N_2214);
and U8665 (N_8665,N_4108,N_2125);
nand U8666 (N_8666,N_3836,N_2072);
or U8667 (N_8667,N_3255,N_4153);
and U8668 (N_8668,N_117,N_757);
nor U8669 (N_8669,N_684,N_920);
or U8670 (N_8670,N_3233,N_4687);
xnor U8671 (N_8671,N_1115,N_2605);
nand U8672 (N_8672,N_839,N_3155);
xnor U8673 (N_8673,N_4992,N_1885);
nand U8674 (N_8674,N_4715,N_3643);
and U8675 (N_8675,N_1,N_2370);
and U8676 (N_8676,N_4987,N_4075);
xor U8677 (N_8677,N_4729,N_220);
xnor U8678 (N_8678,N_878,N_1351);
nor U8679 (N_8679,N_3693,N_1018);
and U8680 (N_8680,N_3576,N_3540);
or U8681 (N_8681,N_4919,N_1483);
or U8682 (N_8682,N_2402,N_2661);
and U8683 (N_8683,N_2651,N_2206);
or U8684 (N_8684,N_1968,N_3233);
or U8685 (N_8685,N_303,N_3483);
and U8686 (N_8686,N_249,N_4258);
xnor U8687 (N_8687,N_3112,N_2797);
and U8688 (N_8688,N_1301,N_2725);
xor U8689 (N_8689,N_12,N_233);
and U8690 (N_8690,N_280,N_126);
and U8691 (N_8691,N_666,N_2463);
or U8692 (N_8692,N_1653,N_661);
and U8693 (N_8693,N_1,N_4003);
and U8694 (N_8694,N_3261,N_4454);
nor U8695 (N_8695,N_431,N_3250);
and U8696 (N_8696,N_476,N_2440);
or U8697 (N_8697,N_1529,N_3785);
nor U8698 (N_8698,N_4325,N_2867);
or U8699 (N_8699,N_3060,N_4997);
xnor U8700 (N_8700,N_833,N_4692);
nand U8701 (N_8701,N_12,N_4311);
or U8702 (N_8702,N_435,N_952);
nand U8703 (N_8703,N_2887,N_2412);
xor U8704 (N_8704,N_1823,N_2030);
nor U8705 (N_8705,N_3879,N_826);
nor U8706 (N_8706,N_1367,N_1048);
nor U8707 (N_8707,N_2970,N_4656);
or U8708 (N_8708,N_4484,N_671);
nand U8709 (N_8709,N_2468,N_1919);
and U8710 (N_8710,N_3868,N_1420);
nand U8711 (N_8711,N_1517,N_756);
nor U8712 (N_8712,N_3595,N_2078);
nand U8713 (N_8713,N_4192,N_613);
or U8714 (N_8714,N_4867,N_2198);
or U8715 (N_8715,N_282,N_3705);
and U8716 (N_8716,N_4928,N_3973);
nand U8717 (N_8717,N_4268,N_564);
nor U8718 (N_8718,N_4539,N_4456);
or U8719 (N_8719,N_4647,N_140);
nor U8720 (N_8720,N_979,N_2123);
and U8721 (N_8721,N_46,N_2864);
and U8722 (N_8722,N_1440,N_1015);
and U8723 (N_8723,N_2675,N_1322);
xnor U8724 (N_8724,N_3486,N_1814);
nand U8725 (N_8725,N_1585,N_4239);
nand U8726 (N_8726,N_1662,N_3729);
xor U8727 (N_8727,N_2646,N_1220);
xnor U8728 (N_8728,N_2554,N_4634);
or U8729 (N_8729,N_4346,N_4084);
nor U8730 (N_8730,N_3627,N_274);
nor U8731 (N_8731,N_1645,N_3279);
xor U8732 (N_8732,N_2733,N_3700);
or U8733 (N_8733,N_1479,N_4306);
nor U8734 (N_8734,N_2763,N_3304);
xnor U8735 (N_8735,N_4354,N_3479);
xor U8736 (N_8736,N_3272,N_972);
and U8737 (N_8737,N_4696,N_3476);
and U8738 (N_8738,N_3997,N_606);
nand U8739 (N_8739,N_1159,N_3615);
or U8740 (N_8740,N_3640,N_4752);
or U8741 (N_8741,N_642,N_1082);
or U8742 (N_8742,N_4873,N_828);
nand U8743 (N_8743,N_181,N_2135);
and U8744 (N_8744,N_3520,N_3277);
xnor U8745 (N_8745,N_1193,N_1897);
xnor U8746 (N_8746,N_50,N_3284);
nand U8747 (N_8747,N_3430,N_2150);
and U8748 (N_8748,N_4120,N_567);
nor U8749 (N_8749,N_1280,N_4082);
xnor U8750 (N_8750,N_1477,N_4122);
nand U8751 (N_8751,N_1368,N_1155);
or U8752 (N_8752,N_1575,N_362);
nand U8753 (N_8753,N_2423,N_4118);
and U8754 (N_8754,N_1845,N_362);
xnor U8755 (N_8755,N_1107,N_516);
nand U8756 (N_8756,N_1720,N_1642);
xor U8757 (N_8757,N_955,N_4168);
and U8758 (N_8758,N_2924,N_4969);
xnor U8759 (N_8759,N_4265,N_2666);
nor U8760 (N_8760,N_1105,N_2384);
or U8761 (N_8761,N_4438,N_536);
or U8762 (N_8762,N_3400,N_4054);
nor U8763 (N_8763,N_4129,N_3123);
nand U8764 (N_8764,N_2129,N_4287);
nand U8765 (N_8765,N_212,N_1603);
xor U8766 (N_8766,N_739,N_2280);
and U8767 (N_8767,N_3609,N_3354);
or U8768 (N_8768,N_2479,N_560);
nor U8769 (N_8769,N_2647,N_1086);
nand U8770 (N_8770,N_466,N_3693);
or U8771 (N_8771,N_2673,N_2358);
nor U8772 (N_8772,N_4678,N_2135);
nand U8773 (N_8773,N_2047,N_4846);
or U8774 (N_8774,N_2630,N_2587);
xnor U8775 (N_8775,N_3060,N_3271);
or U8776 (N_8776,N_982,N_2711);
and U8777 (N_8777,N_173,N_3920);
nand U8778 (N_8778,N_1552,N_994);
nand U8779 (N_8779,N_1449,N_514);
nor U8780 (N_8780,N_70,N_4654);
nor U8781 (N_8781,N_1980,N_1656);
nor U8782 (N_8782,N_947,N_1201);
and U8783 (N_8783,N_3343,N_4380);
or U8784 (N_8784,N_2122,N_2256);
xor U8785 (N_8785,N_3863,N_850);
or U8786 (N_8786,N_814,N_1664);
and U8787 (N_8787,N_4759,N_1378);
nor U8788 (N_8788,N_382,N_1660);
or U8789 (N_8789,N_2083,N_818);
xnor U8790 (N_8790,N_3508,N_707);
xnor U8791 (N_8791,N_2412,N_4679);
nand U8792 (N_8792,N_553,N_3377);
or U8793 (N_8793,N_370,N_1761);
xnor U8794 (N_8794,N_2935,N_3938);
xnor U8795 (N_8795,N_330,N_2269);
nand U8796 (N_8796,N_246,N_39);
nor U8797 (N_8797,N_3653,N_1395);
nand U8798 (N_8798,N_149,N_3137);
or U8799 (N_8799,N_3450,N_484);
or U8800 (N_8800,N_2608,N_4270);
xnor U8801 (N_8801,N_1012,N_1339);
or U8802 (N_8802,N_4181,N_4697);
nand U8803 (N_8803,N_1900,N_2406);
nand U8804 (N_8804,N_4949,N_562);
and U8805 (N_8805,N_1754,N_84);
nor U8806 (N_8806,N_3604,N_4923);
or U8807 (N_8807,N_1448,N_4861);
xnor U8808 (N_8808,N_601,N_79);
or U8809 (N_8809,N_3009,N_271);
xor U8810 (N_8810,N_3518,N_3848);
and U8811 (N_8811,N_462,N_2322);
nand U8812 (N_8812,N_4230,N_540);
or U8813 (N_8813,N_2737,N_1881);
xnor U8814 (N_8814,N_4541,N_3810);
or U8815 (N_8815,N_878,N_3467);
or U8816 (N_8816,N_2287,N_3717);
nand U8817 (N_8817,N_4617,N_4531);
nand U8818 (N_8818,N_4686,N_4112);
nand U8819 (N_8819,N_500,N_4819);
nand U8820 (N_8820,N_3330,N_3620);
or U8821 (N_8821,N_788,N_1423);
nor U8822 (N_8822,N_2751,N_2037);
or U8823 (N_8823,N_1168,N_3827);
nor U8824 (N_8824,N_3505,N_3558);
and U8825 (N_8825,N_4684,N_2567);
nand U8826 (N_8826,N_3628,N_4535);
nor U8827 (N_8827,N_3387,N_4957);
or U8828 (N_8828,N_1830,N_2307);
xor U8829 (N_8829,N_3464,N_4185);
and U8830 (N_8830,N_2145,N_2269);
and U8831 (N_8831,N_2117,N_3110);
nor U8832 (N_8832,N_2732,N_4164);
and U8833 (N_8833,N_1621,N_4478);
xor U8834 (N_8834,N_2155,N_1983);
and U8835 (N_8835,N_4975,N_2276);
nand U8836 (N_8836,N_1557,N_1194);
or U8837 (N_8837,N_758,N_3726);
or U8838 (N_8838,N_1978,N_2069);
or U8839 (N_8839,N_1055,N_861);
or U8840 (N_8840,N_831,N_1236);
nand U8841 (N_8841,N_3559,N_1307);
nand U8842 (N_8842,N_3419,N_1769);
or U8843 (N_8843,N_3007,N_4334);
and U8844 (N_8844,N_3546,N_1890);
xor U8845 (N_8845,N_1515,N_1725);
and U8846 (N_8846,N_812,N_436);
and U8847 (N_8847,N_873,N_3985);
or U8848 (N_8848,N_495,N_2849);
nand U8849 (N_8849,N_1681,N_4237);
or U8850 (N_8850,N_3712,N_4084);
xor U8851 (N_8851,N_4321,N_4071);
nand U8852 (N_8852,N_2780,N_4198);
nand U8853 (N_8853,N_3700,N_511);
or U8854 (N_8854,N_3107,N_348);
nor U8855 (N_8855,N_115,N_2994);
xor U8856 (N_8856,N_274,N_1736);
or U8857 (N_8857,N_4006,N_3331);
nor U8858 (N_8858,N_3246,N_4243);
and U8859 (N_8859,N_3760,N_4949);
and U8860 (N_8860,N_505,N_4641);
or U8861 (N_8861,N_1272,N_147);
nand U8862 (N_8862,N_2749,N_3715);
nor U8863 (N_8863,N_3816,N_2392);
nor U8864 (N_8864,N_1877,N_1022);
and U8865 (N_8865,N_127,N_658);
nor U8866 (N_8866,N_1737,N_237);
or U8867 (N_8867,N_2567,N_1082);
xnor U8868 (N_8868,N_3955,N_584);
or U8869 (N_8869,N_1657,N_3353);
and U8870 (N_8870,N_2025,N_3880);
nand U8871 (N_8871,N_207,N_3130);
and U8872 (N_8872,N_2126,N_3862);
or U8873 (N_8873,N_3323,N_4188);
xor U8874 (N_8874,N_4729,N_2266);
xnor U8875 (N_8875,N_3088,N_1751);
xnor U8876 (N_8876,N_2102,N_1669);
or U8877 (N_8877,N_2421,N_4512);
or U8878 (N_8878,N_2771,N_2431);
nor U8879 (N_8879,N_658,N_911);
or U8880 (N_8880,N_3653,N_2507);
nand U8881 (N_8881,N_4825,N_148);
nor U8882 (N_8882,N_4694,N_284);
and U8883 (N_8883,N_143,N_2360);
and U8884 (N_8884,N_1388,N_4903);
xnor U8885 (N_8885,N_3428,N_3380);
nand U8886 (N_8886,N_3684,N_4433);
or U8887 (N_8887,N_1913,N_3398);
xor U8888 (N_8888,N_1030,N_4353);
and U8889 (N_8889,N_2569,N_3120);
and U8890 (N_8890,N_4211,N_1468);
nand U8891 (N_8891,N_3797,N_2656);
and U8892 (N_8892,N_4723,N_288);
and U8893 (N_8893,N_584,N_500);
or U8894 (N_8894,N_650,N_739);
nand U8895 (N_8895,N_2684,N_4993);
or U8896 (N_8896,N_195,N_4794);
and U8897 (N_8897,N_1193,N_2686);
or U8898 (N_8898,N_1775,N_2174);
or U8899 (N_8899,N_4485,N_3456);
xor U8900 (N_8900,N_4357,N_1848);
and U8901 (N_8901,N_27,N_4073);
xnor U8902 (N_8902,N_2173,N_3375);
or U8903 (N_8903,N_4262,N_1274);
and U8904 (N_8904,N_4809,N_1281);
and U8905 (N_8905,N_4103,N_806);
and U8906 (N_8906,N_3751,N_2834);
nor U8907 (N_8907,N_276,N_3748);
xor U8908 (N_8908,N_3750,N_3633);
or U8909 (N_8909,N_3589,N_799);
nor U8910 (N_8910,N_3745,N_237);
nor U8911 (N_8911,N_1138,N_513);
nor U8912 (N_8912,N_3923,N_3772);
nand U8913 (N_8913,N_4141,N_3888);
nand U8914 (N_8914,N_3278,N_3886);
nor U8915 (N_8915,N_311,N_3166);
nand U8916 (N_8916,N_1330,N_1161);
and U8917 (N_8917,N_4683,N_1726);
nor U8918 (N_8918,N_3610,N_4155);
and U8919 (N_8919,N_4886,N_474);
nand U8920 (N_8920,N_3130,N_311);
xnor U8921 (N_8921,N_4724,N_381);
nor U8922 (N_8922,N_2328,N_3642);
nor U8923 (N_8923,N_4265,N_458);
nand U8924 (N_8924,N_2178,N_221);
and U8925 (N_8925,N_180,N_2550);
and U8926 (N_8926,N_2605,N_2905);
nor U8927 (N_8927,N_1988,N_441);
and U8928 (N_8928,N_1413,N_13);
xor U8929 (N_8929,N_2304,N_4781);
nor U8930 (N_8930,N_4236,N_1938);
xnor U8931 (N_8931,N_2942,N_199);
nor U8932 (N_8932,N_3551,N_4891);
or U8933 (N_8933,N_2031,N_4639);
or U8934 (N_8934,N_265,N_902);
nor U8935 (N_8935,N_4732,N_2844);
or U8936 (N_8936,N_2546,N_1236);
nor U8937 (N_8937,N_2879,N_3613);
and U8938 (N_8938,N_2189,N_1771);
xnor U8939 (N_8939,N_4032,N_1965);
or U8940 (N_8940,N_83,N_2078);
xnor U8941 (N_8941,N_2094,N_276);
nor U8942 (N_8942,N_4953,N_1595);
and U8943 (N_8943,N_1271,N_2281);
and U8944 (N_8944,N_4779,N_3986);
xnor U8945 (N_8945,N_3757,N_3562);
nor U8946 (N_8946,N_3376,N_1847);
and U8947 (N_8947,N_2232,N_3709);
nor U8948 (N_8948,N_234,N_1692);
xnor U8949 (N_8949,N_1478,N_4610);
nand U8950 (N_8950,N_4535,N_1953);
or U8951 (N_8951,N_2466,N_216);
and U8952 (N_8952,N_2694,N_420);
or U8953 (N_8953,N_4218,N_4979);
and U8954 (N_8954,N_786,N_4698);
nand U8955 (N_8955,N_3857,N_3022);
nand U8956 (N_8956,N_3744,N_224);
nand U8957 (N_8957,N_971,N_3086);
or U8958 (N_8958,N_2651,N_4926);
nand U8959 (N_8959,N_2701,N_1649);
or U8960 (N_8960,N_1416,N_1610);
or U8961 (N_8961,N_1044,N_708);
nor U8962 (N_8962,N_653,N_2393);
or U8963 (N_8963,N_1591,N_4545);
or U8964 (N_8964,N_4009,N_1211);
or U8965 (N_8965,N_390,N_1334);
or U8966 (N_8966,N_1767,N_947);
nand U8967 (N_8967,N_3935,N_2372);
or U8968 (N_8968,N_4177,N_1609);
or U8969 (N_8969,N_1948,N_1259);
xnor U8970 (N_8970,N_834,N_1064);
xnor U8971 (N_8971,N_3076,N_4384);
nand U8972 (N_8972,N_673,N_4818);
nor U8973 (N_8973,N_714,N_4083);
xor U8974 (N_8974,N_1698,N_2921);
nand U8975 (N_8975,N_3510,N_134);
xor U8976 (N_8976,N_3464,N_3842);
or U8977 (N_8977,N_2623,N_4750);
nand U8978 (N_8978,N_1714,N_3790);
xnor U8979 (N_8979,N_4217,N_3348);
or U8980 (N_8980,N_1302,N_2959);
and U8981 (N_8981,N_574,N_2807);
xnor U8982 (N_8982,N_4465,N_4742);
nand U8983 (N_8983,N_2949,N_3431);
and U8984 (N_8984,N_3783,N_3162);
xor U8985 (N_8985,N_1007,N_4584);
nor U8986 (N_8986,N_2331,N_860);
and U8987 (N_8987,N_2436,N_4885);
or U8988 (N_8988,N_4539,N_239);
nor U8989 (N_8989,N_43,N_3161);
and U8990 (N_8990,N_338,N_2284);
or U8991 (N_8991,N_1900,N_2699);
xnor U8992 (N_8992,N_4403,N_84);
nor U8993 (N_8993,N_2718,N_3575);
nand U8994 (N_8994,N_2244,N_406);
and U8995 (N_8995,N_35,N_2028);
xnor U8996 (N_8996,N_4061,N_1085);
nand U8997 (N_8997,N_1228,N_3756);
and U8998 (N_8998,N_2344,N_1271);
nand U8999 (N_8999,N_1452,N_1736);
xor U9000 (N_9000,N_291,N_1666);
and U9001 (N_9001,N_4040,N_2531);
nor U9002 (N_9002,N_3305,N_1859);
nor U9003 (N_9003,N_1552,N_1449);
or U9004 (N_9004,N_2581,N_4068);
nor U9005 (N_9005,N_4488,N_2627);
or U9006 (N_9006,N_1229,N_3941);
nand U9007 (N_9007,N_2330,N_1577);
or U9008 (N_9008,N_2335,N_910);
xnor U9009 (N_9009,N_2353,N_1075);
nand U9010 (N_9010,N_179,N_635);
or U9011 (N_9011,N_2970,N_1597);
nor U9012 (N_9012,N_150,N_3314);
nand U9013 (N_9013,N_2914,N_4480);
and U9014 (N_9014,N_2785,N_172);
nor U9015 (N_9015,N_1488,N_4637);
xor U9016 (N_9016,N_3738,N_3016);
or U9017 (N_9017,N_3221,N_124);
and U9018 (N_9018,N_3384,N_3071);
or U9019 (N_9019,N_4871,N_165);
nand U9020 (N_9020,N_2244,N_672);
xnor U9021 (N_9021,N_868,N_4015);
xor U9022 (N_9022,N_3371,N_3085);
nor U9023 (N_9023,N_3515,N_197);
nand U9024 (N_9024,N_1035,N_2923);
nor U9025 (N_9025,N_2686,N_4044);
xor U9026 (N_9026,N_2533,N_4575);
nand U9027 (N_9027,N_4940,N_3378);
xnor U9028 (N_9028,N_3020,N_2207);
nor U9029 (N_9029,N_4686,N_2150);
nor U9030 (N_9030,N_2604,N_61);
or U9031 (N_9031,N_3293,N_3682);
and U9032 (N_9032,N_643,N_2829);
or U9033 (N_9033,N_1364,N_1850);
nor U9034 (N_9034,N_1016,N_4870);
nor U9035 (N_9035,N_4645,N_1955);
or U9036 (N_9036,N_1108,N_4545);
and U9037 (N_9037,N_2601,N_3495);
nand U9038 (N_9038,N_4181,N_3171);
nand U9039 (N_9039,N_4702,N_3161);
xor U9040 (N_9040,N_2407,N_2505);
xnor U9041 (N_9041,N_1474,N_1001);
nand U9042 (N_9042,N_4281,N_777);
and U9043 (N_9043,N_560,N_1905);
nand U9044 (N_9044,N_4004,N_3167);
xnor U9045 (N_9045,N_3419,N_4685);
nand U9046 (N_9046,N_4263,N_441);
nand U9047 (N_9047,N_3203,N_367);
nor U9048 (N_9048,N_4418,N_4408);
nand U9049 (N_9049,N_1647,N_776);
nand U9050 (N_9050,N_1918,N_534);
nor U9051 (N_9051,N_136,N_4657);
nor U9052 (N_9052,N_1760,N_3126);
and U9053 (N_9053,N_1155,N_340);
nand U9054 (N_9054,N_3998,N_3853);
nand U9055 (N_9055,N_1539,N_2343);
nor U9056 (N_9056,N_436,N_4478);
or U9057 (N_9057,N_1847,N_3347);
xor U9058 (N_9058,N_4326,N_2516);
xor U9059 (N_9059,N_712,N_3487);
xnor U9060 (N_9060,N_4690,N_2760);
and U9061 (N_9061,N_804,N_183);
or U9062 (N_9062,N_3715,N_2534);
nand U9063 (N_9063,N_4588,N_1042);
nor U9064 (N_9064,N_4534,N_2691);
xor U9065 (N_9065,N_304,N_1968);
or U9066 (N_9066,N_761,N_2404);
and U9067 (N_9067,N_1446,N_4379);
or U9068 (N_9068,N_1904,N_1936);
nand U9069 (N_9069,N_1217,N_3821);
xor U9070 (N_9070,N_4062,N_4515);
and U9071 (N_9071,N_3931,N_3691);
nand U9072 (N_9072,N_1319,N_4906);
or U9073 (N_9073,N_1640,N_4658);
or U9074 (N_9074,N_1346,N_1528);
xor U9075 (N_9075,N_2219,N_1205);
nand U9076 (N_9076,N_235,N_4301);
or U9077 (N_9077,N_2784,N_924);
or U9078 (N_9078,N_187,N_4044);
nor U9079 (N_9079,N_147,N_2176);
and U9080 (N_9080,N_4475,N_1063);
nor U9081 (N_9081,N_198,N_3675);
or U9082 (N_9082,N_2257,N_4765);
nand U9083 (N_9083,N_1767,N_1804);
or U9084 (N_9084,N_3056,N_1627);
and U9085 (N_9085,N_2791,N_4241);
nand U9086 (N_9086,N_4819,N_2018);
or U9087 (N_9087,N_2855,N_1158);
xor U9088 (N_9088,N_3606,N_1014);
nor U9089 (N_9089,N_3428,N_1070);
nand U9090 (N_9090,N_3766,N_3912);
and U9091 (N_9091,N_3996,N_3774);
nor U9092 (N_9092,N_1323,N_1099);
or U9093 (N_9093,N_4062,N_4384);
or U9094 (N_9094,N_2041,N_827);
nand U9095 (N_9095,N_584,N_2614);
and U9096 (N_9096,N_2764,N_2940);
and U9097 (N_9097,N_2382,N_361);
and U9098 (N_9098,N_2614,N_175);
and U9099 (N_9099,N_497,N_4204);
xor U9100 (N_9100,N_4870,N_1829);
or U9101 (N_9101,N_624,N_773);
or U9102 (N_9102,N_439,N_1139);
nand U9103 (N_9103,N_3948,N_1949);
xor U9104 (N_9104,N_4940,N_2716);
and U9105 (N_9105,N_2678,N_3055);
nand U9106 (N_9106,N_309,N_4476);
nand U9107 (N_9107,N_4009,N_4820);
and U9108 (N_9108,N_1698,N_4239);
and U9109 (N_9109,N_1635,N_383);
nor U9110 (N_9110,N_3692,N_1757);
nor U9111 (N_9111,N_1979,N_1671);
nor U9112 (N_9112,N_3663,N_1499);
nor U9113 (N_9113,N_1160,N_3113);
and U9114 (N_9114,N_3639,N_2570);
nand U9115 (N_9115,N_2682,N_718);
or U9116 (N_9116,N_3883,N_3189);
nand U9117 (N_9117,N_4586,N_4363);
nor U9118 (N_9118,N_2759,N_4156);
nand U9119 (N_9119,N_3418,N_2357);
or U9120 (N_9120,N_3428,N_4751);
and U9121 (N_9121,N_2539,N_4554);
nor U9122 (N_9122,N_1529,N_4270);
or U9123 (N_9123,N_2371,N_2236);
nor U9124 (N_9124,N_742,N_810);
nand U9125 (N_9125,N_1147,N_3477);
and U9126 (N_9126,N_3688,N_1338);
xor U9127 (N_9127,N_4089,N_3108);
nor U9128 (N_9128,N_2669,N_346);
or U9129 (N_9129,N_3133,N_4090);
and U9130 (N_9130,N_514,N_4528);
and U9131 (N_9131,N_3331,N_3457);
nor U9132 (N_9132,N_1316,N_4239);
xnor U9133 (N_9133,N_4057,N_3713);
or U9134 (N_9134,N_1279,N_2718);
and U9135 (N_9135,N_1643,N_1466);
xor U9136 (N_9136,N_2848,N_864);
nor U9137 (N_9137,N_2780,N_726);
xor U9138 (N_9138,N_4383,N_2787);
nor U9139 (N_9139,N_2892,N_1187);
nor U9140 (N_9140,N_375,N_311);
nor U9141 (N_9141,N_131,N_3972);
or U9142 (N_9142,N_4556,N_4585);
xor U9143 (N_9143,N_1253,N_2508);
xnor U9144 (N_9144,N_2350,N_4260);
or U9145 (N_9145,N_1742,N_2893);
or U9146 (N_9146,N_4318,N_2171);
or U9147 (N_9147,N_3255,N_1826);
xor U9148 (N_9148,N_208,N_4963);
nand U9149 (N_9149,N_4925,N_3743);
or U9150 (N_9150,N_4436,N_804);
nor U9151 (N_9151,N_4003,N_362);
xnor U9152 (N_9152,N_4755,N_2507);
nor U9153 (N_9153,N_2474,N_2087);
or U9154 (N_9154,N_997,N_658);
or U9155 (N_9155,N_851,N_4658);
xnor U9156 (N_9156,N_1195,N_1853);
or U9157 (N_9157,N_384,N_4593);
or U9158 (N_9158,N_4835,N_2897);
xnor U9159 (N_9159,N_618,N_2688);
xor U9160 (N_9160,N_1314,N_3704);
and U9161 (N_9161,N_4376,N_986);
or U9162 (N_9162,N_1639,N_4294);
nand U9163 (N_9163,N_275,N_1865);
nor U9164 (N_9164,N_506,N_4153);
nand U9165 (N_9165,N_4756,N_961);
xnor U9166 (N_9166,N_2099,N_2850);
nand U9167 (N_9167,N_3900,N_330);
nand U9168 (N_9168,N_2804,N_1871);
nor U9169 (N_9169,N_587,N_650);
and U9170 (N_9170,N_3385,N_3114);
or U9171 (N_9171,N_3779,N_4926);
nand U9172 (N_9172,N_543,N_1797);
xnor U9173 (N_9173,N_2409,N_4440);
xor U9174 (N_9174,N_2853,N_2010);
nor U9175 (N_9175,N_4511,N_3788);
nor U9176 (N_9176,N_1330,N_3602);
nand U9177 (N_9177,N_1076,N_2173);
and U9178 (N_9178,N_4220,N_3618);
nand U9179 (N_9179,N_1715,N_3537);
nor U9180 (N_9180,N_1673,N_3220);
nor U9181 (N_9181,N_4148,N_378);
nand U9182 (N_9182,N_3106,N_247);
or U9183 (N_9183,N_2523,N_1431);
xor U9184 (N_9184,N_1813,N_2418);
xnor U9185 (N_9185,N_2539,N_2600);
or U9186 (N_9186,N_2119,N_3384);
nand U9187 (N_9187,N_286,N_3750);
nor U9188 (N_9188,N_2279,N_862);
or U9189 (N_9189,N_1245,N_3699);
nand U9190 (N_9190,N_4351,N_4602);
xor U9191 (N_9191,N_4642,N_1216);
xnor U9192 (N_9192,N_242,N_3752);
and U9193 (N_9193,N_4679,N_1004);
nor U9194 (N_9194,N_23,N_1574);
nand U9195 (N_9195,N_1645,N_1254);
nor U9196 (N_9196,N_1571,N_1428);
nand U9197 (N_9197,N_1587,N_3168);
xnor U9198 (N_9198,N_3468,N_1428);
and U9199 (N_9199,N_4569,N_3015);
and U9200 (N_9200,N_4760,N_566);
nand U9201 (N_9201,N_4773,N_3047);
nor U9202 (N_9202,N_1605,N_2100);
nor U9203 (N_9203,N_2328,N_1247);
or U9204 (N_9204,N_2070,N_259);
xor U9205 (N_9205,N_3034,N_4440);
nor U9206 (N_9206,N_1253,N_2680);
and U9207 (N_9207,N_1714,N_4004);
xnor U9208 (N_9208,N_1746,N_303);
nor U9209 (N_9209,N_3541,N_608);
or U9210 (N_9210,N_3402,N_2414);
nand U9211 (N_9211,N_2858,N_2445);
xor U9212 (N_9212,N_3649,N_4967);
nand U9213 (N_9213,N_903,N_3159);
nor U9214 (N_9214,N_1689,N_206);
and U9215 (N_9215,N_1738,N_633);
and U9216 (N_9216,N_1518,N_2613);
and U9217 (N_9217,N_4492,N_3609);
nand U9218 (N_9218,N_4157,N_4049);
nor U9219 (N_9219,N_4831,N_1072);
or U9220 (N_9220,N_822,N_1193);
xor U9221 (N_9221,N_3677,N_666);
xor U9222 (N_9222,N_888,N_2647);
xor U9223 (N_9223,N_1111,N_4015);
nand U9224 (N_9224,N_536,N_4922);
nand U9225 (N_9225,N_3149,N_3322);
nand U9226 (N_9226,N_92,N_2781);
and U9227 (N_9227,N_2425,N_3915);
nand U9228 (N_9228,N_3068,N_3965);
or U9229 (N_9229,N_2008,N_648);
and U9230 (N_9230,N_3836,N_4988);
and U9231 (N_9231,N_80,N_478);
nand U9232 (N_9232,N_601,N_2760);
nand U9233 (N_9233,N_2910,N_3073);
nand U9234 (N_9234,N_2,N_3799);
and U9235 (N_9235,N_3462,N_3946);
xor U9236 (N_9236,N_4993,N_3974);
and U9237 (N_9237,N_3961,N_4090);
nor U9238 (N_9238,N_4318,N_1222);
or U9239 (N_9239,N_4311,N_1987);
and U9240 (N_9240,N_88,N_1709);
and U9241 (N_9241,N_2797,N_189);
or U9242 (N_9242,N_3009,N_3319);
nand U9243 (N_9243,N_4092,N_2633);
or U9244 (N_9244,N_897,N_714);
and U9245 (N_9245,N_4137,N_4395);
or U9246 (N_9246,N_4925,N_3733);
xnor U9247 (N_9247,N_428,N_990);
xnor U9248 (N_9248,N_932,N_538);
and U9249 (N_9249,N_1125,N_2500);
nor U9250 (N_9250,N_4763,N_1665);
xor U9251 (N_9251,N_2103,N_4424);
or U9252 (N_9252,N_2250,N_3105);
nor U9253 (N_9253,N_2161,N_4001);
or U9254 (N_9254,N_4151,N_2762);
nand U9255 (N_9255,N_1403,N_3395);
xnor U9256 (N_9256,N_653,N_2423);
nor U9257 (N_9257,N_3661,N_2956);
nand U9258 (N_9258,N_4181,N_4838);
nand U9259 (N_9259,N_458,N_2832);
xnor U9260 (N_9260,N_2477,N_18);
nor U9261 (N_9261,N_2312,N_1040);
xnor U9262 (N_9262,N_1014,N_2079);
xnor U9263 (N_9263,N_4386,N_1885);
and U9264 (N_9264,N_4999,N_1845);
nand U9265 (N_9265,N_680,N_1720);
and U9266 (N_9266,N_1471,N_3176);
or U9267 (N_9267,N_432,N_4353);
nand U9268 (N_9268,N_4961,N_4041);
or U9269 (N_9269,N_3168,N_1971);
xor U9270 (N_9270,N_1287,N_3657);
or U9271 (N_9271,N_1171,N_782);
and U9272 (N_9272,N_48,N_1900);
nand U9273 (N_9273,N_4576,N_737);
and U9274 (N_9274,N_1651,N_1763);
nor U9275 (N_9275,N_818,N_3165);
nor U9276 (N_9276,N_588,N_2037);
and U9277 (N_9277,N_4940,N_3499);
nor U9278 (N_9278,N_3304,N_3218);
xnor U9279 (N_9279,N_2431,N_3798);
and U9280 (N_9280,N_3669,N_1917);
nor U9281 (N_9281,N_4345,N_2034);
nand U9282 (N_9282,N_1378,N_1597);
nand U9283 (N_9283,N_4469,N_4713);
xor U9284 (N_9284,N_811,N_1143);
nor U9285 (N_9285,N_2493,N_4681);
or U9286 (N_9286,N_2220,N_4950);
or U9287 (N_9287,N_728,N_4603);
and U9288 (N_9288,N_1246,N_91);
nand U9289 (N_9289,N_1960,N_4031);
and U9290 (N_9290,N_644,N_380);
or U9291 (N_9291,N_4395,N_2443);
xnor U9292 (N_9292,N_4820,N_3386);
nand U9293 (N_9293,N_3535,N_748);
xnor U9294 (N_9294,N_4740,N_875);
xnor U9295 (N_9295,N_2517,N_1242);
or U9296 (N_9296,N_2826,N_2501);
nor U9297 (N_9297,N_3605,N_1123);
or U9298 (N_9298,N_4939,N_2283);
and U9299 (N_9299,N_746,N_4729);
xnor U9300 (N_9300,N_1027,N_1033);
nand U9301 (N_9301,N_1351,N_2449);
or U9302 (N_9302,N_655,N_3169);
or U9303 (N_9303,N_1066,N_1392);
xor U9304 (N_9304,N_2304,N_702);
and U9305 (N_9305,N_1028,N_473);
xnor U9306 (N_9306,N_2802,N_388);
nor U9307 (N_9307,N_2202,N_2884);
and U9308 (N_9308,N_3784,N_972);
nand U9309 (N_9309,N_511,N_3734);
nand U9310 (N_9310,N_4043,N_3983);
nand U9311 (N_9311,N_1096,N_3163);
xnor U9312 (N_9312,N_3688,N_1595);
or U9313 (N_9313,N_4682,N_754);
nand U9314 (N_9314,N_4927,N_2782);
or U9315 (N_9315,N_2103,N_4861);
or U9316 (N_9316,N_3502,N_4737);
and U9317 (N_9317,N_194,N_91);
xor U9318 (N_9318,N_2921,N_1211);
and U9319 (N_9319,N_1386,N_2714);
nand U9320 (N_9320,N_4974,N_3851);
xor U9321 (N_9321,N_2389,N_2504);
nor U9322 (N_9322,N_4974,N_438);
nand U9323 (N_9323,N_2255,N_491);
nor U9324 (N_9324,N_3506,N_1848);
and U9325 (N_9325,N_1819,N_3415);
nor U9326 (N_9326,N_4606,N_4653);
xnor U9327 (N_9327,N_2798,N_207);
nand U9328 (N_9328,N_3099,N_2241);
or U9329 (N_9329,N_451,N_2131);
nor U9330 (N_9330,N_1155,N_2260);
nor U9331 (N_9331,N_3725,N_1921);
nor U9332 (N_9332,N_4009,N_2287);
nand U9333 (N_9333,N_3553,N_3182);
or U9334 (N_9334,N_792,N_607);
xnor U9335 (N_9335,N_2983,N_713);
xnor U9336 (N_9336,N_1904,N_136);
nor U9337 (N_9337,N_3072,N_96);
and U9338 (N_9338,N_3504,N_3366);
nor U9339 (N_9339,N_3337,N_1336);
xor U9340 (N_9340,N_59,N_1972);
nor U9341 (N_9341,N_4940,N_635);
xor U9342 (N_9342,N_1850,N_4616);
nor U9343 (N_9343,N_1359,N_1583);
xnor U9344 (N_9344,N_314,N_1593);
xnor U9345 (N_9345,N_2625,N_1757);
xnor U9346 (N_9346,N_2951,N_4708);
xor U9347 (N_9347,N_4536,N_2735);
xor U9348 (N_9348,N_1354,N_616);
or U9349 (N_9349,N_3540,N_1213);
and U9350 (N_9350,N_4573,N_392);
xor U9351 (N_9351,N_205,N_4036);
nor U9352 (N_9352,N_1045,N_1456);
nor U9353 (N_9353,N_872,N_1582);
nor U9354 (N_9354,N_1405,N_3959);
or U9355 (N_9355,N_2312,N_2792);
nor U9356 (N_9356,N_2483,N_163);
nor U9357 (N_9357,N_1225,N_2202);
xnor U9358 (N_9358,N_3258,N_4189);
xor U9359 (N_9359,N_4911,N_2573);
xnor U9360 (N_9360,N_1577,N_4228);
nor U9361 (N_9361,N_4586,N_3108);
or U9362 (N_9362,N_691,N_2008);
and U9363 (N_9363,N_424,N_2664);
nor U9364 (N_9364,N_3556,N_218);
and U9365 (N_9365,N_4426,N_3084);
xnor U9366 (N_9366,N_1311,N_1861);
and U9367 (N_9367,N_1569,N_1560);
and U9368 (N_9368,N_1348,N_4464);
nand U9369 (N_9369,N_3453,N_4358);
and U9370 (N_9370,N_3434,N_3328);
nor U9371 (N_9371,N_1031,N_1067);
or U9372 (N_9372,N_1051,N_1749);
and U9373 (N_9373,N_700,N_3202);
xor U9374 (N_9374,N_4283,N_3640);
and U9375 (N_9375,N_112,N_348);
nand U9376 (N_9376,N_2575,N_2538);
nand U9377 (N_9377,N_4854,N_3866);
or U9378 (N_9378,N_4516,N_60);
nand U9379 (N_9379,N_4718,N_1856);
nand U9380 (N_9380,N_858,N_3444);
and U9381 (N_9381,N_3754,N_3454);
xor U9382 (N_9382,N_1198,N_3052);
nand U9383 (N_9383,N_4272,N_4652);
nor U9384 (N_9384,N_1355,N_3419);
nor U9385 (N_9385,N_4173,N_1097);
nand U9386 (N_9386,N_3692,N_4971);
nor U9387 (N_9387,N_2374,N_2553);
nand U9388 (N_9388,N_1196,N_3153);
or U9389 (N_9389,N_3501,N_2345);
nand U9390 (N_9390,N_4896,N_4509);
nand U9391 (N_9391,N_3845,N_3460);
and U9392 (N_9392,N_3471,N_2104);
and U9393 (N_9393,N_4734,N_1815);
nor U9394 (N_9394,N_72,N_135);
nand U9395 (N_9395,N_2025,N_3891);
nand U9396 (N_9396,N_2268,N_274);
or U9397 (N_9397,N_1436,N_3063);
or U9398 (N_9398,N_1411,N_1347);
and U9399 (N_9399,N_2004,N_3555);
and U9400 (N_9400,N_1391,N_572);
xnor U9401 (N_9401,N_4132,N_2570);
xnor U9402 (N_9402,N_2424,N_2852);
and U9403 (N_9403,N_3399,N_2411);
xnor U9404 (N_9404,N_15,N_286);
xor U9405 (N_9405,N_4922,N_2853);
nand U9406 (N_9406,N_3794,N_2401);
nor U9407 (N_9407,N_4516,N_2858);
or U9408 (N_9408,N_1827,N_2882);
nand U9409 (N_9409,N_4788,N_877);
or U9410 (N_9410,N_878,N_592);
xnor U9411 (N_9411,N_1213,N_239);
nor U9412 (N_9412,N_1382,N_3779);
or U9413 (N_9413,N_4647,N_801);
xor U9414 (N_9414,N_1288,N_1326);
nor U9415 (N_9415,N_1791,N_1996);
xor U9416 (N_9416,N_2165,N_2685);
nor U9417 (N_9417,N_893,N_2754);
nor U9418 (N_9418,N_4918,N_4065);
nand U9419 (N_9419,N_2946,N_3221);
or U9420 (N_9420,N_600,N_1624);
and U9421 (N_9421,N_737,N_2830);
or U9422 (N_9422,N_1832,N_1636);
nand U9423 (N_9423,N_1326,N_4139);
nor U9424 (N_9424,N_977,N_760);
and U9425 (N_9425,N_1160,N_850);
nor U9426 (N_9426,N_3438,N_448);
and U9427 (N_9427,N_3194,N_4035);
or U9428 (N_9428,N_2387,N_10);
or U9429 (N_9429,N_3427,N_4868);
nand U9430 (N_9430,N_3629,N_1288);
and U9431 (N_9431,N_373,N_3358);
or U9432 (N_9432,N_4421,N_3940);
or U9433 (N_9433,N_3372,N_2793);
or U9434 (N_9434,N_3601,N_1723);
or U9435 (N_9435,N_142,N_2394);
nand U9436 (N_9436,N_1166,N_1847);
and U9437 (N_9437,N_1493,N_2036);
nand U9438 (N_9438,N_1159,N_1945);
or U9439 (N_9439,N_967,N_3285);
and U9440 (N_9440,N_1794,N_2900);
nand U9441 (N_9441,N_2528,N_1791);
and U9442 (N_9442,N_2855,N_3305);
and U9443 (N_9443,N_2687,N_2981);
and U9444 (N_9444,N_4297,N_1939);
nand U9445 (N_9445,N_2060,N_2688);
nor U9446 (N_9446,N_390,N_865);
and U9447 (N_9447,N_163,N_1016);
xnor U9448 (N_9448,N_3657,N_312);
xor U9449 (N_9449,N_2988,N_596);
and U9450 (N_9450,N_4361,N_3094);
nand U9451 (N_9451,N_161,N_219);
and U9452 (N_9452,N_1355,N_4442);
nor U9453 (N_9453,N_195,N_2754);
nor U9454 (N_9454,N_1035,N_3637);
xor U9455 (N_9455,N_4068,N_2551);
and U9456 (N_9456,N_2378,N_1069);
and U9457 (N_9457,N_3260,N_4495);
and U9458 (N_9458,N_572,N_2023);
or U9459 (N_9459,N_960,N_4946);
nand U9460 (N_9460,N_4458,N_2401);
xnor U9461 (N_9461,N_2805,N_3547);
xor U9462 (N_9462,N_2018,N_4655);
or U9463 (N_9463,N_1344,N_2162);
and U9464 (N_9464,N_1196,N_1859);
or U9465 (N_9465,N_3171,N_3832);
nand U9466 (N_9466,N_404,N_914);
xnor U9467 (N_9467,N_3731,N_25);
and U9468 (N_9468,N_2065,N_2714);
nand U9469 (N_9469,N_2023,N_1401);
or U9470 (N_9470,N_1953,N_3198);
or U9471 (N_9471,N_1730,N_3682);
xor U9472 (N_9472,N_2839,N_1974);
nor U9473 (N_9473,N_3357,N_887);
and U9474 (N_9474,N_3005,N_58);
xnor U9475 (N_9475,N_2321,N_277);
xnor U9476 (N_9476,N_2720,N_3762);
nand U9477 (N_9477,N_4075,N_3823);
nor U9478 (N_9478,N_491,N_1520);
xor U9479 (N_9479,N_3871,N_1972);
or U9480 (N_9480,N_2228,N_1706);
nor U9481 (N_9481,N_4725,N_1931);
nand U9482 (N_9482,N_3575,N_3847);
and U9483 (N_9483,N_4347,N_609);
nor U9484 (N_9484,N_126,N_2948);
nand U9485 (N_9485,N_1411,N_2698);
nand U9486 (N_9486,N_3935,N_1009);
xnor U9487 (N_9487,N_2523,N_3386);
and U9488 (N_9488,N_3979,N_1762);
nor U9489 (N_9489,N_2712,N_3475);
and U9490 (N_9490,N_1375,N_2243);
nand U9491 (N_9491,N_4460,N_2683);
xor U9492 (N_9492,N_388,N_2674);
and U9493 (N_9493,N_3626,N_4847);
nand U9494 (N_9494,N_3273,N_4777);
xnor U9495 (N_9495,N_981,N_2675);
nand U9496 (N_9496,N_3454,N_3706);
nand U9497 (N_9497,N_4532,N_1676);
xor U9498 (N_9498,N_1805,N_4885);
nor U9499 (N_9499,N_978,N_4666);
or U9500 (N_9500,N_3744,N_519);
nor U9501 (N_9501,N_2721,N_2154);
xnor U9502 (N_9502,N_297,N_913);
or U9503 (N_9503,N_1637,N_3317);
nand U9504 (N_9504,N_1358,N_2769);
and U9505 (N_9505,N_4338,N_1708);
or U9506 (N_9506,N_4487,N_2469);
xor U9507 (N_9507,N_472,N_1866);
nor U9508 (N_9508,N_2529,N_4832);
nand U9509 (N_9509,N_3799,N_1738);
and U9510 (N_9510,N_2723,N_107);
nand U9511 (N_9511,N_812,N_1385);
nor U9512 (N_9512,N_40,N_3147);
nor U9513 (N_9513,N_3232,N_983);
nand U9514 (N_9514,N_4034,N_1623);
nand U9515 (N_9515,N_797,N_3593);
nor U9516 (N_9516,N_1818,N_1116);
and U9517 (N_9517,N_4353,N_2152);
and U9518 (N_9518,N_3024,N_2138);
nor U9519 (N_9519,N_1418,N_4170);
xnor U9520 (N_9520,N_2799,N_657);
xor U9521 (N_9521,N_79,N_1073);
xor U9522 (N_9522,N_3919,N_902);
or U9523 (N_9523,N_3685,N_4118);
or U9524 (N_9524,N_3182,N_3610);
xnor U9525 (N_9525,N_2729,N_230);
nand U9526 (N_9526,N_683,N_493);
xor U9527 (N_9527,N_388,N_1152);
nand U9528 (N_9528,N_159,N_523);
and U9529 (N_9529,N_1985,N_1520);
nor U9530 (N_9530,N_2491,N_431);
or U9531 (N_9531,N_2111,N_2385);
nand U9532 (N_9532,N_3411,N_2665);
nand U9533 (N_9533,N_934,N_4477);
xor U9534 (N_9534,N_3698,N_551);
nand U9535 (N_9535,N_2227,N_1970);
xnor U9536 (N_9536,N_286,N_2850);
nor U9537 (N_9537,N_951,N_964);
xnor U9538 (N_9538,N_1397,N_888);
or U9539 (N_9539,N_3866,N_172);
xnor U9540 (N_9540,N_2173,N_1241);
and U9541 (N_9541,N_253,N_3253);
nand U9542 (N_9542,N_111,N_773);
nand U9543 (N_9543,N_1495,N_371);
nor U9544 (N_9544,N_2162,N_4764);
or U9545 (N_9545,N_246,N_3230);
xnor U9546 (N_9546,N_1622,N_3577);
xnor U9547 (N_9547,N_2793,N_640);
or U9548 (N_9548,N_2898,N_2375);
and U9549 (N_9549,N_143,N_1031);
nor U9550 (N_9550,N_750,N_1426);
or U9551 (N_9551,N_2764,N_1914);
xnor U9552 (N_9552,N_3584,N_709);
nand U9553 (N_9553,N_4415,N_1308);
or U9554 (N_9554,N_332,N_2450);
nand U9555 (N_9555,N_660,N_4490);
xor U9556 (N_9556,N_3033,N_3824);
xnor U9557 (N_9557,N_4651,N_2366);
nand U9558 (N_9558,N_4364,N_843);
xor U9559 (N_9559,N_2832,N_4487);
and U9560 (N_9560,N_4343,N_4906);
or U9561 (N_9561,N_4369,N_1065);
or U9562 (N_9562,N_1520,N_1963);
and U9563 (N_9563,N_1389,N_1873);
nor U9564 (N_9564,N_1068,N_2620);
xor U9565 (N_9565,N_2349,N_2609);
nor U9566 (N_9566,N_4414,N_3315);
nand U9567 (N_9567,N_1744,N_4568);
xnor U9568 (N_9568,N_3749,N_2252);
and U9569 (N_9569,N_4908,N_1243);
nor U9570 (N_9570,N_4053,N_46);
nand U9571 (N_9571,N_3994,N_500);
xor U9572 (N_9572,N_167,N_3490);
and U9573 (N_9573,N_3792,N_4419);
nand U9574 (N_9574,N_3458,N_3122);
xor U9575 (N_9575,N_4976,N_1658);
xnor U9576 (N_9576,N_4340,N_772);
and U9577 (N_9577,N_2095,N_379);
or U9578 (N_9578,N_1775,N_3221);
nand U9579 (N_9579,N_1316,N_1942);
nand U9580 (N_9580,N_2966,N_3294);
xnor U9581 (N_9581,N_646,N_3770);
or U9582 (N_9582,N_2083,N_4164);
xor U9583 (N_9583,N_3004,N_1094);
nor U9584 (N_9584,N_662,N_1470);
xor U9585 (N_9585,N_770,N_1535);
nor U9586 (N_9586,N_2039,N_2489);
xnor U9587 (N_9587,N_3253,N_1966);
xnor U9588 (N_9588,N_3798,N_1253);
nor U9589 (N_9589,N_3418,N_4505);
and U9590 (N_9590,N_4888,N_2711);
nor U9591 (N_9591,N_1032,N_143);
nand U9592 (N_9592,N_3921,N_1624);
or U9593 (N_9593,N_1071,N_4373);
nand U9594 (N_9594,N_1872,N_1562);
nor U9595 (N_9595,N_3996,N_3933);
nor U9596 (N_9596,N_2960,N_2562);
nand U9597 (N_9597,N_3845,N_2585);
nand U9598 (N_9598,N_3841,N_1835);
nand U9599 (N_9599,N_4612,N_3137);
or U9600 (N_9600,N_2749,N_2635);
nor U9601 (N_9601,N_4294,N_4847);
and U9602 (N_9602,N_508,N_4573);
or U9603 (N_9603,N_4375,N_1286);
xnor U9604 (N_9604,N_3460,N_3593);
xnor U9605 (N_9605,N_1673,N_3684);
and U9606 (N_9606,N_1026,N_1912);
nor U9607 (N_9607,N_3682,N_1525);
and U9608 (N_9608,N_1817,N_4188);
and U9609 (N_9609,N_4775,N_3761);
and U9610 (N_9610,N_657,N_1126);
nor U9611 (N_9611,N_4075,N_4327);
and U9612 (N_9612,N_144,N_1103);
and U9613 (N_9613,N_1014,N_646);
nor U9614 (N_9614,N_2087,N_3481);
nand U9615 (N_9615,N_2089,N_2792);
nand U9616 (N_9616,N_1050,N_818);
and U9617 (N_9617,N_2324,N_347);
nor U9618 (N_9618,N_3137,N_2387);
xor U9619 (N_9619,N_2454,N_3588);
xnor U9620 (N_9620,N_3589,N_4027);
nand U9621 (N_9621,N_207,N_2461);
nand U9622 (N_9622,N_3564,N_4870);
or U9623 (N_9623,N_531,N_2075);
nand U9624 (N_9624,N_1778,N_4063);
nor U9625 (N_9625,N_2416,N_815);
and U9626 (N_9626,N_706,N_148);
or U9627 (N_9627,N_1361,N_2384);
and U9628 (N_9628,N_3634,N_1670);
and U9629 (N_9629,N_955,N_3992);
xnor U9630 (N_9630,N_1697,N_2982);
or U9631 (N_9631,N_3851,N_2275);
nor U9632 (N_9632,N_4999,N_1652);
xnor U9633 (N_9633,N_3942,N_3155);
and U9634 (N_9634,N_4452,N_3754);
nand U9635 (N_9635,N_2401,N_1156);
xor U9636 (N_9636,N_1811,N_674);
nand U9637 (N_9637,N_4123,N_2902);
nand U9638 (N_9638,N_4734,N_4333);
nor U9639 (N_9639,N_3405,N_4824);
nor U9640 (N_9640,N_4099,N_4744);
and U9641 (N_9641,N_633,N_923);
nor U9642 (N_9642,N_4929,N_4251);
and U9643 (N_9643,N_4279,N_3144);
nor U9644 (N_9644,N_3656,N_3649);
nor U9645 (N_9645,N_1262,N_1808);
or U9646 (N_9646,N_2029,N_4236);
nor U9647 (N_9647,N_1060,N_1583);
and U9648 (N_9648,N_1890,N_1968);
nor U9649 (N_9649,N_4444,N_3720);
xor U9650 (N_9650,N_592,N_4559);
or U9651 (N_9651,N_3458,N_3528);
xor U9652 (N_9652,N_813,N_573);
and U9653 (N_9653,N_1918,N_2348);
xor U9654 (N_9654,N_2335,N_2323);
and U9655 (N_9655,N_4255,N_573);
or U9656 (N_9656,N_4950,N_2343);
or U9657 (N_9657,N_1129,N_1283);
xor U9658 (N_9658,N_4587,N_2095);
xnor U9659 (N_9659,N_3687,N_4948);
and U9660 (N_9660,N_2651,N_2799);
nor U9661 (N_9661,N_256,N_2310);
xnor U9662 (N_9662,N_2052,N_1164);
xnor U9663 (N_9663,N_3128,N_1443);
and U9664 (N_9664,N_631,N_995);
or U9665 (N_9665,N_2477,N_1064);
or U9666 (N_9666,N_736,N_218);
xnor U9667 (N_9667,N_3431,N_146);
nand U9668 (N_9668,N_1925,N_3319);
nand U9669 (N_9669,N_4632,N_2935);
nor U9670 (N_9670,N_4984,N_3814);
nand U9671 (N_9671,N_2021,N_1470);
nand U9672 (N_9672,N_2809,N_2072);
xnor U9673 (N_9673,N_495,N_1287);
xor U9674 (N_9674,N_3061,N_1703);
and U9675 (N_9675,N_2654,N_2653);
xor U9676 (N_9676,N_1784,N_2545);
xnor U9677 (N_9677,N_4664,N_3214);
xnor U9678 (N_9678,N_4298,N_2193);
xnor U9679 (N_9679,N_2123,N_4902);
xnor U9680 (N_9680,N_4171,N_450);
nor U9681 (N_9681,N_1119,N_1043);
and U9682 (N_9682,N_3784,N_4492);
and U9683 (N_9683,N_4563,N_4809);
and U9684 (N_9684,N_4024,N_235);
xor U9685 (N_9685,N_1375,N_3806);
nand U9686 (N_9686,N_2034,N_3609);
nand U9687 (N_9687,N_3538,N_897);
or U9688 (N_9688,N_3528,N_1218);
xnor U9689 (N_9689,N_163,N_1133);
xnor U9690 (N_9690,N_2858,N_1727);
or U9691 (N_9691,N_3536,N_623);
and U9692 (N_9692,N_2531,N_2449);
xor U9693 (N_9693,N_3542,N_2545);
xor U9694 (N_9694,N_2824,N_94);
nor U9695 (N_9695,N_3598,N_3241);
or U9696 (N_9696,N_3130,N_2526);
and U9697 (N_9697,N_1613,N_1618);
nor U9698 (N_9698,N_4951,N_2974);
and U9699 (N_9699,N_3913,N_4894);
and U9700 (N_9700,N_3156,N_4277);
nand U9701 (N_9701,N_2146,N_1705);
and U9702 (N_9702,N_2391,N_3331);
nand U9703 (N_9703,N_4773,N_1497);
nor U9704 (N_9704,N_2079,N_2688);
nor U9705 (N_9705,N_3318,N_2956);
nand U9706 (N_9706,N_3564,N_568);
and U9707 (N_9707,N_2336,N_3895);
or U9708 (N_9708,N_3252,N_4375);
nor U9709 (N_9709,N_3382,N_73);
nand U9710 (N_9710,N_4525,N_4192);
xnor U9711 (N_9711,N_2639,N_1210);
and U9712 (N_9712,N_708,N_2047);
and U9713 (N_9713,N_1983,N_590);
and U9714 (N_9714,N_2610,N_3469);
nor U9715 (N_9715,N_3800,N_560);
or U9716 (N_9716,N_520,N_3109);
and U9717 (N_9717,N_590,N_4764);
nor U9718 (N_9718,N_3428,N_3419);
nor U9719 (N_9719,N_3909,N_4203);
or U9720 (N_9720,N_1179,N_1747);
nand U9721 (N_9721,N_4267,N_1540);
nor U9722 (N_9722,N_4779,N_435);
nand U9723 (N_9723,N_609,N_2463);
xor U9724 (N_9724,N_547,N_1198);
xnor U9725 (N_9725,N_1942,N_1505);
nand U9726 (N_9726,N_1226,N_650);
nand U9727 (N_9727,N_3701,N_2176);
nand U9728 (N_9728,N_1150,N_3702);
xnor U9729 (N_9729,N_4019,N_684);
xor U9730 (N_9730,N_4011,N_4708);
nor U9731 (N_9731,N_364,N_1075);
nand U9732 (N_9732,N_667,N_3946);
or U9733 (N_9733,N_2617,N_3526);
xnor U9734 (N_9734,N_1437,N_73);
nand U9735 (N_9735,N_718,N_1918);
xor U9736 (N_9736,N_3156,N_1352);
nor U9737 (N_9737,N_1487,N_2110);
and U9738 (N_9738,N_2487,N_1145);
or U9739 (N_9739,N_4211,N_80);
nor U9740 (N_9740,N_1375,N_2188);
nand U9741 (N_9741,N_4742,N_2219);
xor U9742 (N_9742,N_4423,N_1369);
or U9743 (N_9743,N_2969,N_3783);
and U9744 (N_9744,N_2725,N_1916);
xor U9745 (N_9745,N_1130,N_568);
nand U9746 (N_9746,N_1790,N_4919);
nor U9747 (N_9747,N_1171,N_2134);
and U9748 (N_9748,N_2649,N_2371);
and U9749 (N_9749,N_4186,N_1438);
or U9750 (N_9750,N_4801,N_3277);
or U9751 (N_9751,N_1187,N_386);
nor U9752 (N_9752,N_4531,N_905);
or U9753 (N_9753,N_1211,N_541);
nand U9754 (N_9754,N_4332,N_3874);
or U9755 (N_9755,N_2384,N_4252);
nor U9756 (N_9756,N_3878,N_625);
xor U9757 (N_9757,N_3090,N_3983);
xor U9758 (N_9758,N_3743,N_2933);
nor U9759 (N_9759,N_1635,N_400);
or U9760 (N_9760,N_4620,N_4672);
or U9761 (N_9761,N_1281,N_4892);
or U9762 (N_9762,N_2854,N_2469);
xnor U9763 (N_9763,N_4053,N_3526);
nor U9764 (N_9764,N_633,N_4948);
and U9765 (N_9765,N_4406,N_1772);
or U9766 (N_9766,N_3406,N_1338);
nor U9767 (N_9767,N_2520,N_1631);
nand U9768 (N_9768,N_2876,N_3085);
xor U9769 (N_9769,N_2057,N_693);
xnor U9770 (N_9770,N_4665,N_2952);
nor U9771 (N_9771,N_4475,N_3683);
xor U9772 (N_9772,N_730,N_1091);
nor U9773 (N_9773,N_4568,N_2476);
nand U9774 (N_9774,N_1637,N_2405);
nor U9775 (N_9775,N_3276,N_2396);
or U9776 (N_9776,N_4426,N_3668);
or U9777 (N_9777,N_4400,N_4279);
and U9778 (N_9778,N_4816,N_1130);
and U9779 (N_9779,N_2230,N_1721);
or U9780 (N_9780,N_1362,N_1806);
nand U9781 (N_9781,N_3285,N_3598);
or U9782 (N_9782,N_4883,N_696);
nor U9783 (N_9783,N_4940,N_4648);
or U9784 (N_9784,N_2162,N_1806);
nor U9785 (N_9785,N_2664,N_1557);
or U9786 (N_9786,N_2773,N_911);
and U9787 (N_9787,N_3295,N_2443);
or U9788 (N_9788,N_1766,N_3600);
and U9789 (N_9789,N_1268,N_2332);
xnor U9790 (N_9790,N_758,N_2931);
nor U9791 (N_9791,N_3857,N_2848);
or U9792 (N_9792,N_1864,N_45);
nand U9793 (N_9793,N_2253,N_2555);
and U9794 (N_9794,N_1849,N_2684);
and U9795 (N_9795,N_4282,N_833);
nor U9796 (N_9796,N_2791,N_1327);
nand U9797 (N_9797,N_3163,N_180);
nor U9798 (N_9798,N_69,N_4502);
and U9799 (N_9799,N_1380,N_3071);
nand U9800 (N_9800,N_1794,N_128);
and U9801 (N_9801,N_4642,N_4117);
or U9802 (N_9802,N_2766,N_3983);
or U9803 (N_9803,N_3637,N_406);
nand U9804 (N_9804,N_4847,N_3417);
or U9805 (N_9805,N_4325,N_304);
and U9806 (N_9806,N_1465,N_1611);
nor U9807 (N_9807,N_2532,N_2072);
nor U9808 (N_9808,N_3300,N_14);
nor U9809 (N_9809,N_2834,N_2134);
or U9810 (N_9810,N_4607,N_1300);
nor U9811 (N_9811,N_1586,N_2910);
and U9812 (N_9812,N_610,N_414);
and U9813 (N_9813,N_1807,N_756);
nand U9814 (N_9814,N_2606,N_3578);
or U9815 (N_9815,N_2542,N_2623);
nor U9816 (N_9816,N_29,N_1366);
nor U9817 (N_9817,N_1605,N_2748);
and U9818 (N_9818,N_188,N_4166);
nor U9819 (N_9819,N_4314,N_305);
xor U9820 (N_9820,N_2470,N_2728);
and U9821 (N_9821,N_3070,N_1197);
xor U9822 (N_9822,N_1946,N_191);
and U9823 (N_9823,N_1022,N_2530);
and U9824 (N_9824,N_3837,N_1397);
nand U9825 (N_9825,N_2908,N_4063);
xor U9826 (N_9826,N_235,N_2136);
and U9827 (N_9827,N_3148,N_4842);
nor U9828 (N_9828,N_1182,N_4497);
nor U9829 (N_9829,N_3367,N_3352);
or U9830 (N_9830,N_3215,N_4400);
nand U9831 (N_9831,N_958,N_975);
nor U9832 (N_9832,N_2824,N_4988);
nor U9833 (N_9833,N_3717,N_4215);
or U9834 (N_9834,N_3125,N_2230);
or U9835 (N_9835,N_616,N_3525);
and U9836 (N_9836,N_3993,N_3012);
or U9837 (N_9837,N_1113,N_4935);
nand U9838 (N_9838,N_2358,N_3748);
or U9839 (N_9839,N_2834,N_4952);
and U9840 (N_9840,N_3421,N_4890);
and U9841 (N_9841,N_3380,N_3029);
nand U9842 (N_9842,N_1289,N_1342);
nor U9843 (N_9843,N_1795,N_3628);
or U9844 (N_9844,N_3416,N_4772);
xor U9845 (N_9845,N_1331,N_1841);
nor U9846 (N_9846,N_4549,N_3027);
and U9847 (N_9847,N_3875,N_581);
or U9848 (N_9848,N_2887,N_1108);
nand U9849 (N_9849,N_2118,N_1002);
nand U9850 (N_9850,N_2176,N_3562);
nand U9851 (N_9851,N_1488,N_4478);
nand U9852 (N_9852,N_2769,N_3659);
nor U9853 (N_9853,N_4724,N_1827);
and U9854 (N_9854,N_2912,N_4619);
nor U9855 (N_9855,N_1008,N_4921);
xnor U9856 (N_9856,N_1146,N_898);
and U9857 (N_9857,N_4299,N_3618);
nand U9858 (N_9858,N_4563,N_3531);
and U9859 (N_9859,N_2329,N_1712);
xnor U9860 (N_9860,N_2811,N_56);
nor U9861 (N_9861,N_3986,N_2929);
or U9862 (N_9862,N_296,N_2153);
xnor U9863 (N_9863,N_4916,N_1313);
xnor U9864 (N_9864,N_4902,N_4648);
nor U9865 (N_9865,N_1513,N_4309);
and U9866 (N_9866,N_2147,N_4438);
xnor U9867 (N_9867,N_1598,N_573);
nand U9868 (N_9868,N_4267,N_3081);
nor U9869 (N_9869,N_195,N_2521);
nand U9870 (N_9870,N_2488,N_502);
xor U9871 (N_9871,N_3153,N_323);
nand U9872 (N_9872,N_538,N_354);
nand U9873 (N_9873,N_2607,N_675);
and U9874 (N_9874,N_537,N_1241);
nor U9875 (N_9875,N_3700,N_2981);
xnor U9876 (N_9876,N_4933,N_2177);
or U9877 (N_9877,N_1397,N_2469);
and U9878 (N_9878,N_2313,N_4494);
nand U9879 (N_9879,N_2072,N_4429);
xnor U9880 (N_9880,N_157,N_274);
or U9881 (N_9881,N_3136,N_2452);
nor U9882 (N_9882,N_2211,N_1148);
and U9883 (N_9883,N_2331,N_3410);
xnor U9884 (N_9884,N_3792,N_3073);
nand U9885 (N_9885,N_1928,N_1228);
nor U9886 (N_9886,N_2272,N_3038);
or U9887 (N_9887,N_1954,N_3568);
xor U9888 (N_9888,N_1847,N_1817);
or U9889 (N_9889,N_1526,N_2021);
xor U9890 (N_9890,N_3616,N_2365);
nand U9891 (N_9891,N_702,N_2250);
nor U9892 (N_9892,N_2002,N_167);
and U9893 (N_9893,N_2498,N_1865);
nand U9894 (N_9894,N_1307,N_2600);
nor U9895 (N_9895,N_4271,N_1203);
and U9896 (N_9896,N_2442,N_2049);
nand U9897 (N_9897,N_3650,N_2816);
or U9898 (N_9898,N_3244,N_1125);
xnor U9899 (N_9899,N_3698,N_2181);
and U9900 (N_9900,N_3361,N_1504);
or U9901 (N_9901,N_1104,N_3582);
xnor U9902 (N_9902,N_4141,N_81);
nor U9903 (N_9903,N_1892,N_3475);
nor U9904 (N_9904,N_424,N_1146);
nand U9905 (N_9905,N_1436,N_78);
nand U9906 (N_9906,N_1567,N_4711);
xnor U9907 (N_9907,N_1610,N_4631);
and U9908 (N_9908,N_4316,N_2810);
nor U9909 (N_9909,N_386,N_3866);
nor U9910 (N_9910,N_2325,N_2757);
xnor U9911 (N_9911,N_31,N_2854);
nand U9912 (N_9912,N_3624,N_473);
or U9913 (N_9913,N_3462,N_1557);
or U9914 (N_9914,N_2038,N_1651);
nand U9915 (N_9915,N_2789,N_4374);
and U9916 (N_9916,N_3933,N_4191);
nand U9917 (N_9917,N_865,N_652);
xor U9918 (N_9918,N_2732,N_126);
nor U9919 (N_9919,N_599,N_3544);
xnor U9920 (N_9920,N_1755,N_2831);
nor U9921 (N_9921,N_2147,N_4571);
and U9922 (N_9922,N_4041,N_649);
and U9923 (N_9923,N_205,N_778);
or U9924 (N_9924,N_2952,N_2241);
and U9925 (N_9925,N_1132,N_2683);
nand U9926 (N_9926,N_4802,N_1321);
xnor U9927 (N_9927,N_2715,N_1835);
nand U9928 (N_9928,N_3751,N_2308);
nor U9929 (N_9929,N_2112,N_1691);
nand U9930 (N_9930,N_4387,N_106);
or U9931 (N_9931,N_3773,N_4034);
nand U9932 (N_9932,N_4644,N_2933);
or U9933 (N_9933,N_1114,N_4515);
nor U9934 (N_9934,N_3923,N_2450);
or U9935 (N_9935,N_1791,N_3426);
or U9936 (N_9936,N_4433,N_647);
xnor U9937 (N_9937,N_4125,N_703);
xnor U9938 (N_9938,N_3339,N_587);
and U9939 (N_9939,N_2507,N_2571);
nor U9940 (N_9940,N_3420,N_747);
or U9941 (N_9941,N_2037,N_3625);
or U9942 (N_9942,N_1398,N_791);
nor U9943 (N_9943,N_507,N_1264);
and U9944 (N_9944,N_1110,N_790);
nor U9945 (N_9945,N_4475,N_2525);
or U9946 (N_9946,N_3898,N_1213);
nand U9947 (N_9947,N_531,N_3814);
nor U9948 (N_9948,N_344,N_3182);
nor U9949 (N_9949,N_2683,N_2781);
and U9950 (N_9950,N_4065,N_3002);
and U9951 (N_9951,N_3421,N_853);
nand U9952 (N_9952,N_4237,N_1775);
xor U9953 (N_9953,N_4223,N_743);
xor U9954 (N_9954,N_1334,N_4121);
and U9955 (N_9955,N_3728,N_4983);
nor U9956 (N_9956,N_1764,N_800);
and U9957 (N_9957,N_1438,N_1947);
or U9958 (N_9958,N_3888,N_1785);
nor U9959 (N_9959,N_4258,N_1693);
and U9960 (N_9960,N_416,N_2033);
nand U9961 (N_9961,N_2674,N_1267);
nor U9962 (N_9962,N_2690,N_2806);
or U9963 (N_9963,N_3566,N_3853);
and U9964 (N_9964,N_4002,N_4539);
nand U9965 (N_9965,N_4823,N_1341);
nor U9966 (N_9966,N_292,N_17);
or U9967 (N_9967,N_1779,N_2676);
nand U9968 (N_9968,N_2007,N_2148);
and U9969 (N_9969,N_29,N_3601);
xnor U9970 (N_9970,N_3043,N_3069);
nand U9971 (N_9971,N_4204,N_4489);
nor U9972 (N_9972,N_4805,N_206);
nor U9973 (N_9973,N_1627,N_382);
and U9974 (N_9974,N_636,N_1755);
nand U9975 (N_9975,N_3265,N_2741);
xor U9976 (N_9976,N_1038,N_1882);
xnor U9977 (N_9977,N_842,N_4728);
and U9978 (N_9978,N_3777,N_4891);
and U9979 (N_9979,N_1000,N_4830);
nor U9980 (N_9980,N_2361,N_4176);
nand U9981 (N_9981,N_2667,N_4052);
and U9982 (N_9982,N_1076,N_2007);
nand U9983 (N_9983,N_1659,N_840);
or U9984 (N_9984,N_1778,N_2742);
xor U9985 (N_9985,N_3665,N_2564);
nand U9986 (N_9986,N_2687,N_3357);
or U9987 (N_9987,N_3027,N_3212);
xor U9988 (N_9988,N_4263,N_2061);
nor U9989 (N_9989,N_2999,N_516);
and U9990 (N_9990,N_1540,N_2061);
and U9991 (N_9991,N_1887,N_3931);
and U9992 (N_9992,N_842,N_3200);
xor U9993 (N_9993,N_1450,N_2778);
and U9994 (N_9994,N_460,N_4037);
xor U9995 (N_9995,N_2218,N_1930);
nand U9996 (N_9996,N_4620,N_525);
and U9997 (N_9997,N_902,N_109);
nor U9998 (N_9998,N_2504,N_2239);
nand U9999 (N_9999,N_3894,N_3714);
nor U10000 (N_10000,N_7962,N_7961);
and U10001 (N_10001,N_6993,N_9892);
or U10002 (N_10002,N_6429,N_8475);
nand U10003 (N_10003,N_8413,N_5328);
nor U10004 (N_10004,N_5097,N_8619);
and U10005 (N_10005,N_9019,N_5353);
xor U10006 (N_10006,N_8762,N_5699);
nand U10007 (N_10007,N_7578,N_5336);
nor U10008 (N_10008,N_8134,N_7787);
xnor U10009 (N_10009,N_7428,N_5498);
nand U10010 (N_10010,N_9866,N_5108);
nand U10011 (N_10011,N_7856,N_7848);
nor U10012 (N_10012,N_9235,N_6891);
xor U10013 (N_10013,N_8321,N_9407);
or U10014 (N_10014,N_9133,N_7380);
or U10015 (N_10015,N_5305,N_6110);
nor U10016 (N_10016,N_8656,N_7821);
nand U10017 (N_10017,N_6123,N_6660);
and U10018 (N_10018,N_6622,N_8182);
nand U10019 (N_10019,N_8342,N_9279);
nand U10020 (N_10020,N_5303,N_7016);
and U10021 (N_10021,N_5481,N_9004);
or U10022 (N_10022,N_9801,N_8665);
and U10023 (N_10023,N_7599,N_6909);
nor U10024 (N_10024,N_9995,N_8967);
xnor U10025 (N_10025,N_9575,N_5804);
nand U10026 (N_10026,N_8313,N_5258);
and U10027 (N_10027,N_9784,N_6015);
and U10028 (N_10028,N_7191,N_6498);
nand U10029 (N_10029,N_9250,N_9337);
nor U10030 (N_10030,N_7756,N_8568);
and U10031 (N_10031,N_7203,N_5443);
xor U10032 (N_10032,N_5862,N_5206);
or U10033 (N_10033,N_9294,N_8207);
and U10034 (N_10034,N_8708,N_8145);
nand U10035 (N_10035,N_8434,N_8021);
nand U10036 (N_10036,N_7989,N_8565);
or U10037 (N_10037,N_7001,N_6302);
xnor U10038 (N_10038,N_5176,N_6674);
xnor U10039 (N_10039,N_6164,N_7754);
and U10040 (N_10040,N_7995,N_8788);
nor U10041 (N_10041,N_5073,N_6528);
nor U10042 (N_10042,N_5456,N_8871);
xnor U10043 (N_10043,N_8789,N_5789);
or U10044 (N_10044,N_8718,N_9262);
and U10045 (N_10045,N_7321,N_6075);
xnor U10046 (N_10046,N_5806,N_9792);
and U10047 (N_10047,N_9411,N_7815);
nand U10048 (N_10048,N_8080,N_9067);
nand U10049 (N_10049,N_9105,N_7782);
and U10050 (N_10050,N_5900,N_6945);
nor U10051 (N_10051,N_5376,N_7116);
or U10052 (N_10052,N_6409,N_8140);
nor U10053 (N_10053,N_8070,N_6049);
nor U10054 (N_10054,N_5741,N_9198);
xor U10055 (N_10055,N_7274,N_7642);
xnor U10056 (N_10056,N_8770,N_8461);
nor U10057 (N_10057,N_7575,N_8933);
and U10058 (N_10058,N_7547,N_8064);
or U10059 (N_10059,N_6006,N_9335);
or U10060 (N_10060,N_7901,N_8132);
nand U10061 (N_10061,N_5865,N_9480);
xor U10062 (N_10062,N_9841,N_9179);
nand U10063 (N_10063,N_9523,N_9965);
nand U10064 (N_10064,N_5510,N_7381);
xnor U10065 (N_10065,N_9246,N_9372);
and U10066 (N_10066,N_7177,N_6431);
nor U10067 (N_10067,N_7407,N_6316);
and U10068 (N_10068,N_8219,N_6928);
or U10069 (N_10069,N_7216,N_6976);
nor U10070 (N_10070,N_5253,N_6505);
or U10071 (N_10071,N_6981,N_5468);
and U10072 (N_10072,N_9464,N_6056);
and U10073 (N_10073,N_9991,N_5933);
nor U10074 (N_10074,N_9943,N_6307);
nand U10075 (N_10075,N_9795,N_7669);
nor U10076 (N_10076,N_9000,N_9805);
or U10077 (N_10077,N_7509,N_7532);
xor U10078 (N_10078,N_7679,N_6761);
and U10079 (N_10079,N_7730,N_6688);
and U10080 (N_10080,N_6369,N_7793);
or U10081 (N_10081,N_9569,N_5674);
or U10082 (N_10082,N_8947,N_8533);
and U10083 (N_10083,N_7517,N_5539);
nor U10084 (N_10084,N_5534,N_7391);
xnor U10085 (N_10085,N_8977,N_8868);
and U10086 (N_10086,N_6356,N_5999);
and U10087 (N_10087,N_6742,N_9050);
xnor U10088 (N_10088,N_8618,N_8894);
and U10089 (N_10089,N_6522,N_5544);
nand U10090 (N_10090,N_5803,N_7263);
nor U10091 (N_10091,N_7968,N_8778);
nand U10092 (N_10092,N_7617,N_8734);
and U10093 (N_10093,N_7333,N_6400);
or U10094 (N_10094,N_7984,N_7067);
nor U10095 (N_10095,N_6567,N_9616);
nor U10096 (N_10096,N_7893,N_9859);
xnor U10097 (N_10097,N_9488,N_6105);
xnor U10098 (N_10098,N_7163,N_5655);
nor U10099 (N_10099,N_6951,N_8333);
xnor U10100 (N_10100,N_5871,N_6546);
nand U10101 (N_10101,N_7631,N_7506);
xnor U10102 (N_10102,N_8936,N_8640);
and U10103 (N_10103,N_9089,N_6131);
nand U10104 (N_10104,N_7921,N_6325);
or U10105 (N_10105,N_7709,N_9394);
nand U10106 (N_10106,N_6971,N_6843);
or U10107 (N_10107,N_9092,N_7991);
and U10108 (N_10108,N_9743,N_7275);
nand U10109 (N_10109,N_7105,N_9315);
nor U10110 (N_10110,N_5605,N_9899);
or U10111 (N_10111,N_7621,N_5678);
and U10112 (N_10112,N_9257,N_8932);
nor U10113 (N_10113,N_8638,N_8381);
or U10114 (N_10114,N_9111,N_5065);
nor U10115 (N_10115,N_6308,N_6958);
and U10116 (N_10116,N_9256,N_7917);
or U10117 (N_10117,N_6669,N_6575);
or U10118 (N_10118,N_5561,N_8769);
nand U10119 (N_10119,N_5288,N_5799);
nand U10120 (N_10120,N_7450,N_5310);
xnor U10121 (N_10121,N_8004,N_9648);
nand U10122 (N_10122,N_7319,N_7474);
nor U10123 (N_10123,N_7375,N_8858);
and U10124 (N_10124,N_5289,N_6675);
xor U10125 (N_10125,N_6760,N_7472);
nor U10126 (N_10126,N_8751,N_8037);
and U10127 (N_10127,N_9340,N_9309);
xnor U10128 (N_10128,N_7774,N_5026);
nand U10129 (N_10129,N_9532,N_7788);
nor U10130 (N_10130,N_7083,N_5362);
and U10131 (N_10131,N_8469,N_8314);
or U10132 (N_10132,N_8493,N_7336);
or U10133 (N_10133,N_9373,N_5094);
xor U10134 (N_10134,N_9941,N_6747);
nor U10135 (N_10135,N_9145,N_5488);
and U10136 (N_10136,N_5926,N_8567);
or U10137 (N_10137,N_7370,N_7993);
xor U10138 (N_10138,N_6552,N_8485);
or U10139 (N_10139,N_8500,N_6019);
nand U10140 (N_10140,N_7429,N_7181);
nor U10141 (N_10141,N_7422,N_9530);
nor U10142 (N_10142,N_9644,N_9116);
nor U10143 (N_10143,N_7860,N_5323);
xor U10144 (N_10144,N_7889,N_8864);
nand U10145 (N_10145,N_8186,N_5416);
xnor U10146 (N_10146,N_7361,N_9762);
nor U10147 (N_10147,N_6849,N_6905);
nor U10148 (N_10148,N_9932,N_9101);
and U10149 (N_10149,N_7530,N_6236);
or U10150 (N_10150,N_5232,N_7954);
nand U10151 (N_10151,N_7071,N_9420);
and U10152 (N_10152,N_8201,N_7277);
and U10153 (N_10153,N_5837,N_6310);
nor U10154 (N_10154,N_5686,N_6708);
and U10155 (N_10155,N_5922,N_8874);
nand U10156 (N_10156,N_5939,N_9117);
or U10157 (N_10157,N_9700,N_6732);
or U10158 (N_10158,N_6472,N_6919);
xnor U10159 (N_10159,N_9724,N_6658);
xor U10160 (N_10160,N_6806,N_9826);
nand U10161 (N_10161,N_5181,N_8232);
xnor U10162 (N_10162,N_7158,N_8099);
and U10163 (N_10163,N_9576,N_5364);
or U10164 (N_10164,N_6453,N_5371);
xnor U10165 (N_10165,N_9497,N_6288);
nand U10166 (N_10166,N_5370,N_6884);
nand U10167 (N_10167,N_7762,N_6815);
or U10168 (N_10168,N_5742,N_8197);
xor U10169 (N_10169,N_8904,N_7919);
or U10170 (N_10170,N_9357,N_9266);
xor U10171 (N_10171,N_9579,N_6997);
or U10172 (N_10172,N_6375,N_7088);
and U10173 (N_10173,N_8729,N_5902);
nand U10174 (N_10174,N_6046,N_8442);
or U10175 (N_10175,N_7876,N_6141);
and U10176 (N_10176,N_6259,N_8347);
or U10177 (N_10177,N_7715,N_9426);
or U10178 (N_10178,N_9352,N_5893);
nor U10179 (N_10179,N_8206,N_8616);
xnor U10180 (N_10180,N_7455,N_9916);
nand U10181 (N_10181,N_8457,N_5651);
nand U10182 (N_10182,N_8644,N_9330);
and U10183 (N_10183,N_6260,N_5746);
or U10184 (N_10184,N_5142,N_8800);
and U10185 (N_10185,N_7289,N_5598);
nor U10186 (N_10186,N_9147,N_8570);
and U10187 (N_10187,N_9056,N_6706);
nand U10188 (N_10188,N_8170,N_5571);
xnor U10189 (N_10189,N_5188,N_5719);
nor U10190 (N_10190,N_9415,N_7900);
or U10191 (N_10191,N_9127,N_5169);
nand U10192 (N_10192,N_7563,N_7287);
nand U10193 (N_10193,N_8428,N_5850);
nand U10194 (N_10194,N_9209,N_5672);
or U10195 (N_10195,N_7448,N_5795);
xnor U10196 (N_10196,N_5543,N_5815);
and U10197 (N_10197,N_9510,N_7271);
xnor U10198 (N_10198,N_8694,N_7392);
xor U10199 (N_10199,N_9362,N_6309);
and U10200 (N_10200,N_9201,N_6728);
nand U10201 (N_10201,N_8759,N_9516);
nor U10202 (N_10202,N_7923,N_6603);
nand U10203 (N_10203,N_8861,N_9012);
xor U10204 (N_10204,N_6966,N_7233);
nand U10205 (N_10205,N_5961,N_5016);
nor U10206 (N_10206,N_5966,N_6427);
nor U10207 (N_10207,N_9143,N_6959);
nand U10208 (N_10208,N_8209,N_6073);
nand U10209 (N_10209,N_8453,N_9285);
nor U10210 (N_10210,N_8459,N_8642);
or U10211 (N_10211,N_8615,N_6115);
nand U10212 (N_10212,N_5620,N_8014);
nor U10213 (N_10213,N_5852,N_7928);
nand U10214 (N_10214,N_6112,N_5831);
and U10215 (N_10215,N_6490,N_8719);
nor U10216 (N_10216,N_8174,N_9293);
or U10217 (N_10217,N_7916,N_7064);
and U10218 (N_10218,N_8429,N_7930);
xor U10219 (N_10219,N_8312,N_8462);
and U10220 (N_10220,N_5722,N_7784);
xor U10221 (N_10221,N_6512,N_9643);
nor U10222 (N_10222,N_5735,N_9625);
xor U10223 (N_10223,N_8395,N_6821);
xor U10224 (N_10224,N_7082,N_9742);
nor U10225 (N_10225,N_5974,N_5550);
nand U10226 (N_10226,N_9486,N_9825);
xor U10227 (N_10227,N_9430,N_6205);
nand U10228 (N_10228,N_7896,N_9592);
or U10229 (N_10229,N_6101,N_5492);
nor U10230 (N_10230,N_9313,N_6768);
or U10231 (N_10231,N_5942,N_7162);
nand U10232 (N_10232,N_8282,N_8608);
nand U10233 (N_10233,N_9987,N_5327);
or U10234 (N_10234,N_8245,N_8715);
xnor U10235 (N_10235,N_8259,N_6191);
nor U10236 (N_10236,N_8943,N_9493);
xnor U10237 (N_10237,N_8702,N_6229);
nor U10238 (N_10238,N_6014,N_9642);
or U10239 (N_10239,N_9156,N_7008);
and U10240 (N_10240,N_8220,N_9653);
and U10241 (N_10241,N_5827,N_6072);
or U10242 (N_10242,N_7047,N_7851);
nand U10243 (N_10243,N_9986,N_6988);
and U10244 (N_10244,N_5070,N_9698);
nand U10245 (N_10245,N_9354,N_8880);
nand U10246 (N_10246,N_5527,N_7101);
and U10247 (N_10247,N_7383,N_6804);
xnor U10248 (N_10248,N_6537,N_5405);
and U10249 (N_10249,N_6393,N_9386);
xor U10250 (N_10250,N_6084,N_6598);
nand U10251 (N_10251,N_7394,N_6574);
and U10252 (N_10252,N_6315,N_6169);
nand U10253 (N_10253,N_6224,N_5236);
nor U10254 (N_10254,N_6331,N_5104);
nand U10255 (N_10255,N_6285,N_6639);
nor U10256 (N_10256,N_9591,N_8523);
nor U10257 (N_10257,N_9495,N_6947);
xor U10258 (N_10258,N_5355,N_8606);
nor U10259 (N_10259,N_6280,N_9290);
and U10260 (N_10260,N_7938,N_7309);
xnor U10261 (N_10261,N_8155,N_8508);
xnor U10262 (N_10262,N_6594,N_7801);
nor U10263 (N_10263,N_7464,N_8978);
or U10264 (N_10264,N_7701,N_5513);
or U10265 (N_10265,N_6257,N_9728);
xor U10266 (N_10266,N_7926,N_8414);
nand U10267 (N_10267,N_5625,N_8921);
or U10268 (N_10268,N_5201,N_5863);
nand U10269 (N_10269,N_5136,N_6155);
or U10270 (N_10270,N_8077,N_5196);
xnor U10271 (N_10271,N_5830,N_6187);
or U10272 (N_10272,N_9349,N_9476);
xnor U10273 (N_10273,N_5629,N_8798);
or U10274 (N_10274,N_6354,N_7789);
xor U10275 (N_10275,N_9424,N_8412);
and U10276 (N_10276,N_8354,N_5398);
and U10277 (N_10277,N_6055,N_8062);
xor U10278 (N_10278,N_5957,N_5989);
and U10279 (N_10279,N_6385,N_7208);
nand U10280 (N_10280,N_9170,N_8173);
or U10281 (N_10281,N_5182,N_9560);
xnor U10282 (N_10282,N_8760,N_9061);
xnor U10283 (N_10283,N_6436,N_9039);
nand U10284 (N_10284,N_8464,N_5419);
or U10285 (N_10285,N_7122,N_7721);
nor U10286 (N_10286,N_8555,N_7417);
or U10287 (N_10287,N_6077,N_5093);
nand U10288 (N_10288,N_8722,N_6978);
nand U10289 (N_10289,N_8227,N_6138);
or U10290 (N_10290,N_7221,N_5020);
or U10291 (N_10291,N_8228,N_8538);
or U10292 (N_10292,N_8497,N_8558);
and U10293 (N_10293,N_5587,N_9199);
and U10294 (N_10294,N_9097,N_6339);
nor U10295 (N_10295,N_7755,N_9259);
xor U10296 (N_10296,N_9405,N_7904);
xor U10297 (N_10297,N_9777,N_8211);
nor U10298 (N_10298,N_6679,N_5062);
and U10299 (N_10299,N_8052,N_6198);
or U10300 (N_10300,N_9194,N_7684);
nor U10301 (N_10301,N_5436,N_9909);
nand U10302 (N_10302,N_5151,N_7297);
xnor U10303 (N_10303,N_9243,N_6344);
nand U10304 (N_10304,N_6135,N_8042);
nor U10305 (N_10305,N_7457,N_9580);
nor U10306 (N_10306,N_6620,N_7898);
or U10307 (N_10307,N_6185,N_8194);
nand U10308 (N_10308,N_9928,N_7199);
and U10309 (N_10309,N_5532,N_9696);
or U10310 (N_10310,N_8982,N_7590);
and U10311 (N_10311,N_8458,N_7232);
or U10312 (N_10312,N_8624,N_5463);
nand U10313 (N_10313,N_7413,N_7073);
and U10314 (N_10314,N_8513,N_9766);
xor U10315 (N_10315,N_8388,N_9672);
nor U10316 (N_10316,N_6696,N_5347);
or U10317 (N_10317,N_6838,N_7559);
nor U10318 (N_10318,N_7143,N_5111);
or U10319 (N_10319,N_7759,N_9802);
nand U10320 (N_10320,N_9325,N_5015);
nor U10321 (N_10321,N_9190,N_9388);
or U10322 (N_10322,N_9203,N_9462);
or U10323 (N_10323,N_7596,N_5283);
xor U10324 (N_10324,N_7491,N_7920);
nand U10325 (N_10325,N_6443,N_5124);
and U10326 (N_10326,N_6178,N_9297);
nor U10327 (N_10327,N_8940,N_6842);
and U10328 (N_10328,N_8526,N_6426);
nor U10329 (N_10329,N_5464,N_8152);
nand U10330 (N_10330,N_6465,N_7052);
nor U10331 (N_10331,N_5010,N_7732);
nand U10332 (N_10332,N_7724,N_8691);
nand U10333 (N_10333,N_5393,N_7259);
nand U10334 (N_10334,N_6078,N_8217);
or U10335 (N_10335,N_5412,N_5382);
xor U10336 (N_10336,N_5135,N_8536);
and U10337 (N_10337,N_6320,N_7859);
and U10338 (N_10338,N_5307,N_8931);
or U10339 (N_10339,N_8075,N_8974);
and U10340 (N_10340,N_9036,N_7985);
nand U10341 (N_10341,N_6555,N_5220);
nand U10342 (N_10342,N_8191,N_6955);
or U10343 (N_10343,N_9609,N_9224);
or U10344 (N_10344,N_6167,N_5003);
or U10345 (N_10345,N_5851,N_5754);
or U10346 (N_10346,N_8454,N_9554);
nand U10347 (N_10347,N_6441,N_6491);
nand U10348 (N_10348,N_7529,N_8484);
xnor U10349 (N_10349,N_8824,N_9163);
nor U10350 (N_10350,N_8609,N_8580);
or U10351 (N_10351,N_5660,N_7226);
xor U10352 (N_10352,N_9024,N_7145);
xor U10353 (N_10353,N_6968,N_8143);
xnor U10354 (N_10354,N_6486,N_9206);
nand U10355 (N_10355,N_5263,N_5000);
nand U10356 (N_10356,N_6462,N_7691);
xnor U10357 (N_10357,N_5624,N_7890);
nand U10358 (N_10358,N_8131,N_5679);
nand U10359 (N_10359,N_8621,N_8437);
nor U10360 (N_10360,N_8095,N_7946);
nor U10361 (N_10361,N_9834,N_7771);
and U10362 (N_10362,N_6290,N_6351);
nor U10363 (N_10363,N_9214,N_6301);
nor U10364 (N_10364,N_6274,N_8534);
nor U10365 (N_10365,N_9369,N_8287);
xnor U10366 (N_10366,N_9436,N_9824);
and U10367 (N_10367,N_6292,N_6831);
xor U10368 (N_10368,N_9940,N_6044);
and U10369 (N_10369,N_9099,N_7172);
or U10370 (N_10370,N_8058,N_7262);
nor U10371 (N_10371,N_9539,N_9504);
xnor U10372 (N_10372,N_5623,N_5462);
nand U10373 (N_10373,N_5157,N_8877);
nor U10374 (N_10374,N_7875,N_9417);
or U10375 (N_10375,N_8742,N_7054);
and U10376 (N_10376,N_9134,N_6425);
or U10377 (N_10377,N_9468,N_7501);
or U10378 (N_10378,N_7671,N_6935);
nor U10379 (N_10379,N_7841,N_9954);
and U10380 (N_10380,N_7245,N_7924);
and U10381 (N_10381,N_6727,N_7194);
nor U10382 (N_10382,N_8910,N_8264);
nand U10383 (N_10383,N_9073,N_6926);
and U10384 (N_10384,N_8024,N_5163);
and U10385 (N_10385,N_7310,N_7544);
or U10386 (N_10386,N_9267,N_8808);
nand U10387 (N_10387,N_9114,N_7884);
or U10388 (N_10388,N_6041,N_9741);
or U10389 (N_10389,N_7397,N_7553);
and U10390 (N_10390,N_7533,N_9007);
or U10391 (N_10391,N_7009,N_5427);
or U10392 (N_10392,N_7063,N_9612);
nor U10393 (N_10393,N_8183,N_5739);
xnor U10394 (N_10394,N_9229,N_8733);
and U10395 (N_10395,N_5970,N_8404);
xnor U10396 (N_10396,N_9184,N_8905);
nand U10397 (N_10397,N_8806,N_5100);
xor U10398 (N_10398,N_9138,N_5024);
nand U10399 (N_10399,N_5279,N_7167);
or U10400 (N_10400,N_7408,N_8588);
nor U10401 (N_10401,N_7645,N_9861);
nand U10402 (N_10402,N_6237,N_9541);
and U10403 (N_10403,N_6918,N_7185);
and U10404 (N_10404,N_8482,N_5580);
and U10405 (N_10405,N_9720,N_7925);
and U10406 (N_10406,N_6360,N_9773);
nand U10407 (N_10407,N_6153,N_8471);
or U10408 (N_10408,N_6504,N_6298);
nor U10409 (N_10409,N_6312,N_5511);
xor U10410 (N_10410,N_8337,N_6529);
or U10411 (N_10411,N_8892,N_6002);
nor U10412 (N_10412,N_6830,N_8171);
and U10413 (N_10413,N_9967,N_8930);
nand U10414 (N_10414,N_8285,N_6826);
and U10415 (N_10415,N_9974,N_7495);
xnor U10416 (N_10416,N_5442,N_7581);
nor U10417 (N_10417,N_6850,N_8654);
and U10418 (N_10418,N_7393,N_5084);
xor U10419 (N_10419,N_9761,N_5165);
and U10420 (N_10420,N_5213,N_8048);
or U10421 (N_10421,N_6384,N_6651);
xor U10422 (N_10422,N_5964,N_6295);
and U10423 (N_10423,N_7362,N_6720);
and U10424 (N_10424,N_6705,N_5642);
nor U10425 (N_10425,N_8540,N_7668);
nor U10426 (N_10426,N_5428,N_8195);
nor U10427 (N_10427,N_6104,N_7024);
nand U10428 (N_10428,N_9975,N_8231);
xor U10429 (N_10429,N_6765,N_9626);
nor U10430 (N_10430,N_7060,N_7825);
and U10431 (N_10431,N_5568,N_8448);
and U10432 (N_10432,N_5928,N_5844);
and U10433 (N_10433,N_7700,N_9220);
and U10434 (N_10434,N_7286,N_5119);
nand U10435 (N_10435,N_8281,N_8230);
xor U10436 (N_10436,N_6053,N_9453);
and U10437 (N_10437,N_5589,N_8000);
nor U10438 (N_10438,N_6543,N_6799);
or U10439 (N_10439,N_9982,N_7378);
nand U10440 (N_10440,N_7696,N_5794);
nor U10441 (N_10441,N_8463,N_5372);
nand U10442 (N_10442,N_9230,N_5557);
nor U10443 (N_10443,N_8963,N_7029);
nand U10444 (N_10444,N_9065,N_9587);
or U10445 (N_10445,N_8586,N_6210);
nor U10446 (N_10446,N_8271,N_7775);
nor U10447 (N_10447,N_7023,N_6433);
nand U10448 (N_10448,N_7736,N_8834);
xor U10449 (N_10449,N_6481,N_8401);
xnor U10450 (N_10450,N_9113,N_9136);
or U10451 (N_10451,N_6036,N_8820);
xor U10452 (N_10452,N_6940,N_9359);
xor U10453 (N_10453,N_7104,N_6957);
nor U10454 (N_10454,N_5541,N_5234);
or U10455 (N_10455,N_9561,N_7477);
and U10456 (N_10456,N_7750,N_6614);
xnor U10457 (N_10457,N_7880,N_8325);
nand U10458 (N_10458,N_5566,N_5089);
xnor U10459 (N_10459,N_6816,N_9454);
and U10460 (N_10460,N_6701,N_5599);
or U10461 (N_10461,N_6922,N_5096);
and U10462 (N_10462,N_8289,N_9272);
nand U10463 (N_10463,N_8233,N_5845);
xor U10464 (N_10464,N_6069,N_5431);
nand U10465 (N_10465,N_9827,N_5095);
and U10466 (N_10466,N_7997,N_5267);
nand U10467 (N_10467,N_7182,N_8643);
nand U10468 (N_10468,N_5432,N_6083);
nor U10469 (N_10469,N_7792,N_8721);
nand U10470 (N_10470,N_5349,N_7228);
or U10471 (N_10471,N_5663,N_7752);
xnor U10472 (N_10472,N_6663,N_9716);
or U10473 (N_10473,N_9669,N_7249);
nor U10474 (N_10474,N_9810,N_6609);
and U10475 (N_10475,N_7204,N_8677);
or U10476 (N_10476,N_7212,N_7749);
nand U10477 (N_10477,N_9284,N_5407);
nor U10478 (N_10478,N_7514,N_9788);
nand U10479 (N_10479,N_8678,N_5992);
xor U10480 (N_10480,N_6540,N_6779);
or U10481 (N_10481,N_9973,N_5879);
nor U10482 (N_10482,N_5633,N_8854);
nand U10483 (N_10483,N_7630,N_8012);
xnor U10484 (N_10484,N_7291,N_7566);
and U10485 (N_10485,N_7567,N_6618);
or U10486 (N_10486,N_7718,N_6203);
or U10487 (N_10487,N_7883,N_7521);
and U10488 (N_10488,N_9183,N_6763);
or U10489 (N_10489,N_8329,N_5727);
or U10490 (N_10490,N_6973,N_9258);
or U10491 (N_10491,N_7099,N_5471);
nand U10492 (N_10492,N_7433,N_7481);
nor U10493 (N_10493,N_7377,N_5667);
nand U10494 (N_10494,N_5348,N_9508);
xor U10495 (N_10495,N_9251,N_5235);
nand U10496 (N_10496,N_7373,N_7694);
or U10497 (N_10497,N_5164,N_9025);
nand U10498 (N_10498,N_7999,N_6190);
nand U10499 (N_10499,N_7894,N_6704);
xnor U10500 (N_10500,N_8547,N_8782);
xnor U10501 (N_10501,N_6173,N_9200);
nand U10502 (N_10502,N_7225,N_5507);
and U10503 (N_10503,N_8439,N_7356);
nor U10504 (N_10504,N_8650,N_8791);
and U10505 (N_10505,N_5277,N_9692);
nand U10506 (N_10506,N_8291,N_8026);
nor U10507 (N_10507,N_6451,N_9160);
or U10508 (N_10508,N_5848,N_9557);
xor U10509 (N_10509,N_9875,N_6589);
or U10510 (N_10510,N_9389,N_7251);
and U10511 (N_10511,N_7197,N_8441);
xnor U10512 (N_10512,N_9755,N_6738);
and U10513 (N_10513,N_6681,N_6382);
or U10514 (N_10514,N_6042,N_6476);
or U10515 (N_10515,N_8392,N_7807);
nor U10516 (N_10516,N_7400,N_8361);
nor U10517 (N_10517,N_8779,N_9949);
nand U10518 (N_10518,N_6568,N_9747);
nand U10519 (N_10519,N_5202,N_5088);
and U10520 (N_10520,N_9639,N_9942);
xor U10521 (N_10521,N_5317,N_5137);
or U10522 (N_10522,N_7156,N_6936);
and U10523 (N_10523,N_7470,N_9952);
xnor U10524 (N_10524,N_7790,N_8255);
nor U10525 (N_10525,N_5159,N_5351);
nor U10526 (N_10526,N_7745,N_8300);
or U10527 (N_10527,N_7032,N_7248);
and U10528 (N_10528,N_7186,N_8658);
nor U10529 (N_10529,N_5564,N_7065);
or U10530 (N_10530,N_7267,N_8051);
and U10531 (N_10531,N_6114,N_5354);
nand U10532 (N_10532,N_5047,N_9208);
nor U10533 (N_10533,N_5854,N_6599);
or U10534 (N_10534,N_5002,N_8763);
nand U10535 (N_10535,N_5334,N_8850);
nor U10536 (N_10536,N_5391,N_5840);
nor U10537 (N_10537,N_5702,N_6374);
and U10538 (N_10538,N_6080,N_5724);
or U10539 (N_10539,N_9041,N_8917);
or U10540 (N_10540,N_5453,N_5603);
nor U10541 (N_10541,N_7826,N_8541);
xor U10542 (N_10542,N_6347,N_6729);
nand U10543 (N_10543,N_6251,N_8689);
xor U10544 (N_10544,N_7682,N_8277);
xnor U10545 (N_10545,N_5757,N_5683);
and U10546 (N_10546,N_9384,N_5826);
and U10547 (N_10547,N_8754,N_9711);
and U10548 (N_10548,N_5858,N_8637);
nor U10549 (N_10549,N_8670,N_7086);
or U10550 (N_10550,N_5374,N_8929);
nand U10551 (N_10551,N_7828,N_8593);
nor U10552 (N_10552,N_5864,N_8979);
and U10553 (N_10553,N_5256,N_6264);
nand U10554 (N_10554,N_7504,N_9819);
xor U10555 (N_10555,N_6697,N_8888);
or U10556 (N_10556,N_9106,N_5740);
nand U10557 (N_10557,N_7030,N_9549);
xnor U10558 (N_10558,N_5914,N_6854);
nor U10559 (N_10559,N_9475,N_6896);
or U10560 (N_10560,N_7974,N_8362);
or U10561 (N_10561,N_9181,N_6457);
nor U10562 (N_10562,N_7839,N_7576);
and U10563 (N_10563,N_5041,N_9289);
nand U10564 (N_10564,N_9398,N_6814);
nand U10565 (N_10565,N_9647,N_9759);
or U10566 (N_10566,N_9144,N_5594);
nor U10567 (N_10567,N_6977,N_7562);
or U10568 (N_10568,N_9571,N_9045);
nand U10569 (N_10569,N_8965,N_9406);
or U10570 (N_10570,N_7589,N_8149);
and U10571 (N_10571,N_5684,N_7096);
nand U10572 (N_10572,N_9046,N_7643);
nor U10573 (N_10573,N_6306,N_6405);
nand U10574 (N_10574,N_9374,N_9703);
and U10575 (N_10575,N_5285,N_5518);
nand U10576 (N_10576,N_9994,N_9884);
xor U10577 (N_10577,N_7865,N_7935);
xor U10578 (N_10578,N_8717,N_9818);
and U10579 (N_10579,N_8486,N_7577);
and U10580 (N_10580,N_5152,N_9323);
or U10581 (N_10581,N_6653,N_7329);
xor U10582 (N_10582,N_6202,N_7503);
and U10583 (N_10583,N_8870,N_6408);
xor U10584 (N_10584,N_8935,N_8016);
and U10585 (N_10585,N_9378,N_7955);
nor U10586 (N_10586,N_6026,N_8652);
and U10587 (N_10587,N_8073,N_7279);
and U10588 (N_10588,N_7786,N_5441);
and U10589 (N_10589,N_6414,N_9132);
xnor U10590 (N_10590,N_8261,N_7308);
xor U10591 (N_10591,N_9474,N_9353);
and U10592 (N_10592,N_5101,N_8753);
or U10593 (N_10593,N_5075,N_7282);
nand U10594 (N_10594,N_8213,N_5829);
nor U10595 (N_10595,N_5012,N_5472);
nand U10596 (N_10596,N_8275,N_8517);
or U10597 (N_10597,N_5424,N_8262);
nor U10598 (N_10598,N_7741,N_9860);
xnor U10599 (N_10599,N_7943,N_6168);
nand U10600 (N_10600,N_9550,N_7857);
nand U10601 (N_10601,N_5775,N_9676);
or U10602 (N_10602,N_9710,N_5446);
nand U10603 (N_10603,N_7193,N_9880);
nor U10604 (N_10604,N_6031,N_9040);
nor U10605 (N_10605,N_6623,N_5548);
or U10606 (N_10606,N_8135,N_8732);
and U10607 (N_10607,N_6186,N_8088);
nor U10608 (N_10608,N_6244,N_8151);
xor U10609 (N_10609,N_8927,N_7386);
nand U10610 (N_10610,N_8739,N_7772);
and U10611 (N_10611,N_9570,N_5923);
and U10612 (N_10612,N_9253,N_6032);
xnor U10613 (N_10613,N_8772,N_7144);
and U10614 (N_10614,N_8078,N_7100);
and U10615 (N_10615,N_6373,N_6477);
nor U10616 (N_10616,N_5013,N_6987);
nand U10617 (N_10617,N_8273,N_8556);
and U10618 (N_10618,N_6341,N_7372);
and U10619 (N_10619,N_6371,N_8032);
nor U10620 (N_10620,N_9913,N_9205);
or U10621 (N_10621,N_5537,N_7777);
xor U10622 (N_10622,N_9843,N_7298);
and U10623 (N_10623,N_9832,N_6070);
xnor U10624 (N_10624,N_6061,N_5647);
or U10625 (N_10625,N_8554,N_9734);
xor U10626 (N_10626,N_9029,N_9534);
nand U10627 (N_10627,N_8710,N_8641);
and U10628 (N_10628,N_6142,N_6012);
nor U10629 (N_10629,N_7717,N_6268);
nor U10630 (N_10630,N_9964,N_7261);
or U10631 (N_10631,N_8192,N_9128);
and U10632 (N_10632,N_5245,N_9032);
or U10633 (N_10633,N_8630,N_5671);
xor U10634 (N_10634,N_6108,N_7800);
or U10635 (N_10635,N_8743,N_5186);
xnor U10636 (N_10636,N_5546,N_5411);
xor U10637 (N_10637,N_5470,N_5791);
xnor U10638 (N_10638,N_8602,N_5536);
xnor U10639 (N_10639,N_5996,N_5723);
nand U10640 (N_10640,N_9631,N_5043);
nand U10641 (N_10641,N_9494,N_9634);
nor U10642 (N_10642,N_7136,N_5064);
nand U10643 (N_10643,N_8775,N_7219);
nand U10644 (N_10644,N_5278,N_8990);
or U10645 (N_10645,N_8900,N_6921);
nand U10646 (N_10646,N_8968,N_7299);
nand U10647 (N_10647,N_7292,N_5792);
or U10648 (N_10648,N_7432,N_5676);
nand U10649 (N_10649,N_6367,N_9066);
nor U10650 (N_10650,N_5890,N_6827);
xor U10651 (N_10651,N_7037,N_9404);
nand U10652 (N_10652,N_5925,N_6778);
or U10653 (N_10653,N_9757,N_6592);
nor U10654 (N_10654,N_5166,N_9503);
xnor U10655 (N_10655,N_6432,N_8828);
xnor U10656 (N_10656,N_5408,N_5395);
and U10657 (N_10657,N_8885,N_7844);
or U10658 (N_10658,N_6324,N_8443);
nand U10659 (N_10659,N_7153,N_9014);
nand U10660 (N_10660,N_7426,N_5465);
nor U10661 (N_10661,N_6029,N_8937);
and U10662 (N_10662,N_9553,N_6694);
and U10663 (N_10663,N_6329,N_9929);
xnor U10664 (N_10664,N_9685,N_7652);
xnor U10665 (N_10665,N_8224,N_6001);
nor U10666 (N_10666,N_9738,N_7165);
nor U10667 (N_10667,N_7211,N_5916);
xor U10668 (N_10668,N_9277,N_6246);
or U10669 (N_10669,N_8956,N_6045);
nand U10670 (N_10670,N_5981,N_6817);
nor U10671 (N_10671,N_8758,N_6180);
nor U10672 (N_10672,N_9431,N_5756);
nand U10673 (N_10673,N_7421,N_9466);
and U10674 (N_10674,N_8420,N_8253);
nand U10675 (N_10675,N_8477,N_5913);
or U10676 (N_10676,N_9641,N_7902);
and U10677 (N_10677,N_9027,N_7027);
and U10678 (N_10678,N_8607,N_6227);
nand U10679 (N_10679,N_9559,N_6103);
and U10680 (N_10680,N_9191,N_9414);
nand U10681 (N_10681,N_7780,N_9152);
xnor U10682 (N_10682,N_6086,N_5817);
or U10683 (N_10683,N_5401,N_9472);
xor U10684 (N_10684,N_6438,N_6774);
or U10685 (N_10685,N_9957,N_7041);
and U10686 (N_10686,N_6640,N_9816);
and U10687 (N_10687,N_9022,N_9733);
nor U10688 (N_10688,N_9883,N_8802);
or U10689 (N_10689,N_7763,N_9613);
nand U10690 (N_10690,N_6081,N_7950);
nor U10691 (N_10691,N_9470,N_9137);
xnor U10692 (N_10692,N_8863,N_8304);
nand U10693 (N_10693,N_8417,N_8111);
nand U10694 (N_10694,N_6313,N_9112);
or U10695 (N_10695,N_8328,N_6215);
and U10696 (N_10696,N_8845,N_8168);
xnor U10697 (N_10697,N_7719,N_8156);
or U10698 (N_10698,N_6923,N_6368);
xnor U10699 (N_10699,N_6245,N_9162);
nor U10700 (N_10700,N_8664,N_7613);
xor U10701 (N_10701,N_5878,N_9870);
or U10702 (N_10702,N_8339,N_5995);
and U10703 (N_10703,N_8784,N_7256);
and U10704 (N_10704,N_6572,N_6781);
or U10705 (N_10705,N_5313,N_5953);
or U10706 (N_10706,N_9327,N_9707);
xor U10707 (N_10707,N_7611,N_5495);
or U10708 (N_10708,N_5379,N_8218);
or U10709 (N_10709,N_5593,N_9172);
and U10710 (N_10710,N_7250,N_8629);
and U10711 (N_10711,N_9320,N_6444);
xnor U10712 (N_10712,N_5071,N_6645);
xor U10713 (N_10713,N_9338,N_8254);
or U10714 (N_10714,N_9735,N_9467);
nor U10715 (N_10715,N_8119,N_5828);
or U10716 (N_10716,N_7441,N_7190);
or U10717 (N_10717,N_7649,N_7076);
and U10718 (N_10718,N_7123,N_9188);
or U10719 (N_10719,N_5241,N_9629);
and U10720 (N_10720,N_6800,N_5261);
nor U10721 (N_10721,N_6972,N_9797);
xnor U10722 (N_10722,N_8767,N_8489);
nor U10723 (N_10723,N_9807,N_6349);
nand U10724 (N_10724,N_5917,N_6413);
nor U10725 (N_10725,N_9551,N_8436);
xor U10726 (N_10726,N_9740,N_9213);
nor U10727 (N_10727,N_7055,N_6715);
xor U10728 (N_10728,N_8604,N_5045);
xor U10729 (N_10729,N_5429,N_5886);
nand U10730 (N_10730,N_7412,N_5098);
or U10731 (N_10731,N_9611,N_7084);
xor U10732 (N_10732,N_7557,N_6859);
or U10733 (N_10733,N_5643,N_7473);
xnor U10734 (N_10734,N_9211,N_9799);
nor U10735 (N_10735,N_9993,N_6969);
and U10736 (N_10736,N_6638,N_7829);
nand U10737 (N_10737,N_7357,N_5584);
nor U10738 (N_10738,N_9618,N_8407);
or U10739 (N_10739,N_8971,N_5749);
and U10740 (N_10740,N_8406,N_5940);
or U10741 (N_10741,N_6092,N_7672);
nand U10742 (N_10742,N_6591,N_6017);
nand U10743 (N_10743,N_8576,N_6684);
nor U10744 (N_10744,N_7737,N_5315);
nand U10745 (N_10745,N_6550,N_8022);
and U10746 (N_10746,N_5728,N_8649);
and U10747 (N_10747,N_7125,N_5484);
nor U10748 (N_10748,N_7728,N_7035);
xor U10749 (N_10749,N_8409,N_9688);
and U10750 (N_10750,N_9076,N_5895);
and U10751 (N_10751,N_7213,N_6025);
and U10752 (N_10752,N_5237,N_9363);
xnor U10753 (N_10753,N_5588,N_9936);
and U10754 (N_10754,N_5813,N_7527);
or U10755 (N_10755,N_6364,N_5345);
and U10756 (N_10756,N_6106,N_9033);
xor U10757 (N_10757,N_6545,N_9085);
nor U10758 (N_10758,N_5160,N_9772);
and U10759 (N_10759,N_5112,N_5664);
xnor U10760 (N_10760,N_7958,N_6563);
nand U10761 (N_10761,N_7025,N_6882);
nand U10762 (N_10762,N_8476,N_8292);
nor U10763 (N_10763,N_5360,N_6980);
nor U10764 (N_10764,N_7960,N_5079);
nand U10765 (N_10765,N_5375,N_5877);
or U10766 (N_10766,N_5029,N_9008);
nor U10767 (N_10767,N_8013,N_9614);
nor U10768 (N_10768,N_5496,N_8045);
nor U10769 (N_10769,N_5622,N_7091);
xor U10770 (N_10770,N_6897,N_8198);
nor U10771 (N_10771,N_9567,N_9888);
nor U10772 (N_10772,N_7653,N_7847);
xor U10773 (N_10773,N_7931,N_9593);
nor U10774 (N_10774,N_7485,N_5273);
or U10775 (N_10775,N_9247,N_5035);
or U10776 (N_10776,N_9461,N_9649);
nor U10777 (N_10777,N_9699,N_6043);
xor U10778 (N_10778,N_6910,N_8474);
nor U10779 (N_10779,N_5168,N_5761);
and U10780 (N_10780,N_6634,N_5450);
nor U10781 (N_10781,N_6554,N_8699);
nand U10782 (N_10782,N_7051,N_8867);
nor U10783 (N_10783,N_7944,N_7572);
nand U10784 (N_10784,N_9104,N_9894);
and U10785 (N_10785,N_7667,N_5614);
xor U10786 (N_10786,N_6232,N_8247);
or U10787 (N_10787,N_5818,N_5019);
xor U10788 (N_10788,N_7215,N_9197);
or U10789 (N_10789,N_8049,N_7546);
xnor U10790 (N_10790,N_8435,N_8757);
nand U10791 (N_10791,N_5506,N_8915);
xor U10792 (N_10792,N_9109,N_5451);
nand U10793 (N_10793,N_8118,N_5935);
nor U10794 (N_10794,N_7159,N_6327);
or U10795 (N_10795,N_7507,N_8010);
or U10796 (N_10796,N_8089,N_7947);
nor U10797 (N_10797,N_9392,N_8290);
or U10798 (N_10798,N_8176,N_7106);
nand U10799 (N_10799,N_8133,N_6189);
nand U10800 (N_10800,N_6668,N_8488);
and U10801 (N_10801,N_6037,N_5782);
or U10802 (N_10802,N_9347,N_8959);
nor U10803 (N_10803,N_7230,N_5540);
nor U10804 (N_10804,N_7348,N_9896);
or U10805 (N_10805,N_6294,N_7647);
nor U10806 (N_10806,N_5980,N_8449);
or U10807 (N_10807,N_9794,N_5816);
nor U10808 (N_10808,N_6758,N_7726);
xor U10809 (N_10809,N_8276,N_9248);
nand U10810 (N_10810,N_9704,N_8295);
and U10811 (N_10811,N_8882,N_5812);
or U10812 (N_10812,N_7151,N_6759);
and U10813 (N_10813,N_9903,N_6484);
or U10814 (N_10814,N_8635,N_6994);
xnor U10815 (N_10815,N_9822,N_5526);
and U10816 (N_10816,N_8472,N_7097);
nor U10817 (N_10817,N_8114,N_7725);
and U10818 (N_10818,N_8902,N_5167);
nand U10819 (N_10819,N_6829,N_9268);
and U10820 (N_10820,N_6146,N_6753);
xnor U10821 (N_10821,N_8200,N_9070);
and U10822 (N_10822,N_9396,N_5037);
or U10823 (N_10823,N_9790,N_5210);
nand U10824 (N_10824,N_8067,N_7235);
xnor U10825 (N_10825,N_9102,N_8364);
xnor U10826 (N_10826,N_6879,N_9078);
and U10827 (N_10827,N_7892,N_5533);
xor U10828 (N_10828,N_9726,N_9367);
nor U10829 (N_10829,N_5377,N_5570);
nand U10830 (N_10830,N_8663,N_6326);
xnor U10831 (N_10831,N_8383,N_6028);
or U10832 (N_10832,N_8890,N_9361);
or U10833 (N_10833,N_9263,N_6365);
xor U10834 (N_10834,N_5314,N_5240);
and U10835 (N_10835,N_9505,N_7744);
or U10836 (N_10836,N_7411,N_7543);
nand U10837 (N_10837,N_8455,N_7139);
xor U10838 (N_10838,N_5849,N_9187);
or U10839 (N_10839,N_8142,N_8811);
nand U10840 (N_10840,N_6553,N_5641);
nor U10841 (N_10841,N_5449,N_9996);
and U10842 (N_10842,N_5399,N_8355);
nor U10843 (N_10843,N_7641,N_6916);
xnor U10844 (N_10844,N_6782,N_8589);
and U10845 (N_10845,N_6125,N_8700);
and U10846 (N_10846,N_9455,N_7952);
xor U10847 (N_10847,N_6095,N_8875);
and U10848 (N_10848,N_9301,N_7818);
and U10849 (N_10849,N_7816,N_8620);
and U10850 (N_10850,N_6469,N_9155);
nand U10851 (N_10851,N_8020,N_7118);
nand U10852 (N_10852,N_9863,N_7820);
and U10853 (N_10853,N_5982,N_8345);
nand U10854 (N_10854,N_8112,N_7881);
or U10855 (N_10855,N_5887,N_5417);
or U10856 (N_10856,N_5233,N_5932);
or U10857 (N_10857,N_7673,N_7526);
and U10858 (N_10858,N_5030,N_7564);
nand U10859 (N_10859,N_7538,N_9985);
or U10860 (N_10860,N_5759,N_7152);
and U10861 (N_10861,N_9158,N_6844);
xnor U10862 (N_10862,N_9202,N_6956);
nor U10863 (N_10863,N_7794,N_7627);
nor U10864 (N_10864,N_8725,N_9930);
nand U10865 (N_10865,N_9514,N_9440);
nand U10866 (N_10866,N_7368,N_7797);
or U10867 (N_10867,N_6559,N_6074);
nor U10868 (N_10868,N_6119,N_8701);
nand U10869 (N_10869,N_5626,N_9881);
nand U10870 (N_10870,N_8411,N_5426);
or U10871 (N_10871,N_6869,N_8573);
or U10872 (N_10872,N_7742,N_7723);
and U10873 (N_10873,N_9300,N_5777);
and U10874 (N_10874,N_6726,N_8857);
and U10875 (N_10875,N_5617,N_7034);
xor U10876 (N_10876,N_7731,N_9803);
nand U10877 (N_10877,N_7442,N_8076);
xnor U10878 (N_10878,N_5562,N_9376);
nand U10879 (N_10879,N_8115,N_6454);
nand U10880 (N_10880,N_9808,N_5300);
and U10881 (N_10881,N_7360,N_8688);
and U10882 (N_10882,N_5516,N_8823);
or U10883 (N_10883,N_8524,N_6866);
xor U10884 (N_10884,N_8492,N_9026);
xnor U10885 (N_10885,N_8666,N_7555);
or U10886 (N_10886,N_5915,N_9852);
nor U10887 (N_10887,N_7799,N_7906);
and U10888 (N_10888,N_5033,N_5123);
and U10889 (N_10889,N_6878,N_9260);
xnor U10890 (N_10890,N_8528,N_5763);
nand U10891 (N_10891,N_5466,N_8038);
xor U10892 (N_10892,N_8319,N_6934);
xnor U10893 (N_10893,N_9159,N_7511);
and U10894 (N_10894,N_8698,N_9336);
nand U10895 (N_10895,N_8946,N_9661);
nor U10896 (N_10896,N_5610,N_5638);
or U10897 (N_10897,N_7119,N_6514);
and U10898 (N_10898,N_6483,N_5501);
xor U10899 (N_10899,N_6595,N_8223);
nor U10900 (N_10900,N_7595,N_6193);
nand U10901 (N_10901,N_9608,N_7748);
xnor U10902 (N_10902,N_5657,N_5716);
nor U10903 (N_10903,N_6136,N_9342);
nand U10904 (N_10904,N_7831,N_5908);
and U10905 (N_10905,N_9380,N_6497);
nand U10906 (N_10906,N_9120,N_9528);
or U10907 (N_10907,N_8578,N_7346);
or U10908 (N_10908,N_5673,N_6607);
or U10909 (N_10909,N_5006,N_6184);
nand U10910 (N_10910,N_9654,N_7288);
and U10911 (N_10911,N_5148,N_8043);
nand U10912 (N_10912,N_6449,N_8503);
and U10913 (N_10913,N_8130,N_6452);
xor U10914 (N_10914,N_7087,N_7438);
nand U10915 (N_10915,N_7205,N_6871);
and U10916 (N_10916,N_7638,N_9218);
and U10917 (N_10917,N_6488,N_5843);
xor U10918 (N_10918,N_6902,N_6502);
xor U10919 (N_10919,N_5034,N_8822);
xor U10920 (N_10920,N_9918,N_8525);
or U10921 (N_10921,N_5613,N_8922);
xnor U10922 (N_10922,N_5538,N_8033);
nand U10923 (N_10923,N_6798,N_8756);
nand U10924 (N_10924,N_8105,N_8103);
and U10925 (N_10925,N_8376,N_9947);
xor U10926 (N_10926,N_6907,N_8054);
or U10927 (N_10927,N_7247,N_6068);
or U10928 (N_10928,N_7471,N_8374);
nand U10929 (N_10929,N_8110,N_6430);
nand U10930 (N_10930,N_7137,N_9177);
xnor U10931 (N_10931,N_5493,N_8657);
or U10932 (N_10932,N_7644,N_6524);
or U10933 (N_10933,N_5250,N_5198);
nand U10934 (N_10934,N_8349,N_5946);
nand U10935 (N_10935,N_5292,N_7570);
nor U10936 (N_10936,N_7588,N_6158);
nand U10937 (N_10937,N_8127,N_6975);
or U10938 (N_10938,N_7657,N_6508);
nor U10939 (N_10939,N_6493,N_7809);
nand U10940 (N_10940,N_5820,N_8031);
and U10941 (N_10941,N_7281,N_5520);
xor U10942 (N_10942,N_9939,N_5736);
xnor U10943 (N_10943,N_5418,N_5039);
nand U10944 (N_10944,N_9660,N_7791);
nand U10945 (N_10945,N_6172,N_5402);
xnor U10946 (N_10946,N_6394,N_9756);
and U10947 (N_10947,N_5114,N_9166);
and U10948 (N_10948,N_7341,N_8818);
xor U10949 (N_10949,N_9490,N_6788);
xnor U10950 (N_10950,N_8855,N_9091);
and U10951 (N_10951,N_9960,N_9531);
xor U10952 (N_10952,N_8622,N_9907);
xor U10953 (N_10953,N_9577,N_7033);
xnor U10954 (N_10954,N_6111,N_8248);
and U10955 (N_10955,N_6318,N_5855);
and U10956 (N_10956,N_5214,N_9778);
or U10957 (N_10957,N_9410,N_6495);
and U10958 (N_10958,N_9887,N_6358);
or U10959 (N_10959,N_7301,N_5048);
nor U10960 (N_10960,N_6820,N_7210);
and U10961 (N_10961,N_9237,N_5365);
or U10962 (N_10962,N_8060,N_6649);
xnor U10963 (N_10963,N_5130,N_8737);
and U10964 (N_10964,N_5055,N_9387);
nor U10965 (N_10965,N_6557,N_8939);
xnor U10966 (N_10966,N_5264,N_7959);
or U10967 (N_10967,N_8204,N_5776);
or U10968 (N_10968,N_5713,N_8083);
nand U10969 (N_10969,N_6024,N_9023);
nor U10970 (N_10970,N_5359,N_7304);
and U10971 (N_10971,N_9443,N_7940);
nand U10972 (N_10972,N_8545,N_9042);
nor U10973 (N_10973,N_9457,N_5290);
nor U10974 (N_10974,N_7897,N_7604);
xor U10975 (N_10975,N_6500,N_8005);
nand U10976 (N_10976,N_7796,N_8308);
xnor U10977 (N_10977,N_7284,N_7227);
or U10978 (N_10978,N_6390,N_7612);
nor U10979 (N_10979,N_9542,N_8136);
xnor U10980 (N_10980,N_7150,N_6932);
nor U10981 (N_10981,N_5519,N_8773);
or U10982 (N_10982,N_6914,N_6719);
nand U10983 (N_10983,N_6588,N_5997);
nor U10984 (N_10984,N_5529,N_6894);
or U10985 (N_10985,N_5648,N_7040);
or U10986 (N_10986,N_9339,N_7963);
nor U10987 (N_10987,N_9665,N_5977);
or U10988 (N_10988,N_8297,N_5773);
xor U10989 (N_10989,N_7313,N_9189);
nor U10990 (N_10990,N_6323,N_7905);
or U10991 (N_10991,N_6723,N_8787);
or U10992 (N_10992,N_9157,N_5304);
or U10993 (N_10993,N_5195,N_5255);
or U10994 (N_10994,N_8587,N_7114);
and U10995 (N_10995,N_7072,N_8711);
nor U10996 (N_10996,N_5224,N_5909);
nor U10997 (N_10997,N_5549,N_7355);
or U10998 (N_10998,N_8730,N_5984);
or U10999 (N_10999,N_8431,N_9509);
and U11000 (N_11000,N_6345,N_6625);
nand U11001 (N_11001,N_5200,N_6709);
and U11002 (N_11002,N_6143,N_8797);
or U11003 (N_11003,N_9708,N_7452);
nor U11004 (N_11004,N_5087,N_8669);
nand U11005 (N_11005,N_9655,N_9900);
or U11006 (N_11006,N_7195,N_9244);
or U11007 (N_11007,N_7990,N_6003);
xnor U11008 (N_11008,N_8047,N_6992);
or U11009 (N_11009,N_7000,N_7133);
or U11010 (N_11010,N_9233,N_7188);
nor U11011 (N_11011,N_5884,N_6412);
or U11012 (N_11012,N_6130,N_6805);
and U11013 (N_11013,N_7768,N_6152);
nor U11014 (N_11014,N_8592,N_9951);
xnor U11015 (N_11015,N_7878,N_8097);
nand U11016 (N_11016,N_6221,N_6038);
or U11017 (N_11017,N_7327,N_7779);
or U11018 (N_11018,N_9879,N_8086);
xnor U11019 (N_11019,N_6311,N_6810);
or U11020 (N_11020,N_7351,N_8952);
and U11021 (N_11021,N_6632,N_6218);
and U11022 (N_11022,N_8942,N_5082);
xor U11023 (N_11023,N_5042,N_5318);
nor U11024 (N_11024,N_8826,N_6407);
or U11025 (N_11025,N_8280,N_9096);
and U11026 (N_11026,N_8859,N_8094);
nand U11027 (N_11027,N_6370,N_6903);
or U11028 (N_11028,N_5779,N_7970);
nand U11029 (N_11029,N_9314,N_5682);
and U11030 (N_11030,N_9637,N_8344);
xnor U11031 (N_11031,N_6767,N_9823);
nor U11032 (N_11032,N_7141,N_7592);
or U11033 (N_11033,N_9307,N_8046);
nor U11034 (N_11034,N_7601,N_7713);
and U11035 (N_11035,N_5448,N_8061);
and U11036 (N_11036,N_7624,N_8761);
or U11037 (N_11037,N_6602,N_6547);
xnor U11038 (N_11038,N_8373,N_6678);
and U11039 (N_11039,N_5905,N_5298);
xor U11040 (N_11040,N_7109,N_9499);
xor U11041 (N_11041,N_5988,N_8953);
nor U11042 (N_11042,N_6499,N_7131);
and U11043 (N_11043,N_8153,N_8181);
or U11044 (N_11044,N_9425,N_7053);
xnor U11045 (N_11045,N_6635,N_6872);
and U11046 (N_11046,N_7743,N_5109);
nor U11047 (N_11047,N_5325,N_9437);
and U11048 (N_11048,N_7244,N_7584);
nor U11049 (N_11049,N_5696,N_9274);
and U11050 (N_11050,N_6892,N_8844);
or U11051 (N_11051,N_9399,N_7458);
or U11052 (N_11052,N_7490,N_7130);
nor U11053 (N_11053,N_8057,N_6832);
xnor U11054 (N_11054,N_7746,N_6248);
nand U11055 (N_11055,N_7318,N_5569);
xnor U11056 (N_11056,N_7127,N_6272);
and U11057 (N_11057,N_8452,N_8036);
and U11058 (N_11058,N_8841,N_7121);
and U11059 (N_11059,N_7253,N_8551);
nor U11060 (N_11060,N_9924,N_6672);
nor U11061 (N_11061,N_5652,N_9423);
nand U11062 (N_11062,N_7594,N_6841);
nor U11063 (N_11063,N_6016,N_5630);
xor U11064 (N_11064,N_7496,N_8836);
nor U11065 (N_11065,N_8755,N_8306);
nor U11066 (N_11066,N_7046,N_9331);
nand U11067 (N_11067,N_8346,N_8301);
xor U11068 (N_11068,N_5528,N_8817);
nor U11069 (N_11069,N_9400,N_5337);
or U11070 (N_11070,N_7855,N_9176);
nand U11071 (N_11071,N_6424,N_5659);
nor U11072 (N_11072,N_6521,N_8895);
nand U11073 (N_11073,N_6253,N_9958);
and U11074 (N_11074,N_9533,N_5832);
nand U11075 (N_11075,N_5085,N_8187);
or U11076 (N_11076,N_8367,N_7453);
and U11077 (N_11077,N_9774,N_5552);
and U11078 (N_11078,N_9858,N_7942);
and U11079 (N_11079,N_7332,N_9910);
xor U11080 (N_11080,N_8812,N_5138);
nor U11081 (N_11081,N_8278,N_7110);
and U11082 (N_11082,N_9765,N_6328);
xor U11083 (N_11083,N_7945,N_8040);
nand U11084 (N_11084,N_9632,N_7456);
xnor U11085 (N_11085,N_5697,N_7864);
nor U11086 (N_11086,N_5861,N_8371);
nand U11087 (N_11087,N_8379,N_5898);
or U11088 (N_11088,N_8027,N_7569);
or U11089 (N_11089,N_9873,N_8557);
nor U11090 (N_11090,N_9751,N_8969);
nor U11091 (N_11091,N_6949,N_8124);
nand U11092 (N_11092,N_9473,N_8899);
and U11093 (N_11093,N_8833,N_6797);
nor U11094 (N_11094,N_6179,N_8941);
or U11095 (N_11095,N_7908,N_9403);
xnor U11096 (N_11096,N_5338,N_7300);
nor U11097 (N_11097,N_6415,N_9167);
xnor U11098 (N_11098,N_8887,N_8896);
xnor U11099 (N_11099,N_6058,N_7231);
or U11100 (N_11100,N_5718,N_7899);
xor U11101 (N_11101,N_6780,N_9052);
nand U11102 (N_11102,N_8926,N_9961);
nor U11103 (N_11103,N_6322,N_8783);
and U11104 (N_11104,N_7270,N_6699);
nand U11105 (N_11105,N_5415,N_8214);
and U11106 (N_11106,N_7128,N_9908);
xor U11107 (N_11107,N_5627,N_9568);
nand U11108 (N_11108,N_6562,N_5068);
or U11109 (N_11109,N_8847,N_8165);
nand U11110 (N_11110,N_9830,N_6576);
and U11111 (N_11111,N_9972,N_6953);
nand U11112 (N_11112,N_7022,N_8305);
nand U11113 (N_11113,N_8916,N_9598);
and U11114 (N_11114,N_7129,N_8713);
and U11115 (N_11115,N_9601,N_9282);
and U11116 (N_11116,N_7918,N_8569);
nand U11117 (N_11117,N_7061,N_6235);
nor U11118 (N_11118,N_7236,N_8901);
nor U11119 (N_11119,N_8809,N_5578);
or U11120 (N_11120,N_6100,N_5044);
nand U11121 (N_11121,N_6887,N_6749);
xnor U11122 (N_11122,N_9131,N_6991);
and U11123 (N_11123,N_9217,N_8790);
nor U11124 (N_11124,N_9445,N_7364);
xnor U11125 (N_11125,N_7811,N_5906);
and U11126 (N_11126,N_9053,N_6739);
nand U11127 (N_11127,N_8981,N_7462);
nand U11128 (N_11128,N_9677,N_8129);
and U11129 (N_11129,N_9391,N_5004);
and U11130 (N_11130,N_7013,N_8925);
nor U11131 (N_11131,N_6166,N_7628);
and U11132 (N_11132,N_5938,N_6183);
xor U11133 (N_11133,N_9265,N_5810);
nor U11134 (N_11134,N_7415,N_6927);
and U11135 (N_11135,N_7964,N_8087);
xnor U11136 (N_11136,N_6611,N_9346);
and U11137 (N_11137,N_8681,N_7579);
nor U11138 (N_11138,N_6255,N_8368);
xnor U11139 (N_11139,N_6787,N_5246);
xnor U11140 (N_11140,N_8815,N_5342);
nand U11141 (N_11141,N_8307,N_8594);
xor U11142 (N_11142,N_7832,N_7827);
xor U11143 (N_11143,N_6140,N_9130);
or U11144 (N_11144,N_5653,N_8995);
and U11145 (N_11145,N_6181,N_5185);
nand U11146 (N_11146,N_5631,N_9182);
xor U11147 (N_11147,N_8350,N_5772);
nor U11148 (N_11148,N_7385,N_8914);
nand U11149 (N_11149,N_8001,N_5937);
or U11150 (N_11150,N_8928,N_7971);
nand U11151 (N_11151,N_6560,N_6748);
nor U11152 (N_11152,N_5721,N_8338);
and U11153 (N_11153,N_6163,N_9124);
nand U11154 (N_11154,N_5608,N_9379);
or U11155 (N_11155,N_5184,N_9308);
nand U11156 (N_11156,N_5180,N_8205);
nand U11157 (N_11157,N_9071,N_8128);
nand U11158 (N_11158,N_8712,N_9651);
nor U11159 (N_11159,N_8384,N_6223);
nand U11160 (N_11160,N_9828,N_5888);
nand U11161 (N_11161,N_5226,N_7183);
xnor U11162 (N_11162,N_5482,N_7160);
nand U11163 (N_11163,N_8093,N_9409);
nand U11164 (N_11164,N_7056,N_9084);
and U11165 (N_11165,N_9935,N_6082);
nor U11166 (N_11166,N_5308,N_5139);
xor U11167 (N_11167,N_6819,N_9874);
nor U11168 (N_11168,N_7320,N_8816);
or U11169 (N_11169,N_7465,N_5508);
or U11170 (N_11170,N_7849,N_7835);
or U11171 (N_11171,N_9868,N_5122);
nand U11172 (N_11172,N_7460,N_7074);
nor U11173 (N_11173,N_6666,N_6395);
nor U11174 (N_11174,N_5190,N_8150);
nand U11175 (N_11175,N_5692,N_5284);
or U11176 (N_11176,N_5866,N_8499);
xnor U11177 (N_11177,N_9360,N_6149);
or U11178 (N_11178,N_5698,N_5556);
or U11179 (N_11179,N_5259,N_7722);
nand U11180 (N_11180,N_7012,N_9520);
xor U11181 (N_11181,N_6581,N_6396);
xor U11182 (N_11182,N_8365,N_8842);
xor U11183 (N_11183,N_5478,N_8419);
or U11184 (N_11184,N_7981,N_7623);
xor U11185 (N_11185,N_7264,N_7031);
nor U11186 (N_11186,N_5274,N_9923);
or U11187 (N_11187,N_5732,N_6386);
nand U11188 (N_11188,N_6539,N_9971);
nand U11189 (N_11189,N_7957,N_8504);
nor U11190 (N_11190,N_8546,N_5199);
nand U11191 (N_11191,N_5440,N_9281);
xnor U11192 (N_11192,N_9650,N_7049);
nand U11193 (N_11193,N_5545,N_9878);
nor U11194 (N_11194,N_9432,N_9151);
nand U11195 (N_11195,N_6177,N_9006);
nand U11196 (N_11196,N_5694,N_5733);
xnor U11197 (N_11197,N_8125,N_8148);
nand U11198 (N_11198,N_6808,N_8883);
and U11199 (N_11199,N_7686,N_7798);
nor U11200 (N_11200,N_5522,N_7982);
nor U11201 (N_11201,N_9684,N_6733);
xnor U11202 (N_11202,N_5120,N_7039);
xnor U11203 (N_11203,N_5987,N_6752);
nor U11204 (N_11204,N_6501,N_7834);
xor U11205 (N_11205,N_6885,N_5203);
or U11206 (N_11206,N_9481,N_9926);
nand U11207 (N_11207,N_8577,N_9345);
and U11208 (N_11208,N_9627,N_9658);
xnor U11209 (N_11209,N_5726,N_5963);
or U11210 (N_11210,N_5435,N_7518);
or U11211 (N_11211,N_5802,N_9390);
nand U11212 (N_11212,N_9364,N_6109);
nor U11213 (N_11213,N_6990,N_7760);
nand U11214 (N_11214,N_9983,N_9876);
and U11215 (N_11215,N_9578,N_6116);
and U11216 (N_11216,N_5525,N_5352);
or U11217 (N_11217,N_5551,N_6984);
xnor U11218 (N_11218,N_7654,N_5706);
and U11219 (N_11219,N_8391,N_7437);
nand U11220 (N_11220,N_6558,N_5346);
or U11221 (N_11221,N_7425,N_6868);
or U11222 (N_11222,N_7494,N_8303);
or U11223 (N_11223,N_9558,N_5286);
nand U11224 (N_11224,N_9356,N_5958);
nor U11225 (N_11225,N_9051,N_8705);
or U11226 (N_11226,N_9666,N_6612);
xnor U11227 (N_11227,N_5969,N_9311);
and U11228 (N_11228,N_9662,N_5394);
nand U11229 (N_11229,N_7330,N_8535);
xnor U11230 (N_11230,N_7200,N_7479);
nor U11231 (N_11231,N_5612,N_7069);
and U11232 (N_11232,N_7636,N_6544);
xnor U11233 (N_11233,N_8467,N_5591);
nor U11234 (N_11234,N_8632,N_7180);
xor U11235 (N_11235,N_7705,N_9103);
nand U11236 (N_11236,N_9712,N_5162);
or U11237 (N_11237,N_5956,N_7081);
and U11238 (N_11238,N_6093,N_6282);
and U11239 (N_11239,N_7519,N_5930);
nand U11240 (N_11240,N_8911,N_8521);
or U11241 (N_11241,N_7598,N_5500);
and U11242 (N_11242,N_8270,N_6853);
and U11243 (N_11243,N_8706,N_6812);
or U11244 (N_11244,N_8279,N_7126);
xor U11245 (N_11245,N_8628,N_8056);
nand U11246 (N_11246,N_5268,N_5494);
nand U11247 (N_11247,N_5677,N_6154);
xor U11248 (N_11248,N_9544,N_5254);
nor U11249 (N_11249,N_9242,N_6847);
and U11250 (N_11250,N_9689,N_5639);
xnor U11251 (N_11251,N_6435,N_8456);
or U11252 (N_11252,N_6834,N_5406);
nand U11253 (N_11253,N_8852,N_9178);
xor U11254 (N_11254,N_7409,N_8117);
or U11255 (N_11255,N_7574,N_5223);
or U11256 (N_11256,N_9161,N_5217);
xor U11257 (N_11257,N_8614,N_9280);
xnor U11258 (N_11258,N_8445,N_5753);
or U11259 (N_11259,N_5297,N_8495);
or U11260 (N_11260,N_6121,N_8009);
nor U11261 (N_11261,N_5368,N_5363);
nor U11262 (N_11262,N_7382,N_8684);
nand U11263 (N_11263,N_8516,N_8548);
or U11264 (N_11264,N_9984,N_9298);
and U11265 (N_11265,N_9107,N_9781);
or U11266 (N_11266,N_9385,N_5853);
nand U11267 (N_11267,N_6170,N_6862);
xor U11268 (N_11268,N_8479,N_7692);
and U11269 (N_11269,N_9869,N_8238);
nor U11270 (N_11270,N_7689,N_8744);
nor U11271 (N_11271,N_5801,N_6474);
nor U11272 (N_11272,N_5409,N_8161);
nor U11273 (N_11273,N_9002,N_5565);
nand U11274 (N_11274,N_6207,N_7879);
and U11275 (N_11275,N_9839,N_7387);
xor U11276 (N_11276,N_7175,N_6608);
nand U11277 (N_11277,N_9563,N_7994);
nand U11278 (N_11278,N_9402,N_6564);
xor U11279 (N_11279,N_9905,N_6233);
nand U11280 (N_11280,N_5028,N_6124);
nor U11281 (N_11281,N_6541,N_5339);
nor U11282 (N_11282,N_6209,N_7367);
and U11283 (N_11283,N_8144,N_8157);
nand U11284 (N_11284,N_6225,N_6150);
xor U11285 (N_11285,N_5632,N_5717);
nand U11286 (N_11286,N_5031,N_8102);
and U11287 (N_11287,N_5145,N_5381);
xnor U11288 (N_11288,N_6676,N_8661);
nand U11289 (N_11289,N_9292,N_7597);
or U11290 (N_11290,N_9240,N_7342);
xnor U11291 (N_11291,N_6633,N_9925);
and U11292 (N_11292,N_6064,N_6027);
and U11293 (N_11293,N_9075,N_6680);
and U11294 (N_11294,N_9922,N_8906);
nand U11295 (N_11295,N_9959,N_9791);
nand U11296 (N_11296,N_5731,N_9694);
and U11297 (N_11297,N_7418,N_7539);
and U11298 (N_11298,N_9977,N_7552);
and U11299 (N_11299,N_5005,N_5847);
nand U11300 (N_11300,N_6332,N_7335);
nand U11301 (N_11301,N_8799,N_9687);
nand U11302 (N_11302,N_8765,N_9638);
xnor U11303 (N_11303,N_8072,N_8382);
and U11304 (N_11304,N_9451,N_9049);
nor U11305 (N_11305,N_8549,N_7080);
xor U11306 (N_11306,N_5535,N_8537);
and U11307 (N_11307,N_8309,N_5281);
and U11308 (N_11308,N_7716,N_7568);
nor U11309 (N_11309,N_8389,N_8571);
or U11310 (N_11310,N_6637,N_5872);
nand U11311 (N_11311,N_8433,N_6479);
and U11312 (N_11312,N_8408,N_6513);
nand U11313 (N_11313,N_6698,N_8296);
xor U11314 (N_11314,N_5637,N_6117);
and U11315 (N_11315,N_8579,N_5634);
nand U11316 (N_11316,N_6526,N_9442);
and U11317 (N_11317,N_5060,N_9885);
or U11318 (N_11318,N_9232,N_7677);
xor U11319 (N_11319,N_9713,N_9617);
nand U11320 (N_11320,N_9031,N_7164);
nand U11321 (N_11321,N_9833,N_5312);
and U11322 (N_11322,N_9572,N_9667);
or U11323 (N_11323,N_8396,N_9921);
nand U11324 (N_11324,N_9595,N_6464);
or U11325 (N_11325,N_5553,N_5335);
nor U11326 (N_11326,N_8340,N_6391);
or U11327 (N_11327,N_7447,N_5378);
nor U11328 (N_11328,N_9705,N_6714);
and U11329 (N_11329,N_6283,N_9727);
nor U11330 (N_11330,N_9072,N_8175);
or U11331 (N_11331,N_8544,N_7560);
nor U11332 (N_11332,N_8685,N_6456);
xor U11333 (N_11333,N_8651,N_9764);
xnor U11334 (N_11334,N_6220,N_6406);
or U11335 (N_11335,N_6018,N_9806);
nand U11336 (N_11336,N_6398,N_5951);
nand U11337 (N_11337,N_9254,N_6911);
and U11338 (N_11338,N_6641,N_8660);
or U11339 (N_11339,N_9525,N_7618);
nor U11340 (N_11340,N_5809,N_5329);
xnor U11341 (N_11341,N_7358,N_9904);
nand U11342 (N_11342,N_7003,N_6423);
nor U11343 (N_11343,N_9769,N_7112);
nand U11344 (N_11344,N_5475,N_8359);
nand U11345 (N_11345,N_9081,N_5918);
nand U11346 (N_11346,N_9434,N_7404);
nand U11347 (N_11347,N_9173,N_5153);
nor U11348 (N_11348,N_9192,N_6378);
and U11349 (N_11349,N_5521,N_8745);
nor U11350 (N_11350,N_5367,N_6520);
and U11351 (N_11351,N_8390,N_5302);
nand U11352 (N_11352,N_8801,N_8180);
or U11353 (N_11353,N_8438,N_8498);
or U11354 (N_11354,N_5080,N_9978);
nand U11355 (N_11355,N_9210,N_6703);
xnor U11356 (N_11356,N_8352,N_5646);
nor U11357 (N_11357,N_9856,N_8107);
or U11358 (N_11358,N_6208,N_8494);
nand U11359 (N_11359,N_5458,N_9736);
nand U11360 (N_11360,N_9062,N_8518);
or U11361 (N_11361,N_7459,N_9017);
nand U11362 (N_11362,N_8625,N_7523);
nand U11363 (N_11363,N_7103,N_6213);
and U11364 (N_11364,N_6662,N_9358);
or U11365 (N_11365,N_6009,N_9850);
or U11366 (N_11366,N_6091,N_5140);
nor U11367 (N_11367,N_9334,N_6643);
xnor U11368 (N_11368,N_9980,N_5869);
xnor U11369 (N_11369,N_5690,N_6249);
nand U11370 (N_11370,N_8250,N_5656);
nor U11371 (N_11371,N_6596,N_5680);
xnor U11372 (N_11372,N_6089,N_9701);
or U11373 (N_11373,N_7124,N_7007);
nor U11374 (N_11374,N_9316,N_5296);
nor U11375 (N_11375,N_8514,N_6773);
xor U11376 (N_11376,N_7528,N_9670);
nor U11377 (N_11377,N_5125,N_8272);
or U11378 (N_11378,N_5324,N_8697);
nand U11379 (N_11379,N_9034,N_9845);
xnor U11380 (N_11380,N_5170,N_6818);
xor U11381 (N_11381,N_5356,N_7510);
nand U11382 (N_11382,N_8879,N_8423);
nor U11383 (N_11383,N_5640,N_6996);
and U11384 (N_11384,N_6489,N_5825);
nand U11385 (N_11385,N_8302,N_8190);
nor U11386 (N_11386,N_8819,N_8266);
xor U11387 (N_11387,N_6809,N_6908);
xor U11388 (N_11388,N_9511,N_7525);
nand U11389 (N_11389,N_7663,N_7634);
xor U11390 (N_11390,N_7410,N_5216);
nor U11391 (N_11391,N_5072,N_8084);
nor U11392 (N_11392,N_7070,N_6828);
nor U11393 (N_11393,N_7805,N_5322);
nand U11394 (N_11394,N_6238,N_7344);
nor U11395 (N_11395,N_6803,N_5197);
xnor U11396 (N_11396,N_6050,N_9889);
or U11397 (N_11397,N_6419,N_8633);
xnor U11398 (N_11398,N_5993,N_5572);
or U11399 (N_11399,N_7334,N_8529);
nand U11400 (N_11400,N_7583,N_7206);
nor U11401 (N_11401,N_5489,N_5282);
and U11402 (N_11402,N_8944,N_8394);
nor U11403 (N_11403,N_5228,N_6710);
xnor U11404 (N_11404,N_9787,N_9048);
xor U11405 (N_11405,N_5560,N_6954);
xor U11406 (N_11406,N_8617,N_9543);
or U11407 (N_11407,N_7773,N_5615);
nor U11408 (N_11408,N_8323,N_9108);
nand U11409 (N_11409,N_8903,N_6673);
xnor U11410 (N_11410,N_8166,N_7729);
xor U11411 (N_11411,N_7218,N_7019);
nor U11412 (N_11412,N_7992,N_8674);
xnor U11413 (N_11413,N_8317,N_7783);
and U11414 (N_11414,N_9009,N_6901);
nand U11415 (N_11415,N_6942,N_8410);
nand U11416 (N_11416,N_8848,N_8249);
nor U11417 (N_11417,N_7545,N_6387);
nor U11418 (N_11418,N_9540,N_6784);
xor U11419 (N_11419,N_5341,N_8123);
and U11420 (N_11420,N_8720,N_8481);
and U11421 (N_11421,N_9319,N_7326);
or U11422 (N_11422,N_6721,N_6700);
or U11423 (N_11423,N_5058,N_7406);
xnor U11424 (N_11424,N_6783,N_8924);
nand U11425 (N_11425,N_5051,N_6883);
xnor U11426 (N_11426,N_7877,N_7246);
and U11427 (N_11427,N_8962,N_7586);
and U11428 (N_11428,N_9640,N_5798);
xor U11429 (N_11429,N_9418,N_6096);
nand U11430 (N_11430,N_5743,N_9615);
nand U11431 (N_11431,N_7551,N_7956);
nor U11432 (N_11432,N_6776,N_7444);
xor U11433 (N_11433,N_9517,N_7115);
nor U11434 (N_11434,N_6134,N_8162);
xnor U11435 (N_11435,N_6582,N_7629);
nand U11436 (N_11436,N_8473,N_8774);
or U11437 (N_11437,N_5575,N_9678);
nor U11438 (N_11438,N_6630,N_7708);
nor U11439 (N_11439,N_7243,N_9193);
and U11440 (N_11440,N_7939,N_8468);
nand U11441 (N_11441,N_9001,N_7758);
nor U11442 (N_11442,N_7662,N_6523);
nor U11443 (N_11443,N_9011,N_6279);
xor U11444 (N_11444,N_6219,N_9890);
nand U11445 (N_11445,N_6211,N_8583);
xor U11446 (N_11446,N_5410,N_7998);
nand U11447 (N_11447,N_9566,N_5380);
nor U11448 (N_11448,N_9433,N_7238);
nor U11449 (N_11449,N_7044,N_7697);
nor U11450 (N_11450,N_8193,N_5038);
xnor U11451 (N_11451,N_6689,N_7536);
nor U11452 (N_11452,N_8693,N_9911);
nor U11453 (N_11453,N_7224,N_6627);
and U11454 (N_11454,N_9786,N_7951);
and U11455 (N_11455,N_8008,N_9663);
xor U11456 (N_11456,N_7571,N_6963);
or U11457 (N_11457,N_5607,N_7349);
or U11458 (N_11458,N_7606,N_8562);
or U11459 (N_11459,N_5433,N_8912);
nand U11460 (N_11460,N_7934,N_9721);
nor U11461 (N_11461,N_5924,N_5502);
and U11462 (N_11462,N_8840,N_5467);
nor U11463 (N_11463,N_8065,N_5504);
nor U11464 (N_11464,N_9165,N_9383);
xor U11465 (N_11465,N_6471,N_9800);
nand U11466 (N_11466,N_9228,N_8030);
or U11467 (N_11467,N_6652,N_5873);
xor U11468 (N_11468,N_6917,N_5616);
nor U11469 (N_11469,N_9999,N_5705);
nor U11470 (N_11470,N_5821,N_9255);
and U11471 (N_11471,N_6877,N_8226);
or U11472 (N_11472,N_7608,N_9931);
xor U11473 (N_11473,N_9847,N_7484);
and U11474 (N_11474,N_9286,N_5444);
and U11475 (N_11475,N_5056,N_8450);
nor U11476 (N_11476,N_7015,N_9484);
nor U11477 (N_11477,N_8838,N_5714);
nand U11478 (N_11478,N_8478,N_9600);
xnor U11479 (N_11479,N_8222,N_5618);
and U11480 (N_11480,N_5461,N_9427);
nand U11481 (N_11481,N_7307,N_5514);
nand U11482 (N_11482,N_8975,N_7688);
nor U11483 (N_11483,N_8011,N_9079);
nand U11484 (N_11484,N_8768,N_6835);
and U11485 (N_11485,N_9652,N_8872);
nor U11486 (N_11486,N_9548,N_5422);
nor U11487 (N_11487,N_8385,N_8393);
xnor U11488 (N_11488,N_9261,N_8897);
nor U11489 (N_11489,N_6616,N_8137);
nor U11490 (N_11490,N_6590,N_9478);
and U11491 (N_11491,N_5384,N_8235);
or U11492 (N_11492,N_5619,N_6230);
and U11493 (N_11493,N_5396,N_6090);
nand U11494 (N_11494,N_9005,N_6960);
nor U11495 (N_11495,N_8803,N_8676);
xnor U11496 (N_11496,N_8636,N_6346);
xnor U11497 (N_11497,N_7674,N_7948);
or U11498 (N_11498,N_5474,N_5061);
nor U11499 (N_11499,N_5219,N_8240);
nand U11500 (N_11500,N_8210,N_6920);
nand U11501 (N_11501,N_6772,N_7062);
xnor U11502 (N_11502,N_9844,N_6048);
and U11503 (N_11503,N_5133,N_7610);
and U11504 (N_11504,N_9365,N_9288);
nand U11505 (N_11505,N_9635,N_5662);
and U11506 (N_11506,N_6647,N_6825);
and U11507 (N_11507,N_6525,N_5891);
xor U11508 (N_11508,N_9857,N_5790);
or U11509 (N_11509,N_6355,N_5577);
and U11510 (N_11510,N_6600,N_5091);
xnor U11511 (N_11511,N_5252,N_9702);
and U11512 (N_11512,N_9594,N_7419);
nand U11513 (N_11513,N_5725,N_8424);
nand U11514 (N_11514,N_6743,N_9838);
nand U11515 (N_11515,N_6383,N_9234);
or U11516 (N_11516,N_9854,N_6085);
and U11517 (N_11517,N_6654,N_7891);
and U11518 (N_11518,N_6974,N_8908);
or U11519 (N_11519,N_9450,N_6731);
nand U11520 (N_11520,N_5239,N_5141);
and U11521 (N_11521,N_5485,N_6335);
and U11522 (N_11522,N_8716,N_9003);
nand U11523 (N_11523,N_8236,N_5747);
xor U11524 (N_11524,N_7520,N_8846);
and U11525 (N_11525,N_7102,N_6250);
or U11526 (N_11526,N_5077,N_5287);
nor U11527 (N_11527,N_7969,N_8605);
xor U11528 (N_11528,N_6065,N_9371);
xor U11529 (N_11529,N_5912,N_8807);
xor U11530 (N_11530,N_7328,N_6836);
and U11531 (N_11531,N_6813,N_9283);
nand U11532 (N_11532,N_9395,N_7781);
xnor U11533 (N_11533,N_5645,N_6855);
nand U11534 (N_11534,N_5793,N_9519);
nand U11535 (N_11535,N_9760,N_8050);
or U11536 (N_11536,N_7616,N_8101);
and U11537 (N_11537,N_6418,N_6943);
nor U11538 (N_11538,N_9082,N_7757);
and U11539 (N_11539,N_9171,N_5007);
nor U11540 (N_11540,N_9599,N_5207);
xnor U11541 (N_11541,N_8907,N_5161);
nand U11542 (N_11542,N_8889,N_7469);
or U11543 (N_11543,N_5358,N_7607);
nor U11544 (N_11544,N_8322,N_8612);
nor U11545 (N_11545,N_6865,N_9775);
nand U11546 (N_11546,N_9016,N_8727);
and U11547 (N_11547,N_7486,N_6604);
xnor U11548 (N_11548,N_8017,N_9968);
nand U11549 (N_11549,N_9619,N_9413);
and U11550 (N_11550,N_9060,N_8839);
or U11551 (N_11551,N_7852,N_8372);
xnor U11552 (N_11552,N_7006,N_7867);
or U11553 (N_11553,N_9021,N_9090);
nand U11554 (N_11554,N_5230,N_9310);
and U11555 (N_11555,N_9521,N_9057);
xnor U11556 (N_11556,N_7488,N_5875);
or U11557 (N_11557,N_7766,N_5008);
and U11558 (N_11558,N_9118,N_8139);
and U11559 (N_11559,N_8961,N_9456);
and U11560 (N_11560,N_6297,N_6445);
xor U11561 (N_11561,N_6713,N_9393);
nand U11562 (N_11562,N_5819,N_9645);
xor U11563 (N_11563,N_5921,N_7187);
nor U11564 (N_11564,N_5057,N_5099);
nor U11565 (N_11565,N_6686,N_7840);
nor U11566 (N_11566,N_8426,N_6585);
or U11567 (N_11567,N_9604,N_8316);
or U11568 (N_11568,N_5675,N_6863);
or U11569 (N_11569,N_7739,N_7155);
or U11570 (N_11570,N_5839,N_7973);
xnor U11571 (N_11571,N_7258,N_7020);
nor U11572 (N_11572,N_6051,N_7057);
nand U11573 (N_11573,N_8366,N_9583);
xor U11574 (N_11574,N_7217,N_5049);
nor U11575 (N_11575,N_7979,N_5707);
nand U11576 (N_11576,N_9636,N_7229);
and U11577 (N_11577,N_9435,N_5693);
and U11578 (N_11578,N_5102,N_7822);
or U11579 (N_11579,N_6857,N_9512);
nand U11580 (N_11580,N_8918,N_8724);
and U11581 (N_11581,N_9321,N_8960);
xor U11582 (N_11582,N_9448,N_9204);
and U11583 (N_11583,N_7189,N_6845);
nor U11584 (N_11584,N_8106,N_7295);
nor U11585 (N_11585,N_6284,N_6944);
and U11586 (N_11586,N_8318,N_8667);
nand U11587 (N_11587,N_9725,N_9030);
xor U11588 (N_11588,N_7480,N_7085);
nor U11589 (N_11589,N_5330,N_8958);
and U11590 (N_11590,N_9536,N_8265);
xor U11591 (N_11591,N_5187,N_6165);
xor U11592 (N_11592,N_7449,N_8343);
nand U11593 (N_11593,N_7764,N_8849);
and U11594 (N_11594,N_8553,N_7446);
xnor U11595 (N_11595,N_6299,N_8164);
and U11596 (N_11596,N_9458,N_8082);
or U11597 (N_11597,N_6350,N_8288);
nand U11598 (N_11598,N_6948,N_8341);
nand U11599 (N_11599,N_6846,N_6754);
xor U11600 (N_11600,N_8945,N_9054);
xor U11601 (N_11601,N_5262,N_9068);
and U11602 (N_11602,N_7395,N_5272);
nor U11603 (N_11603,N_6889,N_8225);
nor U11604 (N_11604,N_6556,N_9715);
or U11605 (N_11605,N_6337,N_9527);
and U11606 (N_11606,N_8507,N_7895);
or U11607 (N_11607,N_5704,N_7862);
nor U11608 (N_11608,N_7094,N_5927);
or U11609 (N_11609,N_8603,N_7476);
nor U11610 (N_11610,N_5581,N_9937);
nand U11611 (N_11611,N_7869,N_6664);
nor U11612 (N_11612,N_9245,N_5299);
xor U11613 (N_11613,N_9064,N_9829);
nor U11614 (N_11614,N_8771,N_9526);
nand U11615 (N_11615,N_8258,N_8561);
nor U11616 (N_11616,N_5833,N_7664);
nand U11617 (N_11617,N_5834,N_9303);
nor U11618 (N_11618,N_9080,N_5248);
nand U11619 (N_11619,N_9287,N_5209);
nor U11620 (N_11620,N_9732,N_5027);
xor U11621 (N_11621,N_6127,N_7937);
nand U11622 (N_11622,N_5191,N_7451);
xor U11623 (N_11623,N_7661,N_5149);
and U11624 (N_11624,N_7337,N_6010);
nand U11625 (N_11625,N_9992,N_8830);
xor U11626 (N_11626,N_9043,N_5744);
nand U11627 (N_11627,N_7640,N_8357);
nand U11628 (N_11628,N_8543,N_8212);
and U11629 (N_11629,N_6531,N_5636);
nand U11630 (N_11630,N_5505,N_9465);
nor U11631 (N_11631,N_6542,N_5242);
nand U11632 (N_11632,N_7761,N_6054);
xor U11633 (N_11633,N_5968,N_6983);
xnor U11634 (N_11634,N_8955,N_9998);
nor U11635 (N_11635,N_7269,N_9646);
xnor U11636 (N_11636,N_9555,N_9737);
and U11637 (N_11637,N_7339,N_5387);
and U11638 (N_11638,N_5835,N_5249);
and U11639 (N_11639,N_8237,N_5144);
or U11640 (N_11640,N_6342,N_8687);
and U11641 (N_11641,N_7043,N_6796);
and U11642 (N_11642,N_6578,N_8029);
and U11643 (N_11643,N_8752,N_8422);
or U11644 (N_11644,N_7582,N_7615);
xor U11645 (N_11645,N_9348,N_9141);
nand U11646 (N_11646,N_6458,N_5154);
nor U11647 (N_11647,N_6063,N_5943);
and U11648 (N_11648,N_6276,N_8421);
and U11649 (N_11649,N_5767,N_8590);
nand U11650 (N_11650,N_5066,N_8827);
nor U11651 (N_11651,N_7635,N_6286);
xnor U11652 (N_11652,N_5439,N_8202);
or U11653 (N_11653,N_8865,N_6348);
nand U11654 (N_11654,N_5592,N_5868);
xnor U11655 (N_11655,N_9370,N_7416);
nand U11656 (N_11656,N_5438,N_7838);
and U11657 (N_11657,N_5755,N_7912);
and U11658 (N_11658,N_7620,N_9154);
xor U11659 (N_11659,N_6913,N_9814);
xnor U11660 (N_11660,N_6873,N_7704);
and U11661 (N_11661,N_5480,N_5766);
and U11662 (N_11662,N_8284,N_9945);
or U11663 (N_11663,N_7885,N_7077);
xor U11664 (N_11664,N_9241,N_8074);
or U11665 (N_11665,N_8776,N_8299);
xor U11666 (N_11666,N_9893,N_6060);
xnor U11667 (N_11667,N_9963,N_7240);
nor U11668 (N_11668,N_8835,N_9225);
nand U11669 (N_11669,N_8380,N_8970);
and U11670 (N_11670,N_5117,N_6062);
nor U11671 (N_11671,N_9771,N_9485);
or U11672 (N_11672,N_8998,N_9630);
or U11673 (N_11673,N_9719,N_7983);
nand U11674 (N_11674,N_5491,N_8585);
and U11675 (N_11675,N_6159,N_6319);
or U11676 (N_11676,N_9129,N_7846);
nor U11677 (N_11677,N_8334,N_8878);
nand U11678 (N_11678,N_6833,N_7863);
or U11679 (N_11679,N_6712,N_6422);
and U11680 (N_11680,N_5628,N_5611);
and U11681 (N_11681,N_6139,N_8335);
nand U11682 (N_11682,N_7134,N_8356);
or U11683 (N_11683,N_8387,N_9487);
xor U11684 (N_11684,N_8512,N_5025);
nor U11685 (N_11685,N_5067,N_9796);
nor U11686 (N_11686,N_9950,N_6039);
nor U11687 (N_11687,N_6273,N_8163);
nand U11688 (N_11688,N_9529,N_7505);
or U11689 (N_11689,N_7554,N_8403);
nor U11690 (N_11690,N_5204,N_7808);
and U11691 (N_11691,N_6516,N_8386);
nor U11692 (N_11692,N_9969,N_8006);
nand U11693 (N_11693,N_8709,N_6262);
nand U11694 (N_11694,N_5991,N_8987);
xor U11695 (N_11695,N_8172,N_5231);
nor U11696 (N_11696,N_9125,N_7403);
xnor U11697 (N_11697,N_9633,N_7017);
nand U11698 (N_11698,N_7769,N_9351);
or U11699 (N_11699,N_7540,N_5797);
xor U11700 (N_11700,N_7727,N_5668);
and U11701 (N_11701,N_6770,N_8015);
nand U11702 (N_11702,N_8041,N_6930);
or U11703 (N_11703,N_5172,N_5173);
xnor U11704 (N_11704,N_9562,N_6793);
xnor U11705 (N_11705,N_5554,N_6128);
and U11706 (N_11706,N_9780,N_9970);
nand U11707 (N_11707,N_7467,N_8055);
nand U11708 (N_11708,N_6404,N_6059);
nor U11709 (N_11709,N_9507,N_8843);
nor U11710 (N_11710,N_5403,N_9610);
xor U11711 (N_11711,N_7242,N_8269);
and U11712 (N_11712,N_7753,N_5269);
nor U11713 (N_11713,N_6478,N_5301);
and U11714 (N_11714,N_7658,N_7048);
or U11715 (N_11715,N_6549,N_9946);
and U11716 (N_11716,N_6860,N_6794);
nand U11717 (N_11717,N_6671,N_6915);
nand U11718 (N_11718,N_9305,N_8813);
nand U11719 (N_11719,N_6242,N_7241);
xnor U11720 (N_11720,N_8425,N_6303);
nand U11721 (N_11721,N_9565,N_5621);
xor U11722 (N_11722,N_9231,N_7463);
or U11723 (N_11723,N_9872,N_6243);
nor U11724 (N_11724,N_6439,N_6252);
nand U11725 (N_11725,N_9063,N_7556);
xnor U11726 (N_11726,N_9545,N_9447);
xor U11727 (N_11727,N_9813,N_8692);
or U11728 (N_11728,N_7435,N_9901);
nand U11729 (N_11729,N_7888,N_8653);
xnor U11730 (N_11730,N_9344,N_8260);
nand U11731 (N_11731,N_9948,N_6899);
and U11732 (N_11732,N_5941,N_8267);
nand U11733 (N_11733,N_7836,N_6269);
or U11734 (N_11734,N_7585,N_8851);
xnor U11735 (N_11735,N_6538,N_7646);
nor U11736 (N_11736,N_7911,N_6792);
nand U11737 (N_11737,N_9782,N_8402);
xor U11738 (N_11738,N_5856,N_9746);
nand U11739 (N_11739,N_6995,N_5454);
or U11740 (N_11740,N_9821,N_9590);
or U11741 (N_11741,N_7343,N_6839);
and U11742 (N_11742,N_7941,N_9278);
xor U11743 (N_11743,N_6421,N_7933);
nor U11744 (N_11744,N_6837,N_7910);
nor U11745 (N_11745,N_6517,N_6226);
nor U11746 (N_11746,N_5811,N_9537);
xor U11747 (N_11747,N_9586,N_5748);
and U11748 (N_11748,N_6571,N_5579);
or U11749 (N_11749,N_8069,N_5597);
nand U11750 (N_11750,N_9015,N_5585);
and U11751 (N_11751,N_5567,N_5687);
and U11752 (N_11752,N_9350,N_7420);
nand U11753 (N_11753,N_8160,N_5823);
and U11754 (N_11754,N_5107,N_5954);
xor U11755 (N_11755,N_5920,N_7431);
xnor U11756 (N_11756,N_9836,N_7929);
xnor U11757 (N_11757,N_6790,N_5074);
nand U11758 (N_11758,N_7266,N_6296);
nand U11759 (N_11759,N_6380,N_5904);
and U11760 (N_11760,N_7147,N_5390);
or U11761 (N_11761,N_7005,N_7388);
nand U11762 (N_11762,N_9988,N_8416);
and U11763 (N_11763,N_9809,N_7154);
or U11764 (N_11764,N_6052,N_6888);
and U11765 (N_11765,N_6021,N_6659);
xnor U11766 (N_11766,N_7316,N_6442);
nor U11767 (N_11767,N_6300,N_9518);
nor U11768 (N_11768,N_7676,N_5770);
and U11769 (N_11769,N_7148,N_5897);
and U11770 (N_11770,N_6417,N_6533);
and U11771 (N_11771,N_9459,N_8781);
xor U11772 (N_11772,N_7010,N_6007);
nor U11773 (N_11773,N_8310,N_8215);
or U11774 (N_11774,N_9273,N_8059);
nor U11775 (N_11775,N_8154,N_7747);
nor U11776 (N_11776,N_9953,N_9100);
and U11777 (N_11777,N_5788,N_8398);
xnor U11778 (N_11778,N_8465,N_9276);
and U11779 (N_11779,N_7202,N_5078);
xnor U11780 (N_11780,N_6724,N_6702);
and U11781 (N_11781,N_5389,N_6254);
and U11782 (N_11782,N_9312,N_7265);
xnor U11783 (N_11783,N_6670,N_6515);
or U11784 (N_11784,N_5487,N_7276);
nor U11785 (N_11785,N_8234,N_8920);
nand U11786 (N_11786,N_6751,N_9069);
or U11787 (N_11787,N_6446,N_6482);
xnor U11788 (N_11788,N_5894,N_5340);
xor U11789 (N_11789,N_6321,N_6737);
nand U11790 (N_11790,N_6475,N_5086);
and U11791 (N_11791,N_5383,N_8470);
nor U11792 (N_11792,N_6650,N_8723);
nand U11793 (N_11793,N_6867,N_5046);
and U11794 (N_11794,N_5490,N_7108);
nand U11795 (N_11795,N_7142,N_7823);
and U11796 (N_11796,N_7986,N_8598);
xnor U11797 (N_11797,N_9222,N_5880);
xnor U11798 (N_11798,N_9886,N_7089);
xor U11799 (N_11799,N_7179,N_7802);
nand U11800 (N_11800,N_6791,N_5919);
nor U11801 (N_11801,N_5889,N_5882);
nand U11802 (N_11802,N_6194,N_5870);
nor U11803 (N_11803,N_7401,N_7625);
xor U11804 (N_11804,N_7776,N_7171);
nor U11805 (N_11805,N_9758,N_5952);
nand U11806 (N_11806,N_7765,N_9891);
or U11807 (N_11807,N_5413,N_7542);
or U11808 (N_11808,N_6642,N_9848);
xnor U11809 (N_11809,N_7714,N_7436);
nor U11810 (N_11810,N_8596,N_6717);
xor U11811 (N_11811,N_6535,N_6399);
nor U11812 (N_11812,N_5174,N_6473);
nor U11813 (N_11813,N_7614,N_8714);
xor U11814 (N_11814,N_8869,N_8957);
and U11815 (N_11815,N_9422,N_5022);
nand U11816 (N_11816,N_5986,N_7325);
and U11817 (N_11817,N_8951,N_8221);
nand U11818 (N_11818,N_7740,N_8053);
nand U11819 (N_11819,N_6120,N_6133);
nor U11820 (N_11820,N_5781,N_8825);
nand U11821 (N_11821,N_7702,N_5805);
nand U11822 (N_11822,N_6692,N_9620);
nor U11823 (N_11823,N_5208,N_9135);
nor U11824 (N_11824,N_7515,N_6584);
nand U11825 (N_11825,N_9146,N_9585);
and U11826 (N_11826,N_9153,N_7113);
nor U11827 (N_11827,N_7390,N_8353);
and U11828 (N_11828,N_8294,N_6775);
or U11829 (N_11829,N_5115,N_6035);
xnor U11830 (N_11830,N_5867,N_5758);
nor U11831 (N_11831,N_9175,N_6008);
nand U11832 (N_11832,N_6022,N_6258);
and U11833 (N_11833,N_9306,N_9956);
xor U11834 (N_11834,N_5695,N_8672);
nand U11835 (N_11835,N_8141,N_5131);
nor U11836 (N_11836,N_6239,N_7173);
or U11837 (N_11837,N_6094,N_9693);
and U11838 (N_11838,N_8502,N_5229);
or U11839 (N_11839,N_9706,N_7996);
and U11840 (N_11840,N_6261,N_9853);
xor U11841 (N_11841,N_5808,N_6979);
nand U11842 (N_11842,N_5271,N_9087);
nand U11843 (N_11843,N_7138,N_7886);
and U11844 (N_11844,N_7711,N_5729);
nand U11845 (N_11845,N_8873,N_8189);
nand U11846 (N_11846,N_9169,N_5118);
xor U11847 (N_11847,N_9366,N_5083);
xnor U11848 (N_11848,N_5445,N_5244);
or U11849 (N_11849,N_9501,N_7427);
and U11850 (N_11850,N_5103,N_9855);
nand U11851 (N_11851,N_5602,N_9867);
and U11852 (N_11852,N_5215,N_8490);
nand U11853 (N_11853,N_9322,N_8377);
xnor U11854 (N_11854,N_5116,N_8138);
nor U11855 (N_11855,N_8530,N_8081);
or U11856 (N_11856,N_7169,N_5944);
or U11857 (N_11857,N_8611,N_8332);
and U11858 (N_11858,N_9095,N_7036);
nor U11859 (N_11859,N_8972,N_8177);
nand U11860 (N_11860,N_7482,N_8506);
nor U11861 (N_11861,N_7987,N_5734);
nor U11862 (N_11862,N_6171,N_8728);
nand U11863 (N_11863,N_7965,N_8668);
xor U11864 (N_11864,N_6033,N_6822);
nand U11865 (N_11865,N_6372,N_9659);
xnor U11866 (N_11866,N_7843,N_9318);
nand U11867 (N_11867,N_9463,N_9515);
or U11868 (N_11868,N_6151,N_8735);
xor U11869 (N_11869,N_6107,N_9785);
and U11870 (N_11870,N_8327,N_7915);
xnor U11871 (N_11871,N_6122,N_6745);
and U11872 (N_11872,N_8994,N_6200);
nor U11873 (N_11873,N_5990,N_5192);
nand U11874 (N_11874,N_6964,N_6448);
and U11875 (N_11875,N_6340,N_7092);
nor U11876 (N_11876,N_9623,N_6722);
and U11877 (N_11877,N_9831,N_9933);
and U11878 (N_11878,N_9770,N_6880);
nor U11879 (N_11879,N_8563,N_7695);
or U11880 (N_11880,N_7468,N_7434);
nand U11881 (N_11881,N_6352,N_7887);
nand U11882 (N_11882,N_5931,N_7405);
and U11883 (N_11883,N_5156,N_9582);
xor U11884 (N_11884,N_6769,N_6587);
xor U11885 (N_11885,N_7734,N_8634);
xnor U11886 (N_11886,N_8256,N_9270);
xor U11887 (N_11887,N_6403,N_5936);
xnor U11888 (N_11888,N_5601,N_8179);
nand U11889 (N_11889,N_9489,N_5092);
and U11890 (N_11890,N_8856,N_8696);
and U11891 (N_11891,N_7384,N_8483);
nor U11892 (N_11892,N_5896,N_9798);
nor U11893 (N_11893,N_8167,N_7690);
xor U11894 (N_11894,N_6270,N_5737);
nand U11895 (N_11895,N_5309,N_7936);
nor U11896 (N_11896,N_7516,N_8810);
nand U11897 (N_11897,N_6379,N_6470);
or U11898 (N_11898,N_6986,N_5971);
or U11899 (N_11899,N_7767,N_5582);
and U11900 (N_11900,N_8400,N_6132);
xnor U11901 (N_11901,N_8703,N_5590);
and U11902 (N_11902,N_8532,N_9681);
nand U11903 (N_11903,N_7340,N_9864);
nand U11904 (N_11904,N_5670,N_9291);
and U11905 (N_11905,N_5994,N_6683);
nand U11906 (N_11906,N_9264,N_5270);
xnor U11907 (N_11907,N_9675,N_9837);
xor U11908 (N_11908,N_6744,N_8515);
nor U11909 (N_11909,N_9074,N_8263);
or U11910 (N_11910,N_6693,N_6771);
and U11911 (N_11911,N_6188,N_8326);
xnor U11912 (N_11912,N_7140,N_6118);
and U11913 (N_11913,N_6480,N_7565);
or U11914 (N_11914,N_8795,N_7305);
and U11915 (N_11915,N_9452,N_5397);
or U11916 (N_11916,N_8983,N_5661);
nor U11917 (N_11917,N_7278,N_5469);
nor U11918 (N_11918,N_7192,N_9088);
and U11919 (N_11919,N_5040,N_5503);
and U11920 (N_11920,N_8348,N_9324);
xnor U11921 (N_11921,N_6746,N_5596);
nor U11922 (N_11922,N_9333,N_9275);
nor U11923 (N_11923,N_9035,N_8837);
nand U11924 (N_11924,N_9862,N_9588);
nor U11925 (N_11925,N_9219,N_6401);
or U11926 (N_11926,N_6240,N_8293);
nand U11927 (N_11927,N_7285,N_8208);
nor U11928 (N_11928,N_6534,N_8736);
nor U11929 (N_11929,N_6852,N_8246);
xnor U11930 (N_11930,N_5150,N_5814);
or U11931 (N_11931,N_9656,N_5499);
and U11932 (N_11932,N_8360,N_5225);
nor U11933 (N_11933,N_5063,N_9979);
xor U11934 (N_11934,N_6392,N_7550);
or U11935 (N_11935,N_9498,N_7549);
nand U11936 (N_11936,N_6937,N_5477);
xnor U11937 (N_11937,N_8631,N_9212);
xnor U11938 (N_11938,N_8109,N_5110);
and U11939 (N_11939,N_6228,N_6023);
xor U11940 (N_11940,N_5972,N_8601);
nand U11941 (N_11941,N_6317,N_8120);
and U11942 (N_11942,N_5155,N_5011);
and U11943 (N_11943,N_7443,N_7214);
nor U11944 (N_11944,N_9835,N_8999);
nor U11945 (N_11945,N_6201,N_7817);
or U11946 (N_11946,N_9119,N_5542);
xor U11947 (N_11947,N_9709,N_8466);
xnor U11948 (N_11948,N_8510,N_8460);
or U11949 (N_11949,N_6275,N_9748);
xnor U11950 (N_11950,N_5901,N_8113);
and U11951 (N_11951,N_5876,N_8591);
and U11952 (N_11952,N_5316,N_6088);
or U11953 (N_11953,N_9018,N_9185);
and U11954 (N_11954,N_9139,N_9739);
and U11955 (N_11955,N_5960,N_9269);
nor U11956 (N_11956,N_6102,N_9150);
nor U11957 (N_11957,N_7977,N_6099);
nor U11958 (N_11958,N_6137,N_6459);
nand U11959 (N_11959,N_9767,N_8793);
and U11960 (N_11960,N_5344,N_5221);
xor U11961 (N_11961,N_9439,N_7184);
and U11962 (N_11962,N_6718,N_6507);
or U11963 (N_11963,N_8071,N_5911);
xor U11964 (N_11964,N_6626,N_7558);
nor U11965 (N_11965,N_8949,N_7927);
and U11966 (N_11966,N_8682,N_9657);
or U11967 (N_11967,N_5459,N_6020);
or U11968 (N_11968,N_9851,N_7707);
or U11969 (N_11969,N_5128,N_7079);
nand U11970 (N_11970,N_5547,N_6789);
and U11971 (N_11971,N_7324,N_8509);
nand U11972 (N_11972,N_8158,N_7854);
nor U11973 (N_11973,N_5366,N_6197);
and U11974 (N_11974,N_9123,N_6265);
and U11975 (N_11975,N_5280,N_9382);
or U11976 (N_11976,N_7499,N_6851);
nand U11977 (N_11977,N_6527,N_5524);
nand U11978 (N_11978,N_5949,N_5745);
and U11979 (N_11979,N_9236,N_6613);
or U11980 (N_11980,N_6487,N_6113);
nor U11981 (N_11981,N_8704,N_8792);
or U11982 (N_11982,N_5420,N_6661);
xnor U11983 (N_11983,N_5457,N_6577);
xor U11984 (N_11984,N_6485,N_8934);
nor U11985 (N_11985,N_9446,N_6040);
nand U11986 (N_11986,N_9695,N_6938);
nor U11987 (N_11987,N_7703,N_6287);
nor U11988 (N_11988,N_6212,N_6389);
xor U11989 (N_11989,N_5275,N_9299);
nand U11990 (N_11990,N_9180,N_8063);
or U11991 (N_11991,N_5090,N_8003);
nand U11992 (N_11992,N_5720,N_9919);
nor U11993 (N_11993,N_5081,N_6076);
or U11994 (N_11994,N_7157,N_6695);
and U11995 (N_11995,N_6933,N_6881);
xor U11996 (N_11996,N_7178,N_8242);
or U11997 (N_11997,N_7534,N_8491);
or U11998 (N_11998,N_5134,N_7315);
nand U11999 (N_11999,N_8251,N_7454);
or U12000 (N_12000,N_8100,N_8375);
xnor U12001 (N_12001,N_8146,N_5437);
nor U12002 (N_12002,N_6206,N_8440);
or U12003 (N_12003,N_9500,N_9917);
nand U12004 (N_12004,N_5712,N_5009);
and U12005 (N_12005,N_5473,N_9605);
nand U12006 (N_12006,N_5126,N_9010);
and U12007 (N_12007,N_7478,N_8600);
nor U12008 (N_12008,N_9607,N_5147);
xor U12009 (N_12009,N_5014,N_5778);
xnor U12010 (N_12010,N_6175,N_7018);
xnor U12011 (N_12011,N_5609,N_8091);
nand U12012 (N_12012,N_7483,N_9927);
nand U12013 (N_12013,N_5976,N_5979);
nand U12014 (N_12014,N_6079,N_6463);
and U12015 (N_12015,N_7396,N_5604);
xor U12016 (N_12016,N_6161,N_9714);
nor U12017 (N_12017,N_9381,N_5751);
or U12018 (N_12018,N_5998,N_9596);
and U12019 (N_12019,N_5421,N_9603);
and U12020 (N_12020,N_9332,N_5669);
nand U12021 (N_12021,N_6402,N_8985);
nand U12022 (N_12022,N_5357,N_7042);
and U12023 (N_12023,N_7785,N_8919);
or U12024 (N_12024,N_5497,N_6222);
and U12025 (N_12025,N_7050,N_7678);
and U12026 (N_12026,N_7670,N_6434);
xnor U12027 (N_12027,N_8749,N_6900);
xor U12028 (N_12028,N_8766,N_7966);
or U12029 (N_12029,N_6467,N_8973);
or U12030 (N_12030,N_6566,N_9865);
nand U12031 (N_12031,N_9115,N_7633);
nor U12032 (N_12032,N_9934,N_8980);
nor U12033 (N_12033,N_5934,N_7135);
and U12034 (N_12034,N_8659,N_6629);
and U12035 (N_12035,N_5227,N_6898);
xor U12036 (N_12036,N_7861,N_9538);
nand U12037 (N_12037,N_8241,N_6764);
and U12038 (N_12038,N_7028,N_9140);
nand U12039 (N_12039,N_7693,N_8564);
nor U12040 (N_12040,N_5531,N_7914);
nand U12041 (N_12041,N_5260,N_7738);
and U12042 (N_12042,N_6593,N_5291);
or U12043 (N_12043,N_6924,N_9110);
xor U12044 (N_12044,N_9412,N_9730);
nor U12045 (N_12045,N_7548,N_7255);
nor U12046 (N_12046,N_6756,N_7932);
nand U12047 (N_12047,N_7675,N_5666);
and U12048 (N_12048,N_6786,N_9920);
xnor U12049 (N_12049,N_8336,N_8655);
xnor U12050 (N_12050,N_9776,N_6098);
xnor U12051 (N_12051,N_6946,N_5178);
nand U12052 (N_12052,N_8550,N_9296);
xor U12053 (N_12053,N_6685,N_7512);
nor U12054 (N_12054,N_6278,N_5018);
or U12055 (N_12055,N_6848,N_6338);
nand U12056 (N_12056,N_6886,N_7710);
xnor U12057 (N_12057,N_9906,N_7424);
and U12058 (N_12058,N_6965,N_9038);
and U12059 (N_12059,N_5644,N_9668);
and U12060 (N_12060,N_7201,N_9522);
xor U12061 (N_12061,N_5975,N_9524);
nand U12062 (N_12062,N_6801,N_5452);
nor U12063 (N_12063,N_9469,N_6874);
and U12064 (N_12064,N_8159,N_8126);
and U12065 (N_12065,N_5050,N_7632);
or U12066 (N_12066,N_7502,N_7374);
or U12067 (N_12067,N_9223,N_8432);
nor U12068 (N_12068,N_8315,N_8639);
or U12069 (N_12069,N_6231,N_6519);
xor U12070 (N_12070,N_7254,N_8662);
or U12071 (N_12071,N_9752,N_6734);
nand U12072 (N_12072,N_7209,N_9302);
or U12073 (N_12073,N_5129,N_6858);
xor U12074 (N_12074,N_8764,N_5319);
nor U12075 (N_12075,N_7770,N_8096);
and U12076 (N_12076,N_7975,N_7314);
or U12077 (N_12077,N_5430,N_7804);
or U12078 (N_12078,N_6199,N_7290);
and U12079 (N_12079,N_8794,N_5838);
nor U12080 (N_12080,N_5836,N_9428);
or U12081 (N_12081,N_6690,N_7819);
xor U12082 (N_12082,N_8582,N_5730);
or U12083 (N_12083,N_7059,N_8019);
nor U12084 (N_12084,N_9674,N_8741);
xor U12085 (N_12085,N_5785,N_7354);
nor U12086 (N_12086,N_5326,N_5846);
xor U12087 (N_12087,N_8976,N_8531);
or U12088 (N_12088,N_5708,N_9449);
and U12089 (N_12089,N_5691,N_5762);
and U12090 (N_12090,N_6741,N_9944);
nor U12091 (N_12091,N_9602,N_6336);
and U12092 (N_12092,N_6682,N_6904);
nor U12093 (N_12093,N_8185,N_7665);
or U12094 (N_12094,N_9020,N_5559);
and U12095 (N_12095,N_5143,N_9355);
or U12096 (N_12096,N_6766,N_8613);
and U12097 (N_12097,N_7132,N_7972);
or U12098 (N_12098,N_7561,N_6716);
xnor U12099 (N_12099,N_7500,N_9729);
xor U12100 (N_12100,N_7098,N_8679);
and U12101 (N_12101,N_7622,N_6579);
nand U12102 (N_12102,N_5238,N_9840);
nand U12103 (N_12103,N_9990,N_6357);
nand U12104 (N_12104,N_7014,N_7810);
xor U12105 (N_12105,N_7445,N_6912);
and U12106 (N_12106,N_6931,N_7573);
nor U12107 (N_12107,N_9547,N_7312);
nor U12108 (N_12108,N_8581,N_5600);
and U12109 (N_12109,N_8068,N_9492);
nand U12110 (N_12110,N_9717,N_7252);
xnor U12111 (N_12111,N_9421,N_7066);
and U12112 (N_12112,N_8358,N_8750);
nor U12113 (N_12113,N_5573,N_9441);
nand U12114 (N_12114,N_8572,N_7522);
xor U12115 (N_12115,N_6450,N_7402);
nor U12116 (N_12116,N_7350,N_5194);
nand U12117 (N_12117,N_9086,N_5036);
nor U12118 (N_12118,N_9055,N_9817);
and U12119 (N_12119,N_5750,N_9149);
and U12120 (N_12120,N_5423,N_9429);
xnor U12121 (N_12121,N_9226,N_6304);
nand U12122 (N_12122,N_5218,N_6145);
or U12123 (N_12123,N_5689,N_5711);
nor U12124 (N_12124,N_7535,N_7842);
xnor U12125 (N_12125,N_8039,N_9673);
xnor U12126 (N_12126,N_9745,N_7666);
nand U12127 (N_12127,N_5715,N_6677);
nand U12128 (N_12128,N_7870,N_9897);
nand U12129 (N_12129,N_8268,N_6004);
or U12130 (N_12130,N_6148,N_8116);
nand U12131 (N_12131,N_7090,N_9718);
or U12132 (N_12132,N_8829,N_7371);
or U12133 (N_12133,N_8519,N_7004);
and U12134 (N_12134,N_6388,N_5752);
nor U12135 (N_12135,N_5950,N_8777);
or U12136 (N_12136,N_8898,N_6777);
xor U12137 (N_12137,N_8418,N_9552);
nor U12138 (N_12138,N_9624,N_6333);
nand U12139 (N_12139,N_5177,N_9416);
or U12140 (N_12140,N_9686,N_5247);
xnor U12141 (N_12141,N_5700,N_6707);
and U12142 (N_12142,N_6247,N_6636);
and U12143 (N_12143,N_5211,N_6147);
xor U12144 (N_12144,N_5294,N_9846);
or U12145 (N_12145,N_7639,N_7651);
xnor U12146 (N_12146,N_8511,N_6000);
nand U12147 (N_12147,N_9513,N_5784);
nand U12148 (N_12148,N_6840,N_5483);
nor U12149 (N_12149,N_5965,N_7045);
and U12150 (N_12150,N_7967,N_6071);
nor U12151 (N_12151,N_7858,N_5414);
xor U12152 (N_12152,N_5053,N_5113);
and U12153 (N_12153,N_7489,N_8239);
nand U12154 (N_12154,N_7352,N_6967);
nor U12155 (N_12155,N_9597,N_6861);
xnor U12156 (N_12156,N_7903,N_7795);
and U12157 (N_12157,N_7803,N_6047);
nor U12158 (N_12158,N_5205,N_8964);
nor U12159 (N_12159,N_8363,N_9902);
nand U12160 (N_12160,N_5860,N_7650);
nor U12161 (N_12161,N_7359,N_7439);
nand U12162 (N_12162,N_9938,N_5685);
and U12163 (N_12163,N_9239,N_9581);
nor U12164 (N_12164,N_9094,N_7347);
or U12165 (N_12165,N_6362,N_6263);
nor U12166 (N_12166,N_9174,N_6359);
xor U12167 (N_12167,N_5635,N_9622);
or U12168 (N_12168,N_5373,N_6291);
and U12169 (N_12169,N_9142,N_8028);
xor U12170 (N_12170,N_8881,N_6506);
xor U12171 (N_12171,N_7541,N_8997);
and U12172 (N_12172,N_5824,N_8747);
nand U12173 (N_12173,N_6174,N_7317);
nor U12174 (N_12174,N_8673,N_6970);
xor U12175 (N_12175,N_7283,N_8595);
and U12176 (N_12176,N_7980,N_6496);
nor U12177 (N_12177,N_5512,N_7293);
xnor U12178 (N_12178,N_8298,N_9789);
nor U12179 (N_12179,N_5903,N_9126);
and U12180 (N_12180,N_9375,N_6617);
and U12181 (N_12181,N_8487,N_5455);
nand U12182 (N_12182,N_7107,N_6410);
or U12183 (N_12183,N_9013,N_5425);
or U12184 (N_12184,N_6583,N_7093);
and U12185 (N_12185,N_8560,N_6530);
xor U12186 (N_12186,N_7587,N_8002);
and U12187 (N_12187,N_8430,N_7475);
or U12188 (N_12188,N_5032,N_6621);
and U12189 (N_12189,N_5132,N_5059);
xnor U12190 (N_12190,N_6330,N_9573);
nand U12191 (N_12191,N_6656,N_8092);
xor U12192 (N_12192,N_6305,N_8748);
or U12193 (N_12193,N_7306,N_5222);
nor U12194 (N_12194,N_9976,N_8853);
nor U12195 (N_12195,N_6939,N_7845);
nand U12196 (N_12196,N_9483,N_6740);
nor U12197 (N_12197,N_8178,N_7379);
nor U12198 (N_12198,N_8196,N_6030);
nor U12199 (N_12199,N_7733,N_5509);
or U12200 (N_12200,N_8909,N_6518);
nor U12201 (N_12201,N_9680,N_5874);
nand U12202 (N_12202,N_8122,N_8320);
and U12203 (N_12203,N_8780,N_6750);
and U12204 (N_12204,N_9723,N_7874);
xnor U12205 (N_12205,N_7508,N_8496);
nand U12206 (N_12206,N_7497,N_7687);
xnor U12207 (N_12207,N_8324,N_6548);
nor U12208 (N_12208,N_8648,N_9589);
xor U12209 (N_12209,N_9271,N_5574);
nand U12210 (N_12210,N_5243,N_8451);
and U12211 (N_12211,N_5769,N_6437);
nand U12212 (N_12212,N_7487,N_8188);
or U12213 (N_12213,N_5183,N_9295);
or U12214 (N_12214,N_7303,N_7239);
nor U12215 (N_12215,N_7498,N_6293);
or U12216 (N_12216,N_8690,N_9628);
and U12217 (N_12217,N_5523,N_5105);
nand U12218 (N_12218,N_8147,N_7234);
or U12219 (N_12219,N_8832,N_5583);
and U12220 (N_12220,N_9749,N_6363);
and U12221 (N_12221,N_7720,N_6156);
nand U12222 (N_12222,N_9812,N_5023);
xnor U12223 (N_12223,N_6366,N_7680);
and U12224 (N_12224,N_8274,N_5106);
nor U12225 (N_12225,N_9750,N_6503);
nand U12226 (N_12226,N_9438,N_6807);
nor U12227 (N_12227,N_5517,N_5586);
or U12228 (N_12228,N_7513,N_8034);
or U12229 (N_12229,N_6569,N_5486);
or U12230 (N_12230,N_9121,N_6494);
nor U12231 (N_12231,N_5400,N_6461);
nand U12232 (N_12232,N_5807,N_9606);
nor U12233 (N_12233,N_6381,N_7440);
nor U12234 (N_12234,N_6657,N_6182);
and U12235 (N_12235,N_8786,N_5780);
xnor U12236 (N_12236,N_9329,N_6216);
or U12237 (N_12237,N_8680,N_6129);
and U12238 (N_12238,N_5983,N_9341);
or U12239 (N_12239,N_6195,N_6648);
nand U12240 (N_12240,N_6864,N_7398);
xnor U12241 (N_12241,N_9535,N_6256);
nor U12242 (N_12242,N_5350,N_8330);
nand U12243 (N_12243,N_6034,N_9058);
xor U12244 (N_12244,N_6361,N_5369);
nor U12245 (N_12245,N_8584,N_8938);
or U12246 (N_12246,N_8121,N_6573);
and U12247 (N_12247,N_6989,N_7600);
nand U12248 (N_12248,N_8913,N_7146);
xor U12249 (N_12249,N_7681,N_9914);
xnor U12250 (N_12250,N_7605,N_5576);
or U12251 (N_12251,N_8647,N_7872);
and U12252 (N_12252,N_5558,N_5768);
nand U12253 (N_12253,N_7268,N_9697);
nor U12254 (N_12254,N_8599,N_6687);
xor U12255 (N_12255,N_9556,N_7222);
and U12256 (N_12256,N_6536,N_7953);
or U12257 (N_12257,N_7399,N_7260);
or U12258 (N_12258,N_8480,N_5333);
nand U12259 (N_12259,N_9491,N_5555);
nor U12260 (N_12260,N_5962,N_7149);
nor U12261 (N_12261,N_6011,N_8415);
nor U12262 (N_12262,N_8199,N_6655);
nand U12263 (N_12263,N_8893,N_6823);
nor U12264 (N_12264,N_9882,N_5320);
nor U12265 (N_12265,N_9037,N_7273);
xnor U12266 (N_12266,N_5388,N_9690);
nand U12267 (N_12267,N_9077,N_9849);
and U12268 (N_12268,N_6580,N_7002);
xnor U12269 (N_12269,N_9574,N_7011);
xnor U12270 (N_12270,N_8427,N_7683);
nor U12271 (N_12271,N_5447,N_7812);
and U12272 (N_12272,N_6561,N_6509);
xor U12273 (N_12273,N_5311,N_7988);
nor U12274 (N_12274,N_7223,N_9502);
xnor U12275 (N_12275,N_8645,N_9546);
nor U12276 (N_12276,N_9377,N_6097);
nor U12277 (N_12277,N_9682,N_7698);
or U12278 (N_12278,N_8331,N_5386);
nor U12279 (N_12279,N_9047,N_7423);
nor U12280 (N_12280,N_6510,N_6343);
or U12281 (N_12281,N_8731,N_6735);
nor U12282 (N_12282,N_5738,N_7389);
nor U12283 (N_12283,N_7353,N_6204);
xnor U12284 (N_12284,N_7196,N_6420);
nor U12285 (N_12285,N_7580,N_9460);
xor U12286 (N_12286,N_8686,N_9877);
nor U12287 (N_12287,N_8992,N_7176);
xnor U12288 (N_12288,N_5479,N_7166);
nand U12289 (N_12289,N_6925,N_6961);
or U12290 (N_12290,N_8597,N_6160);
and U12291 (N_12291,N_7685,N_9731);
xnor U12292 (N_12292,N_7866,N_8522);
xor U12293 (N_12293,N_7294,N_6875);
nor U12294 (N_12294,N_8986,N_5710);
or U12295 (N_12295,N_9820,N_8996);
nor U12296 (N_12296,N_9989,N_8104);
and U12297 (N_12297,N_7837,N_5760);
or U12298 (N_12298,N_9793,N_8993);
xor U12299 (N_12299,N_7058,N_5654);
or U12300 (N_12300,N_8399,N_6455);
nand U12301 (N_12301,N_7466,N_6811);
and U12302 (N_12302,N_7706,N_6757);
and U12303 (N_12303,N_6214,N_6586);
or U12304 (N_12304,N_6013,N_7302);
xnor U12305 (N_12305,N_5800,N_5332);
or U12306 (N_12306,N_9621,N_9671);
xnor U12307 (N_12307,N_9679,N_9195);
or U12308 (N_12308,N_5765,N_6271);
nand U12309 (N_12309,N_7492,N_6691);
and U12310 (N_12310,N_5771,N_5955);
or U12311 (N_12311,N_5563,N_6802);
or U12312 (N_12312,N_9168,N_5460);
xnor U12313 (N_12313,N_9898,N_6066);
nand U12314 (N_12314,N_6856,N_8821);
nand U12315 (N_12315,N_9804,N_5650);
nor U12316 (N_12316,N_7365,N_9215);
xor U12317 (N_12317,N_7120,N_5251);
nand U12318 (N_12318,N_7655,N_9227);
nor U12319 (N_12319,N_5265,N_6615);
xor U12320 (N_12320,N_8984,N_9962);
or U12321 (N_12321,N_8405,N_8746);
and U12322 (N_12322,N_9691,N_9196);
nand U12323 (N_12323,N_6570,N_5001);
and U12324 (N_12324,N_5069,N_7021);
or U12325 (N_12325,N_9966,N_8216);
xor U12326 (N_12326,N_7751,N_5796);
xnor U12327 (N_12327,N_5021,N_8243);
and U12328 (N_12328,N_6234,N_9779);
and U12329 (N_12329,N_9768,N_5158);
nand U12330 (N_12330,N_8989,N_6376);
and U12331 (N_12331,N_7603,N_8079);
nor U12332 (N_12332,N_9997,N_6870);
nor U12333 (N_12333,N_5945,N_6605);
and U12334 (N_12334,N_8252,N_8025);
xor U12335 (N_12335,N_7871,N_8862);
xor U12336 (N_12336,N_5179,N_8954);
or U12337 (N_12337,N_7868,N_6492);
nand U12338 (N_12338,N_6511,N_9093);
or U12339 (N_12339,N_6440,N_7626);
nor U12340 (N_12340,N_7659,N_6646);
nor U12341 (N_12341,N_7922,N_7656);
xnor U12342 (N_12342,N_7111,N_9419);
or U12343 (N_12343,N_9326,N_5822);
nand U12344 (N_12344,N_7602,N_5857);
nand U12345 (N_12345,N_7824,N_6468);
nor U12346 (N_12346,N_6619,N_8814);
xor U12347 (N_12347,N_6952,N_6157);
nor U12348 (N_12348,N_7280,N_5331);
nand U12349 (N_12349,N_9744,N_9249);
nor U12350 (N_12350,N_8876,N_8574);
xor U12351 (N_12351,N_8501,N_8446);
xnor U12352 (N_12352,N_8203,N_5973);
xnor U12353 (N_12353,N_8886,N_7363);
nand U12354 (N_12354,N_8184,N_7237);
nor U12355 (N_12355,N_6895,N_5764);
or U12356 (N_12356,N_8671,N_6428);
nand U12357 (N_12357,N_7220,N_7026);
or U12358 (N_12358,N_9664,N_7170);
and U12359 (N_12359,N_6377,N_8505);
or U12360 (N_12360,N_9207,N_8090);
nor U12361 (N_12361,N_7850,N_7591);
xor U12362 (N_12362,N_6565,N_8831);
nor U12363 (N_12363,N_7075,N_5658);
or U12364 (N_12364,N_9763,N_9444);
and U12365 (N_12365,N_9479,N_6277);
xnor U12366 (N_12366,N_7493,N_6005);
nor U12367 (N_12367,N_5595,N_5146);
and U12368 (N_12368,N_9722,N_7038);
nor U12369 (N_12369,N_5076,N_7913);
or U12370 (N_12370,N_7907,N_5787);
and U12371 (N_12371,N_8866,N_5321);
and U12372 (N_12372,N_9221,N_5052);
or U12373 (N_12373,N_5892,N_5985);
nor U12374 (N_12374,N_7198,N_6962);
or U12375 (N_12375,N_8447,N_8860);
nand U12376 (N_12376,N_5703,N_5883);
nand U12377 (N_12377,N_7699,N_8695);
or U12378 (N_12378,N_9252,N_5910);
and U12379 (N_12379,N_7366,N_8610);
xnor U12380 (N_12380,N_7331,N_8559);
nor U12381 (N_12381,N_6397,N_6196);
nor U12382 (N_12382,N_6628,N_6144);
nand U12383 (N_12383,N_8229,N_5175);
or U12384 (N_12384,N_8675,N_6711);
and U12385 (N_12385,N_9981,N_5392);
nand U12386 (N_12386,N_6416,N_6267);
or U12387 (N_12387,N_7806,N_5786);
nand U12388 (N_12388,N_9815,N_9059);
nor U12389 (N_12389,N_6057,N_8369);
and U12390 (N_12390,N_7909,N_8626);
or U12391 (N_12391,N_9164,N_8575);
and U12392 (N_12392,N_7882,N_5306);
or U12393 (N_12393,N_5783,N_6982);
or U12394 (N_12394,N_5257,N_9564);
nand U12395 (N_12395,N_7376,N_5899);
nor U12396 (N_12396,N_5476,N_9368);
nand U12397 (N_12397,N_9754,N_6730);
and U12398 (N_12398,N_7322,N_7161);
nand U12399 (N_12399,N_8444,N_8988);
nand U12400 (N_12400,N_5967,N_6281);
or U12401 (N_12401,N_9122,N_8566);
or U12402 (N_12402,N_5841,N_9871);
and U12403 (N_12403,N_8966,N_8950);
and U12404 (N_12404,N_6890,N_7272);
xor U12405 (N_12405,N_5606,N_5361);
and U12406 (N_12406,N_6217,N_5929);
or U12407 (N_12407,N_7369,N_7735);
xnor U12408 (N_12408,N_6411,N_8066);
or U12409 (N_12409,N_6466,N_5121);
and U12410 (N_12410,N_8884,N_8169);
and U12411 (N_12411,N_9186,N_6314);
xor U12412 (N_12412,N_9496,N_7814);
xnor U12413 (N_12413,N_7296,N_5948);
or U12414 (N_12414,N_9811,N_6353);
or U12415 (N_12415,N_6755,N_8520);
nand U12416 (N_12416,N_7207,N_7117);
or U12417 (N_12417,N_7174,N_7648);
nand U12418 (N_12418,N_8785,N_7414);
and U12419 (N_12419,N_5293,N_5959);
and U12420 (N_12420,N_8044,N_6876);
or U12421 (N_12421,N_9683,N_5885);
nand U12422 (N_12422,N_6334,N_5907);
nor U12423 (N_12423,N_6610,N_7619);
xnor U12424 (N_12424,N_6785,N_5701);
nand U12425 (N_12425,N_7430,N_7524);
and U12426 (N_12426,N_9783,N_9328);
nor U12427 (N_12427,N_5665,N_7461);
and U12428 (N_12428,N_9148,N_8740);
nand U12429 (N_12429,N_5212,N_6665);
xnor U12430 (N_12430,N_7537,N_7873);
and U12431 (N_12431,N_7068,N_8286);
and U12432 (N_12432,N_5947,N_9506);
and U12433 (N_12433,N_8552,N_6667);
or U12434 (N_12434,N_8707,N_7095);
nand U12435 (N_12435,N_5404,N_5266);
or U12436 (N_12436,N_8351,N_5859);
and U12437 (N_12437,N_7345,N_9044);
or U12438 (N_12438,N_8623,N_6631);
and U12439 (N_12439,N_6893,N_8023);
or U12440 (N_12440,N_5774,N_9397);
or U12441 (N_12441,N_6906,N_5434);
xor U12442 (N_12442,N_8948,N_6725);
or U12443 (N_12443,N_6824,N_7978);
nor U12444 (N_12444,N_6266,N_5842);
nand U12445 (N_12445,N_5171,N_9408);
and U12446 (N_12446,N_7257,N_7949);
xnor U12447 (N_12447,N_8257,N_6998);
nand U12448 (N_12448,N_9098,N_6460);
xnor U12449 (N_12449,N_5649,N_9304);
and U12450 (N_12450,N_5385,N_9915);
nand U12451 (N_12451,N_6762,N_5017);
and U12452 (N_12452,N_8991,N_8923);
nor U12453 (N_12453,N_9083,N_6176);
nor U12454 (N_12454,N_5054,N_6950);
or U12455 (N_12455,N_8539,N_6126);
nor U12456 (N_12456,N_6289,N_9482);
xnor U12457 (N_12457,N_9477,N_6241);
xor U12458 (N_12458,N_6929,N_6551);
and U12459 (N_12459,N_8098,N_5881);
xnor U12460 (N_12460,N_9238,N_9753);
nor U12461 (N_12461,N_9471,N_5515);
or U12462 (N_12462,N_5189,N_8035);
and U12463 (N_12463,N_8108,N_7637);
xor U12464 (N_12464,N_6087,N_8683);
and U12465 (N_12465,N_6597,N_8007);
nor U12466 (N_12466,N_6624,N_7323);
or U12467 (N_12467,N_7660,N_6644);
nor U12468 (N_12468,N_6736,N_8397);
nor U12469 (N_12469,N_5709,N_6067);
xor U12470 (N_12470,N_7976,N_7078);
or U12471 (N_12471,N_6606,N_9895);
xnor U12472 (N_12472,N_8370,N_8627);
xnor U12473 (N_12473,N_5978,N_8646);
or U12474 (N_12474,N_9912,N_7311);
and U12475 (N_12475,N_8796,N_7338);
and U12476 (N_12476,N_7531,N_7833);
nor U12477 (N_12477,N_9584,N_5530);
xor U12478 (N_12478,N_5295,N_7830);
or U12479 (N_12479,N_6795,N_5127);
nand U12480 (N_12480,N_6601,N_8018);
or U12481 (N_12481,N_5276,N_8085);
or U12482 (N_12482,N_6985,N_5688);
and U12483 (N_12483,N_8891,N_6447);
nor U12484 (N_12484,N_8527,N_7778);
or U12485 (N_12485,N_7813,N_6192);
or U12486 (N_12486,N_7593,N_6999);
xnor U12487 (N_12487,N_5193,N_9955);
or U12488 (N_12488,N_8244,N_7712);
nor U12489 (N_12489,N_8804,N_5681);
or U12490 (N_12490,N_7609,N_8726);
or U12491 (N_12491,N_9343,N_8805);
xnor U12492 (N_12492,N_9401,N_6162);
or U12493 (N_12493,N_8311,N_6941);
nor U12494 (N_12494,N_7853,N_8542);
nand U12495 (N_12495,N_5343,N_9216);
nand U12496 (N_12496,N_7168,N_8378);
nor U12497 (N_12497,N_6532,N_9317);
xor U12498 (N_12498,N_8283,N_9842);
or U12499 (N_12499,N_9028,N_8738);
nand U12500 (N_12500,N_7784,N_6317);
xor U12501 (N_12501,N_6665,N_9760);
xnor U12502 (N_12502,N_5827,N_7622);
or U12503 (N_12503,N_6552,N_5631);
nor U12504 (N_12504,N_6227,N_7681);
nand U12505 (N_12505,N_7487,N_9633);
and U12506 (N_12506,N_5046,N_7491);
and U12507 (N_12507,N_5705,N_6841);
nor U12508 (N_12508,N_6806,N_8153);
and U12509 (N_12509,N_7074,N_9536);
xor U12510 (N_12510,N_9582,N_5717);
nand U12511 (N_12511,N_7362,N_8507);
nand U12512 (N_12512,N_8769,N_6491);
and U12513 (N_12513,N_5625,N_8097);
xnor U12514 (N_12514,N_8009,N_9926);
and U12515 (N_12515,N_6151,N_7344);
or U12516 (N_12516,N_9430,N_9554);
xor U12517 (N_12517,N_8550,N_6704);
and U12518 (N_12518,N_7534,N_7412);
nand U12519 (N_12519,N_8707,N_7767);
or U12520 (N_12520,N_6924,N_9258);
or U12521 (N_12521,N_8176,N_6109);
nor U12522 (N_12522,N_5592,N_5290);
and U12523 (N_12523,N_8091,N_9038);
and U12524 (N_12524,N_9883,N_7089);
and U12525 (N_12525,N_7332,N_8359);
or U12526 (N_12526,N_5432,N_7277);
xnor U12527 (N_12527,N_9793,N_9033);
nor U12528 (N_12528,N_9977,N_6647);
nand U12529 (N_12529,N_6384,N_9765);
xor U12530 (N_12530,N_5007,N_8811);
and U12531 (N_12531,N_5070,N_9144);
and U12532 (N_12532,N_8406,N_9491);
xor U12533 (N_12533,N_9170,N_9357);
nor U12534 (N_12534,N_5343,N_6166);
nand U12535 (N_12535,N_9328,N_5595);
nand U12536 (N_12536,N_5133,N_7575);
xnor U12537 (N_12537,N_8225,N_7901);
and U12538 (N_12538,N_6090,N_5397);
xor U12539 (N_12539,N_9150,N_5996);
nor U12540 (N_12540,N_7043,N_9452);
nor U12541 (N_12541,N_7154,N_9389);
xnor U12542 (N_12542,N_5135,N_8599);
nand U12543 (N_12543,N_7384,N_9990);
nor U12544 (N_12544,N_7337,N_7153);
nand U12545 (N_12545,N_9256,N_9944);
nand U12546 (N_12546,N_8205,N_8235);
or U12547 (N_12547,N_9371,N_8023);
and U12548 (N_12548,N_9155,N_6023);
nor U12549 (N_12549,N_5437,N_7829);
xor U12550 (N_12550,N_8277,N_7065);
xnor U12551 (N_12551,N_5412,N_5827);
xnor U12552 (N_12552,N_9314,N_5582);
and U12553 (N_12553,N_6290,N_7266);
and U12554 (N_12554,N_6644,N_7595);
or U12555 (N_12555,N_9835,N_9697);
or U12556 (N_12556,N_8413,N_7690);
nor U12557 (N_12557,N_8490,N_5982);
xnor U12558 (N_12558,N_6218,N_7649);
nand U12559 (N_12559,N_6656,N_9721);
or U12560 (N_12560,N_6334,N_7859);
and U12561 (N_12561,N_8881,N_6363);
nand U12562 (N_12562,N_7079,N_5696);
or U12563 (N_12563,N_6753,N_6894);
xnor U12564 (N_12564,N_8149,N_8092);
nand U12565 (N_12565,N_9156,N_5977);
nand U12566 (N_12566,N_5456,N_6335);
and U12567 (N_12567,N_6080,N_6464);
xnor U12568 (N_12568,N_8886,N_5411);
nor U12569 (N_12569,N_7180,N_6906);
nor U12570 (N_12570,N_6413,N_7330);
nand U12571 (N_12571,N_8868,N_9825);
nor U12572 (N_12572,N_7803,N_5657);
nor U12573 (N_12573,N_8311,N_9879);
or U12574 (N_12574,N_7723,N_8807);
and U12575 (N_12575,N_6983,N_5729);
xor U12576 (N_12576,N_6047,N_8752);
xnor U12577 (N_12577,N_7304,N_8848);
nor U12578 (N_12578,N_5610,N_6524);
nand U12579 (N_12579,N_9400,N_9457);
or U12580 (N_12580,N_9993,N_8829);
nand U12581 (N_12581,N_7768,N_5650);
and U12582 (N_12582,N_9975,N_5982);
nand U12583 (N_12583,N_6648,N_8396);
xor U12584 (N_12584,N_6190,N_9094);
xor U12585 (N_12585,N_9145,N_7730);
xnor U12586 (N_12586,N_8036,N_7145);
nor U12587 (N_12587,N_7340,N_6505);
and U12588 (N_12588,N_5515,N_9589);
and U12589 (N_12589,N_7588,N_7837);
or U12590 (N_12590,N_7655,N_6293);
or U12591 (N_12591,N_8413,N_5751);
nor U12592 (N_12592,N_7690,N_7759);
nand U12593 (N_12593,N_6180,N_8735);
xor U12594 (N_12594,N_8902,N_7066);
or U12595 (N_12595,N_8688,N_5944);
and U12596 (N_12596,N_5765,N_8054);
or U12597 (N_12597,N_7851,N_9751);
nand U12598 (N_12598,N_9904,N_6196);
and U12599 (N_12599,N_7924,N_6484);
nor U12600 (N_12600,N_7496,N_9658);
nor U12601 (N_12601,N_6136,N_7389);
nand U12602 (N_12602,N_8072,N_8033);
and U12603 (N_12603,N_6031,N_8228);
or U12604 (N_12604,N_5676,N_8689);
nand U12605 (N_12605,N_7261,N_5880);
nor U12606 (N_12606,N_9199,N_5642);
and U12607 (N_12607,N_8236,N_7168);
xnor U12608 (N_12608,N_7631,N_5061);
or U12609 (N_12609,N_6529,N_6912);
nor U12610 (N_12610,N_5554,N_8861);
nand U12611 (N_12611,N_8363,N_9540);
and U12612 (N_12612,N_5527,N_9372);
or U12613 (N_12613,N_7601,N_8533);
xnor U12614 (N_12614,N_6857,N_5378);
or U12615 (N_12615,N_8762,N_6036);
nand U12616 (N_12616,N_5603,N_5206);
and U12617 (N_12617,N_9250,N_9164);
xnor U12618 (N_12618,N_5045,N_9722);
nor U12619 (N_12619,N_9985,N_6700);
nor U12620 (N_12620,N_9966,N_7684);
and U12621 (N_12621,N_6049,N_5305);
and U12622 (N_12622,N_5799,N_7387);
xor U12623 (N_12623,N_7823,N_8789);
nor U12624 (N_12624,N_7222,N_7798);
or U12625 (N_12625,N_5042,N_9137);
nand U12626 (N_12626,N_6442,N_6842);
or U12627 (N_12627,N_6191,N_9338);
xor U12628 (N_12628,N_6260,N_6347);
xor U12629 (N_12629,N_6374,N_8156);
nor U12630 (N_12630,N_5190,N_9804);
and U12631 (N_12631,N_6969,N_6415);
nor U12632 (N_12632,N_9490,N_9286);
and U12633 (N_12633,N_8054,N_9976);
nand U12634 (N_12634,N_7341,N_5892);
nand U12635 (N_12635,N_9250,N_5863);
and U12636 (N_12636,N_5609,N_7472);
xnor U12637 (N_12637,N_7134,N_8852);
or U12638 (N_12638,N_9978,N_5715);
or U12639 (N_12639,N_9054,N_5397);
or U12640 (N_12640,N_9353,N_7415);
or U12641 (N_12641,N_7502,N_5908);
or U12642 (N_12642,N_7103,N_9351);
or U12643 (N_12643,N_7407,N_7744);
and U12644 (N_12644,N_6007,N_8661);
nand U12645 (N_12645,N_8198,N_8951);
nor U12646 (N_12646,N_5062,N_5200);
xnor U12647 (N_12647,N_6381,N_7771);
and U12648 (N_12648,N_9923,N_9636);
and U12649 (N_12649,N_6013,N_9079);
nor U12650 (N_12650,N_6329,N_9926);
xnor U12651 (N_12651,N_8746,N_6200);
xor U12652 (N_12652,N_6953,N_9695);
nand U12653 (N_12653,N_5223,N_7853);
xor U12654 (N_12654,N_6528,N_9016);
nor U12655 (N_12655,N_8491,N_6195);
nor U12656 (N_12656,N_5845,N_6634);
and U12657 (N_12657,N_7894,N_7394);
nand U12658 (N_12658,N_5971,N_7065);
nand U12659 (N_12659,N_6021,N_9857);
nand U12660 (N_12660,N_7818,N_6485);
nand U12661 (N_12661,N_5382,N_8891);
nand U12662 (N_12662,N_5159,N_8690);
or U12663 (N_12663,N_8937,N_9262);
and U12664 (N_12664,N_6357,N_9623);
xnor U12665 (N_12665,N_5092,N_9681);
nor U12666 (N_12666,N_8065,N_7852);
xnor U12667 (N_12667,N_5066,N_7735);
nor U12668 (N_12668,N_6333,N_6709);
and U12669 (N_12669,N_8319,N_6291);
nand U12670 (N_12670,N_5382,N_5751);
and U12671 (N_12671,N_7971,N_5414);
or U12672 (N_12672,N_8643,N_9603);
and U12673 (N_12673,N_7096,N_8394);
or U12674 (N_12674,N_5983,N_8398);
nand U12675 (N_12675,N_5278,N_6808);
nand U12676 (N_12676,N_5200,N_8690);
nand U12677 (N_12677,N_9592,N_6511);
or U12678 (N_12678,N_7789,N_9971);
or U12679 (N_12679,N_8184,N_9886);
nand U12680 (N_12680,N_6688,N_5456);
nand U12681 (N_12681,N_7453,N_8946);
nand U12682 (N_12682,N_9589,N_9970);
or U12683 (N_12683,N_7003,N_8305);
xnor U12684 (N_12684,N_7199,N_7740);
xnor U12685 (N_12685,N_8024,N_5161);
xnor U12686 (N_12686,N_5749,N_9157);
nor U12687 (N_12687,N_8269,N_9405);
and U12688 (N_12688,N_6065,N_6733);
or U12689 (N_12689,N_6722,N_7346);
xor U12690 (N_12690,N_5285,N_5151);
and U12691 (N_12691,N_8673,N_5235);
and U12692 (N_12692,N_9259,N_9426);
nor U12693 (N_12693,N_5605,N_5505);
and U12694 (N_12694,N_5642,N_6851);
xnor U12695 (N_12695,N_8693,N_6909);
nor U12696 (N_12696,N_8674,N_6019);
nand U12697 (N_12697,N_8231,N_9831);
and U12698 (N_12698,N_7291,N_5699);
and U12699 (N_12699,N_9123,N_5867);
nand U12700 (N_12700,N_6962,N_8753);
or U12701 (N_12701,N_7342,N_5979);
and U12702 (N_12702,N_7530,N_5065);
and U12703 (N_12703,N_9227,N_5095);
nor U12704 (N_12704,N_7607,N_6779);
and U12705 (N_12705,N_5529,N_6056);
or U12706 (N_12706,N_5184,N_9485);
xor U12707 (N_12707,N_9739,N_7907);
and U12708 (N_12708,N_8029,N_8962);
or U12709 (N_12709,N_6906,N_6066);
nor U12710 (N_12710,N_6042,N_5120);
nor U12711 (N_12711,N_6235,N_8792);
nor U12712 (N_12712,N_5373,N_5744);
xor U12713 (N_12713,N_5067,N_5262);
nand U12714 (N_12714,N_8808,N_6365);
nor U12715 (N_12715,N_6885,N_7804);
xor U12716 (N_12716,N_7629,N_9495);
nand U12717 (N_12717,N_9971,N_9861);
nor U12718 (N_12718,N_6598,N_6375);
or U12719 (N_12719,N_9472,N_5136);
and U12720 (N_12720,N_5458,N_6181);
nand U12721 (N_12721,N_8282,N_9944);
nand U12722 (N_12722,N_7292,N_5129);
xor U12723 (N_12723,N_9109,N_5153);
xnor U12724 (N_12724,N_8189,N_6773);
xnor U12725 (N_12725,N_6484,N_5183);
nor U12726 (N_12726,N_9983,N_7127);
nand U12727 (N_12727,N_8170,N_7940);
nand U12728 (N_12728,N_9191,N_9518);
and U12729 (N_12729,N_7147,N_9503);
nor U12730 (N_12730,N_6735,N_8515);
nor U12731 (N_12731,N_9379,N_9992);
or U12732 (N_12732,N_6681,N_7277);
and U12733 (N_12733,N_6322,N_8956);
and U12734 (N_12734,N_8230,N_8003);
or U12735 (N_12735,N_9265,N_8028);
xor U12736 (N_12736,N_5228,N_5554);
nand U12737 (N_12737,N_8373,N_6139);
xnor U12738 (N_12738,N_5258,N_8469);
nor U12739 (N_12739,N_8477,N_9281);
nor U12740 (N_12740,N_6470,N_5276);
nor U12741 (N_12741,N_7148,N_9440);
and U12742 (N_12742,N_7793,N_6186);
xor U12743 (N_12743,N_6968,N_7985);
xnor U12744 (N_12744,N_9328,N_9391);
xor U12745 (N_12745,N_9338,N_8651);
and U12746 (N_12746,N_5628,N_8716);
xor U12747 (N_12747,N_6955,N_7567);
xnor U12748 (N_12748,N_9197,N_7232);
xor U12749 (N_12749,N_7345,N_7858);
xor U12750 (N_12750,N_8323,N_8736);
nor U12751 (N_12751,N_7476,N_8899);
nor U12752 (N_12752,N_9154,N_8910);
or U12753 (N_12753,N_8421,N_7319);
xor U12754 (N_12754,N_7516,N_6131);
or U12755 (N_12755,N_7978,N_5324);
nor U12756 (N_12756,N_5133,N_6927);
or U12757 (N_12757,N_9146,N_5897);
nand U12758 (N_12758,N_9414,N_6755);
and U12759 (N_12759,N_9464,N_5680);
xor U12760 (N_12760,N_6211,N_8431);
xor U12761 (N_12761,N_8359,N_8260);
or U12762 (N_12762,N_7792,N_8413);
nor U12763 (N_12763,N_6812,N_5327);
and U12764 (N_12764,N_8920,N_5106);
nand U12765 (N_12765,N_6562,N_6396);
or U12766 (N_12766,N_6425,N_9688);
or U12767 (N_12767,N_8420,N_6642);
and U12768 (N_12768,N_6151,N_9571);
xor U12769 (N_12769,N_8769,N_5504);
or U12770 (N_12770,N_9589,N_5581);
nor U12771 (N_12771,N_9498,N_6199);
and U12772 (N_12772,N_5156,N_8794);
nor U12773 (N_12773,N_8689,N_6237);
nand U12774 (N_12774,N_9875,N_5054);
nand U12775 (N_12775,N_5469,N_9630);
or U12776 (N_12776,N_9318,N_9226);
nor U12777 (N_12777,N_7210,N_7146);
nand U12778 (N_12778,N_9759,N_9051);
or U12779 (N_12779,N_8311,N_5468);
nor U12780 (N_12780,N_7348,N_7622);
nand U12781 (N_12781,N_6573,N_6143);
nor U12782 (N_12782,N_5903,N_6826);
and U12783 (N_12783,N_9938,N_9970);
nand U12784 (N_12784,N_5272,N_8151);
or U12785 (N_12785,N_7477,N_9671);
nor U12786 (N_12786,N_6847,N_9779);
or U12787 (N_12787,N_5312,N_8059);
nor U12788 (N_12788,N_9785,N_8127);
nor U12789 (N_12789,N_9111,N_7853);
nor U12790 (N_12790,N_7167,N_7802);
and U12791 (N_12791,N_5987,N_7648);
and U12792 (N_12792,N_7516,N_8724);
and U12793 (N_12793,N_6063,N_7598);
nor U12794 (N_12794,N_5843,N_6269);
and U12795 (N_12795,N_7602,N_9733);
and U12796 (N_12796,N_7161,N_9728);
xnor U12797 (N_12797,N_5523,N_6114);
or U12798 (N_12798,N_9718,N_9434);
or U12799 (N_12799,N_5357,N_8837);
xnor U12800 (N_12800,N_7513,N_6954);
and U12801 (N_12801,N_5340,N_9725);
nor U12802 (N_12802,N_8931,N_7901);
or U12803 (N_12803,N_6014,N_7785);
nand U12804 (N_12804,N_6773,N_9044);
nor U12805 (N_12805,N_8304,N_6489);
and U12806 (N_12806,N_6226,N_8006);
xor U12807 (N_12807,N_6697,N_5625);
or U12808 (N_12808,N_5525,N_6864);
nor U12809 (N_12809,N_9862,N_6122);
or U12810 (N_12810,N_7123,N_9798);
nor U12811 (N_12811,N_7931,N_5788);
nor U12812 (N_12812,N_8372,N_5891);
or U12813 (N_12813,N_7651,N_7484);
nor U12814 (N_12814,N_9497,N_6195);
xnor U12815 (N_12815,N_7991,N_9490);
and U12816 (N_12816,N_8403,N_6730);
or U12817 (N_12817,N_9917,N_6776);
xor U12818 (N_12818,N_8233,N_7940);
nand U12819 (N_12819,N_8714,N_5807);
nand U12820 (N_12820,N_8497,N_8432);
xnor U12821 (N_12821,N_8580,N_5458);
and U12822 (N_12822,N_5099,N_7050);
nand U12823 (N_12823,N_5675,N_9210);
xnor U12824 (N_12824,N_9622,N_8202);
and U12825 (N_12825,N_9428,N_6988);
and U12826 (N_12826,N_6477,N_8886);
and U12827 (N_12827,N_9955,N_7994);
and U12828 (N_12828,N_8301,N_8123);
nor U12829 (N_12829,N_7815,N_9537);
nand U12830 (N_12830,N_8864,N_5000);
xor U12831 (N_12831,N_8725,N_5975);
and U12832 (N_12832,N_5908,N_9035);
nand U12833 (N_12833,N_8203,N_9604);
nor U12834 (N_12834,N_5703,N_5200);
and U12835 (N_12835,N_8258,N_8832);
or U12836 (N_12836,N_5013,N_6369);
nand U12837 (N_12837,N_9911,N_7976);
and U12838 (N_12838,N_9279,N_8050);
and U12839 (N_12839,N_9622,N_7297);
or U12840 (N_12840,N_7341,N_6569);
and U12841 (N_12841,N_9282,N_8943);
xnor U12842 (N_12842,N_6634,N_7871);
or U12843 (N_12843,N_7865,N_6829);
xor U12844 (N_12844,N_9728,N_7253);
xor U12845 (N_12845,N_5384,N_8039);
nor U12846 (N_12846,N_5475,N_5773);
or U12847 (N_12847,N_9751,N_9209);
xnor U12848 (N_12848,N_9035,N_7217);
and U12849 (N_12849,N_6669,N_7647);
xnor U12850 (N_12850,N_9891,N_6744);
and U12851 (N_12851,N_7329,N_7286);
and U12852 (N_12852,N_8290,N_6635);
nor U12853 (N_12853,N_5301,N_9833);
and U12854 (N_12854,N_9665,N_7207);
nor U12855 (N_12855,N_9993,N_7327);
nor U12856 (N_12856,N_9031,N_5457);
xnor U12857 (N_12857,N_7765,N_6903);
or U12858 (N_12858,N_8947,N_6215);
xor U12859 (N_12859,N_6874,N_8409);
xnor U12860 (N_12860,N_8326,N_7417);
or U12861 (N_12861,N_6232,N_9718);
xnor U12862 (N_12862,N_7215,N_8939);
nand U12863 (N_12863,N_8900,N_5410);
xor U12864 (N_12864,N_7929,N_7320);
or U12865 (N_12865,N_7136,N_9145);
nor U12866 (N_12866,N_8024,N_9916);
nor U12867 (N_12867,N_9835,N_8537);
nor U12868 (N_12868,N_6561,N_6006);
and U12869 (N_12869,N_7847,N_6539);
nor U12870 (N_12870,N_5793,N_5747);
nand U12871 (N_12871,N_8611,N_7197);
and U12872 (N_12872,N_9965,N_7729);
nand U12873 (N_12873,N_5545,N_7711);
xnor U12874 (N_12874,N_9798,N_7740);
nor U12875 (N_12875,N_5799,N_8668);
nor U12876 (N_12876,N_8907,N_8546);
nand U12877 (N_12877,N_8444,N_7496);
nand U12878 (N_12878,N_5006,N_5784);
and U12879 (N_12879,N_5407,N_5652);
and U12880 (N_12880,N_5653,N_7328);
or U12881 (N_12881,N_5664,N_5324);
nor U12882 (N_12882,N_8800,N_6933);
and U12883 (N_12883,N_5456,N_5957);
nor U12884 (N_12884,N_8513,N_8293);
nand U12885 (N_12885,N_8242,N_5242);
or U12886 (N_12886,N_6478,N_6515);
nor U12887 (N_12887,N_7788,N_9072);
nor U12888 (N_12888,N_7500,N_6842);
nor U12889 (N_12889,N_7019,N_8487);
xor U12890 (N_12890,N_8425,N_7778);
nor U12891 (N_12891,N_8432,N_9731);
nand U12892 (N_12892,N_6906,N_6329);
xnor U12893 (N_12893,N_7164,N_6954);
xor U12894 (N_12894,N_8881,N_6704);
or U12895 (N_12895,N_6096,N_9928);
nand U12896 (N_12896,N_9420,N_7130);
nor U12897 (N_12897,N_6146,N_6488);
and U12898 (N_12898,N_7365,N_6034);
nor U12899 (N_12899,N_5194,N_7491);
and U12900 (N_12900,N_7307,N_9795);
or U12901 (N_12901,N_5508,N_6849);
nor U12902 (N_12902,N_5251,N_7339);
or U12903 (N_12903,N_9402,N_6626);
or U12904 (N_12904,N_7992,N_9102);
xnor U12905 (N_12905,N_6804,N_6238);
and U12906 (N_12906,N_8689,N_6922);
nand U12907 (N_12907,N_8132,N_8548);
nand U12908 (N_12908,N_9748,N_9514);
nand U12909 (N_12909,N_6437,N_6335);
or U12910 (N_12910,N_5563,N_6187);
nor U12911 (N_12911,N_5350,N_7411);
nand U12912 (N_12912,N_5685,N_8273);
and U12913 (N_12913,N_8968,N_5784);
nor U12914 (N_12914,N_6627,N_9671);
nor U12915 (N_12915,N_9187,N_8962);
or U12916 (N_12916,N_8261,N_9329);
and U12917 (N_12917,N_8717,N_7742);
and U12918 (N_12918,N_7210,N_7027);
or U12919 (N_12919,N_7049,N_7671);
or U12920 (N_12920,N_5562,N_5412);
xor U12921 (N_12921,N_6391,N_6105);
or U12922 (N_12922,N_5890,N_8123);
or U12923 (N_12923,N_5259,N_7484);
xnor U12924 (N_12924,N_7081,N_5244);
xnor U12925 (N_12925,N_8729,N_6093);
nand U12926 (N_12926,N_7978,N_6700);
nor U12927 (N_12927,N_8392,N_9877);
nor U12928 (N_12928,N_8249,N_6235);
xor U12929 (N_12929,N_6404,N_7171);
nor U12930 (N_12930,N_7001,N_6404);
and U12931 (N_12931,N_7763,N_7438);
or U12932 (N_12932,N_8794,N_9805);
or U12933 (N_12933,N_5420,N_5909);
and U12934 (N_12934,N_5483,N_5571);
nand U12935 (N_12935,N_9968,N_6175);
and U12936 (N_12936,N_9574,N_9053);
nand U12937 (N_12937,N_7199,N_5987);
or U12938 (N_12938,N_7095,N_9117);
and U12939 (N_12939,N_8947,N_7340);
nor U12940 (N_12940,N_7034,N_5684);
xnor U12941 (N_12941,N_6408,N_7646);
and U12942 (N_12942,N_6153,N_5224);
and U12943 (N_12943,N_9872,N_6248);
xnor U12944 (N_12944,N_9409,N_5584);
or U12945 (N_12945,N_7405,N_5143);
and U12946 (N_12946,N_8836,N_6032);
xor U12947 (N_12947,N_9542,N_7559);
or U12948 (N_12948,N_9842,N_9398);
or U12949 (N_12949,N_5219,N_8256);
or U12950 (N_12950,N_6446,N_9347);
or U12951 (N_12951,N_7376,N_6451);
nor U12952 (N_12952,N_8618,N_8037);
nor U12953 (N_12953,N_9488,N_8446);
nand U12954 (N_12954,N_7011,N_9528);
or U12955 (N_12955,N_6441,N_8792);
or U12956 (N_12956,N_6175,N_5307);
xnor U12957 (N_12957,N_7585,N_8406);
nor U12958 (N_12958,N_7361,N_9820);
nand U12959 (N_12959,N_5385,N_9532);
and U12960 (N_12960,N_7184,N_9581);
or U12961 (N_12961,N_6272,N_5721);
nor U12962 (N_12962,N_8222,N_6980);
or U12963 (N_12963,N_6877,N_6243);
and U12964 (N_12964,N_6315,N_8895);
xnor U12965 (N_12965,N_6150,N_9482);
or U12966 (N_12966,N_7534,N_5867);
nor U12967 (N_12967,N_8056,N_6010);
nor U12968 (N_12968,N_8555,N_9139);
nor U12969 (N_12969,N_8868,N_8043);
and U12970 (N_12970,N_5864,N_5242);
nor U12971 (N_12971,N_6091,N_8533);
or U12972 (N_12972,N_9631,N_5706);
nor U12973 (N_12973,N_8348,N_8353);
and U12974 (N_12974,N_9652,N_9440);
nor U12975 (N_12975,N_5884,N_9961);
nand U12976 (N_12976,N_5712,N_7108);
nand U12977 (N_12977,N_9466,N_8316);
or U12978 (N_12978,N_6484,N_6049);
xor U12979 (N_12979,N_5341,N_8221);
nor U12980 (N_12980,N_7336,N_6975);
nand U12981 (N_12981,N_6875,N_6171);
nand U12982 (N_12982,N_8439,N_9773);
and U12983 (N_12983,N_9037,N_8875);
and U12984 (N_12984,N_9774,N_6249);
or U12985 (N_12985,N_8730,N_5903);
nand U12986 (N_12986,N_6926,N_9917);
nand U12987 (N_12987,N_7207,N_6571);
or U12988 (N_12988,N_8002,N_8989);
and U12989 (N_12989,N_8726,N_9344);
nor U12990 (N_12990,N_7617,N_7006);
or U12991 (N_12991,N_7924,N_9523);
nand U12992 (N_12992,N_9371,N_5225);
and U12993 (N_12993,N_5108,N_6108);
nand U12994 (N_12994,N_9514,N_8251);
nand U12995 (N_12995,N_8145,N_6722);
or U12996 (N_12996,N_8927,N_7741);
xor U12997 (N_12997,N_9628,N_5530);
and U12998 (N_12998,N_8314,N_6192);
nor U12999 (N_12999,N_9174,N_9007);
xor U13000 (N_13000,N_8892,N_5188);
xor U13001 (N_13001,N_6157,N_6154);
and U13002 (N_13002,N_5505,N_9387);
nand U13003 (N_13003,N_9025,N_5278);
and U13004 (N_13004,N_5501,N_8125);
or U13005 (N_13005,N_9299,N_9929);
nand U13006 (N_13006,N_6873,N_6943);
nand U13007 (N_13007,N_9037,N_7740);
and U13008 (N_13008,N_6357,N_9343);
or U13009 (N_13009,N_9796,N_9618);
xnor U13010 (N_13010,N_6973,N_9767);
and U13011 (N_13011,N_6039,N_9481);
and U13012 (N_13012,N_7395,N_5205);
and U13013 (N_13013,N_7659,N_6830);
or U13014 (N_13014,N_9853,N_6312);
xor U13015 (N_13015,N_9707,N_9032);
nor U13016 (N_13016,N_5694,N_7162);
nand U13017 (N_13017,N_7165,N_7800);
and U13018 (N_13018,N_8965,N_8603);
and U13019 (N_13019,N_5525,N_7466);
nor U13020 (N_13020,N_7510,N_5450);
and U13021 (N_13021,N_7904,N_9428);
and U13022 (N_13022,N_7932,N_5215);
and U13023 (N_13023,N_5626,N_7639);
xnor U13024 (N_13024,N_8804,N_7791);
xor U13025 (N_13025,N_7697,N_9861);
nor U13026 (N_13026,N_7223,N_8377);
or U13027 (N_13027,N_8349,N_5430);
or U13028 (N_13028,N_7200,N_7786);
nand U13029 (N_13029,N_6090,N_9438);
and U13030 (N_13030,N_7111,N_9610);
xor U13031 (N_13031,N_5166,N_7619);
xnor U13032 (N_13032,N_9144,N_9665);
or U13033 (N_13033,N_5088,N_6338);
nor U13034 (N_13034,N_9569,N_7894);
and U13035 (N_13035,N_6514,N_9548);
nand U13036 (N_13036,N_6877,N_6839);
and U13037 (N_13037,N_5361,N_5271);
or U13038 (N_13038,N_6294,N_6324);
nor U13039 (N_13039,N_9668,N_5235);
and U13040 (N_13040,N_6575,N_5494);
and U13041 (N_13041,N_9358,N_7187);
and U13042 (N_13042,N_5096,N_5898);
or U13043 (N_13043,N_5740,N_5584);
nand U13044 (N_13044,N_5985,N_6076);
nand U13045 (N_13045,N_6852,N_8482);
nor U13046 (N_13046,N_5480,N_7376);
nor U13047 (N_13047,N_6727,N_5473);
nor U13048 (N_13048,N_7924,N_6905);
nand U13049 (N_13049,N_6899,N_6803);
and U13050 (N_13050,N_8392,N_8314);
or U13051 (N_13051,N_9195,N_9478);
nand U13052 (N_13052,N_8094,N_5208);
and U13053 (N_13053,N_6895,N_9705);
xnor U13054 (N_13054,N_7457,N_8152);
nor U13055 (N_13055,N_9602,N_5757);
nor U13056 (N_13056,N_8063,N_7579);
or U13057 (N_13057,N_9796,N_8325);
nor U13058 (N_13058,N_6517,N_6820);
xor U13059 (N_13059,N_6827,N_6533);
or U13060 (N_13060,N_6263,N_8246);
and U13061 (N_13061,N_8897,N_5016);
nand U13062 (N_13062,N_5239,N_9325);
nor U13063 (N_13063,N_7302,N_5959);
nand U13064 (N_13064,N_8857,N_7256);
xor U13065 (N_13065,N_8997,N_6317);
and U13066 (N_13066,N_9481,N_9612);
or U13067 (N_13067,N_9966,N_7878);
nand U13068 (N_13068,N_7790,N_7983);
nand U13069 (N_13069,N_9644,N_7113);
nor U13070 (N_13070,N_5521,N_6745);
nor U13071 (N_13071,N_6559,N_8877);
nor U13072 (N_13072,N_6046,N_6503);
and U13073 (N_13073,N_9332,N_5705);
and U13074 (N_13074,N_6183,N_5309);
nor U13075 (N_13075,N_5291,N_7178);
xor U13076 (N_13076,N_6210,N_8254);
nand U13077 (N_13077,N_9440,N_8481);
nor U13078 (N_13078,N_6641,N_8891);
nand U13079 (N_13079,N_8715,N_8939);
or U13080 (N_13080,N_6888,N_7731);
xor U13081 (N_13081,N_8559,N_5909);
and U13082 (N_13082,N_7779,N_7287);
and U13083 (N_13083,N_6386,N_7703);
or U13084 (N_13084,N_9840,N_8313);
xnor U13085 (N_13085,N_6964,N_7707);
or U13086 (N_13086,N_8634,N_7756);
and U13087 (N_13087,N_6411,N_9596);
nor U13088 (N_13088,N_5720,N_7004);
nor U13089 (N_13089,N_5637,N_9941);
and U13090 (N_13090,N_8730,N_9996);
or U13091 (N_13091,N_5939,N_8627);
or U13092 (N_13092,N_9730,N_5104);
nand U13093 (N_13093,N_8965,N_6246);
and U13094 (N_13094,N_7438,N_5314);
xor U13095 (N_13095,N_6052,N_9403);
xor U13096 (N_13096,N_9047,N_7102);
xnor U13097 (N_13097,N_9437,N_6376);
and U13098 (N_13098,N_6763,N_9447);
nand U13099 (N_13099,N_6587,N_7309);
nand U13100 (N_13100,N_9262,N_6006);
or U13101 (N_13101,N_6392,N_7883);
and U13102 (N_13102,N_6863,N_9380);
nand U13103 (N_13103,N_9668,N_8201);
nor U13104 (N_13104,N_6254,N_6557);
and U13105 (N_13105,N_6366,N_5952);
and U13106 (N_13106,N_5506,N_6222);
xor U13107 (N_13107,N_7560,N_5246);
xnor U13108 (N_13108,N_7787,N_9235);
nand U13109 (N_13109,N_5305,N_8890);
xor U13110 (N_13110,N_5419,N_8159);
nand U13111 (N_13111,N_8217,N_6304);
xor U13112 (N_13112,N_8806,N_6107);
and U13113 (N_13113,N_9569,N_7460);
xnor U13114 (N_13114,N_8216,N_9514);
nand U13115 (N_13115,N_8174,N_5010);
or U13116 (N_13116,N_9108,N_8108);
nor U13117 (N_13117,N_5527,N_6509);
xnor U13118 (N_13118,N_7315,N_8528);
or U13119 (N_13119,N_9823,N_6881);
and U13120 (N_13120,N_7841,N_6821);
xnor U13121 (N_13121,N_7117,N_9593);
or U13122 (N_13122,N_6212,N_6656);
or U13123 (N_13123,N_9098,N_6363);
nand U13124 (N_13124,N_5475,N_8340);
and U13125 (N_13125,N_7654,N_7746);
and U13126 (N_13126,N_5865,N_6497);
nor U13127 (N_13127,N_8275,N_8485);
nor U13128 (N_13128,N_8021,N_8675);
and U13129 (N_13129,N_9429,N_9058);
nand U13130 (N_13130,N_7389,N_9495);
xnor U13131 (N_13131,N_7186,N_6410);
nand U13132 (N_13132,N_6028,N_5291);
or U13133 (N_13133,N_8711,N_6577);
and U13134 (N_13134,N_5586,N_8132);
or U13135 (N_13135,N_9908,N_8938);
or U13136 (N_13136,N_7510,N_9360);
and U13137 (N_13137,N_8559,N_6831);
nor U13138 (N_13138,N_9621,N_9656);
or U13139 (N_13139,N_5685,N_5551);
xor U13140 (N_13140,N_5870,N_6172);
nor U13141 (N_13141,N_8194,N_8838);
nor U13142 (N_13142,N_8435,N_8118);
and U13143 (N_13143,N_7274,N_6512);
and U13144 (N_13144,N_6344,N_5635);
xor U13145 (N_13145,N_5796,N_9421);
nand U13146 (N_13146,N_8116,N_8534);
or U13147 (N_13147,N_6496,N_7182);
nand U13148 (N_13148,N_7514,N_5566);
xor U13149 (N_13149,N_7257,N_6043);
xnor U13150 (N_13150,N_8602,N_9040);
and U13151 (N_13151,N_6709,N_6571);
or U13152 (N_13152,N_7638,N_9806);
nand U13153 (N_13153,N_5801,N_6943);
nand U13154 (N_13154,N_7763,N_8590);
xor U13155 (N_13155,N_9262,N_6240);
and U13156 (N_13156,N_9695,N_7809);
and U13157 (N_13157,N_6453,N_7015);
xor U13158 (N_13158,N_7178,N_6957);
nor U13159 (N_13159,N_7676,N_6153);
nor U13160 (N_13160,N_8667,N_9387);
nor U13161 (N_13161,N_9575,N_5721);
or U13162 (N_13162,N_8666,N_8397);
nand U13163 (N_13163,N_9314,N_7708);
nor U13164 (N_13164,N_5544,N_8349);
xnor U13165 (N_13165,N_6894,N_7857);
nor U13166 (N_13166,N_8950,N_7565);
xnor U13167 (N_13167,N_7787,N_6378);
nand U13168 (N_13168,N_8208,N_6361);
and U13169 (N_13169,N_9484,N_5619);
nor U13170 (N_13170,N_9588,N_9337);
nand U13171 (N_13171,N_8058,N_9460);
xor U13172 (N_13172,N_6093,N_5091);
and U13173 (N_13173,N_9499,N_6493);
or U13174 (N_13174,N_8278,N_6610);
or U13175 (N_13175,N_5375,N_8406);
or U13176 (N_13176,N_5938,N_5551);
or U13177 (N_13177,N_9667,N_7869);
xor U13178 (N_13178,N_7373,N_7670);
xnor U13179 (N_13179,N_7298,N_5327);
or U13180 (N_13180,N_5932,N_7689);
nor U13181 (N_13181,N_7717,N_5059);
xnor U13182 (N_13182,N_7113,N_8438);
nor U13183 (N_13183,N_6005,N_7860);
nand U13184 (N_13184,N_5817,N_9477);
xor U13185 (N_13185,N_7074,N_7556);
nand U13186 (N_13186,N_5305,N_6935);
nor U13187 (N_13187,N_5865,N_9406);
or U13188 (N_13188,N_7545,N_8137);
xnor U13189 (N_13189,N_6466,N_8090);
nor U13190 (N_13190,N_5094,N_6425);
nand U13191 (N_13191,N_9075,N_7673);
or U13192 (N_13192,N_8276,N_5606);
nor U13193 (N_13193,N_8125,N_8355);
nor U13194 (N_13194,N_6844,N_5586);
nand U13195 (N_13195,N_5117,N_8417);
or U13196 (N_13196,N_9139,N_8114);
or U13197 (N_13197,N_6090,N_5148);
xor U13198 (N_13198,N_9169,N_6187);
and U13199 (N_13199,N_5508,N_6045);
nand U13200 (N_13200,N_7314,N_8120);
and U13201 (N_13201,N_8696,N_6203);
xor U13202 (N_13202,N_9340,N_5704);
nand U13203 (N_13203,N_5842,N_6786);
and U13204 (N_13204,N_8039,N_6086);
nor U13205 (N_13205,N_7940,N_9309);
or U13206 (N_13206,N_8105,N_7281);
xor U13207 (N_13207,N_5182,N_6851);
and U13208 (N_13208,N_8839,N_7544);
xor U13209 (N_13209,N_9652,N_5567);
nand U13210 (N_13210,N_9352,N_9001);
and U13211 (N_13211,N_8894,N_6689);
nor U13212 (N_13212,N_5752,N_8564);
nor U13213 (N_13213,N_5768,N_9367);
or U13214 (N_13214,N_9488,N_5189);
nor U13215 (N_13215,N_7969,N_7306);
or U13216 (N_13216,N_5726,N_5323);
nand U13217 (N_13217,N_9922,N_6210);
nand U13218 (N_13218,N_9461,N_9129);
or U13219 (N_13219,N_6455,N_8624);
nand U13220 (N_13220,N_8055,N_7703);
xor U13221 (N_13221,N_5980,N_5391);
and U13222 (N_13222,N_6564,N_5685);
xnor U13223 (N_13223,N_5400,N_5664);
xnor U13224 (N_13224,N_5552,N_7577);
and U13225 (N_13225,N_6729,N_6456);
and U13226 (N_13226,N_8793,N_7423);
and U13227 (N_13227,N_6400,N_8422);
and U13228 (N_13228,N_9387,N_8306);
or U13229 (N_13229,N_6557,N_5388);
or U13230 (N_13230,N_9542,N_9792);
and U13231 (N_13231,N_7740,N_9052);
nor U13232 (N_13232,N_5117,N_9777);
nor U13233 (N_13233,N_5776,N_8106);
xor U13234 (N_13234,N_9311,N_6756);
nor U13235 (N_13235,N_5145,N_9981);
nor U13236 (N_13236,N_7798,N_7850);
and U13237 (N_13237,N_9676,N_8117);
xnor U13238 (N_13238,N_5150,N_9621);
or U13239 (N_13239,N_8131,N_5338);
or U13240 (N_13240,N_8949,N_6046);
and U13241 (N_13241,N_8762,N_6544);
and U13242 (N_13242,N_9993,N_6144);
or U13243 (N_13243,N_9778,N_9402);
or U13244 (N_13244,N_8239,N_6269);
nand U13245 (N_13245,N_9732,N_8157);
xnor U13246 (N_13246,N_5934,N_9834);
nor U13247 (N_13247,N_9930,N_6781);
or U13248 (N_13248,N_7939,N_8938);
or U13249 (N_13249,N_5402,N_7149);
nor U13250 (N_13250,N_8740,N_8419);
nand U13251 (N_13251,N_9983,N_8157);
or U13252 (N_13252,N_9296,N_6017);
nor U13253 (N_13253,N_7242,N_8523);
nand U13254 (N_13254,N_8548,N_9465);
or U13255 (N_13255,N_5596,N_9097);
or U13256 (N_13256,N_8440,N_5193);
xor U13257 (N_13257,N_8866,N_8844);
xor U13258 (N_13258,N_5729,N_8061);
or U13259 (N_13259,N_9092,N_5241);
or U13260 (N_13260,N_5989,N_8265);
nor U13261 (N_13261,N_9900,N_8652);
nand U13262 (N_13262,N_7779,N_6722);
and U13263 (N_13263,N_8956,N_5602);
nand U13264 (N_13264,N_5153,N_8096);
nor U13265 (N_13265,N_8147,N_6912);
xor U13266 (N_13266,N_5454,N_6896);
nand U13267 (N_13267,N_7180,N_5634);
xor U13268 (N_13268,N_6003,N_9328);
and U13269 (N_13269,N_6896,N_8797);
or U13270 (N_13270,N_5562,N_8273);
nand U13271 (N_13271,N_5992,N_9441);
or U13272 (N_13272,N_8368,N_8229);
xor U13273 (N_13273,N_9221,N_6875);
nand U13274 (N_13274,N_5522,N_7974);
or U13275 (N_13275,N_6901,N_7145);
or U13276 (N_13276,N_9449,N_7547);
nor U13277 (N_13277,N_5255,N_5765);
nand U13278 (N_13278,N_6807,N_9265);
nand U13279 (N_13279,N_6429,N_9048);
xor U13280 (N_13280,N_8456,N_5000);
or U13281 (N_13281,N_6012,N_9711);
xor U13282 (N_13282,N_5646,N_5180);
nand U13283 (N_13283,N_9268,N_8479);
xor U13284 (N_13284,N_7779,N_9206);
nor U13285 (N_13285,N_9564,N_5996);
nand U13286 (N_13286,N_9500,N_6731);
nor U13287 (N_13287,N_7103,N_5836);
nand U13288 (N_13288,N_6893,N_7479);
nand U13289 (N_13289,N_6557,N_5811);
nand U13290 (N_13290,N_6939,N_8452);
and U13291 (N_13291,N_9345,N_7128);
or U13292 (N_13292,N_8148,N_9895);
nor U13293 (N_13293,N_5893,N_7216);
and U13294 (N_13294,N_7561,N_9355);
and U13295 (N_13295,N_6567,N_8120);
xor U13296 (N_13296,N_7078,N_9793);
or U13297 (N_13297,N_8602,N_8884);
or U13298 (N_13298,N_7245,N_5318);
and U13299 (N_13299,N_9992,N_7226);
and U13300 (N_13300,N_5178,N_9072);
nor U13301 (N_13301,N_6488,N_6959);
xnor U13302 (N_13302,N_8876,N_6380);
and U13303 (N_13303,N_7771,N_6118);
and U13304 (N_13304,N_8837,N_9143);
and U13305 (N_13305,N_6232,N_5130);
nor U13306 (N_13306,N_9770,N_5293);
nor U13307 (N_13307,N_9846,N_6228);
and U13308 (N_13308,N_7800,N_7194);
and U13309 (N_13309,N_6475,N_7118);
and U13310 (N_13310,N_7875,N_5980);
xor U13311 (N_13311,N_8401,N_7289);
and U13312 (N_13312,N_7958,N_6578);
nand U13313 (N_13313,N_6103,N_7166);
and U13314 (N_13314,N_8118,N_6617);
and U13315 (N_13315,N_9024,N_6999);
and U13316 (N_13316,N_5289,N_9995);
nor U13317 (N_13317,N_6088,N_8428);
or U13318 (N_13318,N_5572,N_5215);
or U13319 (N_13319,N_6566,N_9255);
or U13320 (N_13320,N_9907,N_9634);
xnor U13321 (N_13321,N_5954,N_7156);
or U13322 (N_13322,N_7068,N_6161);
xnor U13323 (N_13323,N_7678,N_7456);
nor U13324 (N_13324,N_7797,N_9338);
nor U13325 (N_13325,N_7024,N_7424);
or U13326 (N_13326,N_6636,N_6737);
nor U13327 (N_13327,N_8147,N_5252);
nor U13328 (N_13328,N_6035,N_5590);
or U13329 (N_13329,N_6383,N_9298);
nor U13330 (N_13330,N_6356,N_8835);
nand U13331 (N_13331,N_9698,N_7263);
and U13332 (N_13332,N_8145,N_8013);
nand U13333 (N_13333,N_6305,N_8839);
xnor U13334 (N_13334,N_7735,N_5487);
nand U13335 (N_13335,N_9677,N_7638);
and U13336 (N_13336,N_9304,N_5696);
or U13337 (N_13337,N_6591,N_6004);
nor U13338 (N_13338,N_5067,N_5255);
and U13339 (N_13339,N_9046,N_6733);
xor U13340 (N_13340,N_7804,N_5334);
nand U13341 (N_13341,N_8108,N_6160);
and U13342 (N_13342,N_7126,N_5722);
xnor U13343 (N_13343,N_8409,N_5612);
xor U13344 (N_13344,N_5249,N_7551);
nand U13345 (N_13345,N_6395,N_7471);
nor U13346 (N_13346,N_6696,N_7087);
nand U13347 (N_13347,N_5352,N_5132);
and U13348 (N_13348,N_6949,N_6182);
and U13349 (N_13349,N_8042,N_8473);
nor U13350 (N_13350,N_8310,N_6272);
xnor U13351 (N_13351,N_9967,N_8733);
nor U13352 (N_13352,N_6420,N_5421);
nor U13353 (N_13353,N_5475,N_7067);
or U13354 (N_13354,N_8993,N_9893);
nand U13355 (N_13355,N_9436,N_6917);
or U13356 (N_13356,N_9206,N_5005);
nor U13357 (N_13357,N_9757,N_9651);
nor U13358 (N_13358,N_9578,N_5263);
xor U13359 (N_13359,N_8894,N_9075);
xor U13360 (N_13360,N_6135,N_8100);
xor U13361 (N_13361,N_7271,N_9997);
nor U13362 (N_13362,N_7204,N_8523);
and U13363 (N_13363,N_8339,N_7729);
nand U13364 (N_13364,N_6214,N_6439);
and U13365 (N_13365,N_7053,N_6467);
or U13366 (N_13366,N_5449,N_9053);
xnor U13367 (N_13367,N_8179,N_8362);
nand U13368 (N_13368,N_7777,N_6291);
or U13369 (N_13369,N_7810,N_5914);
or U13370 (N_13370,N_8441,N_7586);
nand U13371 (N_13371,N_8459,N_7082);
nor U13372 (N_13372,N_8171,N_8605);
nor U13373 (N_13373,N_7440,N_9621);
xnor U13374 (N_13374,N_8993,N_6302);
and U13375 (N_13375,N_6612,N_9660);
nor U13376 (N_13376,N_8532,N_8404);
nand U13377 (N_13377,N_8128,N_8055);
nand U13378 (N_13378,N_8848,N_6738);
xnor U13379 (N_13379,N_5390,N_8005);
nor U13380 (N_13380,N_9110,N_7116);
nand U13381 (N_13381,N_7374,N_6492);
or U13382 (N_13382,N_8939,N_7081);
nor U13383 (N_13383,N_9653,N_9517);
nand U13384 (N_13384,N_9476,N_6422);
xor U13385 (N_13385,N_5737,N_6826);
nor U13386 (N_13386,N_5944,N_7962);
nor U13387 (N_13387,N_7813,N_9117);
and U13388 (N_13388,N_8792,N_8749);
nor U13389 (N_13389,N_9021,N_9467);
or U13390 (N_13390,N_7254,N_7697);
nor U13391 (N_13391,N_9328,N_9451);
nor U13392 (N_13392,N_9689,N_9675);
and U13393 (N_13393,N_9077,N_8682);
nor U13394 (N_13394,N_8990,N_7154);
nand U13395 (N_13395,N_8163,N_7202);
xnor U13396 (N_13396,N_6564,N_6208);
nor U13397 (N_13397,N_5797,N_9346);
xnor U13398 (N_13398,N_9343,N_6280);
xnor U13399 (N_13399,N_9437,N_5782);
nor U13400 (N_13400,N_6575,N_9943);
or U13401 (N_13401,N_8265,N_6384);
or U13402 (N_13402,N_7260,N_5077);
and U13403 (N_13403,N_6336,N_8072);
nand U13404 (N_13404,N_9429,N_8830);
nor U13405 (N_13405,N_8393,N_7494);
and U13406 (N_13406,N_6170,N_9216);
xnor U13407 (N_13407,N_5614,N_7956);
xor U13408 (N_13408,N_9303,N_9398);
nor U13409 (N_13409,N_9665,N_8751);
or U13410 (N_13410,N_9130,N_8848);
and U13411 (N_13411,N_7820,N_8761);
and U13412 (N_13412,N_5354,N_8673);
and U13413 (N_13413,N_7304,N_7087);
nand U13414 (N_13414,N_5975,N_8641);
xnor U13415 (N_13415,N_5029,N_5401);
nand U13416 (N_13416,N_9493,N_7606);
xnor U13417 (N_13417,N_5017,N_9484);
or U13418 (N_13418,N_8209,N_9950);
or U13419 (N_13419,N_8114,N_7160);
and U13420 (N_13420,N_5264,N_8745);
nor U13421 (N_13421,N_9031,N_6065);
nor U13422 (N_13422,N_9242,N_9239);
nor U13423 (N_13423,N_7492,N_8352);
nor U13424 (N_13424,N_7719,N_6592);
nand U13425 (N_13425,N_6599,N_8636);
nor U13426 (N_13426,N_9772,N_5889);
and U13427 (N_13427,N_7814,N_6019);
and U13428 (N_13428,N_5968,N_8976);
nand U13429 (N_13429,N_5925,N_6346);
nor U13430 (N_13430,N_9903,N_8511);
or U13431 (N_13431,N_9471,N_9406);
nor U13432 (N_13432,N_6521,N_6662);
nand U13433 (N_13433,N_8344,N_6261);
nand U13434 (N_13434,N_6465,N_6265);
nor U13435 (N_13435,N_9372,N_8793);
nand U13436 (N_13436,N_6553,N_9750);
nor U13437 (N_13437,N_6966,N_8076);
nand U13438 (N_13438,N_6626,N_5130);
nand U13439 (N_13439,N_5555,N_8858);
nand U13440 (N_13440,N_9813,N_9174);
and U13441 (N_13441,N_7947,N_7937);
or U13442 (N_13442,N_6855,N_9537);
nand U13443 (N_13443,N_6677,N_6984);
nor U13444 (N_13444,N_9462,N_7546);
and U13445 (N_13445,N_8151,N_7804);
nor U13446 (N_13446,N_7755,N_8021);
and U13447 (N_13447,N_7144,N_6090);
nor U13448 (N_13448,N_5108,N_7274);
nand U13449 (N_13449,N_7289,N_7232);
nor U13450 (N_13450,N_7904,N_8279);
xor U13451 (N_13451,N_9008,N_5404);
or U13452 (N_13452,N_5898,N_8200);
and U13453 (N_13453,N_7647,N_6061);
nand U13454 (N_13454,N_7880,N_7883);
nor U13455 (N_13455,N_5801,N_6399);
or U13456 (N_13456,N_6275,N_5827);
xor U13457 (N_13457,N_7289,N_5874);
xnor U13458 (N_13458,N_9288,N_7818);
or U13459 (N_13459,N_7048,N_6489);
xnor U13460 (N_13460,N_7164,N_8193);
xor U13461 (N_13461,N_9484,N_6614);
and U13462 (N_13462,N_5500,N_6068);
nor U13463 (N_13463,N_7755,N_9857);
nand U13464 (N_13464,N_8376,N_7870);
xor U13465 (N_13465,N_6673,N_7945);
nand U13466 (N_13466,N_9700,N_7581);
nand U13467 (N_13467,N_5239,N_5751);
xnor U13468 (N_13468,N_7186,N_8904);
nand U13469 (N_13469,N_5850,N_6563);
or U13470 (N_13470,N_5905,N_9685);
nand U13471 (N_13471,N_6200,N_5761);
nand U13472 (N_13472,N_8312,N_8618);
nor U13473 (N_13473,N_7018,N_8233);
or U13474 (N_13474,N_9767,N_5600);
nand U13475 (N_13475,N_9050,N_9318);
nor U13476 (N_13476,N_9531,N_9608);
nor U13477 (N_13477,N_7841,N_6579);
nor U13478 (N_13478,N_5771,N_5819);
or U13479 (N_13479,N_6558,N_8067);
nor U13480 (N_13480,N_7107,N_9195);
and U13481 (N_13481,N_7516,N_9095);
and U13482 (N_13482,N_8099,N_6403);
xnor U13483 (N_13483,N_8453,N_6336);
nor U13484 (N_13484,N_6201,N_9288);
nand U13485 (N_13485,N_7963,N_5878);
and U13486 (N_13486,N_9468,N_9635);
nand U13487 (N_13487,N_6046,N_7453);
nor U13488 (N_13488,N_5694,N_8482);
or U13489 (N_13489,N_9086,N_9042);
nor U13490 (N_13490,N_8159,N_5525);
xnor U13491 (N_13491,N_7499,N_9067);
or U13492 (N_13492,N_6745,N_9200);
or U13493 (N_13493,N_6001,N_7332);
nand U13494 (N_13494,N_9907,N_9155);
xnor U13495 (N_13495,N_7405,N_8435);
nand U13496 (N_13496,N_5148,N_8668);
and U13497 (N_13497,N_9734,N_9112);
xor U13498 (N_13498,N_8997,N_9477);
nand U13499 (N_13499,N_8930,N_7779);
nand U13500 (N_13500,N_7389,N_9520);
nor U13501 (N_13501,N_9100,N_8481);
xor U13502 (N_13502,N_8034,N_8682);
nand U13503 (N_13503,N_9591,N_8534);
nand U13504 (N_13504,N_8143,N_8756);
and U13505 (N_13505,N_9605,N_8176);
nor U13506 (N_13506,N_6782,N_5579);
nor U13507 (N_13507,N_7322,N_7361);
and U13508 (N_13508,N_9279,N_8165);
xor U13509 (N_13509,N_9832,N_5695);
xnor U13510 (N_13510,N_7531,N_7234);
or U13511 (N_13511,N_9013,N_8802);
or U13512 (N_13512,N_8875,N_8445);
nand U13513 (N_13513,N_5886,N_7750);
nor U13514 (N_13514,N_6487,N_9449);
and U13515 (N_13515,N_9963,N_5114);
xnor U13516 (N_13516,N_9824,N_7990);
and U13517 (N_13517,N_8084,N_5252);
xor U13518 (N_13518,N_7525,N_5104);
nor U13519 (N_13519,N_8029,N_9609);
and U13520 (N_13520,N_6912,N_8020);
nor U13521 (N_13521,N_6459,N_7332);
or U13522 (N_13522,N_5981,N_8104);
and U13523 (N_13523,N_5423,N_6097);
nor U13524 (N_13524,N_7783,N_6354);
xnor U13525 (N_13525,N_9413,N_7573);
or U13526 (N_13526,N_6529,N_7783);
and U13527 (N_13527,N_9067,N_5014);
xnor U13528 (N_13528,N_6779,N_8227);
nor U13529 (N_13529,N_5285,N_8628);
or U13530 (N_13530,N_6932,N_8852);
nor U13531 (N_13531,N_8988,N_9000);
and U13532 (N_13532,N_6533,N_7083);
nand U13533 (N_13533,N_7911,N_9639);
nand U13534 (N_13534,N_7314,N_9595);
and U13535 (N_13535,N_5005,N_9829);
xnor U13536 (N_13536,N_8096,N_8013);
and U13537 (N_13537,N_7481,N_8422);
and U13538 (N_13538,N_7281,N_9614);
or U13539 (N_13539,N_6805,N_9244);
or U13540 (N_13540,N_8306,N_5692);
nand U13541 (N_13541,N_7929,N_7152);
xor U13542 (N_13542,N_5142,N_7083);
or U13543 (N_13543,N_6123,N_6490);
xor U13544 (N_13544,N_8331,N_5225);
nor U13545 (N_13545,N_9260,N_6610);
nor U13546 (N_13546,N_8358,N_5868);
nor U13547 (N_13547,N_8363,N_9925);
nand U13548 (N_13548,N_7207,N_7187);
nor U13549 (N_13549,N_7880,N_8026);
xor U13550 (N_13550,N_7682,N_8156);
nand U13551 (N_13551,N_8621,N_6274);
and U13552 (N_13552,N_9317,N_6727);
nand U13553 (N_13553,N_9257,N_7578);
xor U13554 (N_13554,N_7220,N_5706);
nand U13555 (N_13555,N_8264,N_6308);
nand U13556 (N_13556,N_7733,N_8446);
nor U13557 (N_13557,N_7369,N_9901);
nand U13558 (N_13558,N_7661,N_9167);
xnor U13559 (N_13559,N_5545,N_5882);
nand U13560 (N_13560,N_8266,N_5120);
nor U13561 (N_13561,N_8511,N_7046);
nor U13562 (N_13562,N_5792,N_9603);
xor U13563 (N_13563,N_9371,N_7909);
nor U13564 (N_13564,N_9176,N_5799);
nor U13565 (N_13565,N_9313,N_5479);
nand U13566 (N_13566,N_6427,N_8116);
or U13567 (N_13567,N_6625,N_7519);
xor U13568 (N_13568,N_6835,N_5736);
nor U13569 (N_13569,N_5559,N_5987);
nor U13570 (N_13570,N_5820,N_5279);
nand U13571 (N_13571,N_5869,N_5832);
and U13572 (N_13572,N_5768,N_6208);
or U13573 (N_13573,N_6601,N_5445);
or U13574 (N_13574,N_6079,N_7211);
nand U13575 (N_13575,N_8488,N_8940);
nand U13576 (N_13576,N_8774,N_6279);
xnor U13577 (N_13577,N_6302,N_5542);
nand U13578 (N_13578,N_5534,N_8670);
and U13579 (N_13579,N_9623,N_7629);
and U13580 (N_13580,N_9449,N_8894);
xnor U13581 (N_13581,N_7338,N_7618);
or U13582 (N_13582,N_5474,N_6367);
nor U13583 (N_13583,N_7237,N_7687);
nand U13584 (N_13584,N_5711,N_7184);
nand U13585 (N_13585,N_7428,N_9040);
or U13586 (N_13586,N_6672,N_9879);
nor U13587 (N_13587,N_5353,N_7945);
xor U13588 (N_13588,N_7608,N_8034);
nand U13589 (N_13589,N_9566,N_7811);
nor U13590 (N_13590,N_9905,N_8931);
nand U13591 (N_13591,N_7025,N_7659);
nor U13592 (N_13592,N_9759,N_5957);
nand U13593 (N_13593,N_5722,N_8912);
xor U13594 (N_13594,N_5595,N_8594);
xnor U13595 (N_13595,N_8373,N_6478);
nand U13596 (N_13596,N_8391,N_7076);
xor U13597 (N_13597,N_8371,N_7522);
xnor U13598 (N_13598,N_8732,N_7487);
and U13599 (N_13599,N_5598,N_5632);
nor U13600 (N_13600,N_9462,N_7877);
or U13601 (N_13601,N_7889,N_6484);
nand U13602 (N_13602,N_5280,N_7702);
xnor U13603 (N_13603,N_7332,N_5775);
nor U13604 (N_13604,N_9667,N_8733);
nor U13605 (N_13605,N_6838,N_7965);
nor U13606 (N_13606,N_7263,N_9857);
nand U13607 (N_13607,N_8791,N_5032);
or U13608 (N_13608,N_9042,N_9855);
nor U13609 (N_13609,N_7921,N_9011);
or U13610 (N_13610,N_8381,N_5837);
nor U13611 (N_13611,N_5510,N_6371);
nor U13612 (N_13612,N_6481,N_7261);
nor U13613 (N_13613,N_9451,N_9754);
or U13614 (N_13614,N_5051,N_8537);
or U13615 (N_13615,N_6143,N_5689);
nor U13616 (N_13616,N_7459,N_6351);
nand U13617 (N_13617,N_5515,N_9090);
xor U13618 (N_13618,N_5016,N_6849);
nor U13619 (N_13619,N_5491,N_5454);
or U13620 (N_13620,N_5121,N_7939);
nand U13621 (N_13621,N_6912,N_5249);
nand U13622 (N_13622,N_8204,N_6838);
xnor U13623 (N_13623,N_9741,N_9646);
nor U13624 (N_13624,N_6752,N_6676);
nor U13625 (N_13625,N_8121,N_6159);
xor U13626 (N_13626,N_5005,N_6076);
xor U13627 (N_13627,N_6578,N_6359);
xor U13628 (N_13628,N_6718,N_6473);
nor U13629 (N_13629,N_8710,N_8875);
and U13630 (N_13630,N_5384,N_6676);
and U13631 (N_13631,N_9549,N_9425);
nand U13632 (N_13632,N_8414,N_8200);
or U13633 (N_13633,N_7136,N_9064);
xnor U13634 (N_13634,N_8974,N_5295);
nor U13635 (N_13635,N_6926,N_8406);
nor U13636 (N_13636,N_5663,N_9593);
or U13637 (N_13637,N_5281,N_9995);
xor U13638 (N_13638,N_6341,N_6613);
or U13639 (N_13639,N_7449,N_5620);
and U13640 (N_13640,N_7174,N_5391);
xor U13641 (N_13641,N_8462,N_6649);
and U13642 (N_13642,N_6502,N_6043);
and U13643 (N_13643,N_6860,N_5492);
nor U13644 (N_13644,N_8750,N_9366);
xor U13645 (N_13645,N_6645,N_8983);
and U13646 (N_13646,N_7939,N_8241);
and U13647 (N_13647,N_9821,N_7283);
and U13648 (N_13648,N_9711,N_9790);
nand U13649 (N_13649,N_5675,N_6533);
and U13650 (N_13650,N_9809,N_9211);
nor U13651 (N_13651,N_8258,N_7830);
and U13652 (N_13652,N_6028,N_8994);
nor U13653 (N_13653,N_7016,N_7518);
xnor U13654 (N_13654,N_8732,N_9704);
nand U13655 (N_13655,N_8570,N_8770);
or U13656 (N_13656,N_6313,N_5387);
nand U13657 (N_13657,N_8468,N_7000);
or U13658 (N_13658,N_6725,N_9234);
xnor U13659 (N_13659,N_9704,N_9381);
and U13660 (N_13660,N_5488,N_7433);
and U13661 (N_13661,N_7627,N_8376);
or U13662 (N_13662,N_5541,N_8058);
and U13663 (N_13663,N_9849,N_6685);
and U13664 (N_13664,N_5705,N_6807);
xor U13665 (N_13665,N_5959,N_8211);
xor U13666 (N_13666,N_5402,N_6534);
or U13667 (N_13667,N_5004,N_7876);
nor U13668 (N_13668,N_5746,N_5128);
xor U13669 (N_13669,N_6293,N_5271);
or U13670 (N_13670,N_8505,N_6983);
and U13671 (N_13671,N_8807,N_8402);
nand U13672 (N_13672,N_9138,N_5210);
and U13673 (N_13673,N_7979,N_5440);
nor U13674 (N_13674,N_9402,N_6492);
or U13675 (N_13675,N_5031,N_9132);
nand U13676 (N_13676,N_7789,N_8270);
nor U13677 (N_13677,N_5759,N_8015);
or U13678 (N_13678,N_8592,N_5222);
nor U13679 (N_13679,N_9255,N_5142);
nand U13680 (N_13680,N_5366,N_9953);
xnor U13681 (N_13681,N_7458,N_8251);
xnor U13682 (N_13682,N_7921,N_8469);
nor U13683 (N_13683,N_9253,N_9281);
nand U13684 (N_13684,N_9519,N_5383);
and U13685 (N_13685,N_7101,N_6816);
xnor U13686 (N_13686,N_8299,N_8147);
nand U13687 (N_13687,N_8928,N_7235);
nor U13688 (N_13688,N_6139,N_6608);
xnor U13689 (N_13689,N_6721,N_5571);
xnor U13690 (N_13690,N_9143,N_9920);
xnor U13691 (N_13691,N_8207,N_8760);
nor U13692 (N_13692,N_7098,N_7071);
and U13693 (N_13693,N_9883,N_8613);
xnor U13694 (N_13694,N_9282,N_9094);
nor U13695 (N_13695,N_8841,N_9545);
or U13696 (N_13696,N_9366,N_7174);
nor U13697 (N_13697,N_9214,N_8968);
or U13698 (N_13698,N_9630,N_6286);
or U13699 (N_13699,N_6914,N_6034);
nor U13700 (N_13700,N_9576,N_6541);
nor U13701 (N_13701,N_7041,N_7890);
and U13702 (N_13702,N_5651,N_7028);
nor U13703 (N_13703,N_7823,N_6357);
nand U13704 (N_13704,N_7418,N_5768);
nor U13705 (N_13705,N_5730,N_7830);
nor U13706 (N_13706,N_9211,N_8766);
nand U13707 (N_13707,N_8015,N_9979);
or U13708 (N_13708,N_5083,N_9723);
nand U13709 (N_13709,N_8375,N_7841);
and U13710 (N_13710,N_8966,N_8963);
nor U13711 (N_13711,N_5284,N_8350);
xnor U13712 (N_13712,N_8950,N_8767);
and U13713 (N_13713,N_8064,N_6943);
xnor U13714 (N_13714,N_8008,N_9928);
nand U13715 (N_13715,N_8513,N_5262);
nand U13716 (N_13716,N_9980,N_5827);
and U13717 (N_13717,N_6343,N_6247);
or U13718 (N_13718,N_8740,N_9586);
xor U13719 (N_13719,N_9241,N_7515);
or U13720 (N_13720,N_6290,N_7030);
nand U13721 (N_13721,N_9543,N_5202);
xnor U13722 (N_13722,N_6304,N_5244);
xor U13723 (N_13723,N_7404,N_7872);
xnor U13724 (N_13724,N_9980,N_6782);
nor U13725 (N_13725,N_5632,N_8654);
and U13726 (N_13726,N_7833,N_9797);
nor U13727 (N_13727,N_5605,N_9711);
or U13728 (N_13728,N_8063,N_5433);
nor U13729 (N_13729,N_8813,N_5096);
nand U13730 (N_13730,N_5833,N_8449);
and U13731 (N_13731,N_6320,N_8890);
nand U13732 (N_13732,N_6755,N_5680);
nor U13733 (N_13733,N_5577,N_9120);
nor U13734 (N_13734,N_5236,N_8623);
xnor U13735 (N_13735,N_5981,N_5387);
nor U13736 (N_13736,N_8515,N_9871);
xor U13737 (N_13737,N_9519,N_9772);
or U13738 (N_13738,N_9825,N_9723);
xor U13739 (N_13739,N_6868,N_7115);
and U13740 (N_13740,N_8970,N_6102);
or U13741 (N_13741,N_9167,N_8119);
nor U13742 (N_13742,N_5095,N_9647);
nand U13743 (N_13743,N_9711,N_6606);
nor U13744 (N_13744,N_7976,N_9146);
nand U13745 (N_13745,N_6790,N_8499);
and U13746 (N_13746,N_8263,N_7896);
and U13747 (N_13747,N_8161,N_5962);
nor U13748 (N_13748,N_5336,N_8140);
xor U13749 (N_13749,N_9944,N_5726);
or U13750 (N_13750,N_7992,N_5965);
or U13751 (N_13751,N_5758,N_6166);
or U13752 (N_13752,N_5322,N_8596);
nand U13753 (N_13753,N_9479,N_7421);
nand U13754 (N_13754,N_7555,N_9684);
nor U13755 (N_13755,N_8235,N_7628);
nor U13756 (N_13756,N_8771,N_6718);
xnor U13757 (N_13757,N_6927,N_9274);
xor U13758 (N_13758,N_9291,N_8831);
and U13759 (N_13759,N_6020,N_7526);
nand U13760 (N_13760,N_5000,N_5609);
and U13761 (N_13761,N_6007,N_7406);
xor U13762 (N_13762,N_9169,N_7599);
or U13763 (N_13763,N_9905,N_5030);
nand U13764 (N_13764,N_6401,N_6994);
nor U13765 (N_13765,N_6963,N_7423);
xnor U13766 (N_13766,N_8025,N_6028);
and U13767 (N_13767,N_6023,N_5408);
xor U13768 (N_13768,N_5754,N_5426);
or U13769 (N_13769,N_5134,N_6318);
xnor U13770 (N_13770,N_5716,N_5015);
nor U13771 (N_13771,N_9678,N_8219);
or U13772 (N_13772,N_9732,N_9657);
and U13773 (N_13773,N_6009,N_5390);
nand U13774 (N_13774,N_5801,N_6006);
nand U13775 (N_13775,N_5312,N_6758);
and U13776 (N_13776,N_6764,N_9330);
or U13777 (N_13777,N_7534,N_9604);
nand U13778 (N_13778,N_8773,N_9251);
xnor U13779 (N_13779,N_9968,N_7266);
nor U13780 (N_13780,N_5303,N_7725);
nand U13781 (N_13781,N_8177,N_6617);
nand U13782 (N_13782,N_7405,N_6077);
nor U13783 (N_13783,N_7500,N_9179);
and U13784 (N_13784,N_7422,N_6514);
nor U13785 (N_13785,N_9212,N_7498);
xor U13786 (N_13786,N_8665,N_8418);
nor U13787 (N_13787,N_8491,N_7105);
nand U13788 (N_13788,N_9117,N_5786);
nor U13789 (N_13789,N_7275,N_9144);
or U13790 (N_13790,N_9970,N_5038);
xor U13791 (N_13791,N_6904,N_7579);
and U13792 (N_13792,N_7249,N_7986);
nor U13793 (N_13793,N_7845,N_5117);
xor U13794 (N_13794,N_5920,N_8781);
or U13795 (N_13795,N_9619,N_9989);
and U13796 (N_13796,N_6923,N_7388);
xnor U13797 (N_13797,N_9350,N_8111);
and U13798 (N_13798,N_6716,N_7059);
xnor U13799 (N_13799,N_7419,N_6234);
nor U13800 (N_13800,N_8083,N_9585);
and U13801 (N_13801,N_5992,N_6012);
nor U13802 (N_13802,N_7653,N_8061);
nor U13803 (N_13803,N_7862,N_7162);
xor U13804 (N_13804,N_8468,N_9487);
or U13805 (N_13805,N_9312,N_6816);
nor U13806 (N_13806,N_7816,N_7259);
xnor U13807 (N_13807,N_7008,N_5456);
xnor U13808 (N_13808,N_9074,N_8679);
and U13809 (N_13809,N_7753,N_5044);
xor U13810 (N_13810,N_6327,N_9216);
nor U13811 (N_13811,N_5138,N_9566);
nand U13812 (N_13812,N_6293,N_6784);
or U13813 (N_13813,N_6712,N_9497);
nor U13814 (N_13814,N_9724,N_5664);
and U13815 (N_13815,N_7319,N_9735);
xnor U13816 (N_13816,N_7508,N_5675);
nand U13817 (N_13817,N_8684,N_8705);
and U13818 (N_13818,N_6135,N_5813);
nand U13819 (N_13819,N_8438,N_8714);
nand U13820 (N_13820,N_8967,N_8104);
xor U13821 (N_13821,N_9681,N_7174);
nand U13822 (N_13822,N_5299,N_9006);
nor U13823 (N_13823,N_7757,N_5206);
or U13824 (N_13824,N_7463,N_7315);
nor U13825 (N_13825,N_9055,N_8805);
nand U13826 (N_13826,N_6484,N_5998);
and U13827 (N_13827,N_6420,N_8736);
nor U13828 (N_13828,N_8548,N_7659);
nor U13829 (N_13829,N_9438,N_6030);
nand U13830 (N_13830,N_7029,N_8552);
and U13831 (N_13831,N_5925,N_7135);
xnor U13832 (N_13832,N_9943,N_5705);
nor U13833 (N_13833,N_7191,N_7522);
xnor U13834 (N_13834,N_7331,N_8700);
xor U13835 (N_13835,N_5719,N_5243);
nand U13836 (N_13836,N_8448,N_6221);
nor U13837 (N_13837,N_9914,N_7578);
and U13838 (N_13838,N_9384,N_7310);
or U13839 (N_13839,N_9093,N_9117);
and U13840 (N_13840,N_5854,N_6515);
xnor U13841 (N_13841,N_9676,N_5639);
and U13842 (N_13842,N_9835,N_5085);
or U13843 (N_13843,N_9225,N_5347);
and U13844 (N_13844,N_6661,N_5465);
and U13845 (N_13845,N_7797,N_9962);
nor U13846 (N_13846,N_5329,N_6406);
and U13847 (N_13847,N_5671,N_6956);
or U13848 (N_13848,N_9180,N_8415);
nand U13849 (N_13849,N_7339,N_6699);
xor U13850 (N_13850,N_8426,N_9626);
nand U13851 (N_13851,N_6059,N_8197);
nor U13852 (N_13852,N_5502,N_9459);
and U13853 (N_13853,N_5999,N_7873);
and U13854 (N_13854,N_6317,N_6675);
or U13855 (N_13855,N_8860,N_6308);
or U13856 (N_13856,N_8813,N_7958);
nand U13857 (N_13857,N_8907,N_7268);
and U13858 (N_13858,N_8034,N_7258);
nor U13859 (N_13859,N_8341,N_6631);
or U13860 (N_13860,N_8270,N_9496);
nand U13861 (N_13861,N_8585,N_7907);
xnor U13862 (N_13862,N_6152,N_8821);
nor U13863 (N_13863,N_5908,N_6139);
and U13864 (N_13864,N_7528,N_7684);
nand U13865 (N_13865,N_6626,N_6763);
nand U13866 (N_13866,N_6168,N_6282);
xnor U13867 (N_13867,N_8189,N_6715);
nand U13868 (N_13868,N_6705,N_8769);
or U13869 (N_13869,N_6332,N_7956);
xnor U13870 (N_13870,N_6629,N_9992);
nand U13871 (N_13871,N_9971,N_7274);
and U13872 (N_13872,N_9278,N_9345);
and U13873 (N_13873,N_9709,N_8261);
or U13874 (N_13874,N_6240,N_9956);
nand U13875 (N_13875,N_5654,N_8781);
or U13876 (N_13876,N_8211,N_9256);
xnor U13877 (N_13877,N_9233,N_5507);
or U13878 (N_13878,N_9775,N_8203);
or U13879 (N_13879,N_8290,N_6568);
and U13880 (N_13880,N_6359,N_6524);
xnor U13881 (N_13881,N_5515,N_7172);
or U13882 (N_13882,N_7536,N_5419);
xor U13883 (N_13883,N_9208,N_9710);
nand U13884 (N_13884,N_6755,N_6923);
xnor U13885 (N_13885,N_6900,N_8463);
and U13886 (N_13886,N_7662,N_9892);
nand U13887 (N_13887,N_7776,N_8064);
xor U13888 (N_13888,N_9778,N_5659);
and U13889 (N_13889,N_5854,N_5239);
and U13890 (N_13890,N_9191,N_6891);
or U13891 (N_13891,N_9971,N_8063);
and U13892 (N_13892,N_6046,N_6279);
nor U13893 (N_13893,N_9375,N_9023);
nand U13894 (N_13894,N_8014,N_8131);
or U13895 (N_13895,N_6372,N_8565);
nor U13896 (N_13896,N_7604,N_9395);
and U13897 (N_13897,N_7097,N_8621);
nor U13898 (N_13898,N_5837,N_7936);
xor U13899 (N_13899,N_7766,N_8583);
nand U13900 (N_13900,N_6496,N_5749);
or U13901 (N_13901,N_7479,N_8184);
and U13902 (N_13902,N_5881,N_6832);
or U13903 (N_13903,N_6888,N_8697);
or U13904 (N_13904,N_6095,N_7396);
nor U13905 (N_13905,N_6237,N_6385);
nand U13906 (N_13906,N_8776,N_7526);
nor U13907 (N_13907,N_7496,N_7266);
or U13908 (N_13908,N_7119,N_7283);
and U13909 (N_13909,N_7881,N_9114);
nor U13910 (N_13910,N_5347,N_5346);
nand U13911 (N_13911,N_5570,N_5428);
nor U13912 (N_13912,N_5886,N_7100);
xnor U13913 (N_13913,N_8024,N_8495);
xor U13914 (N_13914,N_7560,N_9247);
and U13915 (N_13915,N_5589,N_8712);
xnor U13916 (N_13916,N_8735,N_6799);
and U13917 (N_13917,N_6210,N_8247);
nand U13918 (N_13918,N_7153,N_9029);
xor U13919 (N_13919,N_8141,N_6555);
or U13920 (N_13920,N_5586,N_7279);
or U13921 (N_13921,N_6223,N_6117);
and U13922 (N_13922,N_5574,N_9867);
nand U13923 (N_13923,N_8835,N_7233);
xor U13924 (N_13924,N_9447,N_6025);
nor U13925 (N_13925,N_6864,N_9427);
and U13926 (N_13926,N_5453,N_6531);
nor U13927 (N_13927,N_7719,N_7661);
nand U13928 (N_13928,N_8627,N_7052);
nor U13929 (N_13929,N_5848,N_5768);
xnor U13930 (N_13930,N_7287,N_9171);
nand U13931 (N_13931,N_8297,N_7449);
and U13932 (N_13932,N_6540,N_5483);
nand U13933 (N_13933,N_5949,N_5174);
or U13934 (N_13934,N_7920,N_6014);
nor U13935 (N_13935,N_6721,N_7354);
nor U13936 (N_13936,N_8390,N_5651);
nand U13937 (N_13937,N_5370,N_6962);
xor U13938 (N_13938,N_6824,N_5560);
nand U13939 (N_13939,N_6513,N_5454);
or U13940 (N_13940,N_7459,N_7456);
xnor U13941 (N_13941,N_8973,N_5393);
and U13942 (N_13942,N_9998,N_5723);
and U13943 (N_13943,N_8514,N_8827);
xnor U13944 (N_13944,N_5084,N_5457);
nand U13945 (N_13945,N_7999,N_9891);
nor U13946 (N_13946,N_5461,N_5873);
nor U13947 (N_13947,N_6931,N_5480);
or U13948 (N_13948,N_8180,N_7364);
and U13949 (N_13949,N_9462,N_5009);
nand U13950 (N_13950,N_9488,N_7570);
and U13951 (N_13951,N_9684,N_8447);
and U13952 (N_13952,N_7598,N_5433);
nor U13953 (N_13953,N_6967,N_9920);
nand U13954 (N_13954,N_6241,N_8534);
xor U13955 (N_13955,N_9750,N_5871);
and U13956 (N_13956,N_5717,N_8772);
xor U13957 (N_13957,N_7844,N_7529);
xnor U13958 (N_13958,N_5487,N_7508);
xor U13959 (N_13959,N_7810,N_8411);
nor U13960 (N_13960,N_8899,N_5046);
or U13961 (N_13961,N_9187,N_6362);
or U13962 (N_13962,N_9283,N_5253);
or U13963 (N_13963,N_5398,N_7141);
nor U13964 (N_13964,N_8073,N_7300);
nand U13965 (N_13965,N_8463,N_5222);
xor U13966 (N_13966,N_8671,N_8040);
nor U13967 (N_13967,N_8365,N_8517);
nand U13968 (N_13968,N_5666,N_8675);
or U13969 (N_13969,N_7310,N_6676);
or U13970 (N_13970,N_7103,N_6206);
nor U13971 (N_13971,N_8129,N_8274);
and U13972 (N_13972,N_5506,N_6674);
nand U13973 (N_13973,N_5496,N_6647);
nand U13974 (N_13974,N_9341,N_8344);
or U13975 (N_13975,N_6359,N_6430);
nand U13976 (N_13976,N_9603,N_9239);
nand U13977 (N_13977,N_8365,N_9346);
xor U13978 (N_13978,N_6157,N_9923);
or U13979 (N_13979,N_5889,N_9421);
xnor U13980 (N_13980,N_7326,N_7835);
nand U13981 (N_13981,N_5143,N_8818);
and U13982 (N_13982,N_8581,N_6588);
nor U13983 (N_13983,N_8869,N_8471);
nor U13984 (N_13984,N_9692,N_7609);
xnor U13985 (N_13985,N_8824,N_9381);
and U13986 (N_13986,N_5149,N_7753);
nand U13987 (N_13987,N_5814,N_9905);
xnor U13988 (N_13988,N_5846,N_5223);
or U13989 (N_13989,N_5532,N_7201);
nand U13990 (N_13990,N_5104,N_8781);
xnor U13991 (N_13991,N_9969,N_8877);
and U13992 (N_13992,N_5184,N_6778);
xnor U13993 (N_13993,N_7723,N_8091);
nand U13994 (N_13994,N_8333,N_7132);
and U13995 (N_13995,N_8840,N_9175);
and U13996 (N_13996,N_9464,N_8199);
xor U13997 (N_13997,N_6720,N_9571);
xnor U13998 (N_13998,N_5630,N_5995);
nand U13999 (N_13999,N_9424,N_6951);
xor U14000 (N_14000,N_6480,N_5983);
or U14001 (N_14001,N_5357,N_9419);
and U14002 (N_14002,N_5671,N_9589);
or U14003 (N_14003,N_9586,N_5423);
xnor U14004 (N_14004,N_7510,N_5071);
nand U14005 (N_14005,N_9673,N_9755);
or U14006 (N_14006,N_9613,N_7512);
or U14007 (N_14007,N_8271,N_9714);
nor U14008 (N_14008,N_9732,N_9268);
nor U14009 (N_14009,N_9640,N_9500);
and U14010 (N_14010,N_8756,N_7028);
and U14011 (N_14011,N_6265,N_7082);
and U14012 (N_14012,N_7248,N_5058);
or U14013 (N_14013,N_5232,N_5039);
xnor U14014 (N_14014,N_9300,N_6571);
nor U14015 (N_14015,N_7255,N_8363);
and U14016 (N_14016,N_9009,N_5659);
nand U14017 (N_14017,N_9153,N_9480);
and U14018 (N_14018,N_7408,N_8710);
nor U14019 (N_14019,N_9997,N_7751);
nor U14020 (N_14020,N_6444,N_5535);
or U14021 (N_14021,N_9138,N_6915);
and U14022 (N_14022,N_8717,N_7345);
or U14023 (N_14023,N_9412,N_5540);
or U14024 (N_14024,N_5995,N_6774);
xnor U14025 (N_14025,N_9483,N_6590);
xor U14026 (N_14026,N_7740,N_8593);
nor U14027 (N_14027,N_7978,N_7498);
or U14028 (N_14028,N_6182,N_7576);
and U14029 (N_14029,N_5310,N_6459);
nand U14030 (N_14030,N_5216,N_6057);
nand U14031 (N_14031,N_9815,N_9774);
and U14032 (N_14032,N_8172,N_9409);
xor U14033 (N_14033,N_6676,N_9370);
nand U14034 (N_14034,N_5809,N_7265);
nor U14035 (N_14035,N_5703,N_5930);
nor U14036 (N_14036,N_8024,N_5830);
nor U14037 (N_14037,N_7084,N_8655);
or U14038 (N_14038,N_5754,N_6734);
nand U14039 (N_14039,N_6207,N_6353);
nor U14040 (N_14040,N_5111,N_5302);
nor U14041 (N_14041,N_9253,N_5445);
or U14042 (N_14042,N_9563,N_6936);
nor U14043 (N_14043,N_7705,N_7902);
nand U14044 (N_14044,N_8264,N_5974);
nand U14045 (N_14045,N_9871,N_7178);
and U14046 (N_14046,N_7758,N_9680);
xor U14047 (N_14047,N_9035,N_8301);
and U14048 (N_14048,N_7031,N_9005);
and U14049 (N_14049,N_7725,N_7698);
nand U14050 (N_14050,N_6520,N_7058);
nor U14051 (N_14051,N_5531,N_8194);
nor U14052 (N_14052,N_5728,N_8837);
xor U14053 (N_14053,N_9617,N_5445);
and U14054 (N_14054,N_7120,N_7032);
xor U14055 (N_14055,N_8589,N_5097);
nand U14056 (N_14056,N_6165,N_9919);
nand U14057 (N_14057,N_9753,N_9695);
or U14058 (N_14058,N_9393,N_5638);
and U14059 (N_14059,N_7863,N_6916);
or U14060 (N_14060,N_8448,N_8855);
and U14061 (N_14061,N_7196,N_8571);
nor U14062 (N_14062,N_7837,N_6701);
xnor U14063 (N_14063,N_8290,N_5461);
nor U14064 (N_14064,N_6181,N_8844);
nor U14065 (N_14065,N_8768,N_6469);
or U14066 (N_14066,N_8320,N_9724);
xor U14067 (N_14067,N_9292,N_8674);
and U14068 (N_14068,N_6828,N_9755);
nor U14069 (N_14069,N_6034,N_6143);
nand U14070 (N_14070,N_8996,N_5409);
or U14071 (N_14071,N_6367,N_9660);
nand U14072 (N_14072,N_9426,N_8809);
and U14073 (N_14073,N_8341,N_7438);
and U14074 (N_14074,N_9460,N_7907);
or U14075 (N_14075,N_7820,N_8108);
nor U14076 (N_14076,N_7377,N_6602);
nor U14077 (N_14077,N_9505,N_5625);
and U14078 (N_14078,N_6865,N_8530);
or U14079 (N_14079,N_8679,N_5085);
or U14080 (N_14080,N_6396,N_7017);
or U14081 (N_14081,N_8212,N_7018);
xnor U14082 (N_14082,N_9038,N_7936);
or U14083 (N_14083,N_6619,N_6023);
nor U14084 (N_14084,N_5388,N_8614);
or U14085 (N_14085,N_7990,N_6415);
nor U14086 (N_14086,N_8917,N_7507);
and U14087 (N_14087,N_7323,N_6108);
or U14088 (N_14088,N_5726,N_8020);
xor U14089 (N_14089,N_8158,N_7057);
nand U14090 (N_14090,N_6377,N_5929);
and U14091 (N_14091,N_8825,N_9040);
xor U14092 (N_14092,N_6456,N_5546);
and U14093 (N_14093,N_7013,N_5561);
and U14094 (N_14094,N_7250,N_6574);
or U14095 (N_14095,N_5846,N_5321);
xnor U14096 (N_14096,N_8837,N_9854);
or U14097 (N_14097,N_6342,N_9036);
or U14098 (N_14098,N_9613,N_6306);
nand U14099 (N_14099,N_5309,N_6260);
xnor U14100 (N_14100,N_9324,N_7711);
nand U14101 (N_14101,N_9194,N_8645);
nor U14102 (N_14102,N_7287,N_7414);
nand U14103 (N_14103,N_7282,N_8747);
and U14104 (N_14104,N_5547,N_8368);
xnor U14105 (N_14105,N_6055,N_8939);
nor U14106 (N_14106,N_9661,N_5768);
nand U14107 (N_14107,N_6242,N_5625);
nor U14108 (N_14108,N_9313,N_5090);
xnor U14109 (N_14109,N_7984,N_6681);
nand U14110 (N_14110,N_7099,N_7524);
nand U14111 (N_14111,N_7090,N_6299);
nand U14112 (N_14112,N_7080,N_8596);
nor U14113 (N_14113,N_5596,N_5256);
and U14114 (N_14114,N_7141,N_8676);
and U14115 (N_14115,N_7129,N_9072);
or U14116 (N_14116,N_8783,N_9143);
xor U14117 (N_14117,N_7954,N_7241);
nor U14118 (N_14118,N_5700,N_5509);
or U14119 (N_14119,N_8091,N_5053);
or U14120 (N_14120,N_8166,N_7457);
nor U14121 (N_14121,N_7689,N_5551);
xor U14122 (N_14122,N_6316,N_5524);
nor U14123 (N_14123,N_7392,N_8682);
xnor U14124 (N_14124,N_6746,N_8373);
and U14125 (N_14125,N_8986,N_5451);
and U14126 (N_14126,N_5268,N_7881);
xor U14127 (N_14127,N_5409,N_6431);
nand U14128 (N_14128,N_9037,N_5797);
nor U14129 (N_14129,N_6114,N_9454);
or U14130 (N_14130,N_5816,N_5703);
xor U14131 (N_14131,N_7176,N_5543);
xor U14132 (N_14132,N_5307,N_9897);
and U14133 (N_14133,N_6667,N_8589);
nand U14134 (N_14134,N_9973,N_7748);
nor U14135 (N_14135,N_5296,N_9454);
nor U14136 (N_14136,N_7956,N_7163);
and U14137 (N_14137,N_7884,N_5031);
or U14138 (N_14138,N_9988,N_9029);
nand U14139 (N_14139,N_6700,N_6875);
xnor U14140 (N_14140,N_7851,N_5346);
and U14141 (N_14141,N_8326,N_7871);
or U14142 (N_14142,N_7238,N_9837);
or U14143 (N_14143,N_8376,N_5296);
nand U14144 (N_14144,N_9518,N_5649);
nor U14145 (N_14145,N_8725,N_9494);
nor U14146 (N_14146,N_9014,N_6622);
or U14147 (N_14147,N_7114,N_9232);
or U14148 (N_14148,N_7436,N_6679);
or U14149 (N_14149,N_5884,N_5973);
and U14150 (N_14150,N_7620,N_8482);
or U14151 (N_14151,N_9280,N_5756);
and U14152 (N_14152,N_5747,N_8425);
or U14153 (N_14153,N_6882,N_8426);
and U14154 (N_14154,N_5031,N_6231);
nor U14155 (N_14155,N_5946,N_7121);
nand U14156 (N_14156,N_9812,N_7081);
xor U14157 (N_14157,N_5572,N_7467);
nand U14158 (N_14158,N_7580,N_6396);
or U14159 (N_14159,N_7544,N_5096);
or U14160 (N_14160,N_6066,N_7748);
or U14161 (N_14161,N_6203,N_6651);
nor U14162 (N_14162,N_7653,N_7409);
nand U14163 (N_14163,N_6895,N_7179);
nor U14164 (N_14164,N_5163,N_7826);
nand U14165 (N_14165,N_7260,N_7710);
and U14166 (N_14166,N_6287,N_7986);
and U14167 (N_14167,N_9071,N_9567);
nand U14168 (N_14168,N_9426,N_7970);
nand U14169 (N_14169,N_8286,N_5814);
xor U14170 (N_14170,N_8724,N_8928);
or U14171 (N_14171,N_9443,N_5023);
nand U14172 (N_14172,N_9136,N_5345);
and U14173 (N_14173,N_7196,N_7358);
or U14174 (N_14174,N_8957,N_9676);
or U14175 (N_14175,N_6995,N_8575);
nor U14176 (N_14176,N_8002,N_9027);
and U14177 (N_14177,N_8753,N_7793);
and U14178 (N_14178,N_8573,N_8365);
and U14179 (N_14179,N_5425,N_7592);
or U14180 (N_14180,N_5752,N_7870);
or U14181 (N_14181,N_6638,N_6266);
xor U14182 (N_14182,N_5648,N_5531);
or U14183 (N_14183,N_7487,N_7360);
nor U14184 (N_14184,N_5886,N_6209);
nor U14185 (N_14185,N_8345,N_7847);
nor U14186 (N_14186,N_6928,N_9893);
or U14187 (N_14187,N_6539,N_7512);
nor U14188 (N_14188,N_5636,N_9687);
xor U14189 (N_14189,N_9551,N_8493);
xor U14190 (N_14190,N_7743,N_6542);
nand U14191 (N_14191,N_6188,N_7705);
nor U14192 (N_14192,N_8390,N_6286);
nor U14193 (N_14193,N_7273,N_7929);
nor U14194 (N_14194,N_5421,N_6388);
or U14195 (N_14195,N_7725,N_8476);
or U14196 (N_14196,N_9770,N_5356);
nand U14197 (N_14197,N_6344,N_5892);
or U14198 (N_14198,N_5138,N_5826);
nand U14199 (N_14199,N_5010,N_9406);
or U14200 (N_14200,N_5602,N_8631);
nor U14201 (N_14201,N_7509,N_7661);
or U14202 (N_14202,N_9180,N_6259);
nand U14203 (N_14203,N_8782,N_6618);
or U14204 (N_14204,N_5236,N_5893);
and U14205 (N_14205,N_9263,N_9955);
or U14206 (N_14206,N_5638,N_9009);
nor U14207 (N_14207,N_8371,N_5653);
or U14208 (N_14208,N_8875,N_5387);
nand U14209 (N_14209,N_6709,N_6828);
nor U14210 (N_14210,N_5189,N_5883);
and U14211 (N_14211,N_9584,N_7499);
or U14212 (N_14212,N_7899,N_9837);
xnor U14213 (N_14213,N_6935,N_9672);
nor U14214 (N_14214,N_7767,N_8605);
xor U14215 (N_14215,N_6695,N_7700);
nor U14216 (N_14216,N_6731,N_7869);
or U14217 (N_14217,N_9235,N_7134);
and U14218 (N_14218,N_8218,N_7380);
or U14219 (N_14219,N_7095,N_7812);
nand U14220 (N_14220,N_6422,N_8002);
nor U14221 (N_14221,N_6869,N_6510);
nor U14222 (N_14222,N_9039,N_6739);
nand U14223 (N_14223,N_6775,N_7140);
nor U14224 (N_14224,N_8937,N_9561);
and U14225 (N_14225,N_7254,N_7544);
xnor U14226 (N_14226,N_8733,N_8113);
and U14227 (N_14227,N_6236,N_8562);
nor U14228 (N_14228,N_9688,N_8846);
nor U14229 (N_14229,N_6572,N_5822);
xnor U14230 (N_14230,N_7583,N_7311);
and U14231 (N_14231,N_6498,N_9210);
xnor U14232 (N_14232,N_6952,N_9584);
or U14233 (N_14233,N_8992,N_5051);
nor U14234 (N_14234,N_5051,N_6338);
xor U14235 (N_14235,N_8846,N_5557);
and U14236 (N_14236,N_8398,N_7788);
nor U14237 (N_14237,N_6180,N_7358);
nand U14238 (N_14238,N_8924,N_9766);
nand U14239 (N_14239,N_9433,N_5606);
nor U14240 (N_14240,N_5568,N_5601);
nor U14241 (N_14241,N_5914,N_9735);
nor U14242 (N_14242,N_8135,N_8419);
and U14243 (N_14243,N_8253,N_9767);
nor U14244 (N_14244,N_9996,N_6562);
and U14245 (N_14245,N_7741,N_9837);
or U14246 (N_14246,N_5083,N_6367);
or U14247 (N_14247,N_7966,N_7917);
nor U14248 (N_14248,N_7348,N_9326);
or U14249 (N_14249,N_6941,N_6491);
nor U14250 (N_14250,N_9825,N_6983);
and U14251 (N_14251,N_7429,N_5792);
or U14252 (N_14252,N_6033,N_8821);
nand U14253 (N_14253,N_6281,N_5507);
nand U14254 (N_14254,N_9457,N_7651);
nor U14255 (N_14255,N_9618,N_8323);
or U14256 (N_14256,N_5356,N_7424);
or U14257 (N_14257,N_6628,N_9796);
xnor U14258 (N_14258,N_6365,N_7632);
or U14259 (N_14259,N_6416,N_5066);
nand U14260 (N_14260,N_9531,N_9185);
and U14261 (N_14261,N_6751,N_7334);
nand U14262 (N_14262,N_6017,N_6108);
nor U14263 (N_14263,N_7297,N_7876);
or U14264 (N_14264,N_7274,N_8356);
and U14265 (N_14265,N_6536,N_9271);
nand U14266 (N_14266,N_8194,N_9932);
nand U14267 (N_14267,N_7683,N_9564);
or U14268 (N_14268,N_6281,N_8708);
or U14269 (N_14269,N_7986,N_8132);
or U14270 (N_14270,N_8779,N_6761);
xor U14271 (N_14271,N_9442,N_7266);
xnor U14272 (N_14272,N_7503,N_6187);
xnor U14273 (N_14273,N_6755,N_7860);
and U14274 (N_14274,N_8065,N_7068);
nand U14275 (N_14275,N_5826,N_6366);
nor U14276 (N_14276,N_5479,N_8747);
nand U14277 (N_14277,N_7650,N_8933);
and U14278 (N_14278,N_8893,N_7419);
and U14279 (N_14279,N_8961,N_5666);
or U14280 (N_14280,N_9209,N_5987);
xnor U14281 (N_14281,N_6866,N_5052);
nor U14282 (N_14282,N_5245,N_6395);
and U14283 (N_14283,N_8276,N_7677);
xor U14284 (N_14284,N_9619,N_7231);
or U14285 (N_14285,N_9328,N_5199);
or U14286 (N_14286,N_5988,N_6147);
and U14287 (N_14287,N_9033,N_8689);
xor U14288 (N_14288,N_5282,N_5156);
nand U14289 (N_14289,N_8055,N_9732);
nor U14290 (N_14290,N_9166,N_6978);
and U14291 (N_14291,N_7273,N_7866);
xnor U14292 (N_14292,N_7796,N_6929);
xor U14293 (N_14293,N_6991,N_8374);
nor U14294 (N_14294,N_8419,N_9575);
and U14295 (N_14295,N_7006,N_7094);
nand U14296 (N_14296,N_8464,N_7709);
xor U14297 (N_14297,N_6564,N_6889);
or U14298 (N_14298,N_6984,N_7226);
nor U14299 (N_14299,N_5670,N_5422);
and U14300 (N_14300,N_6848,N_8479);
or U14301 (N_14301,N_7599,N_9439);
nand U14302 (N_14302,N_7438,N_8700);
or U14303 (N_14303,N_8433,N_9177);
and U14304 (N_14304,N_6401,N_5380);
nand U14305 (N_14305,N_9234,N_8539);
nor U14306 (N_14306,N_6579,N_8833);
and U14307 (N_14307,N_9312,N_5258);
nand U14308 (N_14308,N_5487,N_8550);
nor U14309 (N_14309,N_9278,N_9226);
nor U14310 (N_14310,N_8824,N_8625);
nor U14311 (N_14311,N_5847,N_9673);
or U14312 (N_14312,N_8146,N_7209);
nand U14313 (N_14313,N_5624,N_6640);
nor U14314 (N_14314,N_9021,N_8780);
and U14315 (N_14315,N_8465,N_8358);
or U14316 (N_14316,N_8651,N_8706);
or U14317 (N_14317,N_6018,N_7284);
and U14318 (N_14318,N_9086,N_5544);
or U14319 (N_14319,N_6179,N_5113);
nor U14320 (N_14320,N_9854,N_9041);
xor U14321 (N_14321,N_7898,N_7746);
or U14322 (N_14322,N_6892,N_5235);
or U14323 (N_14323,N_9300,N_7038);
and U14324 (N_14324,N_9230,N_8225);
xnor U14325 (N_14325,N_7187,N_5455);
xor U14326 (N_14326,N_8819,N_8223);
nand U14327 (N_14327,N_7509,N_5743);
nand U14328 (N_14328,N_7259,N_8683);
and U14329 (N_14329,N_9946,N_8676);
xor U14330 (N_14330,N_6096,N_6988);
or U14331 (N_14331,N_5094,N_5026);
or U14332 (N_14332,N_9513,N_5422);
xnor U14333 (N_14333,N_6974,N_5107);
xor U14334 (N_14334,N_7333,N_7974);
or U14335 (N_14335,N_9311,N_5426);
xnor U14336 (N_14336,N_5480,N_9604);
and U14337 (N_14337,N_5301,N_9187);
nor U14338 (N_14338,N_9515,N_7968);
xnor U14339 (N_14339,N_7766,N_9693);
nand U14340 (N_14340,N_6606,N_8428);
and U14341 (N_14341,N_7045,N_9632);
or U14342 (N_14342,N_6172,N_8654);
or U14343 (N_14343,N_9033,N_6336);
nor U14344 (N_14344,N_8680,N_5064);
nand U14345 (N_14345,N_6910,N_6432);
nor U14346 (N_14346,N_6012,N_6975);
xnor U14347 (N_14347,N_7106,N_5001);
nor U14348 (N_14348,N_6066,N_8785);
or U14349 (N_14349,N_6980,N_5405);
xnor U14350 (N_14350,N_6751,N_6201);
nor U14351 (N_14351,N_7683,N_7120);
nand U14352 (N_14352,N_7348,N_7697);
nand U14353 (N_14353,N_7622,N_9737);
nand U14354 (N_14354,N_6063,N_9853);
xor U14355 (N_14355,N_6004,N_7788);
or U14356 (N_14356,N_5006,N_7174);
nor U14357 (N_14357,N_8772,N_8157);
and U14358 (N_14358,N_5085,N_8683);
or U14359 (N_14359,N_5065,N_9071);
nand U14360 (N_14360,N_9936,N_8480);
nor U14361 (N_14361,N_9124,N_8418);
nor U14362 (N_14362,N_6299,N_9877);
nor U14363 (N_14363,N_7014,N_8664);
and U14364 (N_14364,N_7099,N_8112);
and U14365 (N_14365,N_6079,N_8444);
xor U14366 (N_14366,N_9231,N_9824);
nor U14367 (N_14367,N_9061,N_7155);
xnor U14368 (N_14368,N_9256,N_7936);
or U14369 (N_14369,N_9228,N_8387);
or U14370 (N_14370,N_9744,N_8902);
and U14371 (N_14371,N_9697,N_8745);
or U14372 (N_14372,N_8513,N_6716);
nor U14373 (N_14373,N_7814,N_6578);
nand U14374 (N_14374,N_5408,N_5626);
xnor U14375 (N_14375,N_6280,N_5005);
or U14376 (N_14376,N_5814,N_9330);
nand U14377 (N_14377,N_6033,N_7042);
nand U14378 (N_14378,N_8962,N_6194);
and U14379 (N_14379,N_5628,N_8666);
or U14380 (N_14380,N_9848,N_5611);
nand U14381 (N_14381,N_9911,N_8647);
xnor U14382 (N_14382,N_8461,N_8301);
xor U14383 (N_14383,N_6850,N_9375);
or U14384 (N_14384,N_9359,N_8288);
nand U14385 (N_14385,N_7425,N_7668);
or U14386 (N_14386,N_9243,N_8749);
and U14387 (N_14387,N_5869,N_5371);
nand U14388 (N_14388,N_6845,N_9149);
or U14389 (N_14389,N_6847,N_8561);
and U14390 (N_14390,N_7455,N_5891);
or U14391 (N_14391,N_5355,N_8236);
or U14392 (N_14392,N_9840,N_7909);
or U14393 (N_14393,N_8406,N_7401);
xor U14394 (N_14394,N_7555,N_6514);
or U14395 (N_14395,N_9425,N_6663);
and U14396 (N_14396,N_5556,N_5495);
or U14397 (N_14397,N_6134,N_5810);
nand U14398 (N_14398,N_8164,N_7486);
and U14399 (N_14399,N_7725,N_6980);
or U14400 (N_14400,N_9164,N_7439);
or U14401 (N_14401,N_5989,N_5667);
and U14402 (N_14402,N_6867,N_6837);
or U14403 (N_14403,N_7788,N_7185);
or U14404 (N_14404,N_5027,N_8361);
or U14405 (N_14405,N_6265,N_5899);
nand U14406 (N_14406,N_9872,N_6687);
or U14407 (N_14407,N_5136,N_5998);
nor U14408 (N_14408,N_7619,N_8082);
nor U14409 (N_14409,N_8182,N_9699);
nor U14410 (N_14410,N_7239,N_7201);
and U14411 (N_14411,N_5008,N_7674);
and U14412 (N_14412,N_5056,N_8586);
xnor U14413 (N_14413,N_6191,N_8722);
and U14414 (N_14414,N_7132,N_8252);
xor U14415 (N_14415,N_8685,N_5282);
and U14416 (N_14416,N_6627,N_5706);
or U14417 (N_14417,N_8540,N_8829);
nand U14418 (N_14418,N_6674,N_7818);
and U14419 (N_14419,N_9810,N_7157);
and U14420 (N_14420,N_8417,N_9294);
nor U14421 (N_14421,N_8424,N_7686);
nor U14422 (N_14422,N_6798,N_9208);
nand U14423 (N_14423,N_9912,N_7855);
xor U14424 (N_14424,N_5667,N_7648);
and U14425 (N_14425,N_5496,N_7912);
xor U14426 (N_14426,N_6974,N_7488);
nor U14427 (N_14427,N_7299,N_8381);
and U14428 (N_14428,N_9860,N_5988);
nor U14429 (N_14429,N_7762,N_7378);
and U14430 (N_14430,N_6644,N_9018);
or U14431 (N_14431,N_9002,N_8986);
nand U14432 (N_14432,N_8623,N_7579);
and U14433 (N_14433,N_7145,N_7078);
nor U14434 (N_14434,N_7185,N_9959);
nand U14435 (N_14435,N_8161,N_7155);
and U14436 (N_14436,N_7269,N_5401);
nand U14437 (N_14437,N_5427,N_9997);
nor U14438 (N_14438,N_7910,N_5992);
xnor U14439 (N_14439,N_6751,N_7548);
nor U14440 (N_14440,N_7161,N_6006);
nand U14441 (N_14441,N_5992,N_5902);
nor U14442 (N_14442,N_5556,N_5942);
or U14443 (N_14443,N_9046,N_9213);
xor U14444 (N_14444,N_5452,N_6868);
xor U14445 (N_14445,N_7976,N_8038);
and U14446 (N_14446,N_5593,N_8752);
or U14447 (N_14447,N_5013,N_9523);
nor U14448 (N_14448,N_6995,N_5536);
xor U14449 (N_14449,N_9021,N_9851);
and U14450 (N_14450,N_6041,N_7287);
nor U14451 (N_14451,N_7034,N_8516);
or U14452 (N_14452,N_5472,N_9371);
nor U14453 (N_14453,N_9345,N_8346);
or U14454 (N_14454,N_8533,N_6846);
xor U14455 (N_14455,N_9142,N_8380);
xnor U14456 (N_14456,N_8554,N_7792);
nor U14457 (N_14457,N_5154,N_6791);
or U14458 (N_14458,N_8337,N_7823);
xnor U14459 (N_14459,N_7751,N_7668);
nor U14460 (N_14460,N_7454,N_7890);
or U14461 (N_14461,N_8211,N_6179);
nand U14462 (N_14462,N_6502,N_8732);
xor U14463 (N_14463,N_8822,N_7178);
nor U14464 (N_14464,N_5555,N_6026);
nor U14465 (N_14465,N_6158,N_5495);
or U14466 (N_14466,N_6605,N_5278);
nor U14467 (N_14467,N_9391,N_6220);
and U14468 (N_14468,N_6492,N_6659);
nand U14469 (N_14469,N_6170,N_9023);
nand U14470 (N_14470,N_7957,N_5838);
or U14471 (N_14471,N_7540,N_7973);
and U14472 (N_14472,N_9094,N_6653);
or U14473 (N_14473,N_8508,N_9188);
or U14474 (N_14474,N_8157,N_7284);
nor U14475 (N_14475,N_6998,N_5871);
and U14476 (N_14476,N_6377,N_6479);
and U14477 (N_14477,N_8884,N_6700);
or U14478 (N_14478,N_7581,N_8285);
and U14479 (N_14479,N_5439,N_6766);
nand U14480 (N_14480,N_9365,N_8391);
nor U14481 (N_14481,N_6436,N_9587);
and U14482 (N_14482,N_9404,N_7028);
nand U14483 (N_14483,N_5877,N_9097);
and U14484 (N_14484,N_7251,N_8205);
and U14485 (N_14485,N_9562,N_8550);
nor U14486 (N_14486,N_6986,N_5289);
nor U14487 (N_14487,N_6880,N_8447);
nand U14488 (N_14488,N_7575,N_5654);
nand U14489 (N_14489,N_8626,N_7291);
and U14490 (N_14490,N_8999,N_8988);
or U14491 (N_14491,N_9599,N_7335);
nor U14492 (N_14492,N_9637,N_5595);
nor U14493 (N_14493,N_5625,N_8928);
nor U14494 (N_14494,N_6601,N_8460);
and U14495 (N_14495,N_8882,N_8430);
or U14496 (N_14496,N_6144,N_8109);
nor U14497 (N_14497,N_7357,N_6627);
xnor U14498 (N_14498,N_6192,N_8464);
and U14499 (N_14499,N_6939,N_9750);
or U14500 (N_14500,N_5766,N_5447);
and U14501 (N_14501,N_9724,N_7969);
nand U14502 (N_14502,N_8695,N_8387);
xnor U14503 (N_14503,N_9641,N_5153);
or U14504 (N_14504,N_5434,N_7797);
and U14505 (N_14505,N_7722,N_6378);
or U14506 (N_14506,N_9600,N_7082);
xnor U14507 (N_14507,N_5768,N_5832);
and U14508 (N_14508,N_5347,N_6458);
nor U14509 (N_14509,N_7190,N_9977);
or U14510 (N_14510,N_5950,N_6247);
nor U14511 (N_14511,N_6328,N_5124);
and U14512 (N_14512,N_8725,N_6165);
nor U14513 (N_14513,N_8431,N_9096);
nand U14514 (N_14514,N_5479,N_6552);
and U14515 (N_14515,N_5807,N_8279);
or U14516 (N_14516,N_9079,N_7909);
or U14517 (N_14517,N_7541,N_5245);
or U14518 (N_14518,N_7259,N_7880);
nand U14519 (N_14519,N_5351,N_6364);
xor U14520 (N_14520,N_8772,N_8995);
nor U14521 (N_14521,N_5908,N_7660);
nand U14522 (N_14522,N_9612,N_9866);
nand U14523 (N_14523,N_8867,N_6540);
and U14524 (N_14524,N_7854,N_8049);
or U14525 (N_14525,N_9657,N_7745);
nor U14526 (N_14526,N_6018,N_6429);
xnor U14527 (N_14527,N_7219,N_5296);
and U14528 (N_14528,N_8656,N_7613);
and U14529 (N_14529,N_5557,N_9756);
and U14530 (N_14530,N_5063,N_8008);
nor U14531 (N_14531,N_8315,N_6843);
nand U14532 (N_14532,N_7419,N_5337);
nor U14533 (N_14533,N_6064,N_5337);
xnor U14534 (N_14534,N_9922,N_6345);
or U14535 (N_14535,N_8264,N_6052);
xor U14536 (N_14536,N_7106,N_7406);
and U14537 (N_14537,N_9754,N_5731);
and U14538 (N_14538,N_9636,N_8431);
and U14539 (N_14539,N_7006,N_5593);
nor U14540 (N_14540,N_7068,N_9053);
nor U14541 (N_14541,N_7992,N_6584);
and U14542 (N_14542,N_7796,N_7834);
nand U14543 (N_14543,N_7191,N_7365);
xor U14544 (N_14544,N_6805,N_7158);
or U14545 (N_14545,N_9494,N_8200);
xor U14546 (N_14546,N_7913,N_5669);
or U14547 (N_14547,N_6142,N_5718);
nor U14548 (N_14548,N_6103,N_5706);
or U14549 (N_14549,N_6116,N_9927);
and U14550 (N_14550,N_5870,N_8309);
xnor U14551 (N_14551,N_7026,N_5139);
and U14552 (N_14552,N_6825,N_6909);
and U14553 (N_14553,N_6479,N_7642);
and U14554 (N_14554,N_9516,N_9385);
and U14555 (N_14555,N_8175,N_6062);
nand U14556 (N_14556,N_6757,N_5860);
nor U14557 (N_14557,N_5996,N_8920);
or U14558 (N_14558,N_9275,N_9130);
xnor U14559 (N_14559,N_9872,N_5284);
and U14560 (N_14560,N_6567,N_8177);
xnor U14561 (N_14561,N_5426,N_9297);
nand U14562 (N_14562,N_6512,N_8927);
nor U14563 (N_14563,N_9504,N_8483);
xor U14564 (N_14564,N_8116,N_6066);
and U14565 (N_14565,N_9896,N_8196);
or U14566 (N_14566,N_7707,N_5983);
and U14567 (N_14567,N_9048,N_6799);
nor U14568 (N_14568,N_5986,N_6160);
xor U14569 (N_14569,N_8849,N_9301);
xnor U14570 (N_14570,N_5802,N_8373);
and U14571 (N_14571,N_5795,N_9922);
nor U14572 (N_14572,N_7505,N_6408);
nor U14573 (N_14573,N_9582,N_5290);
or U14574 (N_14574,N_7517,N_9654);
and U14575 (N_14575,N_8411,N_9746);
xnor U14576 (N_14576,N_6656,N_5141);
nand U14577 (N_14577,N_7753,N_8222);
nand U14578 (N_14578,N_7318,N_8148);
or U14579 (N_14579,N_5176,N_7564);
xnor U14580 (N_14580,N_9097,N_8692);
nor U14581 (N_14581,N_5159,N_9550);
nor U14582 (N_14582,N_9479,N_8962);
nor U14583 (N_14583,N_6084,N_6384);
and U14584 (N_14584,N_9324,N_7451);
or U14585 (N_14585,N_7487,N_7406);
nor U14586 (N_14586,N_8997,N_6570);
nor U14587 (N_14587,N_9272,N_7162);
or U14588 (N_14588,N_5344,N_9545);
nor U14589 (N_14589,N_8577,N_9945);
nor U14590 (N_14590,N_8858,N_8252);
nand U14591 (N_14591,N_5758,N_6370);
and U14592 (N_14592,N_5547,N_8433);
and U14593 (N_14593,N_5665,N_5072);
xor U14594 (N_14594,N_7102,N_6837);
nor U14595 (N_14595,N_8429,N_8634);
nor U14596 (N_14596,N_6892,N_6566);
nand U14597 (N_14597,N_8120,N_6091);
xor U14598 (N_14598,N_8353,N_8237);
xor U14599 (N_14599,N_8008,N_7085);
nor U14600 (N_14600,N_5120,N_6803);
or U14601 (N_14601,N_7161,N_8389);
and U14602 (N_14602,N_9947,N_7275);
nand U14603 (N_14603,N_7089,N_5008);
nand U14604 (N_14604,N_7862,N_8518);
and U14605 (N_14605,N_7061,N_8002);
xor U14606 (N_14606,N_7136,N_9122);
and U14607 (N_14607,N_8550,N_6066);
or U14608 (N_14608,N_5143,N_6722);
nand U14609 (N_14609,N_8680,N_5267);
nand U14610 (N_14610,N_9101,N_7463);
or U14611 (N_14611,N_6882,N_9002);
and U14612 (N_14612,N_6837,N_5281);
xor U14613 (N_14613,N_6737,N_7719);
or U14614 (N_14614,N_5259,N_6511);
xnor U14615 (N_14615,N_8374,N_9622);
xnor U14616 (N_14616,N_7247,N_7125);
and U14617 (N_14617,N_8801,N_5543);
nor U14618 (N_14618,N_9658,N_6951);
nand U14619 (N_14619,N_5358,N_7414);
and U14620 (N_14620,N_9192,N_9738);
nor U14621 (N_14621,N_7217,N_9449);
nor U14622 (N_14622,N_8195,N_7130);
nand U14623 (N_14623,N_9450,N_8704);
nor U14624 (N_14624,N_7183,N_9318);
xnor U14625 (N_14625,N_5829,N_8051);
nand U14626 (N_14626,N_5949,N_5608);
and U14627 (N_14627,N_5083,N_6003);
xor U14628 (N_14628,N_5835,N_8706);
nor U14629 (N_14629,N_9740,N_5706);
or U14630 (N_14630,N_9742,N_8515);
nor U14631 (N_14631,N_9878,N_7186);
and U14632 (N_14632,N_7705,N_9443);
and U14633 (N_14633,N_6747,N_5777);
nand U14634 (N_14634,N_6218,N_9730);
or U14635 (N_14635,N_7956,N_7521);
and U14636 (N_14636,N_5868,N_6775);
and U14637 (N_14637,N_7906,N_7017);
and U14638 (N_14638,N_7289,N_7487);
and U14639 (N_14639,N_7702,N_7004);
nor U14640 (N_14640,N_6566,N_9019);
or U14641 (N_14641,N_8155,N_9917);
and U14642 (N_14642,N_9546,N_9123);
or U14643 (N_14643,N_8608,N_8882);
nor U14644 (N_14644,N_9706,N_9948);
and U14645 (N_14645,N_8258,N_5305);
nand U14646 (N_14646,N_9820,N_8297);
and U14647 (N_14647,N_5010,N_7463);
or U14648 (N_14648,N_6052,N_6503);
nor U14649 (N_14649,N_7632,N_7122);
or U14650 (N_14650,N_7797,N_8330);
nor U14651 (N_14651,N_5859,N_8461);
xor U14652 (N_14652,N_9272,N_8518);
and U14653 (N_14653,N_9174,N_6723);
nor U14654 (N_14654,N_7690,N_7187);
or U14655 (N_14655,N_5413,N_5193);
or U14656 (N_14656,N_6863,N_8557);
xnor U14657 (N_14657,N_8402,N_8149);
and U14658 (N_14658,N_6105,N_8626);
and U14659 (N_14659,N_5021,N_8847);
nor U14660 (N_14660,N_7888,N_5733);
or U14661 (N_14661,N_6325,N_6204);
nor U14662 (N_14662,N_6058,N_6106);
xor U14663 (N_14663,N_7027,N_6314);
and U14664 (N_14664,N_6439,N_7002);
nand U14665 (N_14665,N_8227,N_6371);
nand U14666 (N_14666,N_5510,N_7136);
nor U14667 (N_14667,N_5080,N_5954);
and U14668 (N_14668,N_9396,N_6101);
xnor U14669 (N_14669,N_9135,N_8569);
and U14670 (N_14670,N_8752,N_5684);
and U14671 (N_14671,N_8343,N_5363);
nand U14672 (N_14672,N_5238,N_5630);
nand U14673 (N_14673,N_8088,N_6453);
nor U14674 (N_14674,N_5964,N_5292);
xor U14675 (N_14675,N_8838,N_7452);
and U14676 (N_14676,N_8972,N_5671);
xnor U14677 (N_14677,N_5684,N_5041);
nand U14678 (N_14678,N_9943,N_6667);
or U14679 (N_14679,N_6031,N_8870);
and U14680 (N_14680,N_5169,N_6876);
or U14681 (N_14681,N_7405,N_6953);
nor U14682 (N_14682,N_6802,N_7982);
xor U14683 (N_14683,N_9192,N_5116);
xnor U14684 (N_14684,N_9269,N_5418);
xor U14685 (N_14685,N_9142,N_7312);
xnor U14686 (N_14686,N_5193,N_9449);
nand U14687 (N_14687,N_9459,N_6109);
or U14688 (N_14688,N_5966,N_5410);
nor U14689 (N_14689,N_5314,N_5284);
and U14690 (N_14690,N_6880,N_5251);
xnor U14691 (N_14691,N_5440,N_8809);
and U14692 (N_14692,N_6170,N_5294);
nand U14693 (N_14693,N_6887,N_7114);
nand U14694 (N_14694,N_8890,N_5156);
or U14695 (N_14695,N_8600,N_7038);
nand U14696 (N_14696,N_7939,N_6099);
xor U14697 (N_14697,N_7634,N_8522);
nand U14698 (N_14698,N_9070,N_6608);
or U14699 (N_14699,N_7099,N_7076);
nor U14700 (N_14700,N_9362,N_9413);
nand U14701 (N_14701,N_9021,N_5082);
or U14702 (N_14702,N_9328,N_9227);
nand U14703 (N_14703,N_7572,N_5404);
and U14704 (N_14704,N_9747,N_5524);
xnor U14705 (N_14705,N_5121,N_8280);
nor U14706 (N_14706,N_7452,N_6458);
or U14707 (N_14707,N_9708,N_7587);
and U14708 (N_14708,N_5888,N_5944);
and U14709 (N_14709,N_9122,N_5417);
and U14710 (N_14710,N_5582,N_9865);
nor U14711 (N_14711,N_8327,N_8390);
or U14712 (N_14712,N_6111,N_8378);
xor U14713 (N_14713,N_9516,N_7409);
xnor U14714 (N_14714,N_7007,N_7380);
or U14715 (N_14715,N_5118,N_7127);
xor U14716 (N_14716,N_5398,N_7092);
and U14717 (N_14717,N_8597,N_7718);
xnor U14718 (N_14718,N_5630,N_8170);
nor U14719 (N_14719,N_5608,N_8268);
and U14720 (N_14720,N_7616,N_6635);
and U14721 (N_14721,N_8051,N_9692);
and U14722 (N_14722,N_7171,N_7439);
and U14723 (N_14723,N_8687,N_7530);
xnor U14724 (N_14724,N_9773,N_9327);
xnor U14725 (N_14725,N_9354,N_7887);
nor U14726 (N_14726,N_7903,N_5741);
and U14727 (N_14727,N_7755,N_8718);
nor U14728 (N_14728,N_9628,N_9886);
xnor U14729 (N_14729,N_5981,N_7879);
xor U14730 (N_14730,N_9639,N_8588);
or U14731 (N_14731,N_6931,N_8197);
nor U14732 (N_14732,N_7098,N_8292);
or U14733 (N_14733,N_7356,N_6316);
nand U14734 (N_14734,N_6965,N_5891);
and U14735 (N_14735,N_9244,N_9888);
and U14736 (N_14736,N_6681,N_9423);
xnor U14737 (N_14737,N_6617,N_6432);
nand U14738 (N_14738,N_7895,N_6472);
xnor U14739 (N_14739,N_9279,N_5190);
and U14740 (N_14740,N_9870,N_5123);
xnor U14741 (N_14741,N_9145,N_5732);
nor U14742 (N_14742,N_5670,N_8175);
and U14743 (N_14743,N_9651,N_8297);
or U14744 (N_14744,N_6004,N_5524);
xor U14745 (N_14745,N_8406,N_9392);
nor U14746 (N_14746,N_9071,N_7678);
nand U14747 (N_14747,N_6254,N_8725);
or U14748 (N_14748,N_5837,N_8505);
and U14749 (N_14749,N_6813,N_8015);
nor U14750 (N_14750,N_5334,N_7576);
xor U14751 (N_14751,N_7886,N_7775);
nand U14752 (N_14752,N_7848,N_7733);
nor U14753 (N_14753,N_6355,N_8703);
nor U14754 (N_14754,N_8925,N_9257);
xor U14755 (N_14755,N_5004,N_9100);
and U14756 (N_14756,N_6965,N_7709);
nand U14757 (N_14757,N_8427,N_6179);
or U14758 (N_14758,N_5027,N_9346);
or U14759 (N_14759,N_5347,N_6270);
and U14760 (N_14760,N_7942,N_6520);
and U14761 (N_14761,N_8427,N_9472);
or U14762 (N_14762,N_5987,N_8771);
nand U14763 (N_14763,N_5568,N_7618);
and U14764 (N_14764,N_6671,N_5298);
xnor U14765 (N_14765,N_8612,N_6923);
or U14766 (N_14766,N_9105,N_8704);
nand U14767 (N_14767,N_9811,N_9711);
xnor U14768 (N_14768,N_9965,N_9725);
nand U14769 (N_14769,N_6059,N_5355);
xor U14770 (N_14770,N_9286,N_7724);
xnor U14771 (N_14771,N_6237,N_7516);
or U14772 (N_14772,N_9088,N_6016);
nand U14773 (N_14773,N_9966,N_7232);
and U14774 (N_14774,N_8609,N_9083);
xor U14775 (N_14775,N_6648,N_9849);
nor U14776 (N_14776,N_6661,N_6672);
xnor U14777 (N_14777,N_6113,N_9586);
nor U14778 (N_14778,N_8700,N_5226);
nor U14779 (N_14779,N_7505,N_7865);
nand U14780 (N_14780,N_6797,N_7095);
nand U14781 (N_14781,N_5987,N_5854);
nand U14782 (N_14782,N_5315,N_8554);
and U14783 (N_14783,N_9266,N_6618);
nor U14784 (N_14784,N_9475,N_9053);
nand U14785 (N_14785,N_7130,N_5067);
nor U14786 (N_14786,N_7850,N_6445);
xor U14787 (N_14787,N_9407,N_9015);
nor U14788 (N_14788,N_8693,N_5893);
and U14789 (N_14789,N_7510,N_6316);
and U14790 (N_14790,N_8565,N_8850);
nor U14791 (N_14791,N_9766,N_7684);
nand U14792 (N_14792,N_6357,N_7051);
and U14793 (N_14793,N_7036,N_5526);
nor U14794 (N_14794,N_6100,N_5066);
and U14795 (N_14795,N_5179,N_9975);
xnor U14796 (N_14796,N_8807,N_7821);
nor U14797 (N_14797,N_6621,N_7912);
and U14798 (N_14798,N_8978,N_6614);
nor U14799 (N_14799,N_7509,N_5804);
nor U14800 (N_14800,N_6441,N_6251);
and U14801 (N_14801,N_5052,N_8370);
nand U14802 (N_14802,N_9599,N_6871);
nor U14803 (N_14803,N_5014,N_8468);
and U14804 (N_14804,N_6218,N_5532);
nor U14805 (N_14805,N_6114,N_7589);
or U14806 (N_14806,N_6696,N_5950);
nand U14807 (N_14807,N_8942,N_5537);
and U14808 (N_14808,N_5811,N_9702);
and U14809 (N_14809,N_5911,N_5374);
or U14810 (N_14810,N_6547,N_9590);
and U14811 (N_14811,N_5989,N_6888);
or U14812 (N_14812,N_5075,N_7189);
or U14813 (N_14813,N_8030,N_8563);
xnor U14814 (N_14814,N_8892,N_8536);
nand U14815 (N_14815,N_8616,N_5588);
xor U14816 (N_14816,N_7460,N_5393);
nand U14817 (N_14817,N_9169,N_6569);
and U14818 (N_14818,N_9747,N_8634);
or U14819 (N_14819,N_9005,N_5844);
and U14820 (N_14820,N_9998,N_9282);
or U14821 (N_14821,N_6723,N_8008);
or U14822 (N_14822,N_6420,N_6739);
nand U14823 (N_14823,N_8010,N_7479);
and U14824 (N_14824,N_7379,N_6049);
xnor U14825 (N_14825,N_8388,N_7493);
xnor U14826 (N_14826,N_8169,N_9883);
xor U14827 (N_14827,N_6485,N_9572);
or U14828 (N_14828,N_8182,N_9254);
nor U14829 (N_14829,N_6984,N_9779);
nor U14830 (N_14830,N_7735,N_9301);
nand U14831 (N_14831,N_7997,N_7834);
xnor U14832 (N_14832,N_6674,N_6314);
nand U14833 (N_14833,N_6022,N_9485);
nor U14834 (N_14834,N_7629,N_7835);
nand U14835 (N_14835,N_5669,N_5021);
nor U14836 (N_14836,N_6996,N_6081);
nor U14837 (N_14837,N_7729,N_7618);
nor U14838 (N_14838,N_7055,N_9760);
and U14839 (N_14839,N_6356,N_6126);
nor U14840 (N_14840,N_8895,N_7305);
and U14841 (N_14841,N_7690,N_5248);
nor U14842 (N_14842,N_5602,N_8551);
and U14843 (N_14843,N_9014,N_7874);
and U14844 (N_14844,N_9927,N_9387);
or U14845 (N_14845,N_6533,N_7486);
xnor U14846 (N_14846,N_7679,N_7811);
and U14847 (N_14847,N_5591,N_9333);
or U14848 (N_14848,N_8577,N_9349);
or U14849 (N_14849,N_5240,N_9548);
or U14850 (N_14850,N_8903,N_9209);
and U14851 (N_14851,N_8582,N_6899);
nor U14852 (N_14852,N_5503,N_8849);
and U14853 (N_14853,N_5320,N_7654);
nand U14854 (N_14854,N_6919,N_9197);
and U14855 (N_14855,N_9524,N_9255);
and U14856 (N_14856,N_9933,N_6072);
nand U14857 (N_14857,N_5663,N_9663);
nor U14858 (N_14858,N_7053,N_8996);
nor U14859 (N_14859,N_8301,N_6522);
nor U14860 (N_14860,N_6835,N_8234);
xnor U14861 (N_14861,N_9326,N_8023);
or U14862 (N_14862,N_6611,N_7085);
xnor U14863 (N_14863,N_6023,N_6345);
xnor U14864 (N_14864,N_8707,N_8602);
nand U14865 (N_14865,N_7527,N_8070);
and U14866 (N_14866,N_7991,N_8121);
nor U14867 (N_14867,N_7420,N_7674);
nor U14868 (N_14868,N_7085,N_5415);
and U14869 (N_14869,N_9469,N_6371);
nand U14870 (N_14870,N_6869,N_9066);
or U14871 (N_14871,N_7890,N_8904);
nand U14872 (N_14872,N_9854,N_7082);
or U14873 (N_14873,N_6025,N_5122);
xnor U14874 (N_14874,N_8624,N_8197);
nand U14875 (N_14875,N_9053,N_5259);
nor U14876 (N_14876,N_5526,N_9541);
and U14877 (N_14877,N_8967,N_8085);
xor U14878 (N_14878,N_9644,N_9082);
or U14879 (N_14879,N_9562,N_7427);
nor U14880 (N_14880,N_7713,N_6724);
or U14881 (N_14881,N_7063,N_9488);
xor U14882 (N_14882,N_7070,N_7489);
or U14883 (N_14883,N_5601,N_8750);
xnor U14884 (N_14884,N_9684,N_6198);
and U14885 (N_14885,N_9427,N_8948);
nor U14886 (N_14886,N_7857,N_6917);
or U14887 (N_14887,N_5639,N_8748);
nor U14888 (N_14888,N_6092,N_8206);
nand U14889 (N_14889,N_5362,N_7001);
nand U14890 (N_14890,N_7116,N_7025);
nor U14891 (N_14891,N_6732,N_9870);
xnor U14892 (N_14892,N_5542,N_8954);
nand U14893 (N_14893,N_7903,N_7637);
xnor U14894 (N_14894,N_9585,N_6692);
and U14895 (N_14895,N_5355,N_7414);
xor U14896 (N_14896,N_5015,N_6789);
nand U14897 (N_14897,N_5851,N_5010);
nand U14898 (N_14898,N_6662,N_5270);
xnor U14899 (N_14899,N_6444,N_9326);
xor U14900 (N_14900,N_7466,N_8025);
nor U14901 (N_14901,N_5183,N_9230);
and U14902 (N_14902,N_6295,N_5489);
nor U14903 (N_14903,N_5157,N_7888);
nand U14904 (N_14904,N_9886,N_5208);
nand U14905 (N_14905,N_6951,N_8424);
or U14906 (N_14906,N_8766,N_8459);
nand U14907 (N_14907,N_8251,N_5911);
nand U14908 (N_14908,N_8750,N_6366);
and U14909 (N_14909,N_8451,N_9674);
or U14910 (N_14910,N_5822,N_6176);
nor U14911 (N_14911,N_6799,N_9126);
and U14912 (N_14912,N_5812,N_6725);
xor U14913 (N_14913,N_5304,N_6300);
xor U14914 (N_14914,N_9970,N_7021);
and U14915 (N_14915,N_8729,N_9415);
xnor U14916 (N_14916,N_8003,N_8694);
nand U14917 (N_14917,N_9283,N_8116);
xor U14918 (N_14918,N_8771,N_6492);
nor U14919 (N_14919,N_9977,N_8862);
and U14920 (N_14920,N_7753,N_7197);
nor U14921 (N_14921,N_9787,N_5324);
xnor U14922 (N_14922,N_8976,N_8643);
or U14923 (N_14923,N_9830,N_6778);
and U14924 (N_14924,N_9793,N_7552);
nor U14925 (N_14925,N_7437,N_5677);
xor U14926 (N_14926,N_8396,N_6382);
nor U14927 (N_14927,N_6738,N_5411);
xnor U14928 (N_14928,N_7277,N_5865);
nor U14929 (N_14929,N_6519,N_9738);
nor U14930 (N_14930,N_8717,N_7695);
nor U14931 (N_14931,N_5947,N_8045);
nand U14932 (N_14932,N_8539,N_5181);
and U14933 (N_14933,N_6297,N_8838);
nand U14934 (N_14934,N_5314,N_5409);
nor U14935 (N_14935,N_5328,N_7625);
nor U14936 (N_14936,N_6468,N_8742);
or U14937 (N_14937,N_8227,N_8225);
or U14938 (N_14938,N_7308,N_7753);
nor U14939 (N_14939,N_8610,N_5631);
xor U14940 (N_14940,N_6097,N_7620);
nor U14941 (N_14941,N_8577,N_8206);
or U14942 (N_14942,N_8846,N_5802);
xnor U14943 (N_14943,N_5163,N_5748);
nand U14944 (N_14944,N_7865,N_8230);
or U14945 (N_14945,N_9021,N_5243);
or U14946 (N_14946,N_9833,N_9888);
and U14947 (N_14947,N_8245,N_9125);
xnor U14948 (N_14948,N_8351,N_9583);
nor U14949 (N_14949,N_9431,N_7595);
and U14950 (N_14950,N_6015,N_8470);
and U14951 (N_14951,N_7624,N_8145);
nand U14952 (N_14952,N_5214,N_5535);
or U14953 (N_14953,N_8925,N_8545);
and U14954 (N_14954,N_9906,N_7780);
nor U14955 (N_14955,N_9480,N_8608);
and U14956 (N_14956,N_8350,N_9025);
and U14957 (N_14957,N_6875,N_5880);
nor U14958 (N_14958,N_7106,N_6322);
xor U14959 (N_14959,N_6061,N_8977);
and U14960 (N_14960,N_8732,N_8314);
nand U14961 (N_14961,N_8633,N_5359);
xor U14962 (N_14962,N_8174,N_7786);
or U14963 (N_14963,N_6477,N_8235);
and U14964 (N_14964,N_9693,N_5745);
or U14965 (N_14965,N_6429,N_6706);
xnor U14966 (N_14966,N_9675,N_8321);
or U14967 (N_14967,N_9334,N_9291);
nand U14968 (N_14968,N_6758,N_8621);
or U14969 (N_14969,N_8269,N_8631);
or U14970 (N_14970,N_7855,N_7298);
nand U14971 (N_14971,N_9923,N_8946);
nand U14972 (N_14972,N_9115,N_5463);
and U14973 (N_14973,N_9806,N_9987);
and U14974 (N_14974,N_7160,N_6879);
and U14975 (N_14975,N_7937,N_7691);
or U14976 (N_14976,N_5234,N_9471);
or U14977 (N_14977,N_6151,N_5610);
or U14978 (N_14978,N_7638,N_5385);
and U14979 (N_14979,N_5233,N_5952);
xnor U14980 (N_14980,N_5769,N_9735);
xor U14981 (N_14981,N_6381,N_9534);
xor U14982 (N_14982,N_7816,N_6934);
nor U14983 (N_14983,N_6948,N_7401);
nand U14984 (N_14984,N_7450,N_8178);
and U14985 (N_14985,N_9901,N_9193);
or U14986 (N_14986,N_7947,N_8745);
nand U14987 (N_14987,N_5387,N_5339);
xor U14988 (N_14988,N_9259,N_5607);
and U14989 (N_14989,N_9147,N_9258);
or U14990 (N_14990,N_6347,N_7003);
nor U14991 (N_14991,N_6278,N_7135);
nor U14992 (N_14992,N_7681,N_8253);
nor U14993 (N_14993,N_9399,N_5971);
nor U14994 (N_14994,N_9936,N_8977);
nand U14995 (N_14995,N_7361,N_5643);
and U14996 (N_14996,N_8532,N_8508);
nor U14997 (N_14997,N_9253,N_8944);
nand U14998 (N_14998,N_5376,N_8233);
or U14999 (N_14999,N_6720,N_9756);
nand UO_0 (O_0,N_12534,N_10013);
xnor UO_1 (O_1,N_13911,N_13636);
nor UO_2 (O_2,N_10432,N_13460);
xnor UO_3 (O_3,N_10969,N_12745);
or UO_4 (O_4,N_13200,N_10728);
nand UO_5 (O_5,N_14206,N_13512);
nor UO_6 (O_6,N_12006,N_12143);
nor UO_7 (O_7,N_14750,N_12062);
xor UO_8 (O_8,N_10441,N_12223);
or UO_9 (O_9,N_13906,N_12997);
xnor UO_10 (O_10,N_14880,N_10972);
or UO_11 (O_11,N_11950,N_11681);
nand UO_12 (O_12,N_12501,N_14705);
nand UO_13 (O_13,N_14566,N_12860);
nor UO_14 (O_14,N_10708,N_13265);
and UO_15 (O_15,N_11511,N_12587);
nor UO_16 (O_16,N_10403,N_12355);
or UO_17 (O_17,N_10007,N_13195);
nand UO_18 (O_18,N_13309,N_11477);
nand UO_19 (O_19,N_13376,N_11402);
or UO_20 (O_20,N_13802,N_10517);
nor UO_21 (O_21,N_12700,N_10292);
or UO_22 (O_22,N_14169,N_11556);
and UO_23 (O_23,N_11945,N_11342);
nor UO_24 (O_24,N_10743,N_10706);
nand UO_25 (O_25,N_12987,N_14247);
or UO_26 (O_26,N_11914,N_13204);
nor UO_27 (O_27,N_10340,N_10511);
or UO_28 (O_28,N_10316,N_10508);
xor UO_29 (O_29,N_12640,N_14622);
nand UO_30 (O_30,N_13100,N_11958);
nand UO_31 (O_31,N_11221,N_11916);
xor UO_32 (O_32,N_11863,N_10137);
or UO_33 (O_33,N_14690,N_14198);
or UO_34 (O_34,N_10850,N_12118);
and UO_35 (O_35,N_12418,N_12089);
and UO_36 (O_36,N_10243,N_11016);
and UO_37 (O_37,N_13050,N_11057);
and UO_38 (O_38,N_13875,N_13912);
and UO_39 (O_39,N_13584,N_11039);
nor UO_40 (O_40,N_14852,N_10874);
or UO_41 (O_41,N_13697,N_13217);
or UO_42 (O_42,N_14898,N_10592);
nand UO_43 (O_43,N_13463,N_13448);
xnor UO_44 (O_44,N_13720,N_13535);
xnor UO_45 (O_45,N_14636,N_13879);
and UO_46 (O_46,N_13898,N_12622);
nor UO_47 (O_47,N_13729,N_14351);
or UO_48 (O_48,N_13160,N_10773);
xor UO_49 (O_49,N_14882,N_10388);
or UO_50 (O_50,N_12232,N_13179);
or UO_51 (O_51,N_13450,N_14340);
or UO_52 (O_52,N_14902,N_14034);
nor UO_53 (O_53,N_14330,N_11272);
nor UO_54 (O_54,N_12486,N_12742);
or UO_55 (O_55,N_12609,N_13829);
nand UO_56 (O_56,N_12617,N_11033);
or UO_57 (O_57,N_10930,N_14248);
nor UO_58 (O_58,N_13387,N_14051);
nor UO_59 (O_59,N_12036,N_10157);
xor UO_60 (O_60,N_14010,N_13411);
nor UO_61 (O_61,N_14105,N_14478);
nand UO_62 (O_62,N_14407,N_13730);
nor UO_63 (O_63,N_10631,N_14551);
nor UO_64 (O_64,N_11220,N_12721);
nor UO_65 (O_65,N_12309,N_12950);
or UO_66 (O_66,N_13055,N_10430);
nor UO_67 (O_67,N_14672,N_14396);
nor UO_68 (O_68,N_14254,N_10778);
xnor UO_69 (O_69,N_14976,N_13023);
nor UO_70 (O_70,N_12770,N_11411);
nand UO_71 (O_71,N_11806,N_11529);
and UO_72 (O_72,N_12560,N_11454);
xnor UO_73 (O_73,N_11331,N_13190);
xnor UO_74 (O_74,N_12951,N_12209);
and UO_75 (O_75,N_13336,N_10270);
nor UO_76 (O_76,N_10088,N_11508);
and UO_77 (O_77,N_12333,N_10181);
or UO_78 (O_78,N_11755,N_14968);
xor UO_79 (O_79,N_12903,N_14320);
nor UO_80 (O_80,N_10990,N_13375);
nor UO_81 (O_81,N_10087,N_13981);
and UO_82 (O_82,N_12169,N_14332);
xor UO_83 (O_83,N_10822,N_14743);
or UO_84 (O_84,N_14797,N_12673);
and UO_85 (O_85,N_13944,N_14932);
xnor UO_86 (O_86,N_12962,N_14553);
and UO_87 (O_87,N_12017,N_10456);
and UO_88 (O_88,N_11191,N_14655);
and UO_89 (O_89,N_11791,N_11427);
or UO_90 (O_90,N_14244,N_12641);
or UO_91 (O_91,N_12156,N_14853);
xnor UO_92 (O_92,N_10010,N_10703);
nand UO_93 (O_93,N_12170,N_10279);
and UO_94 (O_94,N_14303,N_10101);
xnor UO_95 (O_95,N_10847,N_10645);
and UO_96 (O_96,N_10431,N_14980);
nand UO_97 (O_97,N_12286,N_13503);
nor UO_98 (O_98,N_13082,N_14460);
nand UO_99 (O_99,N_12329,N_10956);
xor UO_100 (O_100,N_14466,N_13124);
and UO_101 (O_101,N_12595,N_11086);
xor UO_102 (O_102,N_10662,N_10494);
and UO_103 (O_103,N_14663,N_14574);
or UO_104 (O_104,N_14139,N_13841);
and UO_105 (O_105,N_13533,N_11350);
xor UO_106 (O_106,N_14038,N_10147);
or UO_107 (O_107,N_13915,N_14579);
nor UO_108 (O_108,N_12973,N_13806);
nor UO_109 (O_109,N_14547,N_11224);
xor UO_110 (O_110,N_10421,N_12417);
nand UO_111 (O_111,N_11678,N_11134);
and UO_112 (O_112,N_12437,N_11912);
or UO_113 (O_113,N_10786,N_11404);
nor UO_114 (O_114,N_14243,N_11462);
nor UO_115 (O_115,N_14219,N_12436);
nand UO_116 (O_116,N_12855,N_10218);
xor UO_117 (O_117,N_14421,N_11621);
nand UO_118 (O_118,N_10813,N_12849);
nor UO_119 (O_119,N_13905,N_11204);
or UO_120 (O_120,N_14997,N_14215);
nand UO_121 (O_121,N_11267,N_14720);
nor UO_122 (O_122,N_14497,N_12723);
nor UO_123 (O_123,N_12872,N_13703);
xor UO_124 (O_124,N_12352,N_14369);
xnor UO_125 (O_125,N_12033,N_14052);
or UO_126 (O_126,N_13855,N_12422);
and UO_127 (O_127,N_10638,N_11029);
nand UO_128 (O_128,N_13894,N_12384);
nand UO_129 (O_129,N_14752,N_14209);
xor UO_130 (O_130,N_10378,N_13285);
or UO_131 (O_131,N_10372,N_11734);
nor UO_132 (O_132,N_14920,N_13184);
or UO_133 (O_133,N_13304,N_12345);
and UO_134 (O_134,N_14744,N_10986);
nor UO_135 (O_135,N_14132,N_10958);
or UO_136 (O_136,N_14072,N_10361);
xor UO_137 (O_137,N_12784,N_12407);
or UO_138 (O_138,N_12387,N_11689);
or UO_139 (O_139,N_11657,N_11175);
and UO_140 (O_140,N_12161,N_10798);
or UO_141 (O_141,N_11260,N_14176);
or UO_142 (O_142,N_14003,N_10892);
nor UO_143 (O_143,N_12935,N_13197);
xor UO_144 (O_144,N_14097,N_13850);
and UO_145 (O_145,N_14609,N_12293);
xnor UO_146 (O_146,N_13986,N_12777);
nor UO_147 (O_147,N_14395,N_13079);
nand UO_148 (O_148,N_14266,N_12618);
xor UO_149 (O_149,N_11491,N_10161);
xor UO_150 (O_150,N_10452,N_12996);
nor UO_151 (O_151,N_14722,N_10072);
nor UO_152 (O_152,N_10675,N_10830);
and UO_153 (O_153,N_11707,N_13144);
and UO_154 (O_154,N_11960,N_12659);
xor UO_155 (O_155,N_14725,N_11962);
and UO_156 (O_156,N_10203,N_13340);
or UO_157 (O_157,N_13145,N_14403);
or UO_158 (O_158,N_13102,N_11605);
nor UO_159 (O_159,N_12416,N_11417);
nor UO_160 (O_160,N_14681,N_12061);
or UO_161 (O_161,N_14154,N_12221);
nand UO_162 (O_162,N_13837,N_10916);
xnor UO_163 (O_163,N_14045,N_13922);
nand UO_164 (O_164,N_10647,N_13598);
xnor UO_165 (O_165,N_10887,N_10941);
or UO_166 (O_166,N_12492,N_12994);
nand UO_167 (O_167,N_14513,N_13410);
nor UO_168 (O_168,N_14041,N_12029);
or UO_169 (O_169,N_12471,N_10621);
nor UO_170 (O_170,N_13616,N_11860);
xor UO_171 (O_171,N_10780,N_11751);
and UO_172 (O_172,N_10955,N_12869);
or UO_173 (O_173,N_11559,N_12612);
nor UO_174 (O_174,N_13008,N_13267);
or UO_175 (O_175,N_12045,N_13360);
xnor UO_176 (O_176,N_13115,N_12095);
and UO_177 (O_177,N_10192,N_11059);
and UO_178 (O_178,N_13007,N_14799);
nand UO_179 (O_179,N_11816,N_10918);
nor UO_180 (O_180,N_14572,N_12980);
and UO_181 (O_181,N_13576,N_14433);
xnor UO_182 (O_182,N_10410,N_11058);
and UO_183 (O_183,N_11453,N_14270);
and UO_184 (O_184,N_11773,N_10398);
or UO_185 (O_185,N_10834,N_11156);
nor UO_186 (O_186,N_11470,N_14149);
nand UO_187 (O_187,N_11359,N_14761);
nand UO_188 (O_188,N_11194,N_11155);
or UO_189 (O_189,N_11984,N_13457);
nor UO_190 (O_190,N_10802,N_12875);
nor UO_191 (O_191,N_11262,N_10457);
and UO_192 (O_192,N_10545,N_10596);
or UO_193 (O_193,N_13126,N_11149);
and UO_194 (O_194,N_13796,N_14226);
nor UO_195 (O_195,N_11518,N_12496);
and UO_196 (O_196,N_10745,N_10284);
or UO_197 (O_197,N_13538,N_10566);
nand UO_198 (O_198,N_14739,N_13751);
nand UO_199 (O_199,N_13715,N_14930);
and UO_200 (O_200,N_12172,N_14952);
nand UO_201 (O_201,N_10439,N_14240);
nand UO_202 (O_202,N_11167,N_13578);
and UO_203 (O_203,N_14781,N_11954);
and UO_204 (O_204,N_13579,N_10746);
and UO_205 (O_205,N_11612,N_14691);
or UO_206 (O_206,N_10559,N_14514);
xnor UO_207 (O_207,N_12893,N_11132);
nand UO_208 (O_208,N_12635,N_10362);
and UO_209 (O_209,N_12000,N_14378);
or UO_210 (O_210,N_13640,N_12445);
nor UO_211 (O_211,N_14211,N_14485);
nand UO_212 (O_212,N_10227,N_10648);
xor UO_213 (O_213,N_10384,N_13635);
xor UO_214 (O_214,N_12904,N_10864);
nand UO_215 (O_215,N_13633,N_11487);
nand UO_216 (O_216,N_14987,N_10843);
or UO_217 (O_217,N_12772,N_11759);
or UO_218 (O_218,N_10556,N_12597);
or UO_219 (O_219,N_13081,N_13771);
or UO_220 (O_220,N_11946,N_11205);
or UO_221 (O_221,N_10032,N_12569);
nand UO_222 (O_222,N_13948,N_13878);
and UO_223 (O_223,N_10784,N_14949);
or UO_224 (O_224,N_14922,N_14981);
or UO_225 (O_225,N_14893,N_13994);
or UO_226 (O_226,N_13191,N_13990);
xor UO_227 (O_227,N_10055,N_12555);
xor UO_228 (O_228,N_10018,N_10070);
nand UO_229 (O_229,N_14391,N_12755);
nor UO_230 (O_230,N_12726,N_12761);
nand UO_231 (O_231,N_10985,N_10390);
and UO_232 (O_232,N_12021,N_11679);
nand UO_233 (O_233,N_11226,N_10411);
nor UO_234 (O_234,N_13580,N_13355);
nor UO_235 (O_235,N_11360,N_11070);
nor UO_236 (O_236,N_11300,N_13332);
and UO_237 (O_237,N_14608,N_14540);
nand UO_238 (O_238,N_10610,N_14941);
or UO_239 (O_239,N_12245,N_11721);
and UO_240 (O_240,N_10711,N_12028);
nand UO_241 (O_241,N_10296,N_11624);
or UO_242 (O_242,N_14163,N_11739);
and UO_243 (O_243,N_13161,N_14680);
nand UO_244 (O_244,N_12094,N_12141);
and UO_245 (O_245,N_12923,N_12414);
xnor UO_246 (O_246,N_14212,N_13775);
nor UO_247 (O_247,N_12799,N_12827);
nor UO_248 (O_248,N_14780,N_14625);
and UO_249 (O_249,N_10505,N_11310);
nand UO_250 (O_250,N_14310,N_13478);
nand UO_251 (O_251,N_14683,N_14315);
nor UO_252 (O_252,N_11646,N_14385);
and UO_253 (O_253,N_13617,N_13741);
or UO_254 (O_254,N_10526,N_11436);
xor UO_255 (O_255,N_11562,N_13090);
nand UO_256 (O_256,N_11826,N_14900);
nor UO_257 (O_257,N_14471,N_11422);
or UO_258 (O_258,N_10193,N_11222);
nand UO_259 (O_259,N_11050,N_13354);
nand UO_260 (O_260,N_13298,N_13242);
or UO_261 (O_261,N_13627,N_11682);
nor UO_262 (O_262,N_13388,N_10568);
and UO_263 (O_263,N_10067,N_13809);
and UO_264 (O_264,N_13089,N_13210);
nand UO_265 (O_265,N_10344,N_12203);
and UO_266 (O_266,N_14520,N_10380);
or UO_267 (O_267,N_12984,N_12009);
or UO_268 (O_268,N_10913,N_13710);
nand UO_269 (O_269,N_14665,N_14058);
nand UO_270 (O_270,N_12714,N_12918);
nor UO_271 (O_271,N_12007,N_13726);
and UO_272 (O_272,N_14620,N_12362);
or UO_273 (O_273,N_14737,N_13546);
and UO_274 (O_274,N_13504,N_10179);
and UO_275 (O_275,N_12800,N_10819);
nor UO_276 (O_276,N_11644,N_11534);
nor UO_277 (O_277,N_12686,N_14762);
or UO_278 (O_278,N_11838,N_14441);
nand UO_279 (O_279,N_10690,N_11466);
nand UO_280 (O_280,N_14974,N_11928);
nor UO_281 (O_281,N_14819,N_13493);
or UO_282 (O_282,N_13394,N_10661);
nand UO_283 (O_283,N_10471,N_13468);
or UO_284 (O_284,N_13469,N_12016);
nor UO_285 (O_285,N_11522,N_11504);
nor UO_286 (O_286,N_13446,N_10434);
or UO_287 (O_287,N_11842,N_12544);
nand UO_288 (O_288,N_11120,N_14584);
or UO_289 (O_289,N_11372,N_11238);
xnor UO_290 (O_290,N_10710,N_11066);
xnor UO_291 (O_291,N_12303,N_12024);
and UO_292 (O_292,N_13541,N_11645);
and UO_293 (O_293,N_12656,N_10106);
nand UO_294 (O_294,N_11365,N_12991);
nand UO_295 (O_295,N_14302,N_11715);
and UO_296 (O_296,N_13122,N_10730);
nor UO_297 (O_297,N_14488,N_12732);
nand UO_298 (O_298,N_14530,N_12562);
and UO_299 (O_299,N_12535,N_14029);
nor UO_300 (O_300,N_10182,N_10386);
and UO_301 (O_301,N_10170,N_10250);
nand UO_302 (O_302,N_13947,N_14617);
nor UO_303 (O_303,N_12351,N_10537);
nand UO_304 (O_304,N_14353,N_14641);
nand UO_305 (O_305,N_14552,N_10107);
or UO_306 (O_306,N_13863,N_13490);
nand UO_307 (O_307,N_13816,N_13682);
or UO_308 (O_308,N_10435,N_13329);
nor UO_309 (O_309,N_14603,N_13700);
nand UO_310 (O_310,N_11209,N_13568);
or UO_311 (O_311,N_12528,N_12696);
and UO_312 (O_312,N_13315,N_12750);
and UO_313 (O_313,N_14063,N_11037);
nand UO_314 (O_314,N_14365,N_12411);
nor UO_315 (O_315,N_12782,N_10602);
and UO_316 (O_316,N_13626,N_12294);
nor UO_317 (O_317,N_12888,N_11836);
nor UO_318 (O_318,N_11699,N_10160);
nand UO_319 (O_319,N_10153,N_12960);
and UO_320 (O_320,N_11391,N_11936);
xnor UO_321 (O_321,N_13107,N_12039);
or UO_322 (O_322,N_13880,N_12003);
nand UO_323 (O_323,N_12490,N_12249);
nor UO_324 (O_324,N_12572,N_12119);
nand UO_325 (O_325,N_10809,N_14145);
xor UO_326 (O_326,N_11151,N_10190);
nand UO_327 (O_327,N_12503,N_11351);
and UO_328 (O_328,N_10350,N_12529);
nor UO_329 (O_329,N_12790,N_11561);
nand UO_330 (O_330,N_14524,N_11778);
nor UO_331 (O_331,N_10130,N_13744);
xor UO_332 (O_332,N_11676,N_14660);
or UO_333 (O_333,N_13348,N_10333);
or UO_334 (O_334,N_13241,N_11097);
xnor UO_335 (O_335,N_14137,N_10723);
and UO_336 (O_336,N_10507,N_11203);
xor UO_337 (O_337,N_10673,N_13672);
or UO_338 (O_338,N_14727,N_10712);
nor UO_339 (O_339,N_10173,N_10852);
xnor UO_340 (O_340,N_13754,N_11880);
nor UO_341 (O_341,N_13694,N_12464);
or UO_342 (O_342,N_10312,N_13545);
nand UO_343 (O_343,N_14426,N_13689);
nand UO_344 (O_344,N_13068,N_10205);
nand UO_345 (O_345,N_12959,N_13371);
and UO_346 (O_346,N_13372,N_12844);
nor UO_347 (O_347,N_11975,N_13936);
nand UO_348 (O_348,N_11420,N_12479);
or UO_349 (O_349,N_13508,N_10577);
xor UO_350 (O_350,N_10939,N_10565);
nand UO_351 (O_351,N_14951,N_11512);
or UO_352 (O_352,N_10607,N_13901);
nand UO_353 (O_353,N_12508,N_12914);
nand UO_354 (O_354,N_11396,N_11613);
xnor UO_355 (O_355,N_12727,N_12852);
nor UO_356 (O_356,N_12706,N_12956);
or UO_357 (O_357,N_10014,N_10394);
or UO_358 (O_358,N_14467,N_10628);
and UO_359 (O_359,N_10073,N_11237);
and UO_360 (O_360,N_14228,N_11869);
xor UO_361 (O_361,N_10623,N_12453);
xnor UO_362 (O_362,N_12381,N_11076);
xnor UO_363 (O_363,N_14808,N_12709);
nor UO_364 (O_364,N_12671,N_10321);
or UO_365 (O_365,N_10796,N_12026);
and UO_366 (O_366,N_14972,N_13839);
nor UO_367 (O_367,N_12531,N_11733);
nand UO_368 (O_368,N_14592,N_12967);
and UO_369 (O_369,N_11324,N_11782);
xor UO_370 (O_370,N_13657,N_12275);
xor UO_371 (O_371,N_14025,N_13042);
xor UO_372 (O_372,N_14841,N_12821);
xor UO_373 (O_373,N_12695,N_11851);
or UO_374 (O_374,N_11179,N_11547);
nand UO_375 (O_375,N_10683,N_12741);
or UO_376 (O_376,N_12301,N_13641);
or UO_377 (O_377,N_12248,N_14084);
xnor UO_378 (O_378,N_14943,N_11007);
nand UO_379 (O_379,N_14148,N_13029);
xnor UO_380 (O_380,N_10324,N_14656);
or UO_381 (O_381,N_11948,N_12069);
nor UO_382 (O_382,N_12071,N_12968);
nor UO_383 (O_383,N_14580,N_12715);
or UO_384 (O_384,N_13464,N_13756);
nand UO_385 (O_385,N_10021,N_12005);
xnor UO_386 (O_386,N_11075,N_12720);
and UO_387 (O_387,N_14831,N_11135);
nor UO_388 (O_388,N_11760,N_12198);
nand UO_389 (O_389,N_12150,N_12603);
nand UO_390 (O_390,N_12791,N_14837);
nor UO_391 (O_391,N_10208,N_12495);
xor UO_392 (O_392,N_14939,N_12585);
nor UO_393 (O_393,N_14101,N_11463);
nand UO_394 (O_394,N_12808,N_13249);
and UO_395 (O_395,N_13516,N_12051);
xnor UO_396 (O_396,N_12912,N_12269);
xor UO_397 (O_397,N_14954,N_11458);
nor UO_398 (O_398,N_10256,N_10370);
and UO_399 (O_399,N_14419,N_12180);
nor UO_400 (O_400,N_12015,N_14869);
nand UO_401 (O_401,N_10653,N_10027);
or UO_402 (O_402,N_14521,N_13582);
nor UO_403 (O_403,N_12604,N_11514);
or UO_404 (O_404,N_11978,N_12060);
or UO_405 (O_405,N_12815,N_10831);
nand UO_406 (O_406,N_14963,N_12055);
xnor UO_407 (O_407,N_12450,N_11357);
xnor UO_408 (O_408,N_14539,N_10849);
or UO_409 (O_409,N_13571,N_10385);
nand UO_410 (O_410,N_10950,N_11526);
nand UO_411 (O_411,N_12056,N_12242);
nand UO_412 (O_412,N_13403,N_12974);
nand UO_413 (O_413,N_10853,N_10231);
xnor UO_414 (O_414,N_13345,N_14892);
and UO_415 (O_415,N_13440,N_11459);
and UO_416 (O_416,N_14926,N_10082);
nor UO_417 (O_417,N_12979,N_10151);
and UO_418 (O_418,N_14515,N_13383);
xnor UO_419 (O_419,N_11115,N_13175);
nor UO_420 (O_420,N_12273,N_14158);
nor UO_421 (O_421,N_14109,N_10294);
xor UO_422 (O_422,N_10988,N_14510);
nor UO_423 (O_423,N_11369,N_11874);
nand UO_424 (O_424,N_14545,N_11278);
xor UO_425 (O_425,N_13436,N_12022);
xnor UO_426 (O_426,N_12554,N_10999);
and UO_427 (O_427,N_14785,N_11905);
nor UO_428 (O_428,N_13350,N_14777);
or UO_429 (O_429,N_10981,N_14208);
xnor UO_430 (O_430,N_11544,N_14754);
nor UO_431 (O_431,N_13442,N_14334);
nor UO_432 (O_432,N_13873,N_13224);
or UO_433 (O_433,N_10845,N_11192);
and UO_434 (O_434,N_12530,N_11498);
nor UO_435 (O_435,N_11253,N_11346);
nand UO_436 (O_436,N_14559,N_10677);
or UO_437 (O_437,N_14590,N_14418);
and UO_438 (O_438,N_12404,N_13262);
nor UO_439 (O_439,N_12219,N_11617);
xor UO_440 (O_440,N_10169,N_13114);
and UO_441 (O_441,N_10866,N_11440);
nor UO_442 (O_442,N_10948,N_13595);
nor UO_443 (O_443,N_10469,N_11768);
nand UO_444 (O_444,N_13892,N_12499);
or UO_445 (O_445,N_14278,N_14912);
nor UO_446 (O_446,N_13566,N_10081);
nand UO_447 (O_447,N_11341,N_10038);
nor UO_448 (O_448,N_10929,N_12227);
xnor UO_449 (O_449,N_13473,N_13495);
and UO_450 (O_450,N_10571,N_11152);
nand UO_451 (O_451,N_14253,N_11393);
xor UO_452 (O_452,N_10925,N_13946);
and UO_453 (O_453,N_11071,N_12929);
nand UO_454 (O_454,N_13011,N_13086);
nor UO_455 (O_455,N_13559,N_11573);
xnor UO_456 (O_456,N_10417,N_11724);
nand UO_457 (O_457,N_13925,N_10258);
nand UO_458 (O_458,N_11216,N_11060);
and UO_459 (O_459,N_12965,N_11472);
or UO_460 (O_460,N_12476,N_14492);
or UO_461 (O_461,N_10076,N_10984);
nor UO_462 (O_462,N_13150,N_10156);
nor UO_463 (O_463,N_11703,N_12058);
nor UO_464 (O_464,N_10229,N_14151);
nor UO_465 (O_465,N_11730,N_11720);
and UO_466 (O_466,N_10858,N_11198);
nand UO_467 (O_467,N_13953,N_10189);
nor UO_468 (O_468,N_11375,N_14146);
or UO_469 (O_469,N_10455,N_13035);
nor UO_470 (O_470,N_10837,N_13017);
nor UO_471 (O_471,N_10476,N_10252);
or UO_472 (O_472,N_14450,N_12371);
nor UO_473 (O_473,N_10049,N_14434);
xor UO_474 (O_474,N_13238,N_11542);
or UO_475 (O_475,N_12748,N_14870);
or UO_476 (O_476,N_12430,N_14832);
xnor UO_477 (O_477,N_12916,N_12176);
xor UO_478 (O_478,N_14999,N_11244);
nand UO_479 (O_479,N_13539,N_11792);
and UO_480 (O_480,N_13920,N_10769);
and UO_481 (O_481,N_12307,N_11744);
or UO_482 (O_482,N_10165,N_13166);
and UO_483 (O_483,N_12127,N_13245);
and UO_484 (O_484,N_10318,N_12083);
or UO_485 (O_485,N_13699,N_13876);
or UO_486 (O_486,N_13109,N_14504);
and UO_487 (O_487,N_13531,N_13789);
or UO_488 (O_488,N_12581,N_12885);
nand UO_489 (O_489,N_10009,N_10230);
nand UO_490 (O_490,N_11822,N_10113);
xnor UO_491 (O_491,N_14282,N_10867);
xnor UO_492 (O_492,N_14956,N_12786);
and UO_493 (O_493,N_10932,N_12611);
and UO_494 (O_494,N_12421,N_13337);
or UO_495 (O_495,N_11607,N_10420);
and UO_496 (O_496,N_11231,N_11558);
and UO_497 (O_497,N_10079,N_12336);
or UO_498 (O_498,N_14375,N_12681);
or UO_499 (O_499,N_10040,N_10019);
or UO_500 (O_500,N_11861,N_13459);
xnor UO_501 (O_501,N_12676,N_14599);
nor UO_502 (O_502,N_10716,N_13005);
nor UO_503 (O_503,N_12746,N_10209);
and UO_504 (O_504,N_10375,N_13620);
or UO_505 (O_505,N_13536,N_13519);
xnor UO_506 (O_506,N_13956,N_10314);
and UO_507 (O_507,N_14397,N_14300);
or UO_508 (O_508,N_10625,N_12252);
and UO_509 (O_509,N_11596,N_13407);
xnor UO_510 (O_510,N_11247,N_10149);
xnor UO_511 (O_511,N_11537,N_12757);
nor UO_512 (O_512,N_11002,N_14772);
nor UO_513 (O_513,N_14990,N_11421);
nand UO_514 (O_514,N_13881,N_10288);
or UO_515 (O_515,N_10717,N_13661);
or UO_516 (O_516,N_12949,N_10557);
xor UO_517 (O_517,N_12139,N_10077);
and UO_518 (O_518,N_10221,N_14249);
or UO_519 (O_519,N_10666,N_14577);
or UO_520 (O_520,N_11460,N_12632);
nor UO_521 (O_521,N_14227,N_12027);
xor UO_522 (O_522,N_12523,N_11692);
and UO_523 (O_523,N_10599,N_12097);
or UO_524 (O_524,N_10857,N_13897);
and UO_525 (O_525,N_13019,N_12753);
xor UO_526 (O_526,N_14709,N_12887);
or UO_527 (O_527,N_12472,N_11938);
nand UO_528 (O_528,N_11642,N_10619);
and UO_529 (O_529,N_10907,N_11217);
nand UO_530 (O_530,N_11506,N_14489);
nor UO_531 (O_531,N_14042,N_14381);
nand UO_532 (O_532,N_13844,N_11098);
xor UO_533 (O_533,N_13063,N_13098);
nor UO_534 (O_534,N_11770,N_11479);
nor UO_535 (O_535,N_10612,N_11823);
nand UO_536 (O_536,N_14522,N_12794);
xor UO_537 (O_537,N_14011,N_11318);
and UO_538 (O_538,N_11907,N_13334);
nor UO_539 (O_539,N_10200,N_11122);
nand UO_540 (O_540,N_10686,N_12466);
xnor UO_541 (O_541,N_12579,N_12905);
and UO_542 (O_542,N_13960,N_11233);
nor UO_543 (O_543,N_11541,N_13781);
xor UO_544 (O_544,N_11600,N_14813);
nand UO_545 (O_545,N_12194,N_11668);
nand UO_546 (O_546,N_13513,N_10902);
or UO_547 (O_547,N_12175,N_11304);
or UO_548 (O_548,N_14686,N_13258);
nand UO_549 (O_549,N_14124,N_12913);
or UO_550 (O_550,N_11021,N_14851);
and UO_551 (O_551,N_14131,N_13976);
and UO_552 (O_552,N_12186,N_11234);
nor UO_553 (O_553,N_12266,N_10586);
nor UO_554 (O_554,N_12518,N_14887);
xnor UO_555 (O_555,N_11981,N_10860);
or UO_556 (O_556,N_10691,N_13180);
and UO_557 (O_557,N_11035,N_14836);
and UO_558 (O_558,N_13745,N_13232);
xor UO_559 (O_559,N_10186,N_10870);
nor UO_560 (O_560,N_13804,N_13625);
and UO_561 (O_561,N_12607,N_11650);
and UO_562 (O_562,N_12767,N_12505);
xnor UO_563 (O_563,N_14404,N_12689);
or UO_564 (O_564,N_11982,N_10226);
xnor UO_565 (O_565,N_12730,N_10877);
xor UO_566 (O_566,N_11034,N_10590);
and UO_567 (O_567,N_11387,N_13549);
nand UO_568 (O_568,N_12299,N_14824);
nand UO_569 (O_569,N_11486,N_13938);
xor UO_570 (O_570,N_14060,N_13711);
and UO_571 (O_571,N_11896,N_12813);
and UO_572 (O_572,N_13465,N_14197);
xnor UO_573 (O_573,N_11587,N_12215);
xor UO_574 (O_574,N_11835,N_11432);
nor UO_575 (O_575,N_12773,N_10277);
xnor UO_576 (O_576,N_14499,N_13347);
or UO_577 (O_577,N_12431,N_10397);
nand UO_578 (O_578,N_11985,N_10975);
nand UO_579 (O_579,N_13949,N_14473);
nor UO_580 (O_580,N_10198,N_11523);
and UO_581 (O_581,N_11052,N_13417);
xor UO_582 (O_582,N_14700,N_10052);
nor UO_583 (O_583,N_12105,N_11003);
or UO_584 (O_584,N_13311,N_13105);
xor UO_585 (O_585,N_13324,N_12222);
and UO_586 (O_586,N_10833,N_10474);
and UO_587 (O_587,N_13038,N_12500);
and UO_588 (O_588,N_10523,N_11769);
nor UO_589 (O_589,N_14458,N_14801);
nand UO_590 (O_590,N_11028,N_10366);
nor UO_591 (O_591,N_10206,N_13289);
and UO_592 (O_592,N_13251,N_10735);
nand UO_593 (O_593,N_10896,N_11722);
nand UO_594 (O_594,N_12487,N_10872);
nand UO_595 (O_595,N_11280,N_14127);
xnor UO_596 (O_596,N_13671,N_13762);
and UO_597 (O_597,N_10989,N_10371);
nand UO_598 (O_598,N_14273,N_12549);
nand UO_599 (O_599,N_12877,N_13231);
nand UO_600 (O_600,N_10484,N_12862);
or UO_601 (O_601,N_12953,N_12926);
nor UO_602 (O_602,N_14062,N_12792);
xor UO_603 (O_603,N_12204,N_11434);
nand UO_604 (O_604,N_11030,N_10185);
nand UO_605 (O_605,N_13886,N_12583);
or UO_606 (O_606,N_14563,N_11271);
and UO_607 (O_607,N_13600,N_12151);
nand UO_608 (O_608,N_12292,N_12737);
nand UO_609 (O_609,N_12214,N_11677);
or UO_610 (O_610,N_14490,N_13447);
or UO_611 (O_611,N_10719,N_11102);
and UO_612 (O_612,N_12076,N_10278);
and UO_613 (O_613,N_14507,N_11399);
and UO_614 (O_614,N_12677,N_13444);
and UO_615 (O_615,N_11415,N_12394);
and UO_616 (O_616,N_13968,N_14078);
and UO_617 (O_617,N_10376,N_10879);
nor UO_618 (O_618,N_10309,N_10665);
nand UO_619 (O_619,N_14012,N_14348);
xor UO_620 (O_620,N_10668,N_13036);
or UO_621 (O_621,N_10152,N_13247);
nand UO_622 (O_622,N_10166,N_10470);
nand UO_623 (O_623,N_14322,N_12747);
xnor UO_624 (O_624,N_12826,N_14371);
nand UO_625 (O_625,N_13462,N_13367);
xnor UO_626 (O_626,N_10805,N_14321);
and UO_627 (O_627,N_11313,N_14994);
and UO_628 (O_628,N_11855,N_14867);
nor UO_629 (O_629,N_11858,N_11040);
or UO_630 (O_630,N_13776,N_14349);
nand UO_631 (O_631,N_11236,N_11004);
or UO_632 (O_632,N_11772,N_12341);
xnor UO_633 (O_633,N_14630,N_14770);
or UO_634 (O_634,N_10246,N_12205);
nand UO_635 (O_635,N_12124,N_12280);
nor UO_636 (O_636,N_13416,N_13379);
xor UO_637 (O_637,N_10803,N_12638);
nor UO_638 (O_638,N_11401,N_13831);
and UO_639 (O_639,N_10630,N_13314);
nand UO_640 (O_640,N_14984,N_10132);
nand UO_641 (O_641,N_13865,N_11065);
nand UO_642 (O_642,N_10924,N_14736);
nand UO_643 (O_643,N_13263,N_11001);
nand UO_644 (O_644,N_11616,N_11144);
nor UO_645 (O_645,N_12114,N_12665);
nand UO_646 (O_646,N_14957,N_12405);
nor UO_647 (O_647,N_10083,N_10167);
nand UO_648 (O_648,N_12739,N_10920);
xor UO_649 (O_649,N_13614,N_13544);
nand UO_650 (O_650,N_14483,N_14117);
nand UO_651 (O_651,N_14001,N_11273);
and UO_652 (O_652,N_14377,N_13927);
nor UO_653 (O_653,N_12013,N_12185);
nand UO_654 (O_654,N_12230,N_10751);
nand UO_655 (O_655,N_10003,N_12592);
nand UO_656 (O_656,N_11171,N_13857);
xnor UO_657 (O_657,N_14834,N_12041);
or UO_658 (O_658,N_14099,N_14463);
nand UO_659 (O_659,N_13780,N_14518);
xor UO_660 (O_660,N_14390,N_13666);
nand UO_661 (O_661,N_13608,N_13266);
nor UO_662 (O_662,N_12228,N_11005);
or UO_663 (O_663,N_14714,N_10820);
xor UO_664 (O_664,N_13214,N_14260);
and UO_665 (O_665,N_14346,N_13819);
xnor UO_666 (O_666,N_13013,N_13828);
nand UO_667 (O_667,N_11316,N_13705);
or UO_668 (O_668,N_13366,N_12836);
and UO_669 (O_669,N_14268,N_14694);
nor UO_670 (O_670,N_12361,N_13644);
and UO_671 (O_671,N_10099,N_11490);
xnor UO_672 (O_672,N_12311,N_13733);
and UO_673 (O_673,N_14204,N_11839);
nand UO_674 (O_674,N_12192,N_10755);
or UO_675 (O_675,N_11281,N_13074);
and UO_676 (O_676,N_10821,N_13827);
or UO_677 (O_677,N_14558,N_10102);
and UO_678 (O_678,N_12948,N_11746);
nor UO_679 (O_679,N_14860,N_11540);
and UO_680 (O_680,N_14406,N_12251);
nor UO_681 (O_681,N_11013,N_12386);
or UO_682 (O_682,N_13476,N_12149);
nor UO_683 (O_683,N_13428,N_10789);
or UO_684 (O_684,N_14923,N_13103);
nor UO_685 (O_685,N_11790,N_13001);
xnor UO_686 (O_686,N_14288,N_13615);
or UO_687 (O_687,N_14120,N_12155);
or UO_688 (O_688,N_13413,N_14175);
and UO_689 (O_689,N_11107,N_11825);
nand UO_690 (O_690,N_11879,N_14945);
and UO_691 (O_691,N_11183,N_12731);
xnor UO_692 (O_692,N_12126,N_12473);
xor UO_693 (O_693,N_11339,N_13669);
or UO_694 (O_694,N_12179,N_10996);
or UO_695 (O_695,N_11632,N_12847);
xor UO_696 (O_696,N_14650,N_14894);
nand UO_697 (O_697,N_13280,N_13524);
nor UO_698 (O_698,N_12284,N_10158);
nor UO_699 (O_699,N_10175,N_12557);
xnor UO_700 (O_700,N_10522,N_14874);
and UO_701 (O_701,N_14461,N_12342);
nand UO_702 (O_702,N_10938,N_14468);
nand UO_703 (O_703,N_12220,N_14640);
or UO_704 (O_704,N_14792,N_10635);
and UO_705 (O_705,N_14033,N_13777);
nand UO_706 (O_706,N_10305,N_11197);
nor UO_707 (O_707,N_11344,N_10135);
xor UO_708 (O_708,N_12680,N_11911);
and UO_709 (O_709,N_10991,N_12106);
and UO_710 (O_710,N_11843,N_14075);
or UO_711 (O_711,N_10108,N_11302);
and UO_712 (O_712,N_10404,N_11448);
and UO_713 (O_713,N_14838,N_10337);
xor UO_714 (O_714,N_14654,N_11990);
and UO_715 (O_715,N_10449,N_13077);
or UO_716 (O_716,N_10245,N_10689);
nor UO_717 (O_717,N_11742,N_14871);
and UO_718 (O_718,N_13728,N_11503);
xnor UO_719 (O_719,N_11497,N_12652);
xor UO_720 (O_720,N_12174,N_10228);
and UO_721 (O_721,N_11821,N_10297);
nand UO_722 (O_722,N_14803,N_14835);
nand UO_723 (O_723,N_13832,N_13389);
nor UO_724 (O_724,N_14959,N_11215);
nor UO_725 (O_725,N_13064,N_14054);
nand UO_726 (O_726,N_13443,N_10529);
nor UO_727 (O_727,N_14362,N_14126);
or UO_728 (O_728,N_12484,N_14728);
nand UO_729 (O_729,N_12619,N_14865);
and UO_730 (O_730,N_10777,N_11872);
or UO_731 (O_731,N_13022,N_14436);
nand UO_732 (O_732,N_12474,N_10154);
nor UO_733 (O_733,N_13176,N_10127);
xor UO_734 (O_734,N_11671,N_12563);
xor UO_735 (O_735,N_14080,N_12804);
nor UO_736 (O_736,N_13845,N_14220);
nor UO_737 (O_737,N_14392,N_10022);
xnor UO_738 (O_738,N_12520,N_11022);
or UO_739 (O_739,N_10880,N_11284);
nand UO_740 (O_740,N_13651,N_11832);
or UO_741 (O_741,N_13978,N_13975);
nor UO_742 (O_742,N_13170,N_10883);
and UO_743 (O_743,N_10539,N_11653);
nand UO_744 (O_744,N_14612,N_12010);
xor UO_745 (O_745,N_14818,N_13302);
and UO_746 (O_746,N_12533,N_12839);
xnor UO_747 (O_747,N_11551,N_11410);
nor UO_748 (O_748,N_14241,N_14723);
xor UO_749 (O_749,N_14462,N_10897);
xnor UO_750 (O_750,N_13235,N_12754);
nor UO_751 (O_751,N_11041,N_12831);
xor UO_752 (O_752,N_12271,N_11796);
xor UO_753 (O_753,N_13202,N_14868);
nand UO_754 (O_754,N_13033,N_12070);
xor UO_755 (O_755,N_11922,N_13670);
or UO_756 (O_756,N_10499,N_14039);
and UO_757 (O_757,N_12674,N_14480);
or UO_758 (O_758,N_12296,N_13743);
nand UO_759 (O_759,N_13583,N_13610);
nand UO_760 (O_760,N_12655,N_11296);
or UO_761 (O_761,N_12440,N_11687);
nor UO_762 (O_762,N_10886,N_14796);
and UO_763 (O_763,N_11024,N_10634);
or UO_764 (O_764,N_14596,N_11952);
or UO_765 (O_765,N_11705,N_11213);
xnor UO_766 (O_766,N_10863,N_12035);
nand UO_767 (O_767,N_13003,N_11775);
nor UO_768 (O_768,N_11335,N_10025);
nor UO_769 (O_769,N_10799,N_11148);
or UO_770 (O_770,N_11753,N_10993);
or UO_771 (O_771,N_10667,N_10848);
nand UO_772 (O_772,N_10172,N_12559);
xnor UO_773 (O_773,N_12483,N_11493);
xor UO_774 (O_774,N_10573,N_11136);
nor UO_775 (O_775,N_13732,N_13149);
and UO_776 (O_776,N_11371,N_14624);
nor UO_777 (O_777,N_12090,N_11610);
xor UO_778 (O_778,N_13717,N_13659);
nor UO_779 (O_779,N_10603,N_11188);
nand UO_780 (O_780,N_10133,N_12080);
or UO_781 (O_781,N_11886,N_13606);
nor UO_782 (O_782,N_10535,N_13253);
nand UO_783 (O_783,N_14304,N_11225);
or UO_784 (O_784,N_11875,N_11298);
xor UO_785 (O_785,N_10176,N_13461);
nand UO_786 (O_786,N_12193,N_12123);
xnor UO_787 (O_787,N_11116,N_12552);
xnor UO_788 (O_788,N_10358,N_11580);
and UO_789 (O_789,N_13269,N_11856);
or UO_790 (O_790,N_13141,N_10749);
xnor UO_791 (O_791,N_14717,N_13858);
nor UO_792 (O_792,N_10800,N_12818);
nor UO_793 (O_793,N_12378,N_12895);
nand UO_794 (O_794,N_10396,N_14313);
and UO_795 (O_795,N_10760,N_11900);
and UO_796 (O_796,N_11870,N_13351);
xor UO_797 (O_797,N_12153,N_12216);
xor UO_798 (O_798,N_13621,N_14546);
and UO_799 (O_799,N_11032,N_14787);
nor UO_800 (O_800,N_12054,N_11901);
and UO_801 (O_801,N_10150,N_10480);
nor UO_802 (O_802,N_10759,N_13326);
nand UO_803 (O_803,N_11409,N_13639);
and UO_804 (O_804,N_10854,N_14366);
and UO_805 (O_805,N_12646,N_14048);
xnor UO_806 (O_806,N_10092,N_13268);
xor UO_807 (O_807,N_12295,N_11570);
and UO_808 (O_808,N_14886,N_14159);
and UO_809 (O_809,N_13866,N_14259);
nor UO_810 (O_810,N_11471,N_10467);
nor UO_811 (O_811,N_11695,N_11286);
nand UO_812 (O_812,N_11036,N_10412);
xor UO_813 (O_813,N_12845,N_12349);
and UO_814 (O_814,N_12915,N_12052);
xor UO_815 (O_815,N_12111,N_14019);
and UO_816 (O_816,N_13441,N_14707);
and UO_817 (O_817,N_13052,N_11046);
and UO_818 (O_818,N_10983,N_14104);
nor UO_819 (O_819,N_12899,N_12053);
nor UO_820 (O_820,N_11709,N_10957);
and UO_821 (O_821,N_10921,N_14066);
or UO_822 (O_822,N_10588,N_10594);
xor UO_823 (O_823,N_14602,N_11947);
and UO_824 (O_824,N_14595,N_12586);
and UO_825 (O_825,N_13454,N_10339);
and UO_826 (O_826,N_14564,N_14879);
nor UO_827 (O_827,N_12783,N_12059);
or UO_828 (O_828,N_14256,N_11241);
xnor UO_829 (O_829,N_14782,N_14962);
nor UO_830 (O_830,N_10115,N_12999);
xor UO_831 (O_831,N_13618,N_10828);
and UO_832 (O_832,N_14676,N_10782);
and UO_833 (O_833,N_13164,N_11934);
or UO_834 (O_834,N_14614,N_14555);
or UO_835 (O_835,N_11998,N_12760);
or UO_836 (O_836,N_14308,N_10117);
nand UO_837 (O_837,N_14977,N_13393);
or UO_838 (O_838,N_14167,N_12687);
nand UO_839 (O_839,N_11893,N_12449);
xor UO_840 (O_840,N_13761,N_10121);
xnor UO_841 (O_841,N_14449,N_14847);
or UO_842 (O_842,N_12834,N_11533);
nor UO_843 (O_843,N_13174,N_10548);
nand UO_844 (O_844,N_10275,N_12429);
and UO_845 (O_845,N_12896,N_11353);
or UO_846 (O_846,N_10644,N_14697);
and UO_847 (O_847,N_13940,N_10126);
or UO_848 (O_848,N_11088,N_12438);
nor UO_849 (O_849,N_14153,N_14323);
nor UO_850 (O_850,N_11266,N_10129);
and UO_851 (O_851,N_13330,N_13048);
nand UO_852 (O_852,N_11084,N_10801);
nand UO_853 (O_853,N_13420,N_14698);
nor UO_854 (O_854,N_10720,N_11602);
nor UO_855 (O_855,N_12672,N_10551);
and UO_856 (O_856,N_11164,N_10949);
or UO_857 (O_857,N_11285,N_11548);
and UO_858 (O_858,N_11114,N_13972);
xnor UO_859 (O_859,N_11794,N_10213);
or UO_860 (O_860,N_13664,N_13093);
nor UO_861 (O_861,N_12081,N_14111);
and UO_862 (O_862,N_10695,N_11287);
nor UO_863 (O_863,N_10609,N_11656);
or UO_864 (O_864,N_10961,N_14679);
xor UO_865 (O_865,N_11785,N_10868);
and UO_866 (O_866,N_14098,N_14855);
nand UO_867 (O_867,N_12558,N_13088);
nor UO_868 (O_868,N_13237,N_12762);
nand UO_869 (O_869,N_12541,N_13274);
and UO_870 (O_870,N_10659,N_10144);
nor UO_871 (O_871,N_11691,N_11801);
nand UO_872 (O_872,N_10500,N_14550);
xor UO_873 (O_873,N_13812,N_10197);
nand UO_874 (O_874,N_10680,N_10242);
xnor UO_875 (O_875,N_13148,N_13983);
xor UO_876 (O_876,N_12020,N_13895);
and UO_877 (O_877,N_13642,N_10210);
and UO_878 (O_878,N_11307,N_14895);
nand UO_879 (O_879,N_11550,N_14298);
and UO_880 (O_880,N_12247,N_12261);
xnor UO_881 (O_881,N_13992,N_11535);
nand UO_882 (O_882,N_13721,N_12945);
and UO_883 (O_883,N_11424,N_13851);
nand UO_884 (O_884,N_14783,N_14573);
xnor UO_885 (O_885,N_10795,N_13805);
nand UO_886 (O_886,N_13125,N_12981);
nand UO_887 (O_887,N_12037,N_14583);
xnor UO_888 (O_888,N_13292,N_13787);
nand UO_889 (O_889,N_12864,N_12992);
xor UO_890 (O_890,N_13415,N_13913);
or UO_891 (O_891,N_13856,N_11578);
xnor UO_892 (O_892,N_12246,N_11818);
nand UO_893 (O_893,N_14232,N_13735);
or UO_894 (O_894,N_10936,N_11159);
xnor UO_895 (O_895,N_12122,N_12645);
and UO_896 (O_896,N_14234,N_13290);
or UO_897 (O_897,N_11688,N_10071);
nor UO_898 (O_898,N_11965,N_11124);
nand UO_899 (O_899,N_13279,N_13229);
nand UO_900 (O_900,N_13929,N_14567);
nor UO_901 (O_901,N_13788,N_14110);
or UO_902 (O_902,N_13716,N_12188);
and UO_903 (O_903,N_12838,N_10652);
and UO_904 (O_904,N_10341,N_13031);
xnor UO_905 (O_905,N_13966,N_13426);
and UO_906 (O_906,N_11006,N_13686);
xor UO_907 (O_907,N_14695,N_14866);
xnor UO_908 (O_908,N_11690,N_14944);
or UO_909 (O_909,N_11552,N_11105);
and UO_910 (O_910,N_10823,N_11325);
and UO_911 (O_911,N_11121,N_12769);
xor UO_912 (O_912,N_10598,N_12751);
nand UO_913 (O_913,N_11111,N_13049);
xnor UO_914 (O_914,N_10050,N_14715);
nand UO_915 (O_915,N_10550,N_11150);
nand UO_916 (O_916,N_13909,N_12259);
or UO_917 (O_917,N_13025,N_13058);
xor UO_918 (O_918,N_14857,N_13187);
and UO_919 (O_919,N_10604,N_11662);
xnor UO_920 (O_920,N_13185,N_14306);
or UO_921 (O_921,N_11637,N_14297);
xnor UO_922 (O_922,N_12324,N_14257);
nand UO_923 (O_923,N_10479,N_12439);
and UO_924 (O_924,N_12625,N_10414);
xnor UO_925 (O_925,N_13475,N_12613);
nor UO_926 (O_926,N_14281,N_11468);
or UO_927 (O_927,N_12136,N_12668);
xnor UO_928 (O_928,N_12596,N_14193);
nor UO_929 (O_929,N_14229,N_14457);
xor UO_930 (O_930,N_10440,N_10345);
nor UO_931 (O_931,N_10095,N_12278);
or UO_932 (O_932,N_10894,N_10818);
xnor UO_933 (O_933,N_12593,N_12589);
nor UO_934 (O_934,N_14935,N_13551);
xnor UO_935 (O_935,N_12065,N_14200);
nand UO_936 (O_936,N_11956,N_11018);
nand UO_937 (O_937,N_10369,N_11366);
nand UO_938 (O_938,N_12343,N_14223);
xnor UO_939 (O_939,N_11229,N_11891);
nor UO_940 (O_940,N_13982,N_14382);
and UO_941 (O_941,N_10041,N_11283);
nand UO_942 (O_942,N_11964,N_11831);
or UO_943 (O_943,N_10926,N_10636);
or UO_944 (O_944,N_12331,N_13597);
nor UO_945 (O_945,N_10976,N_10224);
xnor UO_946 (O_946,N_13356,N_14134);
or UO_947 (O_947,N_10521,N_14675);
or UO_948 (O_948,N_13967,N_11502);
xor UO_949 (O_949,N_12023,N_12046);
and UO_950 (O_950,N_12758,N_13097);
xor UO_951 (O_951,N_10247,N_13386);
nand UO_952 (O_952,N_13489,N_10217);
and UO_953 (O_953,N_14456,N_10360);
and UO_954 (O_954,N_12971,N_10761);
xor UO_955 (O_955,N_11452,N_12716);
xor UO_956 (O_956,N_13236,N_10884);
and UO_957 (O_957,N_12465,N_10319);
and UO_958 (O_958,N_12288,N_12458);
nor UO_959 (O_959,N_12075,N_10718);
and UO_960 (O_960,N_11356,N_10583);
xor UO_961 (O_961,N_13527,N_13941);
or UO_962 (O_962,N_12067,N_14508);
xnor UO_963 (O_963,N_13782,N_12374);
nand UO_964 (O_964,N_11626,N_12277);
nor UO_965 (O_965,N_14571,N_10111);
and UO_966 (O_966,N_10622,N_10553);
or UO_967 (O_967,N_11845,N_10142);
or UO_968 (O_968,N_10477,N_14387);
or UO_969 (O_969,N_10554,N_13868);
or UO_970 (O_970,N_13663,N_12705);
xnor UO_971 (O_971,N_13323,N_11403);
nand UO_972 (O_972,N_10660,N_14057);
xor UO_973 (O_973,N_13155,N_11227);
and UO_974 (O_974,N_11866,N_13159);
xnor UO_975 (O_975,N_14704,N_14174);
nand UO_976 (O_976,N_13278,N_13358);
nor UO_977 (O_977,N_13673,N_14135);
or UO_978 (O_978,N_11301,N_12197);
nor UO_979 (O_979,N_13638,N_14484);
xnor UO_980 (O_980,N_11991,N_13510);
nor UO_981 (O_981,N_11887,N_11303);
nor UO_982 (O_982,N_10125,N_14173);
xor UO_983 (O_983,N_11697,N_11405);
xor UO_984 (O_984,N_10323,N_13601);
nand UO_985 (O_985,N_11723,N_10490);
and UO_986 (O_986,N_11143,N_11614);
nand UO_987 (O_987,N_12734,N_13529);
nand UO_988 (O_988,N_12946,N_13365);
nor UO_989 (O_989,N_14703,N_13973);
nor UO_990 (O_990,N_14277,N_10109);
or UO_991 (O_991,N_13104,N_12679);
and UO_992 (O_992,N_11849,N_12942);
or UO_993 (O_993,N_10249,N_10766);
nand UO_994 (O_994,N_10772,N_12853);
and UO_995 (O_995,N_13070,N_10946);
xor UO_996 (O_996,N_12166,N_10608);
xor UO_997 (O_997,N_11549,N_11585);
nand UO_998 (O_998,N_14589,N_14613);
nand UO_999 (O_999,N_10134,N_13002);
or UO_1000 (O_1000,N_14476,N_12250);
nand UO_1001 (O_1001,N_13888,N_13649);
nand UO_1002 (O_1002,N_10696,N_11867);
xor UO_1003 (O_1003,N_14789,N_14862);
xnor UO_1004 (O_1004,N_13136,N_12584);
xor UO_1005 (O_1005,N_12300,N_13813);
xor UO_1006 (O_1006,N_13199,N_12173);
nand UO_1007 (O_1007,N_12778,N_11063);
nand UO_1008 (O_1008,N_10591,N_14255);
nor UO_1009 (O_1009,N_10451,N_10373);
nand UO_1010 (O_1010,N_11480,N_12793);
or UO_1011 (O_1011,N_14271,N_11081);
xor UO_1012 (O_1012,N_10407,N_12079);
nor UO_1013 (O_1013,N_12692,N_10538);
nand UO_1014 (O_1014,N_10744,N_13826);
xnor UO_1015 (O_1015,N_12267,N_14157);
nor UO_1016 (O_1016,N_14967,N_11519);
nor UO_1017 (O_1017,N_11530,N_14205);
or UO_1018 (O_1018,N_13565,N_14934);
nand UO_1019 (O_1019,N_13308,N_10359);
nor UO_1020 (O_1020,N_13902,N_11917);
or UO_1021 (O_1021,N_10048,N_14413);
or UO_1022 (O_1022,N_12477,N_13718);
or UO_1023 (O_1023,N_10141,N_14024);
nor UO_1024 (O_1024,N_11038,N_14162);
or UO_1025 (O_1025,N_12983,N_13084);
nand UO_1026 (O_1026,N_11255,N_14983);
nand UO_1027 (O_1027,N_12506,N_14319);
and UO_1028 (O_1028,N_11783,N_10332);
xor UO_1029 (O_1029,N_10329,N_13053);
nor UO_1030 (O_1030,N_14186,N_14324);
or UO_1031 (O_1031,N_10300,N_11756);
and UO_1032 (O_1032,N_13662,N_14044);
nand UO_1033 (O_1033,N_13167,N_10581);
nand UO_1034 (O_1034,N_13320,N_14150);
and UO_1035 (O_1035,N_14765,N_10317);
xnor UO_1036 (O_1036,N_14758,N_11797);
or UO_1037 (O_1037,N_13939,N_11700);
xor UO_1038 (O_1038,N_10900,N_11087);
nand UO_1039 (O_1039,N_12977,N_13341);
xnor UO_1040 (O_1040,N_14726,N_13993);
nor UO_1041 (O_1041,N_13795,N_10391);
and UO_1042 (O_1042,N_12212,N_12883);
nand UO_1043 (O_1043,N_10062,N_11735);
xnor UO_1044 (O_1044,N_11178,N_13921);
xor UO_1045 (O_1045,N_14606,N_10204);
or UO_1046 (O_1046,N_14702,N_12938);
xor UO_1047 (O_1047,N_12370,N_11334);
or UO_1048 (O_1048,N_11349,N_11259);
xor UO_1049 (O_1049,N_13930,N_12260);
nor UO_1050 (O_1050,N_10075,N_13062);
xnor UO_1051 (O_1051,N_11263,N_10408);
and UO_1052 (O_1052,N_12353,N_11788);
xor UO_1053 (O_1053,N_12084,N_14275);
nor UO_1054 (O_1054,N_14532,N_11803);
nand UO_1055 (O_1055,N_13075,N_13453);
nor UO_1056 (O_1056,N_10582,N_13604);
or UO_1057 (O_1057,N_11814,N_14721);
xnor UO_1058 (O_1058,N_11683,N_11348);
or UO_1059 (O_1059,N_12334,N_14311);
or UO_1060 (O_1060,N_13679,N_10816);
or UO_1061 (O_1061,N_14905,N_11130);
nand UO_1062 (O_1062,N_11902,N_11211);
or UO_1063 (O_1063,N_14689,N_13220);
nor UO_1064 (O_1064,N_14692,N_12002);
nor UO_1065 (O_1065,N_13307,N_10436);
or UO_1066 (O_1066,N_10104,N_10569);
xor UO_1067 (O_1067,N_14846,N_12162);
or UO_1068 (O_1068,N_12442,N_14339);
or UO_1069 (O_1069,N_11890,N_13255);
or UO_1070 (O_1070,N_13037,N_11941);
xnor UO_1071 (O_1071,N_14969,N_12779);
or UO_1072 (O_1072,N_11527,N_10465);
nor UO_1073 (O_1073,N_14748,N_13985);
nor UO_1074 (O_1074,N_11729,N_11414);
nor UO_1075 (O_1075,N_12424,N_10901);
nor UO_1076 (O_1076,N_14928,N_14393);
nor UO_1077 (O_1077,N_12513,N_11805);
nand UO_1078 (O_1078,N_10304,N_10259);
nand UO_1079 (O_1079,N_10978,N_12647);
or UO_1080 (O_1080,N_12086,N_12328);
or UO_1081 (O_1081,N_12708,N_11361);
and UO_1082 (O_1082,N_11015,N_10293);
or UO_1083 (O_1083,N_11218,N_14417);
xnor UO_1084 (O_1084,N_12116,N_14085);
nor UO_1085 (O_1085,N_10215,N_10118);
xnor UO_1086 (O_1086,N_13961,N_11196);
or UO_1087 (O_1087,N_12670,N_10977);
nand UO_1088 (O_1088,N_14989,N_12367);
or UO_1089 (O_1089,N_10684,N_11478);
or UO_1090 (O_1090,N_14500,N_13092);
nand UO_1091 (O_1091,N_10753,N_10905);
and UO_1092 (O_1092,N_10694,N_13917);
nand UO_1093 (O_1093,N_13763,N_13260);
nor UO_1094 (O_1094,N_14942,N_13449);
nor UO_1095 (O_1095,N_12049,N_11629);
or UO_1096 (O_1096,N_13222,N_14059);
nand UO_1097 (O_1097,N_14005,N_13343);
xnor UO_1098 (O_1098,N_14858,N_14793);
nor UO_1099 (O_1099,N_10024,N_12874);
nand UO_1100 (O_1100,N_14883,N_10633);
and UO_1101 (O_1101,N_10838,N_13156);
nand UO_1102 (O_1102,N_12380,N_11568);
or UO_1103 (O_1103,N_11708,N_11702);
or UO_1104 (O_1104,N_14786,N_11949);
and UO_1105 (O_1105,N_11824,N_10462);
nand UO_1106 (O_1106,N_12399,N_11489);
or UO_1107 (O_1107,N_14511,N_11924);
or UO_1108 (O_1108,N_10917,N_11407);
nand UO_1109 (O_1109,N_10968,N_13288);
and UO_1110 (O_1110,N_11895,N_14230);
nand UO_1111 (O_1111,N_11577,N_10875);
nor UO_1112 (O_1112,N_12857,N_13668);
xor UO_1113 (O_1113,N_14305,N_11282);
nand UO_1114 (O_1114,N_13872,N_10552);
or UO_1115 (O_1115,N_10651,N_13338);
or UO_1116 (O_1116,N_11973,N_12488);
nand UO_1117 (O_1117,N_14738,N_11435);
xnor UO_1118 (O_1118,N_10481,N_10112);
nand UO_1119 (O_1119,N_11834,N_13792);
nand UO_1120 (O_1120,N_11312,N_11447);
and UO_1121 (O_1121,N_11064,N_10681);
xor UO_1122 (O_1122,N_11673,N_14802);
or UO_1123 (O_1123,N_14991,N_14106);
and UO_1124 (O_1124,N_14113,N_10308);
xnor UO_1125 (O_1125,N_12653,N_12688);
nand UO_1126 (O_1126,N_10409,N_13273);
nand UO_1127 (O_1127,N_14719,N_12765);
xnor UO_1128 (O_1128,N_11859,N_13759);
or UO_1129 (O_1129,N_13342,N_10265);
nor UO_1130 (O_1130,N_10143,N_13169);
nand UO_1131 (O_1131,N_11093,N_12522);
or UO_1132 (O_1132,N_14307,N_13727);
xnor UO_1133 (O_1133,N_14646,N_11091);
nor UO_1134 (O_1134,N_14233,N_12889);
xor UO_1135 (O_1135,N_14201,N_13215);
xor UO_1136 (O_1136,N_14509,N_14877);
nand UO_1137 (O_1137,N_13952,N_14993);
nand UO_1138 (O_1138,N_10177,N_11049);
or UO_1139 (O_1139,N_12876,N_11482);
nand UO_1140 (O_1140,N_13352,N_10615);
or UO_1141 (O_1141,N_13822,N_14089);
nor UO_1142 (O_1142,N_11987,N_12202);
and UO_1143 (O_1143,N_14644,N_11747);
nor UO_1144 (O_1144,N_10616,N_13399);
or UO_1145 (O_1145,N_13507,N_11660);
xnor UO_1146 (O_1146,N_10054,N_13026);
nand UO_1147 (O_1147,N_12939,N_13438);
xor UO_1148 (O_1148,N_11631,N_11126);
and UO_1149 (O_1149,N_14909,N_10354);
or UO_1150 (O_1150,N_13480,N_13414);
xnor UO_1151 (O_1151,N_12580,N_12616);
and UO_1152 (O_1152,N_14046,N_13305);
nand UO_1153 (O_1153,N_13467,N_13401);
and UO_1154 (O_1154,N_10364,N_12937);
nor UO_1155 (O_1155,N_13121,N_13965);
and UO_1156 (O_1156,N_12812,N_14338);
and UO_1157 (O_1157,N_12337,N_13977);
xor UO_1158 (O_1158,N_14238,N_13988);
xnor UO_1159 (O_1159,N_11451,N_14673);
nor UO_1160 (O_1160,N_10138,N_13439);
xnor UO_1161 (O_1161,N_10904,N_12814);
or UO_1162 (O_1162,N_10618,N_14986);
and UO_1163 (O_1163,N_12759,N_10617);
nor UO_1164 (O_1164,N_14049,N_11305);
nor UO_1165 (O_1165,N_13259,N_13692);
nor UO_1166 (O_1166,N_13325,N_13591);
nor UO_1167 (O_1167,N_10424,N_10428);
and UO_1168 (O_1168,N_11505,N_13747);
xnor UO_1169 (O_1169,N_14618,N_14445);
xor UO_1170 (O_1170,N_14408,N_10001);
or UO_1171 (O_1171,N_14002,N_12733);
nor UO_1172 (O_1172,N_14130,N_10646);
or UO_1173 (O_1173,N_14591,N_14732);
nor UO_1174 (O_1174,N_12825,N_12078);
nor UO_1175 (O_1175,N_13891,N_13843);
and UO_1176 (O_1176,N_13755,N_10458);
nor UO_1177 (O_1177,N_12335,N_12359);
nor UO_1178 (O_1178,N_13131,N_10788);
or UO_1179 (O_1179,N_12134,N_14287);
nor UO_1180 (O_1180,N_14081,N_13807);
nand UO_1181 (O_1181,N_12320,N_11476);
xnor UO_1182 (O_1182,N_12966,N_13119);
or UO_1183 (O_1183,N_12096,N_11269);
nor UO_1184 (O_1184,N_12850,N_14160);
nand UO_1185 (O_1185,N_11363,N_13284);
nand UO_1186 (O_1186,N_12117,N_14014);
xor UO_1187 (O_1187,N_12993,N_11189);
or UO_1188 (O_1188,N_13328,N_14973);
and UO_1189 (O_1189,N_11464,N_12470);
nor UO_1190 (O_1190,N_11146,N_11186);
nor UO_1191 (O_1191,N_11745,N_13418);
nand UO_1192 (O_1192,N_10400,N_11766);
and UO_1193 (O_1193,N_14885,N_11881);
and UO_1194 (O_1194,N_14668,N_14222);
xor UO_1195 (O_1195,N_12774,N_10064);
nand UO_1196 (O_1196,N_11395,N_13979);
or UO_1197 (O_1197,N_12894,N_10676);
xor UO_1198 (O_1198,N_12639,N_13423);
nor UO_1199 (O_1199,N_10352,N_11793);
nor UO_1200 (O_1200,N_11295,N_10722);
or UO_1201 (O_1201,N_14901,N_13402);
and UO_1202 (O_1202,N_12314,N_10164);
nor UO_1203 (O_1203,N_11517,N_10281);
nand UO_1204 (O_1204,N_10600,N_12661);
or UO_1205 (O_1205,N_11651,N_13479);
and UO_1206 (O_1206,N_10012,N_11611);
nor UO_1207 (O_1207,N_10273,N_10236);
nor UO_1208 (O_1208,N_10826,N_10289);
and UO_1209 (O_1209,N_13801,N_11943);
and UO_1210 (O_1210,N_13216,N_12524);
and UO_1211 (O_1211,N_12478,N_10122);
and UO_1212 (O_1212,N_14822,N_14741);
nand UO_1213 (O_1213,N_10146,N_10510);
and UO_1214 (O_1214,N_13059,N_12383);
nand UO_1215 (O_1215,N_11445,N_12863);
xnor UO_1216 (O_1216,N_13590,N_12258);
and UO_1217 (O_1217,N_13835,N_13113);
xor UO_1218 (O_1218,N_12365,N_13233);
or UO_1219 (O_1219,N_11971,N_11743);
xnor UO_1220 (O_1220,N_14430,N_14899);
nand UO_1221 (O_1221,N_12048,N_11200);
xnor UO_1222 (O_1222,N_11698,N_11584);
nand UO_1223 (O_1223,N_10395,N_12744);
or UO_1224 (O_1224,N_10454,N_11166);
xnor UO_1225 (O_1225,N_10168,N_14276);
and UO_1226 (O_1226,N_10466,N_11727);
nand UO_1227 (O_1227,N_14231,N_13605);
nand UO_1228 (O_1228,N_11428,N_13205);
nand UO_1229 (O_1229,N_13183,N_12308);
nand UO_1230 (O_1230,N_10531,N_11995);
nor UO_1231 (O_1231,N_14806,N_12108);
nor UO_1232 (O_1232,N_12290,N_11072);
nor UO_1233 (O_1233,N_14627,N_12886);
or UO_1234 (O_1234,N_10063,N_12302);
or UO_1235 (O_1235,N_14171,N_11125);
nand UO_1236 (O_1236,N_10943,N_12008);
nand UO_1237 (O_1237,N_11625,N_10448);
nor UO_1238 (O_1238,N_12218,N_10433);
or UO_1239 (O_1239,N_14141,N_14469);
xor UO_1240 (O_1240,N_11073,N_12032);
or UO_1241 (O_1241,N_14623,N_12113);
or UO_1242 (O_1242,N_12921,N_11903);
or UO_1243 (O_1243,N_11576,N_11265);
xnor UO_1244 (O_1244,N_13240,N_10051);
nor UO_1245 (O_1245,N_13955,N_13014);
nor UO_1246 (O_1246,N_11390,N_12392);
and UO_1247 (O_1247,N_11162,N_11833);
and UO_1248 (O_1248,N_12433,N_13223);
and UO_1249 (O_1249,N_12690,N_11450);
xor UO_1250 (O_1250,N_11598,N_13172);
xnor UO_1251 (O_1251,N_11669,N_11951);
nand UO_1252 (O_1252,N_14015,N_10587);
nor UO_1253 (O_1253,N_13140,N_11597);
or UO_1254 (O_1254,N_13687,N_13458);
or UO_1255 (O_1255,N_11630,N_10029);
xor UO_1256 (O_1256,N_11935,N_14119);
and UO_1257 (O_1257,N_13118,N_13943);
nor UO_1258 (O_1258,N_13817,N_11583);
nand UO_1259 (O_1259,N_14970,N_14776);
xor UO_1260 (O_1260,N_14713,N_12702);
and UO_1261 (O_1261,N_11484,N_13432);
or UO_1262 (O_1262,N_12373,N_12598);
nand UO_1263 (O_1263,N_14906,N_13974);
and UO_1264 (O_1264,N_14519,N_13316);
nand UO_1265 (O_1265,N_13562,N_11474);
and UO_1266 (O_1266,N_11579,N_13046);
nor UO_1267 (O_1267,N_13581,N_13120);
nand UO_1268 (O_1268,N_10947,N_11347);
nand UO_1269 (O_1269,N_11711,N_14472);
and UO_1270 (O_1270,N_13364,N_10426);
nor UO_1271 (O_1271,N_12125,N_10216);
nor UO_1272 (O_1272,N_14826,N_14217);
and UO_1273 (O_1273,N_12684,N_10764);
and UO_1274 (O_1274,N_14481,N_13080);
nand UO_1275 (O_1275,N_13577,N_10878);
xor UO_1276 (O_1276,N_10687,N_13859);
and UO_1277 (O_1277,N_11817,N_11290);
xnor UO_1278 (O_1278,N_14283,N_10128);
xor UO_1279 (O_1279,N_11525,N_13803);
xnor UO_1280 (O_1280,N_11154,N_12601);
nand UO_1281 (O_1281,N_12703,N_11117);
xor UO_1282 (O_1282,N_14678,N_12257);
nor UO_1283 (O_1283,N_11980,N_12254);
and UO_1284 (O_1284,N_13071,N_14746);
nand UO_1285 (O_1285,N_10524,N_11714);
and UO_1286 (O_1286,N_10348,N_14444);
or UO_1287 (O_1287,N_14289,N_12978);
nand UO_1288 (O_1288,N_13877,N_14292);
xnor UO_1289 (O_1289,N_11538,N_14453);
xnor UO_1290 (O_1290,N_11199,N_12662);
nand UO_1291 (O_1291,N_14161,N_13767);
nor UO_1292 (O_1292,N_10392,N_11389);
nand UO_1293 (O_1293,N_12644,N_12238);
nor UO_1294 (O_1294,N_11174,N_14006);
nand UO_1295 (O_1295,N_13713,N_14405);
xnor UO_1296 (O_1296,N_14309,N_14314);
nor UO_1297 (O_1297,N_11172,N_10445);
or UO_1298 (O_1298,N_14998,N_12031);
and UO_1299 (O_1299,N_12493,N_13034);
nor UO_1300 (O_1300,N_13488,N_13528);
nor UO_1301 (O_1301,N_12934,N_10004);
or UO_1302 (O_1302,N_13353,N_13009);
and UO_1303 (O_1303,N_11898,N_10223);
nand UO_1304 (O_1304,N_14486,N_12764);
or UO_1305 (O_1305,N_13648,N_11619);
and UO_1306 (O_1306,N_14389,N_10489);
nor UO_1307 (O_1307,N_10306,N_13135);
nor UO_1308 (O_1308,N_10244,N_11009);
nand UO_1309 (O_1309,N_12537,N_11096);
xor UO_1310 (O_1310,N_10487,N_14267);
nor UO_1311 (O_1311,N_13723,N_11499);
or UO_1312 (O_1312,N_14100,N_14864);
xor UO_1313 (O_1313,N_10992,N_10672);
or UO_1314 (O_1314,N_10515,N_12459);
or UO_1315 (O_1315,N_13044,N_12842);
nor UO_1316 (O_1316,N_11837,N_14218);
nand UO_1317 (O_1317,N_12631,N_12521);
and UO_1318 (O_1318,N_12724,N_13691);
or UO_1319 (O_1319,N_14007,N_14844);
nor UO_1320 (O_1320,N_12805,N_13425);
xnor UO_1321 (O_1321,N_13152,N_13085);
nand UO_1322 (O_1322,N_10235,N_13192);
nand UO_1323 (O_1323,N_10756,N_14775);
xnor UO_1324 (O_1324,N_13409,N_14203);
nor UO_1325 (O_1325,N_13560,N_10488);
or UO_1326 (O_1326,N_14995,N_12920);
nand UO_1327 (O_1327,N_10871,N_12272);
nand UO_1328 (O_1328,N_14889,N_10283);
or UO_1329 (O_1329,N_12542,N_11970);
nand UO_1330 (O_1330,N_14631,N_13129);
nor UO_1331 (O_1331,N_12171,N_13709);
nor UO_1332 (O_1332,N_10419,N_12434);
nand UO_1333 (O_1333,N_13139,N_10429);
nand UO_1334 (O_1334,N_11661,N_14487);
or UO_1335 (O_1335,N_14516,N_11279);
or UO_1336 (O_1336,N_14523,N_13681);
and UO_1337 (O_1337,N_14383,N_10964);
or UO_1338 (O_1338,N_14946,N_14578);
xnor UO_1339 (O_1339,N_12648,N_11119);
nor UO_1340 (O_1340,N_14767,N_13056);
nor UO_1341 (O_1341,N_13110,N_10100);
nor UO_1342 (O_1342,N_14172,N_12400);
or UO_1343 (O_1343,N_12356,N_11099);
nor UO_1344 (O_1344,N_12810,N_10163);
xnor UO_1345 (O_1345,N_12408,N_10563);
nand UO_1346 (O_1346,N_11865,N_13431);
nand UO_1347 (O_1347,N_12133,N_14666);
and UO_1348 (O_1348,N_14684,N_10933);
nor UO_1349 (O_1349,N_13018,N_11830);
xnor UO_1350 (O_1350,N_14043,N_12620);
and UO_1351 (O_1351,N_14996,N_14262);
xnor UO_1352 (O_1352,N_13849,N_12482);
xnor UO_1353 (O_1353,N_12420,N_11180);
and UO_1354 (O_1354,N_11419,N_11643);
or UO_1355 (O_1355,N_10299,N_13543);
nand UO_1356 (O_1356,N_11608,N_11652);
nand UO_1357 (O_1357,N_12236,N_10779);
or UO_1358 (O_1358,N_13607,N_14773);
and UO_1359 (O_1359,N_13769,N_11377);
or UO_1360 (O_1360,N_14768,N_11910);
nor UO_1361 (O_1361,N_13368,N_10463);
or UO_1362 (O_1362,N_14645,N_11338);
and UO_1363 (O_1363,N_11308,N_12538);
nand UO_1364 (O_1364,N_12650,N_12467);
nand UO_1365 (O_1365,N_14827,N_12728);
nand UO_1366 (O_1366,N_14982,N_14424);
and UO_1367 (O_1367,N_11844,N_14022);
nor UO_1368 (O_1368,N_10806,N_11438);
xor UO_1369 (O_1369,N_11919,N_14107);
nand UO_1370 (O_1370,N_14213,N_11212);
or UO_1371 (O_1371,N_14940,N_11048);
nor UO_1372 (O_1372,N_13890,N_11976);
nor UO_1373 (O_1373,N_14658,N_14166);
or UO_1374 (O_1374,N_11636,N_12909);
nor UO_1375 (O_1375,N_11944,N_14494);
or UO_1376 (O_1376,N_11664,N_11594);
and UO_1377 (O_1377,N_11110,N_11328);
and UO_1378 (O_1378,N_11575,N_10363);
xnor UO_1379 (O_1379,N_14854,N_13958);
nand UO_1380 (O_1380,N_11317,N_13312);
or UO_1381 (O_1381,N_10785,N_13517);
and UO_1382 (O_1382,N_10815,N_10034);
or UO_1383 (O_1383,N_12142,N_10237);
and UO_1384 (O_1384,N_11684,N_11994);
nor UO_1385 (O_1385,N_10023,N_10775);
and UO_1386 (O_1386,N_11289,N_11909);
xor UO_1387 (O_1387,N_13800,N_14454);
or UO_1388 (O_1388,N_13091,N_10923);
xor UO_1389 (O_1389,N_13588,N_12941);
and UO_1390 (O_1390,N_13821,N_10264);
nand UO_1391 (O_1391,N_10987,N_14911);
nor UO_1392 (O_1392,N_14074,N_10191);
nor UO_1393 (O_1393,N_14749,N_11077);
nand UO_1394 (O_1394,N_11095,N_12239);
nand UO_1395 (O_1395,N_13054,N_12224);
nor UO_1396 (O_1396,N_11333,N_10016);
and UO_1397 (O_1397,N_11147,N_11461);
xor UO_1398 (O_1398,N_10045,N_11082);
xnor UO_1399 (O_1399,N_11118,N_12925);
or UO_1400 (O_1400,N_13138,N_11937);
nor UO_1401 (O_1401,N_11079,N_10307);
or UO_1402 (O_1402,N_10757,N_12077);
nor UO_1403 (O_1403,N_13301,N_10287);
nor UO_1404 (O_1404,N_13628,N_11930);
xor UO_1405 (O_1405,N_12318,N_13650);
xor UO_1406 (O_1406,N_13838,N_13530);
or UO_1407 (O_1407,N_12481,N_11685);
and UO_1408 (O_1408,N_12694,N_13319);
or UO_1409 (O_1409,N_12698,N_14542);
or UO_1410 (O_1410,N_14140,N_13532);
xor UO_1411 (O_1411,N_13227,N_13569);
xnor UO_1412 (O_1412,N_14401,N_11750);
xnor UO_1413 (O_1413,N_14733,N_13631);
nand UO_1414 (O_1414,N_10632,N_11802);
or UO_1415 (O_1415,N_14036,N_13296);
or UO_1416 (O_1416,N_11439,N_13908);
xnor UO_1417 (O_1417,N_14731,N_13830);
or UO_1418 (O_1418,N_12539,N_12574);
or UO_1419 (O_1419,N_11761,N_11704);
and UO_1420 (O_1420,N_13765,N_14136);
nand UO_1421 (O_1421,N_10416,N_14195);
xor UO_1422 (O_1422,N_12243,N_14358);
or UO_1423 (O_1423,N_14452,N_14290);
xor UO_1424 (O_1424,N_14643,N_11628);
or UO_1425 (O_1425,N_13612,N_14264);
and UO_1426 (O_1426,N_13061,N_13069);
or UO_1427 (O_1427,N_11807,N_14687);
and UO_1428 (O_1428,N_13869,N_11496);
xor UO_1429 (O_1429,N_14185,N_10783);
nor UO_1430 (O_1430,N_12752,N_11820);
xnor UO_1431 (O_1431,N_12283,N_11804);
or UO_1432 (O_1432,N_14633,N_14517);
xnor UO_1433 (O_1433,N_10516,N_12630);
xor UO_1434 (O_1434,N_10098,N_11888);
nand UO_1435 (O_1435,N_14840,N_13570);
nand UO_1436 (O_1436,N_12412,N_14619);
nand UO_1437 (O_1437,N_12415,N_10959);
and UO_1438 (O_1438,N_12326,N_14992);
nand UO_1439 (O_1439,N_10065,N_10382);
and UO_1440 (O_1440,N_11939,N_13096);
nor UO_1441 (O_1441,N_10846,N_14964);
and UO_1442 (O_1442,N_13634,N_12718);
nor UO_1443 (O_1443,N_13171,N_10140);
nor UO_1444 (O_1444,N_13496,N_11752);
or UO_1445 (O_1445,N_13361,N_12468);
nor UO_1446 (O_1446,N_13404,N_10086);
nand UO_1447 (O_1447,N_10241,N_11501);
or UO_1448 (O_1448,N_12594,N_10011);
or UO_1449 (O_1449,N_13980,N_13485);
and UO_1450 (O_1450,N_13962,N_12879);
nor UO_1451 (O_1451,N_11758,N_13257);
xor UO_1452 (O_1452,N_13708,N_11586);
xor UO_1453 (O_1453,N_14092,N_10733);
or UO_1454 (O_1454,N_14575,N_14295);
or UO_1455 (O_1455,N_10171,N_13861);
nand UO_1456 (O_1456,N_13494,N_11622);
nor UO_1457 (O_1457,N_12044,N_14199);
and UO_1458 (O_1458,N_11588,N_10742);
nor UO_1459 (O_1459,N_14394,N_10767);
nor UO_1460 (O_1460,N_10503,N_11989);
or UO_1461 (O_1461,N_10184,N_11345);
or UO_1462 (O_1462,N_10528,N_10174);
nor UO_1463 (O_1463,N_14662,N_12819);
xor UO_1464 (O_1464,N_11299,N_11398);
xnor UO_1465 (O_1465,N_12602,N_10232);
nor UO_1466 (O_1466,N_11475,N_11667);
xor UO_1467 (O_1467,N_11932,N_14764);
or UO_1468 (O_1468,N_13501,N_10700);
nand UO_1469 (O_1469,N_13020,N_11811);
xnor UO_1470 (O_1470,N_13931,N_11025);
nor UO_1471 (O_1471,N_14380,N_13989);
and UO_1472 (O_1472,N_13203,N_13261);
or UO_1473 (O_1473,N_10136,N_14493);
nand UO_1474 (O_1474,N_14188,N_14839);
and UO_1475 (O_1475,N_13283,N_13963);
and UO_1476 (O_1476,N_12225,N_14008);
nand UO_1477 (O_1477,N_10804,N_13722);
nand UO_1478 (O_1478,N_10861,N_14207);
xnor UO_1479 (O_1479,N_14372,N_14904);
xnor UO_1480 (O_1480,N_14291,N_13557);
or UO_1481 (O_1481,N_12928,N_11899);
and UO_1482 (O_1482,N_13678,N_12843);
nand UO_1483 (O_1483,N_12649,N_10365);
nor UO_1484 (O_1484,N_14914,N_14301);
nand UO_1485 (O_1485,N_10641,N_13919);
xnor UO_1486 (O_1486,N_10895,N_14495);
or UO_1487 (O_1487,N_10393,N_14071);
xnor UO_1488 (O_1488,N_14284,N_14581);
or UO_1489 (O_1489,N_10650,N_10026);
nor UO_1490 (O_1490,N_10074,N_12460);
xnor UO_1491 (O_1491,N_11776,N_13791);
or UO_1492 (O_1492,N_14674,N_10374);
nor UO_1493 (O_1493,N_11968,N_14759);
nand UO_1494 (O_1494,N_11275,N_11131);
nor UO_1495 (O_1495,N_13286,N_13593);
and UO_1496 (O_1496,N_14919,N_13586);
nor UO_1497 (O_1497,N_13111,N_10787);
xor UO_1498 (O_1498,N_13057,N_11264);
nor UO_1499 (O_1499,N_11557,N_13299);
nor UO_1500 (O_1500,N_11967,N_12697);
nand UO_1501 (O_1501,N_12664,N_12109);
xnor UO_1502 (O_1502,N_13239,N_10120);
and UO_1503 (O_1503,N_13548,N_13209);
xnor UO_1504 (O_1504,N_11123,N_12828);
nor UO_1505 (O_1505,N_11732,N_13794);
and UO_1506 (O_1506,N_10310,N_11235);
and UO_1507 (O_1507,N_10035,N_12074);
and UO_1508 (O_1508,N_12525,N_12927);
xnor UO_1509 (O_1509,N_11581,N_12369);
xnor UO_1510 (O_1510,N_13243,N_13542);
nor UO_1511 (O_1511,N_14925,N_14561);
and UO_1512 (O_1512,N_10906,N_12073);
xor UO_1513 (O_1513,N_12274,N_14386);
xnor UO_1514 (O_1514,N_10540,N_11748);
nor UO_1515 (O_1515,N_14020,N_12138);
and UO_1516 (O_1516,N_13684,N_14918);
and UO_1517 (O_1517,N_13815,N_13099);
xnor UO_1518 (O_1518,N_12279,N_12657);
nor UO_1519 (O_1519,N_12568,N_10438);
xor UO_1520 (O_1520,N_11330,N_10017);
nor UO_1521 (O_1521,N_11319,N_12147);
or UO_1522 (O_1522,N_12208,N_10219);
and UO_1523 (O_1523,N_10714,N_10536);
and UO_1524 (O_1524,N_12807,N_13852);
nor UO_1525 (O_1525,N_11242,N_14706);
and UO_1526 (O_1526,N_12553,N_10547);
nor UO_1527 (O_1527,N_14634,N_10688);
or UO_1528 (O_1528,N_11885,N_14535);
nand UO_1529 (O_1529,N_10315,N_10814);
and UO_1530 (O_1530,N_10997,N_11774);
nand UO_1531 (O_1531,N_10178,N_10473);
or UO_1532 (O_1532,N_14133,N_10255);
nor UO_1533 (O_1533,N_14409,N_11731);
or UO_1534 (O_1534,N_11977,N_11494);
xnor UO_1535 (O_1535,N_13550,N_10912);
nand UO_1536 (O_1536,N_14125,N_11106);
nand UO_1537 (O_1537,N_14246,N_13599);
nor UO_1538 (O_1538,N_11853,N_11431);
nand UO_1539 (O_1539,N_14607,N_12231);
and UO_1540 (O_1540,N_14924,N_11219);
nor UO_1541 (O_1541,N_11332,N_12087);
xor UO_1542 (O_1542,N_13230,N_12042);
or UO_1543 (O_1543,N_11394,N_14711);
and UO_1544 (O_1544,N_11864,N_11546);
xnor UO_1545 (O_1545,N_14470,N_12738);
nor UO_1546 (O_1546,N_12088,N_12395);
nor UO_1547 (O_1547,N_12030,N_14370);
xnor UO_1548 (O_1548,N_12564,N_12093);
nor UO_1549 (O_1549,N_12200,N_10842);
and UO_1550 (O_1550,N_11320,N_12475);
and UO_1551 (O_1551,N_10238,N_13282);
and UO_1552 (O_1552,N_12413,N_10446);
and UO_1553 (O_1553,N_12902,N_14459);
xor UO_1554 (O_1554,N_10654,N_14448);
or UO_1555 (O_1555,N_11854,N_14560);
nand UO_1556 (O_1556,N_12806,N_12255);
and UO_1557 (O_1557,N_11566,N_10585);
xor UO_1558 (O_1558,N_13698,N_11749);
nand UO_1559 (O_1559,N_13101,N_10674);
and UO_1560 (O_1560,N_11740,N_10047);
and UO_1561 (O_1561,N_14557,N_14936);
nor UO_1562 (O_1562,N_11663,N_10057);
nor UO_1563 (O_1563,N_12798,N_12457);
xor UO_1564 (O_1564,N_13567,N_11927);
xnor UO_1565 (O_1565,N_11819,N_12829);
xnor UO_1566 (O_1566,N_12577,N_14701);
or UO_1567 (O_1567,N_10953,N_14664);
nand UO_1568 (O_1568,N_13637,N_10762);
or UO_1569 (O_1569,N_14913,N_13484);
and UO_1570 (O_1570,N_12958,N_12358);
and UO_1571 (O_1571,N_12377,N_10212);
or UO_1572 (O_1572,N_11717,N_12184);
nor UO_1573 (O_1573,N_11509,N_11228);
nor UO_1574 (O_1574,N_13213,N_13596);
nand UO_1575 (O_1575,N_11373,N_14800);
nand UO_1576 (O_1576,N_10543,N_13300);
and UO_1577 (O_1577,N_13945,N_13226);
xor UO_1578 (O_1578,N_12947,N_11781);
and UO_1579 (O_1579,N_14144,N_11288);
and UO_1580 (O_1580,N_11473,N_14181);
nor UO_1581 (O_1581,N_13112,N_10835);
nor UO_1582 (O_1582,N_12403,N_10207);
xnor UO_1583 (O_1583,N_10865,N_11659);
xor UO_1584 (O_1584,N_10328,N_11873);
or UO_1585 (O_1585,N_14312,N_11513);
nor UO_1586 (O_1586,N_14152,N_10567);
nor UO_1587 (O_1587,N_14649,N_13252);
xor UO_1588 (O_1588,N_12285,N_13848);
nor UO_1589 (O_1589,N_11061,N_11011);
and UO_1590 (O_1590,N_14979,N_13370);
and UO_1591 (O_1591,N_12469,N_12004);
or UO_1592 (O_1592,N_11926,N_14004);
xor UO_1593 (O_1593,N_12057,N_14202);
nor UO_1594 (O_1594,N_10290,N_10709);
nand UO_1595 (O_1595,N_12489,N_11483);
or UO_1596 (O_1596,N_13652,N_11270);
or UO_1597 (O_1597,N_14061,N_14342);
nand UO_1598 (O_1598,N_14363,N_11649);
or UO_1599 (O_1599,N_13369,N_13421);
or UO_1600 (O_1600,N_12157,N_12425);
and UO_1601 (O_1601,N_14090,N_13344);
or UO_1602 (O_1602,N_11092,N_10994);
and UO_1603 (O_1603,N_10856,N_13024);
nand UO_1604 (O_1604,N_12132,N_10261);
nor UO_1605 (O_1605,N_12310,N_10262);
nor UO_1606 (O_1606,N_13736,N_13482);
nor UO_1607 (O_1607,N_13168,N_11433);
nor UO_1608 (O_1608,N_12497,N_12191);
or UO_1609 (O_1609,N_14896,N_12229);
nand UO_1610 (O_1610,N_10148,N_11641);
nand UO_1611 (O_1611,N_13499,N_10199);
xnor UO_1612 (O_1612,N_14079,N_13483);
and UO_1613 (O_1613,N_11383,N_13487);
and UO_1614 (O_1614,N_10519,N_11963);
and UO_1615 (O_1615,N_13397,N_12623);
or UO_1616 (O_1616,N_12532,N_11090);
nand UO_1617 (O_1617,N_13704,N_10311);
or UO_1618 (O_1618,N_10530,N_12578);
nand UO_1619 (O_1619,N_10496,N_11053);
xor UO_1620 (O_1620,N_13087,N_14064);
or UO_1621 (O_1621,N_11815,N_11674);
or UO_1622 (O_1622,N_12330,N_14009);
and UO_1623 (O_1623,N_13893,N_10841);
nor UO_1624 (O_1624,N_14817,N_14196);
and UO_1625 (O_1625,N_14293,N_12610);
and UO_1626 (O_1626,N_10931,N_14356);
or UO_1627 (O_1627,N_10301,N_13419);
xnor UO_1628 (O_1628,N_11207,N_11654);
or UO_1629 (O_1629,N_12823,N_12128);
nand UO_1630 (O_1630,N_13400,N_11658);
xnor UO_1631 (O_1631,N_12102,N_11141);
xor UO_1632 (O_1632,N_14192,N_13996);
and UO_1633 (O_1633,N_13563,N_10326);
xor UO_1634 (O_1634,N_11728,N_12461);
xnor UO_1635 (O_1635,N_13933,N_13772);
and UO_1636 (O_1636,N_10561,N_14699);
nor UO_1637 (O_1637,N_12771,N_13127);
or UO_1638 (O_1638,N_12693,N_12556);
and UO_1639 (O_1639,N_12725,N_10272);
xnor UO_1640 (O_1640,N_12636,N_14432);
nand UO_1641 (O_1641,N_10699,N_12494);
and UO_1642 (O_1642,N_14070,N_13725);
nor UO_1643 (O_1643,N_10383,N_13907);
nor UO_1644 (O_1644,N_12571,N_11618);
and UO_1645 (O_1645,N_10614,N_10196);
or UO_1646 (O_1646,N_11456,N_14601);
or UO_1647 (O_1647,N_14745,N_11813);
xnor UO_1648 (O_1648,N_13349,N_10002);
or UO_1649 (O_1649,N_10882,N_10389);
xnor UO_1650 (O_1650,N_11925,N_13073);
and UO_1651 (O_1651,N_12627,N_13674);
and UO_1652 (O_1652,N_11384,N_13256);
and UO_1653 (O_1653,N_10721,N_13221);
xor UO_1654 (O_1654,N_12509,N_12435);
and UO_1655 (O_1655,N_11799,N_14279);
or UO_1656 (O_1656,N_13860,N_13321);
xor UO_1657 (O_1657,N_14670,N_10549);
and UO_1658 (O_1658,N_10637,N_12454);
xnor UO_1659 (O_1659,N_13254,N_10399);
nor UO_1660 (O_1660,N_13746,N_12402);
nor UO_1661 (O_1661,N_11103,N_13808);
xor UO_1662 (O_1662,N_14013,N_12064);
nor UO_1663 (O_1663,N_12629,N_12423);
xnor UO_1664 (O_1664,N_13784,N_11592);
nand UO_1665 (O_1665,N_13799,N_11045);
nor UO_1666 (O_1666,N_13882,N_12441);
nand UO_1667 (O_1667,N_10731,N_12101);
or UO_1668 (O_1668,N_12325,N_14355);
nor UO_1669 (O_1669,N_10044,N_12837);
and UO_1670 (O_1670,N_10558,N_10974);
xor UO_1671 (O_1671,N_11847,N_12802);
nand UO_1672 (O_1672,N_12658,N_14425);
xnor UO_1673 (O_1673,N_14605,N_10725);
and UO_1674 (O_1674,N_14531,N_13867);
nor UO_1675 (O_1675,N_12932,N_11385);
xor UO_1676 (O_1676,N_12316,N_14423);
xnor UO_1677 (O_1677,N_13680,N_13552);
xor UO_1678 (O_1678,N_13128,N_10291);
xnor UO_1679 (O_1679,N_12498,N_13889);
or UO_1680 (O_1680,N_10460,N_14328);
nand UO_1681 (O_1681,N_14966,N_12262);
nand UO_1682 (O_1682,N_14712,N_12121);
nor UO_1683 (O_1683,N_11565,N_14184);
or UO_1684 (O_1684,N_10656,N_11516);
nand UO_1685 (O_1685,N_12182,N_14359);
nand UO_1686 (O_1686,N_12924,N_14399);
or UO_1687 (O_1687,N_12930,N_13518);
nand UO_1688 (O_1688,N_12906,N_11056);
and UO_1689 (O_1689,N_11062,N_11961);
nand UO_1690 (O_1690,N_14884,N_13427);
and UO_1691 (O_1691,N_13219,N_12701);
xnor UO_1692 (O_1692,N_13926,N_14414);
and UO_1693 (O_1693,N_14431,N_12797);
xnor UO_1694 (O_1694,N_14760,N_10888);
xor UO_1695 (O_1695,N_10669,N_10793);
xor UO_1696 (O_1696,N_14451,N_10752);
nand UO_1697 (O_1697,N_13602,N_13520);
or UO_1698 (O_1698,N_12504,N_13474);
nand UO_1699 (O_1699,N_10908,N_12600);
nor UO_1700 (O_1700,N_11999,N_14538);
nor UO_1701 (O_1701,N_13748,N_14615);
xnor UO_1702 (O_1702,N_13624,N_10381);
and UO_1703 (O_1703,N_10911,N_14252);
or UO_1704 (O_1704,N_14628,N_14465);
xnor UO_1705 (O_1705,N_11168,N_14373);
or UO_1706 (O_1706,N_11771,N_10084);
nand UO_1707 (O_1707,N_12785,N_12211);
and UO_1708 (O_1708,N_10670,N_10542);
or UO_1709 (O_1709,N_11187,N_12098);
or UO_1710 (O_1710,N_14528,N_14068);
and UO_1711 (O_1711,N_11343,N_12634);
nand UO_1712 (O_1712,N_14143,N_12001);
nand UO_1713 (O_1713,N_11686,N_10998);
nor UO_1714 (O_1714,N_11913,N_14412);
or UO_1715 (O_1715,N_10606,N_13840);
nor UO_1716 (O_1716,N_11457,N_14242);
nand UO_1717 (O_1717,N_14830,N_11137);
nand UO_1718 (O_1718,N_13918,N_13997);
nor UO_1719 (O_1719,N_11252,N_10589);
xor UO_1720 (O_1720,N_14235,N_13181);
or UO_1721 (O_1721,N_14740,N_14629);
nor UO_1722 (O_1722,N_11127,N_11754);
or UO_1723 (O_1723,N_14294,N_12963);
and UO_1724 (O_1724,N_14336,N_13999);
nor UO_1725 (O_1725,N_10437,N_11160);
nand UO_1726 (O_1726,N_14774,N_10327);
and UO_1727 (O_1727,N_12628,N_11425);
nand UO_1728 (O_1728,N_14239,N_13130);
and UO_1729 (O_1729,N_12226,N_11416);
nand UO_1730 (O_1730,N_13182,N_10910);
or UO_1731 (O_1731,N_14621,N_10692);
xnor UO_1732 (O_1732,N_11202,N_11388);
nand UO_1733 (O_1733,N_14682,N_13339);
and UO_1734 (O_1734,N_13509,N_12957);
nand UO_1735 (O_1735,N_12858,N_14347);
and UO_1736 (O_1736,N_10836,N_11430);
or UO_1737 (O_1737,N_13373,N_13942);
nand UO_1738 (O_1738,N_12841,N_12129);
nand UO_1739 (O_1739,N_13731,N_13303);
and UO_1740 (O_1740,N_13778,N_12382);
or UO_1741 (O_1741,N_12217,N_14224);
or UO_1742 (O_1742,N_12131,N_14794);
xnor UO_1743 (O_1743,N_13797,N_11706);
and UO_1744 (O_1744,N_12536,N_12327);
and UO_1745 (O_1745,N_10855,N_14164);
or UO_1746 (O_1746,N_12178,N_11158);
and UO_1747 (O_1747,N_11604,N_10664);
or UO_1748 (O_1748,N_13786,N_11719);
nand UO_1749 (O_1749,N_14420,N_12713);
xnor UO_1750 (O_1750,N_14056,N_12348);
and UO_1751 (O_1751,N_11969,N_14031);
xor UO_1752 (O_1752,N_10952,N_14527);
xor UO_1753 (O_1753,N_13173,N_13244);
and UO_1754 (O_1754,N_14225,N_10031);
nor UO_1755 (O_1755,N_11109,N_14570);
xnor UO_1756 (O_1756,N_11441,N_12159);
xnor UO_1757 (O_1757,N_13016,N_11153);
xnor UO_1758 (O_1758,N_10697,N_12667);
nand UO_1759 (O_1759,N_10509,N_10642);
xnor UO_1760 (O_1760,N_14769,N_12393);
nand UO_1761 (O_1761,N_13250,N_11808);
or UO_1762 (O_1762,N_13422,N_11848);
or UO_1763 (O_1763,N_13294,N_11696);
nand UO_1764 (O_1764,N_14565,N_14479);
nor UO_1765 (O_1765,N_14103,N_12091);
or UO_1766 (O_1766,N_11327,N_12669);
and UO_1767 (O_1767,N_13147,N_11370);
nand UO_1768 (O_1768,N_14562,N_12820);
and UO_1769 (O_1769,N_13158,N_14825);
xor UO_1770 (O_1770,N_13706,N_14053);
and UO_1771 (O_1771,N_12961,N_10211);
nand UO_1772 (O_1772,N_12379,N_11294);
and UO_1773 (O_1773,N_11894,N_12964);
nor UO_1774 (O_1774,N_11959,N_13738);
nand UO_1775 (O_1775,N_10693,N_13218);
or UO_1776 (O_1776,N_12410,N_10555);
xor UO_1777 (O_1777,N_11254,N_12548);
xor UO_1778 (O_1778,N_10145,N_14116);
nor UO_1779 (O_1779,N_12891,N_10286);
or UO_1780 (O_1780,N_12110,N_14400);
or UO_1781 (O_1781,N_11599,N_10091);
nor UO_1782 (O_1782,N_13275,N_10898);
xnor UO_1783 (O_1783,N_10202,N_12181);
nand UO_1784 (O_1784,N_14438,N_10763);
nor UO_1785 (O_1785,N_13916,N_14326);
or UO_1786 (O_1786,N_11412,N_13297);
xnor UO_1787 (O_1787,N_10114,N_10724);
nand UO_1788 (O_1788,N_12297,N_13452);
xnor UO_1789 (O_1789,N_14917,N_11074);
nor UO_1790 (O_1790,N_12735,N_10008);
nand UO_1791 (O_1791,N_10620,N_10829);
nand UO_1792 (O_1792,N_12678,N_12240);
or UO_1793 (O_1793,N_11638,N_14477);
xor UO_1794 (O_1794,N_14948,N_10368);
and UO_1795 (O_1795,N_12749,N_14929);
nor UO_1796 (O_1796,N_13318,N_14907);
nand UO_1797 (O_1797,N_11955,N_14299);
nor UO_1798 (O_1798,N_14876,N_12167);
nor UO_1799 (O_1799,N_12519,N_13406);
nor UO_1800 (O_1800,N_11368,N_14165);
xor UO_1801 (O_1801,N_13424,N_13690);
and UO_1802 (O_1802,N_13212,N_14415);
and UO_1803 (O_1803,N_14076,N_10060);
nor UO_1804 (O_1804,N_11142,N_10771);
or UO_1805 (O_1805,N_13208,N_12158);
or UO_1806 (O_1806,N_12660,N_11931);
nand UO_1807 (O_1807,N_13246,N_11067);
xnor UO_1808 (O_1808,N_10124,N_10765);
and UO_1809 (O_1809,N_14285,N_13526);
xnor UO_1810 (O_1810,N_11640,N_13573);
xnor UO_1811 (O_1811,N_14534,N_10971);
and UO_1812 (O_1812,N_14810,N_12144);
and UO_1813 (O_1813,N_12867,N_12756);
xnor UO_1814 (O_1814,N_12233,N_11113);
nor UO_1815 (O_1815,N_10464,N_12605);
or UO_1816 (O_1816,N_12107,N_11601);
or UO_1817 (O_1817,N_12546,N_13773);
nand UO_1818 (O_1818,N_13153,N_14440);
nor UO_1819 (O_1819,N_13047,N_14258);
xnor UO_1820 (O_1820,N_12817,N_10747);
or UO_1821 (O_1821,N_11000,N_11528);
xnor UO_1822 (O_1822,N_13592,N_10817);
xor UO_1823 (O_1823,N_14384,N_14632);
or UO_1824 (O_1824,N_10472,N_12137);
and UO_1825 (O_1825,N_13825,N_10110);
and UO_1826 (O_1826,N_10520,N_14897);
nor UO_1827 (O_1827,N_14965,N_11634);
xor UO_1828 (O_1828,N_11101,N_10030);
nor UO_1829 (O_1829,N_13987,N_11852);
xor UO_1830 (O_1830,N_12237,N_13611);
or UO_1831 (O_1831,N_12066,N_13724);
or UO_1832 (O_1832,N_10899,N_11449);
xnor UO_1833 (O_1833,N_10405,N_14950);
and UO_1834 (O_1834,N_10059,N_11139);
xnor UO_1835 (O_1835,N_10655,N_11311);
or UO_1836 (O_1836,N_14187,N_11507);
or UO_1837 (O_1837,N_14506,N_11429);
or UO_1838 (O_1838,N_13643,N_10574);
and UO_1839 (O_1839,N_10159,N_12507);
nor UO_1840 (O_1840,N_10162,N_14757);
or UO_1841 (O_1841,N_13177,N_10965);
xor UO_1842 (O_1842,N_11633,N_13357);
nor UO_1843 (O_1843,N_12573,N_10033);
nor UO_1844 (O_1844,N_12323,N_14795);
or UO_1845 (O_1845,N_10827,N_14318);
nand UO_1846 (O_1846,N_12011,N_12154);
nor UO_1847 (O_1847,N_13752,N_12543);
and UO_1848 (O_1848,N_13923,N_11635);
and UO_1849 (O_1849,N_13225,N_13335);
and UO_1850 (O_1850,N_12282,N_12933);
nand UO_1851 (O_1851,N_11741,N_14364);
xor UO_1852 (O_1852,N_10541,N_12615);
nor UO_1853 (O_1853,N_11274,N_10792);
and UO_1854 (O_1854,N_12426,N_12576);
nor UO_1855 (O_1855,N_11531,N_11208);
and UO_1856 (O_1856,N_10330,N_14908);
and UO_1857 (O_1857,N_10705,N_14115);
nor UO_1858 (O_1858,N_10180,N_13378);
or UO_1859 (O_1859,N_12848,N_13971);
or UO_1860 (O_1860,N_13914,N_14978);
nand UO_1861 (O_1861,N_11195,N_11974);
or UO_1862 (O_1862,N_14891,N_12606);
nand UO_1863 (O_1863,N_10351,N_10873);
or UO_1864 (O_1864,N_11315,N_12897);
xor UO_1865 (O_1865,N_11827,N_14533);
and UO_1866 (O_1866,N_14872,N_12298);
or UO_1867 (O_1867,N_11574,N_11019);
nand UO_1868 (O_1868,N_10415,N_12816);
nor UO_1869 (O_1869,N_10094,N_12291);
xor UO_1870 (O_1870,N_14568,N_10322);
or UO_1871 (O_1871,N_14331,N_14357);
and UO_1872 (O_1872,N_11223,N_14416);
xor UO_1873 (O_1873,N_12917,N_13382);
nand UO_1874 (O_1874,N_13766,N_10754);
and UO_1875 (O_1875,N_11672,N_13833);
xnor UO_1876 (O_1876,N_13842,N_14082);
or UO_1877 (O_1877,N_14921,N_10649);
nor UO_1878 (O_1878,N_14017,N_10492);
xor UO_1879 (O_1879,N_12840,N_11140);
or UO_1880 (O_1880,N_14354,N_11492);
xnor UO_1881 (O_1881,N_11850,N_10624);
nand UO_1882 (O_1882,N_10960,N_14102);
or UO_1883 (O_1883,N_14190,N_10006);
nand UO_1884 (O_1884,N_11670,N_13749);
or UO_1885 (O_1885,N_12898,N_11736);
nor UO_1886 (O_1886,N_10534,N_13143);
nor UO_1887 (O_1887,N_11515,N_13630);
nand UO_1888 (O_1888,N_11094,N_14077);
and UO_1889 (O_1889,N_12339,N_13554);
and UO_1890 (O_1890,N_10188,N_10893);
and UO_1891 (O_1891,N_10781,N_13537);
nor UO_1892 (O_1892,N_10851,N_13693);
nand UO_1893 (O_1893,N_12722,N_12201);
nand UO_1894 (O_1894,N_13412,N_12068);
nor UO_1895 (O_1895,N_11716,N_12428);
and UO_1896 (O_1896,N_12510,N_12654);
or UO_1897 (O_1897,N_12270,N_13613);
nor UO_1898 (O_1898,N_10810,N_13032);
or UO_1899 (O_1899,N_12115,N_12717);
nor UO_1900 (O_1900,N_12268,N_13935);
nor UO_1901 (O_1901,N_13398,N_14718);
xor UO_1902 (O_1902,N_10639,N_12931);
and UO_1903 (O_1903,N_12511,N_14179);
or UO_1904 (O_1904,N_14091,N_10347);
and UO_1905 (O_1905,N_12890,N_10056);
and UO_1906 (O_1906,N_14296,N_12892);
xnor UO_1907 (O_1907,N_12626,N_11276);
nor UO_1908 (O_1908,N_14798,N_12719);
xnor UO_1909 (O_1909,N_10601,N_14216);
or UO_1910 (O_1910,N_10562,N_14182);
and UO_1911 (O_1911,N_14536,N_11292);
nand UO_1912 (O_1912,N_10640,N_10979);
nor UO_1913 (O_1913,N_11693,N_11031);
or UO_1914 (O_1914,N_13506,N_12025);
nand UO_1915 (O_1915,N_11358,N_13523);
nor UO_1916 (O_1916,N_10093,N_11181);
nand UO_1917 (O_1917,N_13870,N_11297);
nor UO_1918 (O_1918,N_14805,N_10951);
nor UO_1919 (O_1919,N_12624,N_12366);
and UO_1920 (O_1920,N_12775,N_12789);
and UO_1921 (O_1921,N_12795,N_10876);
xor UO_1922 (O_1922,N_11381,N_13696);
and UO_1923 (O_1923,N_10379,N_13820);
nand UO_1924 (O_1924,N_13995,N_11017);
nand UO_1925 (O_1925,N_14938,N_11277);
xnor UO_1926 (O_1926,N_13885,N_13555);
or UO_1927 (O_1927,N_13587,N_13451);
xnor UO_1928 (O_1928,N_14916,N_11992);
and UO_1929 (O_1929,N_14112,N_14272);
or UO_1930 (O_1930,N_11214,N_14890);
nor UO_1931 (O_1931,N_12195,N_14821);
nand UO_1932 (O_1932,N_11710,N_12882);
and UO_1933 (O_1933,N_11921,N_14724);
or UO_1934 (O_1934,N_14121,N_10726);
nor UO_1935 (O_1935,N_12164,N_14023);
and UO_1936 (O_1936,N_10704,N_12907);
xor UO_1937 (O_1937,N_13408,N_13385);
and UO_1938 (O_1938,N_10482,N_11243);
and UO_1939 (O_1939,N_11354,N_12409);
and UO_1940 (O_1940,N_14667,N_10811);
nor UO_1941 (O_1941,N_14529,N_12357);
xnor UO_1942 (O_1942,N_11326,N_12444);
and UO_1943 (O_1943,N_11108,N_11232);
nand UO_1944 (O_1944,N_11500,N_11780);
and UO_1945 (O_1945,N_11609,N_11539);
xor UO_1946 (O_1946,N_13589,N_13846);
or UO_1947 (O_1947,N_11986,N_12776);
xor UO_1948 (O_1948,N_11883,N_11054);
or UO_1949 (O_1949,N_12633,N_12547);
xnor UO_1950 (O_1950,N_14947,N_11996);
nor UO_1951 (O_1951,N_12244,N_11655);
nand UO_1952 (O_1952,N_12540,N_12976);
nand UO_1953 (O_1953,N_10738,N_11367);
or UO_1954 (O_1954,N_12988,N_14861);
nand UO_1955 (O_1955,N_12452,N_12047);
and UO_1956 (O_1956,N_11798,N_13015);
nand UO_1957 (O_1957,N_12281,N_10698);
xnor UO_1958 (O_1958,N_10768,N_13134);
xor UO_1959 (O_1959,N_11603,N_14548);
nor UO_1960 (O_1960,N_14138,N_10325);
or UO_1961 (O_1961,N_11083,N_14047);
nor UO_1962 (O_1962,N_12712,N_11606);
and UO_1963 (O_1963,N_10097,N_12832);
or UO_1964 (O_1964,N_13381,N_13783);
or UO_1965 (O_1965,N_11564,N_14122);
nor UO_1966 (O_1966,N_13998,N_13041);
nor UO_1967 (O_1967,N_12305,N_12955);
xor UO_1968 (O_1968,N_13010,N_12878);
nor UO_1969 (O_1969,N_13853,N_12551);
nand UO_1970 (O_1970,N_11397,N_10954);
nand UO_1971 (O_1971,N_13959,N_10303);
and UO_1972 (O_1972,N_10741,N_10812);
nand UO_1973 (O_1973,N_10584,N_13437);
nor UO_1974 (O_1974,N_12954,N_14439);
or UO_1975 (O_1975,N_14374,N_11923);
or UO_1976 (O_1976,N_11933,N_11532);
or UO_1977 (O_1977,N_11051,N_13540);
xnor UO_1978 (O_1978,N_14863,N_14250);
nand UO_1979 (O_1979,N_13435,N_12390);
nor UO_1980 (O_1980,N_14503,N_13396);
and UO_1981 (O_1981,N_13271,N_12565);
and UO_1982 (O_1982,N_13392,N_14129);
and UO_1983 (O_1983,N_11510,N_10678);
or UO_1984 (O_1984,N_14069,N_14859);
and UO_1985 (O_1985,N_13317,N_13331);
and UO_1986 (O_1986,N_14685,N_12940);
nand UO_1987 (O_1987,N_13434,N_11250);
and UO_1988 (O_1988,N_10570,N_11012);
or UO_1989 (O_1989,N_14178,N_10909);
and UO_1990 (O_1990,N_11100,N_11306);
xor UO_1991 (O_1991,N_10495,N_14443);
nor UO_1992 (O_1992,N_13739,N_12801);
nor UO_1993 (O_1993,N_14955,N_12092);
nand UO_1994 (O_1994,N_13854,N_11364);
xor UO_1995 (O_1995,N_12146,N_11251);
or UO_1996 (O_1996,N_13675,N_14647);
and UO_1997 (O_1997,N_14086,N_13750);
and UO_1998 (O_1998,N_10713,N_12856);
xnor UO_1999 (O_1999,N_12389,N_10840);
endmodule