module basic_3000_30000_3500_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_2613,In_1774);
or U1 (N_1,In_452,In_2670);
xor U2 (N_2,In_2057,In_1304);
nor U3 (N_3,In_1301,In_1563);
or U4 (N_4,In_1213,In_437);
nor U5 (N_5,In_317,In_494);
xnor U6 (N_6,In_792,In_314);
xnor U7 (N_7,In_2876,In_1222);
or U8 (N_8,In_1165,In_323);
and U9 (N_9,In_1299,In_1977);
nand U10 (N_10,In_1532,In_143);
and U11 (N_11,In_846,In_1620);
and U12 (N_12,In_2986,In_1993);
nand U13 (N_13,In_891,In_775);
nand U14 (N_14,In_1107,In_1290);
nor U15 (N_15,In_2025,In_326);
or U16 (N_16,In_49,In_255);
nor U17 (N_17,In_1007,In_245);
or U18 (N_18,In_496,In_926);
or U19 (N_19,In_2354,In_916);
and U20 (N_20,In_1410,In_1362);
nand U21 (N_21,In_996,In_301);
nand U22 (N_22,In_2940,In_1281);
or U23 (N_23,In_1363,In_2409);
and U24 (N_24,In_2496,In_1258);
xnor U25 (N_25,In_2120,In_2746);
nand U26 (N_26,In_1442,In_2173);
and U27 (N_27,In_1921,In_2256);
nor U28 (N_28,In_666,In_827);
nor U29 (N_29,In_2890,In_1776);
or U30 (N_30,In_1636,In_2930);
nor U31 (N_31,In_1322,In_2901);
xnor U32 (N_32,In_346,In_1238);
xnor U33 (N_33,In_2919,In_1925);
xnor U34 (N_34,In_1690,In_462);
and U35 (N_35,In_1012,In_1973);
and U36 (N_36,In_2547,In_2064);
nor U37 (N_37,In_473,In_431);
nand U38 (N_38,In_2703,In_1495);
xnor U39 (N_39,In_1090,In_2536);
and U40 (N_40,In_119,In_399);
nor U41 (N_41,In_757,In_2880);
and U42 (N_42,In_651,In_116);
nor U43 (N_43,In_2846,In_2101);
xnor U44 (N_44,In_1556,In_1202);
and U45 (N_45,In_1315,In_637);
nor U46 (N_46,In_2809,In_2794);
nor U47 (N_47,In_1338,In_1072);
or U48 (N_48,In_2187,In_1807);
and U49 (N_49,In_1560,In_930);
xor U50 (N_50,In_1276,In_2380);
or U51 (N_51,In_2356,In_2340);
xnor U52 (N_52,In_2068,In_1537);
or U53 (N_53,In_2122,In_244);
or U54 (N_54,In_952,In_2322);
xnor U55 (N_55,In_2648,In_25);
or U56 (N_56,In_2121,In_921);
nand U57 (N_57,In_1475,In_1724);
or U58 (N_58,In_980,In_1573);
nand U59 (N_59,In_2130,In_389);
nor U60 (N_60,In_1637,In_1097);
nand U61 (N_61,In_2126,In_1397);
or U62 (N_62,In_497,In_2820);
xnor U63 (N_63,In_966,In_2338);
xnor U64 (N_64,In_1113,In_773);
or U65 (N_65,In_1520,In_2395);
or U66 (N_66,In_2615,In_36);
nand U67 (N_67,In_285,In_1866);
nand U68 (N_68,In_1132,In_768);
nor U69 (N_69,In_2567,In_2543);
nor U70 (N_70,In_467,In_2574);
nand U71 (N_71,In_228,In_2517);
or U72 (N_72,In_1353,In_1896);
nor U73 (N_73,In_2381,In_531);
and U74 (N_74,In_1590,In_2302);
xnor U75 (N_75,In_1820,In_2365);
xnor U76 (N_76,In_1427,In_2610);
xnor U77 (N_77,In_2294,In_2323);
xnor U78 (N_78,In_2072,In_2956);
or U79 (N_79,In_2359,In_900);
xnor U80 (N_80,In_1508,In_912);
nand U81 (N_81,In_1572,In_1752);
or U82 (N_82,In_733,In_684);
or U83 (N_83,In_129,In_937);
and U84 (N_84,In_587,In_2628);
nand U85 (N_85,In_1576,In_2282);
xnor U86 (N_86,In_483,In_2114);
nor U87 (N_87,In_799,In_2328);
nor U88 (N_88,In_130,In_923);
xor U89 (N_89,In_1310,In_1382);
nor U90 (N_90,In_72,In_753);
xor U91 (N_91,In_2065,In_1792);
or U92 (N_92,In_2784,In_2046);
nor U93 (N_93,In_93,In_974);
or U94 (N_94,In_374,In_2935);
or U95 (N_95,In_2433,In_153);
nor U96 (N_96,In_464,In_1611);
or U97 (N_97,In_2842,In_2324);
xnor U98 (N_98,In_2619,In_226);
xor U99 (N_99,In_1278,In_216);
nand U100 (N_100,In_721,In_85);
xor U101 (N_101,In_2898,In_1340);
or U102 (N_102,In_2688,In_927);
or U103 (N_103,In_298,In_2560);
and U104 (N_104,In_669,In_2894);
and U105 (N_105,In_1229,In_895);
and U106 (N_106,In_1519,In_2806);
nor U107 (N_107,In_2127,In_1142);
xor U108 (N_108,In_1302,In_875);
and U109 (N_109,In_267,In_2247);
and U110 (N_110,In_533,In_2136);
nand U111 (N_111,In_2280,In_199);
nor U112 (N_112,In_2421,In_788);
xor U113 (N_113,In_689,In_466);
nand U114 (N_114,In_2048,In_2822);
xor U115 (N_115,In_99,In_2885);
xnor U116 (N_116,In_1806,In_1504);
xnor U117 (N_117,In_2993,In_2737);
or U118 (N_118,In_2344,In_1974);
xor U119 (N_119,In_2633,In_7);
xor U120 (N_120,In_113,In_2316);
or U121 (N_121,In_140,In_2519);
nor U122 (N_122,In_1393,In_353);
nor U123 (N_123,In_1147,In_1470);
xor U124 (N_124,In_1250,In_1023);
xor U125 (N_125,In_2914,In_370);
nor U126 (N_126,In_260,In_1742);
nor U127 (N_127,In_740,In_1755);
xnor U128 (N_128,In_1188,In_984);
and U129 (N_129,In_273,In_2570);
nand U130 (N_130,In_1610,In_658);
or U131 (N_131,In_2830,In_2755);
xnor U132 (N_132,In_2478,In_627);
and U133 (N_133,In_1145,In_280);
nand U134 (N_134,In_2321,In_2471);
or U135 (N_135,In_2577,In_866);
nand U136 (N_136,In_1359,In_2531);
or U137 (N_137,In_232,In_779);
nand U138 (N_138,In_2873,In_1294);
nor U139 (N_139,In_2699,In_1196);
and U140 (N_140,In_2659,In_2334);
xor U141 (N_141,In_1515,In_201);
and U142 (N_142,In_748,In_1476);
and U143 (N_143,In_1837,In_871);
xor U144 (N_144,In_565,In_1488);
nor U145 (N_145,In_206,In_447);
nor U146 (N_146,In_137,In_2618);
and U147 (N_147,In_547,In_213);
xor U148 (N_148,In_1168,In_536);
nor U149 (N_149,In_215,In_606);
and U150 (N_150,In_1571,In_2936);
nand U151 (N_151,In_2203,In_1986);
xnor U152 (N_152,In_1800,In_2535);
nor U153 (N_153,In_1564,In_2530);
and U154 (N_154,In_2954,In_2129);
and U155 (N_155,In_1779,In_732);
xor U156 (N_156,In_2310,In_2337);
nand U157 (N_157,In_221,In_908);
or U158 (N_158,In_805,In_1935);
xnor U159 (N_159,In_1034,In_1481);
xnor U160 (N_160,In_1371,In_986);
nor U161 (N_161,In_1492,In_1331);
xnor U162 (N_162,In_1005,In_331);
and U163 (N_163,In_697,In_1201);
nand U164 (N_164,In_60,In_582);
and U165 (N_165,In_2398,In_1497);
xnor U166 (N_166,In_2408,In_180);
nand U167 (N_167,In_901,In_1084);
xnor U168 (N_168,In_959,In_870);
xnor U169 (N_169,In_555,In_2874);
nand U170 (N_170,In_537,In_2288);
nand U171 (N_171,In_30,In_205);
xor U172 (N_172,In_120,In_2541);
xnor U173 (N_173,In_2858,In_964);
nor U174 (N_174,In_997,In_2372);
or U175 (N_175,In_2695,In_2027);
nand U176 (N_176,In_2985,In_2386);
and U177 (N_177,In_106,In_1681);
and U178 (N_178,In_1428,In_1711);
or U179 (N_179,In_1098,In_279);
nor U180 (N_180,In_2532,In_806);
nand U181 (N_181,In_1916,In_39);
xnor U182 (N_182,In_1862,In_2810);
and U183 (N_183,In_807,In_1698);
nand U184 (N_184,In_967,In_653);
nand U185 (N_185,In_214,In_2839);
xnor U186 (N_186,In_1295,In_628);
nor U187 (N_187,In_736,In_530);
xnor U188 (N_188,In_1272,In_1691);
xor U189 (N_189,In_1087,In_1646);
nor U190 (N_190,In_1709,In_1255);
and U191 (N_191,In_2815,In_404);
nand U192 (N_192,In_524,In_269);
nor U193 (N_193,In_64,In_29);
and U194 (N_194,In_1618,In_152);
nor U195 (N_195,In_1119,In_2825);
or U196 (N_196,In_1979,In_300);
or U197 (N_197,In_2934,In_1829);
nand U198 (N_198,In_2491,In_2732);
and U199 (N_199,In_2791,In_2616);
or U200 (N_200,In_1326,In_821);
nand U201 (N_201,In_2399,In_763);
xor U202 (N_202,In_1863,In_1642);
or U203 (N_203,In_418,In_1152);
nor U204 (N_204,In_1289,In_1104);
and U205 (N_205,In_1786,In_82);
xnor U206 (N_206,In_1581,In_1805);
or U207 (N_207,In_1163,In_1205);
nand U208 (N_208,In_1040,In_2492);
nor U209 (N_209,In_946,In_1624);
nor U210 (N_210,In_2933,In_2331);
nand U211 (N_211,In_2201,In_321);
nor U212 (N_212,In_1924,In_1670);
or U213 (N_213,In_2745,In_957);
xor U214 (N_214,In_2772,In_2039);
nor U215 (N_215,In_667,In_1985);
nand U216 (N_216,In_1230,In_1035);
xnor U217 (N_217,In_2859,In_2342);
or U218 (N_218,In_713,In_1682);
or U219 (N_219,In_2229,In_892);
xnor U220 (N_220,In_924,In_161);
nor U221 (N_221,In_2812,In_415);
nand U222 (N_222,In_1426,In_2961);
or U223 (N_223,In_1417,In_1419);
or U224 (N_224,In_746,In_1700);
or U225 (N_225,In_2474,In_1489);
xor U226 (N_226,In_74,In_2098);
nor U227 (N_227,In_227,In_2569);
xor U228 (N_228,In_1607,In_434);
and U229 (N_229,In_1844,In_2175);
and U230 (N_230,In_1180,In_1915);
nor U231 (N_231,In_554,In_881);
nor U232 (N_232,In_1514,In_797);
or U233 (N_233,In_737,In_1044);
and U234 (N_234,In_2724,In_1403);
xnor U235 (N_235,In_1297,In_274);
or U236 (N_236,In_936,In_481);
nand U237 (N_237,In_2438,In_1432);
nand U238 (N_238,In_1587,In_802);
or U239 (N_239,In_2587,In_2694);
nand U240 (N_240,In_2414,In_2038);
nor U241 (N_241,In_864,In_249);
nor U242 (N_242,In_499,In_994);
and U243 (N_243,In_1812,In_1178);
nor U244 (N_244,In_2786,In_1194);
and U245 (N_245,In_1365,In_2514);
nand U246 (N_246,In_63,In_1283);
or U247 (N_247,In_1830,In_1968);
nand U248 (N_248,In_1982,In_250);
nand U249 (N_249,In_630,In_2184);
nand U250 (N_250,In_1684,In_508);
and U251 (N_251,In_1341,In_2459);
nand U252 (N_252,In_1370,In_1659);
and U253 (N_253,In_2895,In_687);
nor U254 (N_254,In_822,In_2768);
or U255 (N_255,In_2738,In_2050);
xor U256 (N_256,In_2009,In_2457);
or U257 (N_257,In_2693,In_192);
or U258 (N_258,In_2036,In_789);
and U259 (N_259,In_174,In_2697);
or U260 (N_260,In_1860,In_2000);
xor U261 (N_261,In_1022,In_1274);
xor U262 (N_262,In_2702,In_887);
or U263 (N_263,In_2070,In_2712);
and U264 (N_264,In_634,In_1790);
nand U265 (N_265,In_1667,In_449);
or U266 (N_266,In_1754,In_2405);
or U267 (N_267,In_2219,In_826);
or U268 (N_268,In_294,In_1498);
and U269 (N_269,In_1789,In_1591);
nor U270 (N_270,In_756,In_2726);
or U271 (N_271,In_1686,In_1373);
and U272 (N_272,In_236,In_2634);
xor U273 (N_273,In_1368,In_1533);
xnor U274 (N_274,In_2042,In_1601);
or U275 (N_275,In_445,In_2018);
nor U276 (N_276,In_1028,In_1396);
nor U277 (N_277,In_1160,In_2889);
and U278 (N_278,In_816,In_1893);
or U279 (N_279,In_865,In_2888);
and U280 (N_280,In_1989,In_2540);
nor U281 (N_281,In_2290,In_1017);
xnor U282 (N_282,In_626,In_2100);
or U283 (N_283,In_2720,In_2758);
xnor U284 (N_284,In_296,In_421);
nor U285 (N_285,In_2678,In_2976);
xor U286 (N_286,In_2905,In_81);
nand U287 (N_287,In_411,In_714);
and U288 (N_288,In_2987,In_1004);
nor U289 (N_289,In_2106,In_1019);
or U290 (N_290,In_2581,In_117);
and U291 (N_291,In_1951,In_1816);
or U292 (N_292,In_1437,In_831);
or U293 (N_293,In_904,In_2361);
and U294 (N_294,In_1161,In_334);
and U295 (N_295,In_2411,In_193);
nand U296 (N_296,In_929,In_956);
and U297 (N_297,In_2651,In_1027);
xnor U298 (N_298,In_1981,In_2595);
nand U299 (N_299,In_1286,In_61);
nor U300 (N_300,In_890,In_240);
and U301 (N_301,In_2230,In_278);
xor U302 (N_302,In_2488,In_2146);
nand U303 (N_303,In_1772,In_2379);
xor U304 (N_304,In_69,In_1568);
nand U305 (N_305,In_2441,In_2061);
nor U306 (N_306,In_2447,In_124);
or U307 (N_307,In_2661,In_632);
and U308 (N_308,In_1833,In_1894);
xor U309 (N_309,In_730,In_2892);
nand U310 (N_310,In_2609,In_869);
and U311 (N_311,In_2505,In_1224);
and U312 (N_312,In_585,In_2151);
or U313 (N_313,In_2495,In_2104);
or U314 (N_314,In_2736,In_899);
xnor U315 (N_315,In_1324,In_2960);
nor U316 (N_316,In_1562,In_1386);
or U317 (N_317,In_2824,In_1821);
nand U318 (N_318,In_2979,In_231);
nor U319 (N_319,In_1727,In_2903);
and U320 (N_320,In_151,In_2019);
nand U321 (N_321,In_770,In_1357);
xor U322 (N_322,In_2387,In_2617);
or U323 (N_323,In_2965,In_2705);
and U324 (N_324,In_694,In_2177);
xor U325 (N_325,In_1360,In_1094);
and U326 (N_326,In_1809,In_1057);
nand U327 (N_327,In_2133,In_1333);
nor U328 (N_328,In_1538,In_1268);
nor U329 (N_329,In_862,In_1960);
nand U330 (N_330,In_2152,In_1988);
nor U331 (N_331,In_2029,In_828);
nor U332 (N_332,In_1660,In_2578);
and U333 (N_333,In_903,In_2170);
nand U334 (N_334,In_1192,In_325);
nand U335 (N_335,In_849,In_917);
or U336 (N_336,In_2958,In_87);
nor U337 (N_337,In_1871,In_575);
and U338 (N_338,In_2226,In_1720);
xor U339 (N_339,In_1743,In_928);
xnor U340 (N_340,In_2742,In_1485);
nand U341 (N_341,In_1158,In_1701);
xnor U342 (N_342,In_2805,In_1856);
or U343 (N_343,In_332,In_175);
and U344 (N_344,In_148,In_1190);
nand U345 (N_345,In_2326,In_1053);
or U346 (N_346,In_112,In_600);
nor U347 (N_347,In_2434,In_622);
xor U348 (N_348,In_1950,In_933);
xor U349 (N_349,In_1100,In_1352);
nor U350 (N_350,In_2816,In_2969);
or U351 (N_351,In_2223,In_409);
nand U352 (N_352,In_2545,In_2026);
xnor U353 (N_353,In_2868,In_2924);
or U354 (N_354,In_1399,In_611);
and U355 (N_355,In_2467,In_2483);
xor U356 (N_356,In_97,In_1814);
nand U357 (N_357,In_2708,In_1557);
nor U358 (N_358,In_2717,In_882);
and U359 (N_359,In_2948,In_1630);
and U360 (N_360,In_2573,In_2682);
nor U361 (N_361,In_1101,In_2207);
or U362 (N_362,In_719,In_2067);
and U363 (N_363,In_682,In_2896);
xnor U364 (N_364,In_2358,In_144);
nand U365 (N_365,In_44,In_160);
and U366 (N_366,In_2733,In_1169);
nand U367 (N_367,In_686,In_982);
or U368 (N_368,In_2507,In_659);
and U369 (N_369,In_2729,In_1884);
and U370 (N_370,In_1699,In_454);
nor U371 (N_371,In_2761,In_1995);
and U372 (N_372,In_2611,In_2283);
xnor U373 (N_373,In_413,In_561);
and U374 (N_374,In_2041,In_776);
and U375 (N_375,In_506,In_2240);
nand U376 (N_376,In_2298,In_425);
and U377 (N_377,In_1773,In_2652);
nand U378 (N_378,In_1599,In_1832);
nand U379 (N_379,In_121,In_1957);
or U380 (N_380,In_765,In_2676);
or U381 (N_381,In_2268,In_2900);
xnor U382 (N_382,In_2826,In_2576);
or U383 (N_383,In_1459,In_2266);
xor U384 (N_384,In_1940,In_366);
and U385 (N_385,In_873,In_1211);
xor U386 (N_386,In_1509,In_79);
xnor U387 (N_387,In_2456,In_1140);
nand U388 (N_388,In_2464,In_1579);
nand U389 (N_389,In_2232,In_2345);
nand U390 (N_390,In_1512,In_1947);
xnor U391 (N_391,In_396,In_1273);
and U392 (N_392,In_1962,In_1162);
or U393 (N_393,In_1298,In_1282);
xnor U394 (N_394,In_704,In_2550);
nand U395 (N_395,In_1285,In_1823);
and U396 (N_396,In_975,In_1206);
nor U397 (N_397,In_2202,In_1505);
or U398 (N_398,In_179,In_222);
nor U399 (N_399,In_73,In_2950);
nand U400 (N_400,In_1600,In_2484);
nand U401 (N_401,In_1850,In_2557);
nand U402 (N_402,In_1455,In_1483);
xnor U403 (N_403,In_868,In_344);
xnor U404 (N_404,In_141,In_1409);
nor U405 (N_405,In_2886,In_203);
or U406 (N_406,In_1262,In_2060);
and U407 (N_407,In_968,In_2258);
nor U408 (N_408,In_2730,In_552);
nor U409 (N_409,In_1530,In_1430);
xor U410 (N_410,In_1226,In_1770);
nor U411 (N_411,In_1759,In_2639);
nor U412 (N_412,In_1749,In_126);
and U413 (N_413,In_2123,In_2352);
xnor U414 (N_414,In_2319,In_47);
or U415 (N_415,In_1378,In_2089);
or U416 (N_416,In_1416,In_1625);
or U417 (N_417,In_793,In_2119);
or U418 (N_418,In_2775,In_1737);
nand U419 (N_419,In_2777,In_176);
and U420 (N_420,In_1006,In_2504);
xnor U421 (N_421,In_2533,In_426);
nand U422 (N_422,In_2955,In_2598);
or U423 (N_423,In_476,In_2966);
xnor U424 (N_424,In_2528,In_2147);
nor U425 (N_425,In_1248,In_615);
xor U426 (N_426,In_1083,In_2741);
nor U427 (N_427,In_1942,In_1570);
nor U428 (N_428,In_1835,In_2564);
or U429 (N_429,In_1,In_1640);
or U430 (N_430,In_350,In_1855);
xor U431 (N_431,In_526,In_1078);
or U432 (N_432,In_2887,In_1702);
and U433 (N_433,In_2007,In_1781);
xnor U434 (N_434,In_2602,In_1738);
nand U435 (N_435,In_976,In_54);
nor U436 (N_436,In_2312,In_2743);
xor U437 (N_437,In_2866,In_1010);
nor U438 (N_438,In_340,In_1608);
nand U439 (N_439,In_2711,In_2817);
xor U440 (N_440,In_2862,In_842);
or U441 (N_441,In_2785,In_867);
and U442 (N_442,In_1462,In_1685);
or U443 (N_443,In_23,In_2666);
or U444 (N_444,In_2864,In_2637);
xnor U445 (N_445,In_1653,In_2148);
or U446 (N_446,In_1463,In_724);
xor U447 (N_447,In_1745,In_725);
and U448 (N_448,In_1050,In_1313);
nand U449 (N_449,In_2626,In_2841);
nand U450 (N_450,In_2227,In_1708);
xnor U451 (N_451,In_2453,In_726);
or U452 (N_452,In_610,In_2357);
or U453 (N_453,In_2493,In_1121);
nor U454 (N_454,In_2596,In_1965);
or U455 (N_455,In_391,In_2751);
xnor U456 (N_456,In_1227,In_1677);
nor U457 (N_457,In_1228,In_1267);
nand U458 (N_458,In_1734,In_700);
or U459 (N_459,In_2261,In_1406);
nand U460 (N_460,In_1068,In_2481);
and U461 (N_461,In_517,In_2281);
or U462 (N_462,In_2902,In_31);
xnor U463 (N_463,In_156,In_1042);
nand U464 (N_464,In_1236,In_2460);
nor U465 (N_465,In_2589,In_2325);
nor U466 (N_466,In_2214,In_2506);
nand U467 (N_467,In_2077,In_1972);
nand U468 (N_468,In_1085,In_1051);
nand U469 (N_469,In_897,In_636);
or U470 (N_470,In_388,In_158);
nand U471 (N_471,In_2182,In_248);
nand U472 (N_472,In_2014,In_2165);
or U473 (N_473,In_529,In_744);
and U474 (N_474,In_1834,In_1477);
nor U475 (N_475,In_2154,In_2623);
nor U476 (N_476,In_184,In_1082);
xor U477 (N_477,In_1204,In_1840);
and U478 (N_478,In_111,In_2277);
nand U479 (N_479,In_107,In_1967);
and U480 (N_480,In_678,In_2221);
nand U481 (N_481,In_1259,In_133);
nor U482 (N_482,In_2482,In_2028);
xor U483 (N_483,In_410,In_2675);
and U484 (N_484,In_951,In_2968);
nand U485 (N_485,In_2239,In_2690);
xor U486 (N_486,In_812,In_693);
xnor U487 (N_487,In_1047,In_1364);
nand U488 (N_488,In_638,In_2220);
xnor U489 (N_489,In_1867,In_142);
or U490 (N_490,In_100,In_336);
xor U491 (N_491,In_635,In_306);
nor U492 (N_492,In_2606,In_1308);
xnor U493 (N_493,In_367,In_605);
and U494 (N_494,In_1433,In_2677);
nor U495 (N_495,In_2631,In_154);
and U496 (N_496,In_259,In_641);
nand U497 (N_497,In_1063,In_284);
or U498 (N_498,In_307,In_2142);
or U499 (N_499,In_1252,In_2549);
xnor U500 (N_500,In_2803,In_2516);
and U501 (N_501,In_1937,In_416);
or U502 (N_502,In_1412,In_1105);
nand U503 (N_503,In_701,In_2811);
nand U504 (N_504,In_2899,In_2629);
and U505 (N_505,In_1143,In_2011);
or U506 (N_506,In_1970,In_2719);
xor U507 (N_507,In_2945,In_2622);
nor U508 (N_508,In_2448,In_1181);
and U509 (N_509,In_884,In_2225);
xnor U510 (N_510,In_1344,In_86);
and U511 (N_511,In_2621,In_544);
or U512 (N_512,In_2658,In_2686);
xor U513 (N_513,In_1794,In_2439);
nand U514 (N_514,In_2053,In_1586);
and U515 (N_515,In_699,In_1877);
or U516 (N_516,In_1665,In_1329);
and U517 (N_517,In_2377,In_1548);
or U518 (N_518,In_883,In_1933);
xnor U519 (N_519,In_1448,In_2330);
nor U520 (N_520,In_1390,In_1144);
nor U521 (N_521,In_2423,In_1635);
nand U522 (N_522,In_1059,In_665);
nand U523 (N_523,In_551,In_1439);
xnor U524 (N_524,In_412,In_722);
xnor U525 (N_525,In_1762,In_1927);
and U526 (N_526,In_352,In_1200);
xnor U527 (N_527,In_110,In_2333);
xor U528 (N_528,In_1425,In_2520);
xor U529 (N_529,In_1971,In_570);
nand U530 (N_530,In_1633,In_574);
and U531 (N_531,In_2684,In_1041);
and U532 (N_532,In_752,In_1198);
xnor U533 (N_533,In_2605,In_2292);
and U534 (N_534,In_872,In_1693);
and U535 (N_535,In_433,In_1895);
nand U536 (N_536,In_2999,In_2927);
and U537 (N_537,In_2865,In_503);
nor U538 (N_538,In_486,In_1926);
nor U539 (N_539,In_187,In_2255);
and U540 (N_540,In_523,In_2003);
nor U541 (N_541,In_2537,In_1890);
and U542 (N_542,In_941,In_1712);
nand U543 (N_543,In_1661,In_1355);
xor U544 (N_544,In_440,In_2197);
or U545 (N_545,In_2660,In_2716);
or U546 (N_546,In_1517,In_2020);
xor U547 (N_547,In_322,In_973);
nand U548 (N_548,In_2654,In_1032);
and U549 (N_549,In_513,In_315);
xor U550 (N_550,In_1173,In_1292);
or U551 (N_551,In_790,In_1069);
or U552 (N_552,In_2206,In_2285);
nand U553 (N_553,In_1912,In_2403);
or U554 (N_554,In_1484,In_592);
and U555 (N_555,In_261,In_457);
or U556 (N_556,In_2656,In_2291);
nand U557 (N_557,In_2553,In_1998);
or U558 (N_558,In_2031,In_633);
and U559 (N_559,In_528,In_672);
nor U560 (N_560,In_1987,In_1444);
nand U561 (N_561,In_2818,In_347);
nand U562 (N_562,In_2174,In_2994);
and U563 (N_563,In_2974,In_436);
nand U564 (N_564,In_202,In_2689);
and U565 (N_565,In_1868,In_2244);
nand U566 (N_566,In_590,In_1309);
nor U567 (N_567,In_738,In_894);
nand U568 (N_568,In_2346,In_171);
xor U569 (N_569,In_2662,In_2139);
nand U570 (N_570,In_877,In_1480);
nand U571 (N_571,In_674,In_1824);
or U572 (N_572,In_671,In_2849);
xnor U573 (N_573,In_1117,In_943);
or U574 (N_574,In_1552,In_339);
or U575 (N_575,In_579,In_2799);
and U576 (N_576,In_478,In_1540);
or U577 (N_577,In_2828,In_534);
and U578 (N_578,In_2923,In_1569);
nor U579 (N_579,In_1305,In_1447);
nor U580 (N_580,In_1179,In_204);
and U581 (N_581,In_1149,In_2416);
xor U582 (N_582,In_2115,In_2947);
or U583 (N_583,In_468,In_853);
and U584 (N_584,In_1404,In_1764);
or U585 (N_585,In_1092,In_2066);
nor U586 (N_586,In_2435,In_83);
nor U587 (N_587,In_2160,In_1048);
and U588 (N_588,In_2572,In_2044);
nor U589 (N_589,In_2428,In_1402);
or U590 (N_590,In_1346,In_1407);
nand U591 (N_591,In_2410,In_1025);
and U592 (N_592,In_428,In_1664);
nor U593 (N_593,In_487,In_515);
or U594 (N_594,In_1733,In_28);
and U595 (N_595,In_1164,In_680);
or U596 (N_596,In_2942,In_2728);
xnor U597 (N_597,In_1265,In_1443);
xor U598 (N_598,In_2153,In_844);
nand U599 (N_599,In_2469,In_207);
or U600 (N_600,In_1249,In_1980);
and U601 (N_601,In_837,In_2216);
and U602 (N_602,In_1323,In_987);
nand U603 (N_603,In_422,In_2990);
nand U604 (N_604,In_2315,In_542);
xnor U605 (N_605,In_1802,In_286);
or U606 (N_606,In_1369,In_691);
nor U607 (N_607,In_459,In_1757);
nand U608 (N_608,In_266,In_1534);
or U609 (N_609,In_685,In_277);
nor U610 (N_610,In_2837,In_2253);
and U611 (N_611,In_787,In_2096);
or U612 (N_612,In_1555,In_995);
nand U613 (N_613,In_1075,In_2368);
and U614 (N_614,In_1225,In_597);
nor U615 (N_615,In_104,In_2424);
xnor U616 (N_616,In_2778,In_1030);
or U617 (N_617,In_1920,In_288);
xnor U618 (N_618,In_2731,In_76);
nand U619 (N_619,In_1944,In_944);
or U620 (N_620,In_2362,In_1157);
or U621 (N_621,In_1692,In_2091);
xnor U622 (N_622,In_2672,In_1525);
nand U623 (N_623,In_360,In_349);
nor U624 (N_624,In_40,In_2953);
nor U625 (N_625,In_2137,In_1741);
xor U626 (N_626,In_2722,In_1943);
nand U627 (N_627,In_1680,In_718);
xor U628 (N_628,In_324,In_78);
nand U629 (N_629,In_1605,In_762);
xor U630 (N_630,In_2714,In_1615);
nor U631 (N_631,In_2213,In_960);
nor U632 (N_632,In_1429,In_2565);
and U633 (N_633,In_182,In_24);
nand U634 (N_634,In_1518,In_643);
and U635 (N_635,In_303,In_1851);
nand U636 (N_636,In_612,In_2668);
and U637 (N_637,In_2118,In_304);
and U638 (N_638,In_1014,In_2511);
and U639 (N_639,In_902,In_692);
nor U640 (N_640,In_2363,In_520);
xnor U641 (N_641,In_1349,In_767);
or U642 (N_642,In_1312,In_1865);
nor U643 (N_643,In_1114,In_2320);
or U644 (N_644,In_4,In_1291);
or U645 (N_645,In_115,In_521);
xor U646 (N_646,In_53,In_661);
xnor U647 (N_647,In_1589,In_1054);
xor U648 (N_648,In_609,In_741);
nand U649 (N_649,In_608,In_1109);
and U650 (N_650,In_1843,In_2329);
and U651 (N_651,In_2347,In_1108);
or U652 (N_652,In_1336,In_557);
nand U653 (N_653,In_1456,In_2401);
or U654 (N_654,In_2749,In_373);
xnor U655 (N_655,In_1039,In_2861);
and U656 (N_656,In_1643,In_1765);
nand U657 (N_657,In_1096,In_43);
or U658 (N_658,In_1026,In_2217);
or U659 (N_659,In_2436,In_1061);
nand U660 (N_660,In_1656,In_2238);
and U661 (N_661,In_2855,In_1919);
nand U662 (N_662,In_601,In_386);
nor U663 (N_663,In_1381,In_1888);
nor U664 (N_664,In_229,In_1086);
or U665 (N_665,In_2872,In_312);
or U666 (N_666,In_688,In_2021);
and U667 (N_667,In_91,In_2814);
nand U668 (N_668,In_2124,In_210);
or U669 (N_669,In_939,In_2001);
and U670 (N_670,In_68,In_2748);
xnor U671 (N_671,In_1415,In_9);
xor U672 (N_672,In_92,In_1461);
or U673 (N_673,In_532,In_3);
nor U674 (N_674,In_1649,In_614);
and U675 (N_675,In_1148,In_1220);
xnor U676 (N_676,In_1127,In_1511);
or U677 (N_677,In_138,In_791);
nor U678 (N_678,In_2273,In_2783);
nand U679 (N_679,In_1994,In_1769);
or U680 (N_680,In_1452,In_1076);
and U681 (N_681,In_1908,In_1554);
xor U682 (N_682,In_1457,In_2911);
nor U683 (N_683,In_2391,In_2097);
and U684 (N_684,In_2759,In_1079);
or U685 (N_685,In_1602,In_165);
nand U686 (N_686,In_717,In_2485);
or U687 (N_687,In_502,In_2819);
and U688 (N_688,In_1306,In_538);
and U689 (N_689,In_2248,In_750);
or U690 (N_690,In_2032,In_20);
and U691 (N_691,In_1405,In_950);
xor U692 (N_692,In_1811,In_888);
and U693 (N_693,In_1389,In_771);
or U694 (N_694,In_1787,In_2420);
xor U695 (N_695,In_1574,In_96);
and U696 (N_696,In_364,In_2804);
xnor U697 (N_697,In_580,In_1887);
and U698 (N_698,In_1237,In_2199);
xnor U699 (N_699,In_2107,In_309);
or U700 (N_700,In_1674,In_177);
nor U701 (N_701,In_1436,In_2480);
or U702 (N_702,In_89,In_2792);
xor U703 (N_703,In_1445,In_1150);
nand U704 (N_704,In_2584,In_1502);
and U705 (N_705,In_1966,In_1212);
nand U706 (N_706,In_22,In_1245);
and U707 (N_707,In_2349,In_815);
xor U708 (N_708,In_2556,In_474);
nand U709 (N_709,In_423,In_2552);
or U710 (N_710,In_2692,In_1126);
nand U711 (N_711,In_2171,In_2141);
and U712 (N_712,In_893,In_703);
nor U713 (N_713,In_2432,In_2558);
xnor U714 (N_714,In_493,In_955);
xnor U715 (N_715,In_1377,In_62);
xor U716 (N_716,In_489,In_1760);
and U717 (N_717,In_683,In_1542);
nor U718 (N_718,In_1420,In_2335);
or U719 (N_719,In_660,In_109);
and U720 (N_720,In_2343,In_1597);
nor U721 (N_721,In_1029,In_2838);
nor U722 (N_722,In_1948,In_2375);
nor U723 (N_723,In_1367,In_1694);
and U724 (N_724,In_1706,In_1931);
nand U725 (N_725,In_2299,In_2527);
and U726 (N_726,In_2287,In_2200);
and U727 (N_727,In_1271,In_2706);
nand U728 (N_728,In_696,In_1875);
nor U729 (N_729,In_550,In_2224);
or U730 (N_730,In_2625,In_1136);
nand U731 (N_731,In_525,In_159);
nand U732 (N_732,In_2355,In_2);
and U733 (N_733,In_1652,In_2180);
nor U734 (N_734,In_1886,In_589);
nor U735 (N_735,In_739,In_1631);
or U736 (N_736,In_2696,In_2037);
xor U737 (N_737,In_1687,In_2863);
and U738 (N_738,In_1219,In_1088);
xor U739 (N_739,In_1453,In_1070);
nand U740 (N_740,In_127,In_1154);
nor U741 (N_741,In_1913,In_319);
xor U742 (N_742,In_408,In_1717);
nor U743 (N_743,In_1434,In_2308);
nor U744 (N_744,In_1052,In_2314);
xor U745 (N_745,In_2186,In_1203);
or U746 (N_746,In_1550,In_2272);
or U747 (N_747,In_2024,In_861);
nor U748 (N_748,In_1917,In_1603);
and U749 (N_749,In_1244,In_1595);
nand U750 (N_750,In_1872,In_2012);
nor U751 (N_751,In_1450,In_596);
xor U752 (N_752,In_2981,In_2390);
xnor U753 (N_753,In_1689,In_2973);
and U754 (N_754,In_1751,In_2769);
or U755 (N_755,In_2853,In_2566);
nor U756 (N_756,In_19,In_2191);
nor U757 (N_757,In_2472,In_123);
xnor U758 (N_758,In_2259,In_1379);
nor U759 (N_759,In_2643,In_1766);
or U760 (N_760,In_749,In_1115);
or U761 (N_761,In_1657,In_972);
xor U762 (N_762,In_1130,In_105);
and U763 (N_763,In_2762,In_764);
nor U764 (N_764,In_1883,In_2196);
nor U765 (N_765,In_1314,In_594);
xor U766 (N_766,In_1174,In_1516);
nand U767 (N_767,In_855,In_1932);
or U768 (N_768,In_2262,In_2063);
or U769 (N_769,In_834,In_1898);
or U770 (N_770,In_1936,In_2943);
or U771 (N_771,In_253,In_1822);
xnor U772 (N_772,In_1606,In_2715);
and U773 (N_773,In_1487,In_484);
nand U774 (N_774,In_136,In_2135);
nand U775 (N_775,In_2932,In_1356);
and U776 (N_776,In_1064,In_549);
or U777 (N_777,In_2205,In_668);
or U778 (N_778,In_648,In_395);
or U779 (N_779,In_376,In_1319);
and U780 (N_780,In_2132,In_223);
or U781 (N_781,In_251,In_889);
nand U782 (N_782,In_2062,In_2590);
nand U783 (N_783,In_1260,In_843);
nand U784 (N_784,In_1910,In_369);
nand U785 (N_785,In_1801,In_2274);
nand U786 (N_786,In_103,In_2458);
xor U787 (N_787,In_2181,In_1311);
and U788 (N_788,In_1934,In_1859);
xor U789 (N_789,In_629,In_2848);
nor U790 (N_790,In_1482,In_731);
and U791 (N_791,In_2970,In_1838);
nor U792 (N_792,In_602,In_2270);
and U793 (N_793,In_1683,In_1629);
or U794 (N_794,In_287,In_2721);
or U795 (N_795,In_761,In_2210);
and U796 (N_796,In_1818,In_343);
nand U797 (N_797,In_420,In_2640);
nor U798 (N_798,In_37,In_1719);
nand U799 (N_799,In_2635,In_329);
nand U800 (N_800,In_2242,In_2311);
nor U801 (N_801,In_235,In_1541);
or U802 (N_802,In_1208,In_382);
xor U803 (N_803,In_2407,In_2462);
and U804 (N_804,In_2760,In_2318);
xnor U805 (N_805,In_470,In_1303);
nand U806 (N_806,In_1722,In_1882);
nor U807 (N_807,In_1543,In_2657);
nand U808 (N_808,In_469,In_2002);
or U809 (N_809,In_1008,In_18);
xnor U810 (N_810,In_1923,In_2857);
xor U811 (N_811,In_1696,In_2867);
nor U812 (N_812,In_940,In_1565);
nand U813 (N_813,In_1384,In_356);
nand U814 (N_814,In_354,In_2972);
xnor U815 (N_815,In_963,In_854);
xor U816 (N_816,In_1634,In_281);
xnor U817 (N_817,In_2998,In_1983);
xnor U818 (N_818,In_2486,In_2718);
and U819 (N_819,In_1186,In_1021);
nand U820 (N_820,In_2350,In_2790);
or U821 (N_821,In_2425,In_443);
xor U822 (N_822,In_1031,In_1870);
nand U823 (N_823,In_1112,In_712);
or U824 (N_824,In_2568,In_981);
nor U825 (N_825,In_1388,In_2125);
or U826 (N_826,In_2593,In_1383);
and U827 (N_827,In_348,In_578);
or U828 (N_828,In_801,In_906);
nand U829 (N_829,In_1559,In_2750);
nand U830 (N_830,In_581,In_2601);
xnor U831 (N_831,In_2978,In_427);
or U832 (N_832,In_2402,In_723);
xor U833 (N_833,In_619,In_1122);
nand U834 (N_834,In_1527,In_1714);
or U835 (N_835,In_1791,In_2383);
xor U836 (N_836,In_2627,In_1431);
nor U837 (N_837,In_1949,In_1411);
xnor U838 (N_838,In_1073,In_1782);
nand U839 (N_839,In_337,In_2524);
xor U840 (N_840,In_2376,In_2500);
xor U841 (N_841,In_2787,In_2946);
xnor U842 (N_842,In_558,In_1128);
xor U843 (N_843,In_2515,In_1118);
nor U844 (N_844,In_1327,In_2586);
and U845 (N_845,In_1853,In_2295);
nand U846 (N_846,In_2078,In_1449);
or U847 (N_847,In_2339,In_2928);
nor U848 (N_848,In_2840,In_1500);
and U849 (N_849,In_1473,In_1043);
and U850 (N_850,In_2265,In_1992);
xnor U851 (N_851,In_1907,In_631);
xnor U852 (N_852,In_2301,In_2906);
nand U853 (N_853,In_1414,In_1991);
nand U854 (N_854,In_781,In_168);
nor U855 (N_855,In_2172,In_2641);
or U856 (N_856,In_234,In_1235);
nand U857 (N_857,In_2897,In_1398);
or U858 (N_858,In_1318,In_252);
and U859 (N_859,In_196,In_2254);
nand U860 (N_860,In_2336,In_2499);
or U861 (N_861,In_989,In_1854);
nor U862 (N_862,In_1553,In_2977);
nand U863 (N_863,In_2166,In_1270);
or U864 (N_864,In_1632,In_1077);
nor U865 (N_865,In_1103,In_591);
xnor U866 (N_866,In_2509,In_1561);
nor U867 (N_867,In_1328,In_742);
and U868 (N_868,In_2419,In_1337);
nand U869 (N_869,In_1139,In_1156);
xor U870 (N_870,In_985,In_198);
nand U871 (N_871,In_958,In_1728);
xnor U872 (N_872,In_2884,In_2047);
or U873 (N_873,In_1842,In_2373);
xor U874 (N_874,In_13,In_876);
nand U875 (N_875,In_1460,In_2904);
nand U876 (N_876,In_2518,In_1748);
xnor U877 (N_877,In_1788,In_1466);
and U878 (N_878,In_1189,In_607);
nor U879 (N_879,In_1177,In_2317);
nand U880 (N_880,In_2075,In_435);
xor U881 (N_881,In_1284,In_403);
nor U882 (N_882,In_548,In_1421);
nor U883 (N_883,In_1753,In_51);
and U884 (N_884,In_297,In_1956);
nor U885 (N_885,In_276,In_2211);
nor U886 (N_886,In_2710,In_2740);
xor U887 (N_887,In_755,In_2642);
or U888 (N_888,In_1345,In_1796);
nand U889 (N_889,In_709,In_813);
and U890 (N_890,In_2309,In_559);
and U891 (N_891,In_2208,In_2952);
and U892 (N_892,In_2008,In_1900);
and U893 (N_893,In_999,In_977);
nand U894 (N_894,In_2554,In_1874);
and U895 (N_895,In_108,In_2763);
nand U896 (N_896,In_1731,In_1387);
nand U897 (N_897,In_190,In_1889);
or U898 (N_898,In_2156,In_2525);
nor U899 (N_899,In_992,In_2378);
or U900 (N_900,In_2452,In_2667);
or U901 (N_901,In_2526,In_2465);
nor U902 (N_902,In_863,In_1217);
nand U903 (N_903,In_80,In_1662);
xor U904 (N_904,In_1418,In_2069);
xor U905 (N_905,In_971,In_2869);
nand U906 (N_906,In_710,In_8);
nor U907 (N_907,In_1321,In_1503);
or U908 (N_908,In_275,In_2592);
xor U909 (N_909,In_305,In_835);
xnor U910 (N_910,In_795,In_257);
nand U911 (N_911,In_2967,In_796);
xnor U912 (N_912,In_1424,In_1376);
nor U913 (N_913,In_2275,In_620);
and U914 (N_914,In_172,In_1672);
or U915 (N_915,In_475,In_2204);
or U916 (N_916,In_2231,In_646);
and U917 (N_917,In_2140,In_1638);
and U918 (N_918,In_969,In_194);
and U919 (N_919,In_1067,In_2235);
nand U920 (N_920,In_1780,In_2367);
nand U921 (N_921,In_2246,In_27);
nor U922 (N_922,In_898,In_698);
xor U923 (N_923,In_2951,In_2271);
or U924 (N_924,In_2827,In_915);
or U925 (N_925,In_134,In_2437);
xor U926 (N_926,In_2852,In_1945);
nor U927 (N_927,In_2198,In_2854);
xnor U928 (N_928,In_780,In_1628);
or U929 (N_929,In_2267,In_745);
nand U930 (N_930,In_1535,In_1131);
nor U931 (N_931,In_922,In_1056);
or U932 (N_932,In_2997,In_2297);
xnor U933 (N_933,In_341,In_2081);
xnor U934 (N_934,In_818,In_70);
and U935 (N_935,In_488,In_1941);
or U936 (N_936,In_507,In_1116);
and U937 (N_937,In_225,In_1155);
and U938 (N_938,In_2035,In_2559);
and U939 (N_939,In_564,In_914);
nor U940 (N_940,In_1060,In_2608);
xor U941 (N_941,In_794,In_1521);
or U942 (N_942,In_2263,In_2045);
nand U943 (N_943,In_527,In_2624);
nand U944 (N_944,In_2707,In_1648);
xor U945 (N_945,In_663,In_166);
nand U946 (N_946,In_2701,In_798);
and U947 (N_947,In_2103,In_439);
or U948 (N_948,In_335,In_1575);
nand U949 (N_949,In_1954,In_14);
or U950 (N_950,In_1307,In_1596);
nor U951 (N_951,In_327,In_1876);
or U952 (N_952,In_361,In_1763);
and U953 (N_953,In_1808,In_460);
nand U954 (N_954,In_1080,In_1184);
or U955 (N_955,In_2179,In_1257);
nor U956 (N_956,In_572,In_1676);
or U957 (N_957,In_1197,In_2155);
or U958 (N_958,In_965,In_208);
or U959 (N_959,In_1582,In_291);
xor U960 (N_960,In_729,In_17);
nor U961 (N_961,In_836,In_2369);
xor U962 (N_962,In_2700,In_708);
or U963 (N_963,In_1036,In_571);
xor U964 (N_964,In_1580,In_1486);
xnor U965 (N_965,In_625,In_2796);
or U966 (N_966,In_1350,In_451);
and U967 (N_967,In_230,In_66);
nand U968 (N_968,In_383,In_50);
nor U969 (N_969,In_318,In_1172);
xor U970 (N_970,In_6,In_2871);
and U971 (N_971,In_1380,In_850);
nand U972 (N_972,In_2389,In_2360);
xor U973 (N_973,In_1218,In_1523);
nor U974 (N_974,In_477,In_1650);
and U975 (N_975,In_595,In_1507);
xor U976 (N_976,In_1261,In_1210);
nor U977 (N_977,In_1930,In_617);
xor U978 (N_978,In_1715,In_290);
nor U979 (N_979,In_1506,In_463);
and U980 (N_980,In_1316,In_2443);
nor U981 (N_981,In_2673,In_1015);
and U982 (N_982,In_2798,In_21);
xnor U983 (N_983,In_2023,In_907);
or U984 (N_984,In_219,In_1209);
nor U985 (N_985,In_155,In_1264);
nor U986 (N_986,In_1735,In_1778);
and U987 (N_987,In_2727,In_2192);
and U988 (N_988,In_2475,In_2394);
xor U989 (N_989,In_1458,In_569);
and U990 (N_990,In_16,In_2523);
nand U991 (N_991,In_338,In_264);
nor U992 (N_992,In_2503,In_681);
nor U993 (N_993,In_2157,In_2539);
xnor U994 (N_994,In_2222,In_289);
nor U995 (N_995,In_1996,In_1566);
nand U996 (N_996,In_1726,In_2664);
xor U997 (N_997,In_1846,In_472);
xnor U998 (N_998,In_1551,In_860);
nand U999 (N_999,In_1170,In_2145);
or U1000 (N_1000,In_150,In_543);
xor U1001 (N_1001,In_2404,In_2234);
nand U1002 (N_1002,In_125,In_2860);
nand U1003 (N_1003,In_1001,In_1707);
nor U1004 (N_1004,In_65,In_2744);
or U1005 (N_1005,In_1110,In_2305);
and U1006 (N_1006,In_2674,In_829);
nand U1007 (N_1007,In_2685,In_2644);
or U1008 (N_1008,In_432,In_2194);
nor U1009 (N_1009,In_1775,In_2371);
or U1010 (N_1010,In_1845,In_2788);
or U1011 (N_1011,In_212,In_1817);
nand U1012 (N_1012,In_1744,In_2649);
xor U1013 (N_1013,In_1065,In_743);
nand U1014 (N_1014,In_2588,In_2612);
nand U1015 (N_1015,In_2620,In_2679);
xnor U1016 (N_1016,In_2980,In_2647);
or U1017 (N_1017,In_859,In_1623);
or U1018 (N_1018,In_1732,In_372);
nand U1019 (N_1019,In_262,In_2779);
or U1020 (N_1020,In_2908,In_355);
or U1021 (N_1021,In_1413,In_1467);
and U1022 (N_1022,In_1385,In_1578);
xnor U1023 (N_1023,In_2382,In_1401);
or U1024 (N_1024,In_838,In_2653);
and U1025 (N_1025,In_1592,In_1009);
nand U1026 (N_1026,In_2033,In_934);
and U1027 (N_1027,In_2850,In_311);
or U1028 (N_1028,In_401,In_1669);
nand U1029 (N_1029,In_1666,In_2680);
and U1030 (N_1030,In_2594,In_2161);
or U1031 (N_1031,In_2005,In_841);
nand U1032 (N_1032,In_896,In_778);
nor U1033 (N_1033,In_254,In_32);
nand U1034 (N_1034,In_650,In_948);
nand U1035 (N_1035,In_1240,In_613);
and U1036 (N_1036,In_1946,In_2878);
nand U1037 (N_1037,In_197,In_145);
or U1038 (N_1038,In_858,In_2374);
and U1039 (N_1039,In_1013,In_1847);
xnor U1040 (N_1040,In_1494,In_2218);
xnor U1041 (N_1041,In_1375,In_2845);
nor U1042 (N_1042,In_2522,In_1111);
or U1043 (N_1043,In_2138,In_2445);
or U1044 (N_1044,In_2487,In_1191);
or U1045 (N_1045,In_2384,In_1133);
xor U1046 (N_1046,In_2468,In_603);
or U1047 (N_1047,In_1803,In_654);
and U1048 (N_1048,In_2237,In_1976);
and U1049 (N_1049,In_217,In_840);
nor U1050 (N_1050,In_2236,In_2916);
or U1051 (N_1051,In_2875,In_1038);
nor U1052 (N_1052,In_1394,In_1583);
xor U1053 (N_1053,In_598,In_2215);
nand U1054 (N_1054,In_2807,In_1074);
and U1055 (N_1055,In_2185,In_804);
nand U1056 (N_1056,In_2802,In_662);
xor U1057 (N_1057,In_1496,In_568);
nand U1058 (N_1058,In_2833,In_2086);
and U1059 (N_1059,In_1018,In_1242);
xnor U1060 (N_1060,In_706,In_1066);
xor U1061 (N_1061,In_1626,In_2440);
xnor U1062 (N_1062,In_268,In_448);
xnor U1063 (N_1063,In_1604,In_2427);
nor U1064 (N_1064,In_362,In_2698);
or U1065 (N_1065,In_2489,In_2984);
or U1066 (N_1066,In_247,In_2454);
and U1067 (N_1067,In_2915,In_122);
xor U1068 (N_1068,In_2929,In_2476);
or U1069 (N_1069,In_270,In_1723);
xnor U1070 (N_1070,In_621,In_1831);
nor U1071 (N_1071,In_1903,In_1819);
and U1072 (N_1072,In_1825,In_2397);
and U1073 (N_1073,In_2307,In_2655);
xor U1074 (N_1074,In_2632,In_224);
and U1075 (N_1075,In_1247,In_1358);
and U1076 (N_1076,In_1612,In_2563);
xnor U1077 (N_1077,In_1593,In_2426);
xor U1078 (N_1078,In_461,In_1185);
or U1079 (N_1079,In_1617,In_378);
or U1080 (N_1080,In_1740,In_243);
nand U1081 (N_1081,In_2991,In_1671);
and U1082 (N_1082,In_811,In_239);
and U1083 (N_1083,In_505,In_381);
xnor U1084 (N_1084,In_2084,In_188);
or U1085 (N_1085,In_1468,In_1784);
xor U1086 (N_1086,In_1975,In_2022);
xor U1087 (N_1087,In_358,In_1045);
or U1088 (N_1088,In_211,In_832);
and U1089 (N_1089,In_624,In_2473);
and U1090 (N_1090,In_2971,In_705);
nand U1091 (N_1091,In_2446,In_218);
nor U1092 (N_1092,In_385,In_2851);
nand U1093 (N_1093,In_1167,In_101);
or U1094 (N_1094,In_1588,In_2004);
nand U1095 (N_1095,In_200,In_886);
and U1096 (N_1096,In_2585,In_673);
xor U1097 (N_1097,In_2051,In_604);
nor U1098 (N_1098,In_2521,In_758);
xor U1099 (N_1099,In_1471,In_2111);
xnor U1100 (N_1100,In_874,In_2013);
nor U1101 (N_1101,In_820,In_498);
or U1102 (N_1102,In_2912,In_1577);
nor U1103 (N_1103,In_1614,In_2015);
xnor U1104 (N_1104,In_1864,In_2962);
nor U1105 (N_1105,In_1929,In_1176);
and U1106 (N_1106,In_2245,In_1465);
or U1107 (N_1107,In_1400,In_2417);
and U1108 (N_1108,In_1275,In_2300);
nor U1109 (N_1109,In_2650,In_518);
xor U1110 (N_1110,In_720,In_546);
nand U1111 (N_1111,In_1269,In_2286);
xnor U1112 (N_1112,In_2190,In_2931);
and U1113 (N_1113,In_970,In_2269);
or U1114 (N_1114,In_2010,In_1221);
xnor U1115 (N_1115,In_2836,In_1939);
or U1116 (N_1116,In_438,In_556);
and U1117 (N_1117,In_2284,In_55);
nand U1118 (N_1118,In_2630,In_2555);
nor U1119 (N_1119,In_2364,In_1002);
or U1120 (N_1120,In_618,In_1797);
nand U1121 (N_1121,In_623,In_95);
or U1122 (N_1122,In_1529,In_616);
nand U1123 (N_1123,In_2016,In_991);
and U1124 (N_1124,In_1317,In_52);
or U1125 (N_1125,In_707,In_2988);
or U1126 (N_1126,In_15,In_2891);
and U1127 (N_1127,In_84,In_1241);
nor U1128 (N_1128,In_114,In_1544);
or U1129 (N_1129,In_2939,In_645);
and U1130 (N_1130,In_495,In_2538);
or U1131 (N_1131,In_2580,In_2918);
and U1132 (N_1132,In_417,In_931);
nor U1133 (N_1133,In_2669,In_2043);
or U1134 (N_1134,In_147,In_1287);
and U1135 (N_1135,In_2770,In_2917);
or U1136 (N_1136,In_48,In_308);
nand U1137 (N_1137,In_2102,In_856);
or U1138 (N_1138,In_676,In_1123);
xnor U1139 (N_1139,In_2920,In_1647);
or U1140 (N_1140,In_320,In_2793);
or U1141 (N_1141,In_377,In_2461);
or U1142 (N_1142,In_1151,In_242);
xor U1143 (N_1143,In_784,In_1710);
and U1144 (N_1144,In_2332,In_2113);
and U1145 (N_1145,In_504,In_2109);
nor U1146 (N_1146,In_599,In_1771);
nand U1147 (N_1147,In_1558,In_2882);
nor U1148 (N_1148,In_2781,In_444);
nor U1149 (N_1149,In_185,In_2074);
xor U1150 (N_1150,In_98,In_2877);
and U1151 (N_1151,In_1135,In_2604);
nand U1152 (N_1152,In_735,In_639);
nor U1153 (N_1153,In_342,In_1906);
nand U1154 (N_1154,In_1479,In_1335);
nor U1155 (N_1155,In_1137,In_1214);
nand U1156 (N_1156,In_541,In_1901);
xor U1157 (N_1157,In_783,In_2082);
or U1158 (N_1158,In_2006,In_2430);
and U1159 (N_1159,In_2597,In_947);
nand U1160 (N_1160,In_465,In_1091);
xor U1161 (N_1161,In_1767,In_35);
or U1162 (N_1162,In_2756,In_2542);
and U1163 (N_1163,In_1961,In_810);
nand U1164 (N_1164,In_233,In_139);
and U1165 (N_1165,In_2116,In_1071);
or U1166 (N_1166,In_2963,In_913);
nor U1167 (N_1167,In_2591,In_1446);
xor U1168 (N_1168,In_220,In_2847);
nand U1169 (N_1169,In_26,In_330);
xor U1170 (N_1170,In_1644,In_878);
nand U1171 (N_1171,In_1730,In_727);
nor U1172 (N_1172,In_2054,In_1020);
and U1173 (N_1173,In_1958,In_379);
or U1174 (N_1174,In_1813,In_295);
xor U1175 (N_1175,In_1231,In_2092);
and U1176 (N_1176,In_1253,In_852);
or U1177 (N_1177,In_1024,In_540);
or U1178 (N_1178,In_2169,In_983);
xor U1179 (N_1179,In_368,In_509);
nand U1180 (N_1180,In_1546,In_2143);
xor U1181 (N_1181,In_954,In_1713);
and U1182 (N_1182,In_857,In_519);
and U1183 (N_1183,In_1963,In_2264);
nor U1184 (N_1184,In_162,In_1366);
nand U1185 (N_1185,In_573,In_2767);
xor U1186 (N_1186,In_1675,In_2579);
nand U1187 (N_1187,In_1146,In_514);
nor U1188 (N_1188,In_1869,In_1815);
nor U1189 (N_1189,In_2789,In_405);
xnor U1190 (N_1190,In_918,In_75);
nand U1191 (N_1191,In_2058,In_2470);
and U1192 (N_1192,In_2388,In_715);
xor U1193 (N_1193,In_1522,In_313);
xor U1194 (N_1194,In_1836,In_1609);
nor U1195 (N_1195,In_1858,In_1296);
nand U1196 (N_1196,In_566,In_2250);
or U1197 (N_1197,In_2276,In_2600);
nor U1198 (N_1198,In_1300,In_990);
and U1199 (N_1199,In_2571,In_839);
or U1200 (N_1200,In_2158,In_57);
or U1201 (N_1201,In_1491,In_2548);
or U1202 (N_1202,In_394,In_2582);
and U1203 (N_1203,In_94,In_2776);
or U1204 (N_1204,In_728,In_588);
xnor U1205 (N_1205,In_2385,In_1879);
nor U1206 (N_1206,In_848,In_480);
xor U1207 (N_1207,In_2671,In_670);
nand U1208 (N_1208,In_256,In_2983);
and U1209 (N_1209,In_1746,In_272);
and U1210 (N_1210,In_1524,In_1627);
or U1211 (N_1211,In_1756,In_2306);
nand U1212 (N_1212,In_2094,In_1263);
nor U1213 (N_1213,In_1153,In_2843);
or U1214 (N_1214,In_1081,In_1288);
and U1215 (N_1215,In_1953,In_2351);
and U1216 (N_1216,In_675,In_1089);
nand U1217 (N_1217,In_2502,In_2941);
nor U1218 (N_1218,In_1839,In_1739);
and U1219 (N_1219,In_2683,In_2844);
nor U1220 (N_1220,In_2193,In_2913);
xor U1221 (N_1221,In_1033,In_406);
and U1222 (N_1222,In_2992,In_178);
or U1223 (N_1223,In_384,In_814);
or U1224 (N_1224,In_2212,In_2583);
xnor U1225 (N_1225,In_833,In_2087);
nand U1226 (N_1226,In_169,In_2252);
xnor U1227 (N_1227,In_1585,In_1531);
and U1228 (N_1228,In_1826,In_2429);
and U1229 (N_1229,In_271,In_45);
nor U1230 (N_1230,In_2773,In_2444);
and U1231 (N_1231,In_1348,In_456);
xor U1232 (N_1232,In_1332,In_2099);
and U1233 (N_1233,In_1964,In_1810);
and U1234 (N_1234,In_817,In_1899);
nand U1235 (N_1235,In_2150,In_679);
and U1236 (N_1236,In_1688,In_1695);
xnor U1237 (N_1237,In_1783,In_998);
xor U1238 (N_1238,In_2093,In_1438);
nand U1239 (N_1239,In_2278,In_1351);
and U1240 (N_1240,In_1914,In_1547);
or U1241 (N_1241,In_1878,In_1062);
nor U1242 (N_1242,In_392,In_441);
or U1243 (N_1243,In_1673,In_2293);
and U1244 (N_1244,In_2341,In_2243);
nor U1245 (N_1245,In_2163,In_186);
and U1246 (N_1246,In_2090,In_2989);
or U1247 (N_1247,In_2110,In_2497);
nand U1248 (N_1248,In_962,In_1718);
xor U1249 (N_1249,In_1892,In_545);
or U1250 (N_1250,In_2747,In_1736);
xnor U1251 (N_1251,In_1499,In_1997);
or U1252 (N_1252,In_149,In_2149);
nand U1253 (N_1253,In_146,In_657);
xor U1254 (N_1254,In_2921,In_2691);
and U1255 (N_1255,In_2442,In_128);
and U1256 (N_1256,In_2055,In_33);
and U1257 (N_1257,In_56,In_424);
xor U1258 (N_1258,In_2795,In_1922);
nor U1259 (N_1259,In_2303,In_1703);
or U1260 (N_1260,In_2510,In_455);
or U1261 (N_1261,In_1761,In_1510);
nor U1262 (N_1262,In_879,In_1978);
nor U1263 (N_1263,In_482,In_1747);
nand U1264 (N_1264,In_1938,In_2034);
or U1265 (N_1265,In_2546,In_2233);
and U1266 (N_1266,In_2176,In_586);
xnor U1267 (N_1267,In_1199,In_2910);
xnor U1268 (N_1268,In_1645,In_1911);
xnor U1269 (N_1269,In_2687,In_961);
xor U1270 (N_1270,In_777,In_1613);
xor U1271 (N_1271,In_5,In_1124);
xnor U1272 (N_1272,In_41,In_407);
nand U1273 (N_1273,In_910,In_102);
and U1274 (N_1274,In_429,In_2739);
xor U1275 (N_1275,In_945,In_2893);
xnor U1276 (N_1276,In_1058,In_2681);
and U1277 (N_1277,In_1125,In_293);
xnor U1278 (N_1278,In_446,In_751);
nand U1279 (N_1279,In_1678,In_1904);
or U1280 (N_1280,In_819,In_845);
xor U1281 (N_1281,In_1891,In_785);
nand U1282 (N_1282,In_2645,In_647);
or U1283 (N_1283,In_316,In_167);
nand U1284 (N_1284,In_88,In_979);
nand U1285 (N_1285,In_2498,In_1182);
xor U1286 (N_1286,In_1223,In_1984);
xnor U1287 (N_1287,In_1584,In_351);
nand U1288 (N_1288,In_164,In_2400);
xor U1289 (N_1289,In_345,In_2466);
nor U1290 (N_1290,In_1320,In_387);
nand U1291 (N_1291,In_2059,In_655);
or U1292 (N_1292,In_2832,In_2422);
xor U1293 (N_1293,In_1325,In_67);
nand U1294 (N_1294,In_2575,In_1343);
and U1295 (N_1295,In_390,In_754);
xnor U1296 (N_1296,In_1654,In_181);
and U1297 (N_1297,In_2080,In_2296);
and U1298 (N_1298,In_442,In_2396);
nor U1299 (N_1299,In_2907,In_2646);
xnor U1300 (N_1300,In_173,In_400);
or U1301 (N_1301,In_563,In_2599);
nand U1302 (N_1302,In_157,In_2313);
nand U1303 (N_1303,In_1668,In_2088);
or U1304 (N_1304,In_2834,In_808);
nor U1305 (N_1305,In_644,In_2071);
and U1306 (N_1306,In_2734,In_2095);
nor U1307 (N_1307,In_759,In_2607);
nor U1308 (N_1308,In_1207,In_195);
xnor U1309 (N_1309,In_747,In_2450);
nor U1310 (N_1310,In_1372,In_132);
or U1311 (N_1311,In_2949,In_2167);
nor U1312 (N_1312,In_1857,In_1639);
nor U1313 (N_1313,In_690,In_1037);
and U1314 (N_1314,In_1171,In_10);
xnor U1315 (N_1315,In_2995,In_539);
and U1316 (N_1316,In_2056,In_2406);
xor U1317 (N_1317,In_553,In_560);
or U1318 (N_1318,In_510,In_458);
or U1319 (N_1319,In_935,In_265);
nand U1320 (N_1320,In_1391,In_2835);
and U1321 (N_1321,In_584,In_2883);
or U1322 (N_1322,In_2665,In_46);
xnor U1323 (N_1323,In_191,In_1361);
and U1324 (N_1324,In_1141,In_375);
xor U1325 (N_1325,In_1990,In_2780);
xnor U1326 (N_1326,In_2638,In_237);
or U1327 (N_1327,In_1545,In_491);
xnor U1328 (N_1328,In_851,In_2418);
nor U1329 (N_1329,In_2957,In_2938);
nand U1330 (N_1330,In_1093,In_1134);
or U1331 (N_1331,In_1501,In_2327);
and U1332 (N_1332,In_34,In_1334);
and U1333 (N_1333,In_302,In_90);
nor U1334 (N_1334,In_310,In_2725);
or U1335 (N_1335,In_920,In_2144);
nand U1336 (N_1336,In_2735,In_131);
or U1337 (N_1337,In_58,In_1408);
nand U1338 (N_1338,In_2183,In_1799);
and U1339 (N_1339,In_1828,In_393);
nor U1340 (N_1340,In_760,In_1490);
and U1341 (N_1341,In_1885,In_2164);
xor U1342 (N_1342,In_2289,In_1873);
nand U1343 (N_1343,In_1277,In_949);
or U1344 (N_1344,In_1392,In_2713);
or U1345 (N_1345,In_183,In_1841);
nand U1346 (N_1346,In_1251,In_1000);
xor U1347 (N_1347,In_1049,In_2260);
and U1348 (N_1348,In_1451,In_1454);
and U1349 (N_1349,In_2241,In_1594);
nand U1350 (N_1350,In_1619,In_500);
and U1351 (N_1351,In_2353,In_1918);
nand U1352 (N_1352,In_2512,In_2131);
or U1353 (N_1353,In_512,In_1246);
nor U1354 (N_1354,In_1129,In_118);
xor U1355 (N_1355,In_800,In_932);
and U1356 (N_1356,In_1055,In_716);
and U1357 (N_1357,In_11,In_1469);
nand U1358 (N_1358,In_2451,In_2490);
nor U1359 (N_1359,In_2108,In_1616);
nor U1360 (N_1360,In_1955,In_2508);
nor U1361 (N_1361,In_2392,In_2477);
or U1362 (N_1362,In_953,In_2704);
xnor U1363 (N_1363,In_2249,In_1641);
and U1364 (N_1364,In_1280,In_485);
and U1365 (N_1365,In_772,In_2925);
and U1366 (N_1366,In_2030,In_677);
nand U1367 (N_1367,In_1354,In_2134);
nand U1368 (N_1368,In_1046,In_2189);
nand U1369 (N_1369,In_402,In_2764);
nor U1370 (N_1370,In_1166,In_371);
nor U1371 (N_1371,In_2079,In_1952);
nand U1372 (N_1372,In_2636,In_664);
nor U1373 (N_1373,In_2017,In_2926);
nor U1374 (N_1374,In_880,In_501);
nand U1375 (N_1375,In_2982,In_1016);
xnor U1376 (N_1376,In_1239,In_12);
or U1377 (N_1377,In_2562,In_1658);
and U1378 (N_1378,In_577,In_397);
or U1379 (N_1379,In_1493,In_2975);
nand U1380 (N_1380,In_1721,In_1704);
nor U1381 (N_1381,In_77,In_2603);
xnor U1382 (N_1382,In_2413,In_1011);
or U1383 (N_1383,In_1528,In_1256);
and U1384 (N_1384,In_1159,In_2128);
or U1385 (N_1385,In_479,In_2808);
xor U1386 (N_1386,In_363,In_2052);
nor U1387 (N_1387,In_1536,In_2663);
and U1388 (N_1388,In_292,In_1758);
nand U1389 (N_1389,In_1959,In_1395);
and U1390 (N_1390,In_1848,In_1266);
nand U1391 (N_1391,In_1003,In_522);
nand U1392 (N_1392,In_774,In_1750);
nor U1393 (N_1393,In_1697,In_516);
nor U1394 (N_1394,In_1339,In_1621);
or U1395 (N_1395,In_241,In_567);
or U1396 (N_1396,In_1175,In_2279);
and U1397 (N_1397,In_2162,In_1768);
xnor U1398 (N_1398,In_2774,In_2304);
xor U1399 (N_1399,In_2501,In_911);
or U1400 (N_1400,In_2257,In_357);
xor U1401 (N_1401,In_1651,In_398);
or U1402 (N_1402,In_2449,In_711);
nand U1403 (N_1403,In_2801,In_1234);
xor U1404 (N_1404,In_1106,In_365);
nor U1405 (N_1405,In_2766,In_2159);
xor U1406 (N_1406,In_511,In_2415);
nor U1407 (N_1407,In_1441,In_2195);
xor U1408 (N_1408,In_359,In_2996);
and U1409 (N_1409,In_1102,In_1193);
nand U1410 (N_1410,In_938,In_1705);
nor U1411 (N_1411,In_2771,In_2754);
xnor U1412 (N_1412,In_1622,In_702);
xor U1413 (N_1413,In_2753,In_593);
or U1414 (N_1414,In_825,In_2366);
nor U1415 (N_1415,In_209,In_419);
and U1416 (N_1416,In_2251,In_2076);
or U1417 (N_1417,In_2412,In_1679);
nand U1418 (N_1418,In_656,In_823);
nor U1419 (N_1419,In_649,In_2752);
and U1420 (N_1420,In_1464,In_2757);
xnor U1421 (N_1421,In_2765,In_1293);
nand U1422 (N_1422,In_885,In_1655);
xnor U1423 (N_1423,In_163,In_1374);
or U1424 (N_1424,In_1526,In_490);
nor U1425 (N_1425,In_2831,In_1549);
or U1426 (N_1426,In_2529,In_471);
nand U1427 (N_1427,In_2879,In_2561);
xor U1428 (N_1428,In_2534,In_642);
or U1429 (N_1429,In_909,In_2085);
or U1430 (N_1430,In_71,In_640);
or U1431 (N_1431,In_978,In_1852);
nor U1432 (N_1432,In_1216,In_1233);
nor U1433 (N_1433,In_993,In_450);
nand U1434 (N_1434,In_258,In_1729);
xnor U1435 (N_1435,In_283,In_1330);
or U1436 (N_1436,In_1716,In_925);
and U1437 (N_1437,In_2723,In_2944);
or U1438 (N_1438,In_1902,In_414);
nor U1439 (N_1439,In_2209,In_769);
xnor U1440 (N_1440,In_2431,In_1478);
xor U1441 (N_1441,In_328,In_59);
nand U1442 (N_1442,In_1897,In_1472);
or U1443 (N_1443,In_988,In_1347);
and U1444 (N_1444,In_766,In_0);
nand U1445 (N_1445,In_2821,In_2797);
and U1446 (N_1446,In_2922,In_1598);
nor U1447 (N_1447,In_576,In_1999);
and U1448 (N_1448,In_2709,In_2105);
nor U1449 (N_1449,In_2856,In_1474);
and U1450 (N_1450,In_2829,In_42);
xor U1451 (N_1451,In_2370,In_2479);
nor U1452 (N_1452,In_282,In_2117);
nor U1453 (N_1453,In_919,In_1798);
nand U1454 (N_1454,In_803,In_1215);
or U1455 (N_1455,In_2782,In_734);
xor U1456 (N_1456,In_2168,In_2494);
nor U1457 (N_1457,In_453,In_2937);
nor U1458 (N_1458,In_1254,In_824);
xor U1459 (N_1459,In_1663,In_695);
nand U1460 (N_1460,In_1909,In_1279);
nor U1461 (N_1461,In_1777,In_2959);
or U1462 (N_1462,In_2178,In_1243);
nor U1463 (N_1463,In_562,In_333);
nand U1464 (N_1464,In_905,In_1881);
nand U1465 (N_1465,In_1232,In_2393);
nor U1466 (N_1466,In_238,In_1195);
nor U1467 (N_1467,In_2909,In_299);
and U1468 (N_1468,In_2112,In_2188);
or U1469 (N_1469,In_1138,In_2073);
xnor U1470 (N_1470,In_1099,In_1795);
and U1471 (N_1471,In_782,In_847);
nand U1472 (N_1472,In_2813,In_1440);
nand U1473 (N_1473,In_380,In_2823);
and U1474 (N_1474,In_1928,In_1435);
nor U1475 (N_1475,In_1725,In_1861);
nor U1476 (N_1476,In_2513,In_2228);
xnor U1477 (N_1477,In_1539,In_786);
or U1478 (N_1478,In_263,In_246);
and U1479 (N_1479,In_809,In_1422);
and U1480 (N_1480,In_1804,In_38);
xnor U1481 (N_1481,In_2881,In_652);
and U1482 (N_1482,In_942,In_2614);
and U1483 (N_1483,In_1567,In_2455);
and U1484 (N_1484,In_2040,In_1513);
and U1485 (N_1485,In_135,In_2964);
or U1486 (N_1486,In_1849,In_1120);
xor U1487 (N_1487,In_2870,In_2348);
nand U1488 (N_1488,In_189,In_1342);
xnor U1489 (N_1489,In_1827,In_2083);
xnor U1490 (N_1490,In_170,In_1183);
or U1491 (N_1491,In_1905,In_1793);
or U1492 (N_1492,In_2551,In_583);
nor U1493 (N_1493,In_2800,In_1095);
xnor U1494 (N_1494,In_1880,In_2049);
xnor U1495 (N_1495,In_2544,In_492);
or U1496 (N_1496,In_830,In_1187);
xor U1497 (N_1497,In_1969,In_535);
nor U1498 (N_1498,In_1423,In_430);
and U1499 (N_1499,In_1785,In_2463);
xor U1500 (N_1500,In_67,In_150);
xor U1501 (N_1501,In_556,In_2837);
nand U1502 (N_1502,In_1114,In_459);
xor U1503 (N_1503,In_785,In_2801);
xor U1504 (N_1504,In_2578,In_632);
xnor U1505 (N_1505,In_142,In_2431);
or U1506 (N_1506,In_2526,In_2142);
nand U1507 (N_1507,In_556,In_1122);
and U1508 (N_1508,In_331,In_1938);
and U1509 (N_1509,In_2931,In_1903);
nand U1510 (N_1510,In_1591,In_413);
nand U1511 (N_1511,In_1939,In_1395);
xor U1512 (N_1512,In_633,In_1818);
nand U1513 (N_1513,In_945,In_2760);
or U1514 (N_1514,In_2830,In_104);
and U1515 (N_1515,In_1734,In_2016);
or U1516 (N_1516,In_547,In_91);
or U1517 (N_1517,In_402,In_2455);
xor U1518 (N_1518,In_1019,In_2061);
or U1519 (N_1519,In_2724,In_480);
and U1520 (N_1520,In_1462,In_355);
nor U1521 (N_1521,In_1609,In_1851);
nor U1522 (N_1522,In_1182,In_2151);
or U1523 (N_1523,In_917,In_2819);
nor U1524 (N_1524,In_459,In_1369);
nand U1525 (N_1525,In_2814,In_1104);
xnor U1526 (N_1526,In_1223,In_666);
nor U1527 (N_1527,In_1456,In_265);
or U1528 (N_1528,In_1331,In_535);
xor U1529 (N_1529,In_629,In_2539);
and U1530 (N_1530,In_1330,In_1287);
nand U1531 (N_1531,In_336,In_912);
xor U1532 (N_1532,In_2638,In_1453);
xor U1533 (N_1533,In_946,In_2763);
xnor U1534 (N_1534,In_1549,In_2776);
or U1535 (N_1535,In_1256,In_1009);
and U1536 (N_1536,In_718,In_1777);
and U1537 (N_1537,In_2191,In_1480);
or U1538 (N_1538,In_508,In_1630);
nor U1539 (N_1539,In_1129,In_2799);
or U1540 (N_1540,In_507,In_1925);
nor U1541 (N_1541,In_1427,In_2403);
or U1542 (N_1542,In_1189,In_171);
and U1543 (N_1543,In_1890,In_2200);
xnor U1544 (N_1544,In_264,In_1145);
nand U1545 (N_1545,In_2137,In_2430);
or U1546 (N_1546,In_170,In_2753);
xnor U1547 (N_1547,In_1745,In_567);
and U1548 (N_1548,In_2335,In_296);
nor U1549 (N_1549,In_2605,In_1312);
nand U1550 (N_1550,In_1093,In_1534);
and U1551 (N_1551,In_310,In_2316);
nor U1552 (N_1552,In_828,In_1884);
nand U1553 (N_1553,In_899,In_792);
and U1554 (N_1554,In_352,In_2413);
nand U1555 (N_1555,In_2300,In_2072);
xor U1556 (N_1556,In_310,In_1308);
nor U1557 (N_1557,In_2958,In_1505);
nor U1558 (N_1558,In_2377,In_2061);
nor U1559 (N_1559,In_893,In_527);
xnor U1560 (N_1560,In_2903,In_1564);
or U1561 (N_1561,In_1714,In_106);
nor U1562 (N_1562,In_1244,In_1577);
nor U1563 (N_1563,In_907,In_1195);
and U1564 (N_1564,In_11,In_1573);
nand U1565 (N_1565,In_1525,In_271);
or U1566 (N_1566,In_641,In_121);
nand U1567 (N_1567,In_1535,In_1519);
or U1568 (N_1568,In_255,In_2485);
or U1569 (N_1569,In_2193,In_921);
or U1570 (N_1570,In_1114,In_418);
xor U1571 (N_1571,In_2214,In_169);
xor U1572 (N_1572,In_766,In_561);
nand U1573 (N_1573,In_1653,In_2786);
and U1574 (N_1574,In_223,In_627);
and U1575 (N_1575,In_926,In_2113);
nor U1576 (N_1576,In_1732,In_257);
nand U1577 (N_1577,In_1973,In_1142);
nor U1578 (N_1578,In_2328,In_2424);
and U1579 (N_1579,In_2539,In_2015);
nor U1580 (N_1580,In_1158,In_945);
and U1581 (N_1581,In_2162,In_1691);
and U1582 (N_1582,In_1063,In_310);
nand U1583 (N_1583,In_301,In_2165);
and U1584 (N_1584,In_1767,In_1852);
and U1585 (N_1585,In_1964,In_846);
xnor U1586 (N_1586,In_1261,In_2879);
nand U1587 (N_1587,In_2530,In_2602);
or U1588 (N_1588,In_1371,In_28);
nand U1589 (N_1589,In_1458,In_867);
nand U1590 (N_1590,In_1907,In_2152);
or U1591 (N_1591,In_2042,In_2722);
or U1592 (N_1592,In_500,In_2089);
nand U1593 (N_1593,In_2199,In_2505);
xnor U1594 (N_1594,In_2760,In_638);
and U1595 (N_1595,In_587,In_357);
xor U1596 (N_1596,In_2309,In_158);
or U1597 (N_1597,In_1530,In_791);
and U1598 (N_1598,In_1514,In_1856);
and U1599 (N_1599,In_78,In_345);
or U1600 (N_1600,In_1288,In_1378);
xnor U1601 (N_1601,In_2190,In_2148);
nor U1602 (N_1602,In_911,In_1041);
xor U1603 (N_1603,In_2054,In_814);
and U1604 (N_1604,In_2826,In_447);
nand U1605 (N_1605,In_848,In_2563);
nor U1606 (N_1606,In_1566,In_862);
and U1607 (N_1607,In_211,In_952);
nor U1608 (N_1608,In_1321,In_606);
xnor U1609 (N_1609,In_1380,In_1297);
nor U1610 (N_1610,In_1665,In_2178);
nor U1611 (N_1611,In_1160,In_64);
and U1612 (N_1612,In_2409,In_555);
and U1613 (N_1613,In_1203,In_1691);
nor U1614 (N_1614,In_1422,In_1823);
nand U1615 (N_1615,In_2518,In_1658);
or U1616 (N_1616,In_489,In_1032);
nor U1617 (N_1617,In_2843,In_2853);
nor U1618 (N_1618,In_2345,In_53);
xnor U1619 (N_1619,In_1047,In_2224);
and U1620 (N_1620,In_1703,In_1835);
nand U1621 (N_1621,In_2365,In_2843);
nor U1622 (N_1622,In_2575,In_1586);
xnor U1623 (N_1623,In_576,In_2625);
or U1624 (N_1624,In_1515,In_507);
or U1625 (N_1625,In_2337,In_688);
nor U1626 (N_1626,In_876,In_2646);
nand U1627 (N_1627,In_2228,In_2258);
and U1628 (N_1628,In_1362,In_44);
xor U1629 (N_1629,In_1132,In_2471);
or U1630 (N_1630,In_790,In_2626);
or U1631 (N_1631,In_2302,In_59);
and U1632 (N_1632,In_2244,In_2924);
xnor U1633 (N_1633,In_2843,In_103);
nand U1634 (N_1634,In_981,In_1316);
and U1635 (N_1635,In_724,In_1841);
xnor U1636 (N_1636,In_1132,In_1038);
xnor U1637 (N_1637,In_2353,In_2309);
or U1638 (N_1638,In_1040,In_1725);
or U1639 (N_1639,In_2261,In_2077);
nor U1640 (N_1640,In_2971,In_1665);
xor U1641 (N_1641,In_2222,In_2432);
or U1642 (N_1642,In_2639,In_1514);
or U1643 (N_1643,In_942,In_2167);
and U1644 (N_1644,In_1705,In_2639);
nand U1645 (N_1645,In_1824,In_347);
xor U1646 (N_1646,In_693,In_162);
or U1647 (N_1647,In_134,In_2022);
nand U1648 (N_1648,In_2585,In_1143);
nand U1649 (N_1649,In_2264,In_546);
nand U1650 (N_1650,In_2619,In_2970);
and U1651 (N_1651,In_1010,In_1931);
xor U1652 (N_1652,In_1542,In_2992);
xor U1653 (N_1653,In_1209,In_1401);
nand U1654 (N_1654,In_2934,In_749);
nand U1655 (N_1655,In_2371,In_1346);
and U1656 (N_1656,In_2367,In_1809);
nand U1657 (N_1657,In_418,In_63);
xnor U1658 (N_1658,In_426,In_357);
nor U1659 (N_1659,In_1262,In_140);
or U1660 (N_1660,In_2450,In_1293);
nand U1661 (N_1661,In_921,In_2729);
nand U1662 (N_1662,In_536,In_2823);
or U1663 (N_1663,In_2198,In_415);
or U1664 (N_1664,In_605,In_385);
and U1665 (N_1665,In_1044,In_2285);
and U1666 (N_1666,In_1182,In_441);
nand U1667 (N_1667,In_1340,In_2111);
or U1668 (N_1668,In_750,In_2063);
xor U1669 (N_1669,In_1501,In_501);
xor U1670 (N_1670,In_2454,In_2699);
or U1671 (N_1671,In_2322,In_2901);
nand U1672 (N_1672,In_416,In_1575);
nand U1673 (N_1673,In_1073,In_1525);
or U1674 (N_1674,In_1589,In_565);
nand U1675 (N_1675,In_1482,In_173);
xnor U1676 (N_1676,In_101,In_1775);
or U1677 (N_1677,In_1487,In_1394);
nor U1678 (N_1678,In_2786,In_1050);
nand U1679 (N_1679,In_587,In_2818);
or U1680 (N_1680,In_2445,In_916);
xnor U1681 (N_1681,In_2799,In_2214);
xor U1682 (N_1682,In_1757,In_913);
nor U1683 (N_1683,In_2154,In_2443);
nor U1684 (N_1684,In_834,In_2125);
and U1685 (N_1685,In_2794,In_147);
nand U1686 (N_1686,In_135,In_2536);
and U1687 (N_1687,In_746,In_2557);
xnor U1688 (N_1688,In_2744,In_1432);
and U1689 (N_1689,In_495,In_816);
nor U1690 (N_1690,In_320,In_459);
nor U1691 (N_1691,In_35,In_1412);
xor U1692 (N_1692,In_2551,In_2784);
or U1693 (N_1693,In_2488,In_2798);
nand U1694 (N_1694,In_2220,In_469);
or U1695 (N_1695,In_1826,In_1335);
nor U1696 (N_1696,In_63,In_2180);
xnor U1697 (N_1697,In_282,In_2391);
and U1698 (N_1698,In_881,In_1520);
xnor U1699 (N_1699,In_1643,In_183);
nor U1700 (N_1700,In_2609,In_593);
and U1701 (N_1701,In_835,In_1478);
or U1702 (N_1702,In_884,In_285);
and U1703 (N_1703,In_41,In_2152);
nor U1704 (N_1704,In_614,In_20);
xor U1705 (N_1705,In_586,In_770);
xnor U1706 (N_1706,In_2495,In_343);
and U1707 (N_1707,In_1515,In_1340);
nand U1708 (N_1708,In_2939,In_1651);
or U1709 (N_1709,In_692,In_651);
nand U1710 (N_1710,In_811,In_1793);
nand U1711 (N_1711,In_861,In_406);
and U1712 (N_1712,In_2116,In_1364);
nand U1713 (N_1713,In_1728,In_1832);
nand U1714 (N_1714,In_1075,In_2109);
nand U1715 (N_1715,In_2485,In_2050);
nor U1716 (N_1716,In_2041,In_1382);
and U1717 (N_1717,In_1816,In_555);
or U1718 (N_1718,In_47,In_1606);
xor U1719 (N_1719,In_2700,In_2388);
nand U1720 (N_1720,In_1920,In_2586);
nor U1721 (N_1721,In_2296,In_142);
nor U1722 (N_1722,In_385,In_100);
and U1723 (N_1723,In_2840,In_997);
nand U1724 (N_1724,In_540,In_2299);
nand U1725 (N_1725,In_1675,In_104);
xor U1726 (N_1726,In_2832,In_1057);
and U1727 (N_1727,In_1536,In_233);
and U1728 (N_1728,In_2335,In_2929);
xor U1729 (N_1729,In_332,In_2703);
or U1730 (N_1730,In_2190,In_189);
or U1731 (N_1731,In_2134,In_419);
nand U1732 (N_1732,In_1569,In_2221);
or U1733 (N_1733,In_70,In_1062);
xnor U1734 (N_1734,In_533,In_2460);
xor U1735 (N_1735,In_286,In_531);
and U1736 (N_1736,In_2096,In_1803);
nor U1737 (N_1737,In_1231,In_2223);
and U1738 (N_1738,In_2008,In_638);
xor U1739 (N_1739,In_1187,In_1907);
or U1740 (N_1740,In_289,In_1741);
and U1741 (N_1741,In_1889,In_886);
xor U1742 (N_1742,In_2492,In_14);
or U1743 (N_1743,In_2918,In_182);
nor U1744 (N_1744,In_356,In_1644);
or U1745 (N_1745,In_1265,In_768);
xnor U1746 (N_1746,In_982,In_2187);
nor U1747 (N_1747,In_2965,In_1639);
and U1748 (N_1748,In_1056,In_942);
xnor U1749 (N_1749,In_2300,In_2652);
nor U1750 (N_1750,In_308,In_2581);
xnor U1751 (N_1751,In_519,In_2370);
nand U1752 (N_1752,In_448,In_1991);
and U1753 (N_1753,In_2812,In_2629);
and U1754 (N_1754,In_2749,In_2014);
and U1755 (N_1755,In_2666,In_1920);
nand U1756 (N_1756,In_1573,In_2399);
nor U1757 (N_1757,In_767,In_349);
nor U1758 (N_1758,In_2560,In_750);
nand U1759 (N_1759,In_1075,In_1882);
xnor U1760 (N_1760,In_735,In_408);
xnor U1761 (N_1761,In_153,In_645);
or U1762 (N_1762,In_519,In_1192);
nor U1763 (N_1763,In_498,In_1893);
nand U1764 (N_1764,In_1479,In_2415);
nand U1765 (N_1765,In_1637,In_663);
nand U1766 (N_1766,In_41,In_2958);
nand U1767 (N_1767,In_1942,In_2531);
xor U1768 (N_1768,In_8,In_41);
or U1769 (N_1769,In_2417,In_1013);
nand U1770 (N_1770,In_1811,In_1791);
or U1771 (N_1771,In_1367,In_1426);
and U1772 (N_1772,In_2607,In_491);
nor U1773 (N_1773,In_2767,In_1191);
nor U1774 (N_1774,In_1375,In_2910);
and U1775 (N_1775,In_2079,In_2691);
nor U1776 (N_1776,In_1309,In_2984);
and U1777 (N_1777,In_1154,In_2250);
nand U1778 (N_1778,In_2211,In_1813);
or U1779 (N_1779,In_1408,In_7);
or U1780 (N_1780,In_2965,In_812);
nor U1781 (N_1781,In_66,In_774);
or U1782 (N_1782,In_173,In_620);
nor U1783 (N_1783,In_1501,In_1212);
nand U1784 (N_1784,In_441,In_2587);
and U1785 (N_1785,In_2254,In_2797);
nor U1786 (N_1786,In_598,In_2944);
nand U1787 (N_1787,In_2828,In_1254);
and U1788 (N_1788,In_2366,In_2960);
nor U1789 (N_1789,In_1249,In_343);
and U1790 (N_1790,In_935,In_1871);
nand U1791 (N_1791,In_168,In_80);
xnor U1792 (N_1792,In_646,In_198);
and U1793 (N_1793,In_15,In_1901);
and U1794 (N_1794,In_1298,In_1693);
nor U1795 (N_1795,In_1853,In_2857);
nor U1796 (N_1796,In_1124,In_2713);
xnor U1797 (N_1797,In_140,In_355);
xnor U1798 (N_1798,In_834,In_2648);
nor U1799 (N_1799,In_1428,In_2179);
xnor U1800 (N_1800,In_1207,In_2264);
nor U1801 (N_1801,In_2141,In_2352);
xor U1802 (N_1802,In_1339,In_2598);
and U1803 (N_1803,In_1822,In_1026);
or U1804 (N_1804,In_2,In_563);
and U1805 (N_1805,In_2197,In_2605);
nand U1806 (N_1806,In_325,In_1831);
xor U1807 (N_1807,In_2299,In_2827);
nand U1808 (N_1808,In_2128,In_2948);
or U1809 (N_1809,In_355,In_242);
or U1810 (N_1810,In_1786,In_725);
and U1811 (N_1811,In_941,In_2948);
nor U1812 (N_1812,In_1842,In_1617);
xnor U1813 (N_1813,In_215,In_2175);
nand U1814 (N_1814,In_803,In_185);
xor U1815 (N_1815,In_152,In_1688);
nor U1816 (N_1816,In_2144,In_2493);
nor U1817 (N_1817,In_2570,In_847);
xnor U1818 (N_1818,In_1613,In_1809);
or U1819 (N_1819,In_1757,In_619);
nand U1820 (N_1820,In_261,In_983);
and U1821 (N_1821,In_1675,In_2268);
and U1822 (N_1822,In_835,In_1641);
nand U1823 (N_1823,In_2149,In_2900);
nor U1824 (N_1824,In_808,In_2343);
or U1825 (N_1825,In_1455,In_1961);
nand U1826 (N_1826,In_2197,In_1503);
and U1827 (N_1827,In_1456,In_1498);
nor U1828 (N_1828,In_2302,In_466);
xnor U1829 (N_1829,In_2285,In_2920);
or U1830 (N_1830,In_2978,In_2243);
and U1831 (N_1831,In_1634,In_141);
nor U1832 (N_1832,In_1474,In_654);
nand U1833 (N_1833,In_358,In_587);
and U1834 (N_1834,In_1767,In_14);
or U1835 (N_1835,In_488,In_313);
or U1836 (N_1836,In_173,In_1818);
xnor U1837 (N_1837,In_1383,In_1478);
nand U1838 (N_1838,In_536,In_1803);
and U1839 (N_1839,In_2458,In_1607);
and U1840 (N_1840,In_2978,In_448);
xnor U1841 (N_1841,In_5,In_90);
or U1842 (N_1842,In_2263,In_2624);
and U1843 (N_1843,In_2193,In_1862);
nand U1844 (N_1844,In_2596,In_1349);
nor U1845 (N_1845,In_642,In_2238);
nor U1846 (N_1846,In_1045,In_102);
nand U1847 (N_1847,In_2901,In_1885);
or U1848 (N_1848,In_169,In_2359);
and U1849 (N_1849,In_1002,In_1258);
or U1850 (N_1850,In_672,In_1662);
or U1851 (N_1851,In_919,In_2211);
nor U1852 (N_1852,In_2766,In_2214);
xor U1853 (N_1853,In_1164,In_108);
and U1854 (N_1854,In_2550,In_535);
nand U1855 (N_1855,In_541,In_742);
or U1856 (N_1856,In_635,In_2026);
or U1857 (N_1857,In_2326,In_118);
xnor U1858 (N_1858,In_735,In_1893);
xnor U1859 (N_1859,In_1804,In_279);
or U1860 (N_1860,In_2325,In_2421);
nand U1861 (N_1861,In_159,In_2642);
xor U1862 (N_1862,In_1784,In_1886);
and U1863 (N_1863,In_1082,In_310);
xnor U1864 (N_1864,In_2134,In_1671);
xnor U1865 (N_1865,In_554,In_2242);
or U1866 (N_1866,In_795,In_1039);
and U1867 (N_1867,In_1451,In_1325);
xor U1868 (N_1868,In_2333,In_610);
nor U1869 (N_1869,In_2751,In_1680);
and U1870 (N_1870,In_1656,In_189);
xnor U1871 (N_1871,In_2314,In_1298);
nand U1872 (N_1872,In_542,In_2719);
xnor U1873 (N_1873,In_607,In_340);
or U1874 (N_1874,In_921,In_1002);
nand U1875 (N_1875,In_1114,In_2279);
xnor U1876 (N_1876,In_600,In_432);
nand U1877 (N_1877,In_1293,In_1219);
nor U1878 (N_1878,In_2163,In_2824);
nor U1879 (N_1879,In_2022,In_938);
xnor U1880 (N_1880,In_2908,In_1541);
or U1881 (N_1881,In_1182,In_2280);
or U1882 (N_1882,In_2328,In_2644);
nand U1883 (N_1883,In_197,In_2551);
xnor U1884 (N_1884,In_61,In_2082);
nand U1885 (N_1885,In_471,In_616);
nor U1886 (N_1886,In_1167,In_860);
and U1887 (N_1887,In_1765,In_87);
and U1888 (N_1888,In_1030,In_1824);
nand U1889 (N_1889,In_1732,In_1742);
xor U1890 (N_1890,In_2320,In_709);
xor U1891 (N_1891,In_2783,In_425);
nand U1892 (N_1892,In_1353,In_854);
nand U1893 (N_1893,In_2390,In_2933);
or U1894 (N_1894,In_1366,In_1080);
nor U1895 (N_1895,In_1687,In_195);
nand U1896 (N_1896,In_864,In_2238);
xor U1897 (N_1897,In_2373,In_430);
nand U1898 (N_1898,In_2639,In_1581);
nor U1899 (N_1899,In_2141,In_284);
and U1900 (N_1900,In_560,In_625);
xnor U1901 (N_1901,In_2256,In_2040);
nand U1902 (N_1902,In_1052,In_2479);
xnor U1903 (N_1903,In_1862,In_136);
nand U1904 (N_1904,In_2773,In_2446);
or U1905 (N_1905,In_1937,In_796);
nand U1906 (N_1906,In_991,In_2911);
nor U1907 (N_1907,In_2573,In_1700);
nand U1908 (N_1908,In_253,In_2905);
xor U1909 (N_1909,In_1229,In_283);
nand U1910 (N_1910,In_1870,In_2673);
nor U1911 (N_1911,In_138,In_2899);
and U1912 (N_1912,In_2715,In_1433);
and U1913 (N_1913,In_396,In_2164);
nor U1914 (N_1914,In_2946,In_2510);
xor U1915 (N_1915,In_1769,In_966);
xnor U1916 (N_1916,In_2096,In_1386);
nor U1917 (N_1917,In_2248,In_2331);
and U1918 (N_1918,In_2508,In_2794);
or U1919 (N_1919,In_1900,In_954);
nor U1920 (N_1920,In_2060,In_2470);
or U1921 (N_1921,In_2053,In_55);
nor U1922 (N_1922,In_381,In_94);
nand U1923 (N_1923,In_668,In_152);
or U1924 (N_1924,In_184,In_773);
nand U1925 (N_1925,In_2838,In_2790);
xor U1926 (N_1926,In_2484,In_1140);
or U1927 (N_1927,In_740,In_1282);
xor U1928 (N_1928,In_1568,In_1189);
or U1929 (N_1929,In_15,In_497);
or U1930 (N_1930,In_915,In_361);
xor U1931 (N_1931,In_209,In_588);
and U1932 (N_1932,In_2904,In_1652);
nor U1933 (N_1933,In_2149,In_2659);
nor U1934 (N_1934,In_1224,In_468);
nor U1935 (N_1935,In_2632,In_1958);
nand U1936 (N_1936,In_1881,In_79);
nor U1937 (N_1937,In_806,In_784);
xor U1938 (N_1938,In_28,In_448);
and U1939 (N_1939,In_2587,In_2788);
nor U1940 (N_1940,In_86,In_549);
or U1941 (N_1941,In_2253,In_342);
and U1942 (N_1942,In_110,In_2390);
and U1943 (N_1943,In_2782,In_2599);
or U1944 (N_1944,In_2408,In_68);
or U1945 (N_1945,In_2569,In_221);
or U1946 (N_1946,In_2574,In_1957);
or U1947 (N_1947,In_1316,In_1371);
and U1948 (N_1948,In_1951,In_620);
and U1949 (N_1949,In_2191,In_2625);
nor U1950 (N_1950,In_2687,In_1441);
and U1951 (N_1951,In_1886,In_2252);
and U1952 (N_1952,In_873,In_820);
xnor U1953 (N_1953,In_1390,In_2278);
xnor U1954 (N_1954,In_1265,In_1331);
or U1955 (N_1955,In_195,In_1569);
and U1956 (N_1956,In_638,In_2312);
nor U1957 (N_1957,In_1503,In_1497);
nand U1958 (N_1958,In_7,In_2041);
or U1959 (N_1959,In_687,In_2239);
nor U1960 (N_1960,In_1201,In_2029);
and U1961 (N_1961,In_586,In_2423);
xnor U1962 (N_1962,In_1301,In_191);
xor U1963 (N_1963,In_2501,In_1122);
nand U1964 (N_1964,In_482,In_747);
or U1965 (N_1965,In_1623,In_1150);
xnor U1966 (N_1966,In_1688,In_1923);
nand U1967 (N_1967,In_621,In_2420);
xnor U1968 (N_1968,In_1181,In_2830);
or U1969 (N_1969,In_379,In_2937);
xnor U1970 (N_1970,In_2257,In_1494);
xor U1971 (N_1971,In_375,In_135);
nand U1972 (N_1972,In_2857,In_2601);
nand U1973 (N_1973,In_1474,In_304);
and U1974 (N_1974,In_1251,In_1019);
xor U1975 (N_1975,In_851,In_2649);
or U1976 (N_1976,In_2454,In_1977);
nor U1977 (N_1977,In_498,In_1607);
nor U1978 (N_1978,In_1242,In_495);
nor U1979 (N_1979,In_2331,In_2873);
nand U1980 (N_1980,In_430,In_829);
or U1981 (N_1981,In_0,In_2088);
nor U1982 (N_1982,In_1660,In_1969);
nand U1983 (N_1983,In_1338,In_1489);
xor U1984 (N_1984,In_2126,In_2724);
and U1985 (N_1985,In_777,In_435);
or U1986 (N_1986,In_1118,In_1609);
or U1987 (N_1987,In_24,In_1180);
nand U1988 (N_1988,In_938,In_883);
and U1989 (N_1989,In_344,In_2799);
or U1990 (N_1990,In_1697,In_1557);
and U1991 (N_1991,In_522,In_1966);
and U1992 (N_1992,In_199,In_1166);
or U1993 (N_1993,In_2402,In_1503);
nor U1994 (N_1994,In_2769,In_237);
nand U1995 (N_1995,In_2078,In_2097);
nor U1996 (N_1996,In_2676,In_304);
xor U1997 (N_1997,In_1393,In_1734);
nand U1998 (N_1998,In_1263,In_2572);
or U1999 (N_1999,In_481,In_2221);
or U2000 (N_2000,In_1611,In_2274);
xor U2001 (N_2001,In_2571,In_2599);
xnor U2002 (N_2002,In_1991,In_957);
and U2003 (N_2003,In_1536,In_2120);
xor U2004 (N_2004,In_2545,In_1301);
and U2005 (N_2005,In_605,In_2286);
nor U2006 (N_2006,In_2840,In_272);
nand U2007 (N_2007,In_2628,In_1650);
or U2008 (N_2008,In_1174,In_1415);
and U2009 (N_2009,In_2534,In_2033);
and U2010 (N_2010,In_2165,In_2527);
or U2011 (N_2011,In_2469,In_953);
nor U2012 (N_2012,In_2475,In_1428);
nor U2013 (N_2013,In_575,In_1305);
xnor U2014 (N_2014,In_1536,In_1521);
and U2015 (N_2015,In_310,In_1391);
nand U2016 (N_2016,In_2534,In_317);
and U2017 (N_2017,In_1741,In_503);
and U2018 (N_2018,In_1807,In_2754);
nand U2019 (N_2019,In_1595,In_1628);
nor U2020 (N_2020,In_1716,In_1963);
xnor U2021 (N_2021,In_2210,In_335);
xor U2022 (N_2022,In_393,In_953);
nor U2023 (N_2023,In_1711,In_2228);
and U2024 (N_2024,In_433,In_2919);
nor U2025 (N_2025,In_374,In_2816);
or U2026 (N_2026,In_2784,In_2041);
or U2027 (N_2027,In_1925,In_657);
and U2028 (N_2028,In_52,In_1377);
nor U2029 (N_2029,In_287,In_2645);
nor U2030 (N_2030,In_2380,In_2995);
nor U2031 (N_2031,In_1540,In_828);
or U2032 (N_2032,In_1728,In_1194);
or U2033 (N_2033,In_1809,In_299);
and U2034 (N_2034,In_2893,In_2336);
xor U2035 (N_2035,In_1749,In_2951);
or U2036 (N_2036,In_1252,In_540);
and U2037 (N_2037,In_354,In_2394);
nor U2038 (N_2038,In_434,In_452);
nor U2039 (N_2039,In_2501,In_1634);
or U2040 (N_2040,In_2304,In_2985);
nor U2041 (N_2041,In_2155,In_1237);
and U2042 (N_2042,In_1784,In_1875);
or U2043 (N_2043,In_1018,In_2727);
nand U2044 (N_2044,In_2852,In_2898);
nand U2045 (N_2045,In_2066,In_2247);
nor U2046 (N_2046,In_2624,In_604);
nand U2047 (N_2047,In_2986,In_1470);
or U2048 (N_2048,In_1773,In_2893);
nor U2049 (N_2049,In_201,In_2622);
nor U2050 (N_2050,In_1224,In_2554);
nand U2051 (N_2051,In_1374,In_2756);
nand U2052 (N_2052,In_2382,In_965);
nand U2053 (N_2053,In_2135,In_1797);
nand U2054 (N_2054,In_781,In_2510);
and U2055 (N_2055,In_1607,In_829);
and U2056 (N_2056,In_308,In_2997);
xnor U2057 (N_2057,In_1417,In_1113);
and U2058 (N_2058,In_759,In_332);
nor U2059 (N_2059,In_2942,In_1337);
or U2060 (N_2060,In_1268,In_1699);
or U2061 (N_2061,In_1907,In_1683);
xnor U2062 (N_2062,In_561,In_2342);
nor U2063 (N_2063,In_209,In_789);
or U2064 (N_2064,In_461,In_470);
nand U2065 (N_2065,In_2761,In_1570);
or U2066 (N_2066,In_1021,In_2929);
nand U2067 (N_2067,In_112,In_2557);
and U2068 (N_2068,In_1369,In_953);
or U2069 (N_2069,In_175,In_2439);
or U2070 (N_2070,In_317,In_1852);
and U2071 (N_2071,In_1723,In_2442);
and U2072 (N_2072,In_1047,In_1585);
nor U2073 (N_2073,In_437,In_607);
or U2074 (N_2074,In_1021,In_2920);
or U2075 (N_2075,In_292,In_297);
or U2076 (N_2076,In_613,In_1898);
nor U2077 (N_2077,In_984,In_53);
nor U2078 (N_2078,In_1025,In_2602);
xor U2079 (N_2079,In_2334,In_1211);
nor U2080 (N_2080,In_1620,In_2818);
or U2081 (N_2081,In_2405,In_2708);
and U2082 (N_2082,In_1661,In_356);
and U2083 (N_2083,In_564,In_775);
and U2084 (N_2084,In_1936,In_1091);
xor U2085 (N_2085,In_151,In_2714);
nor U2086 (N_2086,In_2041,In_115);
nor U2087 (N_2087,In_2198,In_499);
and U2088 (N_2088,In_23,In_2499);
nand U2089 (N_2089,In_2460,In_1811);
nand U2090 (N_2090,In_2733,In_1749);
or U2091 (N_2091,In_2969,In_227);
and U2092 (N_2092,In_1961,In_1106);
nor U2093 (N_2093,In_969,In_1323);
nand U2094 (N_2094,In_2530,In_1809);
nand U2095 (N_2095,In_2736,In_925);
or U2096 (N_2096,In_1064,In_246);
xor U2097 (N_2097,In_63,In_1790);
nor U2098 (N_2098,In_1031,In_2538);
and U2099 (N_2099,In_1646,In_800);
nand U2100 (N_2100,In_2637,In_1793);
nor U2101 (N_2101,In_235,In_2238);
and U2102 (N_2102,In_1329,In_1508);
nor U2103 (N_2103,In_791,In_433);
nand U2104 (N_2104,In_1122,In_2723);
or U2105 (N_2105,In_2609,In_2025);
and U2106 (N_2106,In_1722,In_2409);
nand U2107 (N_2107,In_2193,In_507);
and U2108 (N_2108,In_976,In_1929);
or U2109 (N_2109,In_2838,In_907);
and U2110 (N_2110,In_713,In_2776);
and U2111 (N_2111,In_1725,In_1372);
nand U2112 (N_2112,In_2004,In_1085);
nor U2113 (N_2113,In_1589,In_888);
nand U2114 (N_2114,In_167,In_303);
and U2115 (N_2115,In_729,In_1174);
nand U2116 (N_2116,In_2424,In_2504);
and U2117 (N_2117,In_634,In_509);
and U2118 (N_2118,In_1624,In_2191);
xnor U2119 (N_2119,In_2965,In_2573);
nand U2120 (N_2120,In_2151,In_378);
nand U2121 (N_2121,In_1285,In_737);
nand U2122 (N_2122,In_1401,In_2370);
nand U2123 (N_2123,In_2068,In_2733);
nor U2124 (N_2124,In_2739,In_2976);
nand U2125 (N_2125,In_581,In_1462);
and U2126 (N_2126,In_1362,In_1048);
or U2127 (N_2127,In_1000,In_2901);
and U2128 (N_2128,In_1194,In_958);
nor U2129 (N_2129,In_505,In_1463);
nand U2130 (N_2130,In_2281,In_2192);
and U2131 (N_2131,In_820,In_368);
and U2132 (N_2132,In_2622,In_2513);
or U2133 (N_2133,In_2083,In_186);
nand U2134 (N_2134,In_1624,In_777);
nand U2135 (N_2135,In_1895,In_1893);
nand U2136 (N_2136,In_2198,In_1063);
nor U2137 (N_2137,In_2626,In_860);
nand U2138 (N_2138,In_1486,In_278);
or U2139 (N_2139,In_129,In_2079);
nand U2140 (N_2140,In_138,In_2914);
xor U2141 (N_2141,In_414,In_1785);
and U2142 (N_2142,In_1206,In_351);
xnor U2143 (N_2143,In_2347,In_1208);
or U2144 (N_2144,In_1840,In_812);
or U2145 (N_2145,In_2910,In_1934);
and U2146 (N_2146,In_2240,In_1488);
or U2147 (N_2147,In_353,In_2756);
nor U2148 (N_2148,In_2075,In_1894);
nand U2149 (N_2149,In_1491,In_728);
nor U2150 (N_2150,In_174,In_7);
nand U2151 (N_2151,In_2204,In_392);
or U2152 (N_2152,In_2661,In_4);
or U2153 (N_2153,In_574,In_1934);
nor U2154 (N_2154,In_91,In_2543);
and U2155 (N_2155,In_536,In_529);
nand U2156 (N_2156,In_824,In_957);
nand U2157 (N_2157,In_2644,In_1932);
nor U2158 (N_2158,In_2407,In_304);
and U2159 (N_2159,In_1214,In_1160);
xor U2160 (N_2160,In_1876,In_2788);
nand U2161 (N_2161,In_1560,In_1789);
and U2162 (N_2162,In_2402,In_2215);
xor U2163 (N_2163,In_2516,In_2961);
nor U2164 (N_2164,In_637,In_2977);
and U2165 (N_2165,In_2354,In_1912);
nor U2166 (N_2166,In_308,In_2102);
nor U2167 (N_2167,In_970,In_1749);
xnor U2168 (N_2168,In_835,In_1575);
nor U2169 (N_2169,In_1213,In_1125);
nand U2170 (N_2170,In_1533,In_2304);
xnor U2171 (N_2171,In_1978,In_2704);
nand U2172 (N_2172,In_333,In_2061);
and U2173 (N_2173,In_494,In_1505);
and U2174 (N_2174,In_1562,In_2708);
nand U2175 (N_2175,In_538,In_852);
nand U2176 (N_2176,In_2051,In_1750);
and U2177 (N_2177,In_1323,In_2025);
nand U2178 (N_2178,In_650,In_479);
nand U2179 (N_2179,In_426,In_471);
xor U2180 (N_2180,In_1167,In_1362);
and U2181 (N_2181,In_326,In_163);
nand U2182 (N_2182,In_290,In_1365);
xnor U2183 (N_2183,In_2122,In_1366);
nand U2184 (N_2184,In_2303,In_224);
nor U2185 (N_2185,In_36,In_321);
or U2186 (N_2186,In_1862,In_2195);
xor U2187 (N_2187,In_2559,In_569);
nand U2188 (N_2188,In_2443,In_2083);
nor U2189 (N_2189,In_1239,In_1175);
nor U2190 (N_2190,In_1563,In_887);
and U2191 (N_2191,In_2061,In_17);
nor U2192 (N_2192,In_1615,In_910);
nor U2193 (N_2193,In_2509,In_249);
xnor U2194 (N_2194,In_1783,In_2811);
nor U2195 (N_2195,In_1973,In_2163);
nor U2196 (N_2196,In_1907,In_2649);
nand U2197 (N_2197,In_1527,In_2060);
and U2198 (N_2198,In_2021,In_2799);
nand U2199 (N_2199,In_1298,In_2170);
nor U2200 (N_2200,In_1411,In_1424);
xnor U2201 (N_2201,In_2979,In_1915);
xnor U2202 (N_2202,In_1421,In_1355);
and U2203 (N_2203,In_2608,In_756);
nor U2204 (N_2204,In_143,In_300);
xnor U2205 (N_2205,In_913,In_944);
xor U2206 (N_2206,In_2994,In_1717);
nor U2207 (N_2207,In_1506,In_2214);
nand U2208 (N_2208,In_624,In_2186);
xor U2209 (N_2209,In_2708,In_2621);
nand U2210 (N_2210,In_371,In_2492);
or U2211 (N_2211,In_129,In_2129);
nand U2212 (N_2212,In_2471,In_2350);
and U2213 (N_2213,In_366,In_2413);
nor U2214 (N_2214,In_182,In_1597);
and U2215 (N_2215,In_1276,In_1099);
xor U2216 (N_2216,In_715,In_20);
and U2217 (N_2217,In_232,In_999);
and U2218 (N_2218,In_2348,In_1941);
nand U2219 (N_2219,In_2735,In_830);
xnor U2220 (N_2220,In_1714,In_2163);
or U2221 (N_2221,In_2309,In_1434);
nand U2222 (N_2222,In_2747,In_152);
and U2223 (N_2223,In_1484,In_234);
or U2224 (N_2224,In_1523,In_1689);
and U2225 (N_2225,In_819,In_2736);
xnor U2226 (N_2226,In_2212,In_2451);
xnor U2227 (N_2227,In_2496,In_1567);
nor U2228 (N_2228,In_252,In_1666);
or U2229 (N_2229,In_194,In_893);
nand U2230 (N_2230,In_667,In_349);
nand U2231 (N_2231,In_310,In_1643);
xor U2232 (N_2232,In_2983,In_1151);
xor U2233 (N_2233,In_2447,In_1997);
nand U2234 (N_2234,In_1396,In_2482);
or U2235 (N_2235,In_922,In_2689);
or U2236 (N_2236,In_2031,In_1540);
xor U2237 (N_2237,In_1673,In_2695);
nand U2238 (N_2238,In_1211,In_942);
nand U2239 (N_2239,In_2828,In_2664);
or U2240 (N_2240,In_1158,In_2337);
and U2241 (N_2241,In_1999,In_1094);
nand U2242 (N_2242,In_1086,In_1016);
nand U2243 (N_2243,In_2939,In_253);
or U2244 (N_2244,In_2718,In_2659);
and U2245 (N_2245,In_2311,In_2732);
or U2246 (N_2246,In_2126,In_2807);
nor U2247 (N_2247,In_2786,In_2735);
or U2248 (N_2248,In_2864,In_2022);
nand U2249 (N_2249,In_2983,In_2635);
nor U2250 (N_2250,In_250,In_838);
or U2251 (N_2251,In_298,In_1623);
nand U2252 (N_2252,In_2331,In_2076);
or U2253 (N_2253,In_377,In_658);
xor U2254 (N_2254,In_1815,In_1089);
nor U2255 (N_2255,In_1393,In_1334);
nand U2256 (N_2256,In_304,In_750);
nor U2257 (N_2257,In_2793,In_2312);
nor U2258 (N_2258,In_2573,In_631);
and U2259 (N_2259,In_1777,In_1531);
nor U2260 (N_2260,In_2720,In_1893);
nand U2261 (N_2261,In_1657,In_2391);
and U2262 (N_2262,In_516,In_2376);
xnor U2263 (N_2263,In_2042,In_43);
and U2264 (N_2264,In_1084,In_1708);
and U2265 (N_2265,In_438,In_2146);
nand U2266 (N_2266,In_2654,In_2209);
and U2267 (N_2267,In_2125,In_2681);
and U2268 (N_2268,In_1687,In_999);
nor U2269 (N_2269,In_289,In_209);
xor U2270 (N_2270,In_1220,In_2522);
xor U2271 (N_2271,In_2771,In_859);
and U2272 (N_2272,In_612,In_261);
nor U2273 (N_2273,In_236,In_2725);
and U2274 (N_2274,In_1265,In_1039);
and U2275 (N_2275,In_2174,In_2177);
xor U2276 (N_2276,In_2515,In_1570);
xnor U2277 (N_2277,In_2356,In_2226);
or U2278 (N_2278,In_1451,In_1618);
and U2279 (N_2279,In_2995,In_1650);
and U2280 (N_2280,In_319,In_1211);
or U2281 (N_2281,In_2584,In_365);
or U2282 (N_2282,In_502,In_1550);
or U2283 (N_2283,In_2041,In_1994);
xor U2284 (N_2284,In_1413,In_697);
nand U2285 (N_2285,In_1399,In_1910);
nand U2286 (N_2286,In_1336,In_332);
nand U2287 (N_2287,In_1575,In_131);
or U2288 (N_2288,In_565,In_2445);
nor U2289 (N_2289,In_1113,In_459);
nand U2290 (N_2290,In_1618,In_2579);
and U2291 (N_2291,In_2089,In_256);
nor U2292 (N_2292,In_345,In_309);
nor U2293 (N_2293,In_2684,In_1957);
xnor U2294 (N_2294,In_2495,In_1496);
and U2295 (N_2295,In_1379,In_84);
nand U2296 (N_2296,In_2649,In_2921);
xnor U2297 (N_2297,In_2909,In_2805);
nand U2298 (N_2298,In_2176,In_237);
and U2299 (N_2299,In_278,In_2712);
or U2300 (N_2300,In_247,In_703);
nand U2301 (N_2301,In_678,In_2470);
and U2302 (N_2302,In_1366,In_543);
nor U2303 (N_2303,In_383,In_1598);
and U2304 (N_2304,In_1918,In_610);
nand U2305 (N_2305,In_612,In_1573);
xor U2306 (N_2306,In_79,In_1253);
xnor U2307 (N_2307,In_905,In_415);
xnor U2308 (N_2308,In_2204,In_2635);
nor U2309 (N_2309,In_2646,In_1682);
xnor U2310 (N_2310,In_871,In_688);
xor U2311 (N_2311,In_695,In_310);
nor U2312 (N_2312,In_300,In_1671);
nand U2313 (N_2313,In_687,In_2444);
and U2314 (N_2314,In_2594,In_1611);
nor U2315 (N_2315,In_2086,In_1540);
and U2316 (N_2316,In_729,In_1633);
or U2317 (N_2317,In_386,In_1096);
xor U2318 (N_2318,In_1170,In_239);
or U2319 (N_2319,In_409,In_1115);
or U2320 (N_2320,In_1124,In_1008);
xor U2321 (N_2321,In_1558,In_877);
nor U2322 (N_2322,In_2467,In_1770);
nand U2323 (N_2323,In_986,In_2920);
nor U2324 (N_2324,In_2569,In_2130);
and U2325 (N_2325,In_1957,In_2241);
nor U2326 (N_2326,In_536,In_2764);
nor U2327 (N_2327,In_2598,In_686);
nor U2328 (N_2328,In_195,In_383);
nor U2329 (N_2329,In_1225,In_812);
xnor U2330 (N_2330,In_352,In_105);
or U2331 (N_2331,In_2309,In_237);
nor U2332 (N_2332,In_974,In_1081);
or U2333 (N_2333,In_842,In_1023);
and U2334 (N_2334,In_2309,In_574);
nand U2335 (N_2335,In_2440,In_2403);
xor U2336 (N_2336,In_665,In_1915);
or U2337 (N_2337,In_344,In_2839);
nand U2338 (N_2338,In_1255,In_2268);
or U2339 (N_2339,In_47,In_1629);
or U2340 (N_2340,In_2427,In_2733);
and U2341 (N_2341,In_1791,In_2286);
nand U2342 (N_2342,In_965,In_2896);
or U2343 (N_2343,In_1506,In_1649);
or U2344 (N_2344,In_2062,In_2159);
and U2345 (N_2345,In_2462,In_2828);
and U2346 (N_2346,In_173,In_1746);
and U2347 (N_2347,In_2091,In_651);
xnor U2348 (N_2348,In_381,In_308);
nand U2349 (N_2349,In_1391,In_809);
xnor U2350 (N_2350,In_1873,In_2309);
nor U2351 (N_2351,In_1691,In_2157);
and U2352 (N_2352,In_2686,In_1338);
and U2353 (N_2353,In_537,In_1588);
or U2354 (N_2354,In_187,In_388);
and U2355 (N_2355,In_120,In_1463);
and U2356 (N_2356,In_1299,In_1908);
nor U2357 (N_2357,In_2582,In_1589);
or U2358 (N_2358,In_1614,In_1443);
nor U2359 (N_2359,In_2840,In_646);
nor U2360 (N_2360,In_1615,In_1656);
nor U2361 (N_2361,In_2581,In_1569);
and U2362 (N_2362,In_672,In_2145);
and U2363 (N_2363,In_2016,In_1541);
nand U2364 (N_2364,In_1632,In_2355);
nor U2365 (N_2365,In_2771,In_2658);
nand U2366 (N_2366,In_136,In_1078);
nor U2367 (N_2367,In_2769,In_2286);
nor U2368 (N_2368,In_284,In_1513);
nor U2369 (N_2369,In_1403,In_2705);
nand U2370 (N_2370,In_2363,In_2088);
nor U2371 (N_2371,In_1378,In_884);
and U2372 (N_2372,In_1343,In_156);
nand U2373 (N_2373,In_176,In_1245);
nor U2374 (N_2374,In_2774,In_1838);
nor U2375 (N_2375,In_1501,In_1785);
nand U2376 (N_2376,In_1165,In_432);
and U2377 (N_2377,In_1887,In_500);
and U2378 (N_2378,In_1353,In_2566);
nand U2379 (N_2379,In_2621,In_2132);
or U2380 (N_2380,In_2299,In_583);
and U2381 (N_2381,In_2554,In_1964);
and U2382 (N_2382,In_331,In_727);
or U2383 (N_2383,In_295,In_20);
nor U2384 (N_2384,In_2084,In_298);
nand U2385 (N_2385,In_1976,In_2837);
or U2386 (N_2386,In_2066,In_53);
and U2387 (N_2387,In_2948,In_965);
xor U2388 (N_2388,In_2790,In_216);
nor U2389 (N_2389,In_1230,In_2900);
nor U2390 (N_2390,In_429,In_702);
nand U2391 (N_2391,In_2144,In_212);
and U2392 (N_2392,In_1838,In_1615);
xnor U2393 (N_2393,In_1134,In_1532);
xnor U2394 (N_2394,In_914,In_2815);
xor U2395 (N_2395,In_2738,In_2155);
xnor U2396 (N_2396,In_432,In_1259);
or U2397 (N_2397,In_193,In_2270);
or U2398 (N_2398,In_2568,In_2201);
or U2399 (N_2399,In_2413,In_1673);
nor U2400 (N_2400,In_1787,In_1614);
nor U2401 (N_2401,In_407,In_817);
nor U2402 (N_2402,In_865,In_2048);
or U2403 (N_2403,In_690,In_1562);
and U2404 (N_2404,In_962,In_2009);
nand U2405 (N_2405,In_2889,In_2906);
nand U2406 (N_2406,In_183,In_1180);
nor U2407 (N_2407,In_2415,In_2615);
and U2408 (N_2408,In_1779,In_1446);
xnor U2409 (N_2409,In_998,In_1570);
nor U2410 (N_2410,In_2461,In_581);
nor U2411 (N_2411,In_366,In_2944);
xnor U2412 (N_2412,In_1035,In_2862);
nand U2413 (N_2413,In_2092,In_1224);
and U2414 (N_2414,In_1268,In_300);
or U2415 (N_2415,In_2278,In_2846);
nand U2416 (N_2416,In_500,In_709);
nor U2417 (N_2417,In_2321,In_733);
xnor U2418 (N_2418,In_2838,In_2295);
or U2419 (N_2419,In_2262,In_1764);
and U2420 (N_2420,In_243,In_1300);
nand U2421 (N_2421,In_1501,In_1367);
and U2422 (N_2422,In_936,In_367);
or U2423 (N_2423,In_2979,In_295);
or U2424 (N_2424,In_2974,In_2933);
and U2425 (N_2425,In_1652,In_1637);
nand U2426 (N_2426,In_1155,In_1329);
or U2427 (N_2427,In_2055,In_677);
or U2428 (N_2428,In_503,In_2290);
nand U2429 (N_2429,In_1793,In_2808);
or U2430 (N_2430,In_1120,In_2195);
and U2431 (N_2431,In_652,In_800);
nand U2432 (N_2432,In_743,In_1354);
xor U2433 (N_2433,In_2520,In_516);
xnor U2434 (N_2434,In_1277,In_2087);
or U2435 (N_2435,In_1696,In_2178);
nor U2436 (N_2436,In_258,In_880);
and U2437 (N_2437,In_2437,In_1187);
nor U2438 (N_2438,In_212,In_1452);
xor U2439 (N_2439,In_1746,In_1638);
or U2440 (N_2440,In_1077,In_2404);
or U2441 (N_2441,In_1776,In_517);
xnor U2442 (N_2442,In_1454,In_2600);
nor U2443 (N_2443,In_2680,In_1502);
and U2444 (N_2444,In_1254,In_422);
nor U2445 (N_2445,In_2056,In_157);
xor U2446 (N_2446,In_1951,In_150);
xor U2447 (N_2447,In_373,In_1739);
nor U2448 (N_2448,In_2438,In_1567);
or U2449 (N_2449,In_1712,In_436);
and U2450 (N_2450,In_1365,In_784);
or U2451 (N_2451,In_2616,In_2902);
and U2452 (N_2452,In_816,In_1305);
and U2453 (N_2453,In_1287,In_1944);
or U2454 (N_2454,In_1796,In_73);
nor U2455 (N_2455,In_710,In_758);
or U2456 (N_2456,In_1583,In_2374);
and U2457 (N_2457,In_592,In_1414);
and U2458 (N_2458,In_654,In_1920);
nor U2459 (N_2459,In_93,In_2256);
and U2460 (N_2460,In_1251,In_2298);
and U2461 (N_2461,In_2154,In_2303);
and U2462 (N_2462,In_365,In_782);
nor U2463 (N_2463,In_694,In_684);
and U2464 (N_2464,In_142,In_2537);
nand U2465 (N_2465,In_992,In_1601);
and U2466 (N_2466,In_2259,In_1812);
nor U2467 (N_2467,In_624,In_2291);
or U2468 (N_2468,In_701,In_2373);
xnor U2469 (N_2469,In_2719,In_1962);
xnor U2470 (N_2470,In_784,In_1829);
nand U2471 (N_2471,In_2859,In_934);
xor U2472 (N_2472,In_971,In_2949);
xor U2473 (N_2473,In_1914,In_40);
nand U2474 (N_2474,In_863,In_1534);
or U2475 (N_2475,In_1477,In_2833);
nor U2476 (N_2476,In_1717,In_1919);
xnor U2477 (N_2477,In_2969,In_871);
xnor U2478 (N_2478,In_2187,In_1701);
nor U2479 (N_2479,In_1122,In_2239);
nor U2480 (N_2480,In_801,In_2735);
xor U2481 (N_2481,In_2586,In_1148);
or U2482 (N_2482,In_1842,In_2244);
nand U2483 (N_2483,In_1713,In_15);
xnor U2484 (N_2484,In_2418,In_2975);
xor U2485 (N_2485,In_2956,In_229);
xor U2486 (N_2486,In_2112,In_2674);
nand U2487 (N_2487,In_964,In_888);
nand U2488 (N_2488,In_800,In_2998);
nand U2489 (N_2489,In_1303,In_208);
nor U2490 (N_2490,In_2207,In_429);
nand U2491 (N_2491,In_262,In_2535);
nor U2492 (N_2492,In_2591,In_1989);
nor U2493 (N_2493,In_2780,In_622);
and U2494 (N_2494,In_1192,In_778);
and U2495 (N_2495,In_2933,In_221);
xor U2496 (N_2496,In_368,In_2591);
or U2497 (N_2497,In_439,In_2983);
nand U2498 (N_2498,In_1450,In_1098);
nand U2499 (N_2499,In_1612,In_1357);
and U2500 (N_2500,In_1277,In_530);
nor U2501 (N_2501,In_1467,In_538);
xor U2502 (N_2502,In_1440,In_499);
and U2503 (N_2503,In_508,In_1958);
nor U2504 (N_2504,In_259,In_2084);
xor U2505 (N_2505,In_628,In_2031);
nor U2506 (N_2506,In_1588,In_1476);
xnor U2507 (N_2507,In_2095,In_2340);
nor U2508 (N_2508,In_2394,In_1667);
xor U2509 (N_2509,In_2708,In_2508);
and U2510 (N_2510,In_1287,In_376);
xnor U2511 (N_2511,In_251,In_978);
xnor U2512 (N_2512,In_2869,In_1541);
xor U2513 (N_2513,In_2565,In_2881);
xor U2514 (N_2514,In_522,In_1660);
xnor U2515 (N_2515,In_1489,In_1989);
nand U2516 (N_2516,In_831,In_2628);
and U2517 (N_2517,In_1128,In_849);
nor U2518 (N_2518,In_2663,In_606);
nand U2519 (N_2519,In_130,In_421);
nor U2520 (N_2520,In_1846,In_2456);
and U2521 (N_2521,In_453,In_1909);
or U2522 (N_2522,In_289,In_2238);
and U2523 (N_2523,In_946,In_932);
xor U2524 (N_2524,In_772,In_90);
or U2525 (N_2525,In_916,In_208);
xnor U2526 (N_2526,In_2089,In_1513);
nor U2527 (N_2527,In_2970,In_2216);
and U2528 (N_2528,In_256,In_2638);
nor U2529 (N_2529,In_2613,In_171);
and U2530 (N_2530,In_2307,In_1294);
and U2531 (N_2531,In_2098,In_2847);
and U2532 (N_2532,In_746,In_316);
nor U2533 (N_2533,In_2853,In_2318);
nand U2534 (N_2534,In_2114,In_2739);
nand U2535 (N_2535,In_2766,In_2275);
nand U2536 (N_2536,In_767,In_2768);
nor U2537 (N_2537,In_2472,In_2195);
nand U2538 (N_2538,In_2376,In_1995);
nand U2539 (N_2539,In_425,In_2196);
nand U2540 (N_2540,In_2578,In_611);
and U2541 (N_2541,In_2123,In_1337);
and U2542 (N_2542,In_1022,In_569);
nor U2543 (N_2543,In_2862,In_1060);
xor U2544 (N_2544,In_1192,In_1233);
nor U2545 (N_2545,In_1744,In_1595);
and U2546 (N_2546,In_1523,In_585);
nor U2547 (N_2547,In_673,In_1477);
nor U2548 (N_2548,In_2693,In_2175);
and U2549 (N_2549,In_552,In_2287);
nand U2550 (N_2550,In_2009,In_1931);
nor U2551 (N_2551,In_2905,In_1467);
nand U2552 (N_2552,In_267,In_1128);
xnor U2553 (N_2553,In_2439,In_788);
nor U2554 (N_2554,In_608,In_1791);
and U2555 (N_2555,In_1989,In_1864);
or U2556 (N_2556,In_2487,In_1650);
nand U2557 (N_2557,In_1116,In_1129);
nor U2558 (N_2558,In_1503,In_1088);
nand U2559 (N_2559,In_1367,In_808);
nor U2560 (N_2560,In_134,In_2844);
and U2561 (N_2561,In_48,In_2034);
or U2562 (N_2562,In_2628,In_2013);
nand U2563 (N_2563,In_1706,In_2164);
or U2564 (N_2564,In_1015,In_2839);
and U2565 (N_2565,In_2097,In_2407);
nand U2566 (N_2566,In_353,In_563);
xnor U2567 (N_2567,In_7,In_2507);
nor U2568 (N_2568,In_2920,In_1167);
or U2569 (N_2569,In_1064,In_104);
or U2570 (N_2570,In_2056,In_1212);
or U2571 (N_2571,In_411,In_2504);
nor U2572 (N_2572,In_2012,In_1169);
and U2573 (N_2573,In_676,In_2615);
nand U2574 (N_2574,In_1993,In_2890);
xor U2575 (N_2575,In_847,In_278);
xnor U2576 (N_2576,In_1565,In_2037);
xor U2577 (N_2577,In_1393,In_2468);
nor U2578 (N_2578,In_198,In_1054);
nor U2579 (N_2579,In_869,In_1093);
nand U2580 (N_2580,In_1023,In_5);
or U2581 (N_2581,In_1048,In_1619);
nand U2582 (N_2582,In_1784,In_1010);
nand U2583 (N_2583,In_110,In_1610);
xor U2584 (N_2584,In_2729,In_1061);
and U2585 (N_2585,In_2589,In_668);
or U2586 (N_2586,In_972,In_158);
and U2587 (N_2587,In_1845,In_1742);
nand U2588 (N_2588,In_281,In_2845);
and U2589 (N_2589,In_2884,In_1773);
and U2590 (N_2590,In_2840,In_1037);
or U2591 (N_2591,In_693,In_1546);
and U2592 (N_2592,In_1114,In_2635);
nand U2593 (N_2593,In_1145,In_1482);
or U2594 (N_2594,In_1514,In_1022);
nand U2595 (N_2595,In_577,In_528);
nand U2596 (N_2596,In_269,In_789);
or U2597 (N_2597,In_537,In_2223);
and U2598 (N_2598,In_555,In_375);
and U2599 (N_2599,In_343,In_499);
or U2600 (N_2600,In_2678,In_1006);
nand U2601 (N_2601,In_657,In_2391);
or U2602 (N_2602,In_1427,In_1565);
nor U2603 (N_2603,In_1616,In_833);
nor U2604 (N_2604,In_2197,In_2274);
or U2605 (N_2605,In_549,In_463);
xnor U2606 (N_2606,In_2468,In_2117);
nand U2607 (N_2607,In_421,In_351);
nor U2608 (N_2608,In_2861,In_2665);
xnor U2609 (N_2609,In_1316,In_357);
xor U2610 (N_2610,In_1546,In_2089);
nor U2611 (N_2611,In_269,In_1342);
and U2612 (N_2612,In_1129,In_1333);
and U2613 (N_2613,In_2172,In_1868);
nand U2614 (N_2614,In_2769,In_1234);
nor U2615 (N_2615,In_1528,In_1551);
nand U2616 (N_2616,In_1317,In_2388);
or U2617 (N_2617,In_2468,In_276);
nor U2618 (N_2618,In_2552,In_2480);
and U2619 (N_2619,In_1132,In_2090);
nand U2620 (N_2620,In_1662,In_2102);
xnor U2621 (N_2621,In_1439,In_2533);
nor U2622 (N_2622,In_522,In_1518);
and U2623 (N_2623,In_1293,In_2631);
nor U2624 (N_2624,In_162,In_2783);
xnor U2625 (N_2625,In_1800,In_1996);
nand U2626 (N_2626,In_1595,In_12);
xor U2627 (N_2627,In_828,In_1559);
and U2628 (N_2628,In_1597,In_2396);
nand U2629 (N_2629,In_2300,In_1852);
nand U2630 (N_2630,In_992,In_2617);
nand U2631 (N_2631,In_1483,In_2865);
or U2632 (N_2632,In_830,In_282);
xnor U2633 (N_2633,In_1602,In_60);
nand U2634 (N_2634,In_92,In_810);
nand U2635 (N_2635,In_2387,In_488);
xnor U2636 (N_2636,In_2997,In_479);
xor U2637 (N_2637,In_518,In_1914);
and U2638 (N_2638,In_2821,In_209);
xor U2639 (N_2639,In_1604,In_1555);
nand U2640 (N_2640,In_696,In_2669);
nand U2641 (N_2641,In_2348,In_1787);
or U2642 (N_2642,In_450,In_2540);
nand U2643 (N_2643,In_1214,In_2903);
nand U2644 (N_2644,In_2970,In_2367);
nor U2645 (N_2645,In_914,In_1274);
and U2646 (N_2646,In_3,In_1825);
or U2647 (N_2647,In_2090,In_2640);
and U2648 (N_2648,In_1270,In_1221);
xnor U2649 (N_2649,In_1922,In_2833);
and U2650 (N_2650,In_759,In_2187);
or U2651 (N_2651,In_807,In_1355);
xor U2652 (N_2652,In_2882,In_1386);
and U2653 (N_2653,In_310,In_1584);
nand U2654 (N_2654,In_1376,In_1091);
nor U2655 (N_2655,In_2628,In_2248);
and U2656 (N_2656,In_1086,In_2911);
nand U2657 (N_2657,In_283,In_877);
nor U2658 (N_2658,In_2511,In_1572);
xnor U2659 (N_2659,In_293,In_352);
or U2660 (N_2660,In_2256,In_504);
nand U2661 (N_2661,In_1245,In_369);
and U2662 (N_2662,In_406,In_1887);
xnor U2663 (N_2663,In_2275,In_1021);
or U2664 (N_2664,In_879,In_1049);
xor U2665 (N_2665,In_1698,In_2263);
nor U2666 (N_2666,In_884,In_2298);
and U2667 (N_2667,In_2742,In_944);
or U2668 (N_2668,In_2190,In_553);
xor U2669 (N_2669,In_2824,In_1811);
and U2670 (N_2670,In_1286,In_706);
nand U2671 (N_2671,In_2766,In_2591);
xnor U2672 (N_2672,In_62,In_443);
and U2673 (N_2673,In_2723,In_2971);
or U2674 (N_2674,In_1920,In_322);
xor U2675 (N_2675,In_2797,In_1582);
xnor U2676 (N_2676,In_1193,In_2086);
and U2677 (N_2677,In_805,In_283);
xnor U2678 (N_2678,In_2166,In_762);
nor U2679 (N_2679,In_1646,In_2299);
and U2680 (N_2680,In_788,In_301);
nand U2681 (N_2681,In_1029,In_315);
or U2682 (N_2682,In_2607,In_2075);
or U2683 (N_2683,In_2957,In_649);
and U2684 (N_2684,In_756,In_2400);
and U2685 (N_2685,In_463,In_487);
or U2686 (N_2686,In_1051,In_1083);
nor U2687 (N_2687,In_2428,In_2937);
and U2688 (N_2688,In_2301,In_2484);
and U2689 (N_2689,In_2473,In_2465);
or U2690 (N_2690,In_1249,In_2551);
and U2691 (N_2691,In_135,In_2211);
nand U2692 (N_2692,In_85,In_2677);
nand U2693 (N_2693,In_1266,In_789);
nor U2694 (N_2694,In_697,In_1017);
xor U2695 (N_2695,In_2487,In_1311);
nand U2696 (N_2696,In_2279,In_1198);
and U2697 (N_2697,In_1447,In_1322);
or U2698 (N_2698,In_2173,In_2151);
and U2699 (N_2699,In_1940,In_2162);
nor U2700 (N_2700,In_2353,In_1714);
or U2701 (N_2701,In_2289,In_2283);
or U2702 (N_2702,In_2953,In_2384);
or U2703 (N_2703,In_8,In_2843);
xnor U2704 (N_2704,In_2493,In_1444);
and U2705 (N_2705,In_471,In_236);
nand U2706 (N_2706,In_1122,In_613);
nand U2707 (N_2707,In_1503,In_2140);
nor U2708 (N_2708,In_1235,In_842);
and U2709 (N_2709,In_789,In_1093);
or U2710 (N_2710,In_218,In_1356);
or U2711 (N_2711,In_846,In_129);
nand U2712 (N_2712,In_1617,In_2813);
xor U2713 (N_2713,In_1672,In_371);
and U2714 (N_2714,In_1191,In_1460);
nand U2715 (N_2715,In_872,In_783);
nor U2716 (N_2716,In_152,In_364);
nor U2717 (N_2717,In_1892,In_652);
and U2718 (N_2718,In_15,In_2648);
nor U2719 (N_2719,In_689,In_114);
nor U2720 (N_2720,In_509,In_1052);
nand U2721 (N_2721,In_966,In_2607);
and U2722 (N_2722,In_2232,In_2608);
and U2723 (N_2723,In_2938,In_1600);
xor U2724 (N_2724,In_293,In_1533);
or U2725 (N_2725,In_2872,In_1523);
nand U2726 (N_2726,In_1336,In_1233);
or U2727 (N_2727,In_522,In_1958);
and U2728 (N_2728,In_1764,In_512);
nand U2729 (N_2729,In_2824,In_993);
nand U2730 (N_2730,In_2297,In_77);
and U2731 (N_2731,In_560,In_667);
nor U2732 (N_2732,In_1062,In_2761);
and U2733 (N_2733,In_2365,In_1982);
nor U2734 (N_2734,In_1939,In_8);
nand U2735 (N_2735,In_2250,In_83);
and U2736 (N_2736,In_1599,In_166);
xor U2737 (N_2737,In_943,In_2239);
and U2738 (N_2738,In_689,In_1849);
xor U2739 (N_2739,In_461,In_2414);
xnor U2740 (N_2740,In_1603,In_2969);
nor U2741 (N_2741,In_406,In_1617);
nor U2742 (N_2742,In_369,In_737);
and U2743 (N_2743,In_380,In_2435);
and U2744 (N_2744,In_1681,In_493);
nand U2745 (N_2745,In_235,In_1571);
xnor U2746 (N_2746,In_2505,In_1639);
nand U2747 (N_2747,In_382,In_1067);
xor U2748 (N_2748,In_2985,In_1519);
nand U2749 (N_2749,In_139,In_1747);
xor U2750 (N_2750,In_1499,In_1449);
and U2751 (N_2751,In_2286,In_263);
and U2752 (N_2752,In_600,In_1422);
nor U2753 (N_2753,In_1320,In_1697);
or U2754 (N_2754,In_1898,In_1182);
nand U2755 (N_2755,In_2938,In_2040);
or U2756 (N_2756,In_2229,In_1958);
xnor U2757 (N_2757,In_1536,In_199);
and U2758 (N_2758,In_622,In_1533);
xor U2759 (N_2759,In_1353,In_529);
nand U2760 (N_2760,In_1461,In_1330);
or U2761 (N_2761,In_2764,In_2974);
or U2762 (N_2762,In_2518,In_1212);
nor U2763 (N_2763,In_2356,In_2085);
nor U2764 (N_2764,In_1114,In_1590);
nand U2765 (N_2765,In_59,In_1701);
and U2766 (N_2766,In_1460,In_2983);
nand U2767 (N_2767,In_648,In_1626);
xor U2768 (N_2768,In_1256,In_635);
nand U2769 (N_2769,In_518,In_1631);
nand U2770 (N_2770,In_1659,In_1210);
nor U2771 (N_2771,In_1798,In_2611);
xnor U2772 (N_2772,In_161,In_1263);
and U2773 (N_2773,In_108,In_1672);
nand U2774 (N_2774,In_97,In_693);
and U2775 (N_2775,In_819,In_2469);
and U2776 (N_2776,In_2841,In_2013);
xor U2777 (N_2777,In_2103,In_2387);
xnor U2778 (N_2778,In_2127,In_2037);
nor U2779 (N_2779,In_727,In_184);
nand U2780 (N_2780,In_2664,In_2576);
nand U2781 (N_2781,In_2241,In_1485);
xnor U2782 (N_2782,In_2454,In_1479);
nor U2783 (N_2783,In_392,In_920);
nand U2784 (N_2784,In_1878,In_2341);
nor U2785 (N_2785,In_1561,In_2872);
or U2786 (N_2786,In_2981,In_1124);
and U2787 (N_2787,In_541,In_921);
or U2788 (N_2788,In_2463,In_1773);
nand U2789 (N_2789,In_2379,In_906);
and U2790 (N_2790,In_861,In_810);
nand U2791 (N_2791,In_773,In_682);
nor U2792 (N_2792,In_2811,In_650);
nor U2793 (N_2793,In_694,In_1137);
nand U2794 (N_2794,In_904,In_359);
xnor U2795 (N_2795,In_433,In_811);
xor U2796 (N_2796,In_1936,In_2088);
nand U2797 (N_2797,In_2089,In_161);
or U2798 (N_2798,In_1721,In_323);
nand U2799 (N_2799,In_756,In_2437);
or U2800 (N_2800,In_1626,In_191);
or U2801 (N_2801,In_1655,In_1018);
xor U2802 (N_2802,In_491,In_2853);
xnor U2803 (N_2803,In_183,In_614);
nor U2804 (N_2804,In_1973,In_753);
nor U2805 (N_2805,In_1672,In_1323);
or U2806 (N_2806,In_2409,In_678);
and U2807 (N_2807,In_1725,In_821);
nand U2808 (N_2808,In_1007,In_1546);
xor U2809 (N_2809,In_398,In_2641);
and U2810 (N_2810,In_2305,In_310);
nor U2811 (N_2811,In_1935,In_1875);
and U2812 (N_2812,In_648,In_959);
and U2813 (N_2813,In_1279,In_2799);
and U2814 (N_2814,In_1348,In_807);
nor U2815 (N_2815,In_1651,In_514);
and U2816 (N_2816,In_180,In_1599);
and U2817 (N_2817,In_1032,In_1980);
nor U2818 (N_2818,In_1072,In_670);
nand U2819 (N_2819,In_2837,In_1045);
nor U2820 (N_2820,In_517,In_937);
or U2821 (N_2821,In_1145,In_811);
nand U2822 (N_2822,In_1594,In_810);
or U2823 (N_2823,In_2157,In_2600);
nand U2824 (N_2824,In_754,In_2294);
nand U2825 (N_2825,In_2559,In_780);
xor U2826 (N_2826,In_2381,In_2583);
xnor U2827 (N_2827,In_2959,In_1288);
and U2828 (N_2828,In_501,In_1040);
nand U2829 (N_2829,In_2662,In_2937);
nor U2830 (N_2830,In_1305,In_1465);
xnor U2831 (N_2831,In_872,In_1967);
nand U2832 (N_2832,In_1202,In_2307);
nor U2833 (N_2833,In_1818,In_2141);
and U2834 (N_2834,In_421,In_2307);
nor U2835 (N_2835,In_510,In_1499);
xnor U2836 (N_2836,In_565,In_2122);
xor U2837 (N_2837,In_2787,In_1742);
nand U2838 (N_2838,In_901,In_2662);
nor U2839 (N_2839,In_716,In_573);
nand U2840 (N_2840,In_2023,In_1331);
and U2841 (N_2841,In_2747,In_1878);
or U2842 (N_2842,In_2885,In_80);
and U2843 (N_2843,In_114,In_2317);
or U2844 (N_2844,In_1183,In_428);
or U2845 (N_2845,In_245,In_1816);
xor U2846 (N_2846,In_2653,In_1014);
nor U2847 (N_2847,In_1280,In_2599);
xor U2848 (N_2848,In_1172,In_1682);
nand U2849 (N_2849,In_328,In_2998);
xnor U2850 (N_2850,In_2982,In_2874);
or U2851 (N_2851,In_2680,In_901);
and U2852 (N_2852,In_613,In_981);
and U2853 (N_2853,In_664,In_2199);
xor U2854 (N_2854,In_1760,In_2037);
and U2855 (N_2855,In_702,In_268);
nor U2856 (N_2856,In_2472,In_1838);
xnor U2857 (N_2857,In_1291,In_6);
or U2858 (N_2858,In_1809,In_2607);
nor U2859 (N_2859,In_1528,In_1748);
and U2860 (N_2860,In_435,In_539);
xnor U2861 (N_2861,In_110,In_970);
and U2862 (N_2862,In_2531,In_1122);
nor U2863 (N_2863,In_893,In_2146);
nor U2864 (N_2864,In_785,In_245);
nor U2865 (N_2865,In_1804,In_2968);
nand U2866 (N_2866,In_370,In_384);
or U2867 (N_2867,In_1314,In_2910);
nand U2868 (N_2868,In_1196,In_1611);
or U2869 (N_2869,In_1563,In_388);
nor U2870 (N_2870,In_252,In_1523);
or U2871 (N_2871,In_131,In_1839);
nor U2872 (N_2872,In_2567,In_544);
xor U2873 (N_2873,In_83,In_2556);
nand U2874 (N_2874,In_128,In_514);
or U2875 (N_2875,In_1533,In_2847);
xor U2876 (N_2876,In_467,In_1090);
and U2877 (N_2877,In_2660,In_1600);
nand U2878 (N_2878,In_1599,In_2625);
or U2879 (N_2879,In_1149,In_2233);
or U2880 (N_2880,In_981,In_1403);
xnor U2881 (N_2881,In_1756,In_1386);
xnor U2882 (N_2882,In_2366,In_1404);
and U2883 (N_2883,In_1429,In_2885);
nor U2884 (N_2884,In_2611,In_279);
nand U2885 (N_2885,In_1825,In_1118);
nor U2886 (N_2886,In_875,In_1008);
or U2887 (N_2887,In_1661,In_1475);
xnor U2888 (N_2888,In_2435,In_2199);
nand U2889 (N_2889,In_1493,In_313);
and U2890 (N_2890,In_1463,In_50);
and U2891 (N_2891,In_1023,In_1563);
or U2892 (N_2892,In_541,In_1479);
or U2893 (N_2893,In_1940,In_386);
xor U2894 (N_2894,In_1857,In_1975);
xor U2895 (N_2895,In_2585,In_612);
and U2896 (N_2896,In_788,In_1486);
and U2897 (N_2897,In_500,In_2278);
nand U2898 (N_2898,In_2997,In_2065);
xnor U2899 (N_2899,In_2514,In_2344);
nor U2900 (N_2900,In_638,In_2348);
and U2901 (N_2901,In_1298,In_1233);
nor U2902 (N_2902,In_2861,In_1312);
and U2903 (N_2903,In_1734,In_1898);
xnor U2904 (N_2904,In_2292,In_2787);
and U2905 (N_2905,In_1227,In_1207);
nand U2906 (N_2906,In_640,In_678);
nor U2907 (N_2907,In_1469,In_755);
nand U2908 (N_2908,In_286,In_2856);
xor U2909 (N_2909,In_936,In_2077);
nand U2910 (N_2910,In_2537,In_248);
nor U2911 (N_2911,In_1569,In_52);
and U2912 (N_2912,In_254,In_1268);
xor U2913 (N_2913,In_246,In_1301);
or U2914 (N_2914,In_1067,In_2462);
xor U2915 (N_2915,In_2799,In_905);
and U2916 (N_2916,In_949,In_2452);
nand U2917 (N_2917,In_810,In_1764);
or U2918 (N_2918,In_1090,In_367);
xor U2919 (N_2919,In_370,In_1926);
xor U2920 (N_2920,In_2250,In_2390);
xor U2921 (N_2921,In_301,In_1236);
or U2922 (N_2922,In_1442,In_725);
nand U2923 (N_2923,In_2309,In_331);
nand U2924 (N_2924,In_2807,In_1675);
nor U2925 (N_2925,In_2173,In_415);
xor U2926 (N_2926,In_1773,In_136);
nand U2927 (N_2927,In_2005,In_2470);
and U2928 (N_2928,In_2938,In_259);
nor U2929 (N_2929,In_1785,In_1381);
nor U2930 (N_2930,In_1428,In_2093);
and U2931 (N_2931,In_955,In_2094);
or U2932 (N_2932,In_2086,In_2973);
nor U2933 (N_2933,In_2998,In_2085);
nor U2934 (N_2934,In_1954,In_731);
xnor U2935 (N_2935,In_2994,In_2377);
or U2936 (N_2936,In_341,In_2832);
nand U2937 (N_2937,In_2879,In_1197);
or U2938 (N_2938,In_626,In_2290);
nand U2939 (N_2939,In_1529,In_2005);
and U2940 (N_2940,In_1675,In_2865);
or U2941 (N_2941,In_1210,In_26);
nand U2942 (N_2942,In_1520,In_1899);
xnor U2943 (N_2943,In_2708,In_2967);
nor U2944 (N_2944,In_648,In_1629);
and U2945 (N_2945,In_1217,In_2118);
nand U2946 (N_2946,In_604,In_706);
nand U2947 (N_2947,In_2814,In_1539);
and U2948 (N_2948,In_2463,In_589);
nor U2949 (N_2949,In_947,In_1224);
or U2950 (N_2950,In_1486,In_2314);
xnor U2951 (N_2951,In_1878,In_2648);
xnor U2952 (N_2952,In_1546,In_1830);
nand U2953 (N_2953,In_2568,In_193);
and U2954 (N_2954,In_2348,In_1572);
nor U2955 (N_2955,In_2317,In_656);
nor U2956 (N_2956,In_2790,In_2103);
and U2957 (N_2957,In_2717,In_133);
nand U2958 (N_2958,In_2877,In_509);
xor U2959 (N_2959,In_2519,In_115);
xnor U2960 (N_2960,In_2185,In_862);
nor U2961 (N_2961,In_824,In_2942);
nor U2962 (N_2962,In_43,In_2050);
or U2963 (N_2963,In_2900,In_1664);
nor U2964 (N_2964,In_258,In_2462);
or U2965 (N_2965,In_34,In_2077);
nand U2966 (N_2966,In_2387,In_645);
nor U2967 (N_2967,In_74,In_554);
nor U2968 (N_2968,In_1493,In_2244);
or U2969 (N_2969,In_1413,In_1315);
or U2970 (N_2970,In_2210,In_2515);
nor U2971 (N_2971,In_695,In_789);
and U2972 (N_2972,In_301,In_1518);
nand U2973 (N_2973,In_2988,In_822);
or U2974 (N_2974,In_1790,In_2988);
xor U2975 (N_2975,In_2236,In_2402);
or U2976 (N_2976,In_877,In_427);
nor U2977 (N_2977,In_1892,In_185);
and U2978 (N_2978,In_1530,In_111);
xnor U2979 (N_2979,In_654,In_1527);
or U2980 (N_2980,In_341,In_2520);
or U2981 (N_2981,In_834,In_1827);
or U2982 (N_2982,In_1619,In_1342);
nand U2983 (N_2983,In_82,In_915);
xnor U2984 (N_2984,In_1900,In_754);
or U2985 (N_2985,In_710,In_1677);
nand U2986 (N_2986,In_1852,In_692);
nor U2987 (N_2987,In_1620,In_507);
nor U2988 (N_2988,In_1808,In_1371);
nand U2989 (N_2989,In_1623,In_1461);
nor U2990 (N_2990,In_2637,In_2827);
nor U2991 (N_2991,In_2695,In_2289);
and U2992 (N_2992,In_301,In_107);
nor U2993 (N_2993,In_2729,In_1237);
and U2994 (N_2994,In_1280,In_1954);
and U2995 (N_2995,In_768,In_1690);
xnor U2996 (N_2996,In_2831,In_711);
xor U2997 (N_2997,In_1812,In_271);
and U2998 (N_2998,In_667,In_108);
nor U2999 (N_2999,In_1254,In_351);
xnor U3000 (N_3000,In_2795,In_284);
nor U3001 (N_3001,In_2425,In_911);
and U3002 (N_3002,In_132,In_2508);
nand U3003 (N_3003,In_1234,In_195);
nand U3004 (N_3004,In_2419,In_2822);
nand U3005 (N_3005,In_1925,In_2170);
or U3006 (N_3006,In_1241,In_1811);
and U3007 (N_3007,In_168,In_2491);
nand U3008 (N_3008,In_690,In_1);
nor U3009 (N_3009,In_868,In_902);
nor U3010 (N_3010,In_622,In_574);
nor U3011 (N_3011,In_467,In_406);
nand U3012 (N_3012,In_1752,In_325);
xor U3013 (N_3013,In_1551,In_682);
xnor U3014 (N_3014,In_1721,In_847);
and U3015 (N_3015,In_2688,In_1009);
nor U3016 (N_3016,In_884,In_1324);
nand U3017 (N_3017,In_2667,In_1973);
or U3018 (N_3018,In_2125,In_2097);
xor U3019 (N_3019,In_998,In_514);
xnor U3020 (N_3020,In_1915,In_2541);
nand U3021 (N_3021,In_2108,In_2920);
or U3022 (N_3022,In_2454,In_1276);
nor U3023 (N_3023,In_838,In_2667);
nand U3024 (N_3024,In_1474,In_2689);
or U3025 (N_3025,In_1269,In_2835);
or U3026 (N_3026,In_2803,In_2201);
xor U3027 (N_3027,In_2775,In_2375);
nand U3028 (N_3028,In_2234,In_1241);
nand U3029 (N_3029,In_2866,In_2473);
xnor U3030 (N_3030,In_1357,In_1255);
xnor U3031 (N_3031,In_2300,In_2169);
and U3032 (N_3032,In_2615,In_807);
and U3033 (N_3033,In_2163,In_606);
and U3034 (N_3034,In_270,In_1202);
nand U3035 (N_3035,In_1534,In_2190);
and U3036 (N_3036,In_2902,In_653);
xnor U3037 (N_3037,In_1470,In_811);
or U3038 (N_3038,In_1362,In_624);
xor U3039 (N_3039,In_132,In_30);
nor U3040 (N_3040,In_612,In_1017);
and U3041 (N_3041,In_1232,In_2185);
nor U3042 (N_3042,In_1600,In_826);
and U3043 (N_3043,In_628,In_889);
nand U3044 (N_3044,In_2719,In_1862);
xnor U3045 (N_3045,In_2294,In_508);
or U3046 (N_3046,In_2398,In_1548);
nand U3047 (N_3047,In_2277,In_2106);
or U3048 (N_3048,In_1520,In_2721);
nor U3049 (N_3049,In_2691,In_283);
nand U3050 (N_3050,In_2157,In_181);
xor U3051 (N_3051,In_1040,In_349);
nand U3052 (N_3052,In_2780,In_416);
nand U3053 (N_3053,In_2760,In_444);
or U3054 (N_3054,In_1195,In_1869);
xor U3055 (N_3055,In_2203,In_20);
nor U3056 (N_3056,In_982,In_1548);
and U3057 (N_3057,In_171,In_1475);
or U3058 (N_3058,In_66,In_159);
nand U3059 (N_3059,In_2133,In_2800);
nand U3060 (N_3060,In_2820,In_1541);
or U3061 (N_3061,In_317,In_1955);
nand U3062 (N_3062,In_2836,In_1938);
nand U3063 (N_3063,In_1901,In_1249);
and U3064 (N_3064,In_222,In_2641);
or U3065 (N_3065,In_2585,In_760);
or U3066 (N_3066,In_2540,In_2717);
and U3067 (N_3067,In_2895,In_1901);
nand U3068 (N_3068,In_1106,In_1323);
and U3069 (N_3069,In_982,In_2408);
or U3070 (N_3070,In_1956,In_2466);
nand U3071 (N_3071,In_613,In_603);
nand U3072 (N_3072,In_825,In_1275);
xor U3073 (N_3073,In_1723,In_2983);
or U3074 (N_3074,In_2351,In_2703);
xor U3075 (N_3075,In_876,In_2468);
or U3076 (N_3076,In_682,In_1564);
nor U3077 (N_3077,In_664,In_548);
nand U3078 (N_3078,In_1920,In_1836);
nor U3079 (N_3079,In_10,In_1593);
nand U3080 (N_3080,In_1266,In_1035);
nor U3081 (N_3081,In_2091,In_1258);
xor U3082 (N_3082,In_2532,In_1750);
or U3083 (N_3083,In_945,In_2927);
and U3084 (N_3084,In_624,In_2015);
xnor U3085 (N_3085,In_2313,In_256);
xnor U3086 (N_3086,In_800,In_758);
nor U3087 (N_3087,In_1286,In_702);
nor U3088 (N_3088,In_396,In_2149);
and U3089 (N_3089,In_140,In_2078);
nor U3090 (N_3090,In_411,In_1329);
nor U3091 (N_3091,In_2044,In_1009);
and U3092 (N_3092,In_1172,In_1825);
nor U3093 (N_3093,In_1663,In_880);
xnor U3094 (N_3094,In_2774,In_283);
or U3095 (N_3095,In_460,In_259);
nor U3096 (N_3096,In_1751,In_2234);
nand U3097 (N_3097,In_416,In_1928);
xnor U3098 (N_3098,In_1393,In_1763);
nand U3099 (N_3099,In_2643,In_1160);
or U3100 (N_3100,In_1917,In_817);
nor U3101 (N_3101,In_2157,In_1567);
nor U3102 (N_3102,In_962,In_1067);
xor U3103 (N_3103,In_1060,In_1620);
xor U3104 (N_3104,In_549,In_1544);
xnor U3105 (N_3105,In_992,In_447);
nand U3106 (N_3106,In_1488,In_1736);
xnor U3107 (N_3107,In_2122,In_105);
and U3108 (N_3108,In_1736,In_1568);
and U3109 (N_3109,In_1858,In_889);
nor U3110 (N_3110,In_1092,In_362);
and U3111 (N_3111,In_2467,In_1772);
nand U3112 (N_3112,In_701,In_1748);
nand U3113 (N_3113,In_2360,In_362);
nor U3114 (N_3114,In_845,In_467);
nand U3115 (N_3115,In_2987,In_2439);
or U3116 (N_3116,In_2149,In_1622);
nand U3117 (N_3117,In_59,In_1822);
and U3118 (N_3118,In_1381,In_771);
and U3119 (N_3119,In_1083,In_2812);
nand U3120 (N_3120,In_1808,In_2319);
or U3121 (N_3121,In_983,In_1503);
and U3122 (N_3122,In_788,In_2029);
xor U3123 (N_3123,In_1537,In_2287);
xor U3124 (N_3124,In_1041,In_2486);
or U3125 (N_3125,In_1873,In_335);
nand U3126 (N_3126,In_1120,In_2362);
and U3127 (N_3127,In_1907,In_130);
xnor U3128 (N_3128,In_2852,In_1097);
or U3129 (N_3129,In_1306,In_2551);
or U3130 (N_3130,In_1385,In_513);
or U3131 (N_3131,In_693,In_707);
nor U3132 (N_3132,In_1419,In_2681);
or U3133 (N_3133,In_1750,In_2808);
and U3134 (N_3134,In_1992,In_1194);
and U3135 (N_3135,In_1010,In_1203);
or U3136 (N_3136,In_403,In_1622);
or U3137 (N_3137,In_2655,In_1512);
nand U3138 (N_3138,In_2477,In_2859);
nor U3139 (N_3139,In_2102,In_959);
nand U3140 (N_3140,In_2291,In_1098);
nor U3141 (N_3141,In_1022,In_1250);
and U3142 (N_3142,In_2862,In_745);
xor U3143 (N_3143,In_2017,In_447);
xor U3144 (N_3144,In_1950,In_2601);
xor U3145 (N_3145,In_445,In_802);
and U3146 (N_3146,In_2315,In_1969);
xnor U3147 (N_3147,In_1875,In_847);
or U3148 (N_3148,In_2296,In_1226);
nand U3149 (N_3149,In_2722,In_546);
nand U3150 (N_3150,In_1642,In_1472);
xnor U3151 (N_3151,In_2987,In_2401);
and U3152 (N_3152,In_2460,In_93);
nand U3153 (N_3153,In_341,In_2595);
nand U3154 (N_3154,In_175,In_2376);
or U3155 (N_3155,In_2041,In_2524);
or U3156 (N_3156,In_2007,In_647);
nor U3157 (N_3157,In_463,In_1000);
nand U3158 (N_3158,In_1541,In_639);
and U3159 (N_3159,In_2094,In_2376);
xor U3160 (N_3160,In_1890,In_128);
xnor U3161 (N_3161,In_766,In_2163);
or U3162 (N_3162,In_1216,In_1354);
and U3163 (N_3163,In_1397,In_604);
nand U3164 (N_3164,In_1025,In_187);
xor U3165 (N_3165,In_2609,In_1389);
or U3166 (N_3166,In_2474,In_2455);
nand U3167 (N_3167,In_1470,In_886);
nand U3168 (N_3168,In_1830,In_2124);
xnor U3169 (N_3169,In_1220,In_628);
or U3170 (N_3170,In_459,In_1905);
and U3171 (N_3171,In_1159,In_1820);
and U3172 (N_3172,In_113,In_950);
nor U3173 (N_3173,In_1654,In_643);
nor U3174 (N_3174,In_2315,In_1442);
and U3175 (N_3175,In_656,In_1162);
xor U3176 (N_3176,In_1656,In_1893);
or U3177 (N_3177,In_4,In_1600);
xnor U3178 (N_3178,In_1854,In_2385);
nand U3179 (N_3179,In_455,In_2482);
or U3180 (N_3180,In_2421,In_1405);
xnor U3181 (N_3181,In_2463,In_910);
nand U3182 (N_3182,In_546,In_2104);
nand U3183 (N_3183,In_1963,In_2180);
nor U3184 (N_3184,In_1755,In_1178);
and U3185 (N_3185,In_742,In_526);
nor U3186 (N_3186,In_2682,In_2349);
nor U3187 (N_3187,In_130,In_2146);
and U3188 (N_3188,In_1044,In_1351);
nand U3189 (N_3189,In_1296,In_503);
and U3190 (N_3190,In_1572,In_1264);
and U3191 (N_3191,In_416,In_1048);
nand U3192 (N_3192,In_1826,In_2827);
and U3193 (N_3193,In_1944,In_2577);
xor U3194 (N_3194,In_1432,In_2397);
and U3195 (N_3195,In_2135,In_2692);
and U3196 (N_3196,In_502,In_1060);
nand U3197 (N_3197,In_2717,In_2707);
nand U3198 (N_3198,In_1503,In_813);
nor U3199 (N_3199,In_260,In_2399);
and U3200 (N_3200,In_970,In_1109);
nand U3201 (N_3201,In_2811,In_1712);
nand U3202 (N_3202,In_1560,In_254);
nor U3203 (N_3203,In_556,In_1601);
nor U3204 (N_3204,In_2385,In_1187);
nand U3205 (N_3205,In_114,In_836);
xnor U3206 (N_3206,In_168,In_268);
and U3207 (N_3207,In_2119,In_360);
and U3208 (N_3208,In_1625,In_2051);
or U3209 (N_3209,In_566,In_289);
xnor U3210 (N_3210,In_748,In_901);
xor U3211 (N_3211,In_2440,In_2458);
nor U3212 (N_3212,In_472,In_2621);
nand U3213 (N_3213,In_165,In_2061);
or U3214 (N_3214,In_684,In_1735);
nor U3215 (N_3215,In_492,In_494);
nor U3216 (N_3216,In_1572,In_1907);
nand U3217 (N_3217,In_2860,In_2638);
nand U3218 (N_3218,In_555,In_1425);
nand U3219 (N_3219,In_2212,In_2167);
xor U3220 (N_3220,In_2061,In_2730);
xor U3221 (N_3221,In_655,In_1900);
and U3222 (N_3222,In_1934,In_2692);
nand U3223 (N_3223,In_1457,In_1115);
or U3224 (N_3224,In_1108,In_722);
and U3225 (N_3225,In_2523,In_2386);
and U3226 (N_3226,In_2464,In_545);
and U3227 (N_3227,In_722,In_1833);
xnor U3228 (N_3228,In_2478,In_2898);
nor U3229 (N_3229,In_1416,In_2584);
nand U3230 (N_3230,In_730,In_1145);
xnor U3231 (N_3231,In_593,In_983);
nand U3232 (N_3232,In_364,In_149);
nor U3233 (N_3233,In_2970,In_262);
nand U3234 (N_3234,In_2023,In_602);
nand U3235 (N_3235,In_2835,In_1956);
xnor U3236 (N_3236,In_1475,In_2227);
xor U3237 (N_3237,In_2687,In_2376);
nand U3238 (N_3238,In_1948,In_2300);
and U3239 (N_3239,In_1662,In_1602);
and U3240 (N_3240,In_1396,In_2041);
nand U3241 (N_3241,In_1194,In_2840);
nor U3242 (N_3242,In_89,In_1856);
and U3243 (N_3243,In_2475,In_2899);
or U3244 (N_3244,In_488,In_1188);
nand U3245 (N_3245,In_2765,In_2065);
and U3246 (N_3246,In_1431,In_1794);
or U3247 (N_3247,In_956,In_2985);
xor U3248 (N_3248,In_2194,In_2881);
and U3249 (N_3249,In_2637,In_2137);
nor U3250 (N_3250,In_1202,In_1503);
nand U3251 (N_3251,In_2939,In_1811);
or U3252 (N_3252,In_1141,In_2274);
nor U3253 (N_3253,In_988,In_1167);
nor U3254 (N_3254,In_990,In_23);
or U3255 (N_3255,In_1903,In_1466);
or U3256 (N_3256,In_2856,In_465);
nor U3257 (N_3257,In_2956,In_2552);
or U3258 (N_3258,In_1917,In_199);
and U3259 (N_3259,In_2329,In_845);
nand U3260 (N_3260,In_2872,In_1986);
nand U3261 (N_3261,In_160,In_361);
and U3262 (N_3262,In_1910,In_184);
nand U3263 (N_3263,In_340,In_1373);
and U3264 (N_3264,In_2457,In_1234);
and U3265 (N_3265,In_1034,In_1831);
xnor U3266 (N_3266,In_2580,In_320);
nand U3267 (N_3267,In_1906,In_806);
or U3268 (N_3268,In_1608,In_546);
xnor U3269 (N_3269,In_1541,In_1973);
and U3270 (N_3270,In_1990,In_2423);
nor U3271 (N_3271,In_2,In_2023);
nor U3272 (N_3272,In_623,In_2746);
and U3273 (N_3273,In_2949,In_245);
or U3274 (N_3274,In_2186,In_1672);
nor U3275 (N_3275,In_909,In_1628);
nand U3276 (N_3276,In_72,In_2033);
nand U3277 (N_3277,In_171,In_722);
xor U3278 (N_3278,In_2958,In_926);
nor U3279 (N_3279,In_290,In_2167);
nor U3280 (N_3280,In_928,In_1172);
nor U3281 (N_3281,In_2917,In_1793);
and U3282 (N_3282,In_2056,In_2581);
and U3283 (N_3283,In_2679,In_2771);
or U3284 (N_3284,In_2969,In_1074);
nand U3285 (N_3285,In_453,In_2545);
nor U3286 (N_3286,In_1990,In_2081);
or U3287 (N_3287,In_66,In_1340);
or U3288 (N_3288,In_1951,In_11);
or U3289 (N_3289,In_2652,In_2187);
nor U3290 (N_3290,In_2562,In_1178);
or U3291 (N_3291,In_2588,In_1249);
or U3292 (N_3292,In_947,In_1357);
nor U3293 (N_3293,In_224,In_2841);
xor U3294 (N_3294,In_969,In_2790);
nor U3295 (N_3295,In_1846,In_634);
nor U3296 (N_3296,In_2843,In_1219);
nor U3297 (N_3297,In_1992,In_1474);
or U3298 (N_3298,In_1015,In_1256);
nand U3299 (N_3299,In_1066,In_962);
xnor U3300 (N_3300,In_1039,In_639);
nand U3301 (N_3301,In_470,In_1731);
nor U3302 (N_3302,In_2786,In_2367);
and U3303 (N_3303,In_1933,In_2321);
nor U3304 (N_3304,In_778,In_1287);
and U3305 (N_3305,In_483,In_197);
nand U3306 (N_3306,In_196,In_921);
or U3307 (N_3307,In_670,In_2008);
or U3308 (N_3308,In_1086,In_326);
nand U3309 (N_3309,In_2669,In_423);
nand U3310 (N_3310,In_2209,In_1698);
nand U3311 (N_3311,In_2439,In_970);
xnor U3312 (N_3312,In_1070,In_986);
xnor U3313 (N_3313,In_1873,In_2220);
nand U3314 (N_3314,In_2795,In_459);
nor U3315 (N_3315,In_1681,In_307);
nand U3316 (N_3316,In_2631,In_1784);
or U3317 (N_3317,In_2478,In_1144);
and U3318 (N_3318,In_1444,In_2390);
and U3319 (N_3319,In_2864,In_989);
and U3320 (N_3320,In_267,In_2730);
or U3321 (N_3321,In_2062,In_2205);
and U3322 (N_3322,In_162,In_645);
nor U3323 (N_3323,In_23,In_1208);
and U3324 (N_3324,In_2498,In_2390);
nor U3325 (N_3325,In_993,In_248);
or U3326 (N_3326,In_1845,In_2623);
or U3327 (N_3327,In_967,In_1200);
and U3328 (N_3328,In_998,In_1606);
or U3329 (N_3329,In_709,In_620);
nand U3330 (N_3330,In_1744,In_2473);
or U3331 (N_3331,In_2753,In_1956);
or U3332 (N_3332,In_1134,In_2349);
nor U3333 (N_3333,In_188,In_728);
nand U3334 (N_3334,In_580,In_2238);
and U3335 (N_3335,In_2462,In_711);
and U3336 (N_3336,In_2933,In_446);
and U3337 (N_3337,In_1218,In_805);
or U3338 (N_3338,In_1248,In_925);
nand U3339 (N_3339,In_673,In_2766);
xnor U3340 (N_3340,In_882,In_752);
or U3341 (N_3341,In_1582,In_804);
xnor U3342 (N_3342,In_1998,In_1217);
nand U3343 (N_3343,In_1781,In_2914);
nor U3344 (N_3344,In_1006,In_1900);
xor U3345 (N_3345,In_1060,In_2525);
xnor U3346 (N_3346,In_2103,In_2536);
xnor U3347 (N_3347,In_295,In_2003);
xnor U3348 (N_3348,In_2056,In_2111);
nand U3349 (N_3349,In_792,In_695);
or U3350 (N_3350,In_1017,In_1755);
or U3351 (N_3351,In_2348,In_2371);
nor U3352 (N_3352,In_2629,In_1981);
and U3353 (N_3353,In_413,In_2714);
xor U3354 (N_3354,In_987,In_2055);
xor U3355 (N_3355,In_1240,In_2617);
xnor U3356 (N_3356,In_2423,In_1000);
or U3357 (N_3357,In_6,In_1517);
nand U3358 (N_3358,In_2971,In_2820);
or U3359 (N_3359,In_1710,In_862);
nand U3360 (N_3360,In_1986,In_2184);
xor U3361 (N_3361,In_2672,In_177);
nand U3362 (N_3362,In_916,In_141);
nor U3363 (N_3363,In_2694,In_2740);
and U3364 (N_3364,In_1366,In_386);
and U3365 (N_3365,In_1296,In_2003);
and U3366 (N_3366,In_59,In_2392);
nand U3367 (N_3367,In_1930,In_2668);
and U3368 (N_3368,In_2931,In_1511);
xnor U3369 (N_3369,In_1138,In_364);
or U3370 (N_3370,In_432,In_2737);
and U3371 (N_3371,In_1093,In_792);
xor U3372 (N_3372,In_1547,In_1560);
and U3373 (N_3373,In_2380,In_455);
and U3374 (N_3374,In_2329,In_2968);
nor U3375 (N_3375,In_2475,In_1692);
nor U3376 (N_3376,In_2758,In_672);
or U3377 (N_3377,In_2194,In_104);
xor U3378 (N_3378,In_268,In_234);
and U3379 (N_3379,In_1859,In_371);
xor U3380 (N_3380,In_2609,In_1947);
nor U3381 (N_3381,In_814,In_661);
xnor U3382 (N_3382,In_1415,In_1962);
nand U3383 (N_3383,In_1047,In_0);
and U3384 (N_3384,In_2953,In_656);
xor U3385 (N_3385,In_557,In_2634);
xor U3386 (N_3386,In_477,In_463);
nor U3387 (N_3387,In_2036,In_893);
xnor U3388 (N_3388,In_2778,In_941);
or U3389 (N_3389,In_2135,In_616);
xor U3390 (N_3390,In_2111,In_623);
and U3391 (N_3391,In_894,In_187);
xnor U3392 (N_3392,In_1996,In_914);
xnor U3393 (N_3393,In_838,In_1002);
nand U3394 (N_3394,In_201,In_1365);
and U3395 (N_3395,In_148,In_2775);
nor U3396 (N_3396,In_650,In_1118);
xnor U3397 (N_3397,In_298,In_64);
and U3398 (N_3398,In_2986,In_2249);
or U3399 (N_3399,In_2958,In_1467);
nand U3400 (N_3400,In_2731,In_1710);
nor U3401 (N_3401,In_2360,In_2371);
and U3402 (N_3402,In_205,In_2107);
nor U3403 (N_3403,In_417,In_408);
nor U3404 (N_3404,In_1144,In_1582);
xnor U3405 (N_3405,In_200,In_1385);
and U3406 (N_3406,In_1660,In_158);
or U3407 (N_3407,In_168,In_2888);
or U3408 (N_3408,In_1154,In_2607);
nand U3409 (N_3409,In_1973,In_2118);
xnor U3410 (N_3410,In_97,In_1568);
xnor U3411 (N_3411,In_316,In_1677);
or U3412 (N_3412,In_2905,In_239);
nand U3413 (N_3413,In_1564,In_2977);
nand U3414 (N_3414,In_221,In_952);
or U3415 (N_3415,In_1967,In_1209);
or U3416 (N_3416,In_2996,In_2483);
nor U3417 (N_3417,In_2701,In_1661);
nand U3418 (N_3418,In_2948,In_1183);
and U3419 (N_3419,In_465,In_1453);
nor U3420 (N_3420,In_1059,In_407);
and U3421 (N_3421,In_2222,In_2945);
nor U3422 (N_3422,In_1426,In_91);
nor U3423 (N_3423,In_1057,In_2974);
or U3424 (N_3424,In_1935,In_630);
nand U3425 (N_3425,In_2267,In_2183);
xor U3426 (N_3426,In_250,In_1139);
nor U3427 (N_3427,In_1578,In_2071);
xor U3428 (N_3428,In_1974,In_1083);
nand U3429 (N_3429,In_1521,In_393);
xor U3430 (N_3430,In_1818,In_391);
or U3431 (N_3431,In_2673,In_2411);
xnor U3432 (N_3432,In_1106,In_335);
nor U3433 (N_3433,In_1080,In_938);
or U3434 (N_3434,In_554,In_2153);
nor U3435 (N_3435,In_2174,In_874);
nand U3436 (N_3436,In_27,In_2651);
or U3437 (N_3437,In_1338,In_1734);
xnor U3438 (N_3438,In_1105,In_1660);
and U3439 (N_3439,In_1915,In_2320);
nor U3440 (N_3440,In_5,In_894);
xnor U3441 (N_3441,In_2768,In_2462);
or U3442 (N_3442,In_892,In_1949);
nor U3443 (N_3443,In_2562,In_2099);
xor U3444 (N_3444,In_2273,In_565);
and U3445 (N_3445,In_1692,In_1440);
nor U3446 (N_3446,In_1060,In_235);
nor U3447 (N_3447,In_23,In_1192);
nor U3448 (N_3448,In_106,In_215);
and U3449 (N_3449,In_1091,In_894);
and U3450 (N_3450,In_2118,In_788);
xor U3451 (N_3451,In_58,In_928);
and U3452 (N_3452,In_2533,In_1546);
or U3453 (N_3453,In_2531,In_1231);
xnor U3454 (N_3454,In_1866,In_144);
nand U3455 (N_3455,In_664,In_2588);
nor U3456 (N_3456,In_2521,In_410);
or U3457 (N_3457,In_853,In_77);
nand U3458 (N_3458,In_347,In_1350);
and U3459 (N_3459,In_2937,In_2322);
and U3460 (N_3460,In_496,In_2940);
and U3461 (N_3461,In_2671,In_2837);
xor U3462 (N_3462,In_969,In_1696);
or U3463 (N_3463,In_1275,In_1898);
or U3464 (N_3464,In_1238,In_2145);
nor U3465 (N_3465,In_2599,In_2821);
xnor U3466 (N_3466,In_1243,In_385);
nor U3467 (N_3467,In_2711,In_2622);
nor U3468 (N_3468,In_355,In_2209);
or U3469 (N_3469,In_2526,In_331);
nor U3470 (N_3470,In_1640,In_2445);
and U3471 (N_3471,In_1411,In_1279);
and U3472 (N_3472,In_883,In_2403);
nand U3473 (N_3473,In_195,In_2123);
xnor U3474 (N_3474,In_2711,In_0);
and U3475 (N_3475,In_305,In_106);
xor U3476 (N_3476,In_1872,In_1260);
and U3477 (N_3477,In_165,In_1085);
nand U3478 (N_3478,In_2075,In_1271);
or U3479 (N_3479,In_2249,In_149);
nand U3480 (N_3480,In_1462,In_1342);
nand U3481 (N_3481,In_433,In_901);
nand U3482 (N_3482,In_788,In_873);
xor U3483 (N_3483,In_1145,In_1598);
and U3484 (N_3484,In_622,In_979);
xor U3485 (N_3485,In_1570,In_2118);
nand U3486 (N_3486,In_2814,In_2311);
and U3487 (N_3487,In_2072,In_2662);
and U3488 (N_3488,In_952,In_632);
or U3489 (N_3489,In_1772,In_891);
nand U3490 (N_3490,In_858,In_2740);
nor U3491 (N_3491,In_1328,In_344);
and U3492 (N_3492,In_966,In_1635);
and U3493 (N_3493,In_1394,In_186);
nor U3494 (N_3494,In_2095,In_586);
nand U3495 (N_3495,In_2686,In_1921);
xnor U3496 (N_3496,In_283,In_1909);
and U3497 (N_3497,In_824,In_1365);
xor U3498 (N_3498,In_1633,In_2001);
nor U3499 (N_3499,In_577,In_653);
and U3500 (N_3500,In_1260,In_1227);
nor U3501 (N_3501,In_48,In_919);
or U3502 (N_3502,In_1759,In_1310);
nand U3503 (N_3503,In_2328,In_2584);
xor U3504 (N_3504,In_2483,In_468);
and U3505 (N_3505,In_2521,In_1582);
xor U3506 (N_3506,In_1943,In_1884);
nand U3507 (N_3507,In_1089,In_1728);
or U3508 (N_3508,In_2780,In_450);
and U3509 (N_3509,In_2596,In_2374);
and U3510 (N_3510,In_310,In_1759);
nor U3511 (N_3511,In_889,In_2571);
or U3512 (N_3512,In_1231,In_902);
nor U3513 (N_3513,In_2220,In_2473);
xnor U3514 (N_3514,In_25,In_2818);
nor U3515 (N_3515,In_2380,In_387);
nor U3516 (N_3516,In_1,In_1254);
and U3517 (N_3517,In_640,In_2637);
or U3518 (N_3518,In_1414,In_567);
and U3519 (N_3519,In_846,In_996);
nand U3520 (N_3520,In_794,In_1368);
xor U3521 (N_3521,In_1960,In_1934);
nand U3522 (N_3522,In_1198,In_2636);
nand U3523 (N_3523,In_1619,In_2069);
nand U3524 (N_3524,In_2112,In_2315);
xnor U3525 (N_3525,In_714,In_394);
xor U3526 (N_3526,In_2878,In_1861);
nor U3527 (N_3527,In_2927,In_208);
and U3528 (N_3528,In_2533,In_2412);
nand U3529 (N_3529,In_811,In_990);
nor U3530 (N_3530,In_2509,In_1467);
xor U3531 (N_3531,In_149,In_2542);
or U3532 (N_3532,In_687,In_2719);
xor U3533 (N_3533,In_2211,In_1680);
and U3534 (N_3534,In_854,In_342);
nor U3535 (N_3535,In_102,In_1545);
xor U3536 (N_3536,In_2568,In_2513);
or U3537 (N_3537,In_2980,In_2717);
nand U3538 (N_3538,In_917,In_674);
nor U3539 (N_3539,In_1721,In_151);
and U3540 (N_3540,In_1,In_2035);
nor U3541 (N_3541,In_1033,In_2645);
nand U3542 (N_3542,In_1026,In_2146);
or U3543 (N_3543,In_527,In_1273);
or U3544 (N_3544,In_913,In_406);
or U3545 (N_3545,In_529,In_1072);
xnor U3546 (N_3546,In_1818,In_951);
nor U3547 (N_3547,In_1713,In_1030);
nand U3548 (N_3548,In_1103,In_865);
nor U3549 (N_3549,In_1954,In_1309);
xor U3550 (N_3550,In_727,In_2494);
nand U3551 (N_3551,In_2957,In_2960);
xnor U3552 (N_3552,In_1399,In_1589);
nand U3553 (N_3553,In_1514,In_917);
or U3554 (N_3554,In_963,In_1986);
and U3555 (N_3555,In_761,In_1334);
nand U3556 (N_3556,In_346,In_959);
nand U3557 (N_3557,In_944,In_2466);
nand U3558 (N_3558,In_2464,In_611);
or U3559 (N_3559,In_2084,In_1508);
and U3560 (N_3560,In_2771,In_838);
and U3561 (N_3561,In_2778,In_2144);
xnor U3562 (N_3562,In_1802,In_1395);
nand U3563 (N_3563,In_1885,In_214);
xor U3564 (N_3564,In_81,In_1003);
or U3565 (N_3565,In_2989,In_345);
and U3566 (N_3566,In_1867,In_368);
and U3567 (N_3567,In_423,In_1808);
or U3568 (N_3568,In_1076,In_173);
nor U3569 (N_3569,In_1909,In_823);
and U3570 (N_3570,In_1258,In_2168);
xor U3571 (N_3571,In_2033,In_1009);
nor U3572 (N_3572,In_2907,In_133);
and U3573 (N_3573,In_20,In_390);
xor U3574 (N_3574,In_1880,In_1213);
and U3575 (N_3575,In_892,In_422);
nor U3576 (N_3576,In_921,In_997);
nor U3577 (N_3577,In_363,In_2888);
or U3578 (N_3578,In_1300,In_913);
and U3579 (N_3579,In_2613,In_396);
nand U3580 (N_3580,In_675,In_1786);
nand U3581 (N_3581,In_108,In_236);
or U3582 (N_3582,In_2423,In_1285);
nor U3583 (N_3583,In_1635,In_1785);
or U3584 (N_3584,In_2982,In_135);
and U3585 (N_3585,In_595,In_1609);
nand U3586 (N_3586,In_1552,In_1600);
xnor U3587 (N_3587,In_2258,In_906);
or U3588 (N_3588,In_1004,In_2121);
xnor U3589 (N_3589,In_669,In_2194);
or U3590 (N_3590,In_1558,In_702);
and U3591 (N_3591,In_377,In_1832);
xor U3592 (N_3592,In_2098,In_677);
nor U3593 (N_3593,In_498,In_415);
and U3594 (N_3594,In_1514,In_1424);
nor U3595 (N_3595,In_2671,In_2230);
nor U3596 (N_3596,In_697,In_1403);
and U3597 (N_3597,In_1112,In_2670);
or U3598 (N_3598,In_1052,In_178);
and U3599 (N_3599,In_2244,In_1758);
and U3600 (N_3600,In_781,In_1690);
nand U3601 (N_3601,In_2549,In_1832);
nor U3602 (N_3602,In_435,In_1779);
and U3603 (N_3603,In_2611,In_2937);
or U3604 (N_3604,In_2323,In_1098);
nor U3605 (N_3605,In_1392,In_1399);
xnor U3606 (N_3606,In_1900,In_2160);
nor U3607 (N_3607,In_1940,In_471);
nand U3608 (N_3608,In_1496,In_2515);
or U3609 (N_3609,In_48,In_777);
and U3610 (N_3610,In_785,In_2703);
nor U3611 (N_3611,In_2284,In_1448);
nor U3612 (N_3612,In_2614,In_1167);
nor U3613 (N_3613,In_2278,In_1347);
or U3614 (N_3614,In_1082,In_224);
and U3615 (N_3615,In_1239,In_1310);
or U3616 (N_3616,In_569,In_1269);
and U3617 (N_3617,In_1235,In_2357);
and U3618 (N_3618,In_759,In_436);
nor U3619 (N_3619,In_430,In_989);
nand U3620 (N_3620,In_505,In_102);
xnor U3621 (N_3621,In_1732,In_676);
xor U3622 (N_3622,In_663,In_2052);
nand U3623 (N_3623,In_298,In_1787);
xnor U3624 (N_3624,In_2262,In_2436);
and U3625 (N_3625,In_2143,In_866);
and U3626 (N_3626,In_2909,In_719);
nor U3627 (N_3627,In_2223,In_238);
and U3628 (N_3628,In_113,In_574);
nor U3629 (N_3629,In_2891,In_2014);
or U3630 (N_3630,In_2654,In_2396);
and U3631 (N_3631,In_2437,In_1002);
nor U3632 (N_3632,In_917,In_2394);
nand U3633 (N_3633,In_145,In_244);
or U3634 (N_3634,In_1549,In_2260);
xor U3635 (N_3635,In_2061,In_178);
nor U3636 (N_3636,In_2699,In_1323);
xnor U3637 (N_3637,In_2553,In_1708);
nand U3638 (N_3638,In_2596,In_245);
nor U3639 (N_3639,In_1474,In_2715);
xnor U3640 (N_3640,In_662,In_88);
nor U3641 (N_3641,In_2441,In_954);
nor U3642 (N_3642,In_1617,In_434);
or U3643 (N_3643,In_2212,In_670);
nor U3644 (N_3644,In_2350,In_626);
and U3645 (N_3645,In_793,In_891);
xnor U3646 (N_3646,In_1416,In_2351);
or U3647 (N_3647,In_1347,In_2285);
nand U3648 (N_3648,In_1702,In_2020);
xor U3649 (N_3649,In_1807,In_1267);
nor U3650 (N_3650,In_1098,In_93);
and U3651 (N_3651,In_1062,In_2128);
and U3652 (N_3652,In_321,In_61);
or U3653 (N_3653,In_959,In_829);
xnor U3654 (N_3654,In_1835,In_2451);
or U3655 (N_3655,In_1931,In_2162);
xor U3656 (N_3656,In_53,In_1275);
and U3657 (N_3657,In_782,In_2600);
nor U3658 (N_3658,In_2075,In_2009);
and U3659 (N_3659,In_1980,In_2738);
xor U3660 (N_3660,In_63,In_1215);
nor U3661 (N_3661,In_2262,In_893);
and U3662 (N_3662,In_2532,In_450);
or U3663 (N_3663,In_1385,In_2048);
nand U3664 (N_3664,In_2603,In_1660);
and U3665 (N_3665,In_1542,In_11);
and U3666 (N_3666,In_639,In_1792);
and U3667 (N_3667,In_868,In_2481);
and U3668 (N_3668,In_69,In_2662);
nor U3669 (N_3669,In_2263,In_1608);
nor U3670 (N_3670,In_977,In_2732);
or U3671 (N_3671,In_2188,In_1809);
nand U3672 (N_3672,In_2744,In_557);
xor U3673 (N_3673,In_1533,In_853);
and U3674 (N_3674,In_1599,In_1214);
and U3675 (N_3675,In_1711,In_1541);
xnor U3676 (N_3676,In_481,In_2400);
or U3677 (N_3677,In_92,In_1664);
and U3678 (N_3678,In_1047,In_840);
and U3679 (N_3679,In_2846,In_1624);
nor U3680 (N_3680,In_1724,In_2462);
or U3681 (N_3681,In_2407,In_241);
or U3682 (N_3682,In_276,In_2835);
nor U3683 (N_3683,In_2688,In_1952);
xnor U3684 (N_3684,In_21,In_9);
and U3685 (N_3685,In_210,In_160);
nor U3686 (N_3686,In_1711,In_574);
nand U3687 (N_3687,In_86,In_2128);
or U3688 (N_3688,In_1732,In_473);
or U3689 (N_3689,In_2948,In_174);
nor U3690 (N_3690,In_2973,In_2268);
nor U3691 (N_3691,In_2526,In_1720);
nor U3692 (N_3692,In_802,In_2663);
and U3693 (N_3693,In_1658,In_1852);
or U3694 (N_3694,In_1217,In_559);
or U3695 (N_3695,In_1136,In_2631);
or U3696 (N_3696,In_332,In_723);
and U3697 (N_3697,In_432,In_43);
nand U3698 (N_3698,In_944,In_13);
nand U3699 (N_3699,In_29,In_1663);
nor U3700 (N_3700,In_1230,In_721);
and U3701 (N_3701,In_2598,In_532);
or U3702 (N_3702,In_185,In_2881);
xnor U3703 (N_3703,In_2556,In_2121);
and U3704 (N_3704,In_2668,In_1679);
and U3705 (N_3705,In_863,In_2733);
nand U3706 (N_3706,In_534,In_1182);
and U3707 (N_3707,In_1067,In_728);
xor U3708 (N_3708,In_1093,In_2884);
or U3709 (N_3709,In_1889,In_1129);
nor U3710 (N_3710,In_865,In_1257);
nand U3711 (N_3711,In_1310,In_1494);
xnor U3712 (N_3712,In_907,In_1291);
and U3713 (N_3713,In_1155,In_1419);
or U3714 (N_3714,In_1574,In_963);
or U3715 (N_3715,In_2880,In_120);
nor U3716 (N_3716,In_1232,In_815);
and U3717 (N_3717,In_1379,In_233);
nand U3718 (N_3718,In_2853,In_2387);
and U3719 (N_3719,In_1263,In_2767);
or U3720 (N_3720,In_921,In_31);
xnor U3721 (N_3721,In_545,In_1941);
or U3722 (N_3722,In_221,In_2318);
or U3723 (N_3723,In_917,In_1269);
and U3724 (N_3724,In_1891,In_2945);
nor U3725 (N_3725,In_2279,In_1508);
and U3726 (N_3726,In_1460,In_2392);
xnor U3727 (N_3727,In_1716,In_2357);
nand U3728 (N_3728,In_1689,In_384);
or U3729 (N_3729,In_1014,In_1569);
xnor U3730 (N_3730,In_924,In_1551);
nand U3731 (N_3731,In_2692,In_2067);
nand U3732 (N_3732,In_2976,In_2698);
nor U3733 (N_3733,In_302,In_655);
xnor U3734 (N_3734,In_177,In_733);
or U3735 (N_3735,In_1815,In_2064);
nand U3736 (N_3736,In_1111,In_1033);
and U3737 (N_3737,In_2497,In_2389);
nor U3738 (N_3738,In_2996,In_1146);
nand U3739 (N_3739,In_1627,In_2337);
and U3740 (N_3740,In_19,In_147);
or U3741 (N_3741,In_2790,In_99);
nand U3742 (N_3742,In_31,In_838);
nand U3743 (N_3743,In_2482,In_1454);
and U3744 (N_3744,In_1605,In_663);
and U3745 (N_3745,In_504,In_1702);
nor U3746 (N_3746,In_1673,In_2472);
xnor U3747 (N_3747,In_2375,In_644);
nand U3748 (N_3748,In_788,In_988);
xor U3749 (N_3749,In_1765,In_2094);
nand U3750 (N_3750,In_1630,In_2870);
nand U3751 (N_3751,In_1210,In_1434);
nand U3752 (N_3752,In_1215,In_1907);
nor U3753 (N_3753,In_136,In_1700);
nand U3754 (N_3754,In_700,In_1691);
and U3755 (N_3755,In_1479,In_2007);
nand U3756 (N_3756,In_1795,In_1415);
nor U3757 (N_3757,In_155,In_1541);
xor U3758 (N_3758,In_1371,In_1709);
nand U3759 (N_3759,In_353,In_2438);
xnor U3760 (N_3760,In_594,In_268);
xor U3761 (N_3761,In_2360,In_1018);
nor U3762 (N_3762,In_1514,In_2896);
or U3763 (N_3763,In_1837,In_239);
or U3764 (N_3764,In_1923,In_2856);
nor U3765 (N_3765,In_1063,In_1321);
xnor U3766 (N_3766,In_2372,In_2028);
nor U3767 (N_3767,In_77,In_2977);
or U3768 (N_3768,In_2395,In_1899);
or U3769 (N_3769,In_2028,In_2065);
nand U3770 (N_3770,In_2600,In_2411);
xnor U3771 (N_3771,In_513,In_2581);
and U3772 (N_3772,In_1751,In_980);
nand U3773 (N_3773,In_1190,In_2983);
nand U3774 (N_3774,In_1331,In_1434);
nor U3775 (N_3775,In_2799,In_2127);
xor U3776 (N_3776,In_1601,In_2428);
xor U3777 (N_3777,In_2392,In_1347);
xnor U3778 (N_3778,In_637,In_1565);
xor U3779 (N_3779,In_930,In_414);
xnor U3780 (N_3780,In_2230,In_765);
nor U3781 (N_3781,In_105,In_1181);
nor U3782 (N_3782,In_2569,In_916);
and U3783 (N_3783,In_2463,In_2339);
nand U3784 (N_3784,In_510,In_2453);
nor U3785 (N_3785,In_2923,In_253);
nand U3786 (N_3786,In_278,In_2355);
xor U3787 (N_3787,In_2124,In_966);
or U3788 (N_3788,In_2109,In_511);
nand U3789 (N_3789,In_1890,In_1522);
or U3790 (N_3790,In_2241,In_2414);
and U3791 (N_3791,In_1932,In_2095);
nand U3792 (N_3792,In_1200,In_936);
or U3793 (N_3793,In_1442,In_568);
nor U3794 (N_3794,In_1581,In_943);
xor U3795 (N_3795,In_847,In_1319);
nand U3796 (N_3796,In_2069,In_2602);
xnor U3797 (N_3797,In_1297,In_682);
or U3798 (N_3798,In_39,In_945);
nand U3799 (N_3799,In_1649,In_2457);
nor U3800 (N_3800,In_2196,In_399);
or U3801 (N_3801,In_45,In_1657);
or U3802 (N_3802,In_2944,In_1405);
and U3803 (N_3803,In_2451,In_2437);
nor U3804 (N_3804,In_2719,In_532);
nor U3805 (N_3805,In_1404,In_1211);
nand U3806 (N_3806,In_1947,In_2357);
nand U3807 (N_3807,In_502,In_2356);
and U3808 (N_3808,In_1834,In_2021);
nor U3809 (N_3809,In_2433,In_1710);
and U3810 (N_3810,In_2662,In_261);
xnor U3811 (N_3811,In_2355,In_2129);
xnor U3812 (N_3812,In_2291,In_2460);
nand U3813 (N_3813,In_169,In_1925);
nor U3814 (N_3814,In_2788,In_1203);
or U3815 (N_3815,In_2374,In_1929);
nand U3816 (N_3816,In_914,In_2223);
and U3817 (N_3817,In_606,In_1539);
or U3818 (N_3818,In_718,In_2733);
xor U3819 (N_3819,In_1382,In_1257);
and U3820 (N_3820,In_106,In_800);
nand U3821 (N_3821,In_1613,In_1323);
and U3822 (N_3822,In_957,In_1958);
xnor U3823 (N_3823,In_2746,In_1216);
nand U3824 (N_3824,In_689,In_2345);
and U3825 (N_3825,In_340,In_1054);
nor U3826 (N_3826,In_2504,In_752);
nand U3827 (N_3827,In_2517,In_169);
xnor U3828 (N_3828,In_94,In_1232);
nand U3829 (N_3829,In_2367,In_2580);
and U3830 (N_3830,In_2019,In_2349);
or U3831 (N_3831,In_473,In_2600);
nand U3832 (N_3832,In_2868,In_1010);
nand U3833 (N_3833,In_116,In_744);
nand U3834 (N_3834,In_2096,In_1325);
xor U3835 (N_3835,In_2275,In_2823);
and U3836 (N_3836,In_2514,In_1185);
xor U3837 (N_3837,In_1327,In_1664);
xor U3838 (N_3838,In_2664,In_25);
and U3839 (N_3839,In_1778,In_1900);
nor U3840 (N_3840,In_578,In_1213);
or U3841 (N_3841,In_2820,In_108);
or U3842 (N_3842,In_1255,In_894);
xnor U3843 (N_3843,In_2209,In_2573);
xor U3844 (N_3844,In_146,In_2517);
or U3845 (N_3845,In_2409,In_990);
nand U3846 (N_3846,In_1554,In_2014);
or U3847 (N_3847,In_2342,In_2707);
nor U3848 (N_3848,In_774,In_2292);
xor U3849 (N_3849,In_400,In_1766);
and U3850 (N_3850,In_1545,In_558);
or U3851 (N_3851,In_1382,In_2161);
xor U3852 (N_3852,In_2410,In_959);
nor U3853 (N_3853,In_1117,In_397);
or U3854 (N_3854,In_1170,In_685);
nor U3855 (N_3855,In_1705,In_2561);
nor U3856 (N_3856,In_94,In_893);
and U3857 (N_3857,In_536,In_1752);
or U3858 (N_3858,In_104,In_630);
nor U3859 (N_3859,In_435,In_48);
nor U3860 (N_3860,In_1213,In_2876);
nand U3861 (N_3861,In_1068,In_1811);
nand U3862 (N_3862,In_1392,In_2650);
and U3863 (N_3863,In_409,In_2411);
xor U3864 (N_3864,In_681,In_2329);
or U3865 (N_3865,In_2305,In_1936);
nor U3866 (N_3866,In_1295,In_1371);
or U3867 (N_3867,In_1455,In_2699);
nand U3868 (N_3868,In_2859,In_2782);
xnor U3869 (N_3869,In_400,In_588);
or U3870 (N_3870,In_2725,In_597);
and U3871 (N_3871,In_1690,In_966);
or U3872 (N_3872,In_1708,In_1263);
nand U3873 (N_3873,In_2976,In_2798);
and U3874 (N_3874,In_180,In_345);
or U3875 (N_3875,In_221,In_982);
nand U3876 (N_3876,In_1390,In_1245);
and U3877 (N_3877,In_902,In_1979);
nor U3878 (N_3878,In_1336,In_2805);
nand U3879 (N_3879,In_439,In_2444);
or U3880 (N_3880,In_2675,In_2713);
xnor U3881 (N_3881,In_2750,In_1966);
and U3882 (N_3882,In_1603,In_988);
and U3883 (N_3883,In_1294,In_1654);
xnor U3884 (N_3884,In_2024,In_1868);
nand U3885 (N_3885,In_2872,In_169);
and U3886 (N_3886,In_566,In_1552);
xor U3887 (N_3887,In_2788,In_506);
and U3888 (N_3888,In_1070,In_98);
or U3889 (N_3889,In_2166,In_1950);
and U3890 (N_3890,In_565,In_2665);
and U3891 (N_3891,In_304,In_1940);
and U3892 (N_3892,In_767,In_2929);
nand U3893 (N_3893,In_2222,In_1303);
and U3894 (N_3894,In_242,In_833);
nor U3895 (N_3895,In_1961,In_843);
nand U3896 (N_3896,In_2375,In_749);
xnor U3897 (N_3897,In_654,In_2043);
nand U3898 (N_3898,In_598,In_1379);
nor U3899 (N_3899,In_1863,In_47);
and U3900 (N_3900,In_1882,In_1669);
xnor U3901 (N_3901,In_945,In_2758);
nand U3902 (N_3902,In_2368,In_887);
nor U3903 (N_3903,In_2867,In_853);
xnor U3904 (N_3904,In_2216,In_1231);
or U3905 (N_3905,In_1456,In_744);
xnor U3906 (N_3906,In_2287,In_2239);
nand U3907 (N_3907,In_215,In_2569);
xor U3908 (N_3908,In_2246,In_1474);
and U3909 (N_3909,In_352,In_1962);
nor U3910 (N_3910,In_2950,In_1333);
nand U3911 (N_3911,In_1210,In_1073);
xor U3912 (N_3912,In_930,In_639);
nand U3913 (N_3913,In_116,In_961);
nand U3914 (N_3914,In_2678,In_728);
nor U3915 (N_3915,In_2110,In_2672);
xnor U3916 (N_3916,In_1259,In_447);
nand U3917 (N_3917,In_614,In_497);
xnor U3918 (N_3918,In_1088,In_1558);
xor U3919 (N_3919,In_1196,In_1477);
nor U3920 (N_3920,In_593,In_701);
and U3921 (N_3921,In_244,In_2148);
and U3922 (N_3922,In_576,In_1830);
and U3923 (N_3923,In_1746,In_1537);
or U3924 (N_3924,In_755,In_2153);
or U3925 (N_3925,In_1350,In_1564);
and U3926 (N_3926,In_871,In_613);
xor U3927 (N_3927,In_1138,In_161);
nor U3928 (N_3928,In_1071,In_2188);
xnor U3929 (N_3929,In_1021,In_2671);
or U3930 (N_3930,In_979,In_897);
nor U3931 (N_3931,In_232,In_407);
nand U3932 (N_3932,In_1351,In_2475);
nand U3933 (N_3933,In_1763,In_1205);
xor U3934 (N_3934,In_106,In_2408);
xnor U3935 (N_3935,In_1276,In_2946);
xor U3936 (N_3936,In_525,In_1642);
nand U3937 (N_3937,In_1198,In_1625);
and U3938 (N_3938,In_2985,In_2258);
or U3939 (N_3939,In_1041,In_275);
nor U3940 (N_3940,In_2131,In_260);
xnor U3941 (N_3941,In_1243,In_2847);
xnor U3942 (N_3942,In_2838,In_1213);
and U3943 (N_3943,In_968,In_2858);
xnor U3944 (N_3944,In_2142,In_1995);
xnor U3945 (N_3945,In_509,In_2204);
or U3946 (N_3946,In_2652,In_1132);
nor U3947 (N_3947,In_259,In_1731);
xnor U3948 (N_3948,In_2110,In_1977);
xor U3949 (N_3949,In_221,In_2491);
and U3950 (N_3950,In_2620,In_2733);
nor U3951 (N_3951,In_2961,In_506);
xnor U3952 (N_3952,In_2571,In_1223);
xor U3953 (N_3953,In_1892,In_2353);
or U3954 (N_3954,In_1512,In_1934);
or U3955 (N_3955,In_61,In_2151);
and U3956 (N_3956,In_1107,In_2639);
nand U3957 (N_3957,In_1512,In_694);
and U3958 (N_3958,In_2300,In_1858);
nor U3959 (N_3959,In_2555,In_2590);
nand U3960 (N_3960,In_2686,In_278);
xnor U3961 (N_3961,In_2626,In_1001);
xnor U3962 (N_3962,In_2909,In_2286);
xnor U3963 (N_3963,In_1520,In_581);
nor U3964 (N_3964,In_1632,In_2582);
xnor U3965 (N_3965,In_1061,In_364);
nand U3966 (N_3966,In_1734,In_751);
xor U3967 (N_3967,In_1379,In_2052);
or U3968 (N_3968,In_940,In_2906);
nand U3969 (N_3969,In_2993,In_2615);
xor U3970 (N_3970,In_1683,In_2958);
nand U3971 (N_3971,In_2376,In_434);
and U3972 (N_3972,In_2528,In_1181);
nor U3973 (N_3973,In_593,In_1340);
xnor U3974 (N_3974,In_2192,In_2489);
xnor U3975 (N_3975,In_2699,In_1287);
or U3976 (N_3976,In_329,In_1680);
or U3977 (N_3977,In_1919,In_1534);
and U3978 (N_3978,In_2208,In_661);
or U3979 (N_3979,In_1482,In_2430);
and U3980 (N_3980,In_1135,In_2920);
nor U3981 (N_3981,In_1552,In_58);
xnor U3982 (N_3982,In_984,In_293);
and U3983 (N_3983,In_2449,In_1412);
xor U3984 (N_3984,In_250,In_2032);
or U3985 (N_3985,In_2535,In_2938);
xnor U3986 (N_3986,In_1013,In_2451);
nor U3987 (N_3987,In_2026,In_1476);
nor U3988 (N_3988,In_583,In_2859);
or U3989 (N_3989,In_2871,In_861);
or U3990 (N_3990,In_1163,In_1806);
and U3991 (N_3991,In_116,In_2461);
xor U3992 (N_3992,In_203,In_577);
nor U3993 (N_3993,In_2077,In_2848);
and U3994 (N_3994,In_1267,In_1717);
nand U3995 (N_3995,In_575,In_2104);
nand U3996 (N_3996,In_1401,In_2797);
or U3997 (N_3997,In_1413,In_108);
nand U3998 (N_3998,In_1645,In_215);
and U3999 (N_3999,In_563,In_151);
nand U4000 (N_4000,In_1729,In_1557);
nor U4001 (N_4001,In_2733,In_1631);
and U4002 (N_4002,In_1621,In_2172);
xor U4003 (N_4003,In_2669,In_2075);
xor U4004 (N_4004,In_1704,In_2561);
or U4005 (N_4005,In_1232,In_2129);
or U4006 (N_4006,In_1021,In_2168);
xor U4007 (N_4007,In_2077,In_2954);
xor U4008 (N_4008,In_1913,In_2553);
nor U4009 (N_4009,In_2386,In_695);
or U4010 (N_4010,In_1314,In_623);
or U4011 (N_4011,In_1217,In_2544);
and U4012 (N_4012,In_1225,In_2068);
or U4013 (N_4013,In_1256,In_2751);
and U4014 (N_4014,In_1221,In_381);
nor U4015 (N_4015,In_847,In_555);
xor U4016 (N_4016,In_1392,In_2942);
or U4017 (N_4017,In_1765,In_2111);
xor U4018 (N_4018,In_2867,In_1761);
xor U4019 (N_4019,In_1773,In_1654);
xnor U4020 (N_4020,In_847,In_2105);
and U4021 (N_4021,In_469,In_1331);
nor U4022 (N_4022,In_2642,In_2491);
nand U4023 (N_4023,In_1882,In_1755);
and U4024 (N_4024,In_2866,In_2584);
and U4025 (N_4025,In_2757,In_530);
or U4026 (N_4026,In_1522,In_1487);
nor U4027 (N_4027,In_2535,In_687);
or U4028 (N_4028,In_457,In_1365);
nor U4029 (N_4029,In_2538,In_1305);
xor U4030 (N_4030,In_810,In_620);
xor U4031 (N_4031,In_99,In_90);
xor U4032 (N_4032,In_1917,In_2528);
xor U4033 (N_4033,In_2094,In_1297);
nor U4034 (N_4034,In_2327,In_670);
xor U4035 (N_4035,In_638,In_1780);
and U4036 (N_4036,In_2398,In_699);
xnor U4037 (N_4037,In_183,In_1427);
xnor U4038 (N_4038,In_2274,In_2276);
xor U4039 (N_4039,In_1786,In_1036);
or U4040 (N_4040,In_2488,In_2442);
xor U4041 (N_4041,In_2952,In_2333);
nor U4042 (N_4042,In_275,In_1427);
and U4043 (N_4043,In_1907,In_1687);
and U4044 (N_4044,In_857,In_1457);
or U4045 (N_4045,In_828,In_473);
and U4046 (N_4046,In_1509,In_96);
nor U4047 (N_4047,In_1653,In_2456);
nor U4048 (N_4048,In_2998,In_255);
or U4049 (N_4049,In_2344,In_2516);
and U4050 (N_4050,In_2001,In_1218);
nor U4051 (N_4051,In_777,In_1604);
and U4052 (N_4052,In_1633,In_2733);
nand U4053 (N_4053,In_26,In_1276);
and U4054 (N_4054,In_2145,In_741);
nand U4055 (N_4055,In_215,In_59);
xnor U4056 (N_4056,In_2665,In_870);
nand U4057 (N_4057,In_1389,In_2267);
and U4058 (N_4058,In_1128,In_1478);
nand U4059 (N_4059,In_1364,In_1496);
and U4060 (N_4060,In_525,In_1205);
or U4061 (N_4061,In_1096,In_2765);
nor U4062 (N_4062,In_1241,In_677);
nor U4063 (N_4063,In_238,In_261);
and U4064 (N_4064,In_1424,In_2868);
xor U4065 (N_4065,In_2520,In_2607);
nand U4066 (N_4066,In_1824,In_411);
and U4067 (N_4067,In_2902,In_1876);
and U4068 (N_4068,In_135,In_2749);
or U4069 (N_4069,In_1411,In_2147);
nand U4070 (N_4070,In_688,In_683);
or U4071 (N_4071,In_742,In_340);
nor U4072 (N_4072,In_2528,In_1822);
nor U4073 (N_4073,In_313,In_1481);
xnor U4074 (N_4074,In_2804,In_2020);
or U4075 (N_4075,In_1339,In_174);
nor U4076 (N_4076,In_1497,In_2974);
and U4077 (N_4077,In_930,In_1166);
nand U4078 (N_4078,In_811,In_1077);
nand U4079 (N_4079,In_2190,In_1410);
nor U4080 (N_4080,In_798,In_1480);
nor U4081 (N_4081,In_441,In_907);
nor U4082 (N_4082,In_1936,In_1119);
nor U4083 (N_4083,In_483,In_847);
or U4084 (N_4084,In_179,In_932);
nor U4085 (N_4085,In_2618,In_2435);
xnor U4086 (N_4086,In_2758,In_2331);
or U4087 (N_4087,In_1232,In_778);
nor U4088 (N_4088,In_2798,In_926);
xor U4089 (N_4089,In_1252,In_1037);
or U4090 (N_4090,In_732,In_1843);
nand U4091 (N_4091,In_545,In_455);
or U4092 (N_4092,In_2037,In_2900);
or U4093 (N_4093,In_1114,In_2440);
nor U4094 (N_4094,In_763,In_2293);
nor U4095 (N_4095,In_1744,In_2738);
xnor U4096 (N_4096,In_57,In_885);
xor U4097 (N_4097,In_1744,In_2087);
xor U4098 (N_4098,In_1599,In_130);
nor U4099 (N_4099,In_854,In_1451);
xor U4100 (N_4100,In_377,In_962);
nor U4101 (N_4101,In_1446,In_704);
xor U4102 (N_4102,In_64,In_1579);
and U4103 (N_4103,In_652,In_2971);
and U4104 (N_4104,In_1907,In_1894);
nand U4105 (N_4105,In_1211,In_1339);
nand U4106 (N_4106,In_1220,In_2756);
xor U4107 (N_4107,In_2958,In_912);
xor U4108 (N_4108,In_1652,In_2272);
xor U4109 (N_4109,In_2392,In_2820);
nand U4110 (N_4110,In_2954,In_97);
nor U4111 (N_4111,In_1271,In_752);
or U4112 (N_4112,In_2516,In_1403);
nand U4113 (N_4113,In_2278,In_687);
or U4114 (N_4114,In_2240,In_1589);
or U4115 (N_4115,In_852,In_2058);
xnor U4116 (N_4116,In_1366,In_1198);
nor U4117 (N_4117,In_828,In_508);
xor U4118 (N_4118,In_385,In_855);
xnor U4119 (N_4119,In_2625,In_2081);
nor U4120 (N_4120,In_211,In_349);
xor U4121 (N_4121,In_177,In_806);
xor U4122 (N_4122,In_984,In_1126);
nand U4123 (N_4123,In_821,In_890);
nor U4124 (N_4124,In_2456,In_890);
xnor U4125 (N_4125,In_497,In_2978);
and U4126 (N_4126,In_634,In_2414);
nand U4127 (N_4127,In_1240,In_1212);
xnor U4128 (N_4128,In_2836,In_818);
and U4129 (N_4129,In_748,In_1078);
nand U4130 (N_4130,In_2380,In_834);
and U4131 (N_4131,In_2826,In_823);
or U4132 (N_4132,In_2432,In_1617);
xor U4133 (N_4133,In_2482,In_750);
or U4134 (N_4134,In_2938,In_407);
nor U4135 (N_4135,In_1234,In_723);
nor U4136 (N_4136,In_2344,In_257);
xnor U4137 (N_4137,In_437,In_2421);
and U4138 (N_4138,In_1860,In_1404);
xnor U4139 (N_4139,In_2826,In_626);
nand U4140 (N_4140,In_2684,In_2583);
xnor U4141 (N_4141,In_1135,In_2303);
nand U4142 (N_4142,In_510,In_1692);
and U4143 (N_4143,In_2796,In_1265);
and U4144 (N_4144,In_1611,In_1032);
and U4145 (N_4145,In_2390,In_601);
nor U4146 (N_4146,In_979,In_746);
or U4147 (N_4147,In_408,In_2846);
xor U4148 (N_4148,In_2633,In_2469);
xnor U4149 (N_4149,In_20,In_375);
nor U4150 (N_4150,In_987,In_1703);
xnor U4151 (N_4151,In_952,In_1217);
or U4152 (N_4152,In_393,In_949);
nand U4153 (N_4153,In_913,In_2179);
xor U4154 (N_4154,In_1237,In_1225);
nor U4155 (N_4155,In_2961,In_2448);
nand U4156 (N_4156,In_132,In_295);
nand U4157 (N_4157,In_115,In_2841);
and U4158 (N_4158,In_2554,In_646);
xor U4159 (N_4159,In_2352,In_1630);
nand U4160 (N_4160,In_2670,In_741);
and U4161 (N_4161,In_384,In_54);
and U4162 (N_4162,In_1073,In_1502);
or U4163 (N_4163,In_2854,In_56);
xor U4164 (N_4164,In_366,In_2136);
and U4165 (N_4165,In_209,In_1496);
or U4166 (N_4166,In_779,In_2173);
xor U4167 (N_4167,In_2593,In_1999);
nor U4168 (N_4168,In_1880,In_564);
or U4169 (N_4169,In_1068,In_416);
nor U4170 (N_4170,In_2483,In_833);
nand U4171 (N_4171,In_2227,In_406);
and U4172 (N_4172,In_1422,In_2333);
xor U4173 (N_4173,In_411,In_15);
or U4174 (N_4174,In_2543,In_89);
xor U4175 (N_4175,In_2301,In_2208);
nor U4176 (N_4176,In_2118,In_1128);
nand U4177 (N_4177,In_1588,In_2892);
xor U4178 (N_4178,In_638,In_1565);
nand U4179 (N_4179,In_1435,In_912);
and U4180 (N_4180,In_2451,In_2130);
nor U4181 (N_4181,In_2687,In_1887);
nor U4182 (N_4182,In_733,In_1081);
xnor U4183 (N_4183,In_2109,In_1974);
or U4184 (N_4184,In_645,In_1639);
xnor U4185 (N_4185,In_528,In_1335);
or U4186 (N_4186,In_2677,In_1037);
nor U4187 (N_4187,In_1086,In_2698);
xnor U4188 (N_4188,In_2212,In_2386);
nor U4189 (N_4189,In_498,In_2966);
nor U4190 (N_4190,In_2981,In_2105);
nor U4191 (N_4191,In_491,In_2062);
nor U4192 (N_4192,In_209,In_2349);
xor U4193 (N_4193,In_2168,In_2320);
nand U4194 (N_4194,In_1007,In_912);
nor U4195 (N_4195,In_1539,In_2986);
nor U4196 (N_4196,In_597,In_1754);
nor U4197 (N_4197,In_2624,In_2771);
or U4198 (N_4198,In_2852,In_792);
nand U4199 (N_4199,In_1505,In_665);
or U4200 (N_4200,In_801,In_2281);
xor U4201 (N_4201,In_2750,In_1224);
or U4202 (N_4202,In_1572,In_2251);
and U4203 (N_4203,In_1325,In_1739);
and U4204 (N_4204,In_716,In_994);
nand U4205 (N_4205,In_2577,In_528);
xnor U4206 (N_4206,In_2960,In_889);
nor U4207 (N_4207,In_2834,In_1145);
or U4208 (N_4208,In_621,In_922);
nand U4209 (N_4209,In_706,In_752);
xor U4210 (N_4210,In_1384,In_1332);
or U4211 (N_4211,In_2269,In_1275);
and U4212 (N_4212,In_210,In_760);
or U4213 (N_4213,In_1774,In_1666);
xor U4214 (N_4214,In_1940,In_1248);
nor U4215 (N_4215,In_1990,In_1119);
xor U4216 (N_4216,In_131,In_2180);
nor U4217 (N_4217,In_2659,In_419);
and U4218 (N_4218,In_471,In_2523);
or U4219 (N_4219,In_758,In_2700);
nand U4220 (N_4220,In_2890,In_1618);
or U4221 (N_4221,In_1949,In_477);
nand U4222 (N_4222,In_1180,In_408);
and U4223 (N_4223,In_2258,In_227);
and U4224 (N_4224,In_2836,In_2397);
nor U4225 (N_4225,In_478,In_1709);
or U4226 (N_4226,In_16,In_2617);
nor U4227 (N_4227,In_2728,In_2345);
nand U4228 (N_4228,In_1435,In_483);
or U4229 (N_4229,In_1903,In_1634);
nand U4230 (N_4230,In_2452,In_1670);
and U4231 (N_4231,In_432,In_1927);
and U4232 (N_4232,In_2387,In_956);
nor U4233 (N_4233,In_2717,In_2833);
or U4234 (N_4234,In_1493,In_2607);
and U4235 (N_4235,In_2711,In_409);
or U4236 (N_4236,In_846,In_1948);
or U4237 (N_4237,In_2675,In_1794);
nand U4238 (N_4238,In_1654,In_1958);
nand U4239 (N_4239,In_1442,In_603);
nand U4240 (N_4240,In_1490,In_89);
and U4241 (N_4241,In_2439,In_2513);
nand U4242 (N_4242,In_1654,In_949);
nor U4243 (N_4243,In_2270,In_2716);
and U4244 (N_4244,In_117,In_2532);
nor U4245 (N_4245,In_1860,In_822);
xor U4246 (N_4246,In_1770,In_124);
xnor U4247 (N_4247,In_2931,In_2680);
and U4248 (N_4248,In_2533,In_1580);
nor U4249 (N_4249,In_2471,In_1340);
nor U4250 (N_4250,In_2567,In_2529);
xnor U4251 (N_4251,In_2373,In_765);
and U4252 (N_4252,In_2926,In_1136);
xor U4253 (N_4253,In_960,In_1750);
nand U4254 (N_4254,In_991,In_396);
or U4255 (N_4255,In_1283,In_2036);
nor U4256 (N_4256,In_2690,In_1871);
nor U4257 (N_4257,In_1786,In_344);
and U4258 (N_4258,In_245,In_701);
or U4259 (N_4259,In_1172,In_637);
and U4260 (N_4260,In_463,In_2373);
nor U4261 (N_4261,In_807,In_1361);
xnor U4262 (N_4262,In_1466,In_1248);
nor U4263 (N_4263,In_1789,In_730);
or U4264 (N_4264,In_1296,In_2366);
nand U4265 (N_4265,In_1655,In_204);
nand U4266 (N_4266,In_2400,In_1390);
nor U4267 (N_4267,In_954,In_937);
xnor U4268 (N_4268,In_1824,In_2170);
and U4269 (N_4269,In_2003,In_1999);
xnor U4270 (N_4270,In_2168,In_1547);
or U4271 (N_4271,In_599,In_1701);
and U4272 (N_4272,In_1186,In_394);
or U4273 (N_4273,In_1321,In_1829);
xnor U4274 (N_4274,In_2637,In_2660);
and U4275 (N_4275,In_2554,In_182);
and U4276 (N_4276,In_2687,In_1853);
and U4277 (N_4277,In_1659,In_479);
nand U4278 (N_4278,In_1176,In_2892);
xnor U4279 (N_4279,In_2018,In_2787);
nor U4280 (N_4280,In_814,In_766);
and U4281 (N_4281,In_520,In_1714);
nor U4282 (N_4282,In_312,In_433);
nor U4283 (N_4283,In_372,In_835);
nor U4284 (N_4284,In_2002,In_2146);
nor U4285 (N_4285,In_83,In_2596);
xor U4286 (N_4286,In_1177,In_1455);
nand U4287 (N_4287,In_237,In_362);
or U4288 (N_4288,In_671,In_998);
and U4289 (N_4289,In_119,In_1944);
and U4290 (N_4290,In_1406,In_2018);
and U4291 (N_4291,In_2504,In_2388);
xnor U4292 (N_4292,In_744,In_691);
and U4293 (N_4293,In_1889,In_1684);
xor U4294 (N_4294,In_1631,In_629);
or U4295 (N_4295,In_975,In_2791);
xnor U4296 (N_4296,In_655,In_1408);
nand U4297 (N_4297,In_1947,In_915);
xor U4298 (N_4298,In_1013,In_2350);
or U4299 (N_4299,In_2615,In_382);
or U4300 (N_4300,In_2797,In_1893);
nor U4301 (N_4301,In_576,In_1158);
xnor U4302 (N_4302,In_1563,In_1714);
and U4303 (N_4303,In_790,In_200);
or U4304 (N_4304,In_1519,In_170);
nor U4305 (N_4305,In_1211,In_2256);
nand U4306 (N_4306,In_2132,In_1182);
nor U4307 (N_4307,In_576,In_1959);
nand U4308 (N_4308,In_1811,In_1021);
nand U4309 (N_4309,In_35,In_1216);
nor U4310 (N_4310,In_1240,In_809);
or U4311 (N_4311,In_1175,In_1499);
nand U4312 (N_4312,In_2737,In_2533);
nor U4313 (N_4313,In_2773,In_1190);
nand U4314 (N_4314,In_1783,In_2320);
and U4315 (N_4315,In_470,In_52);
nor U4316 (N_4316,In_2806,In_1086);
nor U4317 (N_4317,In_1683,In_682);
nand U4318 (N_4318,In_2156,In_1978);
or U4319 (N_4319,In_2095,In_211);
xnor U4320 (N_4320,In_1283,In_1138);
nand U4321 (N_4321,In_1121,In_1456);
xor U4322 (N_4322,In_332,In_1439);
or U4323 (N_4323,In_2088,In_1098);
or U4324 (N_4324,In_1848,In_2869);
or U4325 (N_4325,In_1560,In_2490);
and U4326 (N_4326,In_185,In_1035);
xor U4327 (N_4327,In_1005,In_1325);
and U4328 (N_4328,In_1991,In_2286);
xor U4329 (N_4329,In_1900,In_1263);
nor U4330 (N_4330,In_2072,In_1384);
xnor U4331 (N_4331,In_2650,In_1646);
and U4332 (N_4332,In_1387,In_2679);
xnor U4333 (N_4333,In_1611,In_2824);
nor U4334 (N_4334,In_1095,In_2911);
and U4335 (N_4335,In_2201,In_2520);
or U4336 (N_4336,In_422,In_2760);
and U4337 (N_4337,In_2119,In_2302);
nand U4338 (N_4338,In_2396,In_1928);
or U4339 (N_4339,In_2795,In_2559);
or U4340 (N_4340,In_1706,In_317);
nor U4341 (N_4341,In_362,In_1290);
nand U4342 (N_4342,In_1421,In_2293);
or U4343 (N_4343,In_1025,In_2815);
nand U4344 (N_4344,In_1136,In_2376);
nor U4345 (N_4345,In_1114,In_1853);
nand U4346 (N_4346,In_483,In_1720);
xnor U4347 (N_4347,In_521,In_617);
and U4348 (N_4348,In_2233,In_1934);
nand U4349 (N_4349,In_875,In_587);
and U4350 (N_4350,In_2377,In_2425);
xor U4351 (N_4351,In_2501,In_2746);
nand U4352 (N_4352,In_356,In_2310);
xor U4353 (N_4353,In_2742,In_1263);
and U4354 (N_4354,In_2961,In_2592);
nor U4355 (N_4355,In_1352,In_2449);
nand U4356 (N_4356,In_1512,In_1531);
xnor U4357 (N_4357,In_631,In_516);
nor U4358 (N_4358,In_2197,In_183);
or U4359 (N_4359,In_1201,In_2112);
nand U4360 (N_4360,In_2501,In_1620);
or U4361 (N_4361,In_1472,In_2435);
nand U4362 (N_4362,In_1632,In_45);
xor U4363 (N_4363,In_339,In_1159);
nand U4364 (N_4364,In_1827,In_635);
nor U4365 (N_4365,In_620,In_307);
xor U4366 (N_4366,In_2497,In_2050);
xnor U4367 (N_4367,In_463,In_1239);
xor U4368 (N_4368,In_1757,In_198);
nand U4369 (N_4369,In_1862,In_2554);
xnor U4370 (N_4370,In_700,In_1809);
or U4371 (N_4371,In_2139,In_216);
nand U4372 (N_4372,In_2709,In_231);
and U4373 (N_4373,In_671,In_2670);
nor U4374 (N_4374,In_896,In_302);
and U4375 (N_4375,In_2864,In_370);
xnor U4376 (N_4376,In_542,In_994);
xnor U4377 (N_4377,In_450,In_2382);
and U4378 (N_4378,In_2788,In_1377);
nand U4379 (N_4379,In_2247,In_2978);
nor U4380 (N_4380,In_1941,In_1211);
or U4381 (N_4381,In_603,In_326);
xnor U4382 (N_4382,In_2503,In_1980);
and U4383 (N_4383,In_629,In_647);
nand U4384 (N_4384,In_1216,In_2026);
nor U4385 (N_4385,In_2250,In_955);
nand U4386 (N_4386,In_2685,In_2151);
xor U4387 (N_4387,In_934,In_2561);
or U4388 (N_4388,In_343,In_451);
or U4389 (N_4389,In_1193,In_1670);
and U4390 (N_4390,In_2887,In_2850);
and U4391 (N_4391,In_503,In_1143);
nor U4392 (N_4392,In_1252,In_2283);
nor U4393 (N_4393,In_965,In_779);
or U4394 (N_4394,In_260,In_4);
nor U4395 (N_4395,In_720,In_1179);
nand U4396 (N_4396,In_1117,In_2299);
nand U4397 (N_4397,In_2109,In_1522);
and U4398 (N_4398,In_855,In_1219);
and U4399 (N_4399,In_670,In_2436);
nor U4400 (N_4400,In_948,In_1405);
or U4401 (N_4401,In_2036,In_2643);
xnor U4402 (N_4402,In_1552,In_1742);
xnor U4403 (N_4403,In_1909,In_2964);
or U4404 (N_4404,In_1138,In_573);
nor U4405 (N_4405,In_56,In_1388);
and U4406 (N_4406,In_532,In_1115);
nor U4407 (N_4407,In_406,In_1037);
xnor U4408 (N_4408,In_313,In_1844);
or U4409 (N_4409,In_2277,In_1720);
xor U4410 (N_4410,In_2317,In_595);
nand U4411 (N_4411,In_1516,In_2164);
nor U4412 (N_4412,In_2432,In_2576);
or U4413 (N_4413,In_737,In_58);
nor U4414 (N_4414,In_592,In_1523);
xnor U4415 (N_4415,In_1364,In_1112);
nand U4416 (N_4416,In_734,In_329);
nor U4417 (N_4417,In_1537,In_107);
nand U4418 (N_4418,In_2086,In_1666);
nor U4419 (N_4419,In_1665,In_1660);
and U4420 (N_4420,In_324,In_2361);
and U4421 (N_4421,In_1476,In_2643);
or U4422 (N_4422,In_1617,In_1500);
and U4423 (N_4423,In_2228,In_2875);
nor U4424 (N_4424,In_2000,In_1652);
and U4425 (N_4425,In_1094,In_2068);
nand U4426 (N_4426,In_1805,In_1548);
xor U4427 (N_4427,In_2296,In_9);
nand U4428 (N_4428,In_2146,In_189);
or U4429 (N_4429,In_2554,In_803);
or U4430 (N_4430,In_692,In_81);
nand U4431 (N_4431,In_2138,In_1580);
xor U4432 (N_4432,In_2247,In_2236);
or U4433 (N_4433,In_1338,In_94);
xnor U4434 (N_4434,In_1371,In_1825);
nor U4435 (N_4435,In_2116,In_1713);
and U4436 (N_4436,In_1600,In_53);
nor U4437 (N_4437,In_1925,In_2449);
xnor U4438 (N_4438,In_2700,In_2529);
nand U4439 (N_4439,In_56,In_1605);
or U4440 (N_4440,In_846,In_205);
nor U4441 (N_4441,In_2785,In_2189);
xnor U4442 (N_4442,In_362,In_2420);
xor U4443 (N_4443,In_2427,In_2378);
xor U4444 (N_4444,In_2426,In_1982);
nand U4445 (N_4445,In_1259,In_2314);
xnor U4446 (N_4446,In_2144,In_974);
nand U4447 (N_4447,In_2685,In_515);
nand U4448 (N_4448,In_2891,In_2693);
xnor U4449 (N_4449,In_1112,In_1965);
and U4450 (N_4450,In_309,In_362);
xnor U4451 (N_4451,In_1055,In_1618);
nand U4452 (N_4452,In_35,In_2753);
and U4453 (N_4453,In_488,In_1086);
nand U4454 (N_4454,In_548,In_565);
nor U4455 (N_4455,In_2344,In_606);
nand U4456 (N_4456,In_1409,In_1847);
xnor U4457 (N_4457,In_258,In_1694);
nor U4458 (N_4458,In_2368,In_641);
and U4459 (N_4459,In_1335,In_2456);
or U4460 (N_4460,In_1548,In_1463);
or U4461 (N_4461,In_531,In_639);
xnor U4462 (N_4462,In_1784,In_1422);
xnor U4463 (N_4463,In_1052,In_2792);
or U4464 (N_4464,In_1483,In_994);
and U4465 (N_4465,In_2468,In_2812);
and U4466 (N_4466,In_458,In_1598);
xor U4467 (N_4467,In_2791,In_668);
xnor U4468 (N_4468,In_909,In_812);
nand U4469 (N_4469,In_1497,In_799);
and U4470 (N_4470,In_1318,In_1663);
or U4471 (N_4471,In_2066,In_330);
xor U4472 (N_4472,In_2946,In_2898);
nand U4473 (N_4473,In_1905,In_762);
or U4474 (N_4474,In_2718,In_1083);
nor U4475 (N_4475,In_206,In_51);
or U4476 (N_4476,In_2946,In_1408);
nor U4477 (N_4477,In_1730,In_961);
nand U4478 (N_4478,In_995,In_1806);
xnor U4479 (N_4479,In_98,In_182);
nand U4480 (N_4480,In_1539,In_2421);
or U4481 (N_4481,In_413,In_390);
xnor U4482 (N_4482,In_692,In_2919);
nand U4483 (N_4483,In_139,In_2150);
nor U4484 (N_4484,In_1476,In_1209);
nor U4485 (N_4485,In_1540,In_2944);
or U4486 (N_4486,In_1428,In_2867);
nor U4487 (N_4487,In_478,In_327);
xor U4488 (N_4488,In_1219,In_1358);
nand U4489 (N_4489,In_2717,In_1860);
and U4490 (N_4490,In_2821,In_2735);
nor U4491 (N_4491,In_2820,In_1787);
and U4492 (N_4492,In_516,In_748);
nor U4493 (N_4493,In_710,In_1275);
nor U4494 (N_4494,In_2577,In_1058);
nand U4495 (N_4495,In_2296,In_1239);
nand U4496 (N_4496,In_224,In_541);
nand U4497 (N_4497,In_90,In_474);
nand U4498 (N_4498,In_302,In_2476);
or U4499 (N_4499,In_2957,In_2579);
and U4500 (N_4500,In_1095,In_1042);
xor U4501 (N_4501,In_2848,In_1860);
nor U4502 (N_4502,In_2759,In_1236);
nand U4503 (N_4503,In_1739,In_2677);
nor U4504 (N_4504,In_2713,In_1860);
or U4505 (N_4505,In_836,In_2066);
nand U4506 (N_4506,In_1492,In_347);
or U4507 (N_4507,In_1961,In_2913);
xor U4508 (N_4508,In_211,In_878);
nor U4509 (N_4509,In_1332,In_2131);
or U4510 (N_4510,In_978,In_647);
nor U4511 (N_4511,In_1094,In_1612);
or U4512 (N_4512,In_2861,In_454);
xnor U4513 (N_4513,In_2568,In_2224);
nand U4514 (N_4514,In_498,In_2915);
or U4515 (N_4515,In_2521,In_1852);
and U4516 (N_4516,In_312,In_1768);
or U4517 (N_4517,In_1516,In_2870);
nor U4518 (N_4518,In_1338,In_2885);
or U4519 (N_4519,In_780,In_33);
and U4520 (N_4520,In_2314,In_2071);
or U4521 (N_4521,In_638,In_103);
or U4522 (N_4522,In_1892,In_575);
nor U4523 (N_4523,In_2400,In_241);
and U4524 (N_4524,In_2909,In_2816);
nand U4525 (N_4525,In_1266,In_2889);
xnor U4526 (N_4526,In_2059,In_515);
nand U4527 (N_4527,In_1473,In_1825);
or U4528 (N_4528,In_588,In_22);
xnor U4529 (N_4529,In_812,In_1829);
and U4530 (N_4530,In_435,In_883);
nand U4531 (N_4531,In_1139,In_1553);
or U4532 (N_4532,In_129,In_745);
and U4533 (N_4533,In_168,In_505);
nor U4534 (N_4534,In_2326,In_578);
nand U4535 (N_4535,In_2460,In_1956);
xnor U4536 (N_4536,In_72,In_1232);
xor U4537 (N_4537,In_1636,In_32);
nor U4538 (N_4538,In_828,In_1591);
or U4539 (N_4539,In_2471,In_942);
nand U4540 (N_4540,In_1869,In_2834);
nand U4541 (N_4541,In_2373,In_254);
xor U4542 (N_4542,In_718,In_372);
and U4543 (N_4543,In_63,In_2759);
or U4544 (N_4544,In_1659,In_515);
or U4545 (N_4545,In_63,In_2598);
nand U4546 (N_4546,In_2163,In_720);
xor U4547 (N_4547,In_2621,In_80);
xor U4548 (N_4548,In_769,In_1056);
nand U4549 (N_4549,In_2149,In_1682);
xnor U4550 (N_4550,In_210,In_1733);
or U4551 (N_4551,In_2470,In_961);
nor U4552 (N_4552,In_15,In_2172);
or U4553 (N_4553,In_2436,In_814);
or U4554 (N_4554,In_786,In_218);
xor U4555 (N_4555,In_2073,In_347);
xor U4556 (N_4556,In_2640,In_387);
xnor U4557 (N_4557,In_838,In_1160);
nand U4558 (N_4558,In_1718,In_2194);
nor U4559 (N_4559,In_159,In_1367);
and U4560 (N_4560,In_1121,In_139);
nor U4561 (N_4561,In_576,In_2320);
xor U4562 (N_4562,In_714,In_686);
or U4563 (N_4563,In_685,In_2224);
nor U4564 (N_4564,In_1717,In_1951);
and U4565 (N_4565,In_2793,In_1172);
nor U4566 (N_4566,In_2216,In_491);
and U4567 (N_4567,In_819,In_2482);
xnor U4568 (N_4568,In_1513,In_2663);
or U4569 (N_4569,In_1163,In_927);
nand U4570 (N_4570,In_1136,In_1463);
xor U4571 (N_4571,In_760,In_2192);
and U4572 (N_4572,In_434,In_115);
xor U4573 (N_4573,In_2838,In_1558);
or U4574 (N_4574,In_1509,In_2245);
nand U4575 (N_4575,In_495,In_1112);
or U4576 (N_4576,In_514,In_905);
or U4577 (N_4577,In_1286,In_2990);
and U4578 (N_4578,In_1330,In_385);
nand U4579 (N_4579,In_923,In_779);
and U4580 (N_4580,In_2787,In_2745);
and U4581 (N_4581,In_2777,In_929);
nor U4582 (N_4582,In_310,In_2450);
nor U4583 (N_4583,In_2257,In_292);
nor U4584 (N_4584,In_1800,In_70);
or U4585 (N_4585,In_418,In_535);
nand U4586 (N_4586,In_2284,In_1577);
and U4587 (N_4587,In_2606,In_1128);
or U4588 (N_4588,In_1665,In_1411);
nand U4589 (N_4589,In_1707,In_1925);
xor U4590 (N_4590,In_2061,In_2596);
xnor U4591 (N_4591,In_2431,In_1805);
nor U4592 (N_4592,In_1159,In_241);
and U4593 (N_4593,In_2519,In_601);
nand U4594 (N_4594,In_281,In_1921);
nand U4595 (N_4595,In_2619,In_613);
nor U4596 (N_4596,In_2501,In_1382);
nand U4597 (N_4597,In_792,In_501);
nand U4598 (N_4598,In_1445,In_1837);
xor U4599 (N_4599,In_2520,In_1942);
nand U4600 (N_4600,In_1674,In_1708);
nand U4601 (N_4601,In_2297,In_2983);
nand U4602 (N_4602,In_70,In_689);
nor U4603 (N_4603,In_1759,In_552);
or U4604 (N_4604,In_567,In_721);
and U4605 (N_4605,In_1222,In_583);
nor U4606 (N_4606,In_1992,In_771);
and U4607 (N_4607,In_1667,In_465);
and U4608 (N_4608,In_2197,In_36);
or U4609 (N_4609,In_2663,In_411);
xor U4610 (N_4610,In_1026,In_320);
and U4611 (N_4611,In_466,In_2185);
or U4612 (N_4612,In_1273,In_2109);
xnor U4613 (N_4613,In_2027,In_828);
nand U4614 (N_4614,In_1721,In_133);
nor U4615 (N_4615,In_24,In_1923);
nor U4616 (N_4616,In_380,In_1301);
nor U4617 (N_4617,In_592,In_487);
nor U4618 (N_4618,In_598,In_923);
xor U4619 (N_4619,In_465,In_2951);
xnor U4620 (N_4620,In_1568,In_533);
and U4621 (N_4621,In_2068,In_2746);
xor U4622 (N_4622,In_318,In_2464);
xnor U4623 (N_4623,In_578,In_69);
nor U4624 (N_4624,In_1567,In_1759);
nand U4625 (N_4625,In_715,In_2586);
or U4626 (N_4626,In_201,In_1012);
or U4627 (N_4627,In_1294,In_1558);
nor U4628 (N_4628,In_867,In_2794);
or U4629 (N_4629,In_802,In_2840);
xnor U4630 (N_4630,In_1250,In_2211);
and U4631 (N_4631,In_894,In_1896);
and U4632 (N_4632,In_605,In_734);
or U4633 (N_4633,In_710,In_1858);
and U4634 (N_4634,In_989,In_2952);
and U4635 (N_4635,In_980,In_427);
nand U4636 (N_4636,In_1816,In_2554);
or U4637 (N_4637,In_2851,In_1486);
nor U4638 (N_4638,In_2807,In_838);
and U4639 (N_4639,In_1965,In_501);
xnor U4640 (N_4640,In_2678,In_1808);
and U4641 (N_4641,In_1048,In_2082);
nor U4642 (N_4642,In_2589,In_1448);
or U4643 (N_4643,In_1893,In_2411);
or U4644 (N_4644,In_887,In_2213);
or U4645 (N_4645,In_2009,In_1188);
xor U4646 (N_4646,In_1176,In_1669);
nor U4647 (N_4647,In_674,In_2083);
and U4648 (N_4648,In_2227,In_354);
nor U4649 (N_4649,In_363,In_1072);
nand U4650 (N_4650,In_1721,In_500);
and U4651 (N_4651,In_206,In_331);
and U4652 (N_4652,In_400,In_1262);
nand U4653 (N_4653,In_1873,In_1021);
nand U4654 (N_4654,In_1524,In_251);
or U4655 (N_4655,In_1032,In_2494);
or U4656 (N_4656,In_755,In_571);
nand U4657 (N_4657,In_88,In_2211);
xnor U4658 (N_4658,In_1117,In_2158);
and U4659 (N_4659,In_1764,In_2642);
nor U4660 (N_4660,In_321,In_2676);
or U4661 (N_4661,In_1170,In_2189);
or U4662 (N_4662,In_1348,In_514);
nor U4663 (N_4663,In_926,In_1382);
nor U4664 (N_4664,In_309,In_2795);
and U4665 (N_4665,In_585,In_2695);
nor U4666 (N_4666,In_901,In_1102);
nand U4667 (N_4667,In_2040,In_2776);
and U4668 (N_4668,In_893,In_2504);
nand U4669 (N_4669,In_2704,In_339);
nand U4670 (N_4670,In_1126,In_2417);
xnor U4671 (N_4671,In_2517,In_1344);
or U4672 (N_4672,In_2331,In_2467);
and U4673 (N_4673,In_1870,In_1285);
nor U4674 (N_4674,In_815,In_1870);
xnor U4675 (N_4675,In_1847,In_687);
or U4676 (N_4676,In_334,In_1751);
nand U4677 (N_4677,In_2251,In_1442);
or U4678 (N_4678,In_1694,In_3);
nor U4679 (N_4679,In_1150,In_2708);
xnor U4680 (N_4680,In_1190,In_2235);
xnor U4681 (N_4681,In_2980,In_2732);
xnor U4682 (N_4682,In_2554,In_732);
xnor U4683 (N_4683,In_1544,In_1507);
nor U4684 (N_4684,In_474,In_1845);
nand U4685 (N_4685,In_2685,In_2866);
or U4686 (N_4686,In_873,In_267);
nand U4687 (N_4687,In_2150,In_1388);
nand U4688 (N_4688,In_1431,In_2287);
or U4689 (N_4689,In_111,In_1726);
nor U4690 (N_4690,In_883,In_2342);
nor U4691 (N_4691,In_806,In_1038);
nor U4692 (N_4692,In_2376,In_112);
or U4693 (N_4693,In_1348,In_944);
xnor U4694 (N_4694,In_618,In_2714);
nand U4695 (N_4695,In_808,In_1499);
nor U4696 (N_4696,In_2204,In_812);
xnor U4697 (N_4697,In_2564,In_2605);
and U4698 (N_4698,In_947,In_2906);
nand U4699 (N_4699,In_2649,In_2934);
and U4700 (N_4700,In_1347,In_1464);
or U4701 (N_4701,In_2307,In_1374);
nor U4702 (N_4702,In_1121,In_1901);
and U4703 (N_4703,In_2199,In_1451);
xnor U4704 (N_4704,In_82,In_467);
and U4705 (N_4705,In_2426,In_1909);
nand U4706 (N_4706,In_1581,In_1060);
nand U4707 (N_4707,In_615,In_1594);
or U4708 (N_4708,In_1897,In_134);
xnor U4709 (N_4709,In_957,In_612);
nand U4710 (N_4710,In_652,In_2660);
xor U4711 (N_4711,In_540,In_1129);
nand U4712 (N_4712,In_110,In_109);
xor U4713 (N_4713,In_453,In_1940);
or U4714 (N_4714,In_2246,In_597);
and U4715 (N_4715,In_569,In_585);
or U4716 (N_4716,In_1667,In_2558);
nand U4717 (N_4717,In_55,In_2088);
nand U4718 (N_4718,In_1791,In_1542);
xnor U4719 (N_4719,In_583,In_1706);
xnor U4720 (N_4720,In_1523,In_2498);
nor U4721 (N_4721,In_1119,In_1438);
nand U4722 (N_4722,In_691,In_2684);
or U4723 (N_4723,In_1765,In_2747);
and U4724 (N_4724,In_2140,In_518);
nand U4725 (N_4725,In_2075,In_2522);
xor U4726 (N_4726,In_1867,In_1123);
and U4727 (N_4727,In_676,In_2838);
or U4728 (N_4728,In_1508,In_594);
xor U4729 (N_4729,In_1488,In_1928);
and U4730 (N_4730,In_98,In_1281);
nor U4731 (N_4731,In_2393,In_2832);
nand U4732 (N_4732,In_2786,In_2849);
nor U4733 (N_4733,In_2238,In_2019);
or U4734 (N_4734,In_2885,In_1717);
or U4735 (N_4735,In_555,In_2796);
or U4736 (N_4736,In_2409,In_1040);
and U4737 (N_4737,In_1082,In_2122);
xnor U4738 (N_4738,In_2479,In_641);
nand U4739 (N_4739,In_1320,In_2327);
or U4740 (N_4740,In_2024,In_2291);
nor U4741 (N_4741,In_2022,In_1926);
or U4742 (N_4742,In_2439,In_667);
nor U4743 (N_4743,In_2170,In_1024);
nand U4744 (N_4744,In_2835,In_2521);
xnor U4745 (N_4745,In_1111,In_760);
nand U4746 (N_4746,In_2283,In_2640);
or U4747 (N_4747,In_2742,In_2394);
nand U4748 (N_4748,In_1917,In_1417);
nor U4749 (N_4749,In_1485,In_2191);
and U4750 (N_4750,In_652,In_2772);
and U4751 (N_4751,In_1767,In_1588);
and U4752 (N_4752,In_1230,In_2227);
xnor U4753 (N_4753,In_736,In_1044);
and U4754 (N_4754,In_195,In_2816);
xnor U4755 (N_4755,In_1865,In_2018);
nand U4756 (N_4756,In_36,In_2887);
nand U4757 (N_4757,In_1727,In_1972);
or U4758 (N_4758,In_2733,In_613);
xnor U4759 (N_4759,In_1210,In_1341);
xnor U4760 (N_4760,In_1029,In_328);
xor U4761 (N_4761,In_1666,In_518);
and U4762 (N_4762,In_1887,In_906);
and U4763 (N_4763,In_1636,In_326);
nor U4764 (N_4764,In_912,In_1044);
and U4765 (N_4765,In_1612,In_1758);
and U4766 (N_4766,In_1447,In_2043);
nor U4767 (N_4767,In_896,In_2205);
and U4768 (N_4768,In_2696,In_1571);
and U4769 (N_4769,In_2417,In_674);
xor U4770 (N_4770,In_1564,In_1773);
xnor U4771 (N_4771,In_791,In_707);
nor U4772 (N_4772,In_2546,In_727);
or U4773 (N_4773,In_1451,In_2347);
or U4774 (N_4774,In_1519,In_797);
and U4775 (N_4775,In_1729,In_1738);
xnor U4776 (N_4776,In_2582,In_2758);
xnor U4777 (N_4777,In_560,In_2634);
or U4778 (N_4778,In_460,In_2800);
xnor U4779 (N_4779,In_2983,In_2806);
and U4780 (N_4780,In_2837,In_781);
nand U4781 (N_4781,In_1282,In_2804);
and U4782 (N_4782,In_122,In_1617);
or U4783 (N_4783,In_2270,In_2538);
and U4784 (N_4784,In_2903,In_807);
or U4785 (N_4785,In_387,In_622);
nor U4786 (N_4786,In_1563,In_2879);
nor U4787 (N_4787,In_56,In_2563);
xnor U4788 (N_4788,In_239,In_566);
nor U4789 (N_4789,In_1846,In_239);
xor U4790 (N_4790,In_1980,In_2185);
or U4791 (N_4791,In_2587,In_2906);
or U4792 (N_4792,In_2647,In_2528);
xor U4793 (N_4793,In_1093,In_1462);
or U4794 (N_4794,In_2597,In_2314);
or U4795 (N_4795,In_2112,In_1610);
and U4796 (N_4796,In_2911,In_2267);
or U4797 (N_4797,In_883,In_156);
nor U4798 (N_4798,In_653,In_184);
nand U4799 (N_4799,In_2873,In_1481);
nor U4800 (N_4800,In_116,In_1870);
nor U4801 (N_4801,In_562,In_881);
xor U4802 (N_4802,In_1162,In_1927);
and U4803 (N_4803,In_586,In_2800);
nand U4804 (N_4804,In_385,In_1061);
and U4805 (N_4805,In_2261,In_126);
xor U4806 (N_4806,In_2636,In_2545);
and U4807 (N_4807,In_1569,In_1324);
nand U4808 (N_4808,In_785,In_1123);
xor U4809 (N_4809,In_1024,In_2216);
and U4810 (N_4810,In_2379,In_2451);
xor U4811 (N_4811,In_2053,In_2778);
and U4812 (N_4812,In_2667,In_565);
or U4813 (N_4813,In_626,In_663);
nand U4814 (N_4814,In_1492,In_842);
or U4815 (N_4815,In_1489,In_1116);
and U4816 (N_4816,In_981,In_872);
nor U4817 (N_4817,In_1326,In_456);
and U4818 (N_4818,In_2808,In_1026);
and U4819 (N_4819,In_2654,In_2448);
and U4820 (N_4820,In_1712,In_1406);
or U4821 (N_4821,In_1352,In_2153);
or U4822 (N_4822,In_1386,In_1939);
nand U4823 (N_4823,In_976,In_2623);
nor U4824 (N_4824,In_1421,In_1764);
xnor U4825 (N_4825,In_2179,In_783);
nand U4826 (N_4826,In_862,In_442);
nor U4827 (N_4827,In_920,In_2941);
and U4828 (N_4828,In_1290,In_2986);
or U4829 (N_4829,In_1644,In_2698);
nor U4830 (N_4830,In_2579,In_2674);
nand U4831 (N_4831,In_81,In_574);
or U4832 (N_4832,In_2280,In_1676);
xor U4833 (N_4833,In_737,In_2054);
nand U4834 (N_4834,In_2470,In_1480);
nor U4835 (N_4835,In_2656,In_1846);
and U4836 (N_4836,In_2254,In_2890);
or U4837 (N_4837,In_56,In_1361);
or U4838 (N_4838,In_571,In_1927);
or U4839 (N_4839,In_2134,In_1484);
xnor U4840 (N_4840,In_1415,In_705);
nor U4841 (N_4841,In_1002,In_2288);
or U4842 (N_4842,In_2691,In_1295);
xor U4843 (N_4843,In_481,In_1116);
and U4844 (N_4844,In_675,In_832);
or U4845 (N_4845,In_1580,In_1397);
xnor U4846 (N_4846,In_2743,In_507);
xor U4847 (N_4847,In_2353,In_498);
xor U4848 (N_4848,In_2759,In_156);
nor U4849 (N_4849,In_426,In_1916);
or U4850 (N_4850,In_2716,In_2145);
nand U4851 (N_4851,In_383,In_2387);
nand U4852 (N_4852,In_754,In_1826);
or U4853 (N_4853,In_2273,In_1206);
and U4854 (N_4854,In_2988,In_1855);
and U4855 (N_4855,In_1581,In_1910);
and U4856 (N_4856,In_1692,In_1296);
or U4857 (N_4857,In_60,In_1808);
nand U4858 (N_4858,In_2672,In_2009);
xor U4859 (N_4859,In_1764,In_599);
nor U4860 (N_4860,In_2745,In_2453);
or U4861 (N_4861,In_2817,In_253);
nand U4862 (N_4862,In_1488,In_2353);
xor U4863 (N_4863,In_1669,In_2059);
nor U4864 (N_4864,In_2661,In_58);
and U4865 (N_4865,In_2446,In_40);
or U4866 (N_4866,In_890,In_797);
or U4867 (N_4867,In_1808,In_2699);
and U4868 (N_4868,In_2563,In_2210);
xor U4869 (N_4869,In_392,In_1150);
or U4870 (N_4870,In_2333,In_107);
nand U4871 (N_4871,In_270,In_1403);
or U4872 (N_4872,In_2481,In_385);
nand U4873 (N_4873,In_553,In_538);
xor U4874 (N_4874,In_856,In_486);
nor U4875 (N_4875,In_2777,In_2917);
xnor U4876 (N_4876,In_291,In_1185);
or U4877 (N_4877,In_2365,In_296);
or U4878 (N_4878,In_50,In_62);
and U4879 (N_4879,In_2820,In_1383);
and U4880 (N_4880,In_58,In_1903);
or U4881 (N_4881,In_1567,In_2181);
xor U4882 (N_4882,In_334,In_2667);
nor U4883 (N_4883,In_2877,In_410);
or U4884 (N_4884,In_2810,In_2665);
nor U4885 (N_4885,In_577,In_226);
nand U4886 (N_4886,In_627,In_2017);
nand U4887 (N_4887,In_2304,In_1966);
nor U4888 (N_4888,In_226,In_2287);
nor U4889 (N_4889,In_1525,In_788);
and U4890 (N_4890,In_1134,In_826);
or U4891 (N_4891,In_2835,In_1595);
and U4892 (N_4892,In_1779,In_361);
xnor U4893 (N_4893,In_1903,In_2110);
or U4894 (N_4894,In_1297,In_456);
nor U4895 (N_4895,In_2672,In_2103);
xor U4896 (N_4896,In_1574,In_2092);
and U4897 (N_4897,In_2315,In_1746);
xor U4898 (N_4898,In_2025,In_2068);
nor U4899 (N_4899,In_2020,In_1912);
or U4900 (N_4900,In_868,In_0);
xor U4901 (N_4901,In_1447,In_590);
nor U4902 (N_4902,In_2591,In_2961);
nor U4903 (N_4903,In_1254,In_640);
nand U4904 (N_4904,In_813,In_1239);
nor U4905 (N_4905,In_638,In_2152);
nand U4906 (N_4906,In_725,In_353);
xor U4907 (N_4907,In_214,In_1849);
nand U4908 (N_4908,In_2899,In_2900);
and U4909 (N_4909,In_2588,In_2731);
and U4910 (N_4910,In_2384,In_2889);
and U4911 (N_4911,In_724,In_2099);
nand U4912 (N_4912,In_953,In_220);
xnor U4913 (N_4913,In_897,In_1527);
or U4914 (N_4914,In_982,In_1519);
or U4915 (N_4915,In_1313,In_2468);
xor U4916 (N_4916,In_1116,In_208);
or U4917 (N_4917,In_680,In_2211);
or U4918 (N_4918,In_1124,In_1660);
nor U4919 (N_4919,In_310,In_2071);
and U4920 (N_4920,In_2222,In_2865);
or U4921 (N_4921,In_1944,In_1575);
or U4922 (N_4922,In_1122,In_410);
and U4923 (N_4923,In_2484,In_361);
xnor U4924 (N_4924,In_284,In_2424);
nor U4925 (N_4925,In_1150,In_1962);
or U4926 (N_4926,In_1276,In_2391);
and U4927 (N_4927,In_1069,In_2676);
xnor U4928 (N_4928,In_2245,In_941);
xnor U4929 (N_4929,In_1269,In_1279);
xor U4930 (N_4930,In_2375,In_1955);
and U4931 (N_4931,In_202,In_1721);
or U4932 (N_4932,In_914,In_197);
xnor U4933 (N_4933,In_1377,In_2915);
nor U4934 (N_4934,In_1773,In_2122);
nand U4935 (N_4935,In_718,In_2259);
or U4936 (N_4936,In_1249,In_1421);
nor U4937 (N_4937,In_220,In_2949);
nand U4938 (N_4938,In_2887,In_1320);
nor U4939 (N_4939,In_299,In_1583);
or U4940 (N_4940,In_2883,In_2652);
or U4941 (N_4941,In_1078,In_746);
nor U4942 (N_4942,In_362,In_134);
xor U4943 (N_4943,In_1729,In_179);
or U4944 (N_4944,In_2920,In_2339);
and U4945 (N_4945,In_2959,In_372);
nand U4946 (N_4946,In_328,In_488);
or U4947 (N_4947,In_2866,In_1471);
or U4948 (N_4948,In_2348,In_2323);
nor U4949 (N_4949,In_1812,In_2373);
and U4950 (N_4950,In_2915,In_2852);
xnor U4951 (N_4951,In_1707,In_281);
xor U4952 (N_4952,In_639,In_2236);
xor U4953 (N_4953,In_1830,In_1722);
and U4954 (N_4954,In_2315,In_1597);
nor U4955 (N_4955,In_1589,In_1265);
nor U4956 (N_4956,In_341,In_1465);
nor U4957 (N_4957,In_653,In_1173);
xnor U4958 (N_4958,In_2874,In_484);
and U4959 (N_4959,In_2933,In_438);
nand U4960 (N_4960,In_472,In_499);
or U4961 (N_4961,In_2478,In_136);
nand U4962 (N_4962,In_1031,In_1216);
nand U4963 (N_4963,In_1076,In_2286);
or U4964 (N_4964,In_1513,In_998);
and U4965 (N_4965,In_1957,In_2243);
or U4966 (N_4966,In_358,In_1880);
nor U4967 (N_4967,In_733,In_330);
nor U4968 (N_4968,In_2318,In_1034);
and U4969 (N_4969,In_1288,In_354);
nor U4970 (N_4970,In_2394,In_2623);
nand U4971 (N_4971,In_995,In_606);
nor U4972 (N_4972,In_5,In_2897);
and U4973 (N_4973,In_183,In_1792);
nor U4974 (N_4974,In_416,In_1317);
nand U4975 (N_4975,In_332,In_2008);
and U4976 (N_4976,In_685,In_2851);
xnor U4977 (N_4977,In_1462,In_419);
nand U4978 (N_4978,In_2121,In_2388);
nand U4979 (N_4979,In_1779,In_1080);
nand U4980 (N_4980,In_261,In_2510);
or U4981 (N_4981,In_1741,In_937);
xor U4982 (N_4982,In_834,In_2104);
nor U4983 (N_4983,In_1321,In_192);
xor U4984 (N_4984,In_934,In_951);
and U4985 (N_4985,In_1811,In_107);
nor U4986 (N_4986,In_1975,In_1112);
nand U4987 (N_4987,In_802,In_1783);
and U4988 (N_4988,In_887,In_572);
or U4989 (N_4989,In_2354,In_1402);
nor U4990 (N_4990,In_1584,In_514);
xnor U4991 (N_4991,In_2303,In_2894);
nand U4992 (N_4992,In_2073,In_2982);
xnor U4993 (N_4993,In_554,In_1608);
or U4994 (N_4994,In_1771,In_255);
nor U4995 (N_4995,In_2415,In_676);
or U4996 (N_4996,In_2416,In_598);
nand U4997 (N_4997,In_1135,In_1695);
nand U4998 (N_4998,In_2013,In_316);
nor U4999 (N_4999,In_1115,In_2647);
nor U5000 (N_5000,In_1427,In_0);
xor U5001 (N_5001,In_2050,In_1362);
nor U5002 (N_5002,In_2809,In_1330);
nor U5003 (N_5003,In_1485,In_1090);
nor U5004 (N_5004,In_1569,In_2403);
xnor U5005 (N_5005,In_2666,In_1630);
and U5006 (N_5006,In_1130,In_83);
nand U5007 (N_5007,In_1131,In_402);
and U5008 (N_5008,In_2002,In_2337);
nand U5009 (N_5009,In_2975,In_1444);
nor U5010 (N_5010,In_2130,In_199);
or U5011 (N_5011,In_1540,In_778);
xor U5012 (N_5012,In_1143,In_1254);
nor U5013 (N_5013,In_181,In_563);
nand U5014 (N_5014,In_1212,In_1256);
or U5015 (N_5015,In_62,In_1754);
and U5016 (N_5016,In_1687,In_2010);
nor U5017 (N_5017,In_1076,In_2062);
nand U5018 (N_5018,In_2360,In_2982);
and U5019 (N_5019,In_2689,In_2045);
and U5020 (N_5020,In_676,In_389);
xor U5021 (N_5021,In_530,In_2080);
or U5022 (N_5022,In_1060,In_2843);
or U5023 (N_5023,In_2429,In_2626);
nand U5024 (N_5024,In_945,In_1596);
nand U5025 (N_5025,In_1562,In_2787);
and U5026 (N_5026,In_367,In_2734);
or U5027 (N_5027,In_2416,In_480);
or U5028 (N_5028,In_292,In_1799);
nand U5029 (N_5029,In_796,In_1631);
nor U5030 (N_5030,In_2264,In_1280);
xor U5031 (N_5031,In_2515,In_2837);
xnor U5032 (N_5032,In_556,In_272);
nor U5033 (N_5033,In_604,In_647);
and U5034 (N_5034,In_707,In_1827);
and U5035 (N_5035,In_1823,In_619);
and U5036 (N_5036,In_1859,In_2149);
or U5037 (N_5037,In_2174,In_1516);
nor U5038 (N_5038,In_558,In_2653);
nor U5039 (N_5039,In_1520,In_160);
nor U5040 (N_5040,In_1873,In_1047);
nor U5041 (N_5041,In_1205,In_1929);
nor U5042 (N_5042,In_849,In_2713);
nand U5043 (N_5043,In_2762,In_1699);
nor U5044 (N_5044,In_2015,In_489);
or U5045 (N_5045,In_1387,In_697);
or U5046 (N_5046,In_1296,In_2518);
xor U5047 (N_5047,In_1506,In_780);
xor U5048 (N_5048,In_1795,In_2044);
nand U5049 (N_5049,In_1658,In_1421);
and U5050 (N_5050,In_2476,In_2169);
nor U5051 (N_5051,In_1464,In_2240);
or U5052 (N_5052,In_1125,In_2173);
xnor U5053 (N_5053,In_1100,In_1477);
nand U5054 (N_5054,In_1596,In_2533);
xnor U5055 (N_5055,In_913,In_1079);
and U5056 (N_5056,In_261,In_529);
nand U5057 (N_5057,In_2065,In_2821);
nand U5058 (N_5058,In_1504,In_625);
nor U5059 (N_5059,In_1414,In_331);
nand U5060 (N_5060,In_248,In_1019);
or U5061 (N_5061,In_443,In_723);
or U5062 (N_5062,In_1012,In_1570);
nand U5063 (N_5063,In_1754,In_1788);
nor U5064 (N_5064,In_929,In_775);
or U5065 (N_5065,In_2991,In_616);
and U5066 (N_5066,In_2206,In_623);
and U5067 (N_5067,In_1861,In_475);
and U5068 (N_5068,In_1748,In_785);
xor U5069 (N_5069,In_2364,In_2273);
and U5070 (N_5070,In_297,In_1152);
nor U5071 (N_5071,In_2254,In_2143);
or U5072 (N_5072,In_499,In_1747);
nor U5073 (N_5073,In_944,In_1458);
or U5074 (N_5074,In_254,In_550);
nand U5075 (N_5075,In_1508,In_1928);
nand U5076 (N_5076,In_2381,In_2458);
xor U5077 (N_5077,In_1672,In_2656);
xor U5078 (N_5078,In_2993,In_2811);
or U5079 (N_5079,In_781,In_2650);
or U5080 (N_5080,In_2669,In_2041);
nor U5081 (N_5081,In_2442,In_246);
or U5082 (N_5082,In_2087,In_632);
and U5083 (N_5083,In_1847,In_2729);
or U5084 (N_5084,In_837,In_516);
xor U5085 (N_5085,In_836,In_1360);
and U5086 (N_5086,In_902,In_2066);
nand U5087 (N_5087,In_691,In_1519);
nand U5088 (N_5088,In_1658,In_2467);
nor U5089 (N_5089,In_2923,In_180);
and U5090 (N_5090,In_152,In_1684);
or U5091 (N_5091,In_1925,In_1391);
nand U5092 (N_5092,In_895,In_1728);
and U5093 (N_5093,In_862,In_1341);
or U5094 (N_5094,In_2727,In_2345);
or U5095 (N_5095,In_1592,In_1262);
and U5096 (N_5096,In_634,In_384);
nand U5097 (N_5097,In_557,In_244);
or U5098 (N_5098,In_288,In_844);
nand U5099 (N_5099,In_1156,In_2279);
nor U5100 (N_5100,In_604,In_610);
xnor U5101 (N_5101,In_856,In_1573);
and U5102 (N_5102,In_376,In_1058);
and U5103 (N_5103,In_2311,In_1574);
and U5104 (N_5104,In_2723,In_390);
and U5105 (N_5105,In_1690,In_1269);
nor U5106 (N_5106,In_2528,In_1456);
nand U5107 (N_5107,In_1217,In_629);
or U5108 (N_5108,In_2963,In_1957);
xnor U5109 (N_5109,In_1367,In_271);
nor U5110 (N_5110,In_2796,In_922);
or U5111 (N_5111,In_1663,In_418);
and U5112 (N_5112,In_338,In_243);
nor U5113 (N_5113,In_2478,In_2573);
nand U5114 (N_5114,In_2979,In_2468);
and U5115 (N_5115,In_1098,In_576);
nand U5116 (N_5116,In_1632,In_1638);
nand U5117 (N_5117,In_2602,In_75);
or U5118 (N_5118,In_1878,In_140);
or U5119 (N_5119,In_393,In_1437);
nand U5120 (N_5120,In_478,In_793);
xor U5121 (N_5121,In_1091,In_2102);
and U5122 (N_5122,In_2309,In_612);
xor U5123 (N_5123,In_1592,In_2180);
xnor U5124 (N_5124,In_2351,In_404);
xor U5125 (N_5125,In_2077,In_2117);
xnor U5126 (N_5126,In_2215,In_1052);
nand U5127 (N_5127,In_2091,In_419);
or U5128 (N_5128,In_1803,In_2730);
nand U5129 (N_5129,In_35,In_639);
xor U5130 (N_5130,In_2012,In_2096);
or U5131 (N_5131,In_2377,In_1516);
and U5132 (N_5132,In_2621,In_2703);
xnor U5133 (N_5133,In_361,In_1175);
nand U5134 (N_5134,In_2684,In_2199);
and U5135 (N_5135,In_1766,In_1067);
xor U5136 (N_5136,In_1711,In_43);
xor U5137 (N_5137,In_978,In_1517);
nor U5138 (N_5138,In_498,In_573);
xor U5139 (N_5139,In_2889,In_1427);
or U5140 (N_5140,In_1004,In_1639);
nor U5141 (N_5141,In_2171,In_1948);
nor U5142 (N_5142,In_1055,In_2736);
nor U5143 (N_5143,In_1079,In_1318);
and U5144 (N_5144,In_1077,In_1137);
nor U5145 (N_5145,In_2529,In_1507);
and U5146 (N_5146,In_2414,In_29);
nor U5147 (N_5147,In_1722,In_2913);
or U5148 (N_5148,In_1095,In_1739);
xnor U5149 (N_5149,In_2548,In_17);
and U5150 (N_5150,In_1731,In_1937);
xnor U5151 (N_5151,In_1386,In_1246);
nor U5152 (N_5152,In_2960,In_2713);
xnor U5153 (N_5153,In_2101,In_1382);
and U5154 (N_5154,In_2969,In_976);
nand U5155 (N_5155,In_1739,In_2104);
xor U5156 (N_5156,In_2747,In_2878);
nand U5157 (N_5157,In_212,In_1695);
nor U5158 (N_5158,In_880,In_2704);
xnor U5159 (N_5159,In_572,In_2059);
nand U5160 (N_5160,In_1001,In_1773);
or U5161 (N_5161,In_174,In_2760);
nor U5162 (N_5162,In_120,In_1710);
or U5163 (N_5163,In_2444,In_1252);
or U5164 (N_5164,In_2941,In_811);
or U5165 (N_5165,In_1359,In_55);
nand U5166 (N_5166,In_2344,In_1285);
xor U5167 (N_5167,In_2151,In_2421);
nor U5168 (N_5168,In_74,In_1321);
and U5169 (N_5169,In_2388,In_139);
xor U5170 (N_5170,In_1507,In_2956);
nor U5171 (N_5171,In_2392,In_2350);
nand U5172 (N_5172,In_39,In_1526);
or U5173 (N_5173,In_1590,In_1385);
or U5174 (N_5174,In_1273,In_2524);
xnor U5175 (N_5175,In_1402,In_2681);
nor U5176 (N_5176,In_1537,In_2856);
nor U5177 (N_5177,In_2222,In_1566);
and U5178 (N_5178,In_2701,In_2659);
and U5179 (N_5179,In_1854,In_344);
xor U5180 (N_5180,In_2314,In_797);
and U5181 (N_5181,In_2979,In_290);
nor U5182 (N_5182,In_376,In_2623);
and U5183 (N_5183,In_1606,In_262);
nor U5184 (N_5184,In_659,In_166);
or U5185 (N_5185,In_2203,In_2282);
nor U5186 (N_5186,In_2553,In_1414);
nor U5187 (N_5187,In_1155,In_1754);
and U5188 (N_5188,In_1926,In_211);
and U5189 (N_5189,In_1723,In_763);
xnor U5190 (N_5190,In_1672,In_1688);
and U5191 (N_5191,In_2917,In_142);
and U5192 (N_5192,In_1116,In_261);
xor U5193 (N_5193,In_2740,In_267);
nand U5194 (N_5194,In_450,In_44);
nand U5195 (N_5195,In_288,In_1939);
and U5196 (N_5196,In_2467,In_2385);
nand U5197 (N_5197,In_188,In_850);
xor U5198 (N_5198,In_2017,In_838);
nor U5199 (N_5199,In_1808,In_2313);
or U5200 (N_5200,In_737,In_2508);
nor U5201 (N_5201,In_1028,In_2170);
nor U5202 (N_5202,In_2116,In_34);
nor U5203 (N_5203,In_2498,In_2708);
nand U5204 (N_5204,In_1564,In_2622);
xnor U5205 (N_5205,In_2282,In_475);
and U5206 (N_5206,In_1387,In_2517);
nor U5207 (N_5207,In_1101,In_1896);
or U5208 (N_5208,In_2777,In_903);
and U5209 (N_5209,In_994,In_770);
nor U5210 (N_5210,In_1160,In_1479);
xnor U5211 (N_5211,In_767,In_2910);
nand U5212 (N_5212,In_2946,In_2742);
and U5213 (N_5213,In_858,In_769);
or U5214 (N_5214,In_552,In_2670);
or U5215 (N_5215,In_456,In_2752);
nand U5216 (N_5216,In_1875,In_1538);
and U5217 (N_5217,In_2517,In_735);
nand U5218 (N_5218,In_2222,In_2838);
xor U5219 (N_5219,In_1349,In_1309);
xnor U5220 (N_5220,In_471,In_237);
or U5221 (N_5221,In_1773,In_1350);
nand U5222 (N_5222,In_2544,In_845);
and U5223 (N_5223,In_2471,In_2200);
nand U5224 (N_5224,In_1766,In_83);
and U5225 (N_5225,In_2857,In_501);
and U5226 (N_5226,In_910,In_1481);
nand U5227 (N_5227,In_1173,In_1259);
and U5228 (N_5228,In_231,In_2548);
xnor U5229 (N_5229,In_1259,In_283);
xnor U5230 (N_5230,In_720,In_1581);
and U5231 (N_5231,In_2263,In_2236);
xnor U5232 (N_5232,In_1947,In_2445);
nor U5233 (N_5233,In_780,In_27);
and U5234 (N_5234,In_2486,In_381);
xnor U5235 (N_5235,In_1655,In_1614);
xnor U5236 (N_5236,In_1784,In_2309);
xnor U5237 (N_5237,In_1580,In_2570);
nand U5238 (N_5238,In_2437,In_2604);
or U5239 (N_5239,In_222,In_1190);
xor U5240 (N_5240,In_1680,In_364);
and U5241 (N_5241,In_2866,In_1281);
xor U5242 (N_5242,In_2462,In_2338);
nor U5243 (N_5243,In_228,In_976);
nand U5244 (N_5244,In_1357,In_101);
and U5245 (N_5245,In_720,In_1684);
nor U5246 (N_5246,In_1379,In_2787);
xor U5247 (N_5247,In_2574,In_2512);
or U5248 (N_5248,In_2402,In_1311);
and U5249 (N_5249,In_1623,In_953);
or U5250 (N_5250,In_1671,In_1921);
nor U5251 (N_5251,In_598,In_2848);
and U5252 (N_5252,In_1730,In_1771);
nor U5253 (N_5253,In_532,In_2966);
nand U5254 (N_5254,In_1805,In_2674);
or U5255 (N_5255,In_986,In_1673);
nand U5256 (N_5256,In_2582,In_631);
and U5257 (N_5257,In_1573,In_2943);
and U5258 (N_5258,In_2560,In_311);
xor U5259 (N_5259,In_425,In_2972);
or U5260 (N_5260,In_1795,In_1095);
xnor U5261 (N_5261,In_1380,In_630);
and U5262 (N_5262,In_2805,In_740);
xor U5263 (N_5263,In_2067,In_1021);
and U5264 (N_5264,In_1586,In_2798);
or U5265 (N_5265,In_1802,In_1838);
or U5266 (N_5266,In_1439,In_1304);
and U5267 (N_5267,In_1353,In_2506);
or U5268 (N_5268,In_2469,In_1426);
nand U5269 (N_5269,In_1698,In_1453);
or U5270 (N_5270,In_1103,In_2254);
or U5271 (N_5271,In_385,In_1872);
and U5272 (N_5272,In_2083,In_2103);
xor U5273 (N_5273,In_1279,In_2733);
and U5274 (N_5274,In_416,In_2621);
or U5275 (N_5275,In_150,In_2159);
or U5276 (N_5276,In_952,In_896);
and U5277 (N_5277,In_2843,In_2242);
and U5278 (N_5278,In_1385,In_2482);
or U5279 (N_5279,In_1034,In_2491);
and U5280 (N_5280,In_2919,In_1198);
nand U5281 (N_5281,In_2001,In_2279);
nand U5282 (N_5282,In_1941,In_2243);
and U5283 (N_5283,In_1245,In_816);
nand U5284 (N_5284,In_692,In_1799);
or U5285 (N_5285,In_2354,In_1505);
nor U5286 (N_5286,In_2126,In_1921);
or U5287 (N_5287,In_1339,In_1571);
xor U5288 (N_5288,In_1662,In_1384);
nor U5289 (N_5289,In_2286,In_2114);
and U5290 (N_5290,In_389,In_950);
and U5291 (N_5291,In_2123,In_2149);
and U5292 (N_5292,In_2560,In_743);
nor U5293 (N_5293,In_74,In_2231);
nand U5294 (N_5294,In_2588,In_2614);
nand U5295 (N_5295,In_2156,In_120);
nor U5296 (N_5296,In_366,In_1129);
and U5297 (N_5297,In_1446,In_344);
or U5298 (N_5298,In_2978,In_2069);
and U5299 (N_5299,In_841,In_1762);
or U5300 (N_5300,In_2526,In_151);
and U5301 (N_5301,In_2092,In_547);
nor U5302 (N_5302,In_1394,In_2283);
and U5303 (N_5303,In_1001,In_104);
xnor U5304 (N_5304,In_2457,In_1396);
nand U5305 (N_5305,In_1485,In_1046);
nand U5306 (N_5306,In_74,In_2166);
or U5307 (N_5307,In_2465,In_2805);
and U5308 (N_5308,In_2881,In_402);
nand U5309 (N_5309,In_43,In_2260);
and U5310 (N_5310,In_829,In_876);
xnor U5311 (N_5311,In_693,In_1618);
nand U5312 (N_5312,In_2888,In_1653);
nor U5313 (N_5313,In_2216,In_2955);
and U5314 (N_5314,In_386,In_138);
nand U5315 (N_5315,In_1994,In_13);
nand U5316 (N_5316,In_2667,In_2355);
or U5317 (N_5317,In_1305,In_906);
xor U5318 (N_5318,In_16,In_1372);
or U5319 (N_5319,In_1816,In_2555);
xnor U5320 (N_5320,In_1008,In_2768);
xor U5321 (N_5321,In_38,In_1183);
and U5322 (N_5322,In_2676,In_2649);
nor U5323 (N_5323,In_2693,In_886);
nand U5324 (N_5324,In_1647,In_460);
nor U5325 (N_5325,In_1428,In_692);
and U5326 (N_5326,In_662,In_1553);
nand U5327 (N_5327,In_2000,In_2920);
xnor U5328 (N_5328,In_1642,In_2851);
xor U5329 (N_5329,In_855,In_2236);
or U5330 (N_5330,In_2469,In_1757);
nand U5331 (N_5331,In_1452,In_1854);
nand U5332 (N_5332,In_1268,In_328);
nand U5333 (N_5333,In_636,In_1064);
nor U5334 (N_5334,In_2148,In_1533);
or U5335 (N_5335,In_1562,In_623);
xnor U5336 (N_5336,In_2863,In_379);
nand U5337 (N_5337,In_2923,In_1027);
and U5338 (N_5338,In_2536,In_1042);
and U5339 (N_5339,In_871,In_704);
and U5340 (N_5340,In_258,In_531);
or U5341 (N_5341,In_1216,In_235);
nand U5342 (N_5342,In_2470,In_484);
and U5343 (N_5343,In_1646,In_1410);
nand U5344 (N_5344,In_2401,In_1736);
and U5345 (N_5345,In_2425,In_218);
and U5346 (N_5346,In_1841,In_1125);
or U5347 (N_5347,In_251,In_1001);
or U5348 (N_5348,In_712,In_2170);
nand U5349 (N_5349,In_2908,In_2971);
or U5350 (N_5350,In_2088,In_2806);
and U5351 (N_5351,In_1870,In_1036);
and U5352 (N_5352,In_1506,In_502);
and U5353 (N_5353,In_1890,In_2636);
nor U5354 (N_5354,In_1791,In_802);
and U5355 (N_5355,In_2154,In_2854);
or U5356 (N_5356,In_1533,In_2068);
or U5357 (N_5357,In_240,In_2498);
and U5358 (N_5358,In_1339,In_838);
xnor U5359 (N_5359,In_1705,In_568);
xnor U5360 (N_5360,In_2520,In_25);
nand U5361 (N_5361,In_2484,In_2060);
and U5362 (N_5362,In_701,In_562);
nor U5363 (N_5363,In_2072,In_2874);
or U5364 (N_5364,In_1895,In_754);
or U5365 (N_5365,In_2873,In_102);
nand U5366 (N_5366,In_385,In_2082);
and U5367 (N_5367,In_1563,In_208);
and U5368 (N_5368,In_2107,In_2684);
or U5369 (N_5369,In_2530,In_1383);
or U5370 (N_5370,In_931,In_249);
nand U5371 (N_5371,In_2538,In_1809);
nor U5372 (N_5372,In_275,In_2713);
xnor U5373 (N_5373,In_1990,In_574);
or U5374 (N_5374,In_2194,In_484);
xor U5375 (N_5375,In_196,In_429);
and U5376 (N_5376,In_1606,In_2388);
and U5377 (N_5377,In_2156,In_2503);
and U5378 (N_5378,In_2926,In_915);
or U5379 (N_5379,In_1422,In_2027);
nand U5380 (N_5380,In_2226,In_2503);
xor U5381 (N_5381,In_2625,In_2370);
xor U5382 (N_5382,In_107,In_1918);
nor U5383 (N_5383,In_649,In_566);
nor U5384 (N_5384,In_135,In_2566);
nand U5385 (N_5385,In_900,In_1066);
or U5386 (N_5386,In_2167,In_602);
or U5387 (N_5387,In_1574,In_1368);
and U5388 (N_5388,In_2950,In_1993);
nor U5389 (N_5389,In_1389,In_1849);
xor U5390 (N_5390,In_491,In_900);
xnor U5391 (N_5391,In_2681,In_1216);
or U5392 (N_5392,In_2818,In_2576);
nor U5393 (N_5393,In_2895,In_11);
nor U5394 (N_5394,In_495,In_350);
nand U5395 (N_5395,In_789,In_1435);
and U5396 (N_5396,In_2909,In_2731);
xnor U5397 (N_5397,In_341,In_220);
and U5398 (N_5398,In_190,In_1226);
and U5399 (N_5399,In_1189,In_2023);
xor U5400 (N_5400,In_281,In_1644);
nand U5401 (N_5401,In_2284,In_528);
xor U5402 (N_5402,In_1285,In_2396);
xnor U5403 (N_5403,In_498,In_833);
nor U5404 (N_5404,In_444,In_1719);
and U5405 (N_5405,In_1535,In_440);
nor U5406 (N_5406,In_2323,In_314);
nor U5407 (N_5407,In_1000,In_688);
and U5408 (N_5408,In_1275,In_2496);
nor U5409 (N_5409,In_203,In_2041);
or U5410 (N_5410,In_624,In_1384);
and U5411 (N_5411,In_30,In_1665);
xnor U5412 (N_5412,In_2972,In_2026);
xnor U5413 (N_5413,In_2845,In_1284);
or U5414 (N_5414,In_1314,In_1531);
xnor U5415 (N_5415,In_252,In_912);
nand U5416 (N_5416,In_2399,In_2421);
nand U5417 (N_5417,In_1695,In_2372);
nand U5418 (N_5418,In_1198,In_2766);
or U5419 (N_5419,In_1602,In_1185);
or U5420 (N_5420,In_173,In_495);
xor U5421 (N_5421,In_2157,In_2045);
or U5422 (N_5422,In_1216,In_465);
and U5423 (N_5423,In_2591,In_1700);
and U5424 (N_5424,In_2175,In_2869);
nand U5425 (N_5425,In_2527,In_177);
xnor U5426 (N_5426,In_1518,In_2424);
xnor U5427 (N_5427,In_2822,In_1488);
nand U5428 (N_5428,In_2596,In_2336);
nand U5429 (N_5429,In_2551,In_1678);
nand U5430 (N_5430,In_2223,In_319);
nor U5431 (N_5431,In_2883,In_2724);
nand U5432 (N_5432,In_410,In_176);
nor U5433 (N_5433,In_1282,In_1563);
nand U5434 (N_5434,In_1440,In_1296);
or U5435 (N_5435,In_2833,In_954);
or U5436 (N_5436,In_1537,In_1144);
nand U5437 (N_5437,In_439,In_922);
and U5438 (N_5438,In_1086,In_1960);
nor U5439 (N_5439,In_679,In_841);
xor U5440 (N_5440,In_1268,In_73);
xor U5441 (N_5441,In_1930,In_2664);
xor U5442 (N_5442,In_159,In_2554);
nor U5443 (N_5443,In_208,In_2706);
or U5444 (N_5444,In_2289,In_166);
and U5445 (N_5445,In_2107,In_726);
nand U5446 (N_5446,In_1004,In_732);
nand U5447 (N_5447,In_1234,In_1264);
xnor U5448 (N_5448,In_650,In_223);
nor U5449 (N_5449,In_2287,In_1768);
and U5450 (N_5450,In_2628,In_2603);
nor U5451 (N_5451,In_656,In_523);
or U5452 (N_5452,In_2151,In_2634);
and U5453 (N_5453,In_1122,In_2593);
nor U5454 (N_5454,In_341,In_2246);
and U5455 (N_5455,In_268,In_1024);
nand U5456 (N_5456,In_884,In_2107);
xnor U5457 (N_5457,In_1502,In_2523);
xor U5458 (N_5458,In_1113,In_2455);
or U5459 (N_5459,In_1979,In_874);
nor U5460 (N_5460,In_1683,In_497);
or U5461 (N_5461,In_2511,In_1354);
or U5462 (N_5462,In_2174,In_271);
xnor U5463 (N_5463,In_1400,In_2089);
nor U5464 (N_5464,In_2507,In_831);
or U5465 (N_5465,In_2081,In_1641);
and U5466 (N_5466,In_2481,In_2657);
nor U5467 (N_5467,In_1501,In_1358);
nand U5468 (N_5468,In_1325,In_82);
nand U5469 (N_5469,In_2607,In_66);
and U5470 (N_5470,In_1939,In_2940);
nand U5471 (N_5471,In_1838,In_1131);
xnor U5472 (N_5472,In_1439,In_1963);
or U5473 (N_5473,In_2008,In_820);
xor U5474 (N_5474,In_2222,In_1139);
xnor U5475 (N_5475,In_1381,In_2026);
and U5476 (N_5476,In_2753,In_358);
nand U5477 (N_5477,In_892,In_875);
and U5478 (N_5478,In_2412,In_497);
or U5479 (N_5479,In_1788,In_2830);
and U5480 (N_5480,In_1643,In_814);
xor U5481 (N_5481,In_1656,In_88);
xor U5482 (N_5482,In_710,In_1650);
nand U5483 (N_5483,In_882,In_1385);
and U5484 (N_5484,In_1850,In_764);
nand U5485 (N_5485,In_2495,In_180);
and U5486 (N_5486,In_1142,In_768);
and U5487 (N_5487,In_2979,In_590);
xor U5488 (N_5488,In_1412,In_1814);
xor U5489 (N_5489,In_344,In_1471);
and U5490 (N_5490,In_1000,In_784);
xnor U5491 (N_5491,In_1937,In_480);
and U5492 (N_5492,In_2851,In_790);
xnor U5493 (N_5493,In_1008,In_323);
or U5494 (N_5494,In_284,In_253);
nor U5495 (N_5495,In_168,In_1407);
or U5496 (N_5496,In_1474,In_1856);
or U5497 (N_5497,In_2113,In_1084);
nor U5498 (N_5498,In_2033,In_1731);
and U5499 (N_5499,In_235,In_1744);
nor U5500 (N_5500,In_546,In_1032);
xor U5501 (N_5501,In_1148,In_56);
or U5502 (N_5502,In_2548,In_2257);
nor U5503 (N_5503,In_2215,In_927);
or U5504 (N_5504,In_764,In_57);
or U5505 (N_5505,In_2787,In_171);
xnor U5506 (N_5506,In_317,In_1520);
nand U5507 (N_5507,In_354,In_2457);
nand U5508 (N_5508,In_1454,In_2957);
nand U5509 (N_5509,In_891,In_542);
and U5510 (N_5510,In_451,In_29);
xor U5511 (N_5511,In_2549,In_1369);
and U5512 (N_5512,In_2463,In_318);
or U5513 (N_5513,In_883,In_2601);
nand U5514 (N_5514,In_959,In_1909);
xor U5515 (N_5515,In_2261,In_235);
and U5516 (N_5516,In_1733,In_62);
and U5517 (N_5517,In_362,In_2171);
and U5518 (N_5518,In_2187,In_1406);
and U5519 (N_5519,In_733,In_2556);
or U5520 (N_5520,In_1610,In_1576);
nor U5521 (N_5521,In_1877,In_1067);
and U5522 (N_5522,In_2741,In_503);
xor U5523 (N_5523,In_2623,In_990);
and U5524 (N_5524,In_978,In_1988);
or U5525 (N_5525,In_2466,In_839);
nor U5526 (N_5526,In_2809,In_818);
and U5527 (N_5527,In_2238,In_415);
or U5528 (N_5528,In_1589,In_929);
nor U5529 (N_5529,In_2181,In_124);
and U5530 (N_5530,In_2314,In_2288);
or U5531 (N_5531,In_2162,In_2342);
nor U5532 (N_5532,In_2548,In_2456);
or U5533 (N_5533,In_1704,In_1744);
nor U5534 (N_5534,In_706,In_889);
and U5535 (N_5535,In_833,In_271);
nor U5536 (N_5536,In_1523,In_1056);
xnor U5537 (N_5537,In_2321,In_385);
nor U5538 (N_5538,In_2012,In_2188);
or U5539 (N_5539,In_1183,In_610);
nand U5540 (N_5540,In_1071,In_112);
xor U5541 (N_5541,In_1641,In_798);
or U5542 (N_5542,In_961,In_1208);
xnor U5543 (N_5543,In_565,In_2309);
or U5544 (N_5544,In_1970,In_8);
nor U5545 (N_5545,In_1018,In_30);
and U5546 (N_5546,In_2173,In_2685);
or U5547 (N_5547,In_863,In_2267);
nor U5548 (N_5548,In_1330,In_1927);
nand U5549 (N_5549,In_1486,In_2423);
nand U5550 (N_5550,In_2627,In_2734);
nand U5551 (N_5551,In_717,In_258);
nor U5552 (N_5552,In_1848,In_784);
nor U5553 (N_5553,In_1927,In_190);
nand U5554 (N_5554,In_1252,In_58);
and U5555 (N_5555,In_654,In_223);
and U5556 (N_5556,In_1092,In_2964);
and U5557 (N_5557,In_1555,In_493);
or U5558 (N_5558,In_1577,In_2463);
or U5559 (N_5559,In_376,In_1956);
and U5560 (N_5560,In_267,In_853);
or U5561 (N_5561,In_108,In_580);
or U5562 (N_5562,In_2188,In_2213);
or U5563 (N_5563,In_666,In_137);
xor U5564 (N_5564,In_1574,In_1556);
or U5565 (N_5565,In_1187,In_2815);
nand U5566 (N_5566,In_858,In_1055);
and U5567 (N_5567,In_1138,In_2771);
and U5568 (N_5568,In_821,In_856);
or U5569 (N_5569,In_1646,In_1325);
nand U5570 (N_5570,In_2726,In_2949);
and U5571 (N_5571,In_2540,In_107);
nand U5572 (N_5572,In_773,In_2895);
or U5573 (N_5573,In_1883,In_2269);
or U5574 (N_5574,In_2610,In_2351);
or U5575 (N_5575,In_1658,In_2676);
nor U5576 (N_5576,In_1177,In_719);
and U5577 (N_5577,In_2658,In_1403);
and U5578 (N_5578,In_99,In_2375);
nand U5579 (N_5579,In_1836,In_86);
or U5580 (N_5580,In_2455,In_1919);
and U5581 (N_5581,In_2074,In_391);
xnor U5582 (N_5582,In_497,In_1416);
nor U5583 (N_5583,In_1263,In_1279);
or U5584 (N_5584,In_1377,In_1120);
nand U5585 (N_5585,In_2866,In_127);
or U5586 (N_5586,In_2314,In_1849);
nand U5587 (N_5587,In_413,In_2777);
or U5588 (N_5588,In_2259,In_1254);
or U5589 (N_5589,In_1105,In_207);
nor U5590 (N_5590,In_2176,In_2829);
nand U5591 (N_5591,In_1420,In_2610);
and U5592 (N_5592,In_1392,In_2861);
and U5593 (N_5593,In_2145,In_1759);
or U5594 (N_5594,In_1401,In_2399);
nor U5595 (N_5595,In_1690,In_872);
xnor U5596 (N_5596,In_1801,In_1193);
nor U5597 (N_5597,In_892,In_1933);
or U5598 (N_5598,In_1141,In_657);
xnor U5599 (N_5599,In_2905,In_2589);
and U5600 (N_5600,In_414,In_442);
xnor U5601 (N_5601,In_1689,In_179);
xnor U5602 (N_5602,In_2805,In_2423);
and U5603 (N_5603,In_1926,In_1048);
xor U5604 (N_5604,In_66,In_2289);
or U5605 (N_5605,In_486,In_1352);
nor U5606 (N_5606,In_1163,In_1780);
nand U5607 (N_5607,In_148,In_423);
xor U5608 (N_5608,In_1557,In_505);
nor U5609 (N_5609,In_2583,In_2662);
nor U5610 (N_5610,In_886,In_918);
nand U5611 (N_5611,In_1829,In_868);
xor U5612 (N_5612,In_144,In_371);
nor U5613 (N_5613,In_2947,In_287);
and U5614 (N_5614,In_2017,In_486);
nand U5615 (N_5615,In_2254,In_2948);
or U5616 (N_5616,In_2263,In_1252);
xnor U5617 (N_5617,In_1714,In_1053);
nor U5618 (N_5618,In_2225,In_2202);
or U5619 (N_5619,In_88,In_2453);
and U5620 (N_5620,In_2049,In_208);
or U5621 (N_5621,In_340,In_1906);
xnor U5622 (N_5622,In_7,In_618);
and U5623 (N_5623,In_1121,In_2735);
or U5624 (N_5624,In_318,In_1608);
nor U5625 (N_5625,In_2500,In_1175);
xor U5626 (N_5626,In_779,In_2642);
and U5627 (N_5627,In_2815,In_1435);
nor U5628 (N_5628,In_1970,In_2074);
xor U5629 (N_5629,In_595,In_2238);
nor U5630 (N_5630,In_2290,In_1);
and U5631 (N_5631,In_2549,In_768);
xor U5632 (N_5632,In_2415,In_851);
nor U5633 (N_5633,In_1099,In_2296);
and U5634 (N_5634,In_1723,In_30);
or U5635 (N_5635,In_2408,In_802);
nor U5636 (N_5636,In_690,In_911);
nor U5637 (N_5637,In_2420,In_327);
or U5638 (N_5638,In_2764,In_2214);
nor U5639 (N_5639,In_2563,In_1367);
nor U5640 (N_5640,In_879,In_2135);
nor U5641 (N_5641,In_975,In_277);
and U5642 (N_5642,In_464,In_2773);
nor U5643 (N_5643,In_2185,In_2780);
nor U5644 (N_5644,In_1261,In_2095);
nor U5645 (N_5645,In_1199,In_2156);
xnor U5646 (N_5646,In_1815,In_1244);
and U5647 (N_5647,In_244,In_1957);
xor U5648 (N_5648,In_2869,In_1746);
nand U5649 (N_5649,In_902,In_2273);
or U5650 (N_5650,In_291,In_689);
and U5651 (N_5651,In_1274,In_111);
and U5652 (N_5652,In_108,In_2272);
xnor U5653 (N_5653,In_415,In_1091);
nand U5654 (N_5654,In_1334,In_300);
or U5655 (N_5655,In_1747,In_1057);
nand U5656 (N_5656,In_1347,In_997);
nor U5657 (N_5657,In_843,In_401);
and U5658 (N_5658,In_372,In_2928);
or U5659 (N_5659,In_1776,In_2144);
nor U5660 (N_5660,In_806,In_1344);
xor U5661 (N_5661,In_1768,In_610);
or U5662 (N_5662,In_686,In_113);
or U5663 (N_5663,In_1226,In_2097);
or U5664 (N_5664,In_2401,In_209);
or U5665 (N_5665,In_2758,In_2336);
nand U5666 (N_5666,In_816,In_1441);
xnor U5667 (N_5667,In_1316,In_2818);
xor U5668 (N_5668,In_1046,In_1482);
and U5669 (N_5669,In_2889,In_2716);
nor U5670 (N_5670,In_466,In_845);
and U5671 (N_5671,In_2032,In_2912);
nor U5672 (N_5672,In_1717,In_1430);
nand U5673 (N_5673,In_761,In_1492);
xor U5674 (N_5674,In_932,In_297);
xnor U5675 (N_5675,In_2834,In_1751);
and U5676 (N_5676,In_1903,In_51);
nor U5677 (N_5677,In_217,In_460);
and U5678 (N_5678,In_2463,In_1714);
or U5679 (N_5679,In_1539,In_1065);
xnor U5680 (N_5680,In_2136,In_1934);
xor U5681 (N_5681,In_600,In_765);
nand U5682 (N_5682,In_2551,In_2105);
nor U5683 (N_5683,In_908,In_1515);
and U5684 (N_5684,In_1704,In_1802);
nand U5685 (N_5685,In_2195,In_103);
and U5686 (N_5686,In_835,In_898);
xor U5687 (N_5687,In_854,In_84);
nand U5688 (N_5688,In_2449,In_256);
or U5689 (N_5689,In_523,In_833);
xor U5690 (N_5690,In_2600,In_1528);
nor U5691 (N_5691,In_1583,In_1244);
nand U5692 (N_5692,In_2244,In_1683);
xnor U5693 (N_5693,In_2738,In_2274);
nand U5694 (N_5694,In_488,In_1008);
or U5695 (N_5695,In_539,In_1608);
nand U5696 (N_5696,In_143,In_1970);
nor U5697 (N_5697,In_16,In_1593);
or U5698 (N_5698,In_2074,In_2329);
and U5699 (N_5699,In_573,In_2009);
and U5700 (N_5700,In_2195,In_1180);
or U5701 (N_5701,In_2289,In_289);
and U5702 (N_5702,In_1005,In_2701);
and U5703 (N_5703,In_2887,In_132);
and U5704 (N_5704,In_636,In_348);
nor U5705 (N_5705,In_710,In_913);
nor U5706 (N_5706,In_2167,In_2493);
or U5707 (N_5707,In_1890,In_1667);
or U5708 (N_5708,In_2689,In_538);
nor U5709 (N_5709,In_2483,In_776);
nor U5710 (N_5710,In_962,In_2012);
nand U5711 (N_5711,In_1283,In_999);
and U5712 (N_5712,In_1547,In_2271);
xor U5713 (N_5713,In_1555,In_1714);
and U5714 (N_5714,In_2507,In_134);
xor U5715 (N_5715,In_2482,In_1341);
nand U5716 (N_5716,In_1635,In_2572);
xnor U5717 (N_5717,In_1699,In_1720);
or U5718 (N_5718,In_800,In_1478);
xnor U5719 (N_5719,In_2302,In_2012);
xnor U5720 (N_5720,In_180,In_1987);
or U5721 (N_5721,In_160,In_102);
and U5722 (N_5722,In_1857,In_2366);
nor U5723 (N_5723,In_1367,In_386);
nand U5724 (N_5724,In_806,In_2972);
xnor U5725 (N_5725,In_1636,In_173);
nand U5726 (N_5726,In_2127,In_839);
and U5727 (N_5727,In_206,In_1601);
nor U5728 (N_5728,In_859,In_234);
or U5729 (N_5729,In_2911,In_2722);
xor U5730 (N_5730,In_2627,In_2750);
nor U5731 (N_5731,In_2820,In_569);
nor U5732 (N_5732,In_2314,In_1871);
nand U5733 (N_5733,In_2902,In_1016);
xnor U5734 (N_5734,In_2194,In_1400);
xnor U5735 (N_5735,In_1503,In_2863);
and U5736 (N_5736,In_2068,In_1451);
xor U5737 (N_5737,In_2154,In_2055);
nor U5738 (N_5738,In_2371,In_2958);
nand U5739 (N_5739,In_2984,In_622);
and U5740 (N_5740,In_2024,In_487);
or U5741 (N_5741,In_288,In_2508);
or U5742 (N_5742,In_1389,In_1099);
nand U5743 (N_5743,In_1321,In_868);
nand U5744 (N_5744,In_1373,In_1898);
and U5745 (N_5745,In_440,In_2216);
and U5746 (N_5746,In_261,In_2850);
or U5747 (N_5747,In_1138,In_402);
xor U5748 (N_5748,In_2525,In_61);
or U5749 (N_5749,In_1041,In_1082);
and U5750 (N_5750,In_2639,In_2107);
xor U5751 (N_5751,In_1724,In_460);
and U5752 (N_5752,In_828,In_321);
nand U5753 (N_5753,In_266,In_1521);
and U5754 (N_5754,In_2811,In_697);
or U5755 (N_5755,In_1738,In_571);
or U5756 (N_5756,In_1120,In_62);
nor U5757 (N_5757,In_1254,In_2844);
nand U5758 (N_5758,In_1607,In_2913);
nor U5759 (N_5759,In_1832,In_592);
or U5760 (N_5760,In_517,In_1490);
nand U5761 (N_5761,In_218,In_1947);
nand U5762 (N_5762,In_45,In_2392);
nand U5763 (N_5763,In_1843,In_2704);
nand U5764 (N_5764,In_2058,In_2513);
nand U5765 (N_5765,In_2146,In_1994);
xnor U5766 (N_5766,In_690,In_844);
nand U5767 (N_5767,In_433,In_536);
xnor U5768 (N_5768,In_1625,In_198);
nand U5769 (N_5769,In_1884,In_1484);
or U5770 (N_5770,In_2243,In_2496);
xor U5771 (N_5771,In_2554,In_1486);
and U5772 (N_5772,In_2369,In_452);
xor U5773 (N_5773,In_2044,In_663);
nor U5774 (N_5774,In_78,In_2428);
and U5775 (N_5775,In_756,In_1658);
and U5776 (N_5776,In_2370,In_791);
and U5777 (N_5777,In_2063,In_752);
nor U5778 (N_5778,In_794,In_1440);
nor U5779 (N_5779,In_2818,In_1195);
nor U5780 (N_5780,In_1629,In_854);
nor U5781 (N_5781,In_2341,In_1123);
and U5782 (N_5782,In_1675,In_1644);
nor U5783 (N_5783,In_2395,In_432);
xor U5784 (N_5784,In_354,In_1267);
or U5785 (N_5785,In_709,In_860);
nor U5786 (N_5786,In_1973,In_1656);
xor U5787 (N_5787,In_501,In_1768);
nand U5788 (N_5788,In_113,In_1515);
nand U5789 (N_5789,In_613,In_835);
nor U5790 (N_5790,In_976,In_1016);
and U5791 (N_5791,In_1667,In_2361);
xnor U5792 (N_5792,In_1179,In_18);
nand U5793 (N_5793,In_2967,In_1753);
nand U5794 (N_5794,In_2275,In_112);
nor U5795 (N_5795,In_2233,In_637);
or U5796 (N_5796,In_2233,In_1604);
nor U5797 (N_5797,In_1456,In_1848);
nor U5798 (N_5798,In_1355,In_27);
nand U5799 (N_5799,In_673,In_608);
and U5800 (N_5800,In_321,In_450);
nor U5801 (N_5801,In_868,In_2627);
xnor U5802 (N_5802,In_1490,In_1470);
nor U5803 (N_5803,In_1508,In_1371);
xor U5804 (N_5804,In_2016,In_1739);
nand U5805 (N_5805,In_116,In_2335);
xnor U5806 (N_5806,In_2791,In_2549);
xor U5807 (N_5807,In_2206,In_2019);
or U5808 (N_5808,In_1559,In_1775);
xnor U5809 (N_5809,In_2288,In_1300);
and U5810 (N_5810,In_465,In_1390);
or U5811 (N_5811,In_2267,In_1571);
and U5812 (N_5812,In_94,In_2289);
and U5813 (N_5813,In_1858,In_1917);
or U5814 (N_5814,In_400,In_2448);
and U5815 (N_5815,In_2190,In_750);
nand U5816 (N_5816,In_285,In_827);
nor U5817 (N_5817,In_1157,In_1714);
nor U5818 (N_5818,In_967,In_1561);
and U5819 (N_5819,In_2601,In_221);
or U5820 (N_5820,In_2311,In_1319);
or U5821 (N_5821,In_483,In_690);
xor U5822 (N_5822,In_2093,In_698);
or U5823 (N_5823,In_2129,In_2961);
and U5824 (N_5824,In_1532,In_1318);
nor U5825 (N_5825,In_1823,In_1120);
xor U5826 (N_5826,In_1514,In_540);
xnor U5827 (N_5827,In_2075,In_280);
and U5828 (N_5828,In_2920,In_542);
or U5829 (N_5829,In_2199,In_2519);
and U5830 (N_5830,In_499,In_2418);
xor U5831 (N_5831,In_2173,In_1434);
nor U5832 (N_5832,In_2731,In_2338);
nor U5833 (N_5833,In_426,In_2297);
or U5834 (N_5834,In_136,In_2786);
or U5835 (N_5835,In_916,In_214);
or U5836 (N_5836,In_1063,In_2385);
nor U5837 (N_5837,In_1987,In_2193);
and U5838 (N_5838,In_1958,In_518);
and U5839 (N_5839,In_2882,In_277);
and U5840 (N_5840,In_1540,In_2724);
nor U5841 (N_5841,In_72,In_26);
and U5842 (N_5842,In_1776,In_1313);
or U5843 (N_5843,In_2856,In_796);
xor U5844 (N_5844,In_2758,In_1103);
and U5845 (N_5845,In_1409,In_2381);
and U5846 (N_5846,In_154,In_2525);
or U5847 (N_5847,In_1904,In_675);
and U5848 (N_5848,In_2317,In_931);
or U5849 (N_5849,In_1321,In_2108);
and U5850 (N_5850,In_1969,In_2464);
and U5851 (N_5851,In_1789,In_850);
and U5852 (N_5852,In_2201,In_1088);
nor U5853 (N_5853,In_1848,In_524);
xor U5854 (N_5854,In_869,In_434);
xnor U5855 (N_5855,In_1532,In_265);
nand U5856 (N_5856,In_2892,In_953);
xor U5857 (N_5857,In_1743,In_1461);
xnor U5858 (N_5858,In_2306,In_1722);
or U5859 (N_5859,In_1652,In_2715);
or U5860 (N_5860,In_2163,In_46);
and U5861 (N_5861,In_2271,In_1341);
nor U5862 (N_5862,In_1842,In_1939);
xnor U5863 (N_5863,In_193,In_1121);
nor U5864 (N_5864,In_558,In_133);
xnor U5865 (N_5865,In_2598,In_1590);
or U5866 (N_5866,In_1563,In_47);
xnor U5867 (N_5867,In_2872,In_1519);
xor U5868 (N_5868,In_1472,In_2089);
nor U5869 (N_5869,In_2011,In_920);
nand U5870 (N_5870,In_1827,In_1565);
and U5871 (N_5871,In_361,In_1791);
and U5872 (N_5872,In_2976,In_264);
xor U5873 (N_5873,In_1021,In_2367);
xor U5874 (N_5874,In_2177,In_962);
nor U5875 (N_5875,In_1564,In_1045);
nand U5876 (N_5876,In_2075,In_1714);
nand U5877 (N_5877,In_2476,In_344);
nor U5878 (N_5878,In_1983,In_487);
nor U5879 (N_5879,In_664,In_126);
nor U5880 (N_5880,In_1127,In_2816);
nand U5881 (N_5881,In_2557,In_2203);
xor U5882 (N_5882,In_1099,In_2902);
and U5883 (N_5883,In_1422,In_1074);
and U5884 (N_5884,In_1754,In_2586);
nand U5885 (N_5885,In_1212,In_1253);
and U5886 (N_5886,In_27,In_2852);
nor U5887 (N_5887,In_1530,In_1209);
nand U5888 (N_5888,In_2204,In_902);
or U5889 (N_5889,In_1838,In_2884);
nand U5890 (N_5890,In_2887,In_325);
xor U5891 (N_5891,In_901,In_2681);
nor U5892 (N_5892,In_1185,In_2859);
and U5893 (N_5893,In_2566,In_614);
and U5894 (N_5894,In_2373,In_392);
nor U5895 (N_5895,In_1431,In_1554);
or U5896 (N_5896,In_831,In_2108);
xnor U5897 (N_5897,In_1858,In_493);
or U5898 (N_5898,In_2049,In_1927);
nand U5899 (N_5899,In_312,In_1976);
or U5900 (N_5900,In_1488,In_434);
nor U5901 (N_5901,In_2182,In_2073);
xor U5902 (N_5902,In_2828,In_522);
xnor U5903 (N_5903,In_619,In_2760);
nor U5904 (N_5904,In_2921,In_502);
xnor U5905 (N_5905,In_2562,In_2551);
xnor U5906 (N_5906,In_2770,In_2613);
xnor U5907 (N_5907,In_947,In_950);
nor U5908 (N_5908,In_87,In_1241);
nand U5909 (N_5909,In_2294,In_2469);
and U5910 (N_5910,In_843,In_1875);
nor U5911 (N_5911,In_77,In_2643);
xnor U5912 (N_5912,In_220,In_2425);
nor U5913 (N_5913,In_1907,In_1083);
nand U5914 (N_5914,In_459,In_1205);
or U5915 (N_5915,In_1698,In_1083);
xnor U5916 (N_5916,In_2872,In_1736);
nor U5917 (N_5917,In_194,In_1988);
xor U5918 (N_5918,In_839,In_2156);
nand U5919 (N_5919,In_2584,In_846);
and U5920 (N_5920,In_703,In_843);
nand U5921 (N_5921,In_854,In_380);
or U5922 (N_5922,In_1417,In_1402);
and U5923 (N_5923,In_2379,In_1257);
and U5924 (N_5924,In_621,In_1663);
nand U5925 (N_5925,In_2042,In_1871);
or U5926 (N_5926,In_708,In_1087);
nor U5927 (N_5927,In_2276,In_1334);
nor U5928 (N_5928,In_2838,In_2144);
or U5929 (N_5929,In_1756,In_2011);
and U5930 (N_5930,In_2687,In_1732);
nor U5931 (N_5931,In_1003,In_70);
and U5932 (N_5932,In_2842,In_1450);
and U5933 (N_5933,In_2276,In_216);
nand U5934 (N_5934,In_1493,In_2430);
and U5935 (N_5935,In_2833,In_1220);
or U5936 (N_5936,In_2507,In_1118);
or U5937 (N_5937,In_1880,In_1712);
or U5938 (N_5938,In_2315,In_1190);
nand U5939 (N_5939,In_1103,In_1460);
nor U5940 (N_5940,In_454,In_1971);
nand U5941 (N_5941,In_1115,In_193);
nor U5942 (N_5942,In_165,In_2639);
nand U5943 (N_5943,In_601,In_192);
or U5944 (N_5944,In_718,In_1799);
xor U5945 (N_5945,In_2361,In_2562);
and U5946 (N_5946,In_2605,In_2233);
or U5947 (N_5947,In_680,In_1242);
nor U5948 (N_5948,In_87,In_1653);
nand U5949 (N_5949,In_182,In_2010);
xor U5950 (N_5950,In_1681,In_1095);
nand U5951 (N_5951,In_2906,In_117);
nor U5952 (N_5952,In_1302,In_2265);
xnor U5953 (N_5953,In_1544,In_1381);
nand U5954 (N_5954,In_2333,In_2381);
or U5955 (N_5955,In_499,In_787);
nand U5956 (N_5956,In_697,In_1890);
xor U5957 (N_5957,In_2671,In_848);
nor U5958 (N_5958,In_2597,In_931);
nand U5959 (N_5959,In_950,In_1258);
nor U5960 (N_5960,In_2290,In_348);
or U5961 (N_5961,In_950,In_2319);
nor U5962 (N_5962,In_154,In_1043);
or U5963 (N_5963,In_1617,In_1291);
nand U5964 (N_5964,In_76,In_231);
nor U5965 (N_5965,In_1942,In_746);
nor U5966 (N_5966,In_244,In_1284);
xnor U5967 (N_5967,In_1731,In_2523);
nor U5968 (N_5968,In_1752,In_1654);
nor U5969 (N_5969,In_2189,In_87);
nand U5970 (N_5970,In_2516,In_2595);
nand U5971 (N_5971,In_1180,In_711);
and U5972 (N_5972,In_2568,In_23);
nand U5973 (N_5973,In_2486,In_1372);
nand U5974 (N_5974,In_1181,In_2592);
or U5975 (N_5975,In_836,In_2893);
nor U5976 (N_5976,In_2917,In_1807);
nand U5977 (N_5977,In_1694,In_2748);
nor U5978 (N_5978,In_671,In_2508);
or U5979 (N_5979,In_2201,In_2642);
and U5980 (N_5980,In_2792,In_1997);
nand U5981 (N_5981,In_1999,In_2982);
and U5982 (N_5982,In_1502,In_872);
nand U5983 (N_5983,In_1510,In_121);
nand U5984 (N_5984,In_1800,In_1504);
or U5985 (N_5985,In_2585,In_2808);
nand U5986 (N_5986,In_2282,In_1884);
nor U5987 (N_5987,In_322,In_1154);
or U5988 (N_5988,In_462,In_1233);
xor U5989 (N_5989,In_380,In_332);
nor U5990 (N_5990,In_2442,In_363);
nor U5991 (N_5991,In_2103,In_2918);
xor U5992 (N_5992,In_514,In_2637);
or U5993 (N_5993,In_2069,In_1956);
and U5994 (N_5994,In_2846,In_714);
nor U5995 (N_5995,In_1087,In_1907);
nor U5996 (N_5996,In_970,In_2492);
nor U5997 (N_5997,In_2626,In_299);
and U5998 (N_5998,In_2613,In_1983);
and U5999 (N_5999,In_281,In_399);
and U6000 (N_6000,N_2915,N_3773);
nand U6001 (N_6001,N_5518,N_5388);
nor U6002 (N_6002,N_5231,N_3612);
or U6003 (N_6003,N_3272,N_4930);
nand U6004 (N_6004,N_2424,N_741);
xnor U6005 (N_6005,N_334,N_4120);
or U6006 (N_6006,N_1573,N_5995);
nor U6007 (N_6007,N_4287,N_302);
and U6008 (N_6008,N_1193,N_1532);
and U6009 (N_6009,N_766,N_3838);
xor U6010 (N_6010,N_221,N_269);
xnor U6011 (N_6011,N_3069,N_5959);
or U6012 (N_6012,N_2907,N_2906);
and U6013 (N_6013,N_3168,N_1274);
nor U6014 (N_6014,N_3389,N_1671);
nand U6015 (N_6015,N_5200,N_4663);
nor U6016 (N_6016,N_4311,N_1004);
and U6017 (N_6017,N_4366,N_73);
or U6018 (N_6018,N_3932,N_465);
xnor U6019 (N_6019,N_1826,N_5536);
nand U6020 (N_6020,N_950,N_1798);
and U6021 (N_6021,N_3712,N_831);
nand U6022 (N_6022,N_644,N_2607);
nor U6023 (N_6023,N_4561,N_4625);
nand U6024 (N_6024,N_5177,N_3258);
and U6025 (N_6025,N_1737,N_354);
xnor U6026 (N_6026,N_3697,N_2379);
or U6027 (N_6027,N_419,N_5159);
or U6028 (N_6028,N_1149,N_3792);
nor U6029 (N_6029,N_3294,N_1281);
and U6030 (N_6030,N_3056,N_3031);
and U6031 (N_6031,N_117,N_1621);
or U6032 (N_6032,N_3666,N_725);
nand U6033 (N_6033,N_1914,N_518);
or U6034 (N_6034,N_2034,N_1981);
nand U6035 (N_6035,N_5358,N_5857);
or U6036 (N_6036,N_49,N_5769);
and U6037 (N_6037,N_4227,N_2478);
nand U6038 (N_6038,N_4341,N_413);
xnor U6039 (N_6039,N_4602,N_2974);
nor U6040 (N_6040,N_2949,N_296);
xor U6041 (N_6041,N_1039,N_3300);
xnor U6042 (N_6042,N_5607,N_29);
nand U6043 (N_6043,N_245,N_4749);
or U6044 (N_6044,N_3109,N_5268);
and U6045 (N_6045,N_1369,N_5160);
nand U6046 (N_6046,N_5026,N_5611);
nand U6047 (N_6047,N_3367,N_832);
and U6048 (N_6048,N_1508,N_4556);
nand U6049 (N_6049,N_2099,N_1044);
and U6050 (N_6050,N_5736,N_5529);
nand U6051 (N_6051,N_2246,N_2313);
and U6052 (N_6052,N_4989,N_349);
or U6053 (N_6053,N_1611,N_5632);
xnor U6054 (N_6054,N_861,N_1427);
nand U6055 (N_6055,N_1748,N_1591);
or U6056 (N_6056,N_1645,N_2914);
and U6057 (N_6057,N_4736,N_1046);
xnor U6058 (N_6058,N_732,N_1372);
or U6059 (N_6059,N_3671,N_4442);
nand U6060 (N_6060,N_2315,N_3581);
and U6061 (N_6061,N_415,N_2119);
nor U6062 (N_6062,N_2941,N_4215);
xor U6063 (N_6063,N_2882,N_4462);
or U6064 (N_6064,N_4002,N_4516);
and U6065 (N_6065,N_5920,N_4975);
nand U6066 (N_6066,N_5092,N_772);
or U6067 (N_6067,N_1391,N_712);
nor U6068 (N_6068,N_1343,N_4844);
and U6069 (N_6069,N_693,N_4134);
and U6070 (N_6070,N_4780,N_1927);
or U6071 (N_6071,N_1416,N_1505);
nand U6072 (N_6072,N_5139,N_5561);
nor U6073 (N_6073,N_1772,N_2171);
nor U6074 (N_6074,N_3055,N_2999);
nand U6075 (N_6075,N_5773,N_3394);
nand U6076 (N_6076,N_134,N_3079);
xor U6077 (N_6077,N_5605,N_3696);
xnor U6078 (N_6078,N_781,N_1992);
or U6079 (N_6079,N_1426,N_4132);
nand U6080 (N_6080,N_3788,N_2748);
nor U6081 (N_6081,N_2660,N_513);
nor U6082 (N_6082,N_3165,N_1523);
or U6083 (N_6083,N_5306,N_1052);
nand U6084 (N_6084,N_408,N_1098);
nor U6085 (N_6085,N_913,N_3372);
xnor U6086 (N_6086,N_1673,N_1678);
nor U6087 (N_6087,N_2729,N_577);
or U6088 (N_6088,N_155,N_2904);
nor U6089 (N_6089,N_3014,N_181);
nor U6090 (N_6090,N_4440,N_2816);
or U6091 (N_6091,N_5325,N_676);
nor U6092 (N_6092,N_5712,N_78);
and U6093 (N_6093,N_5861,N_1395);
nor U6094 (N_6094,N_3204,N_1447);
and U6095 (N_6095,N_864,N_5292);
nand U6096 (N_6096,N_4347,N_4138);
and U6097 (N_6097,N_850,N_1531);
xor U6098 (N_6098,N_5474,N_3175);
or U6099 (N_6099,N_2429,N_651);
nor U6100 (N_6100,N_640,N_2516);
xnor U6101 (N_6101,N_3002,N_3116);
xnor U6102 (N_6102,N_5706,N_530);
nor U6103 (N_6103,N_3340,N_1928);
and U6104 (N_6104,N_4616,N_2537);
xnor U6105 (N_6105,N_2322,N_4713);
or U6106 (N_6106,N_1939,N_3929);
or U6107 (N_6107,N_1709,N_213);
xnor U6108 (N_6108,N_2704,N_2262);
xor U6109 (N_6109,N_4517,N_2894);
nor U6110 (N_6110,N_4093,N_873);
and U6111 (N_6111,N_5310,N_5990);
xnor U6112 (N_6112,N_5244,N_4340);
nand U6113 (N_6113,N_3651,N_2370);
nand U6114 (N_6114,N_880,N_4637);
or U6115 (N_6115,N_343,N_2659);
xnor U6116 (N_6116,N_4084,N_1490);
and U6117 (N_6117,N_2445,N_4251);
nor U6118 (N_6118,N_249,N_1830);
or U6119 (N_6119,N_297,N_309);
and U6120 (N_6120,N_5431,N_5707);
xor U6121 (N_6121,N_1997,N_5994);
nand U6122 (N_6122,N_2554,N_1225);
xnor U6123 (N_6123,N_2135,N_4902);
and U6124 (N_6124,N_339,N_409);
nand U6125 (N_6125,N_3802,N_5782);
or U6126 (N_6126,N_3660,N_5692);
xor U6127 (N_6127,N_5441,N_4451);
xnor U6128 (N_6128,N_1493,N_546);
nor U6129 (N_6129,N_4004,N_4995);
xnor U6130 (N_6130,N_4784,N_4789);
xor U6131 (N_6131,N_4095,N_234);
or U6132 (N_6132,N_5524,N_1796);
xor U6133 (N_6133,N_737,N_2721);
nor U6134 (N_6134,N_188,N_556);
nor U6135 (N_6135,N_5223,N_847);
and U6136 (N_6136,N_4015,N_822);
xnor U6137 (N_6137,N_5479,N_3267);
nor U6138 (N_6138,N_939,N_5364);
or U6139 (N_6139,N_1326,N_3829);
nand U6140 (N_6140,N_3642,N_3879);
nand U6141 (N_6141,N_4179,N_2337);
or U6142 (N_6142,N_5229,N_3713);
or U6143 (N_6143,N_799,N_3661);
xnor U6144 (N_6144,N_2408,N_1419);
and U6145 (N_6145,N_2284,N_4535);
nor U6146 (N_6146,N_2899,N_3304);
nand U6147 (N_6147,N_1957,N_3871);
nor U6148 (N_6148,N_2489,N_3209);
and U6149 (N_6149,N_171,N_2067);
or U6150 (N_6150,N_1204,N_3479);
and U6151 (N_6151,N_3489,N_886);
or U6152 (N_6152,N_5901,N_1937);
or U6153 (N_6153,N_434,N_2897);
nand U6154 (N_6154,N_3286,N_5045);
or U6155 (N_6155,N_2339,N_4186);
or U6156 (N_6156,N_1509,N_5987);
xor U6157 (N_6157,N_4671,N_4401);
or U6158 (N_6158,N_4747,N_5234);
nand U6159 (N_6159,N_215,N_5932);
or U6160 (N_6160,N_3968,N_2425);
and U6161 (N_6161,N_1173,N_1541);
and U6162 (N_6162,N_2958,N_386);
nand U6163 (N_6163,N_3921,N_1468);
and U6164 (N_6164,N_3466,N_5401);
xnor U6165 (N_6165,N_787,N_2368);
or U6166 (N_6166,N_922,N_5854);
or U6167 (N_6167,N_2685,N_690);
xnor U6168 (N_6168,N_798,N_69);
or U6169 (N_6169,N_2084,N_646);
nor U6170 (N_6170,N_632,N_1050);
or U6171 (N_6171,N_4042,N_4221);
xnor U6172 (N_6172,N_2299,N_3742);
nor U6173 (N_6173,N_323,N_1983);
xor U6174 (N_6174,N_5294,N_961);
nand U6175 (N_6175,N_745,N_2943);
nand U6176 (N_6176,N_2416,N_167);
and U6177 (N_6177,N_4801,N_2919);
nand U6178 (N_6178,N_1243,N_3910);
nor U6179 (N_6179,N_675,N_1269);
nand U6180 (N_6180,N_619,N_3373);
and U6181 (N_6181,N_1745,N_5766);
or U6182 (N_6182,N_1985,N_4222);
nor U6183 (N_6183,N_4653,N_3893);
nand U6184 (N_6184,N_3032,N_5287);
xnor U6185 (N_6185,N_371,N_2675);
xor U6186 (N_6186,N_5565,N_3768);
and U6187 (N_6187,N_1970,N_4825);
and U6188 (N_6188,N_264,N_5943);
nor U6189 (N_6189,N_1151,N_2727);
nand U6190 (N_6190,N_2263,N_754);
or U6191 (N_6191,N_2216,N_1564);
or U6192 (N_6192,N_1279,N_156);
nor U6193 (N_6193,N_1306,N_391);
xnor U6194 (N_6194,N_4140,N_1952);
nor U6195 (N_6195,N_1248,N_252);
nor U6196 (N_6196,N_5228,N_3140);
xnor U6197 (N_6197,N_4726,N_1239);
nor U6198 (N_6198,N_2106,N_4238);
xor U6199 (N_6199,N_4342,N_5825);
xor U6200 (N_6200,N_4803,N_658);
nor U6201 (N_6201,N_4731,N_2072);
nand U6202 (N_6202,N_656,N_150);
nand U6203 (N_6203,N_3428,N_1922);
nor U6204 (N_6204,N_974,N_3176);
and U6205 (N_6205,N_2640,N_2808);
xnor U6206 (N_6206,N_1887,N_2775);
and U6207 (N_6207,N_843,N_5935);
nor U6208 (N_6208,N_4675,N_2650);
nor U6209 (N_6209,N_5853,N_3155);
or U6210 (N_6210,N_1018,N_931);
nor U6211 (N_6211,N_295,N_4005);
and U6212 (N_6212,N_510,N_5184);
or U6213 (N_6213,N_3104,N_14);
and U6214 (N_6214,N_1191,N_1030);
nand U6215 (N_6215,N_1246,N_1456);
or U6216 (N_6216,N_3866,N_2580);
nor U6217 (N_6217,N_5044,N_424);
and U6218 (N_6218,N_907,N_3611);
nand U6219 (N_6219,N_4551,N_1754);
and U6220 (N_6220,N_92,N_1055);
nand U6221 (N_6221,N_3542,N_5350);
xnor U6222 (N_6222,N_340,N_2735);
nand U6223 (N_6223,N_4428,N_4934);
or U6224 (N_6224,N_3515,N_2964);
nor U6225 (N_6225,N_4685,N_3602);
nand U6226 (N_6226,N_3120,N_5725);
xor U6227 (N_6227,N_202,N_1504);
xor U6228 (N_6228,N_5690,N_3010);
xor U6229 (N_6229,N_972,N_1428);
nand U6230 (N_6230,N_3644,N_3208);
or U6231 (N_6231,N_205,N_436);
or U6232 (N_6232,N_3881,N_2638);
and U6233 (N_6233,N_5275,N_5297);
xor U6234 (N_6234,N_5392,N_4098);
and U6235 (N_6235,N_2080,N_2527);
nand U6236 (N_6236,N_5339,N_3678);
or U6237 (N_6237,N_4509,N_1265);
or U6238 (N_6238,N_2991,N_1876);
or U6239 (N_6239,N_1261,N_5459);
nor U6240 (N_6240,N_161,N_1605);
or U6241 (N_6241,N_2750,N_5273);
nand U6242 (N_6242,N_3673,N_1787);
or U6243 (N_6243,N_375,N_730);
nor U6244 (N_6244,N_1143,N_3814);
nand U6245 (N_6245,N_1875,N_614);
nand U6246 (N_6246,N_277,N_5601);
or U6247 (N_6247,N_2366,N_5227);
and U6248 (N_6248,N_4330,N_2855);
nand U6249 (N_6249,N_1756,N_4312);
xor U6250 (N_6250,N_4184,N_1587);
or U6251 (N_6251,N_5371,N_4835);
and U6252 (N_6252,N_4261,N_5923);
nor U6253 (N_6253,N_877,N_875);
xor U6254 (N_6254,N_4557,N_2854);
or U6255 (N_6255,N_3989,N_3571);
nor U6256 (N_6256,N_1513,N_1585);
and U6257 (N_6257,N_5154,N_4069);
nand U6258 (N_6258,N_1302,N_2962);
nor U6259 (N_6259,N_1827,N_728);
nand U6260 (N_6260,N_2030,N_3302);
or U6261 (N_6261,N_2197,N_671);
and U6262 (N_6262,N_3689,N_884);
nor U6263 (N_6263,N_3582,N_1370);
xor U6264 (N_6264,N_4226,N_3156);
nor U6265 (N_6265,N_3486,N_1312);
or U6266 (N_6266,N_2963,N_3454);
xnor U6267 (N_6267,N_2118,N_3927);
or U6268 (N_6268,N_3698,N_3095);
nor U6269 (N_6269,N_4748,N_5352);
and U6270 (N_6270,N_1618,N_5694);
nor U6271 (N_6271,N_2207,N_1069);
and U6272 (N_6272,N_4046,N_2485);
nor U6273 (N_6273,N_5105,N_4281);
or U6274 (N_6274,N_1501,N_1620);
nor U6275 (N_6275,N_3243,N_2670);
nand U6276 (N_6276,N_1567,N_3822);
or U6277 (N_6277,N_2059,N_2512);
xor U6278 (N_6278,N_1637,N_1940);
nand U6279 (N_6279,N_5402,N_3532);
nor U6280 (N_6280,N_3003,N_4709);
and U6281 (N_6281,N_400,N_4772);
xnor U6282 (N_6282,N_3040,N_1879);
xnor U6283 (N_6283,N_4031,N_492);
or U6284 (N_6284,N_3448,N_1314);
nor U6285 (N_6285,N_5300,N_4303);
xor U6286 (N_6286,N_3455,N_1470);
xor U6287 (N_6287,N_4687,N_2020);
nand U6288 (N_6288,N_266,N_5313);
nand U6289 (N_6289,N_3270,N_3562);
or U6290 (N_6290,N_4396,N_4730);
xor U6291 (N_6291,N_2846,N_3291);
nor U6292 (N_6292,N_1554,N_5801);
xor U6293 (N_6293,N_3081,N_1211);
xor U6294 (N_6294,N_3752,N_4012);
xnor U6295 (N_6295,N_4842,N_789);
or U6296 (N_6296,N_2063,N_4110);
xnor U6297 (N_6297,N_2686,N_284);
nand U6298 (N_6298,N_2394,N_1662);
or U6299 (N_6299,N_5075,N_2167);
or U6300 (N_6300,N_724,N_5215);
or U6301 (N_6301,N_5206,N_2317);
or U6302 (N_6302,N_2893,N_668);
and U6303 (N_6303,N_2481,N_4529);
xnor U6304 (N_6304,N_1562,N_3203);
xor U6305 (N_6305,N_5233,N_1330);
or U6306 (N_6306,N_4061,N_3569);
or U6307 (N_6307,N_3797,N_5116);
or U6308 (N_6308,N_1946,N_2222);
or U6309 (N_6309,N_2507,N_4092);
or U6310 (N_6310,N_5548,N_5426);
nor U6311 (N_6311,N_5243,N_1675);
xor U6312 (N_6312,N_5531,N_2708);
xnor U6313 (N_6313,N_4790,N_3833);
nor U6314 (N_6314,N_1921,N_793);
and U6315 (N_6315,N_3135,N_4230);
or U6316 (N_6316,N_4866,N_22);
nor U6317 (N_6317,N_4111,N_4849);
or U6318 (N_6318,N_1335,N_2279);
nor U6319 (N_6319,N_4695,N_563);
nand U6320 (N_6320,N_5936,N_2792);
or U6321 (N_6321,N_5783,N_4394);
and U6322 (N_6322,N_5048,N_2751);
xor U6323 (N_6323,N_5757,N_623);
nand U6324 (N_6324,N_3146,N_809);
and U6325 (N_6325,N_520,N_2468);
or U6326 (N_6326,N_4562,N_5203);
nand U6327 (N_6327,N_4066,N_5682);
xnor U6328 (N_6328,N_5169,N_1008);
nor U6329 (N_6329,N_2352,N_226);
or U6330 (N_6330,N_2053,N_4197);
and U6331 (N_6331,N_2649,N_258);
and U6332 (N_6332,N_5865,N_3269);
xor U6333 (N_6333,N_1929,N_5014);
and U6334 (N_6334,N_4104,N_3526);
nor U6335 (N_6335,N_270,N_332);
or U6336 (N_6336,N_85,N_2048);
nor U6337 (N_6337,N_5511,N_2155);
xor U6338 (N_6338,N_2078,N_5503);
nor U6339 (N_6339,N_2225,N_1682);
nor U6340 (N_6340,N_3595,N_1188);
and U6341 (N_6341,N_4463,N_4980);
xor U6342 (N_6342,N_4958,N_543);
xnor U6343 (N_6343,N_2699,N_4635);
or U6344 (N_6344,N_2297,N_2567);
xnor U6345 (N_6345,N_3262,N_2229);
nor U6346 (N_6346,N_2978,N_4245);
or U6347 (N_6347,N_2192,N_4411);
nor U6348 (N_6348,N_2283,N_2264);
xor U6349 (N_6349,N_4553,N_5571);
and U6350 (N_6350,N_2139,N_2144);
nand U6351 (N_6351,N_1487,N_2228);
nand U6352 (N_6352,N_1938,N_4160);
xnor U6353 (N_6353,N_350,N_3132);
or U6354 (N_6354,N_2060,N_3151);
nor U6355 (N_6355,N_4371,N_722);
xnor U6356 (N_6356,N_5674,N_4755);
nor U6357 (N_6357,N_4,N_5817);
nor U6358 (N_6358,N_5097,N_2492);
nor U6359 (N_6359,N_2270,N_3255);
nand U6360 (N_6360,N_5367,N_5558);
nor U6361 (N_6361,N_5831,N_3108);
nand U6362 (N_6362,N_3379,N_3388);
nor U6363 (N_6363,N_3757,N_3008);
nand U6364 (N_6364,N_493,N_1206);
and U6365 (N_6365,N_5957,N_727);
nor U6366 (N_6366,N_702,N_5182);
and U6367 (N_6367,N_2097,N_2049);
or U6368 (N_6368,N_2023,N_2872);
or U6369 (N_6369,N_114,N_3567);
or U6370 (N_6370,N_3853,N_13);
nand U6371 (N_6371,N_2116,N_4715);
nor U6372 (N_6372,N_5620,N_1334);
or U6373 (N_6373,N_2095,N_2188);
nand U6374 (N_6374,N_4961,N_18);
xnor U6375 (N_6375,N_3877,N_3387);
xnor U6376 (N_6376,N_3362,N_1147);
nand U6377 (N_6377,N_4149,N_4128);
xor U6378 (N_6378,N_1873,N_2460);
nor U6379 (N_6379,N_1361,N_3230);
nor U6380 (N_6380,N_2134,N_2702);
nand U6381 (N_6381,N_5684,N_2160);
or U6382 (N_6382,N_4912,N_2050);
and U6383 (N_6383,N_5830,N_2956);
nor U6384 (N_6384,N_5179,N_1578);
xnor U6385 (N_6385,N_2609,N_3981);
nor U6386 (N_6386,N_1804,N_4478);
nor U6387 (N_6387,N_3826,N_3358);
nor U6388 (N_6388,N_1867,N_333);
nor U6389 (N_6389,N_1894,N_254);
nor U6390 (N_6390,N_292,N_692);
nand U6391 (N_6391,N_5096,N_2795);
nor U6392 (N_6392,N_3809,N_5509);
or U6393 (N_6393,N_3527,N_5634);
nor U6394 (N_6394,N_5157,N_4419);
nor U6395 (N_6395,N_151,N_1668);
nor U6396 (N_6396,N_5951,N_4286);
xor U6397 (N_6397,N_2223,N_25);
and U6398 (N_6398,N_3986,N_5285);
nand U6399 (N_6399,N_3561,N_743);
xor U6400 (N_6400,N_1175,N_4178);
nand U6401 (N_6401,N_1015,N_5213);
nand U6402 (N_6402,N_657,N_2151);
and U6403 (N_6403,N_4870,N_4720);
or U6404 (N_6404,N_608,N_1064);
or U6405 (N_6405,N_1625,N_2186);
xnor U6406 (N_6406,N_1010,N_2009);
nor U6407 (N_6407,N_2083,N_4358);
xor U6408 (N_6408,N_2498,N_1485);
or U6409 (N_6409,N_5492,N_5756);
nor U6410 (N_6410,N_3213,N_3891);
or U6411 (N_6411,N_3653,N_1994);
nor U6412 (N_6412,N_3898,N_15);
nor U6413 (N_6413,N_1974,N_1953);
nor U6414 (N_6414,N_3310,N_2327);
and U6415 (N_6415,N_4624,N_1719);
xor U6416 (N_6416,N_1534,N_4464);
xnor U6417 (N_6417,N_1838,N_4009);
or U6418 (N_6418,N_4025,N_2469);
xor U6419 (N_6419,N_1423,N_5286);
and U6420 (N_6420,N_3657,N_4156);
nand U6421 (N_6421,N_3508,N_1999);
xnor U6422 (N_6422,N_3122,N_3401);
nand U6423 (N_6423,N_97,N_2726);
nand U6424 (N_6424,N_780,N_2700);
or U6425 (N_6425,N_920,N_3261);
or U6426 (N_6426,N_1222,N_5860);
nand U6427 (N_6427,N_3077,N_3613);
xor U6428 (N_6428,N_5342,N_3519);
or U6429 (N_6429,N_4224,N_5644);
nand U6430 (N_6430,N_4815,N_3831);
and U6431 (N_6431,N_3297,N_1237);
nor U6432 (N_6432,N_5086,N_1349);
nand U6433 (N_6433,N_1840,N_4363);
and U6434 (N_6434,N_609,N_2071);
xnor U6435 (N_6435,N_5451,N_3381);
nand U6436 (N_6436,N_426,N_3632);
nor U6437 (N_6437,N_243,N_5653);
or U6438 (N_6438,N_3574,N_5667);
nor U6439 (N_6439,N_2844,N_3784);
nand U6440 (N_6440,N_1973,N_5758);
xor U6441 (N_6441,N_5813,N_5595);
and U6442 (N_6442,N_4689,N_4620);
xor U6443 (N_6443,N_1448,N_1063);
or U6444 (N_6444,N_678,N_3775);
and U6445 (N_6445,N_4548,N_1860);
and U6446 (N_6446,N_1371,N_1475);
nand U6447 (N_6447,N_3333,N_1162);
xnor U6448 (N_6448,N_1431,N_1676);
nor U6449 (N_6449,N_3864,N_1223);
or U6450 (N_6450,N_3969,N_2903);
and U6451 (N_6451,N_3392,N_3460);
xnor U6452 (N_6452,N_2086,N_929);
nor U6453 (N_6453,N_3395,N_1300);
nand U6454 (N_6454,N_1833,N_3872);
and U6455 (N_6455,N_372,N_4099);
nand U6456 (N_6456,N_2931,N_2680);
or U6457 (N_6457,N_1105,N_3559);
and U6458 (N_6458,N_853,N_341);
nor U6459 (N_6459,N_5021,N_2892);
xnor U6460 (N_6460,N_2574,N_4900);
or U6461 (N_6461,N_4883,N_5738);
nor U6462 (N_6462,N_3162,N_3021);
xnor U6463 (N_6463,N_12,N_1762);
or U6464 (N_6464,N_2169,N_2693);
or U6465 (N_6465,N_3498,N_3937);
nand U6466 (N_6466,N_1085,N_4267);
nor U6467 (N_6467,N_4094,N_4368);
or U6468 (N_6468,N_5618,N_5158);
xor U6469 (N_6469,N_3933,N_3365);
nand U6470 (N_6470,N_2719,N_2399);
nor U6471 (N_6471,N_3427,N_4594);
and U6472 (N_6472,N_5365,N_4543);
and U6473 (N_6473,N_3157,N_2570);
nor U6474 (N_6474,N_184,N_3072);
nor U6475 (N_6475,N_3206,N_411);
nand U6476 (N_6476,N_2005,N_1165);
or U6477 (N_6477,N_1022,N_4862);
nor U6478 (N_6478,N_3551,N_4847);
xor U6479 (N_6479,N_4356,N_1823);
xor U6480 (N_6480,N_2551,N_4169);
xnor U6481 (N_6481,N_3271,N_1872);
and U6482 (N_6482,N_3247,N_3347);
xor U6483 (N_6483,N_5452,N_5785);
xnor U6484 (N_6484,N_4484,N_1932);
xnor U6485 (N_6485,N_140,N_1473);
xnor U6486 (N_6486,N_768,N_3942);
and U6487 (N_6487,N_5551,N_4680);
or U6488 (N_6488,N_1956,N_2576);
xor U6489 (N_6489,N_2471,N_5448);
nand U6490 (N_6490,N_4113,N_4017);
and U6491 (N_6491,N_1515,N_673);
nand U6492 (N_6492,N_3563,N_2170);
and U6493 (N_6493,N_1776,N_4758);
xor U6494 (N_6494,N_536,N_4280);
nor U6495 (N_6495,N_4505,N_2515);
and U6496 (N_6496,N_2154,N_4203);
and U6497 (N_6497,N_306,N_4474);
nand U6498 (N_6498,N_4235,N_3540);
or U6499 (N_6499,N_1364,N_248);
xor U6500 (N_6500,N_1348,N_3659);
nand U6501 (N_6501,N_3134,N_1936);
nand U6502 (N_6502,N_1420,N_735);
xnor U6503 (N_6503,N_5323,N_2984);
xor U6504 (N_6504,N_1980,N_5335);
and U6505 (N_6505,N_5559,N_4622);
nand U6506 (N_6506,N_1111,N_462);
xnor U6507 (N_6507,N_3702,N_4418);
xnor U6508 (N_6508,N_4333,N_1380);
xor U6509 (N_6509,N_5752,N_4940);
xor U6510 (N_6510,N_5878,N_5557);
and U6511 (N_6511,N_2275,N_2790);
or U6512 (N_6512,N_5336,N_630);
and U6513 (N_6513,N_3861,N_4389);
xnor U6514 (N_6514,N_995,N_863);
and U6515 (N_6515,N_4170,N_4865);
xor U6516 (N_6516,N_1021,N_4465);
and U6517 (N_6517,N_666,N_5404);
nand U6518 (N_6518,N_5100,N_1026);
nand U6519 (N_6519,N_2837,N_5053);
or U6520 (N_6520,N_895,N_5669);
nand U6521 (N_6521,N_5319,N_3416);
nor U6522 (N_6522,N_5988,N_4941);
and U6523 (N_6523,N_1446,N_2004);
and U6524 (N_6524,N_4381,N_792);
or U6525 (N_6525,N_5163,N_5687);
xnor U6526 (N_6526,N_2874,N_2138);
xnor U6527 (N_6527,N_4804,N_2226);
or U6528 (N_6528,N_1901,N_4984);
nor U6529 (N_6529,N_4010,N_3609);
and U6530 (N_6530,N_1545,N_1898);
nand U6531 (N_6531,N_2809,N_4600);
nand U6532 (N_6532,N_1703,N_696);
nor U6533 (N_6533,N_3817,N_541);
or U6534 (N_6534,N_5855,N_3688);
and U6535 (N_6535,N_1402,N_2419);
xor U6536 (N_6536,N_942,N_5708);
xor U6537 (N_6537,N_3450,N_1077);
nand U6538 (N_6538,N_3890,N_352);
or U6539 (N_6539,N_4210,N_3004);
nor U6540 (N_6540,N_912,N_4558);
and U6541 (N_6541,N_960,N_2657);
nand U6542 (N_6542,N_3159,N_2662);
and U6543 (N_6543,N_5444,N_2762);
nand U6544 (N_6544,N_4829,N_4519);
and U6545 (N_6545,N_1292,N_4798);
nand U6546 (N_6546,N_4979,N_3399);
nor U6547 (N_6547,N_3528,N_4157);
xnor U6548 (N_6548,N_2233,N_1989);
xor U6549 (N_6549,N_3950,N_5577);
xnor U6550 (N_6550,N_5279,N_473);
xor U6551 (N_6551,N_3828,N_1263);
or U6552 (N_6552,N_3393,N_3723);
nor U6553 (N_6553,N_4182,N_2141);
and U6554 (N_6554,N_5333,N_4615);
or U6555 (N_6555,N_5337,N_5080);
xnor U6556 (N_6556,N_5038,N_5408);
xnor U6557 (N_6557,N_5574,N_3493);
nor U6558 (N_6558,N_1768,N_767);
xor U6559 (N_6559,N_4933,N_836);
or U6560 (N_6560,N_1230,N_4124);
and U6561 (N_6561,N_4511,N_2629);
xnor U6562 (N_6562,N_1839,N_1971);
and U6563 (N_6563,N_5711,N_220);
and U6564 (N_6564,N_1601,N_2453);
nor U6565 (N_6565,N_4151,N_3905);
and U6566 (N_6566,N_1096,N_1099);
nor U6567 (N_6567,N_4691,N_5061);
nand U6568 (N_6568,N_2959,N_3041);
and U6569 (N_6569,N_5081,N_303);
nand U6570 (N_6570,N_3832,N_882);
and U6571 (N_6571,N_4256,N_3068);
and U6572 (N_6572,N_1651,N_4088);
and U6573 (N_6573,N_5852,N_1492);
and U6574 (N_6574,N_4422,N_2426);
or U6575 (N_6575,N_4180,N_3800);
and U6576 (N_6576,N_2810,N_387);
and U6577 (N_6577,N_2029,N_2884);
or U6578 (N_6578,N_268,N_2746);
nor U6579 (N_6579,N_2993,N_3640);
nor U6580 (N_6580,N_888,N_4370);
and U6581 (N_6581,N_4827,N_5152);
nor U6582 (N_6582,N_1114,N_3959);
xor U6583 (N_6583,N_3918,N_2761);
or U6584 (N_6584,N_5905,N_4998);
nand U6585 (N_6585,N_2695,N_1495);
and U6586 (N_6586,N_4792,N_5960);
xnor U6587 (N_6587,N_653,N_2749);
or U6588 (N_6588,N_4921,N_218);
nor U6589 (N_6589,N_401,N_5360);
or U6590 (N_6590,N_2442,N_2143);
or U6591 (N_6591,N_1033,N_4860);
nand U6592 (N_6592,N_4288,N_3254);
xor U6593 (N_6593,N_1663,N_4284);
and U6594 (N_6594,N_5985,N_2488);
and U6595 (N_6595,N_5191,N_2383);
xor U6596 (N_6596,N_4839,N_3544);
or U6597 (N_6597,N_4444,N_2147);
nor U6598 (N_6598,N_4114,N_1128);
nand U6599 (N_6599,N_2616,N_3231);
or U6600 (N_6600,N_5750,N_466);
or U6601 (N_6601,N_5554,N_2281);
and U6602 (N_6602,N_2672,N_2921);
xor U6603 (N_6603,N_271,N_1242);
nor U6604 (N_6604,N_5018,N_3424);
and U6605 (N_6605,N_5390,N_2724);
nand U6606 (N_6606,N_2376,N_3430);
xnor U6607 (N_6607,N_2599,N_1569);
xor U6608 (N_6608,N_3583,N_287);
nand U6609 (N_6609,N_5435,N_5593);
nor U6610 (N_6610,N_112,N_4190);
nand U6611 (N_6611,N_3217,N_5777);
xnor U6612 (N_6612,N_4676,N_592);
nand U6613 (N_6613,N_4499,N_5296);
nand U6614 (N_6614,N_2025,N_3516);
nand U6615 (N_6615,N_4705,N_3180);
and U6616 (N_6616,N_4056,N_2948);
nand U6617 (N_6617,N_5373,N_4103);
nor U6618 (N_6618,N_3049,N_2158);
or U6619 (N_6619,N_5443,N_5991);
and U6620 (N_6620,N_4920,N_4577);
nor U6621 (N_6621,N_5487,N_4619);
or U6622 (N_6622,N_5355,N_1005);
nor U6623 (N_6623,N_3006,N_3188);
nand U6624 (N_6624,N_5120,N_4071);
nand U6625 (N_6625,N_3351,N_738);
xnor U6626 (N_6626,N_5519,N_4372);
xor U6627 (N_6627,N_2538,N_2258);
and U6628 (N_6628,N_2026,N_4324);
and U6629 (N_6629,N_2477,N_163);
xnor U6630 (N_6630,N_2996,N_141);
xnor U6631 (N_6631,N_4030,N_1036);
nand U6632 (N_6632,N_3639,N_2595);
or U6633 (N_6633,N_892,N_5874);
and U6634 (N_6634,N_4105,N_4096);
nand U6635 (N_6635,N_3573,N_1182);
or U6636 (N_6636,N_1907,N_3762);
or U6637 (N_6637,N_839,N_2979);
or U6638 (N_6638,N_1782,N_1480);
nor U6639 (N_6639,N_2927,N_2371);
xnor U6640 (N_6640,N_5931,N_4917);
and U6641 (N_6641,N_1852,N_4032);
nor U6642 (N_6642,N_5915,N_118);
xor U6643 (N_6643,N_5465,N_1385);
and U6644 (N_6644,N_2412,N_4116);
and U6645 (N_6645,N_1123,N_4734);
xnor U6646 (N_6646,N_5695,N_5123);
nand U6647 (N_6647,N_3945,N_3860);
xnor U6648 (N_6648,N_4608,N_1890);
or U6649 (N_6649,N_2864,N_1287);
or U6650 (N_6650,N_2760,N_5762);
or U6651 (N_6651,N_481,N_1016);
nor U6652 (N_6652,N_438,N_4550);
or U6653 (N_6653,N_935,N_4024);
and U6654 (N_6654,N_2888,N_4951);
nand U6655 (N_6655,N_122,N_4699);
xor U6656 (N_6656,N_5822,N_56);
nand U6657 (N_6657,N_1259,N_4846);
nand U6658 (N_6658,N_612,N_1220);
xnor U6659 (N_6659,N_128,N_2980);
nand U6660 (N_6660,N_5436,N_2862);
nor U6661 (N_6661,N_3601,N_4656);
or U6662 (N_6662,N_4014,N_1712);
xnor U6663 (N_6663,N_2335,N_1403);
and U6664 (N_6664,N_103,N_982);
xnor U6665 (N_6665,N_5262,N_2035);
nor U6666 (N_6666,N_5084,N_3221);
or U6667 (N_6667,N_5395,N_1822);
xnor U6668 (N_6668,N_2788,N_5614);
or U6669 (N_6669,N_4701,N_4432);
nand U6670 (N_6670,N_4966,N_539);
and U6671 (N_6671,N_4818,N_1667);
nor U6672 (N_6672,N_2619,N_107);
nor U6673 (N_6673,N_4399,N_1577);
xnor U6674 (N_6674,N_3494,N_3845);
nor U6675 (N_6675,N_774,N_976);
xor U6676 (N_6676,N_177,N_5794);
nand U6677 (N_6677,N_1340,N_27);
nor U6678 (N_6678,N_538,N_2678);
nand U6679 (N_6679,N_679,N_1177);
or U6680 (N_6680,N_5604,N_5305);
and U6681 (N_6681,N_2351,N_4173);
nand U6682 (N_6682,N_2887,N_237);
nand U6683 (N_6683,N_4437,N_4916);
xnor U6684 (N_6684,N_764,N_3652);
xnor U6685 (N_6685,N_763,N_4601);
or U6686 (N_6686,N_3345,N_3523);
or U6687 (N_6687,N_2861,N_715);
nand U6688 (N_6688,N_2304,N_5391);
and U6689 (N_6689,N_3949,N_5237);
or U6690 (N_6690,N_3998,N_582);
xor U6691 (N_6691,N_2689,N_5412);
nor U6692 (N_6692,N_1474,N_1797);
xnor U6693 (N_6693,N_5863,N_5074);
nor U6694 (N_6694,N_821,N_365);
or U6695 (N_6695,N_3324,N_3026);
nand U6696 (N_6696,N_4426,N_1895);
and U6697 (N_6697,N_4159,N_4021);
nor U6698 (N_6698,N_3767,N_902);
nand U6699 (N_6699,N_2950,N_5368);
nor U6700 (N_6700,N_627,N_4717);
or U6701 (N_6701,N_3662,N_5523);
or U6702 (N_6702,N_4800,N_483);
or U6703 (N_6703,N_5755,N_3524);
and U6704 (N_6704,N_2321,N_1628);
xnor U6705 (N_6705,N_1595,N_940);
nor U6706 (N_6706,N_1647,N_4327);
or U6707 (N_6707,N_3093,N_2627);
nor U6708 (N_6708,N_1140,N_4640);
nand U6709 (N_6709,N_3190,N_2784);
nand U6710 (N_6710,N_2153,N_5517);
and U6711 (N_6711,N_978,N_3722);
nand U6712 (N_6712,N_2336,N_1394);
xor U6713 (N_6713,N_1790,N_2543);
nor U6714 (N_6714,N_132,N_2786);
nor U6715 (N_6715,N_2441,N_1029);
and U6716 (N_6716,N_1104,N_4192);
or U6717 (N_6717,N_5575,N_878);
nand U6718 (N_6718,N_903,N_2036);
or U6719 (N_6719,N_5066,N_1961);
nand U6720 (N_6720,N_3730,N_1616);
nor U6721 (N_6721,N_1749,N_4321);
nand U6722 (N_6722,N_3403,N_3411);
or U6723 (N_6723,N_2123,N_3755);
and U6724 (N_6724,N_1295,N_2343);
nand U6725 (N_6725,N_3483,N_445);
and U6726 (N_6726,N_1159,N_1430);
nand U6727 (N_6727,N_967,N_4604);
nor U6728 (N_6728,N_2230,N_1299);
xnor U6729 (N_6729,N_5666,N_3887);
and U6730 (N_6730,N_5696,N_2390);
and U6731 (N_6731,N_642,N_4313);
or U6732 (N_6732,N_3630,N_5133);
or U6733 (N_6733,N_1392,N_4064);
nand U6734 (N_6734,N_2377,N_1650);
or U6735 (N_6735,N_2413,N_879);
nor U6736 (N_6736,N_4826,N_969);
nand U6737 (N_6737,N_5007,N_2210);
xor U6738 (N_6738,N_2125,N_1806);
or U6739 (N_6739,N_4580,N_3223);
nand U6740 (N_6740,N_4045,N_4946);
nor U6741 (N_6741,N_5972,N_4296);
or U6742 (N_6742,N_2038,N_1900);
nor U6743 (N_6743,N_815,N_5457);
or U6744 (N_6744,N_3149,N_1683);
xnor U6745 (N_6745,N_5043,N_2017);
or U6746 (N_6746,N_2933,N_1028);
nand U6747 (N_6747,N_4927,N_4201);
nor U6748 (N_6748,N_1103,N_4345);
and U6749 (N_6749,N_2504,N_335);
nand U6750 (N_6750,N_2720,N_1666);
and U6751 (N_6751,N_1194,N_1500);
and U6752 (N_6752,N_4174,N_4714);
nor U6753 (N_6753,N_448,N_2466);
and U6754 (N_6754,N_1245,N_5211);
and U6755 (N_6755,N_1674,N_389);
xnor U6756 (N_6756,N_502,N_1633);
nand U6757 (N_6757,N_1451,N_3716);
or U6758 (N_6758,N_4949,N_484);
xnor U6759 (N_6759,N_4722,N_4466);
xor U6760 (N_6760,N_3714,N_4131);
nor U6761 (N_6761,N_933,N_2818);
nand U6762 (N_6762,N_3169,N_4850);
xor U6763 (N_6763,N_1415,N_1437);
nor U6764 (N_6764,N_5840,N_72);
nor U6765 (N_6765,N_2372,N_3869);
nor U6766 (N_6766,N_4320,N_4922);
xor U6767 (N_6767,N_5502,N_4364);
or U6768 (N_6768,N_4412,N_4008);
nand U6769 (N_6769,N_1284,N_3770);
xor U6770 (N_6770,N_2273,N_1506);
or U6771 (N_6771,N_475,N_2873);
xor U6772 (N_6772,N_3305,N_1047);
xnor U6773 (N_6773,N_2467,N_585);
or U6774 (N_6774,N_3538,N_5851);
and U6775 (N_6775,N_1917,N_1439);
nand U6776 (N_6776,N_1831,N_3211);
or U6777 (N_6777,N_3110,N_4322);
nor U6778 (N_6778,N_3975,N_1353);
or U6779 (N_6779,N_5774,N_1384);
nor U6780 (N_6780,N_1449,N_3667);
nor U6781 (N_6781,N_5354,N_3139);
or U6782 (N_6782,N_1160,N_2573);
or U6783 (N_6783,N_5041,N_2651);
and U6784 (N_6784,N_1298,N_4643);
or U6785 (N_6785,N_3600,N_2665);
nor U6786 (N_6786,N_4799,N_4053);
xnor U6787 (N_6787,N_373,N_3699);
xnor U6788 (N_6788,N_238,N_2310);
xor U6789 (N_6789,N_3674,N_4168);
and U6790 (N_6790,N_3693,N_5630);
or U6791 (N_6791,N_3462,N_5848);
or U6792 (N_6792,N_584,N_4282);
nor U6793 (N_6793,N_4023,N_3774);
nor U6794 (N_6794,N_212,N_1608);
xnor U6795 (N_6795,N_3402,N_5137);
or U6796 (N_6796,N_1412,N_1286);
and U6797 (N_6797,N_2462,N_4497);
nor U6798 (N_6798,N_82,N_5625);
nor U6799 (N_6799,N_5188,N_3793);
xnor U6800 (N_6800,N_3064,N_5222);
nor U6801 (N_6801,N_91,N_1548);
and U6802 (N_6802,N_4654,N_2043);
and U6803 (N_6803,N_1816,N_4337);
or U6804 (N_6804,N_3592,N_2799);
xnor U6805 (N_6805,N_1945,N_4219);
nand U6806 (N_6806,N_3888,N_1213);
nand U6807 (N_6807,N_4036,N_346);
nor U6808 (N_6808,N_2598,N_5578);
nor U6809 (N_6809,N_5149,N_917);
nand U6810 (N_6810,N_5330,N_4369);
nor U6811 (N_6811,N_1087,N_4814);
xor U6812 (N_6812,N_1869,N_760);
xnor U6813 (N_6813,N_5673,N_4386);
nand U6814 (N_6814,N_924,N_3280);
nor U6815 (N_6815,N_1978,N_265);
nand U6816 (N_6816,N_5090,N_4277);
or U6817 (N_6817,N_4038,N_1466);
and U6818 (N_6818,N_3930,N_222);
and U6819 (N_6819,N_1592,N_2777);
nor U6820 (N_6820,N_1092,N_3121);
xor U6821 (N_6821,N_5082,N_394);
nand U6822 (N_6822,N_2296,N_5635);
nor U6823 (N_6823,N_1109,N_3744);
or U6824 (N_6824,N_2714,N_3240);
or U6825 (N_6825,N_88,N_552);
xnor U6826 (N_6826,N_230,N_5387);
nand U6827 (N_6827,N_3249,N_3625);
or U6828 (N_6828,N_3505,N_5343);
nand U6829 (N_6829,N_2961,N_4319);
and U6830 (N_6830,N_3326,N_3951);
nand U6831 (N_6831,N_2358,N_5909);
or U6832 (N_6832,N_5425,N_1471);
and U6833 (N_6833,N_4493,N_5937);
nor U6834 (N_6834,N_2251,N_2753);
or U6835 (N_6835,N_4896,N_1387);
xor U6836 (N_6836,N_2248,N_5017);
nor U6837 (N_6837,N_1305,N_3327);
or U6838 (N_6838,N_3431,N_5439);
nand U6839 (N_6839,N_5533,N_1863);
or U6840 (N_6840,N_4515,N_2531);
and U6841 (N_6841,N_3323,N_377);
nor U6842 (N_6842,N_4295,N_4770);
and U6843 (N_6843,N_4914,N_5582);
xnor U6844 (N_6844,N_5741,N_4571);
or U6845 (N_6845,N_307,N_1832);
and U6846 (N_6846,N_1309,N_1656);
and U6847 (N_6847,N_1716,N_4945);
nand U6848 (N_6848,N_2387,N_4293);
nand U6849 (N_6849,N_4593,N_4063);
and U6850 (N_6850,N_316,N_5585);
and U6851 (N_6851,N_273,N_4585);
and U6852 (N_6852,N_2745,N_3154);
nand U6853 (N_6853,N_4181,N_3470);
or U6854 (N_6854,N_4665,N_276);
nand U6855 (N_6855,N_3173,N_4040);
nor U6856 (N_6856,N_938,N_5315);
or U6857 (N_6857,N_3459,N_2316);
xnor U6858 (N_6858,N_1774,N_5729);
or U6859 (N_6859,N_3163,N_2723);
or U6860 (N_6860,N_4085,N_1701);
xor U6861 (N_6861,N_3398,N_1037);
xor U6862 (N_6862,N_1915,N_4876);
and U6863 (N_6863,N_5515,N_649);
or U6864 (N_6864,N_2569,N_23);
xnor U6865 (N_6865,N_1934,N_718);
nand U6866 (N_6866,N_4531,N_4048);
nand U6867 (N_6867,N_3913,N_2731);
xor U6868 (N_6868,N_5001,N_1942);
xor U6869 (N_6869,N_2645,N_4774);
and U6870 (N_6870,N_3065,N_3199);
or U6871 (N_6871,N_1424,N_2089);
nor U6872 (N_6872,N_1781,N_4884);
or U6873 (N_6873,N_2869,N_765);
or U6874 (N_6874,N_5584,N_3502);
nor U6875 (N_6875,N_1750,N_3840);
nand U6876 (N_6876,N_516,N_5570);
and U6877 (N_6877,N_5224,N_1583);
and U6878 (N_6878,N_4575,N_4275);
xnor U6879 (N_6879,N_5064,N_5178);
or U6880 (N_6880,N_4161,N_1568);
and U6881 (N_6881,N_980,N_5269);
nor U6882 (N_6882,N_5616,N_5136);
nor U6883 (N_6883,N_1584,N_4485);
xor U6884 (N_6884,N_2212,N_4067);
xor U6885 (N_6885,N_717,N_3115);
and U6886 (N_6886,N_3239,N_5265);
or U6887 (N_6887,N_665,N_4274);
xor U6888 (N_6888,N_219,N_4962);
and U6889 (N_6889,N_2600,N_5396);
nand U6890 (N_6890,N_5259,N_5088);
or U6891 (N_6891,N_5913,N_5140);
nand U6892 (N_6892,N_5784,N_3100);
xor U6893 (N_6893,N_66,N_849);
nor U6894 (N_6894,N_1916,N_5545);
and U6895 (N_6895,N_589,N_3390);
nor U6896 (N_6896,N_2910,N_3289);
xor U6897 (N_6897,N_379,N_178);
and U6898 (N_6898,N_2006,N_3908);
and U6899 (N_6899,N_392,N_2449);
xnor U6900 (N_6900,N_4403,N_1697);
and U6901 (N_6901,N_3033,N_5349);
and U6902 (N_6902,N_564,N_3664);
or U6903 (N_6903,N_2938,N_4125);
and U6904 (N_6904,N_2916,N_1976);
or U6905 (N_6905,N_1120,N_533);
nand U6906 (N_6906,N_637,N_487);
or U6907 (N_6907,N_1253,N_4447);
or U6908 (N_6908,N_5514,N_5288);
nand U6909 (N_6909,N_1374,N_3279);
xnor U6910 (N_6910,N_5006,N_953);
nand U6911 (N_6911,N_1073,N_3186);
nand U6912 (N_6912,N_2402,N_881);
and U6913 (N_6913,N_1828,N_2000);
xor U6914 (N_6914,N_5952,N_1195);
nand U6915 (N_6915,N_1229,N_4874);
nor U6916 (N_6916,N_2360,N_3303);
nor U6917 (N_6917,N_4854,N_3482);
nand U6918 (N_6918,N_5870,N_2847);
nor U6919 (N_6919,N_272,N_1171);
nand U6920 (N_6920,N_324,N_5345);
nor U6921 (N_6921,N_101,N_2875);
nor U6922 (N_6922,N_244,N_2114);
nor U6923 (N_6923,N_5087,N_751);
and U6924 (N_6924,N_2267,N_1122);
or U6925 (N_6925,N_3971,N_5624);
and U6926 (N_6926,N_3445,N_837);
nand U6927 (N_6927,N_611,N_1700);
xnor U6928 (N_6928,N_4861,N_755);
nand U6929 (N_6929,N_5594,N_4795);
nor U6930 (N_6930,N_1761,N_4929);
nor U6931 (N_6931,N_603,N_1158);
or U6932 (N_6932,N_3556,N_5146);
xor U6933 (N_6933,N_5398,N_5648);
xor U6934 (N_6934,N_5257,N_771);
and U6935 (N_6935,N_3123,N_3996);
xor U6936 (N_6936,N_4054,N_1924);
or U6937 (N_6937,N_109,N_4377);
nor U6938 (N_6938,N_5793,N_3511);
nand U6939 (N_6939,N_315,N_1979);
or U6940 (N_6940,N_2112,N_2539);
nor U6941 (N_6941,N_4621,N_3669);
nor U6942 (N_6942,N_4903,N_5819);
nor U6943 (N_6943,N_383,N_1256);
and U6944 (N_6944,N_2577,N_3803);
and U6945 (N_6945,N_2870,N_2093);
xor U6946 (N_6946,N_1905,N_5338);
and U6947 (N_6947,N_855,N_4049);
xor U6948 (N_6948,N_1236,N_1483);
xor U6949 (N_6949,N_214,N_169);
xnor U6950 (N_6950,N_2022,N_2181);
nor U6951 (N_6951,N_4317,N_2989);
nand U6952 (N_6952,N_110,N_3313);
and U6953 (N_6953,N_4693,N_138);
xor U6954 (N_6954,N_374,N_3499);
nor U6955 (N_6955,N_2163,N_81);
nand U6956 (N_6956,N_229,N_566);
xnor U6957 (N_6957,N_3435,N_2990);
xnor U6958 (N_6958,N_3958,N_5964);
xnor U6959 (N_6959,N_1622,N_2821);
xnor U6960 (N_6960,N_1386,N_5326);
nand U6961 (N_6961,N_3576,N_4055);
xnor U6962 (N_6962,N_119,N_3970);
or U6963 (N_6963,N_2074,N_968);
nor U6964 (N_6964,N_4398,N_5919);
and U6965 (N_6965,N_4909,N_1404);
and U6966 (N_6966,N_1785,N_4905);
and U6967 (N_6967,N_2494,N_19);
nor U6968 (N_6968,N_476,N_4833);
or U6969 (N_6969,N_2540,N_4988);
nand U6970 (N_6970,N_5812,N_4202);
and U6971 (N_6971,N_442,N_3046);
and U6972 (N_6972,N_1488,N_1753);
xnor U6973 (N_6973,N_687,N_2464);
nand U6974 (N_6974,N_3627,N_5929);
nand U6975 (N_6975,N_3558,N_2866);
or U6976 (N_6976,N_1572,N_5382);
and U6977 (N_6977,N_3276,N_1892);
nand U6978 (N_6978,N_2314,N_1432);
and U6979 (N_6979,N_4147,N_2817);
nand U6980 (N_6980,N_748,N_955);
nor U6981 (N_6981,N_595,N_729);
nor U6982 (N_6982,N_3637,N_1714);
xnor U6983 (N_6983,N_3252,N_4538);
nand U6984 (N_6984,N_3566,N_5566);
xnor U6985 (N_6985,N_5636,N_3618);
xor U6986 (N_6986,N_2863,N_5900);
and U6987 (N_6987,N_1954,N_4737);
nor U6988 (N_6988,N_4360,N_928);
nand U6989 (N_6989,N_1732,N_5779);
or U6990 (N_6990,N_485,N_2002);
nor U6991 (N_6991,N_5534,N_5835);
or U6992 (N_6992,N_1718,N_5849);
or U6993 (N_6993,N_129,N_1570);
or U6994 (N_6994,N_2631,N_183);
nor U6995 (N_6995,N_2977,N_5581);
or U6996 (N_6996,N_1695,N_3638);
or U6997 (N_6997,N_148,N_5885);
xnor U6998 (N_6998,N_1738,N_1769);
and U6999 (N_6999,N_5726,N_1835);
nand U7000 (N_7000,N_1076,N_5740);
or U7001 (N_7001,N_4549,N_3197);
xor U7002 (N_7002,N_846,N_2266);
xor U7003 (N_7003,N_2493,N_2013);
and U7004 (N_7004,N_1691,N_3839);
or U7005 (N_7005,N_1356,N_5410);
xor U7006 (N_7006,N_5641,N_723);
nand U7007 (N_7007,N_5328,N_4880);
xor U7008 (N_7008,N_4475,N_2935);
and U7009 (N_7009,N_399,N_2214);
nor U7010 (N_7010,N_3038,N_3220);
nand U7011 (N_7011,N_547,N_3848);
nand U7012 (N_7012,N_2911,N_3275);
xnor U7013 (N_7013,N_4207,N_1636);
nand U7014 (N_7014,N_5976,N_1115);
nor U7015 (N_7015,N_4651,N_227);
nor U7016 (N_7016,N_41,N_2825);
nand U7017 (N_7017,N_3903,N_5904);
nor U7018 (N_7018,N_3229,N_370);
nand U7019 (N_7019,N_4890,N_2191);
and U7020 (N_7020,N_5236,N_4193);
or U7021 (N_7021,N_180,N_1006);
nor U7022 (N_7022,N_2966,N_647);
or U7023 (N_7023,N_298,N_2280);
nor U7024 (N_7024,N_807,N_2204);
nand U7025 (N_7025,N_2265,N_4126);
and U7026 (N_7026,N_3902,N_5576);
or U7027 (N_7027,N_3091,N_4074);
nor U7028 (N_7028,N_327,N_1313);
and U7029 (N_7029,N_4539,N_3956);
nor U7030 (N_7030,N_4259,N_5504);
and U7031 (N_7031,N_5389,N_2410);
or U7032 (N_7032,N_5884,N_786);
nor U7033 (N_7033,N_2867,N_4978);
or U7034 (N_7034,N_2446,N_3034);
nand U7035 (N_7035,N_3195,N_4824);
or U7036 (N_7036,N_512,N_443);
nor U7037 (N_7037,N_1303,N_4294);
nand U7038 (N_7038,N_4143,N_3846);
and U7039 (N_7039,N_3580,N_4583);
nor U7040 (N_7040,N_985,N_2756);
nor U7041 (N_7041,N_4595,N_3189);
nand U7042 (N_7042,N_4666,N_5645);
xnor U7043 (N_7043,N_5295,N_318);
nand U7044 (N_7044,N_94,N_1034);
xnor U7045 (N_7045,N_1228,N_1351);
nand U7046 (N_7046,N_1375,N_4521);
nor U7047 (N_7047,N_2560,N_3740);
nor U7048 (N_7048,N_1877,N_5427);
nor U7049 (N_7049,N_5749,N_1072);
or U7050 (N_7050,N_5748,N_4932);
nor U7051 (N_7051,N_209,N_4993);
nor U7052 (N_7052,N_4688,N_5709);
and U7053 (N_7053,N_3533,N_1596);
nor U7054 (N_7054,N_2771,N_3400);
or U7055 (N_7055,N_5714,N_53);
or U7056 (N_7056,N_4289,N_2587);
xor U7057 (N_7057,N_3315,N_975);
or U7058 (N_7058,N_4997,N_2732);
nor U7059 (N_7059,N_4926,N_1558);
xnor U7060 (N_7060,N_4765,N_1987);
nor U7061 (N_7061,N_5800,N_5580);
or U7062 (N_7062,N_3579,N_2917);
nand U7063 (N_7063,N_3745,N_3421);
and U7064 (N_7064,N_3138,N_5637);
nand U7065 (N_7065,N_480,N_3474);
nand U7066 (N_7066,N_4694,N_4001);
nand U7067 (N_7067,N_1154,N_1208);
nor U7068 (N_7068,N_3312,N_2789);
and U7069 (N_7069,N_5746,N_2692);
xnor U7070 (N_7070,N_5,N_2472);
nor U7071 (N_7071,N_3359,N_1996);
or U7072 (N_7072,N_3232,N_3278);
and U7073 (N_7073,N_2432,N_3185);
nor U7074 (N_7074,N_3635,N_716);
nand U7075 (N_7075,N_3193,N_5118);
or U7076 (N_7076,N_2518,N_4649);
or U7077 (N_7077,N_2016,N_4247);
nor U7078 (N_7078,N_4020,N_4400);
or U7079 (N_7079,N_5589,N_1332);
and U7080 (N_7080,N_2261,N_2632);
nand U7081 (N_7081,N_1227,N_5650);
and U7082 (N_7082,N_217,N_3993);
or U7083 (N_7083,N_2033,N_4254);
nand U7084 (N_7084,N_3736,N_4065);
nand U7085 (N_7085,N_5803,N_5065);
nor U7086 (N_7086,N_5837,N_2409);
nand U7087 (N_7087,N_1221,N_4563);
nor U7088 (N_7088,N_5921,N_2798);
xor U7089 (N_7089,N_1062,N_2758);
nand U7090 (N_7090,N_3329,N_5446);
nand U7091 (N_7091,N_2535,N_3422);
or U7092 (N_7092,N_2148,N_201);
nand U7093 (N_7093,N_3143,N_4338);
nand U7094 (N_7094,N_747,N_3308);
or U7095 (N_7095,N_3607,N_1820);
or U7096 (N_7096,N_4100,N_2508);
xnor U7097 (N_7097,N_1642,N_5596);
xnor U7098 (N_7098,N_1884,N_5486);
or U7099 (N_7099,N_641,N_3676);
xnor U7100 (N_7100,N_99,N_3724);
xor U7101 (N_7101,N_5672,N_1170);
xnor U7102 (N_7102,N_2012,N_2198);
nor U7103 (N_7103,N_1187,N_5383);
and U7104 (N_7104,N_2547,N_3628);
nor U7105 (N_7105,N_3374,N_3753);
or U7106 (N_7106,N_3548,N_4664);
xor U7107 (N_7107,N_3804,N_5161);
or U7108 (N_7108,N_176,N_601);
and U7109 (N_7109,N_2465,N_4212);
nand U7110 (N_7110,N_4310,N_1741);
and U7111 (N_7111,N_2939,N_364);
nor U7112 (N_7112,N_2286,N_593);
nor U7113 (N_7113,N_2625,N_4834);
nand U7114 (N_7114,N_98,N_1846);
xor U7115 (N_7115,N_2374,N_779);
and U7116 (N_7116,N_4976,N_5406);
nor U7117 (N_7117,N_5483,N_1012);
or U7118 (N_7118,N_1549,N_639);
nor U7119 (N_7119,N_3811,N_3080);
xnor U7120 (N_7120,N_2655,N_2590);
nand U7121 (N_7121,N_3330,N_5882);
xnor U7122 (N_7122,N_5807,N_1189);
and U7123 (N_7123,N_240,N_2276);
or U7124 (N_7124,N_2031,N_1881);
xor U7125 (N_7125,N_32,N_2364);
nor U7126 (N_7126,N_1593,N_1805);
nor U7127 (N_7127,N_3575,N_2302);
xor U7128 (N_7128,N_752,N_819);
nand U7129 (N_7129,N_3105,N_1947);
and U7130 (N_7130,N_2428,N_1153);
or U7131 (N_7131,N_1733,N_5485);
and U7132 (N_7132,N_2988,N_549);
nor U7133 (N_7133,N_1218,N_4242);
xnor U7134 (N_7134,N_1352,N_2525);
xor U7135 (N_7135,N_5628,N_1378);
nand U7136 (N_7136,N_2256,N_1793);
and U7137 (N_7137,N_4152,N_616);
and U7138 (N_7138,N_4410,N_5283);
or U7139 (N_7139,N_3732,N_2868);
nor U7140 (N_7140,N_5417,N_5556);
nor U7141 (N_7141,N_1454,N_3886);
xor U7142 (N_7142,N_714,N_4969);
xor U7143 (N_7143,N_200,N_838);
nand U7144 (N_7144,N_3737,N_1704);
nor U7145 (N_7145,N_5083,N_353);
and U7146 (N_7146,N_482,N_1547);
nand U7147 (N_7147,N_3160,N_2734);
or U7148 (N_7148,N_5151,N_1457);
or U7149 (N_7149,N_4376,N_3238);
nor U7150 (N_7150,N_4109,N_3);
nor U7151 (N_7151,N_5608,N_899);
and U7152 (N_7152,N_2885,N_5129);
or U7153 (N_7153,N_3626,N_5810);
or U7154 (N_7154,N_3061,N_800);
and U7155 (N_7155,N_2208,N_3955);
or U7156 (N_7156,N_2422,N_2291);
nor U7157 (N_7157,N_4506,N_1735);
xnor U7158 (N_7158,N_5029,N_1156);
or U7159 (N_7159,N_3044,N_4565);
nor U7160 (N_7160,N_3663,N_449);
and U7161 (N_7161,N_5495,N_4657);
xor U7162 (N_7162,N_2688,N_488);
nor U7163 (N_7163,N_2300,N_4425);
xnor U7164 (N_7164,N_2986,N_5539);
nor U7165 (N_7165,N_3405,N_2385);
nand U7166 (N_7166,N_2245,N_1054);
nand U7167 (N_7167,N_5181,N_3578);
and U7168 (N_7168,N_3426,N_5030);
nand U7169 (N_7169,N_5805,N_2826);
nor U7170 (N_7170,N_5489,N_2787);
nor U7171 (N_7171,N_2132,N_4241);
nand U7172 (N_7172,N_5530,N_2663);
and U7173 (N_7173,N_803,N_820);
nand U7174 (N_7174,N_90,N_4325);
and U7175 (N_7175,N_2386,N_3439);
and U7176 (N_7176,N_4872,N_3099);
and U7177 (N_7177,N_2111,N_685);
xnor U7178 (N_7178,N_422,N_3076);
nand U7179 (N_7179,N_5047,N_1337);
and U7180 (N_7180,N_720,N_3019);
nor U7181 (N_7181,N_1858,N_3456);
and U7182 (N_7182,N_4472,N_2736);
xor U7183 (N_7183,N_1435,N_5961);
and U7184 (N_7184,N_2312,N_2463);
nor U7185 (N_7185,N_906,N_425);
xnor U7186 (N_7186,N_4552,N_5190);
nand U7187 (N_7187,N_4209,N_3549);
xnor U7188 (N_7188,N_5411,N_801);
or U7189 (N_7189,N_1777,N_5790);
and U7190 (N_7190,N_20,N_2744);
nand U7191 (N_7191,N_2090,N_5036);
xor U7192 (N_7192,N_1100,N_2340);
or U7193 (N_7193,N_5003,N_2857);
or U7194 (N_7194,N_3184,N_28);
nor U7195 (N_7195,N_5059,N_5828);
nand U7196 (N_7196,N_5691,N_1725);
and U7197 (N_7197,N_3074,N_2985);
or U7198 (N_7198,N_3172,N_2764);
xnor U7199 (N_7199,N_4265,N_4564);
nor U7200 (N_7200,N_199,N_3920);
nor U7201 (N_7201,N_2113,N_5037);
and U7202 (N_7202,N_5070,N_3370);
or U7203 (N_7203,N_5309,N_3414);
xor U7204 (N_7204,N_2562,N_5772);
or U7205 (N_7205,N_1639,N_966);
nor U7206 (N_7206,N_1359,N_1874);
nand U7207 (N_7207,N_2513,N_3434);
or U7208 (N_7208,N_5418,N_1411);
nand U7209 (N_7209,N_1450,N_4379);
xor U7210 (N_7210,N_1893,N_5145);
or U7211 (N_7211,N_1376,N_4467);
and U7212 (N_7212,N_2687,N_3118);
nor U7213 (N_7213,N_5507,N_3687);
nor U7214 (N_7214,N_3629,N_2417);
or U7215 (N_7215,N_4544,N_3130);
or U7216 (N_7216,N_5107,N_4336);
and U7217 (N_7217,N_5277,N_2774);
nand U7218 (N_7218,N_3622,N_1861);
and U7219 (N_7219,N_2556,N_709);
xor U7220 (N_7220,N_4429,N_5676);
xor U7221 (N_7221,N_2967,N_2614);
nand U7222 (N_7222,N_4354,N_4913);
nor U7223 (N_7223,N_908,N_5240);
or U7224 (N_7224,N_2568,N_3152);
xnor U7225 (N_7225,N_2202,N_4458);
and U7226 (N_7226,N_1654,N_5815);
nor U7227 (N_7227,N_1619,N_45);
nor U7228 (N_7228,N_3472,N_501);
and U7229 (N_7229,N_3510,N_288);
nand U7230 (N_7230,N_185,N_1752);
nand U7231 (N_7231,N_703,N_5428);
xor U7232 (N_7232,N_5763,N_3726);
nor U7233 (N_7233,N_1516,N_3895);
nor U7234 (N_7234,N_5464,N_100);
and U7235 (N_7235,N_5056,N_699);
and U7236 (N_7236,N_5883,N_1904);
xor U7237 (N_7237,N_5117,N_2982);
nand U7238 (N_7238,N_2328,N_5496);
nor U7239 (N_7239,N_1614,N_5572);
nand U7240 (N_7240,N_3306,N_3789);
or U7241 (N_7241,N_1443,N_697);
nand U7242 (N_7242,N_3237,N_5458);
nand U7243 (N_7243,N_1736,N_3042);
or U7244 (N_7244,N_4263,N_1550);
nand U7245 (N_7245,N_2319,N_5743);
xnor U7246 (N_7246,N_3086,N_2260);
nand U7247 (N_7247,N_60,N_5329);
or U7248 (N_7248,N_3363,N_1685);
nand U7249 (N_7249,N_4501,N_1250);
or U7250 (N_7250,N_934,N_4567);
and U7251 (N_7251,N_2182,N_758);
xor U7252 (N_7252,N_575,N_3236);
or U7253 (N_7253,N_2247,N_4936);
nand U7254 (N_7254,N_3734,N_1275);
nor U7255 (N_7255,N_4627,N_625);
nor U7256 (N_7256,N_1941,N_1267);
and U7257 (N_7257,N_4427,N_2881);
xor U7258 (N_7258,N_1706,N_356);
or U7259 (N_7259,N_3341,N_5833);
or U7260 (N_7260,N_396,N_5023);
and U7261 (N_7261,N_1731,N_70);
nand U7262 (N_7262,N_1043,N_3916);
xnor U7263 (N_7263,N_4768,N_4503);
nor U7264 (N_7264,N_5015,N_1702);
or U7265 (N_7265,N_275,N_1818);
nand U7266 (N_7266,N_5013,N_1686);
and U7267 (N_7267,N_5180,N_5981);
nor U7268 (N_7268,N_1812,N_5612);
or U7269 (N_7269,N_1551,N_598);
and U7270 (N_7270,N_804,N_3377);
nor U7271 (N_7271,N_310,N_2338);
xor U7272 (N_7272,N_2165,N_5944);
or U7273 (N_7273,N_4119,N_2524);
or U7274 (N_7274,N_1142,N_1882);
nor U7275 (N_7275,N_1135,N_826);
or U7276 (N_7276,N_2382,N_4591);
or U7277 (N_7277,N_4033,N_2564);
nor U7278 (N_7278,N_3856,N_1968);
xnor U7279 (N_7279,N_367,N_388);
xor U7280 (N_7280,N_867,N_1291);
and U7281 (N_7281,N_223,N_2831);
nand U7282 (N_7282,N_2952,N_1254);
or U7283 (N_7283,N_1984,N_1814);
nand U7284 (N_7284,N_1401,N_2285);
xnor U7285 (N_7285,N_916,N_1933);
or U7286 (N_7286,N_3656,N_4335);
nand U7287 (N_7287,N_5114,N_4942);
and U7288 (N_7288,N_2618,N_4083);
and U7289 (N_7289,N_4968,N_2405);
or U7290 (N_7290,N_3694,N_4214);
and U7291 (N_7291,N_4439,N_4253);
xnor U7292 (N_7292,N_5540,N_3098);
nor U7293 (N_7293,N_5327,N_5235);
and U7294 (N_7294,N_4525,N_4130);
xnor U7295 (N_7295,N_1013,N_3938);
nor U7296 (N_7296,N_1011,N_2838);
xnor U7297 (N_7297,N_2126,N_3001);
and U7298 (N_7298,N_812,N_4332);
nand U7299 (N_7299,N_2440,N_4495);
xnor U7300 (N_7300,N_3586,N_2592);
nor U7301 (N_7301,N_5463,N_1252);
nor U7302 (N_7302,N_4823,N_5992);
nand U7303 (N_7303,N_2803,N_2594);
or U7304 (N_7304,N_4016,N_5416);
or U7305 (N_7305,N_4176,N_2953);
and U7306 (N_7306,N_5888,N_858);
nor U7307 (N_7307,N_4188,N_4027);
or U7308 (N_7308,N_2028,N_1635);
or U7309 (N_7309,N_4659,N_5429);
and U7310 (N_7310,N_823,N_2484);
or U7311 (N_7311,N_2209,N_2454);
or U7312 (N_7312,N_2858,N_5553);
xnor U7313 (N_7313,N_3919,N_4959);
nor U7314 (N_7314,N_4187,N_1878);
or U7315 (N_7315,N_1383,N_5176);
or U7316 (N_7316,N_918,N_1381);
nand U7317 (N_7317,N_4729,N_2487);
or U7318 (N_7318,N_3787,N_4070);
and U7319 (N_7319,N_5528,N_5664);
xnor U7320 (N_7320,N_4767,N_1166);
and U7321 (N_7321,N_2896,N_1677);
nand U7322 (N_7322,N_5063,N_1118);
nor U7323 (N_7323,N_3316,N_1053);
and U7324 (N_7324,N_4719,N_4301);
nand U7325 (N_7325,N_1093,N_299);
and U7326 (N_7326,N_503,N_4154);
xnor U7327 (N_7327,N_4956,N_550);
nor U7328 (N_7328,N_4856,N_5911);
and U7329 (N_7329,N_3500,N_3219);
xnor U7330 (N_7330,N_2062,N_2173);
nor U7331 (N_7331,N_517,N_508);
nor U7332 (N_7332,N_2365,N_5049);
xor U7333 (N_7333,N_3127,N_3083);
and U7334 (N_7334,N_433,N_3911);
and U7335 (N_7335,N_1630,N_3311);
nand U7336 (N_7336,N_5497,N_3825);
nor U7337 (N_7337,N_203,N_535);
or U7338 (N_7338,N_3593,N_3087);
nor U7339 (N_7339,N_5930,N_5488);
nor U7340 (N_7340,N_1511,N_5346);
nand U7341 (N_7341,N_5902,N_1594);
nor U7342 (N_7342,N_2928,N_4481);
nand U7343 (N_7343,N_5654,N_2972);
nand U7344 (N_7344,N_1421,N_655);
nor U7345 (N_7345,N_3885,N_504);
nand U7346 (N_7346,N_973,N_5659);
nor U7347 (N_7347,N_500,N_1851);
nor U7348 (N_7348,N_3777,N_236);
or U7349 (N_7349,N_2740,N_4639);
or U7350 (N_7350,N_1530,N_4153);
nor U7351 (N_7351,N_663,N_1367);
xor U7352 (N_7352,N_5560,N_2589);
nor U7353 (N_7353,N_2820,N_3727);
xor U7354 (N_7354,N_3710,N_71);
xnor U7355 (N_7355,N_454,N_3268);
nand U7356 (N_7356,N_4761,N_1948);
or U7357 (N_7357,N_4597,N_2473);
or U7358 (N_7358,N_3137,N_2542);
or U7359 (N_7359,N_971,N_3022);
xnor U7360 (N_7360,N_136,N_1576);
and U7361 (N_7361,N_2623,N_963);
or U7362 (N_7362,N_1489,N_1476);
nor U7363 (N_7363,N_2224,N_2835);
nand U7364 (N_7364,N_4610,N_4127);
nand U7365 (N_7365,N_5197,N_3962);
or U7366 (N_7366,N_4586,N_3171);
and U7367 (N_7367,N_5765,N_2981);
xor U7368 (N_7368,N_1888,N_4520);
and U7369 (N_7369,N_3909,N_4762);
nand U7370 (N_7370,N_2010,N_4397);
or U7371 (N_7371,N_5953,N_2140);
and U7372 (N_7372,N_1760,N_842);
or U7373 (N_7373,N_1232,N_2509);
and U7374 (N_7374,N_2051,N_1268);
or U7375 (N_7375,N_5933,N_4455);
nand U7376 (N_7376,N_344,N_2849);
or U7377 (N_7377,N_1845,N_1272);
or U7378 (N_7378,N_3961,N_1842);
or U7379 (N_7379,N_4011,N_2534);
or U7380 (N_7380,N_2443,N_3075);
or U7381 (N_7381,N_3301,N_5280);
or U7382 (N_7382,N_2066,N_3148);
xnor U7383 (N_7383,N_5340,N_2288);
nor U7384 (N_7384,N_3997,N_778);
nand U7385 (N_7385,N_624,N_1472);
and U7386 (N_7386,N_580,N_945);
or U7387 (N_7387,N_4838,N_17);
nand U7388 (N_7388,N_2770,N_4269);
xnor U7389 (N_7389,N_131,N_3633);
nand U7390 (N_7390,N_479,N_102);
nand U7391 (N_7391,N_2661,N_3906);
or U7392 (N_7392,N_467,N_4537);
and U7393 (N_7393,N_1078,N_5724);
and U7394 (N_7394,N_794,N_4579);
xor U7395 (N_7395,N_4299,N_827);
nand U7396 (N_7396,N_4783,N_5974);
nand U7397 (N_7397,N_3488,N_2529);
or U7398 (N_7398,N_2759,N_2769);
or U7399 (N_7399,N_1689,N_3475);
xor U7400 (N_7400,N_2333,N_5823);
nand U7401 (N_7401,N_2971,N_5039);
nand U7402 (N_7402,N_2215,N_3287);
nor U7403 (N_7403,N_430,N_2571);
xor U7404 (N_7404,N_3816,N_4003);
and U7405 (N_7405,N_5886,N_3824);
xor U7406 (N_7406,N_3225,N_2523);
or U7407 (N_7407,N_2602,N_1624);
xor U7408 (N_7408,N_2221,N_1002);
or U7409 (N_7409,N_4387,N_2052);
xnor U7410 (N_7410,N_1767,N_1146);
nor U7411 (N_7411,N_4972,N_1257);
and U7412 (N_7412,N_4264,N_583);
nand U7413 (N_7413,N_2120,N_1522);
and U7414 (N_7414,N_1201,N_5590);
or U7415 (N_7415,N_2269,N_5914);
and U7416 (N_7416,N_526,N_4786);
nand U7417 (N_7417,N_127,N_5722);
and U7418 (N_7418,N_1990,N_5627);
nor U7419 (N_7419,N_1467,N_740);
nand U7420 (N_7420,N_5962,N_2701);
nor U7421 (N_7421,N_5353,N_1219);
nor U7422 (N_7422,N_2563,N_3603);
nand U7423 (N_7423,N_3991,N_395);
nor U7424 (N_7424,N_5660,N_4351);
nand U7425 (N_7425,N_3648,N_4348);
nand U7426 (N_7426,N_1444,N_4524);
nand U7427 (N_7427,N_3819,N_1408);
nor U7428 (N_7428,N_290,N_4532);
and U7429 (N_7429,N_5663,N_2878);
nand U7430 (N_7430,N_3980,N_3935);
and U7431 (N_7431,N_5239,N_4573);
nor U7432 (N_7432,N_5899,N_4089);
nand U7433 (N_7433,N_534,N_4155);
xor U7434 (N_7434,N_511,N_1139);
and U7435 (N_7435,N_5544,N_1885);
nor U7436 (N_7436,N_2522,N_1857);
or U7437 (N_7437,N_2334,N_4650);
or U7438 (N_7438,N_3917,N_4383);
and U7439 (N_7439,N_2127,N_3599);
nand U7440 (N_7440,N_568,N_1084);
nand U7441 (N_7441,N_684,N_1925);
and U7442 (N_7442,N_4712,N_5868);
nand U7443 (N_7443,N_5376,N_2348);
xor U7444 (N_7444,N_5568,N_5263);
and U7445 (N_7445,N_876,N_4603);
xnor U7446 (N_7446,N_5093,N_2196);
or U7447 (N_7447,N_3277,N_1544);
and U7448 (N_7448,N_3396,N_2969);
nand U7449 (N_7449,N_1462,N_3701);
and U7450 (N_7450,N_360,N_5125);
xor U7451 (N_7451,N_3446,N_5356);
or U7452 (N_7452,N_615,N_74);
xor U7453 (N_7453,N_3741,N_3353);
nand U7454 (N_7454,N_1615,N_932);
or U7455 (N_7455,N_3106,N_562);
nand U7456 (N_7456,N_121,N_4636);
xor U7457 (N_7457,N_5925,N_811);
nand U7458 (N_7458,N_5348,N_3325);
or U7459 (N_7459,N_4300,N_1764);
nand U7460 (N_7460,N_4177,N_2369);
and U7461 (N_7461,N_5947,N_695);
xor U7462 (N_7462,N_5997,N_4043);
and U7463 (N_7463,N_3425,N_1581);
xnor U7464 (N_7464,N_5226,N_3681);
nand U7465 (N_7465,N_782,N_3568);
xnor U7466 (N_7466,N_3158,N_4086);
nand U7467 (N_7467,N_869,N_3205);
xor U7468 (N_7468,N_3251,N_5917);
nand U7469 (N_7469,N_3650,N_667);
and U7470 (N_7470,N_4867,N_5103);
or U7471 (N_7471,N_2103,N_2287);
and U7472 (N_7472,N_3780,N_1080);
nand U7473 (N_7473,N_105,N_3539);
and U7474 (N_7474,N_3057,N_4994);
and U7475 (N_7475,N_464,N_3813);
xnor U7476 (N_7476,N_5606,N_3779);
and U7477 (N_7477,N_3812,N_958);
xnor U7478 (N_7478,N_2669,N_4572);
and U7479 (N_7479,N_5217,N_4491);
nor U7480 (N_7480,N_1308,N_3790);
xnor U7481 (N_7481,N_5623,N_4185);
nand U7482 (N_7482,N_2496,N_1553);
and U7483 (N_7483,N_4606,N_5713);
xnor U7484 (N_7484,N_896,N_1164);
and U7485 (N_7485,N_3530,N_50);
or U7486 (N_7486,N_3682,N_1231);
xnor U7487 (N_7487,N_1068,N_2142);
and U7488 (N_7488,N_1020,N_5767);
nand U7489 (N_7489,N_4660,N_75);
and U7490 (N_7490,N_2898,N_5867);
xnor U7491 (N_7491,N_2301,N_405);
nand U7492 (N_7492,N_3196,N_1244);
xnor U7493 (N_7493,N_186,N_2558);
or U7494 (N_7494,N_3018,N_3691);
nand U7495 (N_7495,N_1690,N_16);
and U7496 (N_7496,N_5622,N_591);
or U7497 (N_7497,N_2741,N_1155);
nand U7498 (N_7498,N_5378,N_1405);
nor U7499 (N_7499,N_1599,N_3706);
nand U7500 (N_7500,N_941,N_1680);
or U7501 (N_7501,N_3859,N_4453);
and U7502 (N_7502,N_4741,N_2500);
nand U7503 (N_7503,N_5821,N_1744);
and U7504 (N_7504,N_4262,N_871);
nand U7505 (N_7505,N_4218,N_638);
nand U7506 (N_7506,N_5110,N_2346);
nand U7507 (N_7507,N_2326,N_1721);
nand U7508 (N_7508,N_5631,N_1746);
xor U7509 (N_7509,N_2944,N_948);
and U7510 (N_7510,N_677,N_5171);
or U7511 (N_7511,N_3082,N_362);
nor U7512 (N_7512,N_5998,N_61);
and U7513 (N_7513,N_4022,N_1289);
xor U7514 (N_7514,N_2363,N_3070);
nand U7515 (N_7515,N_1664,N_321);
or U7516 (N_7516,N_5407,N_911);
nand U7517 (N_7517,N_1203,N_3835);
and U7518 (N_7518,N_55,N_2183);
or U7519 (N_7519,N_1116,N_4512);
nor U7520 (N_7520,N_5034,N_470);
and U7521 (N_7521,N_197,N_1707);
xor U7522 (N_7522,N_3005,N_2707);
xor U7523 (N_7523,N_4807,N_3346);
and U7524 (N_7524,N_3892,N_5291);
or U7525 (N_7525,N_1747,N_5950);
or U7526 (N_7526,N_2646,N_770);
xnor U7527 (N_7527,N_3977,N_5317);
nor U7528 (N_7528,N_3507,N_5308);
and U7529 (N_7529,N_5989,N_4970);
and U7530 (N_7530,N_2937,N_1285);
xor U7531 (N_7531,N_325,N_2110);
nand U7532 (N_7532,N_1083,N_634);
nand U7533 (N_7533,N_2677,N_3865);
or U7534 (N_7534,N_2447,N_5968);
nor U7535 (N_7535,N_2253,N_3419);
or U7536 (N_7536,N_719,N_1315);
xor U7537 (N_7537,N_521,N_3423);
and U7538 (N_7538,N_5894,N_3166);
nor U7539 (N_7539,N_1655,N_6);
or U7540 (N_7540,N_5954,N_3433);
nand U7541 (N_7541,N_2098,N_4392);
and U7542 (N_7542,N_1610,N_208);
nor U7543 (N_7543,N_4240,N_4954);
nor U7544 (N_7544,N_3615,N_5282);
nand U7545 (N_7545,N_1388,N_2983);
nor U7546 (N_7546,N_4568,N_5357);
nand U7547 (N_7547,N_579,N_418);
nor U7548 (N_7548,N_10,N_4200);
and U7549 (N_7549,N_2490,N_602);
or U7550 (N_7550,N_5662,N_3588);
or U7551 (N_7551,N_38,N_952);
nor U7552 (N_7552,N_5652,N_2889);
or U7553 (N_7553,N_5864,N_4148);
nor U7554 (N_7554,N_3320,N_3295);
nand U7555 (N_7555,N_5839,N_4721);
and U7556 (N_7556,N_4191,N_5266);
nor U7557 (N_7557,N_2929,N_5301);
xnor U7558 (N_7558,N_1066,N_915);
or U7559 (N_7559,N_3924,N_5681);
and U7560 (N_7560,N_2145,N_2845);
and U7561 (N_7561,N_381,N_681);
or U7562 (N_7562,N_1975,N_2642);
nand U7563 (N_7563,N_3749,N_2389);
and U7564 (N_7564,N_1296,N_1328);
and U7565 (N_7565,N_1923,N_5751);
or U7566 (N_7566,N_3224,N_4843);
xnor U7567 (N_7567,N_5866,N_3658);
xnor U7568 (N_7568,N_111,N_1425);
and U7569 (N_7569,N_600,N_241);
nor U7570 (N_7570,N_5423,N_4232);
and U7571 (N_7571,N_5307,N_3807);
and U7572 (N_7572,N_1943,N_2920);
nand U7573 (N_7573,N_4408,N_2605);
nor U7574 (N_7574,N_2705,N_2122);
xnor U7575 (N_7575,N_3550,N_5054);
xor U7576 (N_7576,N_1566,N_4413);
nor U7577 (N_7577,N_2497,N_1734);
xnor U7578 (N_7578,N_2355,N_1920);
and U7579 (N_7579,N_351,N_4050);
and U7580 (N_7580,N_3931,N_3849);
nand U7581 (N_7581,N_421,N_5132);
nand U7582 (N_7582,N_3940,N_844);
xor U7583 (N_7583,N_1465,N_2514);
nand U7584 (N_7584,N_4559,N_5256);
xnor U7585 (N_7585,N_1382,N_5173);
or U7586 (N_7586,N_1717,N_1200);
and U7587 (N_7587,N_5984,N_3703);
xnor U7588 (N_7588,N_3016,N_2624);
or U7589 (N_7589,N_2960,N_4144);
and U7590 (N_7590,N_1181,N_5903);
or U7591 (N_7591,N_680,N_1132);
or U7592 (N_7592,N_4414,N_1786);
xnor U7593 (N_7593,N_5099,N_3128);
or U7594 (N_7594,N_4869,N_3314);
nor U7595 (N_7595,N_5260,N_3202);
or U7596 (N_7596,N_2479,N_4981);
or U7597 (N_7597,N_5626,N_2639);
and U7598 (N_7598,N_749,N_1344);
nor U7599 (N_7599,N_2290,N_3795);
nor U7600 (N_7600,N_3557,N_1993);
or U7601 (N_7601,N_2709,N_5258);
nor U7602 (N_7602,N_2973,N_1247);
nand U7603 (N_7603,N_4060,N_813);
xor U7604 (N_7604,N_1543,N_2205);
and U7605 (N_7605,N_4669,N_3700);
or U7606 (N_7606,N_5697,N_115);
nor U7607 (N_7607,N_468,N_3063);
and U7608 (N_7608,N_5499,N_4837);
and U7609 (N_7609,N_1398,N_5252);
xnor U7610 (N_7610,N_4469,N_5834);
or U7611 (N_7611,N_5918,N_991);
or U7612 (N_7612,N_5004,N_5678);
nor U7613 (N_7613,N_1260,N_2436);
xor U7614 (N_7614,N_3447,N_5005);
nand U7615 (N_7615,N_4923,N_3096);
and U7616 (N_7616,N_2676,N_5809);
or U7617 (N_7617,N_2305,N_3051);
nor U7618 (N_7618,N_4034,N_4871);
nor U7619 (N_7619,N_4039,N_1499);
xnor U7620 (N_7620,N_4633,N_3728);
nor U7621 (N_7621,N_384,N_1362);
or U7622 (N_7622,N_2840,N_1779);
nor U7623 (N_7623,N_225,N_5095);
and U7624 (N_7624,N_4707,N_5646);
nor U7625 (N_7625,N_4857,N_795);
nor U7626 (N_7626,N_2439,N_2001);
nor U7627 (N_7627,N_618,N_4513);
nand U7628 (N_7628,N_2232,N_3776);
or U7629 (N_7629,N_5538,N_4686);
xnor U7630 (N_7630,N_5508,N_3901);
nand U7631 (N_7631,N_2992,N_2801);
or U7632 (N_7632,N_1722,N_4460);
nor U7633 (N_7633,N_1095,N_2780);
nor U7634 (N_7634,N_3735,N_4476);
xor U7635 (N_7635,N_1007,N_943);
and U7636 (N_7636,N_289,N_5324);
nand U7637 (N_7637,N_3007,N_4682);
and U7638 (N_7638,N_1293,N_2068);
or U7639 (N_7639,N_1965,N_3641);
nor U7640 (N_7640,N_733,N_1307);
or U7641 (N_7641,N_1389,N_3504);
nor U7642 (N_7642,N_143,N_5617);
or U7643 (N_7643,N_1580,N_4158);
nand U7644 (N_7644,N_2528,N_2344);
nand U7645 (N_7645,N_1986,N_3771);
xnor U7646 (N_7646,N_48,N_2696);
or U7647 (N_7647,N_4776,N_5153);
nand U7648 (N_7648,N_3228,N_5370);
nor U7649 (N_7649,N_5128,N_578);
or U7650 (N_7650,N_4810,N_2073);
nor U7651 (N_7651,N_1951,N_4479);
or U7652 (N_7652,N_984,N_5238);
nor U7653 (N_7653,N_5649,N_170);
xnor U7654 (N_7654,N_3497,N_5113);
nand U7655 (N_7655,N_2819,N_2830);
or U7656 (N_7656,N_5600,N_3850);
or U7657 (N_7657,N_2647,N_1660);
nor U7658 (N_7658,N_494,N_3721);
nor U7659 (N_7659,N_1518,N_2597);
and U7660 (N_7660,N_1783,N_4613);
xnor U7661 (N_7661,N_5009,N_1038);
xnor U7662 (N_7662,N_1278,N_2499);
nand U7663 (N_7663,N_569,N_5366);
or U7664 (N_7664,N_554,N_5946);
nand U7665 (N_7665,N_4367,N_890);
or U7666 (N_7666,N_3264,N_5072);
and U7667 (N_7667,N_2572,N_5270);
nor U7668 (N_7668,N_5381,N_3645);
and U7669 (N_7669,N_4117,N_320);
and U7670 (N_7670,N_3178,N_4908);
or U7671 (N_7671,N_3974,N_198);
and U7672 (N_7672,N_5847,N_4018);
nand U7673 (N_7673,N_5175,N_3761);
nand U7674 (N_7674,N_2274,N_1919);
xor U7675 (N_7675,N_4724,N_2620);
nand U7676 (N_7676,N_263,N_1429);
or U7677 (N_7677,N_5826,N_4250);
and U7678 (N_7678,N_3765,N_1463);
xor U7679 (N_7679,N_1183,N_108);
and U7680 (N_7680,N_5591,N_429);
nand U7681 (N_7681,N_2329,N_5209);
nand U7682 (N_7682,N_1442,N_5170);
nand U7683 (N_7683,N_2832,N_1176);
or U7684 (N_7684,N_5973,N_3129);
nand U7685 (N_7685,N_5657,N_4189);
nand U7686 (N_7686,N_308,N_179);
nor U7687 (N_7687,N_1014,N_5619);
and U7688 (N_7688,N_753,N_4171);
nand U7689 (N_7689,N_762,N_5661);
xor U7690 (N_7690,N_910,N_3554);
or U7691 (N_7691,N_4373,N_3907);
xor U7692 (N_7692,N_981,N_437);
nand U7693 (N_7693,N_4498,N_3332);
nor U7694 (N_7694,N_3680,N_5079);
xor U7695 (N_7695,N_3141,N_4196);
nand U7696 (N_7696,N_1788,N_4611);
xor U7697 (N_7697,N_3614,N_5060);
nor U7698 (N_7698,N_1258,N_2042);
nand U7699 (N_7699,N_4329,N_856);
xnor U7700 (N_7700,N_4931,N_3649);
and U7701 (N_7701,N_5877,N_1174);
and U7702 (N_7702,N_4894,N_3364);
nand U7703 (N_7703,N_5542,N_4797);
nor U7704 (N_7704,N_3382,N_4468);
or U7705 (N_7705,N_3545,N_2526);
and U7706 (N_7706,N_5587,N_5453);
or U7707 (N_7707,N_4888,N_5671);
nor U7708 (N_7708,N_5537,N_3915);
xor U7709 (N_7709,N_361,N_4566);
or U7710 (N_7710,N_3690,N_1575);
nand U7711 (N_7711,N_5796,N_1486);
and U7712 (N_7712,N_1889,N_1693);
nand U7713 (N_7713,N_4302,N_750);
xor U7714 (N_7714,N_1324,N_2880);
nand U7715 (N_7715,N_4307,N_4091);
or U7716 (N_7716,N_1461,N_4249);
xor U7717 (N_7717,N_5501,N_4991);
or U7718 (N_7718,N_4107,N_509);
or U7719 (N_7719,N_3309,N_137);
or U7720 (N_7720,N_1740,N_3553);
or U7721 (N_7721,N_5042,N_4668);
xnor U7722 (N_7722,N_2357,N_1561);
nor U7723 (N_7723,N_1355,N_2859);
or U7724 (N_7724,N_4198,N_4919);
xor U7725 (N_7725,N_1346,N_797);
xnor U7726 (N_7726,N_5647,N_5478);
xnor U7727 (N_7727,N_2585,N_1510);
and U7728 (N_7728,N_196,N_708);
and U7729 (N_7729,N_1477,N_459);
xnor U7730 (N_7730,N_1521,N_1333);
xnor U7731 (N_7731,N_2434,N_3796);
and U7732 (N_7732,N_4258,N_4452);
and U7733 (N_7733,N_3413,N_3317);
or U7734 (N_7734,N_4343,N_3200);
nand U7735 (N_7735,N_5248,N_3851);
nand U7736 (N_7736,N_5101,N_604);
xnor U7737 (N_7737,N_1559,N_3621);
nor U7738 (N_7738,N_2121,N_2128);
and U7739 (N_7739,N_1045,N_4388);
or U7740 (N_7740,N_576,N_3409);
nor U7741 (N_7741,N_3043,N_5057);
and U7742 (N_7742,N_4233,N_2330);
and U7743 (N_7743,N_2955,N_326);
nor U7744 (N_7744,N_1234,N_2003);
nor U7745 (N_7745,N_5934,N_3781);
or U7746 (N_7746,N_3150,N_1538);
and U7747 (N_7747,N_4974,N_841);
xor U7748 (N_7748,N_4097,N_5247);
xor U7749 (N_7749,N_4220,N_4421);
nand U7750 (N_7750,N_5475,N_2679);
xor U7751 (N_7751,N_242,N_1780);
and U7752 (N_7752,N_3281,N_126);
xor U7753 (N_7753,N_3782,N_5735);
xnor U7754 (N_7754,N_1345,N_5778);
nand U7755 (N_7755,N_5069,N_2332);
and U7756 (N_7756,N_3477,N_1003);
xnor U7757 (N_7757,N_2851,N_2668);
or U7758 (N_7758,N_2,N_4937);
nand U7759 (N_7759,N_3253,N_988);
or U7760 (N_7760,N_57,N_3868);
or U7761 (N_7761,N_1687,N_1964);
or U7762 (N_7762,N_3591,N_860);
nand U7763 (N_7763,N_4315,N_4276);
and U7764 (N_7764,N_3212,N_4906);
and U7765 (N_7765,N_857,N_2307);
nor U7766 (N_7766,N_1196,N_5775);
or U7767 (N_7767,N_1546,N_893);
or U7768 (N_7768,N_1502,N_1);
or U7769 (N_7769,N_139,N_1393);
and U7770 (N_7770,N_1458,N_2976);
or U7771 (N_7771,N_2241,N_4739);
nand U7772 (N_7772,N_2767,N_2418);
nor U7773 (N_7773,N_989,N_4764);
and U7774 (N_7774,N_3979,N_2037);
nand U7775 (N_7775,N_1626,N_901);
xnor U7776 (N_7776,N_1795,N_42);
and U7777 (N_7777,N_363,N_2378);
nor U7778 (N_7778,N_5284,N_3260);
or U7779 (N_7779,N_4848,N_331);
nor U7780 (N_7780,N_2674,N_565);
and U7781 (N_7781,N_2673,N_1912);
xnor U7782 (N_7782,N_570,N_5579);
nor U7783 (N_7783,N_2833,N_5983);
nand U7784 (N_7784,N_4239,N_887);
nand U7785 (N_7785,N_4059,N_555);
nand U7786 (N_7786,N_2865,N_3541);
nor U7787 (N_7787,N_2295,N_5424);
xor U7788 (N_7788,N_1848,N_769);
nor U7789 (N_7789,N_366,N_1870);
nand U7790 (N_7790,N_5035,N_2396);
xnor U7791 (N_7791,N_3384,N_2536);
nand U7792 (N_7792,N_2292,N_1692);
nand U7793 (N_7793,N_1871,N_5958);
and U7794 (N_7794,N_376,N_4483);
nand U7795 (N_7795,N_3654,N_909);
nor U7796 (N_7796,N_4384,N_3994);
and U7797 (N_7797,N_4514,N_3015);
and U7798 (N_7798,N_5500,N_1074);
or U7799 (N_7799,N_2058,N_3957);
and U7800 (N_7800,N_4952,N_4677);
xor U7801 (N_7801,N_2323,N_4788);
or U7802 (N_7802,N_5792,N_1775);
and U7803 (N_7803,N_3375,N_3094);
nor U7804 (N_7804,N_256,N_2811);
nand U7805 (N_7805,N_3995,N_2596);
nor U7806 (N_7806,N_3078,N_3923);
and U7807 (N_7807,N_4314,N_5744);
nor U7808 (N_7808,N_1438,N_146);
or U7809 (N_7809,N_4992,N_959);
or U7810 (N_7810,N_4423,N_5969);
nand U7811 (N_7811,N_4702,N_410);
or U7812 (N_7812,N_5824,N_4522);
nand U7813 (N_7813,N_3912,N_505);
nand U7814 (N_7814,N_4950,N_617);
nor U7815 (N_7815,N_33,N_1507);
xnor U7816 (N_7816,N_1649,N_1048);
nor U7817 (N_7817,N_191,N_5106);
nor U7818 (N_7818,N_3836,N_5347);
and U7819 (N_7819,N_3818,N_3124);
nand U7820 (N_7820,N_1824,N_3605);
xor U7821 (N_7821,N_3142,N_231);
and U7822 (N_7822,N_4416,N_5150);
nor U7823 (N_7823,N_5192,N_834);
and U7824 (N_7824,N_4213,N_2331);
or U7825 (N_7825,N_2217,N_2444);
nor U7826 (N_7826,N_1918,N_2533);
and U7827 (N_7827,N_4290,N_3133);
nor U7828 (N_7828,N_3339,N_5668);
or U7829 (N_7829,N_990,N_2306);
and U7830 (N_7830,N_4273,N_2213);
and U7831 (N_7831,N_4618,N_3496);
xnor U7832 (N_7832,N_5312,N_1911);
or U7833 (N_7833,N_4745,N_281);
and U7834 (N_7834,N_3058,N_689);
and U7835 (N_7835,N_3465,N_457);
nor U7836 (N_7836,N_1317,N_1528);
nor U7837 (N_7837,N_3738,N_5730);
or U7838 (N_7838,N_2754,N_193);
nor U7839 (N_7839,N_4292,N_889);
or U7840 (N_7840,N_5022,N_2544);
xnor U7841 (N_7841,N_4756,N_4684);
xor U7842 (N_7842,N_3298,N_3412);
nand U7843 (N_7843,N_5085,N_2211);
and U7844 (N_7844,N_3407,N_2860);
xor U7845 (N_7845,N_491,N_1794);
nand U7846 (N_7846,N_1512,N_2805);
or U7847 (N_7847,N_5156,N_4609);
nand U7848 (N_7848,N_2548,N_2530);
or U7849 (N_7849,N_3265,N_233);
nor U7850 (N_7850,N_3604,N_830);
and U7851 (N_7851,N_2710,N_5198);
and U7852 (N_7852,N_4718,N_2913);
nor U7853 (N_7853,N_3668,N_2393);
or U7854 (N_7854,N_1341,N_925);
nand U7855 (N_7855,N_2852,N_2294);
nand U7856 (N_7856,N_4285,N_897);
and U7857 (N_7857,N_2637,N_4775);
xor U7858 (N_7858,N_4375,N_2193);
nand U7859 (N_7859,N_4431,N_1855);
nor U7860 (N_7860,N_2448,N_235);
and U7861 (N_7861,N_5020,N_4629);
nor U7862 (N_7862,N_5168,N_1214);
nand U7863 (N_7863,N_5261,N_2546);
nand U7864 (N_7864,N_3805,N_557);
xnor U7865 (N_7865,N_2643,N_158);
xor U7866 (N_7866,N_845,N_2782);
nand U7867 (N_7867,N_2644,N_2968);
nor U7868 (N_7868,N_835,N_2785);
nor U7869 (N_7869,N_1071,N_2671);
nand U7870 (N_7870,N_4057,N_5201);
nand U7871 (N_7871,N_3972,N_3876);
nor U7872 (N_7872,N_5555,N_5130);
xnor U7873 (N_7873,N_829,N_992);
xnor U7874 (N_7874,N_2839,N_2923);
or U7875 (N_7875,N_3429,N_1708);
nand U7876 (N_7876,N_1696,N_2252);
or U7877 (N_7877,N_1040,N_5610);
nand U7878 (N_7878,N_123,N_4614);
nand U7879 (N_7879,N_3725,N_5467);
nand U7880 (N_7880,N_5321,N_1070);
xnor U7881 (N_7881,N_133,N_5272);
nand U7882 (N_7882,N_5051,N_4306);
or U7883 (N_7883,N_187,N_1400);
and U7884 (N_7884,N_4490,N_4077);
and U7885 (N_7885,N_545,N_5753);
nor U7886 (N_7886,N_1357,N_3318);
xor U7887 (N_7887,N_5639,N_784);
nand U7888 (N_7888,N_1629,N_1552);
and U7889 (N_7889,N_311,N_3854);
and U7890 (N_7890,N_4323,N_2722);
xor U7891 (N_7891,N_2195,N_3492);
nor U7892 (N_7892,N_1623,N_4112);
and U7893 (N_7893,N_5745,N_3683);
and U7894 (N_7894,N_4228,N_3273);
nand U7895 (N_7895,N_3522,N_1283);
and U7896 (N_7896,N_706,N_1238);
nand U7897 (N_7897,N_1184,N_423);
nor U7898 (N_7898,N_3073,N_5583);
or U7899 (N_7899,N_1803,N_1843);
xor U7900 (N_7900,N_5520,N_1896);
or U7901 (N_7901,N_682,N_3406);
nor U7902 (N_7902,N_4763,N_4754);
or U7903 (N_7903,N_3531,N_3089);
nand U7904 (N_7904,N_5999,N_926);
nand U7905 (N_7905,N_962,N_3181);
xor U7906 (N_7906,N_125,N_1316);
and U7907 (N_7907,N_4996,N_5789);
or U7908 (N_7908,N_4000,N_4482);
xnor U7909 (N_7909,N_2877,N_4391);
or U7910 (N_7910,N_3187,N_1031);
xnor U7911 (N_7911,N_5274,N_1715);
nor U7912 (N_7912,N_1834,N_523);
xor U7913 (N_7913,N_1909,N_3112);
xnor U7914 (N_7914,N_1027,N_4853);
nor U7915 (N_7915,N_359,N_1757);
and U7916 (N_7916,N_2250,N_3584);
nand U7917 (N_7917,N_3733,N_2199);
nor U7918 (N_7918,N_145,N_3348);
nor U7919 (N_7919,N_2231,N_5776);
nor U7920 (N_7920,N_629,N_2658);
or U7921 (N_7921,N_291,N_4901);
xnor U7922 (N_7922,N_3867,N_1339);
nor U7923 (N_7923,N_5535,N_2431);
and U7924 (N_7924,N_432,N_3964);
xnor U7925 (N_7925,N_4101,N_4449);
or U7926 (N_7926,N_7,N_4631);
nor U7927 (N_7927,N_1669,N_5788);
nand U7928 (N_7928,N_2694,N_3144);
and U7929 (N_7929,N_451,N_5399);
or U7930 (N_7930,N_4052,N_1773);
or U7931 (N_7931,N_707,N_5460);
nor U7932 (N_7932,N_247,N_5165);
nor U7933 (N_7933,N_4136,N_5975);
and U7934 (N_7934,N_5033,N_5906);
nand U7935 (N_7935,N_5907,N_1321);
nor U7936 (N_7936,N_852,N_2350);
and U7937 (N_7937,N_5850,N_796);
or U7938 (N_7938,N_3708,N_5385);
and U7939 (N_7939,N_4644,N_5377);
nand U7940 (N_7940,N_1125,N_4634);
nor U7941 (N_7941,N_4162,N_3729);
and U7942 (N_7942,N_2039,N_2957);
xor U7943 (N_7943,N_1273,N_1350);
or U7944 (N_7944,N_2603,N_4199);
or U7945 (N_7945,N_3299,N_2325);
nand U7946 (N_7946,N_2891,N_2130);
nor U7947 (N_7947,N_1770,N_3090);
and U7948 (N_7948,N_662,N_5875);
and U7949 (N_7949,N_1081,N_5705);
nor U7950 (N_7950,N_4584,N_1755);
and U7951 (N_7951,N_783,N_5220);
nand U7952 (N_7952,N_5586,N_5471);
nand U7953 (N_7953,N_2361,N_3338);
nor U7954 (N_7954,N_2747,N_5856);
nand U7955 (N_7955,N_4626,N_1602);
and U7956 (N_7956,N_1241,N_635);
or U7957 (N_7957,N_628,N_5512);
xor U7958 (N_7958,N_77,N_1172);
and U7959 (N_7959,N_286,N_519);
xor U7960 (N_7960,N_2087,N_3050);
xnor U7961 (N_7961,N_87,N_4244);
nor U7962 (N_7962,N_4518,N_2584);
and U7963 (N_7963,N_3889,N_5119);
and U7964 (N_7964,N_1397,N_3783);
or U7965 (N_7965,N_2309,N_3842);
or U7966 (N_7966,N_626,N_1124);
nand U7967 (N_7967,N_65,N_5701);
nor U7968 (N_7968,N_5480,N_1758);
nor U7969 (N_7969,N_2853,N_5147);
nand U7970 (N_7970,N_5869,N_5629);
xor U7971 (N_7971,N_3634,N_5980);
and U7972 (N_7972,N_5303,N_2730);
and U7973 (N_7973,N_721,N_4887);
nor U7974 (N_7974,N_1360,N_5208);
and U7975 (N_7975,N_4560,N_3321);
nand U7976 (N_7976,N_2697,N_3944);
or U7977 (N_7977,N_2450,N_4404);
nand U7978 (N_7978,N_5963,N_2553);
and U7979 (N_7979,N_195,N_2268);
nand U7980 (N_7980,N_937,N_1897);
nand U7981 (N_7981,N_34,N_5450);
nand U7982 (N_7982,N_3415,N_4231);
and U7983 (N_7983,N_1607,N_3480);
or U7984 (N_7984,N_431,N_4855);
xnor U7985 (N_7985,N_1815,N_5609);
and U7986 (N_7986,N_3293,N_1524);
xor U7987 (N_7987,N_3053,N_1148);
and U7988 (N_7988,N_1950,N_1297);
xor U7989 (N_7989,N_4977,N_1102);
nor U7990 (N_7990,N_3354,N_3596);
xor U7991 (N_7991,N_1150,N_581);
and U7992 (N_7992,N_4965,N_5798);
nor U7993 (N_7993,N_4771,N_3939);
xor U7994 (N_7994,N_594,N_5174);
nand U7995 (N_7995,N_669,N_5267);
and U7996 (N_7996,N_4817,N_5000);
xor U7997 (N_7997,N_4840,N_773);
and U7998 (N_7998,N_994,N_1821);
nand U7999 (N_7999,N_3535,N_3748);
nand U8000 (N_8000,N_2070,N_3288);
and U8001 (N_8001,N_808,N_5716);
xnor U8002 (N_8002,N_402,N_2470);
or U8003 (N_8003,N_5721,N_4374);
or U8004 (N_8004,N_2392,N_3207);
or U8005 (N_8005,N_8,N_2683);
nand U8006 (N_8006,N_5588,N_412);
and U8007 (N_8007,N_3509,N_3711);
nand U8008 (N_8008,N_854,N_4526);
xor U8009 (N_8009,N_3525,N_5134);
nor U8010 (N_8010,N_2218,N_1358);
nor U8011 (N_8011,N_1958,N_328);
and U8012 (N_8012,N_4473,N_3983);
xor U8013 (N_8013,N_5419,N_2359);
xnor U8014 (N_8014,N_5397,N_3113);
or U8015 (N_8015,N_5898,N_1533);
and U8016 (N_8016,N_1366,N_964);
xor U8017 (N_8017,N_5498,N_1491);
xor U8018 (N_8018,N_1434,N_285);
xnor U8019 (N_8019,N_5186,N_4137);
xor U8020 (N_8020,N_1137,N_2200);
and U8021 (N_8021,N_337,N_2930);
or U8022 (N_8022,N_5563,N_3947);
nand U8023 (N_8023,N_4357,N_4588);
nor U8024 (N_8024,N_2459,N_3925);
and U8025 (N_8025,N_5723,N_791);
and U8026 (N_8026,N_5302,N_4732);
and U8027 (N_8027,N_3884,N_1526);
xor U8028 (N_8028,N_1643,N_2101);
nor U8029 (N_8029,N_5289,N_5071);
or U8030 (N_8030,N_5432,N_3670);
xnor U8031 (N_8031,N_744,N_3319);
xnor U8032 (N_8032,N_2951,N_1061);
nor U8033 (N_8033,N_5194,N_4298);
xor U8034 (N_8034,N_2257,N_2604);
and U8035 (N_8035,N_5094,N_1646);
and U8036 (N_8036,N_2021,N_2617);
nor U8037 (N_8037,N_3215,N_5761);
xnor U8038 (N_8038,N_1598,N_3084);
nor U8039 (N_8039,N_2713,N_4944);
xor U8040 (N_8040,N_4781,N_2902);
nor U8041 (N_8041,N_1460,N_5112);
nor U8042 (N_8042,N_1886,N_5897);
or U8043 (N_8043,N_3125,N_3438);
and U8044 (N_8044,N_919,N_2715);
nor U8045 (N_8045,N_1960,N_1571);
and U8046 (N_8046,N_1329,N_5155);
nor U8047 (N_8047,N_870,N_5073);
xnor U8048 (N_8048,N_3476,N_3988);
nor U8049 (N_8049,N_587,N_239);
nor U8050 (N_8050,N_1579,N_4461);
xnor U8051 (N_8051,N_2886,N_790);
nor U8052 (N_8052,N_4450,N_5781);
nand U8053 (N_8053,N_590,N_5862);
nor U8054 (N_8054,N_1233,N_1766);
nor U8055 (N_8055,N_2946,N_5979);
xnor U8056 (N_8056,N_5786,N_3759);
nor U8057 (N_8057,N_704,N_4796);
nand U8058 (N_8058,N_1525,N_5760);
xor U8059 (N_8059,N_987,N_2586);
nor U8060 (N_8060,N_4773,N_4907);
nor U8061 (N_8061,N_2776,N_5683);
xor U8062 (N_8062,N_2778,N_726);
nand U8063 (N_8063,N_382,N_3216);
nor U8064 (N_8064,N_1342,N_9);
and U8065 (N_8065,N_1445,N_998);
and U8066 (N_8066,N_2945,N_5820);
and U8067 (N_8067,N_2828,N_317);
nor U8068 (N_8068,N_5144,N_5698);
or U8069 (N_8069,N_5521,N_5567);
nor U8070 (N_8070,N_4973,N_4206);
nand U8071 (N_8071,N_5359,N_4246);
and U8072 (N_8072,N_862,N_1112);
and U8073 (N_8073,N_742,N_2308);
nand U8074 (N_8074,N_2501,N_5010);
or U8075 (N_8075,N_1459,N_4106);
or U8076 (N_8076,N_1422,N_5727);
xnor U8077 (N_8077,N_1606,N_4648);
or U8078 (N_8078,N_228,N_2451);
nand U8079 (N_8079,N_4402,N_4750);
xor U8080 (N_8080,N_3914,N_3201);
xor U8081 (N_8081,N_5892,N_4889);
and U8082 (N_8082,N_5468,N_469);
or U8083 (N_8083,N_3060,N_996);
xnor U8084 (N_8084,N_4703,N_3292);
or U8085 (N_8085,N_5939,N_2345);
and U8086 (N_8086,N_2391,N_5799);
nor U8087 (N_8087,N_3283,N_5680);
nand U8088 (N_8088,N_4928,N_5027);
nand U8089 (N_8089,N_4013,N_4915);
or U8090 (N_8090,N_4448,N_2349);
or U8091 (N_8091,N_5759,N_4456);
nand U8092 (N_8092,N_453,N_2954);
or U8093 (N_8093,N_1094,N_4470);
nor U8094 (N_8094,N_1484,N_5196);
and U8095 (N_8095,N_2579,N_4735);
and U8096 (N_8096,N_3934,N_5409);
xor U8097 (N_8097,N_5361,N_3410);
and U8098 (N_8098,N_3799,N_1542);
xor U8099 (N_8099,N_3368,N_1464);
or U8100 (N_8100,N_1399,N_4641);
or U8101 (N_8101,N_5420,N_2806);
nor U8102 (N_8102,N_4435,N_2311);
or U8103 (N_8103,N_450,N_3436);
nand U8104 (N_8104,N_4139,N_2318);
nand U8105 (N_8105,N_4555,N_1217);
nor U8106 (N_8106,N_3214,N_1310);
xnor U8107 (N_8107,N_3097,N_2157);
xor U8108 (N_8108,N_4129,N_5955);
and U8109 (N_8109,N_1688,N_3463);
or U8110 (N_8110,N_3636,N_76);
nand U8111 (N_8111,N_1711,N_4897);
nand U8112 (N_8112,N_2555,N_3025);
or U8113 (N_8113,N_650,N_1612);
or U8114 (N_8114,N_824,N_1414);
xor U8115 (N_8115,N_977,N_1995);
nand U8116 (N_8116,N_4271,N_1589);
nor U8117 (N_8117,N_2057,N_532);
nor U8118 (N_8118,N_3823,N_5967);
nand U8119 (N_8119,N_3218,N_596);
nand U8120 (N_8120,N_3491,N_2712);
or U8121 (N_8121,N_2381,N_116);
or U8122 (N_8122,N_5477,N_5599);
nor U8123 (N_8123,N_3307,N_3597);
and U8124 (N_8124,N_2435,N_172);
nand U8125 (N_8125,N_3242,N_1850);
and U8126 (N_8126,N_810,N_2277);
or U8127 (N_8127,N_162,N_5494);
nand U8128 (N_8128,N_5613,N_5922);
or U8129 (N_8129,N_2011,N_558);
or U8130 (N_8130,N_5912,N_1481);
xnor U8131 (N_8131,N_4662,N_4590);
and U8132 (N_8132,N_4963,N_4349);
nand U8133 (N_8133,N_5770,N_497);
and U8134 (N_8134,N_5162,N_2452);
or U8135 (N_8135,N_1090,N_3904);
nand U8136 (N_8136,N_2690,N_1136);
nor U8137 (N_8137,N_1771,N_1212);
and U8138 (N_8138,N_3355,N_1865);
nor U8139 (N_8139,N_894,N_3437);
and U8140 (N_8140,N_4393,N_4385);
or U8141 (N_8141,N_5638,N_3897);
nand U8142 (N_8142,N_496,N_4028);
and U8143 (N_8143,N_4283,N_3383);
xnor U8144 (N_8144,N_3285,N_3862);
xnor U8145 (N_8145,N_3560,N_3843);
or U8146 (N_8146,N_5710,N_4308);
and U8147 (N_8147,N_5413,N_2652);
xor U8148 (N_8148,N_3457,N_1810);
nor U8149 (N_8149,N_357,N_2922);
xor U8150 (N_8150,N_3815,N_1658);
or U8151 (N_8151,N_5971,N_2398);
xnor U8152 (N_8152,N_5318,N_4547);
and U8153 (N_8153,N_3878,N_1631);
nor U8154 (N_8154,N_2773,N_1277);
nor U8155 (N_8155,N_2320,N_3844);
or U8156 (N_8156,N_3263,N_1056);
nor U8157 (N_8157,N_2520,N_4291);
xnor U8158 (N_8158,N_4851,N_5091);
xnor U8159 (N_8159,N_1641,N_4234);
xor U8160 (N_8160,N_2924,N_1868);
nor U8161 (N_8161,N_3469,N_2055);
nand U8162 (N_8162,N_5199,N_5525);
nor U8163 (N_8163,N_5440,N_553);
xnor U8164 (N_8164,N_5747,N_4628);
and U8165 (N_8165,N_3577,N_5205);
or U8166 (N_8166,N_1652,N_1724);
nand U8167 (N_8167,N_5219,N_175);
nor U8168 (N_8168,N_3808,N_3764);
nor U8169 (N_8169,N_2342,N_3967);
nand U8170 (N_8170,N_4812,N_825);
nand U8171 (N_8171,N_954,N_5068);
nor U8172 (N_8172,N_1727,N_5527);
or U8173 (N_8173,N_2380,N_2879);
nor U8174 (N_8174,N_489,N_1728);
nand U8175 (N_8175,N_3453,N_3873);
xor U8176 (N_8176,N_643,N_4268);
and U8177 (N_8177,N_1977,N_5314);
xor U8178 (N_8178,N_4692,N_2895);
xnor U8179 (N_8179,N_3360,N_5893);
nand U8180 (N_8180,N_5369,N_3458);
and U8181 (N_8181,N_1496,N_37);
nor U8182 (N_8182,N_5225,N_701);
nor U8183 (N_8183,N_4146,N_1216);
and U8184 (N_8184,N_5276,N_1991);
xor U8185 (N_8185,N_3717,N_336);
nand U8186 (N_8186,N_3852,N_2180);
nand U8187 (N_8187,N_4911,N_3564);
nand U8188 (N_8188,N_1169,N_4652);
nor U8189 (N_8189,N_3290,N_3992);
nand U8190 (N_8190,N_206,N_3589);
and U8191 (N_8191,N_5858,N_3758);
and U8192 (N_8192,N_2503,N_1613);
nand U8193 (N_8193,N_3976,N_816);
nand U8194 (N_8194,N_3366,N_157);
nand U8195 (N_8195,N_3874,N_2856);
xor U8196 (N_8196,N_3785,N_417);
or U8197 (N_8197,N_1967,N_3503);
nand U8198 (N_8198,N_4545,N_5656);
or U8199 (N_8199,N_4805,N_4204);
xor U8200 (N_8200,N_1079,N_3565);
xor U8201 (N_8201,N_2293,N_4819);
nor U8202 (N_8202,N_1844,N_1998);
and U8203 (N_8203,N_3751,N_2177);
or U8204 (N_8204,N_1270,N_1453);
and U8205 (N_8205,N_3731,N_645);
xnor U8206 (N_8206,N_2716,N_3739);
nand U8207 (N_8207,N_2271,N_2027);
nor U8208 (N_8208,N_4123,N_3585);
and U8209 (N_8209,N_255,N_1829);
nor U8210 (N_8210,N_3164,N_1262);
and U8211 (N_8211,N_2475,N_2681);
nor U8212 (N_8212,N_4711,N_2041);
xor U8213 (N_8213,N_4390,N_4727);
xnor U8214 (N_8214,N_144,N_818);
xnor U8215 (N_8215,N_688,N_5394);
nand U8216 (N_8216,N_4217,N_2519);
xnor U8217 (N_8217,N_322,N_3259);
nor U8218 (N_8218,N_52,N_1705);
nor U8219 (N_8219,N_1617,N_1157);
and U8220 (N_8220,N_2813,N_1320);
or U8221 (N_8221,N_446,N_5871);
nand U8222 (N_8222,N_3101,N_3234);
nand U8223 (N_8223,N_1698,N_1529);
nor U8224 (N_8224,N_5689,N_606);
nor U8225 (N_8225,N_3071,N_4326);
and U8226 (N_8226,N_2622,N_1778);
and U8227 (N_8227,N_898,N_923);
nor U8228 (N_8228,N_2108,N_3177);
xor U8229 (N_8229,N_2187,N_2800);
xnor U8230 (N_8230,N_586,N_4062);
nor U8231 (N_8231,N_5522,N_4822);
or U8232 (N_8232,N_2149,N_2545);
nand U8233 (N_8233,N_5733,N_540);
and U8234 (N_8234,N_1539,N_1325);
and U8235 (N_8235,N_5688,N_1440);
or U8236 (N_8236,N_674,N_463);
nand U8237 (N_8237,N_2137,N_2423);
nor U8238 (N_8238,N_4630,N_2172);
xnor U8239 (N_8239,N_168,N_5651);
nor U8240 (N_8240,N_4679,N_1751);
or U8241 (N_8241,N_2814,N_2107);
and U8242 (N_8242,N_802,N_4494);
nand U8243 (N_8243,N_4297,N_710);
and U8244 (N_8244,N_5942,N_1075);
nand U8245 (N_8245,N_279,N_2168);
xor U8246 (N_8246,N_1322,N_280);
and U8247 (N_8247,N_3361,N_805);
or U8248 (N_8248,N_2565,N_3028);
nor U8249 (N_8249,N_5264,N_951);
or U8250 (N_8250,N_4541,N_5293);
and U8251 (N_8251,N_4670,N_567);
nor U8252 (N_8252,N_2064,N_921);
or U8253 (N_8253,N_4037,N_3791);
nor U8254 (N_8254,N_2094,N_3045);
nand U8255 (N_8255,N_4769,N_1057);
xor U8256 (N_8256,N_5562,N_4489);
or U8257 (N_8257,N_5699,N_2763);
nor U8258 (N_8258,N_4820,N_1017);
xnor U8259 (N_8259,N_4706,N_4904);
nand U8260 (N_8260,N_5254,N_3546);
xnor U8261 (N_8261,N_2635,N_5700);
or U8262 (N_8262,N_672,N_5462);
or U8263 (N_8263,N_2612,N_2044);
and U8264 (N_8264,N_3954,N_1240);
nand U8265 (N_8265,N_3111,N_355);
or U8266 (N_8266,N_4047,N_2483);
nand U8267 (N_8267,N_3936,N_4879);
and U8268 (N_8268,N_1249,N_5665);
nand U8269 (N_8269,N_3183,N_5771);
xor U8270 (N_8270,N_5493,N_4971);
or U8271 (N_8271,N_274,N_30);
xnor U8272 (N_8272,N_4436,N_1479);
xor U8273 (N_8273,N_2666,N_4924);
nand U8274 (N_8274,N_1517,N_3606);
or U8275 (N_8275,N_4683,N_4309);
and U8276 (N_8276,N_456,N_2802);
and U8277 (N_8277,N_759,N_4115);
nand U8278 (N_8278,N_756,N_905);
nand U8279 (N_8279,N_885,N_1634);
nand U8280 (N_8280,N_253,N_2239);
xor U8281 (N_8281,N_5811,N_2289);
and U8282 (N_8282,N_3179,N_3778);
xnor U8283 (N_8283,N_3610,N_1129);
and U8284 (N_8284,N_5311,N_2354);
nor U8285 (N_8285,N_2812,N_84);
nand U8286 (N_8286,N_4777,N_3241);
nand U8287 (N_8287,N_957,N_4406);
xnor U8288 (N_8288,N_4948,N_1001);
or U8289 (N_8289,N_5461,N_5797);
nor U8290 (N_8290,N_5384,N_1665);
xor U8291 (N_8291,N_1854,N_461);
xor U8292 (N_8292,N_4570,N_2698);
and U8293 (N_8293,N_4183,N_4141);
and U8294 (N_8294,N_3643,N_1301);
xor U8295 (N_8295,N_4794,N_4304);
nand U8296 (N_8296,N_3987,N_1179);
xnor U8297 (N_8297,N_2081,N_661);
or U8298 (N_8298,N_1041,N_4243);
xnor U8299 (N_8299,N_5896,N_486);
xnor U8300 (N_8300,N_3029,N_1935);
and U8301 (N_8301,N_3982,N_2834);
and U8302 (N_8302,N_3023,N_5490);
xnor U8303 (N_8303,N_1730,N_2510);
and U8304 (N_8304,N_2400,N_149);
xnor U8305 (N_8305,N_3624,N_5430);
or U8306 (N_8306,N_2621,N_5108);
nand U8307 (N_8307,N_1089,N_4508);
or U8308 (N_8308,N_1282,N_1802);
and U8309 (N_8309,N_3672,N_3746);
and U8310 (N_8310,N_1418,N_3512);
nand U8311 (N_8311,N_2150,N_3875);
and U8312 (N_8312,N_1759,N_5415);
nor U8313 (N_8313,N_2174,N_3246);
and U8314 (N_8314,N_5949,N_3161);
or U8315 (N_8315,N_700,N_2601);
nand U8316 (N_8316,N_5104,N_3417);
and U8317 (N_8317,N_5245,N_997);
and U8318 (N_8318,N_4346,N_3880);
nor U8319 (N_8319,N_304,N_3103);
nor U8320 (N_8320,N_4587,N_224);
nor U8321 (N_8321,N_5926,N_2373);
or U8322 (N_8322,N_5281,N_407);
and U8323 (N_8323,N_5221,N_1503);
nor U8324 (N_8324,N_1582,N_5806);
nand U8325 (N_8325,N_3391,N_2046);
nand U8326 (N_8326,N_4208,N_5876);
nand U8327 (N_8327,N_1413,N_305);
or U8328 (N_8328,N_3529,N_2995);
xnor U8329 (N_8329,N_1765,N_1024);
nor U8330 (N_8330,N_2240,N_1931);
nand U8331 (N_8331,N_2566,N_660);
nor U8332 (N_8332,N_2737,N_35);
nand U8333 (N_8333,N_1088,N_3378);
or U8334 (N_8334,N_5011,N_3335);
xor U8335 (N_8335,N_4704,N_2940);
and U8336 (N_8336,N_4845,N_106);
nand U8337 (N_8337,N_3256,N_1379);
nor U8338 (N_8338,N_5164,N_3766);
and U8339 (N_8339,N_5322,N_3266);
nand U8340 (N_8340,N_817,N_2430);
xor U8341 (N_8341,N_4828,N_2583);
or U8342 (N_8342,N_166,N_607);
or U8343 (N_8343,N_2827,N_1280);
nand U8344 (N_8344,N_2201,N_3334);
and U8345 (N_8345,N_5978,N_3054);
and U8346 (N_8346,N_490,N_5379);
xor U8347 (N_8347,N_4809,N_970);
and U8348 (N_8348,N_1679,N_528);
xnor U8349 (N_8349,N_3810,N_4395);
xor U8350 (N_8350,N_4678,N_814);
or U8351 (N_8351,N_588,N_4216);
and U8352 (N_8352,N_1025,N_1808);
nor U8353 (N_8353,N_5127,N_3331);
and U8354 (N_8354,N_2403,N_4830);
nand U8355 (N_8355,N_152,N_5167);
nand U8356 (N_8356,N_2703,N_1799);
xnor U8357 (N_8357,N_1891,N_4642);
nor U8358 (N_8358,N_4446,N_2552);
nor U8359 (N_8359,N_5331,N_474);
and U8360 (N_8360,N_1556,N_477);
nand U8361 (N_8361,N_3963,N_1825);
or U8362 (N_8362,N_3965,N_43);
or U8363 (N_8363,N_4223,N_524);
nor U8364 (N_8364,N_1266,N_3017);
and U8365 (N_8365,N_2178,N_2411);
nand U8366 (N_8366,N_4868,N_1969);
xnor U8367 (N_8367,N_278,N_1108);
nand U8368 (N_8368,N_4236,N_3000);
and U8369 (N_8369,N_3257,N_5484);
xor U8370 (N_8370,N_2578,N_1600);
or U8371 (N_8371,N_5719,N_5299);
nor U8372 (N_8372,N_2367,N_5728);
or U8373 (N_8373,N_1729,N_3899);
xor U8374 (N_8374,N_1789,N_2793);
nand U8375 (N_8375,N_3274,N_5887);
and U8376 (N_8376,N_4507,N_5603);
nor U8377 (N_8377,N_2511,N_1086);
and U8378 (N_8378,N_2075,N_4740);
nand U8379 (N_8379,N_1290,N_3369);
and U8380 (N_8380,N_4646,N_5808);
xor U8381 (N_8381,N_2615,N_5372);
nand U8382 (N_8382,N_4420,N_3513);
or U8383 (N_8383,N_3794,N_1982);
nor U8384 (N_8384,N_5804,N_1110);
and U8385 (N_8385,N_2303,N_380);
nor U8386 (N_8386,N_1417,N_5829);
nand U8387 (N_8387,N_4655,N_3088);
xnor U8388 (N_8388,N_5993,N_11);
nand U8389 (N_8389,N_5941,N_3943);
nor U8390 (N_8390,N_3420,N_5881);
or U8391 (N_8391,N_2032,N_1131);
nor U8392 (N_8392,N_4617,N_1251);
nor U8393 (N_8393,N_4510,N_3894);
xor U8394 (N_8394,N_3858,N_4359);
or U8395 (N_8395,N_5124,N_5449);
or U8396 (N_8396,N_3481,N_47);
nand U8397 (N_8397,N_548,N_2890);
and U8398 (N_8398,N_2752,N_447);
nor U8399 (N_8399,N_2610,N_2457);
nor U8400 (N_8400,N_5434,N_5351);
nand U8401 (N_8401,N_4035,N_868);
or U8402 (N_8402,N_5019,N_999);
nor U8403 (N_8403,N_4006,N_5442);
nand U8404 (N_8404,N_4793,N_5742);
or U8405 (N_8405,N_1264,N_3820);
nor U8406 (N_8406,N_2823,N_1365);
nand U8407 (N_8407,N_3534,N_39);
nand U8408 (N_8408,N_2557,N_4895);
xor U8409 (N_8409,N_159,N_1186);
or U8410 (N_8410,N_3009,N_3841);
xnor U8411 (N_8411,N_2136,N_4589);
or U8412 (N_8412,N_63,N_5278);
nand U8413 (N_8413,N_4873,N_5249);
nor U8414 (N_8414,N_4350,N_3616);
nor U8415 (N_8415,N_3011,N_5473);
and U8416 (N_8416,N_5513,N_1555);
or U8417 (N_8417,N_2244,N_2164);
or U8418 (N_8418,N_2733,N_4248);
nand U8419 (N_8419,N_904,N_4528);
or U8420 (N_8420,N_4328,N_3855);
xnor U8421 (N_8421,N_3182,N_210);
nor U8422 (N_8422,N_3167,N_4445);
or U8423 (N_8423,N_5472,N_1327);
nor U8424 (N_8424,N_1519,N_3371);
xnor U8425 (N_8425,N_4352,N_368);
and U8426 (N_8426,N_4967,N_1537);
and U8427 (N_8427,N_930,N_648);
nor U8428 (N_8428,N_4457,N_5362);
nor U8429 (N_8429,N_3245,N_2077);
and U8430 (N_8430,N_1859,N_4266);
or U8431 (N_8431,N_2506,N_4339);
or U8432 (N_8432,N_1657,N_300);
nand U8433 (N_8433,N_3145,N_2206);
nand U8434 (N_8434,N_2397,N_54);
nor U8435 (N_8435,N_4477,N_2056);
nor U8436 (N_8436,N_1763,N_2234);
and U8437 (N_8437,N_5077,N_478);
nor U8438 (N_8438,N_1819,N_5642);
or U8439 (N_8439,N_698,N_2461);
nand U8440 (N_8440,N_5506,N_3520);
nor U8441 (N_8441,N_3485,N_872);
nand U8442 (N_8442,N_1792,N_1955);
nand U8443 (N_8443,N_5908,N_1988);
nor U8444 (N_8444,N_173,N_2883);
and U8445 (N_8445,N_2641,N_2076);
nand U8446 (N_8446,N_927,N_993);
or U8447 (N_8447,N_865,N_4344);
nor U8448 (N_8448,N_561,N_5195);
xor U8449 (N_8449,N_3501,N_1527);
nor U8450 (N_8450,N_1373,N_514);
xnor U8451 (N_8451,N_1672,N_3686);
xor U8452 (N_8452,N_1207,N_3594);
nand U8453 (N_8453,N_59,N_5685);
xnor U8454 (N_8454,N_1255,N_1141);
and U8455 (N_8455,N_2807,N_3754);
or U8456 (N_8456,N_3131,N_2061);
or U8457 (N_8457,N_2162,N_5363);
or U8458 (N_8458,N_2175,N_3471);
or U8459 (N_8459,N_3210,N_4832);
nor U8460 (N_8460,N_5025,N_5602);
and U8461 (N_8461,N_1318,N_1648);
xnor U8462 (N_8462,N_3973,N_2738);
nand U8463 (N_8463,N_3646,N_1209);
nand U8464 (N_8464,N_246,N_3847);
nor U8465 (N_8465,N_2791,N_4438);
and U8466 (N_8466,N_734,N_120);
nand U8467 (N_8467,N_4252,N_2908);
or U8468 (N_8468,N_5643,N_1535);
or U8469 (N_8469,N_124,N_4938);
and U8470 (N_8470,N_3948,N_883);
or U8471 (N_8471,N_1880,N_3608);
nor U8472 (N_8472,N_859,N_5253);
nand U8473 (N_8473,N_3039,N_261);
nand U8474 (N_8474,N_5109,N_2781);
and U8475 (N_8475,N_1817,N_3386);
or U8476 (N_8476,N_4075,N_5841);
xor U8477 (N_8477,N_1847,N_2559);
or U8478 (N_8478,N_2415,N_5768);
and U8479 (N_8479,N_3024,N_5055);
nand U8480 (N_8480,N_4305,N_1436);
nand U8481 (N_8481,N_153,N_1407);
nand U8482 (N_8482,N_4864,N_2456);
or U8483 (N_8483,N_4500,N_4076);
or U8484 (N_8484,N_5422,N_5255);
nor U8485 (N_8485,N_1319,N_5754);
or U8486 (N_8486,N_3999,N_2757);
and U8487 (N_8487,N_1338,N_398);
and U8488 (N_8488,N_4361,N_3233);
nand U8489 (N_8489,N_2190,N_1134);
or U8490 (N_8490,N_4752,N_4424);
or U8491 (N_8491,N_5832,N_3136);
nor U8492 (N_8492,N_560,N_2591);
or U8493 (N_8493,N_965,N_3052);
and U8494 (N_8494,N_2628,N_5679);
and U8495 (N_8495,N_1377,N_1586);
and U8496 (N_8496,N_4875,N_2947);
nor U8497 (N_8497,N_947,N_5447);
nand U8498 (N_8498,N_1944,N_3198);
nand U8499 (N_8499,N_3514,N_3282);
and U8500 (N_8500,N_4738,N_1638);
nand U8501 (N_8501,N_1930,N_5734);
nor U8502 (N_8502,N_3750,N_3978);
or U8503 (N_8503,N_3037,N_3521);
or U8504 (N_8504,N_5466,N_36);
or U8505 (N_8505,N_4527,N_949);
nand U8506 (N_8506,N_1161,N_345);
and U8507 (N_8507,N_3085,N_3328);
xor U8508 (N_8508,N_2505,N_4135);
nor U8509 (N_8509,N_5400,N_1841);
nor U8510 (N_8510,N_5210,N_1368);
xnor U8511 (N_8511,N_2656,N_51);
or U8512 (N_8512,N_1837,N_2092);
xnor U8513 (N_8513,N_4891,N_1659);
nor U8514 (N_8514,N_2613,N_5141);
nand U8515 (N_8515,N_5795,N_874);
nor U8516 (N_8516,N_5028,N_5982);
nor U8517 (N_8517,N_5189,N_761);
or U8518 (N_8518,N_3707,N_4753);
xnor U8519 (N_8519,N_3013,N_5615);
nand U8520 (N_8520,N_2255,N_5046);
or U8521 (N_8521,N_2581,N_80);
or U8522 (N_8522,N_3357,N_4766);
and U8523 (N_8523,N_4672,N_4441);
and U8524 (N_8524,N_1574,N_1949);
xnor U8525 (N_8525,N_1051,N_5677);
or U8526 (N_8526,N_2611,N_2783);
and U8527 (N_8527,N_691,N_3349);
nor U8528 (N_8528,N_5818,N_4378);
xor U8529 (N_8529,N_2324,N_3114);
xnor U8530 (N_8530,N_2433,N_4983);
nand U8531 (N_8531,N_2124,N_3756);
nor U8532 (N_8532,N_5393,N_1809);
or U8533 (N_8533,N_5717,N_5549);
nor U8534 (N_8534,N_4725,N_2829);
and U8535 (N_8535,N_194,N_1019);
and U8536 (N_8536,N_1271,N_2079);
xnor U8537 (N_8537,N_4504,N_3695);
and U8538 (N_8538,N_3798,N_189);
nand U8539 (N_8539,N_312,N_4910);
xnor U8540 (N_8540,N_2104,N_4598);
xnor U8541 (N_8541,N_828,N_3344);
xor U8542 (N_8542,N_5491,N_5550);
xor U8543 (N_8543,N_1023,N_68);
or U8544 (N_8544,N_5846,N_3153);
or U8545 (N_8545,N_2932,N_1133);
and U8546 (N_8546,N_4987,N_3451);
nand U8547 (N_8547,N_79,N_5040);
xnor U8548 (N_8548,N_348,N_986);
nor U8549 (N_8549,N_1557,N_89);
or U8550 (N_8550,N_2706,N_1813);
nor U8551 (N_8551,N_2353,N_293);
nand U8552 (N_8552,N_5703,N_5640);
and U8553 (N_8553,N_2684,N_2356);
xor U8554 (N_8554,N_4831,N_2634);
nand U8555 (N_8555,N_2648,N_775);
and U8556 (N_8556,N_5845,N_1082);
nor U8557 (N_8557,N_5986,N_4316);
nor U8558 (N_8558,N_4279,N_2176);
nand U8559 (N_8559,N_3468,N_2965);
or U8560 (N_8560,N_1963,N_428);
nor U8561 (N_8561,N_3543,N_5405);
or U8562 (N_8562,N_1185,N_3619);
xor U8563 (N_8563,N_2437,N_3631);
or U8564 (N_8564,N_3336,N_2007);
or U8565 (N_8565,N_5076,N_5569);
and U8566 (N_8566,N_5089,N_262);
and U8567 (N_8567,N_5880,N_3461);
nand U8568 (N_8568,N_4733,N_5732);
xor U8569 (N_8569,N_458,N_4918);
or U8570 (N_8570,N_204,N_4947);
nor U8571 (N_8571,N_711,N_378);
or U8572 (N_8572,N_164,N_5715);
nor U8573 (N_8573,N_5505,N_1801);
nand U8574 (N_8574,N_5948,N_1720);
or U8575 (N_8575,N_1276,N_2131);
xor U8576 (N_8576,N_4175,N_5516);
or U8577 (N_8577,N_319,N_4728);
nand U8578 (N_8578,N_4082,N_1694);
nor U8579 (N_8579,N_1106,N_1127);
nor U8580 (N_8580,N_3870,N_3685);
and U8581 (N_8581,N_620,N_4982);
or U8582 (N_8582,N_427,N_314);
nor U8583 (N_8583,N_5956,N_5966);
nor U8584 (N_8584,N_757,N_207);
nor U8585 (N_8585,N_4592,N_5374);
xor U8586 (N_8586,N_2455,N_5780);
or U8587 (N_8587,N_2220,N_2298);
and U8588 (N_8588,N_4007,N_3432);
xnor U8589 (N_8589,N_4487,N_4638);
or U8590 (N_8590,N_4782,N_776);
and U8591 (N_8591,N_4051,N_621);
and U8592 (N_8592,N_4554,N_4759);
or U8593 (N_8593,N_24,N_5290);
nand U8594 (N_8594,N_1107,N_1710);
and U8595 (N_8595,N_4697,N_3506);
nor U8596 (N_8596,N_4488,N_1478);
xor U8597 (N_8597,N_3984,N_4623);
or U8598 (N_8598,N_1145,N_3322);
or U8599 (N_8599,N_2401,N_369);
or U8600 (N_8600,N_4723,N_2243);
xor U8601 (N_8601,N_1862,N_1590);
or U8602 (N_8602,N_4569,N_5916);
nor U8603 (N_8603,N_4118,N_4632);
and U8604 (N_8604,N_1192,N_5148);
nor U8605 (N_8605,N_1565,N_2942);
and U8606 (N_8606,N_4142,N_2040);
xor U8607 (N_8607,N_397,N_5316);
nand U8608 (N_8608,N_5658,N_5078);
xor U8609 (N_8609,N_3408,N_4821);
nand U8610 (N_8610,N_1410,N_1198);
xor U8611 (N_8611,N_3397,N_390);
nand U8612 (N_8612,N_4935,N_4612);
or U8613 (N_8613,N_1065,N_5185);
xnor U8614 (N_8614,N_4645,N_4751);
or U8615 (N_8615,N_4811,N_4471);
nor U8616 (N_8616,N_1494,N_2766);
and U8617 (N_8617,N_5172,N_338);
or U8618 (N_8618,N_435,N_1742);
nor U8619 (N_8619,N_5438,N_3117);
xor U8620 (N_8620,N_1899,N_739);
xnor U8621 (N_8621,N_5541,N_5102);
nand U8622 (N_8622,N_2249,N_5250);
xor U8623 (N_8623,N_3718,N_4957);
and U8624 (N_8624,N_5791,N_5996);
nand U8625 (N_8625,N_4986,N_5334);
and U8626 (N_8626,N_5024,N_3655);
or U8627 (N_8627,N_4576,N_3715);
nand U8628 (N_8628,N_2474,N_5879);
nor U8629 (N_8629,N_2815,N_851);
or U8630 (N_8630,N_2166,N_5838);
or U8631 (N_8631,N_95,N_3067);
or U8632 (N_8632,N_537,N_1167);
nor U8633 (N_8633,N_2797,N_3806);
nor U8634 (N_8634,N_3147,N_5470);
xnor U8635 (N_8635,N_2018,N_848);
nor U8636 (N_8636,N_1849,N_4574);
nand U8637 (N_8637,N_4878,N_250);
nor U8638 (N_8638,N_1347,N_2970);
and U8639 (N_8639,N_444,N_664);
xnor U8640 (N_8640,N_2100,N_329);
and U8641 (N_8641,N_5543,N_347);
xor U8642 (N_8642,N_2541,N_5526);
xnor U8643 (N_8643,N_2608,N_4443);
and U8644 (N_8644,N_62,N_1117);
or U8645 (N_8645,N_5977,N_5970);
and U8646 (N_8646,N_2636,N_5218);
and U8647 (N_8647,N_4785,N_1058);
or U8648 (N_8648,N_5597,N_1035);
or U8649 (N_8649,N_3704,N_1609);
nand U8650 (N_8650,N_2725,N_4272);
or U8651 (N_8651,N_1959,N_1049);
nand U8652 (N_8652,N_2272,N_83);
or U8653 (N_8653,N_5456,N_2561);
xor U8654 (N_8654,N_3623,N_5445);
and U8655 (N_8655,N_2667,N_0);
and U8656 (N_8656,N_2765,N_2159);
nand U8657 (N_8657,N_3590,N_5433);
or U8658 (N_8658,N_3900,N_654);
nand U8659 (N_8659,N_5814,N_542);
xor U8660 (N_8660,N_2015,N_282);
or U8661 (N_8661,N_2375,N_1294);
or U8662 (N_8662,N_2517,N_2421);
nand U8663 (N_8663,N_3452,N_216);
nand U8664 (N_8664,N_2203,N_572);
nor U8665 (N_8665,N_4582,N_2717);
or U8666 (N_8666,N_900,N_1390);
nand U8667 (N_8667,N_3960,N_1119);
nor U8668 (N_8668,N_4073,N_232);
xnor U8669 (N_8669,N_147,N_257);
xor U8670 (N_8670,N_2238,N_5573);
nor U8671 (N_8671,N_472,N_4661);
nor U8672 (N_8672,N_1363,N_4255);
and U8673 (N_8673,N_5938,N_1000);
or U8674 (N_8674,N_4090,N_1791);
nand U8675 (N_8675,N_3837,N_3719);
or U8676 (N_8676,N_5298,N_2476);
xnor U8677 (N_8677,N_2796,N_5693);
or U8678 (N_8678,N_4540,N_1498);
or U8679 (N_8679,N_3552,N_5193);
or U8680 (N_8680,N_5836,N_4885);
xnor U8681 (N_8681,N_4102,N_3222);
nand U8682 (N_8682,N_4029,N_113);
nor U8683 (N_8683,N_1202,N_946);
nand U8684 (N_8684,N_5510,N_559);
or U8685 (N_8685,N_2404,N_2912);
and U8686 (N_8686,N_3684,N_2156);
nand U8687 (N_8687,N_5469,N_4365);
nand U8688 (N_8688,N_4334,N_5050);
or U8689 (N_8689,N_956,N_4882);
nand U8690 (N_8690,N_5910,N_2606);
nor U8691 (N_8691,N_633,N_4237);
or U8692 (N_8692,N_944,N_3035);
and U8693 (N_8693,N_2905,N_4939);
xor U8694 (N_8694,N_460,N_3048);
xor U8695 (N_8695,N_4068,N_294);
or U8696 (N_8696,N_1784,N_914);
or U8697 (N_8697,N_414,N_2235);
xnor U8698 (N_8698,N_3985,N_1908);
nand U8699 (N_8699,N_2282,N_4041);
nor U8700 (N_8700,N_3194,N_4859);
or U8701 (N_8701,N_4454,N_4409);
nand U8702 (N_8702,N_3342,N_5843);
or U8703 (N_8703,N_4150,N_4257);
nor U8704 (N_8704,N_4044,N_1190);
xnor U8705 (N_8705,N_441,N_1853);
nand U8706 (N_8706,N_46,N_2088);
nand U8707 (N_8707,N_5552,N_2179);
xnor U8708 (N_8708,N_4778,N_3547);
nor U8709 (N_8709,N_2876,N_1864);
nor U8710 (N_8710,N_165,N_1336);
nand U8711 (N_8711,N_3966,N_2779);
and U8712 (N_8712,N_705,N_2115);
or U8713 (N_8713,N_2936,N_551);
nand U8714 (N_8714,N_1304,N_777);
and U8715 (N_8715,N_1452,N_1661);
xnor U8716 (N_8716,N_58,N_2414);
nor U8717 (N_8717,N_3517,N_5731);
xor U8718 (N_8718,N_1962,N_5251);
nand U8719 (N_8719,N_2804,N_5702);
xnor U8720 (N_8720,N_3679,N_4985);
nand U8721 (N_8721,N_4581,N_2069);
and U8722 (N_8722,N_313,N_4415);
nand U8723 (N_8723,N_1126,N_2014);
nor U8724 (N_8724,N_3675,N_1433);
nor U8725 (N_8725,N_2848,N_2482);
nand U8726 (N_8726,N_2194,N_4205);
or U8727 (N_8727,N_3952,N_5058);
or U8728 (N_8728,N_2768,N_4836);
or U8729 (N_8729,N_1699,N_2822);
or U8730 (N_8730,N_5739,N_3747);
and U8731 (N_8731,N_4605,N_979);
or U8732 (N_8732,N_1514,N_471);
and U8733 (N_8733,N_4534,N_2521);
or U8734 (N_8734,N_683,N_5131);
and U8735 (N_8735,N_2739,N_3922);
nand U8736 (N_8736,N_2925,N_4599);
or U8737 (N_8737,N_3665,N_251);
nand U8738 (N_8738,N_455,N_4696);
nor U8739 (N_8739,N_3821,N_2836);
and U8740 (N_8740,N_631,N_3946);
or U8741 (N_8741,N_2934,N_3062);
nand U8742 (N_8742,N_840,N_5216);
nor U8743 (N_8743,N_610,N_4278);
or U8744 (N_8744,N_2926,N_3352);
nor U8745 (N_8745,N_3926,N_2347);
or U8746 (N_8746,N_5945,N_3786);
or U8747 (N_8747,N_4087,N_5476);
and U8748 (N_8748,N_1520,N_4841);
nand U8749 (N_8749,N_5454,N_4886);
xor U8750 (N_8750,N_4430,N_64);
and U8751 (N_8751,N_2117,N_3418);
nand U8752 (N_8752,N_5002,N_5202);
or U8753 (N_8753,N_5437,N_2582);
xor U8754 (N_8754,N_3020,N_1354);
and U8755 (N_8755,N_3444,N_1163);
xor U8756 (N_8756,N_3027,N_4019);
and U8757 (N_8757,N_5380,N_1972);
xnor U8758 (N_8758,N_713,N_527);
and U8759 (N_8759,N_2146,N_4690);
and U8760 (N_8760,N_515,N_4133);
xor U8761 (N_8761,N_2794,N_495);
nor U8762 (N_8762,N_267,N_1902);
or U8763 (N_8763,N_1144,N_522);
nand U8764 (N_8764,N_2550,N_5214);
xnor U8765 (N_8765,N_788,N_1653);
and U8766 (N_8766,N_636,N_5532);
nand U8767 (N_8767,N_4925,N_4163);
nand U8768 (N_8768,N_3248,N_96);
nor U8769 (N_8769,N_2237,N_3467);
nand U8770 (N_8770,N_5670,N_4667);
xnor U8771 (N_8771,N_4596,N_3617);
xnor U8772 (N_8772,N_2549,N_4674);
nor U8773 (N_8773,N_1644,N_2909);
and U8774 (N_8774,N_4108,N_5386);
xnor U8775 (N_8775,N_5031,N_4999);
nor U8776 (N_8776,N_3720,N_1807);
xnor U8777 (N_8777,N_4081,N_4407);
or U8778 (N_8778,N_5016,N_4673);
nor U8779 (N_8779,N_597,N_4079);
and U8780 (N_8780,N_3857,N_3827);
xor U8781 (N_8781,N_5111,N_5844);
nand U8782 (N_8782,N_3692,N_3343);
or U8783 (N_8783,N_3769,N_652);
nand U8784 (N_8784,N_86,N_3490);
xnor U8785 (N_8785,N_4813,N_3473);
nand U8786 (N_8786,N_4496,N_393);
or U8787 (N_8787,N_406,N_3834);
or U8788 (N_8788,N_4434,N_1032);
nand U8789 (N_8789,N_4195,N_3296);
nor U8790 (N_8790,N_5965,N_4698);
and U8791 (N_8791,N_2438,N_3536);
xnor U8792 (N_8792,N_4708,N_4270);
xnor U8793 (N_8793,N_5126,N_1604);
or U8794 (N_8794,N_403,N_142);
xnor U8795 (N_8795,N_1926,N_4492);
and U8796 (N_8796,N_5895,N_4858);
and U8797 (N_8797,N_544,N_4355);
and U8798 (N_8798,N_2395,N_1323);
xnor U8799 (N_8799,N_4362,N_3443);
nor U8800 (N_8800,N_154,N_4578);
nand U8801 (N_8801,N_5928,N_2871);
and U8802 (N_8802,N_5230,N_3990);
nor U8803 (N_8803,N_2227,N_2420);
and U8804 (N_8804,N_4523,N_4852);
nor U8805 (N_8805,N_1441,N_2024);
xor U8806 (N_8806,N_5633,N_5842);
nand U8807 (N_8807,N_4953,N_2085);
nand U8808 (N_8808,N_2654,N_5320);
and U8809 (N_8809,N_1913,N_2133);
or U8810 (N_8810,N_4480,N_4536);
nor U8811 (N_8811,N_5121,N_1455);
and U8812 (N_8812,N_4607,N_5802);
nand U8813 (N_8813,N_3830,N_3883);
nor U8814 (N_8814,N_182,N_5375);
xnor U8815 (N_8815,N_3953,N_1288);
or U8816 (N_8816,N_3760,N_4893);
nand U8817 (N_8817,N_3012,N_440);
nor U8818 (N_8818,N_5032,N_3376);
nand U8819 (N_8819,N_2742,N_283);
nor U8820 (N_8820,N_1178,N_301);
xor U8821 (N_8821,N_5927,N_1903);
nand U8822 (N_8822,N_2664,N_4806);
and U8823 (N_8823,N_4964,N_5008);
xnor U8824 (N_8824,N_259,N_1723);
xor U8825 (N_8825,N_416,N_3555);
xor U8826 (N_8826,N_5421,N_4700);
nor U8827 (N_8827,N_613,N_4166);
nand U8828 (N_8828,N_4121,N_1536);
nand U8829 (N_8829,N_2653,N_659);
xnor U8830 (N_8830,N_3941,N_1197);
nand U8831 (N_8831,N_507,N_936);
and U8832 (N_8832,N_4260,N_3337);
and U8833 (N_8833,N_5872,N_5052);
nand U8834 (N_8834,N_385,N_2129);
and U8835 (N_8835,N_2054,N_404);
nor U8836 (N_8836,N_670,N_4353);
and U8837 (N_8837,N_4802,N_5924);
and U8838 (N_8838,N_3119,N_5787);
or U8839 (N_8839,N_2842,N_2219);
nand U8840 (N_8840,N_1469,N_1138);
and U8841 (N_8841,N_3174,N_1597);
or U8842 (N_8842,N_3863,N_1726);
or U8843 (N_8843,N_1670,N_3047);
nand U8844 (N_8844,N_4743,N_1406);
xor U8845 (N_8845,N_4026,N_3598);
xor U8846 (N_8846,N_3882,N_4533);
nand U8847 (N_8847,N_1067,N_4892);
and U8848 (N_8848,N_5598,N_1199);
nand U8849 (N_8849,N_67,N_3928);
xnor U8850 (N_8850,N_5720,N_4080);
nand U8851 (N_8851,N_40,N_5012);
and U8852 (N_8852,N_3478,N_3235);
xor U8853 (N_8853,N_5062,N_5143);
and U8854 (N_8854,N_531,N_5737);
or U8855 (N_8855,N_420,N_358);
nor U8856 (N_8856,N_3350,N_1739);
xnor U8857 (N_8857,N_3441,N_4078);
or U8858 (N_8858,N_5142,N_1121);
nor U8859 (N_8859,N_1713,N_2532);
nand U8860 (N_8860,N_2755,N_93);
nand U8861 (N_8861,N_1396,N_3570);
nand U8862 (N_8862,N_4058,N_4225);
or U8863 (N_8863,N_2008,N_2491);
nor U8864 (N_8864,N_3647,N_5889);
nor U8865 (N_8865,N_5204,N_3244);
nor U8866 (N_8866,N_2994,N_4433);
and U8867 (N_8867,N_2384,N_1152);
nand U8868 (N_8868,N_3772,N_3743);
nor U8869 (N_8869,N_2728,N_2843);
and U8870 (N_8870,N_2711,N_4072);
or U8871 (N_8871,N_2458,N_4746);
or U8872 (N_8872,N_1226,N_3226);
and U8873 (N_8873,N_5704,N_190);
and U8874 (N_8874,N_1224,N_1811);
xor U8875 (N_8875,N_2388,N_5891);
xnor U8876 (N_8876,N_5212,N_5827);
and U8877 (N_8877,N_2019,N_2841);
nor U8878 (N_8878,N_5873,N_5067);
nor U8879 (N_8879,N_605,N_5242);
xnor U8880 (N_8880,N_3170,N_1009);
or U8881 (N_8881,N_3587,N_1210);
xor U8882 (N_8882,N_5764,N_1059);
or U8883 (N_8883,N_5655,N_5547);
nor U8884 (N_8884,N_1603,N_3464);
nor U8885 (N_8885,N_686,N_130);
and U8886 (N_8886,N_4779,N_525);
nand U8887 (N_8887,N_571,N_806);
nor U8888 (N_8888,N_174,N_2278);
xnor U8889 (N_8889,N_4681,N_5859);
nor U8890 (N_8890,N_622,N_5414);
nor U8891 (N_8891,N_1497,N_2626);
nand U8892 (N_8892,N_3356,N_4122);
nand U8893 (N_8893,N_2236,N_5138);
or U8894 (N_8894,N_4229,N_2047);
xor U8895 (N_8895,N_3250,N_2189);
xnor U8896 (N_8896,N_891,N_4898);
and U8897 (N_8897,N_1910,N_330);
xnor U8898 (N_8898,N_31,N_736);
nand U8899 (N_8899,N_5183,N_2691);
or U8900 (N_8900,N_4816,N_5304);
nor U8901 (N_8901,N_1331,N_2480);
xnor U8902 (N_8902,N_44,N_574);
xor U8903 (N_8903,N_2743,N_2987);
xnor U8904 (N_8904,N_2185,N_529);
xor U8905 (N_8905,N_2998,N_5675);
and U8906 (N_8906,N_5098,N_5246);
nor U8907 (N_8907,N_1836,N_5166);
and U8908 (N_8908,N_3059,N_1681);
xnor U8909 (N_8909,N_3572,N_5122);
nand U8910 (N_8910,N_4710,N_2082);
or U8911 (N_8911,N_5241,N_1097);
or U8912 (N_8912,N_1215,N_1042);
xor U8913 (N_8913,N_4167,N_1101);
nor U8914 (N_8914,N_4757,N_785);
or U8915 (N_8915,N_3763,N_1130);
xnor U8916 (N_8916,N_26,N_5482);
nand U8917 (N_8917,N_1966,N_2102);
or U8918 (N_8918,N_4542,N_2161);
xnor U8919 (N_8919,N_3092,N_5232);
nand U8920 (N_8920,N_5481,N_694);
or U8921 (N_8921,N_3537,N_2682);
nand U8922 (N_8922,N_731,N_3107);
nand U8923 (N_8923,N_5564,N_5718);
and U8924 (N_8924,N_2184,N_3126);
nor U8925 (N_8925,N_5592,N_5135);
or U8926 (N_8926,N_4716,N_866);
nor U8927 (N_8927,N_4211,N_2975);
or U8928 (N_8928,N_2633,N_4405);
nand U8929 (N_8929,N_4955,N_3484);
nor U8930 (N_8930,N_3404,N_2901);
or U8931 (N_8931,N_260,N_104);
xor U8932 (N_8932,N_5271,N_3495);
xnor U8933 (N_8933,N_5816,N_1640);
or U8934 (N_8934,N_2486,N_1800);
xor U8935 (N_8935,N_1235,N_2341);
xor U8936 (N_8936,N_135,N_439);
and U8937 (N_8937,N_4172,N_192);
nor U8938 (N_8938,N_498,N_5403);
and U8939 (N_8939,N_4165,N_2824);
nand U8940 (N_8940,N_2045,N_2900);
nor U8941 (N_8941,N_983,N_1906);
xnor U8942 (N_8942,N_3192,N_21);
and U8943 (N_8943,N_4899,N_1113);
nor U8944 (N_8944,N_1743,N_2850);
and U8945 (N_8945,N_5546,N_4658);
or U8946 (N_8946,N_1883,N_2593);
nor U8947 (N_8947,N_3102,N_3440);
and U8948 (N_8948,N_2575,N_4742);
nor U8949 (N_8949,N_1168,N_5621);
nand U8950 (N_8950,N_4881,N_2406);
nor U8951 (N_8951,N_2152,N_1180);
nor U8952 (N_8952,N_1856,N_599);
nand U8953 (N_8953,N_573,N_1684);
nand U8954 (N_8954,N_211,N_3487);
nor U8955 (N_8955,N_5207,N_1563);
and U8956 (N_8956,N_2362,N_2109);
nor U8957 (N_8957,N_3518,N_2495);
or U8958 (N_8958,N_4417,N_1482);
and U8959 (N_8959,N_4331,N_2588);
and U8960 (N_8960,N_3896,N_3801);
xor U8961 (N_8961,N_1632,N_160);
and U8962 (N_8962,N_3620,N_4990);
and U8963 (N_8963,N_3709,N_4546);
nor U8964 (N_8964,N_2091,N_4486);
xor U8965 (N_8965,N_1091,N_3449);
and U8966 (N_8966,N_4145,N_833);
nor U8967 (N_8967,N_5332,N_2718);
xnor U8968 (N_8968,N_499,N_3705);
xor U8969 (N_8969,N_2427,N_5686);
or U8970 (N_8970,N_4960,N_1866);
or U8971 (N_8971,N_5344,N_4318);
xor U8972 (N_8972,N_4459,N_4808);
or U8973 (N_8973,N_4382,N_2242);
nor U8974 (N_8974,N_5890,N_4164);
xor U8975 (N_8975,N_3191,N_4791);
and U8976 (N_8976,N_4380,N_3385);
nand U8977 (N_8977,N_2254,N_746);
xnor U8978 (N_8978,N_2105,N_1560);
or U8979 (N_8979,N_4530,N_4863);
nor U8980 (N_8980,N_4787,N_3036);
xnor U8981 (N_8981,N_4877,N_1409);
nor U8982 (N_8982,N_3380,N_2502);
xor U8983 (N_8983,N_5187,N_3030);
or U8984 (N_8984,N_342,N_2630);
nor U8985 (N_8985,N_2997,N_1205);
xnor U8986 (N_8986,N_506,N_5341);
or U8987 (N_8987,N_5940,N_4744);
nand U8988 (N_8988,N_452,N_1627);
nor U8989 (N_8989,N_4943,N_2918);
and U8990 (N_8990,N_3227,N_5455);
xnor U8991 (N_8991,N_1311,N_3677);
or U8992 (N_8992,N_5115,N_3284);
or U8993 (N_8993,N_3066,N_2259);
nand U8994 (N_8994,N_2096,N_2772);
and U8995 (N_8995,N_4647,N_4194);
and U8996 (N_8996,N_4502,N_2065);
nand U8997 (N_8997,N_1540,N_3442);
xor U8998 (N_8998,N_2407,N_1060);
nor U8999 (N_8999,N_1588,N_4760);
nand U9000 (N_9000,N_44,N_4513);
or U9001 (N_9001,N_2911,N_2866);
nor U9002 (N_9002,N_4092,N_5468);
xor U9003 (N_9003,N_2522,N_73);
nor U9004 (N_9004,N_1043,N_3448);
and U9005 (N_9005,N_5695,N_4597);
nand U9006 (N_9006,N_2711,N_1218);
or U9007 (N_9007,N_5268,N_1629);
nand U9008 (N_9008,N_3374,N_5027);
xor U9009 (N_9009,N_752,N_4569);
xnor U9010 (N_9010,N_2247,N_5285);
and U9011 (N_9011,N_334,N_5592);
nor U9012 (N_9012,N_5899,N_400);
or U9013 (N_9013,N_1254,N_3173);
xor U9014 (N_9014,N_1879,N_1064);
xnor U9015 (N_9015,N_1813,N_4312);
nand U9016 (N_9016,N_2420,N_2624);
nor U9017 (N_9017,N_3976,N_3305);
or U9018 (N_9018,N_2687,N_3049);
xnor U9019 (N_9019,N_2744,N_1379);
and U9020 (N_9020,N_867,N_2073);
nand U9021 (N_9021,N_4918,N_2701);
xnor U9022 (N_9022,N_2643,N_5195);
nand U9023 (N_9023,N_2490,N_1658);
nor U9024 (N_9024,N_5938,N_3790);
nand U9025 (N_9025,N_2452,N_4960);
nor U9026 (N_9026,N_4724,N_319);
nor U9027 (N_9027,N_4012,N_3958);
nand U9028 (N_9028,N_4234,N_83);
nor U9029 (N_9029,N_4808,N_889);
or U9030 (N_9030,N_5525,N_1719);
nor U9031 (N_9031,N_354,N_3104);
nor U9032 (N_9032,N_1974,N_5814);
nand U9033 (N_9033,N_5905,N_2167);
nand U9034 (N_9034,N_250,N_4822);
or U9035 (N_9035,N_2024,N_3593);
nand U9036 (N_9036,N_2964,N_3327);
nor U9037 (N_9037,N_4646,N_3839);
xnor U9038 (N_9038,N_203,N_5382);
nor U9039 (N_9039,N_1248,N_4311);
or U9040 (N_9040,N_4748,N_4345);
nor U9041 (N_9041,N_617,N_4885);
xor U9042 (N_9042,N_2440,N_2652);
or U9043 (N_9043,N_2448,N_2721);
nand U9044 (N_9044,N_2579,N_5700);
nor U9045 (N_9045,N_3109,N_5538);
and U9046 (N_9046,N_4725,N_2951);
xor U9047 (N_9047,N_1238,N_2471);
and U9048 (N_9048,N_3650,N_2884);
nand U9049 (N_9049,N_1704,N_537);
nand U9050 (N_9050,N_408,N_1377);
xor U9051 (N_9051,N_1227,N_1130);
and U9052 (N_9052,N_2661,N_3413);
nor U9053 (N_9053,N_5673,N_285);
xor U9054 (N_9054,N_3965,N_2558);
nand U9055 (N_9055,N_1847,N_1142);
nor U9056 (N_9056,N_4235,N_2763);
and U9057 (N_9057,N_679,N_543);
and U9058 (N_9058,N_3664,N_4864);
nand U9059 (N_9059,N_296,N_462);
xnor U9060 (N_9060,N_4770,N_3307);
and U9061 (N_9061,N_3111,N_1561);
nand U9062 (N_9062,N_2719,N_3144);
and U9063 (N_9063,N_4105,N_5402);
nand U9064 (N_9064,N_2548,N_2588);
nor U9065 (N_9065,N_4901,N_3353);
or U9066 (N_9066,N_3541,N_3504);
xor U9067 (N_9067,N_1542,N_5528);
nand U9068 (N_9068,N_1724,N_990);
xor U9069 (N_9069,N_3439,N_2108);
xnor U9070 (N_9070,N_2753,N_211);
nor U9071 (N_9071,N_2096,N_3669);
nor U9072 (N_9072,N_4801,N_1922);
xnor U9073 (N_9073,N_316,N_467);
nor U9074 (N_9074,N_4072,N_4728);
nor U9075 (N_9075,N_4496,N_3184);
nor U9076 (N_9076,N_1366,N_2446);
or U9077 (N_9077,N_544,N_2828);
or U9078 (N_9078,N_2561,N_5903);
nor U9079 (N_9079,N_3800,N_418);
nor U9080 (N_9080,N_1736,N_3073);
xor U9081 (N_9081,N_5001,N_4009);
nor U9082 (N_9082,N_1799,N_3854);
or U9083 (N_9083,N_4240,N_3045);
nand U9084 (N_9084,N_2264,N_4173);
or U9085 (N_9085,N_1499,N_4023);
and U9086 (N_9086,N_1860,N_417);
or U9087 (N_9087,N_5135,N_5193);
nor U9088 (N_9088,N_2658,N_1163);
nor U9089 (N_9089,N_4440,N_1478);
or U9090 (N_9090,N_3066,N_1766);
and U9091 (N_9091,N_1737,N_5014);
xnor U9092 (N_9092,N_2775,N_36);
nor U9093 (N_9093,N_2037,N_107);
nand U9094 (N_9094,N_2480,N_2731);
xor U9095 (N_9095,N_5839,N_4258);
xor U9096 (N_9096,N_4447,N_1645);
nor U9097 (N_9097,N_5583,N_4038);
nor U9098 (N_9098,N_5817,N_5919);
xor U9099 (N_9099,N_4062,N_4789);
nor U9100 (N_9100,N_1345,N_3434);
nor U9101 (N_9101,N_2853,N_528);
or U9102 (N_9102,N_5655,N_2129);
or U9103 (N_9103,N_5950,N_2916);
xnor U9104 (N_9104,N_4468,N_1028);
nor U9105 (N_9105,N_4970,N_2687);
nand U9106 (N_9106,N_743,N_4377);
or U9107 (N_9107,N_4206,N_2487);
nor U9108 (N_9108,N_2060,N_5156);
and U9109 (N_9109,N_1284,N_5473);
nand U9110 (N_9110,N_5237,N_4829);
xor U9111 (N_9111,N_1186,N_5655);
or U9112 (N_9112,N_154,N_5682);
or U9113 (N_9113,N_590,N_3843);
or U9114 (N_9114,N_1745,N_1921);
nor U9115 (N_9115,N_2269,N_269);
nand U9116 (N_9116,N_4144,N_703);
nor U9117 (N_9117,N_4253,N_3623);
nand U9118 (N_9118,N_2914,N_5941);
nor U9119 (N_9119,N_1031,N_2072);
or U9120 (N_9120,N_4549,N_1539);
xor U9121 (N_9121,N_1624,N_749);
nor U9122 (N_9122,N_5178,N_487);
and U9123 (N_9123,N_4056,N_697);
nor U9124 (N_9124,N_3800,N_3190);
xnor U9125 (N_9125,N_2549,N_4198);
and U9126 (N_9126,N_2894,N_751);
and U9127 (N_9127,N_2442,N_193);
xnor U9128 (N_9128,N_974,N_5315);
nand U9129 (N_9129,N_1198,N_2049);
and U9130 (N_9130,N_2015,N_4746);
nand U9131 (N_9131,N_4746,N_592);
nand U9132 (N_9132,N_4716,N_3974);
nor U9133 (N_9133,N_1601,N_264);
and U9134 (N_9134,N_2992,N_4625);
nor U9135 (N_9135,N_1481,N_158);
xor U9136 (N_9136,N_803,N_1057);
nand U9137 (N_9137,N_3278,N_2855);
nor U9138 (N_9138,N_3179,N_455);
xnor U9139 (N_9139,N_3119,N_1183);
or U9140 (N_9140,N_1553,N_5709);
xnor U9141 (N_9141,N_755,N_3861);
nor U9142 (N_9142,N_2588,N_1534);
xnor U9143 (N_9143,N_3061,N_3997);
nand U9144 (N_9144,N_170,N_4104);
nor U9145 (N_9145,N_3624,N_3922);
nand U9146 (N_9146,N_4727,N_787);
nor U9147 (N_9147,N_3091,N_3967);
nor U9148 (N_9148,N_1716,N_4873);
xor U9149 (N_9149,N_2838,N_1929);
xnor U9150 (N_9150,N_3363,N_4155);
xor U9151 (N_9151,N_3201,N_1382);
nor U9152 (N_9152,N_3591,N_4259);
or U9153 (N_9153,N_3612,N_1062);
and U9154 (N_9154,N_4655,N_803);
and U9155 (N_9155,N_784,N_5451);
or U9156 (N_9156,N_2896,N_3612);
nor U9157 (N_9157,N_558,N_488);
or U9158 (N_9158,N_241,N_1402);
or U9159 (N_9159,N_1640,N_3172);
nor U9160 (N_9160,N_3930,N_4868);
xor U9161 (N_9161,N_3388,N_1504);
nor U9162 (N_9162,N_3537,N_2647);
xor U9163 (N_9163,N_4638,N_658);
or U9164 (N_9164,N_2631,N_5179);
and U9165 (N_9165,N_1602,N_575);
or U9166 (N_9166,N_35,N_3130);
or U9167 (N_9167,N_3599,N_2612);
nor U9168 (N_9168,N_3838,N_5911);
or U9169 (N_9169,N_4297,N_255);
nand U9170 (N_9170,N_2095,N_2760);
and U9171 (N_9171,N_698,N_2762);
nand U9172 (N_9172,N_5140,N_3642);
or U9173 (N_9173,N_1903,N_413);
nor U9174 (N_9174,N_5788,N_5096);
and U9175 (N_9175,N_5647,N_5172);
nand U9176 (N_9176,N_3221,N_296);
and U9177 (N_9177,N_4176,N_3728);
nand U9178 (N_9178,N_2751,N_5310);
nand U9179 (N_9179,N_2207,N_2111);
nand U9180 (N_9180,N_4157,N_720);
xor U9181 (N_9181,N_995,N_5611);
or U9182 (N_9182,N_3602,N_4195);
and U9183 (N_9183,N_5467,N_4305);
or U9184 (N_9184,N_2202,N_4881);
and U9185 (N_9185,N_5910,N_5552);
or U9186 (N_9186,N_143,N_5181);
and U9187 (N_9187,N_4703,N_5396);
xnor U9188 (N_9188,N_3827,N_2664);
or U9189 (N_9189,N_2980,N_2664);
or U9190 (N_9190,N_5785,N_5026);
and U9191 (N_9191,N_2655,N_2642);
nor U9192 (N_9192,N_5054,N_3536);
nand U9193 (N_9193,N_4526,N_2132);
and U9194 (N_9194,N_4836,N_2855);
xor U9195 (N_9195,N_5055,N_1971);
or U9196 (N_9196,N_2175,N_4057);
and U9197 (N_9197,N_2467,N_3476);
nor U9198 (N_9198,N_859,N_5189);
xor U9199 (N_9199,N_276,N_2001);
and U9200 (N_9200,N_5914,N_1094);
nand U9201 (N_9201,N_29,N_3412);
nor U9202 (N_9202,N_5876,N_4117);
nand U9203 (N_9203,N_5087,N_5562);
xor U9204 (N_9204,N_4598,N_3113);
nand U9205 (N_9205,N_1779,N_848);
and U9206 (N_9206,N_2719,N_2000);
nor U9207 (N_9207,N_5729,N_1294);
xnor U9208 (N_9208,N_85,N_2538);
xor U9209 (N_9209,N_4177,N_934);
or U9210 (N_9210,N_5835,N_2242);
xnor U9211 (N_9211,N_4810,N_151);
nand U9212 (N_9212,N_1477,N_826);
and U9213 (N_9213,N_2692,N_5979);
xnor U9214 (N_9214,N_5809,N_3879);
or U9215 (N_9215,N_1158,N_467);
and U9216 (N_9216,N_5415,N_5379);
xnor U9217 (N_9217,N_4782,N_811);
and U9218 (N_9218,N_366,N_89);
nor U9219 (N_9219,N_1078,N_4107);
or U9220 (N_9220,N_4087,N_1403);
or U9221 (N_9221,N_4027,N_5066);
nor U9222 (N_9222,N_1418,N_4813);
xor U9223 (N_9223,N_931,N_3458);
or U9224 (N_9224,N_5690,N_3060);
xor U9225 (N_9225,N_1005,N_1433);
nor U9226 (N_9226,N_5894,N_1067);
nor U9227 (N_9227,N_1051,N_3448);
nand U9228 (N_9228,N_1083,N_1978);
xor U9229 (N_9229,N_1540,N_2171);
or U9230 (N_9230,N_3092,N_3494);
nand U9231 (N_9231,N_2650,N_5570);
nand U9232 (N_9232,N_2457,N_4307);
nand U9233 (N_9233,N_2492,N_1386);
nand U9234 (N_9234,N_3633,N_4557);
and U9235 (N_9235,N_2751,N_4285);
nand U9236 (N_9236,N_982,N_3760);
or U9237 (N_9237,N_1578,N_3077);
nor U9238 (N_9238,N_918,N_5135);
and U9239 (N_9239,N_811,N_3743);
nand U9240 (N_9240,N_1967,N_1289);
nor U9241 (N_9241,N_717,N_5358);
and U9242 (N_9242,N_3075,N_609);
nor U9243 (N_9243,N_2218,N_2327);
nor U9244 (N_9244,N_1251,N_2554);
and U9245 (N_9245,N_351,N_1758);
and U9246 (N_9246,N_3967,N_1313);
xor U9247 (N_9247,N_5095,N_5776);
xor U9248 (N_9248,N_5963,N_1978);
nor U9249 (N_9249,N_3589,N_4388);
and U9250 (N_9250,N_547,N_861);
nor U9251 (N_9251,N_2790,N_3040);
nor U9252 (N_9252,N_4999,N_1448);
nor U9253 (N_9253,N_2211,N_1464);
and U9254 (N_9254,N_1919,N_5144);
nor U9255 (N_9255,N_2230,N_5711);
nand U9256 (N_9256,N_5300,N_2149);
xnor U9257 (N_9257,N_1853,N_3922);
nor U9258 (N_9258,N_3783,N_3140);
and U9259 (N_9259,N_2887,N_4170);
nand U9260 (N_9260,N_4886,N_3338);
nor U9261 (N_9261,N_5708,N_4855);
and U9262 (N_9262,N_3587,N_3602);
nand U9263 (N_9263,N_3415,N_196);
nand U9264 (N_9264,N_1145,N_149);
nor U9265 (N_9265,N_3152,N_5835);
nand U9266 (N_9266,N_3826,N_5397);
or U9267 (N_9267,N_4392,N_2650);
nor U9268 (N_9268,N_4424,N_4288);
xnor U9269 (N_9269,N_282,N_1174);
and U9270 (N_9270,N_2590,N_170);
nand U9271 (N_9271,N_1658,N_4882);
or U9272 (N_9272,N_2983,N_2984);
or U9273 (N_9273,N_5197,N_2431);
and U9274 (N_9274,N_5570,N_670);
or U9275 (N_9275,N_1490,N_2184);
or U9276 (N_9276,N_1271,N_4485);
or U9277 (N_9277,N_2492,N_4653);
and U9278 (N_9278,N_5139,N_4360);
or U9279 (N_9279,N_3991,N_4551);
and U9280 (N_9280,N_3584,N_586);
and U9281 (N_9281,N_5510,N_2254);
or U9282 (N_9282,N_1179,N_691);
or U9283 (N_9283,N_4862,N_703);
and U9284 (N_9284,N_3774,N_812);
nor U9285 (N_9285,N_3197,N_4945);
nand U9286 (N_9286,N_4832,N_1986);
and U9287 (N_9287,N_5389,N_1155);
nor U9288 (N_9288,N_2776,N_2596);
or U9289 (N_9289,N_1681,N_4281);
nand U9290 (N_9290,N_340,N_3167);
nor U9291 (N_9291,N_3923,N_444);
xor U9292 (N_9292,N_240,N_2803);
xnor U9293 (N_9293,N_4135,N_4198);
or U9294 (N_9294,N_1981,N_3220);
nand U9295 (N_9295,N_3538,N_3708);
xnor U9296 (N_9296,N_1230,N_4610);
and U9297 (N_9297,N_5588,N_5930);
or U9298 (N_9298,N_465,N_4120);
and U9299 (N_9299,N_1102,N_1987);
xor U9300 (N_9300,N_5283,N_3207);
nor U9301 (N_9301,N_664,N_1045);
nor U9302 (N_9302,N_3496,N_1444);
nand U9303 (N_9303,N_4313,N_1502);
xnor U9304 (N_9304,N_4288,N_2254);
xor U9305 (N_9305,N_5586,N_4186);
or U9306 (N_9306,N_2777,N_3625);
and U9307 (N_9307,N_2301,N_3800);
nor U9308 (N_9308,N_2101,N_4696);
nor U9309 (N_9309,N_4341,N_2855);
xor U9310 (N_9310,N_2207,N_4931);
nand U9311 (N_9311,N_1687,N_2305);
nand U9312 (N_9312,N_5727,N_2664);
nand U9313 (N_9313,N_1714,N_329);
nand U9314 (N_9314,N_5691,N_227);
nor U9315 (N_9315,N_1238,N_1456);
and U9316 (N_9316,N_2035,N_3737);
xor U9317 (N_9317,N_1233,N_966);
xnor U9318 (N_9318,N_1925,N_5477);
and U9319 (N_9319,N_3279,N_4160);
and U9320 (N_9320,N_1439,N_2292);
xor U9321 (N_9321,N_4253,N_3612);
and U9322 (N_9322,N_3063,N_3851);
xor U9323 (N_9323,N_4052,N_2086);
and U9324 (N_9324,N_5339,N_5637);
or U9325 (N_9325,N_3662,N_5951);
xnor U9326 (N_9326,N_737,N_2230);
or U9327 (N_9327,N_1534,N_5355);
nor U9328 (N_9328,N_5014,N_2500);
xor U9329 (N_9329,N_3856,N_2090);
nor U9330 (N_9330,N_3460,N_1018);
nand U9331 (N_9331,N_2334,N_2884);
or U9332 (N_9332,N_1390,N_2461);
nor U9333 (N_9333,N_1504,N_9);
xor U9334 (N_9334,N_4374,N_2656);
or U9335 (N_9335,N_2685,N_79);
xor U9336 (N_9336,N_4106,N_5409);
nand U9337 (N_9337,N_1501,N_1231);
and U9338 (N_9338,N_2777,N_4659);
xor U9339 (N_9339,N_3162,N_1277);
and U9340 (N_9340,N_3444,N_2457);
nand U9341 (N_9341,N_1185,N_2226);
or U9342 (N_9342,N_1986,N_3810);
and U9343 (N_9343,N_2998,N_5395);
and U9344 (N_9344,N_5076,N_4963);
and U9345 (N_9345,N_4879,N_5902);
nor U9346 (N_9346,N_776,N_3176);
xnor U9347 (N_9347,N_5834,N_3392);
nand U9348 (N_9348,N_1531,N_5226);
or U9349 (N_9349,N_2417,N_4906);
nand U9350 (N_9350,N_3422,N_212);
and U9351 (N_9351,N_4266,N_5111);
nor U9352 (N_9352,N_5825,N_3097);
xor U9353 (N_9353,N_5445,N_121);
xor U9354 (N_9354,N_5416,N_4516);
nand U9355 (N_9355,N_3284,N_489);
and U9356 (N_9356,N_2965,N_1313);
xor U9357 (N_9357,N_767,N_1733);
xnor U9358 (N_9358,N_4549,N_4293);
nor U9359 (N_9359,N_3765,N_4488);
xnor U9360 (N_9360,N_4639,N_1426);
nand U9361 (N_9361,N_589,N_4593);
xor U9362 (N_9362,N_5659,N_1998);
nor U9363 (N_9363,N_683,N_1940);
nor U9364 (N_9364,N_4748,N_2855);
nand U9365 (N_9365,N_5607,N_424);
nand U9366 (N_9366,N_3709,N_1694);
nor U9367 (N_9367,N_1587,N_4941);
and U9368 (N_9368,N_4282,N_5233);
or U9369 (N_9369,N_5006,N_4977);
xnor U9370 (N_9370,N_5090,N_1606);
or U9371 (N_9371,N_5869,N_1366);
and U9372 (N_9372,N_3683,N_1762);
or U9373 (N_9373,N_3597,N_4425);
and U9374 (N_9374,N_4817,N_532);
and U9375 (N_9375,N_5090,N_2107);
xnor U9376 (N_9376,N_3713,N_171);
and U9377 (N_9377,N_4409,N_5571);
xor U9378 (N_9378,N_4224,N_5129);
xor U9379 (N_9379,N_4093,N_3250);
nand U9380 (N_9380,N_1737,N_4974);
nor U9381 (N_9381,N_3764,N_4068);
nand U9382 (N_9382,N_1651,N_5345);
nor U9383 (N_9383,N_1132,N_86);
or U9384 (N_9384,N_928,N_5280);
or U9385 (N_9385,N_214,N_1060);
nor U9386 (N_9386,N_2604,N_534);
nand U9387 (N_9387,N_3984,N_3817);
nand U9388 (N_9388,N_1226,N_5457);
or U9389 (N_9389,N_1107,N_3648);
xnor U9390 (N_9390,N_4246,N_266);
or U9391 (N_9391,N_448,N_5369);
nor U9392 (N_9392,N_2994,N_3047);
xnor U9393 (N_9393,N_2851,N_1168);
and U9394 (N_9394,N_1036,N_1792);
or U9395 (N_9395,N_99,N_3436);
and U9396 (N_9396,N_5502,N_4604);
and U9397 (N_9397,N_5341,N_629);
xor U9398 (N_9398,N_5430,N_4791);
xor U9399 (N_9399,N_5170,N_5147);
and U9400 (N_9400,N_4092,N_3691);
nand U9401 (N_9401,N_3340,N_2942);
nand U9402 (N_9402,N_3834,N_2194);
nor U9403 (N_9403,N_2914,N_1112);
nor U9404 (N_9404,N_584,N_4458);
or U9405 (N_9405,N_1412,N_4859);
nor U9406 (N_9406,N_2370,N_2801);
nand U9407 (N_9407,N_276,N_5369);
nand U9408 (N_9408,N_5509,N_4493);
nor U9409 (N_9409,N_4185,N_4942);
xor U9410 (N_9410,N_1320,N_2395);
nand U9411 (N_9411,N_2408,N_4676);
nor U9412 (N_9412,N_3749,N_3362);
xnor U9413 (N_9413,N_1055,N_4149);
xnor U9414 (N_9414,N_995,N_1049);
or U9415 (N_9415,N_5497,N_297);
nor U9416 (N_9416,N_5179,N_4119);
nor U9417 (N_9417,N_4378,N_822);
or U9418 (N_9418,N_5421,N_5098);
and U9419 (N_9419,N_5383,N_4213);
xor U9420 (N_9420,N_933,N_3882);
xor U9421 (N_9421,N_5159,N_709);
or U9422 (N_9422,N_3635,N_5136);
nor U9423 (N_9423,N_8,N_2491);
nand U9424 (N_9424,N_2464,N_5175);
or U9425 (N_9425,N_3558,N_1933);
nand U9426 (N_9426,N_3935,N_623);
nand U9427 (N_9427,N_1719,N_1535);
xnor U9428 (N_9428,N_751,N_2600);
and U9429 (N_9429,N_3090,N_2935);
or U9430 (N_9430,N_949,N_1483);
or U9431 (N_9431,N_1820,N_1981);
nand U9432 (N_9432,N_1710,N_5558);
nor U9433 (N_9433,N_4216,N_2278);
nand U9434 (N_9434,N_3690,N_1757);
or U9435 (N_9435,N_1184,N_5332);
nor U9436 (N_9436,N_1313,N_758);
nand U9437 (N_9437,N_3396,N_190);
xor U9438 (N_9438,N_5433,N_2500);
xnor U9439 (N_9439,N_3159,N_2853);
or U9440 (N_9440,N_4399,N_1180);
nor U9441 (N_9441,N_5784,N_1468);
or U9442 (N_9442,N_1569,N_5048);
or U9443 (N_9443,N_4555,N_5897);
and U9444 (N_9444,N_2456,N_662);
xnor U9445 (N_9445,N_2073,N_5107);
nor U9446 (N_9446,N_408,N_3661);
nand U9447 (N_9447,N_84,N_2710);
nor U9448 (N_9448,N_4656,N_3543);
xor U9449 (N_9449,N_4450,N_1184);
and U9450 (N_9450,N_2190,N_3576);
and U9451 (N_9451,N_119,N_220);
xnor U9452 (N_9452,N_407,N_2785);
or U9453 (N_9453,N_1307,N_1155);
or U9454 (N_9454,N_5463,N_2135);
xor U9455 (N_9455,N_4713,N_3310);
or U9456 (N_9456,N_2291,N_1436);
or U9457 (N_9457,N_5695,N_1375);
nor U9458 (N_9458,N_3095,N_2493);
or U9459 (N_9459,N_2392,N_2693);
and U9460 (N_9460,N_5250,N_2182);
or U9461 (N_9461,N_2308,N_3430);
xnor U9462 (N_9462,N_3296,N_1829);
xnor U9463 (N_9463,N_5299,N_4202);
and U9464 (N_9464,N_4410,N_489);
nor U9465 (N_9465,N_1779,N_1261);
nor U9466 (N_9466,N_1770,N_4264);
nand U9467 (N_9467,N_4985,N_855);
nand U9468 (N_9468,N_5497,N_3810);
xor U9469 (N_9469,N_5586,N_5484);
or U9470 (N_9470,N_2289,N_1168);
nand U9471 (N_9471,N_4025,N_1402);
or U9472 (N_9472,N_3992,N_3635);
xnor U9473 (N_9473,N_819,N_4612);
nand U9474 (N_9474,N_3248,N_2971);
or U9475 (N_9475,N_2732,N_4066);
or U9476 (N_9476,N_791,N_738);
or U9477 (N_9477,N_171,N_3737);
nand U9478 (N_9478,N_1435,N_3698);
nand U9479 (N_9479,N_4015,N_1641);
or U9480 (N_9480,N_1553,N_954);
and U9481 (N_9481,N_3265,N_3970);
xnor U9482 (N_9482,N_1836,N_1772);
or U9483 (N_9483,N_1235,N_4713);
nor U9484 (N_9484,N_4259,N_5398);
and U9485 (N_9485,N_1209,N_230);
xor U9486 (N_9486,N_5283,N_0);
nor U9487 (N_9487,N_2122,N_2078);
and U9488 (N_9488,N_4025,N_4557);
or U9489 (N_9489,N_5581,N_4983);
nor U9490 (N_9490,N_3088,N_1944);
xor U9491 (N_9491,N_5004,N_2791);
and U9492 (N_9492,N_909,N_3310);
or U9493 (N_9493,N_3249,N_2712);
nor U9494 (N_9494,N_13,N_4234);
and U9495 (N_9495,N_815,N_2046);
or U9496 (N_9496,N_3075,N_652);
or U9497 (N_9497,N_1060,N_5913);
xnor U9498 (N_9498,N_1258,N_1563);
xnor U9499 (N_9499,N_2554,N_5272);
nor U9500 (N_9500,N_3639,N_3939);
nor U9501 (N_9501,N_3297,N_5243);
nor U9502 (N_9502,N_3818,N_5806);
or U9503 (N_9503,N_3358,N_1275);
nand U9504 (N_9504,N_449,N_4934);
nor U9505 (N_9505,N_2304,N_1801);
or U9506 (N_9506,N_5251,N_2739);
xnor U9507 (N_9507,N_4990,N_4414);
or U9508 (N_9508,N_5160,N_4818);
nand U9509 (N_9509,N_2868,N_2213);
and U9510 (N_9510,N_3046,N_3182);
xnor U9511 (N_9511,N_536,N_3843);
nor U9512 (N_9512,N_5350,N_3184);
and U9513 (N_9513,N_2669,N_4325);
and U9514 (N_9514,N_1643,N_509);
xor U9515 (N_9515,N_3429,N_2572);
and U9516 (N_9516,N_807,N_3074);
xor U9517 (N_9517,N_3331,N_1479);
nor U9518 (N_9518,N_5583,N_900);
or U9519 (N_9519,N_4717,N_3236);
or U9520 (N_9520,N_2470,N_3560);
nor U9521 (N_9521,N_626,N_5282);
nand U9522 (N_9522,N_4824,N_1947);
or U9523 (N_9523,N_2821,N_5617);
xor U9524 (N_9524,N_2004,N_2076);
nand U9525 (N_9525,N_3459,N_5087);
nor U9526 (N_9526,N_2017,N_2243);
nor U9527 (N_9527,N_3379,N_4150);
nor U9528 (N_9528,N_788,N_427);
or U9529 (N_9529,N_1333,N_1370);
and U9530 (N_9530,N_63,N_5130);
xnor U9531 (N_9531,N_2873,N_5801);
nand U9532 (N_9532,N_2223,N_2409);
nand U9533 (N_9533,N_1245,N_3452);
or U9534 (N_9534,N_32,N_5973);
nor U9535 (N_9535,N_4681,N_4583);
and U9536 (N_9536,N_2771,N_1986);
xnor U9537 (N_9537,N_2385,N_4603);
nor U9538 (N_9538,N_1931,N_1614);
nor U9539 (N_9539,N_1905,N_4324);
nor U9540 (N_9540,N_257,N_60);
nor U9541 (N_9541,N_4318,N_699);
or U9542 (N_9542,N_5433,N_1583);
or U9543 (N_9543,N_1427,N_1751);
xor U9544 (N_9544,N_1267,N_4527);
nor U9545 (N_9545,N_4732,N_4286);
nor U9546 (N_9546,N_171,N_541);
nand U9547 (N_9547,N_4871,N_3435);
nor U9548 (N_9548,N_654,N_5120);
or U9549 (N_9549,N_3614,N_5338);
or U9550 (N_9550,N_5303,N_3964);
or U9551 (N_9551,N_3539,N_3921);
nor U9552 (N_9552,N_3488,N_4894);
and U9553 (N_9553,N_1083,N_5152);
xnor U9554 (N_9554,N_2855,N_5350);
or U9555 (N_9555,N_2582,N_3);
nand U9556 (N_9556,N_2985,N_5813);
nand U9557 (N_9557,N_5205,N_5501);
nor U9558 (N_9558,N_251,N_1028);
xor U9559 (N_9559,N_570,N_2655);
or U9560 (N_9560,N_1754,N_1618);
nor U9561 (N_9561,N_1747,N_1146);
or U9562 (N_9562,N_4987,N_3908);
nor U9563 (N_9563,N_2536,N_1432);
nor U9564 (N_9564,N_5156,N_4087);
and U9565 (N_9565,N_4030,N_683);
and U9566 (N_9566,N_4256,N_962);
and U9567 (N_9567,N_669,N_2633);
nand U9568 (N_9568,N_1941,N_1473);
nand U9569 (N_9569,N_4604,N_4456);
nor U9570 (N_9570,N_3829,N_2455);
nand U9571 (N_9571,N_52,N_647);
or U9572 (N_9572,N_433,N_5347);
nor U9573 (N_9573,N_2021,N_3135);
and U9574 (N_9574,N_103,N_1887);
nand U9575 (N_9575,N_3700,N_4754);
nor U9576 (N_9576,N_150,N_3977);
nor U9577 (N_9577,N_3799,N_1653);
nor U9578 (N_9578,N_4819,N_3454);
nor U9579 (N_9579,N_1182,N_1013);
xor U9580 (N_9580,N_2370,N_508);
xnor U9581 (N_9581,N_1563,N_466);
or U9582 (N_9582,N_3019,N_806);
and U9583 (N_9583,N_5136,N_996);
nor U9584 (N_9584,N_5658,N_4213);
or U9585 (N_9585,N_3311,N_5088);
or U9586 (N_9586,N_2769,N_5125);
and U9587 (N_9587,N_2250,N_3922);
nand U9588 (N_9588,N_5526,N_536);
nor U9589 (N_9589,N_1269,N_2064);
xor U9590 (N_9590,N_3371,N_2035);
xor U9591 (N_9591,N_5276,N_988);
nand U9592 (N_9592,N_145,N_3331);
and U9593 (N_9593,N_93,N_2182);
nor U9594 (N_9594,N_20,N_75);
xnor U9595 (N_9595,N_232,N_403);
nor U9596 (N_9596,N_4617,N_2028);
or U9597 (N_9597,N_4842,N_4896);
nor U9598 (N_9598,N_1176,N_1919);
xor U9599 (N_9599,N_1477,N_2780);
xor U9600 (N_9600,N_3529,N_4509);
nand U9601 (N_9601,N_448,N_237);
nand U9602 (N_9602,N_4618,N_2240);
nor U9603 (N_9603,N_849,N_4199);
and U9604 (N_9604,N_851,N_4857);
xnor U9605 (N_9605,N_832,N_3281);
xor U9606 (N_9606,N_2364,N_444);
xnor U9607 (N_9607,N_527,N_2437);
or U9608 (N_9608,N_4222,N_897);
nor U9609 (N_9609,N_501,N_1318);
nor U9610 (N_9610,N_4305,N_5917);
nand U9611 (N_9611,N_2367,N_5251);
nand U9612 (N_9612,N_1427,N_4832);
or U9613 (N_9613,N_4750,N_2189);
or U9614 (N_9614,N_4273,N_4509);
xor U9615 (N_9615,N_1045,N_2095);
xor U9616 (N_9616,N_3158,N_2956);
nand U9617 (N_9617,N_1877,N_5303);
nor U9618 (N_9618,N_1987,N_2737);
nor U9619 (N_9619,N_4336,N_5676);
and U9620 (N_9620,N_1294,N_3215);
and U9621 (N_9621,N_3090,N_4424);
nor U9622 (N_9622,N_5928,N_2899);
and U9623 (N_9623,N_5699,N_2084);
nand U9624 (N_9624,N_3287,N_5963);
nor U9625 (N_9625,N_5047,N_351);
or U9626 (N_9626,N_4940,N_5414);
or U9627 (N_9627,N_3027,N_5767);
and U9628 (N_9628,N_3497,N_4531);
nand U9629 (N_9629,N_623,N_1993);
and U9630 (N_9630,N_3386,N_1894);
or U9631 (N_9631,N_350,N_2464);
or U9632 (N_9632,N_385,N_5460);
nor U9633 (N_9633,N_1681,N_3813);
nand U9634 (N_9634,N_3151,N_810);
or U9635 (N_9635,N_4449,N_1520);
and U9636 (N_9636,N_5840,N_4501);
or U9637 (N_9637,N_4482,N_2152);
nor U9638 (N_9638,N_2943,N_3802);
and U9639 (N_9639,N_4550,N_355);
and U9640 (N_9640,N_549,N_4148);
xnor U9641 (N_9641,N_5673,N_3088);
xor U9642 (N_9642,N_279,N_2795);
nor U9643 (N_9643,N_4866,N_1780);
xnor U9644 (N_9644,N_3652,N_9);
and U9645 (N_9645,N_4027,N_3340);
nor U9646 (N_9646,N_4383,N_5573);
xnor U9647 (N_9647,N_3452,N_5115);
nor U9648 (N_9648,N_3898,N_5239);
nand U9649 (N_9649,N_4359,N_3685);
xor U9650 (N_9650,N_1716,N_4851);
and U9651 (N_9651,N_4778,N_2188);
nand U9652 (N_9652,N_3898,N_1152);
nor U9653 (N_9653,N_1986,N_1966);
and U9654 (N_9654,N_149,N_1817);
or U9655 (N_9655,N_49,N_992);
and U9656 (N_9656,N_3998,N_2685);
and U9657 (N_9657,N_5014,N_1462);
and U9658 (N_9658,N_1665,N_2628);
nand U9659 (N_9659,N_3419,N_2721);
nor U9660 (N_9660,N_1531,N_3683);
xor U9661 (N_9661,N_2313,N_877);
nor U9662 (N_9662,N_4908,N_4217);
or U9663 (N_9663,N_1987,N_3781);
and U9664 (N_9664,N_1488,N_471);
nor U9665 (N_9665,N_1189,N_3728);
nand U9666 (N_9666,N_4255,N_1644);
nand U9667 (N_9667,N_2975,N_5186);
nor U9668 (N_9668,N_5997,N_4185);
xnor U9669 (N_9669,N_4077,N_1164);
nand U9670 (N_9670,N_103,N_1297);
xnor U9671 (N_9671,N_5242,N_2866);
and U9672 (N_9672,N_5959,N_847);
or U9673 (N_9673,N_1283,N_2407);
or U9674 (N_9674,N_3003,N_5438);
nor U9675 (N_9675,N_5283,N_1905);
xnor U9676 (N_9676,N_1336,N_990);
xnor U9677 (N_9677,N_5664,N_2162);
nand U9678 (N_9678,N_2738,N_1579);
nand U9679 (N_9679,N_1657,N_1268);
nor U9680 (N_9680,N_1441,N_672);
and U9681 (N_9681,N_4001,N_2703);
nand U9682 (N_9682,N_567,N_247);
nor U9683 (N_9683,N_1132,N_2942);
or U9684 (N_9684,N_1189,N_668);
nand U9685 (N_9685,N_2821,N_1988);
and U9686 (N_9686,N_1836,N_3484);
nor U9687 (N_9687,N_2613,N_4943);
xnor U9688 (N_9688,N_4514,N_5725);
and U9689 (N_9689,N_2048,N_2966);
or U9690 (N_9690,N_5858,N_2712);
or U9691 (N_9691,N_5798,N_5292);
xnor U9692 (N_9692,N_3380,N_765);
nand U9693 (N_9693,N_5179,N_2801);
nor U9694 (N_9694,N_2774,N_576);
xnor U9695 (N_9695,N_1557,N_1586);
xnor U9696 (N_9696,N_1231,N_5517);
or U9697 (N_9697,N_780,N_803);
and U9698 (N_9698,N_5516,N_3987);
or U9699 (N_9699,N_3250,N_2758);
nand U9700 (N_9700,N_5218,N_5656);
nor U9701 (N_9701,N_1775,N_5344);
and U9702 (N_9702,N_2189,N_692);
or U9703 (N_9703,N_172,N_25);
nor U9704 (N_9704,N_2272,N_2257);
or U9705 (N_9705,N_4866,N_5023);
nand U9706 (N_9706,N_5325,N_1889);
and U9707 (N_9707,N_2516,N_713);
xnor U9708 (N_9708,N_2647,N_5281);
and U9709 (N_9709,N_3078,N_5300);
and U9710 (N_9710,N_2288,N_1317);
or U9711 (N_9711,N_5795,N_83);
and U9712 (N_9712,N_2574,N_5283);
nand U9713 (N_9713,N_2307,N_4101);
nor U9714 (N_9714,N_3560,N_3700);
xor U9715 (N_9715,N_5906,N_92);
nor U9716 (N_9716,N_2217,N_4744);
nand U9717 (N_9717,N_5459,N_923);
xnor U9718 (N_9718,N_1093,N_1555);
xnor U9719 (N_9719,N_1158,N_3922);
xor U9720 (N_9720,N_307,N_3193);
and U9721 (N_9721,N_5839,N_2209);
nor U9722 (N_9722,N_300,N_3755);
xnor U9723 (N_9723,N_5581,N_267);
nor U9724 (N_9724,N_3029,N_4387);
nor U9725 (N_9725,N_2311,N_3805);
nand U9726 (N_9726,N_5362,N_1593);
nand U9727 (N_9727,N_1191,N_4607);
nand U9728 (N_9728,N_1219,N_2202);
and U9729 (N_9729,N_3110,N_2625);
nand U9730 (N_9730,N_2144,N_5555);
or U9731 (N_9731,N_3922,N_2770);
nand U9732 (N_9732,N_3937,N_4675);
or U9733 (N_9733,N_2690,N_4693);
nor U9734 (N_9734,N_3341,N_377);
nand U9735 (N_9735,N_1709,N_1903);
nand U9736 (N_9736,N_4347,N_332);
or U9737 (N_9737,N_2245,N_397);
nor U9738 (N_9738,N_1395,N_2263);
xnor U9739 (N_9739,N_1257,N_15);
nand U9740 (N_9740,N_15,N_2197);
nor U9741 (N_9741,N_478,N_1199);
xor U9742 (N_9742,N_3078,N_2299);
nor U9743 (N_9743,N_3170,N_3512);
and U9744 (N_9744,N_1449,N_2003);
or U9745 (N_9745,N_5144,N_1336);
nor U9746 (N_9746,N_5733,N_4169);
and U9747 (N_9747,N_1000,N_4692);
xor U9748 (N_9748,N_45,N_3423);
and U9749 (N_9749,N_5909,N_1124);
nor U9750 (N_9750,N_5316,N_3391);
nor U9751 (N_9751,N_2849,N_2127);
nand U9752 (N_9752,N_2798,N_4988);
xnor U9753 (N_9753,N_2364,N_5081);
nand U9754 (N_9754,N_392,N_2239);
nor U9755 (N_9755,N_5990,N_3110);
and U9756 (N_9756,N_1414,N_1902);
and U9757 (N_9757,N_1051,N_3210);
and U9758 (N_9758,N_835,N_4430);
nor U9759 (N_9759,N_666,N_2697);
or U9760 (N_9760,N_2716,N_1038);
or U9761 (N_9761,N_4135,N_753);
and U9762 (N_9762,N_4006,N_2987);
nand U9763 (N_9763,N_3819,N_5460);
or U9764 (N_9764,N_34,N_5477);
xor U9765 (N_9765,N_4301,N_70);
nand U9766 (N_9766,N_3384,N_3366);
nand U9767 (N_9767,N_2144,N_611);
nor U9768 (N_9768,N_4097,N_5908);
and U9769 (N_9769,N_2984,N_1901);
and U9770 (N_9770,N_2566,N_313);
xor U9771 (N_9771,N_3511,N_4531);
nor U9772 (N_9772,N_293,N_5847);
nor U9773 (N_9773,N_5145,N_2099);
nand U9774 (N_9774,N_12,N_517);
nor U9775 (N_9775,N_2799,N_359);
and U9776 (N_9776,N_3399,N_4648);
xor U9777 (N_9777,N_3150,N_4758);
xor U9778 (N_9778,N_1872,N_5578);
or U9779 (N_9779,N_979,N_3355);
nand U9780 (N_9780,N_5861,N_5057);
or U9781 (N_9781,N_153,N_4731);
nand U9782 (N_9782,N_1280,N_1066);
nor U9783 (N_9783,N_5605,N_1627);
and U9784 (N_9784,N_3164,N_2352);
or U9785 (N_9785,N_3172,N_1804);
or U9786 (N_9786,N_3202,N_323);
nor U9787 (N_9787,N_3869,N_1839);
or U9788 (N_9788,N_4440,N_2383);
xor U9789 (N_9789,N_4002,N_3363);
nand U9790 (N_9790,N_5671,N_887);
nor U9791 (N_9791,N_1150,N_2275);
nor U9792 (N_9792,N_1870,N_3100);
or U9793 (N_9793,N_5659,N_5216);
xnor U9794 (N_9794,N_2440,N_4863);
and U9795 (N_9795,N_2977,N_3721);
and U9796 (N_9796,N_5145,N_3309);
nand U9797 (N_9797,N_5695,N_1966);
nand U9798 (N_9798,N_5776,N_4312);
nand U9799 (N_9799,N_4734,N_1649);
nand U9800 (N_9800,N_4670,N_1611);
nor U9801 (N_9801,N_4961,N_3840);
or U9802 (N_9802,N_5588,N_2430);
xor U9803 (N_9803,N_4054,N_5158);
xor U9804 (N_9804,N_5810,N_1966);
and U9805 (N_9805,N_4758,N_4461);
or U9806 (N_9806,N_1222,N_4689);
nand U9807 (N_9807,N_4202,N_3127);
xnor U9808 (N_9808,N_4651,N_4114);
nand U9809 (N_9809,N_1291,N_8);
nor U9810 (N_9810,N_4149,N_30);
nand U9811 (N_9811,N_1785,N_2001);
nand U9812 (N_9812,N_3889,N_3088);
xnor U9813 (N_9813,N_2560,N_153);
nor U9814 (N_9814,N_2789,N_5583);
and U9815 (N_9815,N_2400,N_5114);
or U9816 (N_9816,N_3795,N_4871);
nand U9817 (N_9817,N_963,N_4232);
nor U9818 (N_9818,N_3674,N_5668);
or U9819 (N_9819,N_4622,N_5760);
or U9820 (N_9820,N_555,N_300);
nor U9821 (N_9821,N_5347,N_4250);
or U9822 (N_9822,N_2629,N_5798);
and U9823 (N_9823,N_5222,N_5592);
xnor U9824 (N_9824,N_357,N_460);
and U9825 (N_9825,N_1794,N_5628);
or U9826 (N_9826,N_5633,N_3586);
and U9827 (N_9827,N_5702,N_687);
xor U9828 (N_9828,N_1987,N_5426);
nor U9829 (N_9829,N_2742,N_2595);
nand U9830 (N_9830,N_2632,N_86);
or U9831 (N_9831,N_402,N_1482);
or U9832 (N_9832,N_4281,N_2817);
or U9833 (N_9833,N_5405,N_4650);
or U9834 (N_9834,N_425,N_4421);
and U9835 (N_9835,N_4837,N_3600);
nand U9836 (N_9836,N_5118,N_459);
and U9837 (N_9837,N_2404,N_3254);
nand U9838 (N_9838,N_3343,N_4546);
nand U9839 (N_9839,N_3310,N_1747);
nor U9840 (N_9840,N_1266,N_5374);
nor U9841 (N_9841,N_5605,N_3672);
xor U9842 (N_9842,N_3405,N_3205);
nand U9843 (N_9843,N_131,N_1539);
xnor U9844 (N_9844,N_4768,N_5985);
and U9845 (N_9845,N_998,N_1002);
or U9846 (N_9846,N_964,N_624);
or U9847 (N_9847,N_1715,N_1677);
nand U9848 (N_9848,N_2413,N_4838);
or U9849 (N_9849,N_4188,N_2339);
or U9850 (N_9850,N_506,N_608);
nand U9851 (N_9851,N_2293,N_2283);
and U9852 (N_9852,N_2677,N_3450);
nand U9853 (N_9853,N_3684,N_674);
nor U9854 (N_9854,N_159,N_1915);
nor U9855 (N_9855,N_614,N_4339);
nand U9856 (N_9856,N_3891,N_5866);
xnor U9857 (N_9857,N_1616,N_3926);
xnor U9858 (N_9858,N_5230,N_283);
xnor U9859 (N_9859,N_5563,N_3881);
nand U9860 (N_9860,N_1651,N_1894);
nor U9861 (N_9861,N_1551,N_720);
nand U9862 (N_9862,N_4481,N_2203);
and U9863 (N_9863,N_4393,N_2277);
and U9864 (N_9864,N_2050,N_3485);
xnor U9865 (N_9865,N_3147,N_1837);
nand U9866 (N_9866,N_1690,N_420);
and U9867 (N_9867,N_552,N_2558);
and U9868 (N_9868,N_2175,N_4062);
or U9869 (N_9869,N_4949,N_4018);
and U9870 (N_9870,N_2035,N_2884);
and U9871 (N_9871,N_853,N_963);
or U9872 (N_9872,N_647,N_1203);
nor U9873 (N_9873,N_2864,N_4700);
xor U9874 (N_9874,N_1913,N_3191);
nand U9875 (N_9875,N_5214,N_2389);
and U9876 (N_9876,N_868,N_2725);
nor U9877 (N_9877,N_5437,N_412);
nand U9878 (N_9878,N_3907,N_997);
nor U9879 (N_9879,N_414,N_2486);
or U9880 (N_9880,N_3766,N_5738);
nor U9881 (N_9881,N_4726,N_4412);
xor U9882 (N_9882,N_4577,N_4301);
and U9883 (N_9883,N_988,N_3402);
and U9884 (N_9884,N_106,N_4548);
nand U9885 (N_9885,N_5295,N_3827);
or U9886 (N_9886,N_1546,N_1084);
nand U9887 (N_9887,N_872,N_3607);
xor U9888 (N_9888,N_5023,N_4232);
and U9889 (N_9889,N_720,N_1519);
nand U9890 (N_9890,N_1076,N_52);
or U9891 (N_9891,N_2044,N_4116);
xor U9892 (N_9892,N_5501,N_1096);
and U9893 (N_9893,N_428,N_5958);
and U9894 (N_9894,N_565,N_232);
or U9895 (N_9895,N_2193,N_3076);
or U9896 (N_9896,N_3430,N_5054);
nand U9897 (N_9897,N_2034,N_70);
or U9898 (N_9898,N_948,N_802);
nor U9899 (N_9899,N_2644,N_205);
xnor U9900 (N_9900,N_1470,N_3264);
or U9901 (N_9901,N_3738,N_752);
nor U9902 (N_9902,N_4984,N_1987);
and U9903 (N_9903,N_63,N_5703);
and U9904 (N_9904,N_2150,N_2063);
xor U9905 (N_9905,N_1492,N_385);
and U9906 (N_9906,N_5592,N_5839);
nor U9907 (N_9907,N_1219,N_4980);
and U9908 (N_9908,N_3354,N_1369);
or U9909 (N_9909,N_307,N_1248);
nand U9910 (N_9910,N_2785,N_2488);
nor U9911 (N_9911,N_2008,N_2753);
nand U9912 (N_9912,N_5392,N_5699);
and U9913 (N_9913,N_3099,N_1253);
or U9914 (N_9914,N_262,N_688);
xnor U9915 (N_9915,N_1170,N_2479);
nor U9916 (N_9916,N_3305,N_4511);
nor U9917 (N_9917,N_3564,N_5376);
or U9918 (N_9918,N_4430,N_1744);
xor U9919 (N_9919,N_5529,N_2303);
xor U9920 (N_9920,N_4852,N_5874);
nand U9921 (N_9921,N_3463,N_2557);
nor U9922 (N_9922,N_1114,N_4952);
nand U9923 (N_9923,N_2425,N_431);
or U9924 (N_9924,N_2340,N_4280);
xor U9925 (N_9925,N_2737,N_94);
nor U9926 (N_9926,N_720,N_5580);
or U9927 (N_9927,N_5663,N_2403);
nor U9928 (N_9928,N_5549,N_3076);
nand U9929 (N_9929,N_1746,N_2754);
and U9930 (N_9930,N_3143,N_1885);
or U9931 (N_9931,N_3591,N_3156);
or U9932 (N_9932,N_859,N_803);
nand U9933 (N_9933,N_4813,N_4730);
nand U9934 (N_9934,N_4994,N_1766);
nor U9935 (N_9935,N_2481,N_1118);
nor U9936 (N_9936,N_681,N_1919);
nand U9937 (N_9937,N_2829,N_372);
nor U9938 (N_9938,N_2487,N_2191);
or U9939 (N_9939,N_3312,N_5461);
and U9940 (N_9940,N_732,N_2201);
nor U9941 (N_9941,N_3463,N_1933);
nand U9942 (N_9942,N_3725,N_3036);
xor U9943 (N_9943,N_2467,N_5756);
nor U9944 (N_9944,N_3448,N_5527);
and U9945 (N_9945,N_2774,N_1726);
nand U9946 (N_9946,N_2606,N_2662);
or U9947 (N_9947,N_5051,N_618);
nor U9948 (N_9948,N_5497,N_5996);
xor U9949 (N_9949,N_597,N_1906);
nand U9950 (N_9950,N_1351,N_4497);
and U9951 (N_9951,N_4892,N_3079);
or U9952 (N_9952,N_3538,N_2815);
or U9953 (N_9953,N_3142,N_5039);
and U9954 (N_9954,N_150,N_1760);
and U9955 (N_9955,N_4235,N_449);
and U9956 (N_9956,N_331,N_2427);
nand U9957 (N_9957,N_4817,N_3296);
nor U9958 (N_9958,N_5395,N_1601);
or U9959 (N_9959,N_5374,N_2675);
or U9960 (N_9960,N_4290,N_3031);
nor U9961 (N_9961,N_5779,N_2269);
and U9962 (N_9962,N_3643,N_1520);
and U9963 (N_9963,N_3970,N_5778);
and U9964 (N_9964,N_5065,N_4023);
nand U9965 (N_9965,N_5580,N_2375);
and U9966 (N_9966,N_2482,N_5851);
nand U9967 (N_9967,N_5474,N_3980);
and U9968 (N_9968,N_2958,N_1125);
nor U9969 (N_9969,N_1021,N_3268);
nor U9970 (N_9970,N_326,N_5233);
xnor U9971 (N_9971,N_1410,N_3458);
nand U9972 (N_9972,N_5882,N_1796);
xnor U9973 (N_9973,N_4353,N_2317);
nand U9974 (N_9974,N_4719,N_1698);
nor U9975 (N_9975,N_3244,N_453);
nand U9976 (N_9976,N_662,N_2453);
and U9977 (N_9977,N_1707,N_1853);
xnor U9978 (N_9978,N_2938,N_1636);
xor U9979 (N_9979,N_5162,N_5774);
or U9980 (N_9980,N_1862,N_4600);
nor U9981 (N_9981,N_1157,N_2501);
xnor U9982 (N_9982,N_108,N_4395);
nand U9983 (N_9983,N_4117,N_4603);
xnor U9984 (N_9984,N_3388,N_915);
or U9985 (N_9985,N_4244,N_1935);
nor U9986 (N_9986,N_2065,N_3095);
nand U9987 (N_9987,N_4760,N_741);
and U9988 (N_9988,N_665,N_3478);
or U9989 (N_9989,N_2087,N_242);
nor U9990 (N_9990,N_1873,N_1);
or U9991 (N_9991,N_1702,N_1258);
nor U9992 (N_9992,N_1415,N_5376);
xor U9993 (N_9993,N_2847,N_2005);
or U9994 (N_9994,N_5775,N_2335);
xor U9995 (N_9995,N_1663,N_1345);
or U9996 (N_9996,N_4904,N_3562);
and U9997 (N_9997,N_4139,N_5811);
and U9998 (N_9998,N_903,N_5877);
and U9999 (N_9999,N_3545,N_4442);
nand U10000 (N_10000,N_5499,N_66);
xnor U10001 (N_10001,N_4617,N_283);
or U10002 (N_10002,N_2228,N_1327);
and U10003 (N_10003,N_10,N_4478);
and U10004 (N_10004,N_5451,N_5241);
and U10005 (N_10005,N_2661,N_2372);
xor U10006 (N_10006,N_4525,N_74);
nor U10007 (N_10007,N_3798,N_891);
xor U10008 (N_10008,N_823,N_4785);
or U10009 (N_10009,N_538,N_2486);
or U10010 (N_10010,N_345,N_0);
and U10011 (N_10011,N_5448,N_4431);
xor U10012 (N_10012,N_5682,N_2328);
nor U10013 (N_10013,N_4868,N_4735);
nor U10014 (N_10014,N_863,N_3341);
or U10015 (N_10015,N_2927,N_1727);
nor U10016 (N_10016,N_5657,N_1122);
or U10017 (N_10017,N_3739,N_3053);
nor U10018 (N_10018,N_831,N_3300);
nor U10019 (N_10019,N_3438,N_4132);
nor U10020 (N_10020,N_4775,N_5403);
nand U10021 (N_10021,N_3803,N_5900);
or U10022 (N_10022,N_3973,N_3617);
or U10023 (N_10023,N_2680,N_1358);
nor U10024 (N_10024,N_3771,N_820);
and U10025 (N_10025,N_2652,N_190);
and U10026 (N_10026,N_2370,N_10);
xor U10027 (N_10027,N_3990,N_5450);
or U10028 (N_10028,N_1196,N_2678);
xnor U10029 (N_10029,N_5105,N_1871);
and U10030 (N_10030,N_5866,N_4026);
nor U10031 (N_10031,N_5998,N_634);
or U10032 (N_10032,N_3780,N_3457);
and U10033 (N_10033,N_5488,N_3191);
nor U10034 (N_10034,N_2720,N_5786);
and U10035 (N_10035,N_159,N_1980);
and U10036 (N_10036,N_4046,N_2606);
nor U10037 (N_10037,N_1923,N_3296);
nand U10038 (N_10038,N_1812,N_3662);
and U10039 (N_10039,N_3705,N_3630);
and U10040 (N_10040,N_1458,N_1028);
nor U10041 (N_10041,N_3468,N_3901);
xor U10042 (N_10042,N_2071,N_321);
and U10043 (N_10043,N_2779,N_4012);
nor U10044 (N_10044,N_2263,N_1275);
xnor U10045 (N_10045,N_1728,N_537);
xor U10046 (N_10046,N_1998,N_3671);
nor U10047 (N_10047,N_5149,N_1905);
nand U10048 (N_10048,N_5937,N_1192);
or U10049 (N_10049,N_1390,N_1557);
and U10050 (N_10050,N_4347,N_1529);
and U10051 (N_10051,N_3877,N_5617);
nor U10052 (N_10052,N_2900,N_4750);
nor U10053 (N_10053,N_4636,N_553);
xor U10054 (N_10054,N_1278,N_8);
xnor U10055 (N_10055,N_4751,N_5521);
nor U10056 (N_10056,N_2068,N_3842);
and U10057 (N_10057,N_5651,N_4177);
nand U10058 (N_10058,N_2534,N_5308);
or U10059 (N_10059,N_5236,N_390);
xor U10060 (N_10060,N_5889,N_5446);
nand U10061 (N_10061,N_5146,N_1324);
nand U10062 (N_10062,N_142,N_5296);
or U10063 (N_10063,N_1090,N_2513);
xnor U10064 (N_10064,N_2514,N_2253);
nor U10065 (N_10065,N_4060,N_1681);
nor U10066 (N_10066,N_3738,N_3585);
and U10067 (N_10067,N_2393,N_1810);
nand U10068 (N_10068,N_1817,N_1871);
nor U10069 (N_10069,N_3300,N_5949);
nand U10070 (N_10070,N_3562,N_1548);
nand U10071 (N_10071,N_5524,N_1673);
nor U10072 (N_10072,N_50,N_567);
nand U10073 (N_10073,N_5819,N_168);
or U10074 (N_10074,N_4160,N_17);
xnor U10075 (N_10075,N_2940,N_2972);
or U10076 (N_10076,N_2995,N_4329);
xor U10077 (N_10077,N_5907,N_2643);
nor U10078 (N_10078,N_2816,N_2265);
or U10079 (N_10079,N_5767,N_2830);
xor U10080 (N_10080,N_4208,N_1136);
nor U10081 (N_10081,N_626,N_1130);
nand U10082 (N_10082,N_5772,N_3922);
or U10083 (N_10083,N_2891,N_5322);
or U10084 (N_10084,N_1848,N_2838);
nand U10085 (N_10085,N_1425,N_2623);
xor U10086 (N_10086,N_2000,N_2654);
and U10087 (N_10087,N_1732,N_873);
and U10088 (N_10088,N_3192,N_5644);
or U10089 (N_10089,N_2084,N_4720);
and U10090 (N_10090,N_4184,N_5587);
and U10091 (N_10091,N_1495,N_5884);
and U10092 (N_10092,N_105,N_4602);
nor U10093 (N_10093,N_702,N_5201);
nor U10094 (N_10094,N_677,N_4680);
nand U10095 (N_10095,N_2774,N_3761);
xnor U10096 (N_10096,N_274,N_3784);
and U10097 (N_10097,N_185,N_2210);
or U10098 (N_10098,N_4718,N_5541);
nand U10099 (N_10099,N_2020,N_3717);
xor U10100 (N_10100,N_2879,N_3598);
and U10101 (N_10101,N_2311,N_4426);
and U10102 (N_10102,N_609,N_2323);
xor U10103 (N_10103,N_5232,N_5043);
and U10104 (N_10104,N_3980,N_5528);
xnor U10105 (N_10105,N_3690,N_2852);
xor U10106 (N_10106,N_1500,N_1709);
nor U10107 (N_10107,N_1834,N_176);
or U10108 (N_10108,N_5060,N_120);
or U10109 (N_10109,N_1202,N_3572);
nor U10110 (N_10110,N_1885,N_5789);
xnor U10111 (N_10111,N_3369,N_4350);
xor U10112 (N_10112,N_373,N_2199);
and U10113 (N_10113,N_1958,N_2908);
or U10114 (N_10114,N_3468,N_3613);
nand U10115 (N_10115,N_4588,N_2296);
nor U10116 (N_10116,N_4152,N_5274);
xor U10117 (N_10117,N_4423,N_5919);
or U10118 (N_10118,N_2790,N_2258);
and U10119 (N_10119,N_4616,N_4683);
nor U10120 (N_10120,N_4325,N_436);
or U10121 (N_10121,N_3070,N_5608);
or U10122 (N_10122,N_5939,N_2806);
nand U10123 (N_10123,N_3079,N_570);
or U10124 (N_10124,N_1845,N_2466);
nand U10125 (N_10125,N_4274,N_1266);
nand U10126 (N_10126,N_1795,N_5063);
and U10127 (N_10127,N_2135,N_248);
xnor U10128 (N_10128,N_1128,N_173);
nand U10129 (N_10129,N_1334,N_1942);
xor U10130 (N_10130,N_4940,N_3994);
xor U10131 (N_10131,N_2652,N_898);
nor U10132 (N_10132,N_4725,N_2374);
or U10133 (N_10133,N_371,N_659);
nand U10134 (N_10134,N_3325,N_974);
nand U10135 (N_10135,N_279,N_798);
or U10136 (N_10136,N_2571,N_4667);
xor U10137 (N_10137,N_3647,N_3895);
nor U10138 (N_10138,N_4337,N_1846);
and U10139 (N_10139,N_1610,N_2091);
nor U10140 (N_10140,N_1351,N_5757);
or U10141 (N_10141,N_1574,N_1385);
or U10142 (N_10142,N_832,N_4269);
and U10143 (N_10143,N_5699,N_3607);
and U10144 (N_10144,N_5600,N_5556);
or U10145 (N_10145,N_4456,N_5970);
xnor U10146 (N_10146,N_5005,N_3522);
nand U10147 (N_10147,N_657,N_2373);
nor U10148 (N_10148,N_1571,N_1645);
nand U10149 (N_10149,N_2735,N_3183);
or U10150 (N_10150,N_1739,N_5581);
xor U10151 (N_10151,N_4858,N_2848);
xnor U10152 (N_10152,N_2423,N_325);
nor U10153 (N_10153,N_3118,N_3180);
nor U10154 (N_10154,N_1400,N_4855);
nor U10155 (N_10155,N_4117,N_3816);
nor U10156 (N_10156,N_5638,N_4027);
or U10157 (N_10157,N_1923,N_5519);
or U10158 (N_10158,N_3333,N_2531);
nand U10159 (N_10159,N_1927,N_4537);
xnor U10160 (N_10160,N_5767,N_3488);
and U10161 (N_10161,N_2479,N_1887);
and U10162 (N_10162,N_4245,N_5215);
or U10163 (N_10163,N_4957,N_2617);
nand U10164 (N_10164,N_4130,N_370);
and U10165 (N_10165,N_2535,N_3506);
and U10166 (N_10166,N_3945,N_4123);
nand U10167 (N_10167,N_3135,N_1473);
or U10168 (N_10168,N_5677,N_268);
xnor U10169 (N_10169,N_2679,N_1806);
nor U10170 (N_10170,N_3988,N_160);
and U10171 (N_10171,N_1561,N_1802);
xor U10172 (N_10172,N_2198,N_2160);
xnor U10173 (N_10173,N_237,N_3756);
and U10174 (N_10174,N_2290,N_5334);
nand U10175 (N_10175,N_2968,N_3998);
nor U10176 (N_10176,N_63,N_4525);
nand U10177 (N_10177,N_5045,N_1170);
and U10178 (N_10178,N_1547,N_1137);
xor U10179 (N_10179,N_688,N_3479);
or U10180 (N_10180,N_1389,N_5973);
nand U10181 (N_10181,N_1680,N_1392);
nor U10182 (N_10182,N_1602,N_1712);
xor U10183 (N_10183,N_4624,N_92);
and U10184 (N_10184,N_4848,N_2392);
nor U10185 (N_10185,N_5294,N_3405);
nand U10186 (N_10186,N_3283,N_2209);
and U10187 (N_10187,N_1300,N_2845);
or U10188 (N_10188,N_1602,N_2022);
and U10189 (N_10189,N_460,N_2954);
or U10190 (N_10190,N_81,N_2275);
nor U10191 (N_10191,N_2595,N_1847);
and U10192 (N_10192,N_721,N_3996);
nor U10193 (N_10193,N_4848,N_3770);
nand U10194 (N_10194,N_614,N_2653);
xnor U10195 (N_10195,N_2770,N_161);
and U10196 (N_10196,N_3846,N_1997);
nor U10197 (N_10197,N_926,N_2551);
and U10198 (N_10198,N_3813,N_2372);
or U10199 (N_10199,N_5924,N_2813);
xnor U10200 (N_10200,N_4729,N_3281);
or U10201 (N_10201,N_3262,N_2058);
xnor U10202 (N_10202,N_964,N_565);
xor U10203 (N_10203,N_4219,N_5319);
or U10204 (N_10204,N_1479,N_3915);
nor U10205 (N_10205,N_3485,N_209);
xnor U10206 (N_10206,N_3980,N_1077);
and U10207 (N_10207,N_3410,N_4028);
nor U10208 (N_10208,N_1757,N_1210);
nor U10209 (N_10209,N_209,N_5950);
or U10210 (N_10210,N_594,N_5481);
nor U10211 (N_10211,N_4060,N_4799);
xnor U10212 (N_10212,N_5731,N_2383);
or U10213 (N_10213,N_4684,N_3471);
and U10214 (N_10214,N_5148,N_5459);
and U10215 (N_10215,N_4790,N_4694);
and U10216 (N_10216,N_2076,N_7);
nand U10217 (N_10217,N_2912,N_3297);
or U10218 (N_10218,N_2816,N_5212);
xor U10219 (N_10219,N_1437,N_1420);
and U10220 (N_10220,N_1074,N_2596);
nand U10221 (N_10221,N_4250,N_2470);
nor U10222 (N_10222,N_1421,N_3630);
nor U10223 (N_10223,N_5042,N_822);
nand U10224 (N_10224,N_834,N_3225);
nand U10225 (N_10225,N_944,N_5413);
nor U10226 (N_10226,N_5315,N_477);
or U10227 (N_10227,N_5331,N_347);
or U10228 (N_10228,N_3860,N_3088);
or U10229 (N_10229,N_242,N_3897);
or U10230 (N_10230,N_189,N_4029);
nor U10231 (N_10231,N_3920,N_2119);
nor U10232 (N_10232,N_5806,N_4700);
nand U10233 (N_10233,N_2943,N_1524);
nor U10234 (N_10234,N_769,N_4542);
xor U10235 (N_10235,N_3987,N_2292);
nor U10236 (N_10236,N_38,N_3707);
nand U10237 (N_10237,N_4179,N_3362);
nand U10238 (N_10238,N_3026,N_1076);
and U10239 (N_10239,N_380,N_2505);
or U10240 (N_10240,N_724,N_5328);
or U10241 (N_10241,N_563,N_1586);
xnor U10242 (N_10242,N_5454,N_1336);
or U10243 (N_10243,N_5465,N_3267);
nand U10244 (N_10244,N_3649,N_3421);
nor U10245 (N_10245,N_5886,N_1730);
nor U10246 (N_10246,N_1710,N_5584);
nor U10247 (N_10247,N_4541,N_5438);
and U10248 (N_10248,N_4422,N_4304);
nor U10249 (N_10249,N_4227,N_2629);
nor U10250 (N_10250,N_1594,N_367);
nand U10251 (N_10251,N_1621,N_4773);
nor U10252 (N_10252,N_4601,N_3949);
and U10253 (N_10253,N_519,N_5289);
and U10254 (N_10254,N_365,N_2404);
nor U10255 (N_10255,N_583,N_2958);
nand U10256 (N_10256,N_2806,N_1166);
nand U10257 (N_10257,N_2240,N_1924);
or U10258 (N_10258,N_3461,N_5075);
and U10259 (N_10259,N_2532,N_5553);
nand U10260 (N_10260,N_5648,N_5750);
or U10261 (N_10261,N_4986,N_4946);
and U10262 (N_10262,N_4222,N_5717);
xor U10263 (N_10263,N_4016,N_4964);
xor U10264 (N_10264,N_3926,N_5110);
or U10265 (N_10265,N_2104,N_1922);
or U10266 (N_10266,N_107,N_5158);
nor U10267 (N_10267,N_878,N_4733);
xnor U10268 (N_10268,N_2722,N_3243);
nand U10269 (N_10269,N_5668,N_1641);
nand U10270 (N_10270,N_5182,N_1844);
nor U10271 (N_10271,N_5576,N_727);
nand U10272 (N_10272,N_2508,N_1492);
xor U10273 (N_10273,N_5515,N_4064);
xnor U10274 (N_10274,N_535,N_2252);
or U10275 (N_10275,N_3493,N_3176);
nand U10276 (N_10276,N_3557,N_5869);
nor U10277 (N_10277,N_4165,N_1304);
or U10278 (N_10278,N_117,N_5914);
nor U10279 (N_10279,N_3141,N_1866);
nand U10280 (N_10280,N_5650,N_8);
xor U10281 (N_10281,N_2735,N_3473);
nand U10282 (N_10282,N_1481,N_1245);
and U10283 (N_10283,N_4550,N_4298);
nor U10284 (N_10284,N_1935,N_5434);
nor U10285 (N_10285,N_1780,N_558);
nand U10286 (N_10286,N_2847,N_2426);
nand U10287 (N_10287,N_4301,N_3508);
xnor U10288 (N_10288,N_4184,N_1976);
nand U10289 (N_10289,N_2548,N_1463);
nand U10290 (N_10290,N_5179,N_2755);
nor U10291 (N_10291,N_1216,N_1018);
xor U10292 (N_10292,N_5100,N_3940);
nand U10293 (N_10293,N_4695,N_2998);
and U10294 (N_10294,N_3358,N_5123);
nor U10295 (N_10295,N_2974,N_4560);
nor U10296 (N_10296,N_2350,N_5675);
nor U10297 (N_10297,N_745,N_4984);
nor U10298 (N_10298,N_4302,N_749);
or U10299 (N_10299,N_2975,N_559);
nor U10300 (N_10300,N_642,N_458);
or U10301 (N_10301,N_3783,N_4583);
nor U10302 (N_10302,N_2424,N_4469);
and U10303 (N_10303,N_553,N_1275);
and U10304 (N_10304,N_3158,N_1744);
nor U10305 (N_10305,N_1364,N_2533);
and U10306 (N_10306,N_2040,N_5282);
or U10307 (N_10307,N_4235,N_528);
xor U10308 (N_10308,N_1743,N_2126);
or U10309 (N_10309,N_3619,N_1746);
and U10310 (N_10310,N_5046,N_2736);
xnor U10311 (N_10311,N_5735,N_2821);
nand U10312 (N_10312,N_313,N_1333);
nand U10313 (N_10313,N_5014,N_444);
xnor U10314 (N_10314,N_3690,N_3149);
xor U10315 (N_10315,N_4095,N_1385);
nor U10316 (N_10316,N_5717,N_4525);
xnor U10317 (N_10317,N_1443,N_3335);
nor U10318 (N_10318,N_1010,N_1696);
nor U10319 (N_10319,N_1807,N_4513);
or U10320 (N_10320,N_2432,N_5441);
nand U10321 (N_10321,N_2661,N_1474);
or U10322 (N_10322,N_771,N_1315);
and U10323 (N_10323,N_3738,N_5697);
xor U10324 (N_10324,N_2693,N_1967);
or U10325 (N_10325,N_778,N_566);
xnor U10326 (N_10326,N_2610,N_2347);
or U10327 (N_10327,N_2846,N_5082);
nand U10328 (N_10328,N_304,N_1944);
nor U10329 (N_10329,N_3412,N_39);
and U10330 (N_10330,N_289,N_2818);
xnor U10331 (N_10331,N_5070,N_4552);
xnor U10332 (N_10332,N_2111,N_4093);
nand U10333 (N_10333,N_3338,N_1141);
xnor U10334 (N_10334,N_3709,N_3170);
nand U10335 (N_10335,N_4701,N_4440);
and U10336 (N_10336,N_5306,N_1474);
or U10337 (N_10337,N_4133,N_5211);
or U10338 (N_10338,N_2284,N_1934);
nor U10339 (N_10339,N_2031,N_5835);
xnor U10340 (N_10340,N_2882,N_1398);
nor U10341 (N_10341,N_4523,N_818);
nor U10342 (N_10342,N_1578,N_589);
xor U10343 (N_10343,N_2594,N_3804);
nor U10344 (N_10344,N_3486,N_5455);
or U10345 (N_10345,N_2322,N_2887);
or U10346 (N_10346,N_3292,N_4260);
and U10347 (N_10347,N_4885,N_4016);
or U10348 (N_10348,N_5684,N_2406);
nor U10349 (N_10349,N_5391,N_1332);
nor U10350 (N_10350,N_2049,N_591);
nor U10351 (N_10351,N_503,N_4383);
nor U10352 (N_10352,N_3620,N_1365);
nand U10353 (N_10353,N_4856,N_4217);
nor U10354 (N_10354,N_2183,N_422);
or U10355 (N_10355,N_3223,N_4318);
xor U10356 (N_10356,N_591,N_4850);
nand U10357 (N_10357,N_1639,N_4807);
nand U10358 (N_10358,N_3296,N_208);
nor U10359 (N_10359,N_5181,N_3566);
and U10360 (N_10360,N_3109,N_5647);
xnor U10361 (N_10361,N_379,N_1133);
nand U10362 (N_10362,N_4833,N_2481);
nand U10363 (N_10363,N_4936,N_3275);
xor U10364 (N_10364,N_958,N_5987);
nor U10365 (N_10365,N_4645,N_2291);
or U10366 (N_10366,N_3241,N_5147);
and U10367 (N_10367,N_3010,N_4053);
nand U10368 (N_10368,N_1868,N_1298);
nand U10369 (N_10369,N_3598,N_3956);
and U10370 (N_10370,N_2641,N_5474);
and U10371 (N_10371,N_5851,N_5317);
nor U10372 (N_10372,N_1263,N_4051);
nand U10373 (N_10373,N_1539,N_380);
nand U10374 (N_10374,N_2445,N_1956);
nand U10375 (N_10375,N_3526,N_435);
or U10376 (N_10376,N_4851,N_953);
or U10377 (N_10377,N_3687,N_4671);
or U10378 (N_10378,N_5068,N_1579);
and U10379 (N_10379,N_9,N_1854);
nor U10380 (N_10380,N_5039,N_3079);
nand U10381 (N_10381,N_415,N_5187);
xor U10382 (N_10382,N_1688,N_2583);
or U10383 (N_10383,N_5385,N_5926);
nor U10384 (N_10384,N_3975,N_2353);
or U10385 (N_10385,N_2557,N_3437);
xor U10386 (N_10386,N_2630,N_4286);
nand U10387 (N_10387,N_4685,N_1603);
and U10388 (N_10388,N_5116,N_644);
xnor U10389 (N_10389,N_909,N_726);
or U10390 (N_10390,N_2823,N_4157);
nor U10391 (N_10391,N_3968,N_2665);
nor U10392 (N_10392,N_727,N_4391);
xnor U10393 (N_10393,N_5161,N_3923);
or U10394 (N_10394,N_1647,N_818);
and U10395 (N_10395,N_722,N_4550);
or U10396 (N_10396,N_2694,N_2257);
nand U10397 (N_10397,N_2648,N_698);
nor U10398 (N_10398,N_5597,N_4193);
nand U10399 (N_10399,N_983,N_23);
nand U10400 (N_10400,N_5771,N_611);
and U10401 (N_10401,N_2773,N_668);
and U10402 (N_10402,N_3874,N_3950);
nand U10403 (N_10403,N_5493,N_1378);
nor U10404 (N_10404,N_4196,N_5323);
nor U10405 (N_10405,N_257,N_2969);
and U10406 (N_10406,N_996,N_5892);
nor U10407 (N_10407,N_245,N_3157);
or U10408 (N_10408,N_2257,N_5974);
and U10409 (N_10409,N_4520,N_1911);
nor U10410 (N_10410,N_3017,N_4633);
nor U10411 (N_10411,N_548,N_5164);
nand U10412 (N_10412,N_5126,N_5670);
or U10413 (N_10413,N_3016,N_3766);
or U10414 (N_10414,N_344,N_4790);
xor U10415 (N_10415,N_1465,N_5731);
and U10416 (N_10416,N_3662,N_2535);
or U10417 (N_10417,N_302,N_2783);
or U10418 (N_10418,N_1576,N_210);
xor U10419 (N_10419,N_3771,N_2167);
and U10420 (N_10420,N_1501,N_3676);
nand U10421 (N_10421,N_930,N_372);
or U10422 (N_10422,N_3232,N_4450);
and U10423 (N_10423,N_789,N_4975);
nand U10424 (N_10424,N_2353,N_5369);
xnor U10425 (N_10425,N_437,N_2538);
and U10426 (N_10426,N_197,N_2619);
and U10427 (N_10427,N_5701,N_1886);
and U10428 (N_10428,N_2485,N_3340);
xnor U10429 (N_10429,N_3042,N_845);
nor U10430 (N_10430,N_5150,N_2498);
nand U10431 (N_10431,N_5466,N_2928);
xor U10432 (N_10432,N_5122,N_4227);
or U10433 (N_10433,N_5789,N_2336);
nor U10434 (N_10434,N_1124,N_5368);
or U10435 (N_10435,N_2883,N_4211);
xor U10436 (N_10436,N_4383,N_2837);
and U10437 (N_10437,N_1088,N_1027);
nand U10438 (N_10438,N_5633,N_433);
xor U10439 (N_10439,N_5994,N_2853);
or U10440 (N_10440,N_850,N_4959);
nor U10441 (N_10441,N_4515,N_4800);
or U10442 (N_10442,N_103,N_173);
nand U10443 (N_10443,N_2403,N_5392);
or U10444 (N_10444,N_4698,N_2298);
xor U10445 (N_10445,N_5714,N_35);
nor U10446 (N_10446,N_774,N_5732);
and U10447 (N_10447,N_2367,N_2881);
nor U10448 (N_10448,N_1192,N_315);
or U10449 (N_10449,N_5092,N_3947);
or U10450 (N_10450,N_2075,N_4958);
nand U10451 (N_10451,N_597,N_4748);
nand U10452 (N_10452,N_3677,N_2002);
nor U10453 (N_10453,N_2695,N_5933);
or U10454 (N_10454,N_2608,N_1731);
nand U10455 (N_10455,N_5931,N_3059);
xnor U10456 (N_10456,N_3411,N_1563);
or U10457 (N_10457,N_3242,N_2234);
nor U10458 (N_10458,N_3843,N_5360);
nor U10459 (N_10459,N_3413,N_4809);
and U10460 (N_10460,N_5666,N_1977);
and U10461 (N_10461,N_419,N_1083);
or U10462 (N_10462,N_874,N_5119);
xor U10463 (N_10463,N_3240,N_380);
xor U10464 (N_10464,N_5621,N_740);
nand U10465 (N_10465,N_5933,N_1619);
and U10466 (N_10466,N_683,N_5485);
xnor U10467 (N_10467,N_4126,N_1887);
or U10468 (N_10468,N_3660,N_778);
xnor U10469 (N_10469,N_4530,N_5917);
xor U10470 (N_10470,N_5222,N_1198);
nor U10471 (N_10471,N_3184,N_1777);
nand U10472 (N_10472,N_181,N_3058);
xor U10473 (N_10473,N_555,N_5605);
and U10474 (N_10474,N_5555,N_958);
nor U10475 (N_10475,N_2122,N_2404);
nand U10476 (N_10476,N_5435,N_2601);
nor U10477 (N_10477,N_1684,N_1744);
nor U10478 (N_10478,N_3113,N_299);
or U10479 (N_10479,N_4054,N_1062);
or U10480 (N_10480,N_2250,N_2086);
nor U10481 (N_10481,N_2402,N_4908);
xnor U10482 (N_10482,N_227,N_4138);
nor U10483 (N_10483,N_4999,N_4523);
or U10484 (N_10484,N_5099,N_377);
nor U10485 (N_10485,N_5219,N_2113);
and U10486 (N_10486,N_2599,N_5176);
and U10487 (N_10487,N_1999,N_4788);
and U10488 (N_10488,N_5974,N_4386);
nor U10489 (N_10489,N_1123,N_1148);
and U10490 (N_10490,N_5343,N_510);
or U10491 (N_10491,N_4745,N_874);
nand U10492 (N_10492,N_1694,N_4214);
nand U10493 (N_10493,N_756,N_3888);
nand U10494 (N_10494,N_3519,N_3657);
or U10495 (N_10495,N_1664,N_583);
xnor U10496 (N_10496,N_4223,N_5122);
xor U10497 (N_10497,N_5966,N_326);
or U10498 (N_10498,N_777,N_2533);
xor U10499 (N_10499,N_4483,N_1982);
xor U10500 (N_10500,N_190,N_3573);
or U10501 (N_10501,N_4546,N_3854);
and U10502 (N_10502,N_2674,N_4854);
nand U10503 (N_10503,N_4297,N_4083);
or U10504 (N_10504,N_5009,N_4915);
xnor U10505 (N_10505,N_4544,N_5370);
xor U10506 (N_10506,N_2508,N_4052);
nand U10507 (N_10507,N_2042,N_3994);
or U10508 (N_10508,N_1452,N_4383);
and U10509 (N_10509,N_887,N_4548);
or U10510 (N_10510,N_121,N_18);
nand U10511 (N_10511,N_5333,N_2073);
and U10512 (N_10512,N_4795,N_1664);
and U10513 (N_10513,N_1657,N_3619);
or U10514 (N_10514,N_3883,N_5353);
or U10515 (N_10515,N_342,N_4671);
nand U10516 (N_10516,N_9,N_5473);
and U10517 (N_10517,N_1831,N_4241);
xor U10518 (N_10518,N_2837,N_4727);
nand U10519 (N_10519,N_5444,N_4410);
or U10520 (N_10520,N_2465,N_1807);
and U10521 (N_10521,N_5006,N_78);
and U10522 (N_10522,N_2597,N_1060);
nand U10523 (N_10523,N_2002,N_1857);
xnor U10524 (N_10524,N_4128,N_528);
nor U10525 (N_10525,N_1815,N_5208);
and U10526 (N_10526,N_4573,N_1441);
and U10527 (N_10527,N_2582,N_5506);
nor U10528 (N_10528,N_3846,N_2902);
and U10529 (N_10529,N_3737,N_1565);
nor U10530 (N_10530,N_2346,N_5202);
nor U10531 (N_10531,N_1776,N_2328);
and U10532 (N_10532,N_4247,N_5910);
or U10533 (N_10533,N_448,N_3860);
and U10534 (N_10534,N_2048,N_5240);
nand U10535 (N_10535,N_4266,N_4240);
and U10536 (N_10536,N_1923,N_1194);
and U10537 (N_10537,N_5668,N_3279);
xor U10538 (N_10538,N_2255,N_129);
nor U10539 (N_10539,N_3453,N_4139);
nor U10540 (N_10540,N_3031,N_4319);
xor U10541 (N_10541,N_5362,N_1864);
nand U10542 (N_10542,N_402,N_2829);
or U10543 (N_10543,N_4730,N_3238);
xnor U10544 (N_10544,N_5021,N_3674);
or U10545 (N_10545,N_1078,N_875);
and U10546 (N_10546,N_5028,N_5799);
and U10547 (N_10547,N_4251,N_1983);
xnor U10548 (N_10548,N_3571,N_1484);
and U10549 (N_10549,N_1245,N_5502);
nor U10550 (N_10550,N_4573,N_531);
nand U10551 (N_10551,N_5933,N_1);
or U10552 (N_10552,N_5248,N_860);
nor U10553 (N_10553,N_3949,N_5311);
nand U10554 (N_10554,N_5474,N_2124);
nor U10555 (N_10555,N_2660,N_5899);
xnor U10556 (N_10556,N_4106,N_5446);
xor U10557 (N_10557,N_4221,N_3055);
nor U10558 (N_10558,N_3352,N_2290);
and U10559 (N_10559,N_3086,N_2251);
nor U10560 (N_10560,N_2175,N_2298);
nor U10561 (N_10561,N_4531,N_1916);
and U10562 (N_10562,N_1511,N_5741);
or U10563 (N_10563,N_90,N_1637);
xor U10564 (N_10564,N_3774,N_3746);
or U10565 (N_10565,N_1333,N_5458);
xor U10566 (N_10566,N_4843,N_3681);
nor U10567 (N_10567,N_3817,N_3972);
xor U10568 (N_10568,N_914,N_4467);
xnor U10569 (N_10569,N_5609,N_4494);
xor U10570 (N_10570,N_3828,N_969);
or U10571 (N_10571,N_3013,N_1411);
xnor U10572 (N_10572,N_2699,N_2420);
xor U10573 (N_10573,N_4080,N_2118);
or U10574 (N_10574,N_5105,N_4230);
nor U10575 (N_10575,N_3551,N_953);
and U10576 (N_10576,N_359,N_820);
nor U10577 (N_10577,N_5465,N_3850);
and U10578 (N_10578,N_2923,N_2637);
or U10579 (N_10579,N_5992,N_1297);
and U10580 (N_10580,N_3196,N_5086);
xor U10581 (N_10581,N_3413,N_4220);
nand U10582 (N_10582,N_3848,N_4889);
and U10583 (N_10583,N_2538,N_3708);
nand U10584 (N_10584,N_1083,N_4051);
nor U10585 (N_10585,N_2774,N_5549);
nor U10586 (N_10586,N_2146,N_4770);
nand U10587 (N_10587,N_2805,N_586);
and U10588 (N_10588,N_4751,N_2204);
and U10589 (N_10589,N_3888,N_2600);
xnor U10590 (N_10590,N_3511,N_3209);
xnor U10591 (N_10591,N_3094,N_1583);
nor U10592 (N_10592,N_1462,N_437);
nand U10593 (N_10593,N_5314,N_1412);
nand U10594 (N_10594,N_3756,N_5728);
xnor U10595 (N_10595,N_4484,N_4486);
and U10596 (N_10596,N_5486,N_2451);
nor U10597 (N_10597,N_2218,N_2431);
and U10598 (N_10598,N_817,N_2855);
nor U10599 (N_10599,N_1066,N_1568);
nand U10600 (N_10600,N_173,N_5919);
xnor U10601 (N_10601,N_1135,N_4770);
nor U10602 (N_10602,N_2374,N_444);
nand U10603 (N_10603,N_2425,N_1666);
nor U10604 (N_10604,N_2721,N_5893);
and U10605 (N_10605,N_915,N_4299);
nor U10606 (N_10606,N_4425,N_4549);
nand U10607 (N_10607,N_5013,N_5737);
xnor U10608 (N_10608,N_2661,N_638);
or U10609 (N_10609,N_2548,N_2334);
nand U10610 (N_10610,N_5959,N_1088);
xor U10611 (N_10611,N_4412,N_1498);
nor U10612 (N_10612,N_2946,N_969);
nor U10613 (N_10613,N_3836,N_746);
xor U10614 (N_10614,N_2263,N_1889);
and U10615 (N_10615,N_915,N_465);
nor U10616 (N_10616,N_874,N_2246);
xor U10617 (N_10617,N_600,N_2017);
and U10618 (N_10618,N_5286,N_799);
nand U10619 (N_10619,N_4835,N_2676);
or U10620 (N_10620,N_1852,N_3649);
and U10621 (N_10621,N_3811,N_1296);
or U10622 (N_10622,N_2873,N_144);
xnor U10623 (N_10623,N_4872,N_631);
and U10624 (N_10624,N_5922,N_1422);
nor U10625 (N_10625,N_3966,N_1426);
nand U10626 (N_10626,N_2466,N_770);
nor U10627 (N_10627,N_4725,N_5499);
and U10628 (N_10628,N_5828,N_889);
nor U10629 (N_10629,N_4229,N_5180);
nor U10630 (N_10630,N_1445,N_1223);
or U10631 (N_10631,N_5470,N_4469);
nor U10632 (N_10632,N_2840,N_5185);
and U10633 (N_10633,N_5210,N_2453);
xnor U10634 (N_10634,N_4471,N_3952);
nand U10635 (N_10635,N_2099,N_4091);
nand U10636 (N_10636,N_3431,N_2706);
nor U10637 (N_10637,N_768,N_1869);
nand U10638 (N_10638,N_4236,N_5650);
nand U10639 (N_10639,N_3138,N_3859);
and U10640 (N_10640,N_2828,N_2431);
nand U10641 (N_10641,N_3038,N_5413);
nor U10642 (N_10642,N_43,N_3962);
xor U10643 (N_10643,N_3805,N_1389);
nand U10644 (N_10644,N_4020,N_2514);
nor U10645 (N_10645,N_4155,N_2844);
and U10646 (N_10646,N_2877,N_4406);
nor U10647 (N_10647,N_1125,N_5903);
nor U10648 (N_10648,N_2275,N_3231);
and U10649 (N_10649,N_4441,N_908);
or U10650 (N_10650,N_5656,N_2484);
xor U10651 (N_10651,N_3024,N_4458);
and U10652 (N_10652,N_2553,N_232);
nor U10653 (N_10653,N_131,N_698);
xor U10654 (N_10654,N_1118,N_4008);
or U10655 (N_10655,N_765,N_1243);
xor U10656 (N_10656,N_5097,N_4312);
or U10657 (N_10657,N_2530,N_4349);
xor U10658 (N_10658,N_2867,N_5247);
xor U10659 (N_10659,N_5792,N_2023);
xnor U10660 (N_10660,N_1304,N_2352);
nor U10661 (N_10661,N_1037,N_1765);
and U10662 (N_10662,N_2946,N_3830);
nor U10663 (N_10663,N_1161,N_1662);
and U10664 (N_10664,N_2727,N_331);
nand U10665 (N_10665,N_2689,N_5361);
and U10666 (N_10666,N_2441,N_2985);
xor U10667 (N_10667,N_3865,N_3192);
and U10668 (N_10668,N_1447,N_1606);
nor U10669 (N_10669,N_966,N_59);
nor U10670 (N_10670,N_586,N_4295);
or U10671 (N_10671,N_990,N_3681);
xor U10672 (N_10672,N_5843,N_1823);
nor U10673 (N_10673,N_2042,N_3407);
or U10674 (N_10674,N_515,N_2128);
or U10675 (N_10675,N_4013,N_4956);
and U10676 (N_10676,N_3269,N_5390);
or U10677 (N_10677,N_2072,N_4475);
nor U10678 (N_10678,N_1993,N_949);
nor U10679 (N_10679,N_280,N_1283);
nand U10680 (N_10680,N_3089,N_112);
xor U10681 (N_10681,N_3286,N_5598);
or U10682 (N_10682,N_1879,N_1020);
nor U10683 (N_10683,N_5422,N_1928);
and U10684 (N_10684,N_5343,N_1278);
or U10685 (N_10685,N_27,N_1669);
xnor U10686 (N_10686,N_4329,N_2736);
xnor U10687 (N_10687,N_2017,N_5019);
or U10688 (N_10688,N_808,N_5087);
xor U10689 (N_10689,N_1161,N_443);
and U10690 (N_10690,N_820,N_5405);
nor U10691 (N_10691,N_2539,N_1684);
xor U10692 (N_10692,N_1602,N_5770);
nor U10693 (N_10693,N_4707,N_1540);
or U10694 (N_10694,N_717,N_2753);
or U10695 (N_10695,N_420,N_242);
xor U10696 (N_10696,N_767,N_42);
xnor U10697 (N_10697,N_5568,N_5233);
or U10698 (N_10698,N_1706,N_5116);
xor U10699 (N_10699,N_3400,N_5367);
and U10700 (N_10700,N_4857,N_800);
xnor U10701 (N_10701,N_191,N_1147);
xnor U10702 (N_10702,N_5408,N_861);
xnor U10703 (N_10703,N_1534,N_3416);
nor U10704 (N_10704,N_1995,N_2024);
and U10705 (N_10705,N_267,N_630);
and U10706 (N_10706,N_2602,N_4533);
nor U10707 (N_10707,N_2797,N_583);
xnor U10708 (N_10708,N_3281,N_4473);
nor U10709 (N_10709,N_687,N_4203);
nor U10710 (N_10710,N_1288,N_1889);
nand U10711 (N_10711,N_110,N_4755);
xnor U10712 (N_10712,N_954,N_3664);
or U10713 (N_10713,N_5814,N_5664);
xor U10714 (N_10714,N_3560,N_1641);
nand U10715 (N_10715,N_3268,N_2491);
and U10716 (N_10716,N_582,N_2325);
and U10717 (N_10717,N_1211,N_5858);
nand U10718 (N_10718,N_3377,N_1492);
xnor U10719 (N_10719,N_1497,N_654);
nor U10720 (N_10720,N_1521,N_2373);
nand U10721 (N_10721,N_334,N_836);
and U10722 (N_10722,N_2539,N_1306);
nand U10723 (N_10723,N_1595,N_3432);
nand U10724 (N_10724,N_2896,N_2961);
nand U10725 (N_10725,N_3462,N_167);
nor U10726 (N_10726,N_4874,N_1673);
or U10727 (N_10727,N_1587,N_2532);
nand U10728 (N_10728,N_853,N_5141);
and U10729 (N_10729,N_3433,N_584);
or U10730 (N_10730,N_2806,N_3516);
and U10731 (N_10731,N_5866,N_5344);
or U10732 (N_10732,N_5956,N_4044);
nand U10733 (N_10733,N_934,N_1141);
nand U10734 (N_10734,N_5441,N_4215);
or U10735 (N_10735,N_5990,N_199);
or U10736 (N_10736,N_5358,N_4274);
nor U10737 (N_10737,N_4180,N_2147);
nor U10738 (N_10738,N_3202,N_252);
nor U10739 (N_10739,N_2373,N_5304);
xnor U10740 (N_10740,N_5019,N_4249);
or U10741 (N_10741,N_5435,N_5908);
and U10742 (N_10742,N_3129,N_1612);
xnor U10743 (N_10743,N_4503,N_775);
nand U10744 (N_10744,N_12,N_1515);
nand U10745 (N_10745,N_5785,N_51);
xnor U10746 (N_10746,N_1061,N_1238);
xor U10747 (N_10747,N_3578,N_548);
nand U10748 (N_10748,N_5617,N_1227);
xor U10749 (N_10749,N_3068,N_453);
or U10750 (N_10750,N_3979,N_3404);
nor U10751 (N_10751,N_2494,N_3673);
and U10752 (N_10752,N_1965,N_4716);
nor U10753 (N_10753,N_873,N_955);
or U10754 (N_10754,N_2416,N_1095);
or U10755 (N_10755,N_917,N_1612);
xnor U10756 (N_10756,N_4861,N_848);
xor U10757 (N_10757,N_733,N_788);
nand U10758 (N_10758,N_3341,N_5493);
and U10759 (N_10759,N_225,N_289);
nor U10760 (N_10760,N_5782,N_5216);
and U10761 (N_10761,N_5108,N_5275);
nand U10762 (N_10762,N_2531,N_5129);
xor U10763 (N_10763,N_2491,N_1055);
and U10764 (N_10764,N_3332,N_5484);
xnor U10765 (N_10765,N_269,N_3891);
nor U10766 (N_10766,N_4959,N_5113);
nor U10767 (N_10767,N_4810,N_785);
nand U10768 (N_10768,N_3615,N_4911);
xnor U10769 (N_10769,N_2873,N_4911);
and U10770 (N_10770,N_1227,N_890);
xor U10771 (N_10771,N_3347,N_3892);
xor U10772 (N_10772,N_633,N_4853);
nand U10773 (N_10773,N_602,N_4444);
xnor U10774 (N_10774,N_5055,N_60);
and U10775 (N_10775,N_2547,N_896);
xor U10776 (N_10776,N_5495,N_3158);
and U10777 (N_10777,N_1977,N_2833);
and U10778 (N_10778,N_4884,N_4651);
or U10779 (N_10779,N_3881,N_3214);
or U10780 (N_10780,N_1994,N_5503);
nor U10781 (N_10781,N_2110,N_3217);
nand U10782 (N_10782,N_3022,N_2643);
nor U10783 (N_10783,N_946,N_2865);
nor U10784 (N_10784,N_2663,N_4797);
or U10785 (N_10785,N_5060,N_549);
nand U10786 (N_10786,N_1190,N_995);
and U10787 (N_10787,N_2095,N_4199);
xor U10788 (N_10788,N_5527,N_5141);
or U10789 (N_10789,N_866,N_3274);
and U10790 (N_10790,N_3698,N_2479);
or U10791 (N_10791,N_349,N_5889);
or U10792 (N_10792,N_2998,N_2104);
and U10793 (N_10793,N_165,N_1737);
and U10794 (N_10794,N_4531,N_4461);
or U10795 (N_10795,N_5892,N_3581);
xnor U10796 (N_10796,N_2927,N_1407);
nor U10797 (N_10797,N_4287,N_5641);
and U10798 (N_10798,N_5318,N_481);
nor U10799 (N_10799,N_48,N_5459);
or U10800 (N_10800,N_2029,N_1352);
nor U10801 (N_10801,N_1250,N_3558);
nor U10802 (N_10802,N_4611,N_2973);
or U10803 (N_10803,N_3842,N_4214);
nand U10804 (N_10804,N_2561,N_2255);
nor U10805 (N_10805,N_5416,N_2374);
nor U10806 (N_10806,N_1513,N_502);
nand U10807 (N_10807,N_4377,N_2986);
xor U10808 (N_10808,N_4220,N_5441);
nand U10809 (N_10809,N_4252,N_4543);
nand U10810 (N_10810,N_5595,N_2003);
nand U10811 (N_10811,N_4904,N_3253);
nor U10812 (N_10812,N_3389,N_3040);
nand U10813 (N_10813,N_1286,N_1902);
nor U10814 (N_10814,N_5466,N_5219);
nor U10815 (N_10815,N_2179,N_3564);
and U10816 (N_10816,N_220,N_2959);
xor U10817 (N_10817,N_5403,N_5576);
nor U10818 (N_10818,N_1132,N_3458);
and U10819 (N_10819,N_283,N_312);
and U10820 (N_10820,N_2773,N_4251);
xnor U10821 (N_10821,N_5851,N_1607);
nor U10822 (N_10822,N_4342,N_325);
nand U10823 (N_10823,N_3297,N_3290);
xnor U10824 (N_10824,N_420,N_5110);
and U10825 (N_10825,N_927,N_2006);
and U10826 (N_10826,N_1563,N_4227);
and U10827 (N_10827,N_2682,N_3263);
or U10828 (N_10828,N_1093,N_5158);
or U10829 (N_10829,N_3248,N_3296);
nor U10830 (N_10830,N_2424,N_4546);
nor U10831 (N_10831,N_2455,N_1777);
nor U10832 (N_10832,N_3937,N_2245);
or U10833 (N_10833,N_49,N_4218);
and U10834 (N_10834,N_5737,N_3131);
nor U10835 (N_10835,N_1281,N_5901);
nand U10836 (N_10836,N_5252,N_4554);
xnor U10837 (N_10837,N_1472,N_1499);
xnor U10838 (N_10838,N_5991,N_1376);
xnor U10839 (N_10839,N_2087,N_2906);
xnor U10840 (N_10840,N_4860,N_1259);
or U10841 (N_10841,N_5773,N_2865);
nand U10842 (N_10842,N_5414,N_4231);
or U10843 (N_10843,N_490,N_2496);
nor U10844 (N_10844,N_5720,N_3535);
xor U10845 (N_10845,N_16,N_1087);
and U10846 (N_10846,N_2420,N_1172);
nand U10847 (N_10847,N_3504,N_4592);
nand U10848 (N_10848,N_2668,N_4697);
and U10849 (N_10849,N_2330,N_5906);
or U10850 (N_10850,N_2116,N_1965);
xor U10851 (N_10851,N_5583,N_4002);
and U10852 (N_10852,N_4381,N_796);
xor U10853 (N_10853,N_5159,N_5394);
nand U10854 (N_10854,N_3079,N_5728);
nand U10855 (N_10855,N_455,N_508);
xnor U10856 (N_10856,N_5327,N_3761);
and U10857 (N_10857,N_4931,N_5336);
nor U10858 (N_10858,N_776,N_1213);
xnor U10859 (N_10859,N_4980,N_2127);
and U10860 (N_10860,N_2955,N_2336);
or U10861 (N_10861,N_3748,N_2523);
xnor U10862 (N_10862,N_5980,N_2816);
and U10863 (N_10863,N_2458,N_3482);
xor U10864 (N_10864,N_2161,N_2578);
xor U10865 (N_10865,N_49,N_5595);
nor U10866 (N_10866,N_2722,N_5721);
or U10867 (N_10867,N_230,N_1183);
and U10868 (N_10868,N_3318,N_4802);
xor U10869 (N_10869,N_1829,N_4436);
and U10870 (N_10870,N_4813,N_3979);
or U10871 (N_10871,N_1590,N_4458);
xnor U10872 (N_10872,N_83,N_3460);
xor U10873 (N_10873,N_3248,N_3677);
nor U10874 (N_10874,N_1220,N_2725);
xnor U10875 (N_10875,N_22,N_219);
nand U10876 (N_10876,N_4733,N_5516);
xor U10877 (N_10877,N_3619,N_3409);
or U10878 (N_10878,N_2567,N_1940);
xor U10879 (N_10879,N_3842,N_342);
nand U10880 (N_10880,N_2712,N_3725);
or U10881 (N_10881,N_1549,N_1936);
nand U10882 (N_10882,N_358,N_5465);
and U10883 (N_10883,N_5854,N_4683);
and U10884 (N_10884,N_3451,N_2185);
nand U10885 (N_10885,N_4702,N_3633);
nor U10886 (N_10886,N_4432,N_675);
nor U10887 (N_10887,N_4943,N_1642);
and U10888 (N_10888,N_1266,N_4022);
or U10889 (N_10889,N_1554,N_4362);
nand U10890 (N_10890,N_272,N_4914);
or U10891 (N_10891,N_2400,N_5333);
and U10892 (N_10892,N_5925,N_4603);
nand U10893 (N_10893,N_1277,N_570);
nand U10894 (N_10894,N_850,N_5260);
xnor U10895 (N_10895,N_5284,N_1538);
xnor U10896 (N_10896,N_2619,N_4439);
xnor U10897 (N_10897,N_2226,N_655);
nand U10898 (N_10898,N_1905,N_1447);
nand U10899 (N_10899,N_178,N_3524);
and U10900 (N_10900,N_3321,N_3241);
nor U10901 (N_10901,N_4393,N_3573);
and U10902 (N_10902,N_164,N_1133);
nor U10903 (N_10903,N_2064,N_4438);
and U10904 (N_10904,N_2831,N_4727);
xnor U10905 (N_10905,N_3545,N_3387);
or U10906 (N_10906,N_251,N_1024);
nand U10907 (N_10907,N_1132,N_2991);
xnor U10908 (N_10908,N_2552,N_5682);
nand U10909 (N_10909,N_1057,N_672);
or U10910 (N_10910,N_5925,N_352);
and U10911 (N_10911,N_2333,N_4690);
and U10912 (N_10912,N_5868,N_2385);
or U10913 (N_10913,N_2041,N_2855);
nand U10914 (N_10914,N_5088,N_2234);
nor U10915 (N_10915,N_2086,N_1096);
xnor U10916 (N_10916,N_625,N_3222);
or U10917 (N_10917,N_951,N_1143);
or U10918 (N_10918,N_1392,N_2731);
nor U10919 (N_10919,N_556,N_5601);
xnor U10920 (N_10920,N_4748,N_2870);
nand U10921 (N_10921,N_5088,N_3190);
or U10922 (N_10922,N_207,N_1858);
nor U10923 (N_10923,N_4487,N_5284);
or U10924 (N_10924,N_3047,N_1586);
xor U10925 (N_10925,N_4299,N_3320);
xor U10926 (N_10926,N_243,N_3003);
or U10927 (N_10927,N_4787,N_1279);
nor U10928 (N_10928,N_2451,N_3062);
and U10929 (N_10929,N_3106,N_3834);
and U10930 (N_10930,N_4704,N_3188);
nor U10931 (N_10931,N_27,N_2074);
or U10932 (N_10932,N_3279,N_4002);
xor U10933 (N_10933,N_4889,N_1307);
xnor U10934 (N_10934,N_2028,N_61);
nand U10935 (N_10935,N_2136,N_1757);
xor U10936 (N_10936,N_647,N_3690);
or U10937 (N_10937,N_2964,N_3880);
nor U10938 (N_10938,N_3074,N_4171);
nor U10939 (N_10939,N_5649,N_4492);
or U10940 (N_10940,N_5221,N_1620);
and U10941 (N_10941,N_4879,N_4891);
nand U10942 (N_10942,N_532,N_175);
nor U10943 (N_10943,N_5625,N_2553);
xor U10944 (N_10944,N_4029,N_194);
nor U10945 (N_10945,N_3938,N_170);
and U10946 (N_10946,N_945,N_851);
xnor U10947 (N_10947,N_3850,N_4063);
or U10948 (N_10948,N_1964,N_3020);
or U10949 (N_10949,N_2464,N_5451);
and U10950 (N_10950,N_4212,N_5948);
and U10951 (N_10951,N_3081,N_2143);
and U10952 (N_10952,N_1312,N_2078);
nand U10953 (N_10953,N_3457,N_1404);
xnor U10954 (N_10954,N_579,N_1682);
xnor U10955 (N_10955,N_201,N_1694);
or U10956 (N_10956,N_465,N_5841);
xnor U10957 (N_10957,N_2522,N_165);
xor U10958 (N_10958,N_3588,N_3608);
nand U10959 (N_10959,N_5544,N_5499);
and U10960 (N_10960,N_5743,N_2296);
nor U10961 (N_10961,N_3111,N_4181);
and U10962 (N_10962,N_4512,N_5695);
and U10963 (N_10963,N_4595,N_3699);
or U10964 (N_10964,N_4428,N_4134);
xnor U10965 (N_10965,N_796,N_4444);
nand U10966 (N_10966,N_1713,N_2669);
and U10967 (N_10967,N_1267,N_1120);
nor U10968 (N_10968,N_3845,N_2534);
or U10969 (N_10969,N_4023,N_2157);
and U10970 (N_10970,N_5278,N_2096);
xor U10971 (N_10971,N_2353,N_3213);
nand U10972 (N_10972,N_3417,N_2292);
or U10973 (N_10973,N_855,N_5960);
nand U10974 (N_10974,N_475,N_5332);
nand U10975 (N_10975,N_993,N_5819);
nand U10976 (N_10976,N_1590,N_3983);
or U10977 (N_10977,N_1128,N_3241);
and U10978 (N_10978,N_5441,N_399);
nor U10979 (N_10979,N_2376,N_3784);
or U10980 (N_10980,N_379,N_125);
nor U10981 (N_10981,N_3902,N_3478);
or U10982 (N_10982,N_5477,N_2194);
nand U10983 (N_10983,N_2245,N_439);
or U10984 (N_10984,N_3784,N_1909);
nor U10985 (N_10985,N_2885,N_969);
and U10986 (N_10986,N_7,N_246);
nor U10987 (N_10987,N_2241,N_455);
nand U10988 (N_10988,N_4416,N_456);
nand U10989 (N_10989,N_5883,N_2690);
or U10990 (N_10990,N_4249,N_5270);
xnor U10991 (N_10991,N_3703,N_3412);
and U10992 (N_10992,N_4118,N_4687);
or U10993 (N_10993,N_3735,N_5995);
or U10994 (N_10994,N_4800,N_3388);
and U10995 (N_10995,N_79,N_4998);
and U10996 (N_10996,N_1093,N_5387);
nor U10997 (N_10997,N_5320,N_510);
and U10998 (N_10998,N_1682,N_450);
nand U10999 (N_10999,N_3470,N_5318);
nor U11000 (N_11000,N_5536,N_4645);
nor U11001 (N_11001,N_145,N_5718);
nor U11002 (N_11002,N_2903,N_1801);
nor U11003 (N_11003,N_1867,N_3484);
nor U11004 (N_11004,N_2972,N_3053);
and U11005 (N_11005,N_4225,N_1527);
xor U11006 (N_11006,N_2936,N_2302);
nand U11007 (N_11007,N_3557,N_933);
and U11008 (N_11008,N_705,N_2291);
xor U11009 (N_11009,N_3708,N_4294);
nand U11010 (N_11010,N_2818,N_1422);
and U11011 (N_11011,N_241,N_4797);
nand U11012 (N_11012,N_4568,N_303);
or U11013 (N_11013,N_1284,N_2086);
nor U11014 (N_11014,N_5511,N_1946);
nor U11015 (N_11015,N_4056,N_516);
and U11016 (N_11016,N_5005,N_5964);
nand U11017 (N_11017,N_2456,N_5501);
nor U11018 (N_11018,N_1478,N_310);
nand U11019 (N_11019,N_4221,N_5099);
or U11020 (N_11020,N_1250,N_5631);
or U11021 (N_11021,N_4438,N_3006);
xnor U11022 (N_11022,N_1741,N_754);
xnor U11023 (N_11023,N_1895,N_3276);
and U11024 (N_11024,N_3870,N_4995);
xor U11025 (N_11025,N_824,N_423);
nor U11026 (N_11026,N_1893,N_2898);
and U11027 (N_11027,N_4592,N_5226);
and U11028 (N_11028,N_5479,N_2405);
and U11029 (N_11029,N_1515,N_1922);
nor U11030 (N_11030,N_5860,N_4631);
nor U11031 (N_11031,N_5634,N_3887);
nor U11032 (N_11032,N_5822,N_1188);
nor U11033 (N_11033,N_1537,N_2741);
xnor U11034 (N_11034,N_916,N_4830);
nand U11035 (N_11035,N_3286,N_4592);
and U11036 (N_11036,N_3675,N_5262);
nand U11037 (N_11037,N_394,N_850);
nand U11038 (N_11038,N_5510,N_4146);
nor U11039 (N_11039,N_2576,N_3100);
or U11040 (N_11040,N_2731,N_4841);
nor U11041 (N_11041,N_3367,N_2941);
nor U11042 (N_11042,N_495,N_49);
xor U11043 (N_11043,N_621,N_4191);
xnor U11044 (N_11044,N_4586,N_2390);
and U11045 (N_11045,N_4045,N_2711);
nand U11046 (N_11046,N_1713,N_5184);
nand U11047 (N_11047,N_1963,N_3871);
nor U11048 (N_11048,N_4858,N_3646);
nor U11049 (N_11049,N_1845,N_5376);
and U11050 (N_11050,N_3393,N_2803);
nor U11051 (N_11051,N_1920,N_2120);
or U11052 (N_11052,N_1830,N_4345);
xor U11053 (N_11053,N_5875,N_5062);
xor U11054 (N_11054,N_1152,N_103);
nor U11055 (N_11055,N_4938,N_2331);
or U11056 (N_11056,N_936,N_1291);
xnor U11057 (N_11057,N_2367,N_4839);
and U11058 (N_11058,N_2992,N_5680);
and U11059 (N_11059,N_3207,N_4723);
and U11060 (N_11060,N_423,N_542);
or U11061 (N_11061,N_3264,N_949);
and U11062 (N_11062,N_3445,N_1335);
xor U11063 (N_11063,N_4990,N_952);
xnor U11064 (N_11064,N_3683,N_1298);
nor U11065 (N_11065,N_3584,N_295);
and U11066 (N_11066,N_2199,N_1524);
nor U11067 (N_11067,N_5103,N_876);
nand U11068 (N_11068,N_5458,N_3242);
and U11069 (N_11069,N_2964,N_2433);
nor U11070 (N_11070,N_369,N_4192);
and U11071 (N_11071,N_5256,N_5372);
and U11072 (N_11072,N_5672,N_3044);
xor U11073 (N_11073,N_4559,N_1921);
or U11074 (N_11074,N_2799,N_3636);
and U11075 (N_11075,N_2789,N_5571);
nor U11076 (N_11076,N_353,N_1337);
and U11077 (N_11077,N_2172,N_1011);
xor U11078 (N_11078,N_5724,N_3781);
nand U11079 (N_11079,N_3675,N_4391);
nand U11080 (N_11080,N_1169,N_4661);
and U11081 (N_11081,N_3917,N_4423);
or U11082 (N_11082,N_4059,N_937);
nand U11083 (N_11083,N_5324,N_325);
nand U11084 (N_11084,N_3758,N_416);
nand U11085 (N_11085,N_3459,N_4696);
xnor U11086 (N_11086,N_2747,N_1219);
or U11087 (N_11087,N_5724,N_1288);
and U11088 (N_11088,N_3894,N_5322);
nand U11089 (N_11089,N_3372,N_2610);
or U11090 (N_11090,N_3551,N_414);
xnor U11091 (N_11091,N_4111,N_3546);
xor U11092 (N_11092,N_2783,N_4195);
and U11093 (N_11093,N_2611,N_1971);
or U11094 (N_11094,N_5389,N_4976);
xnor U11095 (N_11095,N_5712,N_3834);
nor U11096 (N_11096,N_576,N_5809);
or U11097 (N_11097,N_540,N_1498);
xor U11098 (N_11098,N_1034,N_277);
nand U11099 (N_11099,N_2854,N_2546);
and U11100 (N_11100,N_1450,N_5011);
nor U11101 (N_11101,N_3747,N_3839);
or U11102 (N_11102,N_195,N_3979);
nor U11103 (N_11103,N_733,N_3096);
nor U11104 (N_11104,N_3253,N_5533);
nand U11105 (N_11105,N_712,N_5315);
or U11106 (N_11106,N_4009,N_4338);
or U11107 (N_11107,N_1819,N_2689);
xnor U11108 (N_11108,N_4572,N_3795);
xor U11109 (N_11109,N_1442,N_2376);
nand U11110 (N_11110,N_5061,N_2723);
or U11111 (N_11111,N_3017,N_2566);
nand U11112 (N_11112,N_3112,N_5829);
nor U11113 (N_11113,N_3149,N_1107);
xnor U11114 (N_11114,N_330,N_3144);
or U11115 (N_11115,N_1112,N_3505);
nand U11116 (N_11116,N_2256,N_2059);
nor U11117 (N_11117,N_5974,N_2772);
nor U11118 (N_11118,N_2746,N_3706);
nand U11119 (N_11119,N_5987,N_5332);
nand U11120 (N_11120,N_305,N_2005);
nor U11121 (N_11121,N_3936,N_3299);
xor U11122 (N_11122,N_2333,N_4506);
or U11123 (N_11123,N_669,N_4513);
and U11124 (N_11124,N_2574,N_2661);
xor U11125 (N_11125,N_3988,N_5590);
or U11126 (N_11126,N_807,N_2177);
nor U11127 (N_11127,N_3594,N_4244);
and U11128 (N_11128,N_3125,N_2784);
nand U11129 (N_11129,N_5239,N_2867);
nor U11130 (N_11130,N_5231,N_3756);
xnor U11131 (N_11131,N_4969,N_57);
or U11132 (N_11132,N_2045,N_4598);
or U11133 (N_11133,N_1192,N_2050);
or U11134 (N_11134,N_5934,N_840);
nand U11135 (N_11135,N_1131,N_2953);
nor U11136 (N_11136,N_1630,N_4854);
or U11137 (N_11137,N_1950,N_1669);
xnor U11138 (N_11138,N_2436,N_281);
and U11139 (N_11139,N_4290,N_1467);
or U11140 (N_11140,N_2664,N_1867);
nor U11141 (N_11141,N_5961,N_5525);
or U11142 (N_11142,N_3868,N_5805);
nor U11143 (N_11143,N_4656,N_4460);
or U11144 (N_11144,N_1776,N_4057);
nor U11145 (N_11145,N_205,N_2546);
xor U11146 (N_11146,N_3083,N_3469);
and U11147 (N_11147,N_2666,N_1913);
nor U11148 (N_11148,N_4131,N_1485);
nand U11149 (N_11149,N_464,N_5540);
nor U11150 (N_11150,N_526,N_2980);
nand U11151 (N_11151,N_1348,N_1728);
nor U11152 (N_11152,N_2664,N_5058);
nand U11153 (N_11153,N_5632,N_3521);
and U11154 (N_11154,N_4985,N_2904);
xor U11155 (N_11155,N_396,N_5273);
nor U11156 (N_11156,N_2552,N_1587);
or U11157 (N_11157,N_983,N_3842);
and U11158 (N_11158,N_3277,N_149);
and U11159 (N_11159,N_2663,N_5494);
nor U11160 (N_11160,N_579,N_877);
and U11161 (N_11161,N_274,N_5838);
and U11162 (N_11162,N_1945,N_1162);
and U11163 (N_11163,N_3524,N_2289);
xnor U11164 (N_11164,N_3018,N_5804);
and U11165 (N_11165,N_3453,N_809);
nor U11166 (N_11166,N_3655,N_4267);
nor U11167 (N_11167,N_3343,N_5544);
nand U11168 (N_11168,N_5877,N_5787);
nor U11169 (N_11169,N_2246,N_3100);
xor U11170 (N_11170,N_4727,N_4620);
or U11171 (N_11171,N_1269,N_961);
nand U11172 (N_11172,N_5609,N_723);
nor U11173 (N_11173,N_306,N_125);
nor U11174 (N_11174,N_3877,N_3917);
xnor U11175 (N_11175,N_5142,N_3421);
or U11176 (N_11176,N_4548,N_4810);
or U11177 (N_11177,N_4526,N_3170);
nor U11178 (N_11178,N_4648,N_4994);
or U11179 (N_11179,N_2957,N_5397);
or U11180 (N_11180,N_2263,N_724);
nor U11181 (N_11181,N_2497,N_5119);
nor U11182 (N_11182,N_3776,N_4998);
nand U11183 (N_11183,N_5277,N_4532);
and U11184 (N_11184,N_480,N_2565);
nor U11185 (N_11185,N_5799,N_4192);
xor U11186 (N_11186,N_606,N_262);
or U11187 (N_11187,N_1311,N_5768);
or U11188 (N_11188,N_3818,N_3778);
nor U11189 (N_11189,N_5556,N_5186);
nor U11190 (N_11190,N_3538,N_3068);
nor U11191 (N_11191,N_5656,N_3994);
nand U11192 (N_11192,N_5989,N_3513);
nand U11193 (N_11193,N_5573,N_3473);
and U11194 (N_11194,N_244,N_1647);
xnor U11195 (N_11195,N_319,N_297);
and U11196 (N_11196,N_78,N_519);
nand U11197 (N_11197,N_2167,N_2725);
and U11198 (N_11198,N_3359,N_3672);
and U11199 (N_11199,N_4279,N_3617);
nor U11200 (N_11200,N_2092,N_4833);
nand U11201 (N_11201,N_2967,N_3861);
and U11202 (N_11202,N_4737,N_5202);
or U11203 (N_11203,N_2007,N_1264);
or U11204 (N_11204,N_1738,N_1771);
nor U11205 (N_11205,N_3315,N_198);
nand U11206 (N_11206,N_1255,N_2856);
nand U11207 (N_11207,N_5112,N_589);
and U11208 (N_11208,N_2631,N_2889);
nor U11209 (N_11209,N_991,N_4568);
nor U11210 (N_11210,N_4536,N_4447);
xnor U11211 (N_11211,N_4913,N_4210);
and U11212 (N_11212,N_5279,N_4987);
xnor U11213 (N_11213,N_3154,N_706);
xor U11214 (N_11214,N_2613,N_28);
nor U11215 (N_11215,N_572,N_5302);
nand U11216 (N_11216,N_1504,N_4832);
xnor U11217 (N_11217,N_2447,N_707);
nor U11218 (N_11218,N_1901,N_4684);
or U11219 (N_11219,N_1438,N_3502);
or U11220 (N_11220,N_2239,N_5663);
and U11221 (N_11221,N_1352,N_2463);
nand U11222 (N_11222,N_5516,N_4646);
or U11223 (N_11223,N_3749,N_4303);
or U11224 (N_11224,N_4407,N_136);
or U11225 (N_11225,N_4601,N_3508);
nand U11226 (N_11226,N_2635,N_4747);
xor U11227 (N_11227,N_5741,N_410);
and U11228 (N_11228,N_978,N_5295);
and U11229 (N_11229,N_2397,N_1554);
nand U11230 (N_11230,N_3624,N_4075);
nor U11231 (N_11231,N_4188,N_1517);
nand U11232 (N_11232,N_4718,N_1292);
and U11233 (N_11233,N_4431,N_1616);
and U11234 (N_11234,N_4578,N_498);
nand U11235 (N_11235,N_1080,N_4961);
nand U11236 (N_11236,N_0,N_1027);
xor U11237 (N_11237,N_3188,N_5544);
and U11238 (N_11238,N_2821,N_4149);
or U11239 (N_11239,N_5840,N_811);
nor U11240 (N_11240,N_4625,N_3843);
xnor U11241 (N_11241,N_2237,N_4371);
nand U11242 (N_11242,N_2540,N_2203);
nand U11243 (N_11243,N_2253,N_5510);
or U11244 (N_11244,N_3822,N_365);
xor U11245 (N_11245,N_3663,N_2565);
xor U11246 (N_11246,N_3181,N_5943);
nor U11247 (N_11247,N_1454,N_1050);
and U11248 (N_11248,N_339,N_4258);
nor U11249 (N_11249,N_992,N_3773);
nand U11250 (N_11250,N_1449,N_3446);
nor U11251 (N_11251,N_4065,N_3931);
xnor U11252 (N_11252,N_4808,N_1099);
nor U11253 (N_11253,N_1409,N_3863);
or U11254 (N_11254,N_36,N_715);
xnor U11255 (N_11255,N_3663,N_2511);
and U11256 (N_11256,N_4226,N_1459);
nand U11257 (N_11257,N_2771,N_2037);
xnor U11258 (N_11258,N_1620,N_3688);
and U11259 (N_11259,N_2734,N_1265);
or U11260 (N_11260,N_5253,N_1802);
nor U11261 (N_11261,N_1735,N_4633);
or U11262 (N_11262,N_4742,N_1517);
nor U11263 (N_11263,N_4262,N_517);
and U11264 (N_11264,N_3769,N_4700);
xnor U11265 (N_11265,N_3733,N_3724);
nand U11266 (N_11266,N_5900,N_2623);
nand U11267 (N_11267,N_5044,N_3523);
and U11268 (N_11268,N_3717,N_169);
nor U11269 (N_11269,N_5068,N_3174);
xnor U11270 (N_11270,N_688,N_5119);
nor U11271 (N_11271,N_2594,N_2226);
and U11272 (N_11272,N_2368,N_5533);
nor U11273 (N_11273,N_850,N_5876);
and U11274 (N_11274,N_3569,N_4184);
and U11275 (N_11275,N_2070,N_235);
xor U11276 (N_11276,N_2929,N_4109);
or U11277 (N_11277,N_5255,N_1396);
nand U11278 (N_11278,N_5974,N_2149);
or U11279 (N_11279,N_4032,N_1345);
nor U11280 (N_11280,N_4646,N_3354);
or U11281 (N_11281,N_1539,N_3818);
or U11282 (N_11282,N_593,N_2985);
nor U11283 (N_11283,N_629,N_15);
nand U11284 (N_11284,N_5709,N_1206);
nor U11285 (N_11285,N_2347,N_2718);
xnor U11286 (N_11286,N_4909,N_3671);
or U11287 (N_11287,N_4948,N_325);
nand U11288 (N_11288,N_3967,N_794);
or U11289 (N_11289,N_2584,N_2169);
or U11290 (N_11290,N_2344,N_2982);
and U11291 (N_11291,N_4841,N_3184);
nand U11292 (N_11292,N_2241,N_4535);
and U11293 (N_11293,N_4129,N_1824);
nand U11294 (N_11294,N_2726,N_630);
nand U11295 (N_11295,N_3160,N_2060);
or U11296 (N_11296,N_3176,N_4366);
or U11297 (N_11297,N_5925,N_619);
nor U11298 (N_11298,N_271,N_4028);
nor U11299 (N_11299,N_311,N_4813);
or U11300 (N_11300,N_2743,N_4689);
or U11301 (N_11301,N_2515,N_4051);
nor U11302 (N_11302,N_3292,N_2943);
nor U11303 (N_11303,N_1702,N_1502);
nor U11304 (N_11304,N_2123,N_4460);
nand U11305 (N_11305,N_2016,N_4299);
or U11306 (N_11306,N_170,N_1120);
xor U11307 (N_11307,N_4167,N_3278);
nand U11308 (N_11308,N_2559,N_3662);
and U11309 (N_11309,N_5580,N_4218);
xnor U11310 (N_11310,N_115,N_462);
nor U11311 (N_11311,N_11,N_2732);
xnor U11312 (N_11312,N_5694,N_241);
or U11313 (N_11313,N_3349,N_3687);
and U11314 (N_11314,N_2426,N_2990);
nor U11315 (N_11315,N_652,N_1922);
nor U11316 (N_11316,N_5832,N_5774);
and U11317 (N_11317,N_5481,N_4272);
nor U11318 (N_11318,N_5667,N_1655);
xor U11319 (N_11319,N_3639,N_5802);
nor U11320 (N_11320,N_2059,N_270);
and U11321 (N_11321,N_5463,N_2479);
xor U11322 (N_11322,N_182,N_790);
or U11323 (N_11323,N_4138,N_3548);
nand U11324 (N_11324,N_5662,N_2733);
xor U11325 (N_11325,N_1574,N_3002);
nor U11326 (N_11326,N_504,N_1676);
nor U11327 (N_11327,N_3866,N_4145);
or U11328 (N_11328,N_4223,N_3755);
nor U11329 (N_11329,N_5678,N_136);
nor U11330 (N_11330,N_4412,N_3879);
nand U11331 (N_11331,N_4139,N_2309);
or U11332 (N_11332,N_2986,N_2198);
nor U11333 (N_11333,N_415,N_5904);
and U11334 (N_11334,N_4536,N_4341);
and U11335 (N_11335,N_4344,N_4121);
or U11336 (N_11336,N_5740,N_2215);
nor U11337 (N_11337,N_676,N_5829);
and U11338 (N_11338,N_3676,N_66);
and U11339 (N_11339,N_4621,N_1867);
nand U11340 (N_11340,N_3552,N_2968);
nand U11341 (N_11341,N_508,N_2779);
nor U11342 (N_11342,N_1817,N_938);
xor U11343 (N_11343,N_2984,N_3796);
and U11344 (N_11344,N_150,N_1625);
xnor U11345 (N_11345,N_3314,N_1631);
nand U11346 (N_11346,N_3820,N_5979);
nor U11347 (N_11347,N_1064,N_2093);
and U11348 (N_11348,N_3727,N_5713);
or U11349 (N_11349,N_586,N_3952);
or U11350 (N_11350,N_1684,N_4208);
nand U11351 (N_11351,N_1277,N_5227);
nor U11352 (N_11352,N_4713,N_3885);
or U11353 (N_11353,N_5479,N_1755);
nand U11354 (N_11354,N_1105,N_1998);
nand U11355 (N_11355,N_5265,N_2540);
and U11356 (N_11356,N_1955,N_5178);
or U11357 (N_11357,N_4935,N_2430);
and U11358 (N_11358,N_1591,N_750);
xor U11359 (N_11359,N_459,N_5980);
or U11360 (N_11360,N_3768,N_5361);
nand U11361 (N_11361,N_4766,N_4474);
xnor U11362 (N_11362,N_4039,N_4916);
or U11363 (N_11363,N_4669,N_4951);
nor U11364 (N_11364,N_5110,N_1912);
nand U11365 (N_11365,N_2015,N_1824);
or U11366 (N_11366,N_4206,N_1586);
xnor U11367 (N_11367,N_4349,N_3120);
and U11368 (N_11368,N_2908,N_1154);
nor U11369 (N_11369,N_5762,N_3185);
nor U11370 (N_11370,N_5527,N_20);
nand U11371 (N_11371,N_1320,N_3773);
xor U11372 (N_11372,N_2107,N_2178);
xor U11373 (N_11373,N_2167,N_4883);
nor U11374 (N_11374,N_951,N_3648);
or U11375 (N_11375,N_4635,N_1949);
or U11376 (N_11376,N_1384,N_770);
or U11377 (N_11377,N_4881,N_1212);
or U11378 (N_11378,N_775,N_43);
nand U11379 (N_11379,N_5775,N_745);
or U11380 (N_11380,N_659,N_1823);
nand U11381 (N_11381,N_2969,N_3886);
nand U11382 (N_11382,N_5519,N_430);
xor U11383 (N_11383,N_2463,N_5377);
or U11384 (N_11384,N_1093,N_5417);
xor U11385 (N_11385,N_4226,N_2289);
xnor U11386 (N_11386,N_1115,N_2360);
or U11387 (N_11387,N_5086,N_3064);
or U11388 (N_11388,N_5863,N_4586);
nand U11389 (N_11389,N_4917,N_1546);
or U11390 (N_11390,N_246,N_4807);
or U11391 (N_11391,N_1174,N_5303);
nand U11392 (N_11392,N_3083,N_1704);
and U11393 (N_11393,N_1405,N_1261);
nand U11394 (N_11394,N_523,N_632);
or U11395 (N_11395,N_2052,N_5135);
or U11396 (N_11396,N_2697,N_3190);
nand U11397 (N_11397,N_1742,N_597);
or U11398 (N_11398,N_3353,N_373);
and U11399 (N_11399,N_5296,N_753);
or U11400 (N_11400,N_3327,N_5457);
and U11401 (N_11401,N_301,N_1537);
nor U11402 (N_11402,N_1178,N_5471);
and U11403 (N_11403,N_4352,N_1252);
or U11404 (N_11404,N_2497,N_5306);
xnor U11405 (N_11405,N_1784,N_4131);
nand U11406 (N_11406,N_1344,N_3916);
nand U11407 (N_11407,N_2598,N_5236);
and U11408 (N_11408,N_942,N_450);
or U11409 (N_11409,N_3397,N_543);
nor U11410 (N_11410,N_1096,N_4489);
or U11411 (N_11411,N_905,N_4796);
xor U11412 (N_11412,N_2528,N_1014);
nand U11413 (N_11413,N_1595,N_463);
or U11414 (N_11414,N_4494,N_1452);
xor U11415 (N_11415,N_2103,N_3672);
xnor U11416 (N_11416,N_127,N_1857);
nand U11417 (N_11417,N_991,N_1584);
nor U11418 (N_11418,N_2397,N_2350);
xnor U11419 (N_11419,N_1275,N_3236);
nand U11420 (N_11420,N_1480,N_4392);
and U11421 (N_11421,N_5372,N_5388);
or U11422 (N_11422,N_2570,N_47);
or U11423 (N_11423,N_1792,N_5801);
xor U11424 (N_11424,N_5713,N_3736);
and U11425 (N_11425,N_395,N_4386);
nand U11426 (N_11426,N_1220,N_3745);
and U11427 (N_11427,N_5749,N_4634);
and U11428 (N_11428,N_3471,N_4756);
and U11429 (N_11429,N_3148,N_4486);
xor U11430 (N_11430,N_2027,N_2208);
nor U11431 (N_11431,N_2343,N_4041);
nand U11432 (N_11432,N_1824,N_1316);
nand U11433 (N_11433,N_3531,N_4133);
and U11434 (N_11434,N_2797,N_3201);
nand U11435 (N_11435,N_627,N_470);
nor U11436 (N_11436,N_4919,N_2324);
nand U11437 (N_11437,N_2384,N_5993);
nor U11438 (N_11438,N_807,N_2873);
or U11439 (N_11439,N_2970,N_4647);
nor U11440 (N_11440,N_1255,N_5148);
xnor U11441 (N_11441,N_2402,N_2043);
xnor U11442 (N_11442,N_5852,N_806);
or U11443 (N_11443,N_5768,N_3497);
and U11444 (N_11444,N_977,N_2218);
nand U11445 (N_11445,N_4594,N_2016);
or U11446 (N_11446,N_2481,N_2823);
xnor U11447 (N_11447,N_312,N_424);
and U11448 (N_11448,N_3759,N_4133);
nand U11449 (N_11449,N_829,N_1061);
nand U11450 (N_11450,N_1849,N_5418);
and U11451 (N_11451,N_2470,N_3208);
and U11452 (N_11452,N_4785,N_1915);
and U11453 (N_11453,N_942,N_5339);
or U11454 (N_11454,N_5022,N_1261);
nor U11455 (N_11455,N_5289,N_1000);
or U11456 (N_11456,N_681,N_1553);
or U11457 (N_11457,N_2488,N_893);
nand U11458 (N_11458,N_736,N_5975);
nor U11459 (N_11459,N_2101,N_224);
nand U11460 (N_11460,N_3778,N_5032);
and U11461 (N_11461,N_5031,N_1540);
and U11462 (N_11462,N_5337,N_2059);
or U11463 (N_11463,N_606,N_4724);
and U11464 (N_11464,N_3073,N_2761);
nand U11465 (N_11465,N_2579,N_3330);
nand U11466 (N_11466,N_4123,N_5136);
and U11467 (N_11467,N_1973,N_5361);
nand U11468 (N_11468,N_5303,N_1782);
and U11469 (N_11469,N_719,N_1861);
xor U11470 (N_11470,N_5144,N_1248);
xor U11471 (N_11471,N_5928,N_5948);
nor U11472 (N_11472,N_2956,N_5825);
nor U11473 (N_11473,N_4475,N_4272);
and U11474 (N_11474,N_4542,N_4418);
and U11475 (N_11475,N_2739,N_3144);
nand U11476 (N_11476,N_952,N_2090);
or U11477 (N_11477,N_5148,N_5153);
xnor U11478 (N_11478,N_4493,N_401);
and U11479 (N_11479,N_2622,N_5073);
or U11480 (N_11480,N_283,N_4877);
nand U11481 (N_11481,N_4981,N_1570);
nor U11482 (N_11482,N_5495,N_5757);
or U11483 (N_11483,N_5645,N_3057);
nand U11484 (N_11484,N_593,N_1360);
nor U11485 (N_11485,N_1190,N_756);
and U11486 (N_11486,N_4392,N_3233);
xor U11487 (N_11487,N_4535,N_5013);
nand U11488 (N_11488,N_3785,N_356);
and U11489 (N_11489,N_3466,N_851);
xor U11490 (N_11490,N_816,N_2825);
or U11491 (N_11491,N_5577,N_4559);
and U11492 (N_11492,N_1369,N_2127);
nor U11493 (N_11493,N_2550,N_2259);
nand U11494 (N_11494,N_5740,N_4575);
nand U11495 (N_11495,N_3602,N_2601);
nor U11496 (N_11496,N_4272,N_5715);
and U11497 (N_11497,N_5508,N_5104);
nor U11498 (N_11498,N_4335,N_4736);
nor U11499 (N_11499,N_4861,N_2764);
nor U11500 (N_11500,N_18,N_4883);
or U11501 (N_11501,N_1735,N_2224);
and U11502 (N_11502,N_2762,N_2232);
or U11503 (N_11503,N_1656,N_3280);
nor U11504 (N_11504,N_5577,N_3751);
xnor U11505 (N_11505,N_2705,N_3495);
and U11506 (N_11506,N_575,N_1518);
nand U11507 (N_11507,N_5812,N_5461);
xor U11508 (N_11508,N_1721,N_2560);
or U11509 (N_11509,N_3825,N_5918);
nor U11510 (N_11510,N_174,N_3119);
nand U11511 (N_11511,N_5796,N_3720);
xor U11512 (N_11512,N_5071,N_3675);
or U11513 (N_11513,N_3096,N_2277);
nor U11514 (N_11514,N_3614,N_2429);
and U11515 (N_11515,N_1069,N_3693);
or U11516 (N_11516,N_4114,N_434);
and U11517 (N_11517,N_2659,N_5756);
nor U11518 (N_11518,N_3383,N_1061);
nor U11519 (N_11519,N_1248,N_183);
and U11520 (N_11520,N_35,N_2385);
nand U11521 (N_11521,N_4735,N_4452);
nand U11522 (N_11522,N_2867,N_3773);
and U11523 (N_11523,N_5040,N_5138);
nor U11524 (N_11524,N_2062,N_2464);
or U11525 (N_11525,N_3503,N_32);
nor U11526 (N_11526,N_1492,N_1054);
xor U11527 (N_11527,N_4813,N_5585);
xnor U11528 (N_11528,N_5802,N_2013);
xor U11529 (N_11529,N_2483,N_2424);
and U11530 (N_11530,N_2753,N_3283);
nand U11531 (N_11531,N_1764,N_4676);
and U11532 (N_11532,N_694,N_5729);
nor U11533 (N_11533,N_4852,N_1221);
nand U11534 (N_11534,N_372,N_5700);
nor U11535 (N_11535,N_3901,N_156);
xor U11536 (N_11536,N_2745,N_4106);
nor U11537 (N_11537,N_5693,N_1168);
and U11538 (N_11538,N_2416,N_3462);
nor U11539 (N_11539,N_2473,N_4324);
and U11540 (N_11540,N_4982,N_4770);
xnor U11541 (N_11541,N_4244,N_4701);
xnor U11542 (N_11542,N_3933,N_3009);
nand U11543 (N_11543,N_1793,N_3817);
and U11544 (N_11544,N_235,N_1868);
nand U11545 (N_11545,N_5047,N_1478);
xnor U11546 (N_11546,N_5774,N_5158);
xnor U11547 (N_11547,N_5460,N_1463);
xnor U11548 (N_11548,N_4214,N_279);
or U11549 (N_11549,N_3353,N_2962);
nor U11550 (N_11550,N_4512,N_5775);
and U11551 (N_11551,N_5764,N_2526);
or U11552 (N_11552,N_1944,N_2155);
nand U11553 (N_11553,N_1194,N_385);
and U11554 (N_11554,N_3752,N_4274);
and U11555 (N_11555,N_607,N_4151);
or U11556 (N_11556,N_4503,N_2426);
and U11557 (N_11557,N_1410,N_1195);
nor U11558 (N_11558,N_1864,N_2122);
nor U11559 (N_11559,N_4702,N_5322);
nand U11560 (N_11560,N_3263,N_736);
and U11561 (N_11561,N_5442,N_854);
or U11562 (N_11562,N_1827,N_5401);
or U11563 (N_11563,N_3873,N_3114);
nand U11564 (N_11564,N_5589,N_619);
xnor U11565 (N_11565,N_1623,N_4563);
xor U11566 (N_11566,N_3889,N_2961);
and U11567 (N_11567,N_3406,N_4587);
xor U11568 (N_11568,N_75,N_5601);
xor U11569 (N_11569,N_4845,N_1104);
xor U11570 (N_11570,N_900,N_1216);
and U11571 (N_11571,N_172,N_5256);
and U11572 (N_11572,N_4451,N_4380);
and U11573 (N_11573,N_3541,N_5499);
and U11574 (N_11574,N_3462,N_220);
or U11575 (N_11575,N_4776,N_3478);
nor U11576 (N_11576,N_2108,N_151);
nand U11577 (N_11577,N_3035,N_4651);
nand U11578 (N_11578,N_2926,N_1480);
and U11579 (N_11579,N_5699,N_1979);
xnor U11580 (N_11580,N_4618,N_1248);
nand U11581 (N_11581,N_2350,N_1283);
nand U11582 (N_11582,N_2075,N_3967);
or U11583 (N_11583,N_5873,N_3635);
and U11584 (N_11584,N_2509,N_2090);
and U11585 (N_11585,N_4950,N_5941);
nor U11586 (N_11586,N_774,N_3585);
and U11587 (N_11587,N_4754,N_1835);
or U11588 (N_11588,N_2870,N_4296);
xor U11589 (N_11589,N_4888,N_3672);
nor U11590 (N_11590,N_5844,N_1170);
and U11591 (N_11591,N_4310,N_4125);
and U11592 (N_11592,N_4944,N_2165);
or U11593 (N_11593,N_5566,N_410);
nor U11594 (N_11594,N_4418,N_3560);
nor U11595 (N_11595,N_4519,N_3446);
nand U11596 (N_11596,N_3246,N_5591);
and U11597 (N_11597,N_1441,N_640);
or U11598 (N_11598,N_992,N_2218);
or U11599 (N_11599,N_210,N_4317);
nor U11600 (N_11600,N_1688,N_3997);
and U11601 (N_11601,N_4809,N_5282);
and U11602 (N_11602,N_3514,N_4454);
nand U11603 (N_11603,N_5762,N_5854);
nand U11604 (N_11604,N_2983,N_4778);
or U11605 (N_11605,N_3785,N_1810);
nand U11606 (N_11606,N_4883,N_1016);
xor U11607 (N_11607,N_2085,N_785);
and U11608 (N_11608,N_5533,N_2233);
nor U11609 (N_11609,N_295,N_96);
xor U11610 (N_11610,N_4712,N_1913);
xnor U11611 (N_11611,N_81,N_5227);
or U11612 (N_11612,N_4479,N_2724);
nor U11613 (N_11613,N_2027,N_3300);
nor U11614 (N_11614,N_3566,N_5789);
or U11615 (N_11615,N_2038,N_5894);
nor U11616 (N_11616,N_2387,N_1289);
and U11617 (N_11617,N_904,N_4719);
nand U11618 (N_11618,N_1107,N_922);
nor U11619 (N_11619,N_3767,N_584);
xnor U11620 (N_11620,N_2893,N_3843);
and U11621 (N_11621,N_4180,N_466);
and U11622 (N_11622,N_5234,N_686);
or U11623 (N_11623,N_1180,N_1617);
nand U11624 (N_11624,N_4445,N_3516);
or U11625 (N_11625,N_3959,N_91);
and U11626 (N_11626,N_3732,N_4189);
xor U11627 (N_11627,N_5876,N_4560);
or U11628 (N_11628,N_4621,N_5221);
and U11629 (N_11629,N_48,N_660);
and U11630 (N_11630,N_983,N_2907);
or U11631 (N_11631,N_3139,N_4170);
or U11632 (N_11632,N_2749,N_4831);
and U11633 (N_11633,N_5057,N_5392);
xor U11634 (N_11634,N_4463,N_4830);
nor U11635 (N_11635,N_3335,N_3473);
or U11636 (N_11636,N_5521,N_1804);
nor U11637 (N_11637,N_2387,N_3423);
or U11638 (N_11638,N_3288,N_4254);
nand U11639 (N_11639,N_3388,N_2600);
nor U11640 (N_11640,N_4123,N_3165);
or U11641 (N_11641,N_2118,N_1459);
or U11642 (N_11642,N_1167,N_5361);
xnor U11643 (N_11643,N_3876,N_2564);
xnor U11644 (N_11644,N_2167,N_5933);
nor U11645 (N_11645,N_1770,N_739);
nor U11646 (N_11646,N_547,N_5713);
or U11647 (N_11647,N_3019,N_336);
nand U11648 (N_11648,N_252,N_5718);
and U11649 (N_11649,N_5573,N_1893);
and U11650 (N_11650,N_4053,N_5091);
and U11651 (N_11651,N_139,N_1232);
or U11652 (N_11652,N_2978,N_3300);
xor U11653 (N_11653,N_1557,N_5966);
and U11654 (N_11654,N_962,N_3635);
and U11655 (N_11655,N_997,N_2621);
nand U11656 (N_11656,N_1611,N_1835);
nand U11657 (N_11657,N_3476,N_5007);
or U11658 (N_11658,N_1011,N_4446);
nor U11659 (N_11659,N_1411,N_4060);
and U11660 (N_11660,N_348,N_2701);
nand U11661 (N_11661,N_4050,N_3848);
nand U11662 (N_11662,N_1440,N_5788);
or U11663 (N_11663,N_5822,N_5306);
nand U11664 (N_11664,N_3389,N_3602);
nor U11665 (N_11665,N_1406,N_1750);
nor U11666 (N_11666,N_4097,N_5710);
or U11667 (N_11667,N_3447,N_3754);
or U11668 (N_11668,N_1371,N_5266);
xnor U11669 (N_11669,N_4070,N_5199);
xor U11670 (N_11670,N_3931,N_5492);
xnor U11671 (N_11671,N_2036,N_2272);
nand U11672 (N_11672,N_3771,N_786);
or U11673 (N_11673,N_596,N_5831);
nand U11674 (N_11674,N_4244,N_357);
nor U11675 (N_11675,N_4174,N_2220);
and U11676 (N_11676,N_5738,N_2786);
nand U11677 (N_11677,N_4953,N_237);
nor U11678 (N_11678,N_5651,N_96);
xor U11679 (N_11679,N_4708,N_76);
nor U11680 (N_11680,N_363,N_527);
nand U11681 (N_11681,N_1866,N_5792);
nor U11682 (N_11682,N_5218,N_5515);
xor U11683 (N_11683,N_2544,N_4407);
nand U11684 (N_11684,N_1317,N_3927);
nor U11685 (N_11685,N_4530,N_5380);
nor U11686 (N_11686,N_4406,N_5617);
and U11687 (N_11687,N_307,N_826);
or U11688 (N_11688,N_2091,N_1413);
or U11689 (N_11689,N_5629,N_3811);
xor U11690 (N_11690,N_474,N_2470);
and U11691 (N_11691,N_1674,N_3428);
xor U11692 (N_11692,N_5287,N_3078);
and U11693 (N_11693,N_2299,N_309);
and U11694 (N_11694,N_1824,N_604);
or U11695 (N_11695,N_2963,N_806);
nand U11696 (N_11696,N_992,N_1451);
nand U11697 (N_11697,N_2169,N_4393);
and U11698 (N_11698,N_3389,N_2892);
and U11699 (N_11699,N_3264,N_243);
nand U11700 (N_11700,N_2349,N_4547);
nand U11701 (N_11701,N_1405,N_3146);
nor U11702 (N_11702,N_5610,N_1249);
xnor U11703 (N_11703,N_5131,N_3710);
nand U11704 (N_11704,N_5097,N_4949);
or U11705 (N_11705,N_2700,N_3604);
nor U11706 (N_11706,N_325,N_5753);
and U11707 (N_11707,N_3049,N_469);
xnor U11708 (N_11708,N_173,N_4353);
xor U11709 (N_11709,N_674,N_4363);
nand U11710 (N_11710,N_5326,N_977);
nand U11711 (N_11711,N_1576,N_2814);
or U11712 (N_11712,N_5961,N_2809);
and U11713 (N_11713,N_2817,N_5784);
xnor U11714 (N_11714,N_3184,N_3603);
nor U11715 (N_11715,N_1587,N_5329);
or U11716 (N_11716,N_2487,N_2319);
or U11717 (N_11717,N_5126,N_2683);
or U11718 (N_11718,N_356,N_2075);
or U11719 (N_11719,N_5250,N_3203);
nor U11720 (N_11720,N_5665,N_2920);
or U11721 (N_11721,N_3914,N_240);
and U11722 (N_11722,N_203,N_1702);
and U11723 (N_11723,N_834,N_5715);
nand U11724 (N_11724,N_2615,N_2485);
nor U11725 (N_11725,N_4282,N_2222);
or U11726 (N_11726,N_225,N_3356);
nor U11727 (N_11727,N_2722,N_744);
xor U11728 (N_11728,N_4317,N_155);
nand U11729 (N_11729,N_2743,N_36);
xnor U11730 (N_11730,N_1867,N_5123);
nand U11731 (N_11731,N_1635,N_477);
nand U11732 (N_11732,N_5409,N_4126);
or U11733 (N_11733,N_3749,N_2525);
or U11734 (N_11734,N_853,N_1057);
and U11735 (N_11735,N_2478,N_5683);
nor U11736 (N_11736,N_3480,N_3507);
nand U11737 (N_11737,N_2928,N_5051);
xor U11738 (N_11738,N_5394,N_4724);
and U11739 (N_11739,N_2190,N_5254);
or U11740 (N_11740,N_515,N_2365);
xor U11741 (N_11741,N_351,N_4154);
xnor U11742 (N_11742,N_1645,N_1591);
nor U11743 (N_11743,N_5040,N_3587);
nor U11744 (N_11744,N_5321,N_2902);
nand U11745 (N_11745,N_30,N_939);
nand U11746 (N_11746,N_1566,N_3399);
nor U11747 (N_11747,N_2352,N_5811);
and U11748 (N_11748,N_1322,N_2428);
xor U11749 (N_11749,N_4077,N_4471);
xnor U11750 (N_11750,N_4680,N_680);
and U11751 (N_11751,N_3372,N_3517);
or U11752 (N_11752,N_1756,N_4878);
xnor U11753 (N_11753,N_4320,N_2269);
xnor U11754 (N_11754,N_1290,N_1784);
and U11755 (N_11755,N_2693,N_2225);
or U11756 (N_11756,N_3462,N_4382);
nor U11757 (N_11757,N_2457,N_2744);
or U11758 (N_11758,N_2149,N_2124);
nand U11759 (N_11759,N_22,N_4215);
and U11760 (N_11760,N_3718,N_5998);
or U11761 (N_11761,N_2514,N_5546);
and U11762 (N_11762,N_5486,N_5110);
xnor U11763 (N_11763,N_2483,N_384);
or U11764 (N_11764,N_5415,N_499);
nor U11765 (N_11765,N_3768,N_5045);
and U11766 (N_11766,N_3271,N_4458);
and U11767 (N_11767,N_5806,N_3534);
nand U11768 (N_11768,N_5569,N_492);
nand U11769 (N_11769,N_3755,N_3856);
or U11770 (N_11770,N_2943,N_2959);
xor U11771 (N_11771,N_384,N_4499);
xnor U11772 (N_11772,N_3737,N_4922);
and U11773 (N_11773,N_1550,N_4024);
nand U11774 (N_11774,N_1571,N_2731);
xor U11775 (N_11775,N_1605,N_3817);
and U11776 (N_11776,N_5051,N_5303);
xor U11777 (N_11777,N_1434,N_602);
nand U11778 (N_11778,N_3419,N_2900);
and U11779 (N_11779,N_1084,N_2363);
xnor U11780 (N_11780,N_4272,N_1686);
nor U11781 (N_11781,N_577,N_4147);
nor U11782 (N_11782,N_2681,N_4973);
nand U11783 (N_11783,N_5351,N_667);
and U11784 (N_11784,N_937,N_1733);
or U11785 (N_11785,N_5277,N_5489);
or U11786 (N_11786,N_1295,N_2);
xor U11787 (N_11787,N_210,N_5480);
xnor U11788 (N_11788,N_2841,N_2030);
xnor U11789 (N_11789,N_2246,N_2025);
xor U11790 (N_11790,N_336,N_3667);
and U11791 (N_11791,N_4930,N_1608);
nand U11792 (N_11792,N_5452,N_1386);
nand U11793 (N_11793,N_4251,N_582);
and U11794 (N_11794,N_4723,N_4816);
nand U11795 (N_11795,N_2937,N_429);
and U11796 (N_11796,N_4738,N_4818);
and U11797 (N_11797,N_4894,N_1489);
nand U11798 (N_11798,N_1252,N_5318);
and U11799 (N_11799,N_1063,N_2792);
or U11800 (N_11800,N_2277,N_1677);
nor U11801 (N_11801,N_5180,N_5614);
or U11802 (N_11802,N_2844,N_3298);
xnor U11803 (N_11803,N_1985,N_4562);
or U11804 (N_11804,N_1218,N_5371);
xnor U11805 (N_11805,N_1596,N_3449);
xnor U11806 (N_11806,N_1147,N_4922);
and U11807 (N_11807,N_2192,N_2512);
and U11808 (N_11808,N_4774,N_2228);
and U11809 (N_11809,N_4736,N_2355);
or U11810 (N_11810,N_3016,N_5587);
and U11811 (N_11811,N_2685,N_434);
nand U11812 (N_11812,N_4852,N_5720);
xor U11813 (N_11813,N_5083,N_2245);
xnor U11814 (N_11814,N_5513,N_1722);
or U11815 (N_11815,N_4774,N_3974);
nand U11816 (N_11816,N_2811,N_2621);
xnor U11817 (N_11817,N_272,N_4833);
xor U11818 (N_11818,N_3011,N_2085);
xor U11819 (N_11819,N_3395,N_1465);
xor U11820 (N_11820,N_257,N_5613);
nand U11821 (N_11821,N_3552,N_2551);
and U11822 (N_11822,N_5684,N_4225);
xnor U11823 (N_11823,N_3415,N_1280);
nor U11824 (N_11824,N_3019,N_3940);
or U11825 (N_11825,N_2806,N_5821);
xor U11826 (N_11826,N_5118,N_1750);
and U11827 (N_11827,N_143,N_4888);
and U11828 (N_11828,N_4259,N_2720);
and U11829 (N_11829,N_824,N_4206);
or U11830 (N_11830,N_1028,N_2653);
and U11831 (N_11831,N_5512,N_1638);
or U11832 (N_11832,N_2181,N_5120);
nand U11833 (N_11833,N_5059,N_3537);
or U11834 (N_11834,N_2833,N_3926);
and U11835 (N_11835,N_1519,N_2490);
and U11836 (N_11836,N_625,N_5662);
and U11837 (N_11837,N_1413,N_2689);
nand U11838 (N_11838,N_2370,N_4060);
nand U11839 (N_11839,N_2539,N_4658);
and U11840 (N_11840,N_4056,N_1456);
and U11841 (N_11841,N_3347,N_3276);
and U11842 (N_11842,N_1975,N_4706);
or U11843 (N_11843,N_373,N_5101);
or U11844 (N_11844,N_5119,N_144);
or U11845 (N_11845,N_3653,N_4555);
and U11846 (N_11846,N_5708,N_105);
nand U11847 (N_11847,N_3755,N_255);
and U11848 (N_11848,N_619,N_1396);
xor U11849 (N_11849,N_759,N_2846);
and U11850 (N_11850,N_3263,N_5221);
and U11851 (N_11851,N_1860,N_5545);
xnor U11852 (N_11852,N_2040,N_3311);
xor U11853 (N_11853,N_3619,N_1878);
and U11854 (N_11854,N_5521,N_1611);
or U11855 (N_11855,N_3165,N_1094);
and U11856 (N_11856,N_5315,N_707);
or U11857 (N_11857,N_3783,N_3537);
xor U11858 (N_11858,N_5475,N_5366);
xnor U11859 (N_11859,N_3919,N_4951);
or U11860 (N_11860,N_5402,N_4322);
nand U11861 (N_11861,N_3758,N_1933);
nor U11862 (N_11862,N_2214,N_5307);
xnor U11863 (N_11863,N_2701,N_913);
and U11864 (N_11864,N_3237,N_1696);
xor U11865 (N_11865,N_3238,N_5269);
nor U11866 (N_11866,N_5440,N_5846);
nor U11867 (N_11867,N_3702,N_4985);
or U11868 (N_11868,N_592,N_417);
or U11869 (N_11869,N_4917,N_5842);
or U11870 (N_11870,N_3088,N_5196);
nor U11871 (N_11871,N_2887,N_3345);
or U11872 (N_11872,N_1014,N_268);
nand U11873 (N_11873,N_3789,N_1614);
nand U11874 (N_11874,N_606,N_5882);
nand U11875 (N_11875,N_5682,N_4220);
or U11876 (N_11876,N_1843,N_4896);
xor U11877 (N_11877,N_88,N_5116);
xor U11878 (N_11878,N_11,N_2838);
nor U11879 (N_11879,N_679,N_722);
nor U11880 (N_11880,N_3352,N_1051);
nand U11881 (N_11881,N_784,N_1754);
nor U11882 (N_11882,N_1820,N_2665);
nor U11883 (N_11883,N_1468,N_4185);
xor U11884 (N_11884,N_1875,N_3286);
and U11885 (N_11885,N_4778,N_876);
nand U11886 (N_11886,N_4662,N_1611);
nor U11887 (N_11887,N_2005,N_2394);
nor U11888 (N_11888,N_4077,N_3956);
or U11889 (N_11889,N_5219,N_43);
and U11890 (N_11890,N_4108,N_3095);
nand U11891 (N_11891,N_5539,N_2628);
xor U11892 (N_11892,N_2766,N_1916);
nor U11893 (N_11893,N_5323,N_158);
and U11894 (N_11894,N_1582,N_4213);
and U11895 (N_11895,N_5532,N_476);
or U11896 (N_11896,N_2809,N_872);
nand U11897 (N_11897,N_4250,N_230);
and U11898 (N_11898,N_4993,N_748);
or U11899 (N_11899,N_5583,N_3146);
xor U11900 (N_11900,N_4880,N_2051);
xor U11901 (N_11901,N_2051,N_5868);
xor U11902 (N_11902,N_4942,N_1214);
xor U11903 (N_11903,N_250,N_4022);
nand U11904 (N_11904,N_463,N_3920);
xnor U11905 (N_11905,N_301,N_4496);
or U11906 (N_11906,N_778,N_112);
and U11907 (N_11907,N_4868,N_1243);
and U11908 (N_11908,N_5671,N_645);
or U11909 (N_11909,N_343,N_3186);
nand U11910 (N_11910,N_4594,N_5697);
nor U11911 (N_11911,N_5513,N_2688);
or U11912 (N_11912,N_3285,N_2831);
nand U11913 (N_11913,N_4165,N_867);
xnor U11914 (N_11914,N_3316,N_3896);
or U11915 (N_11915,N_1562,N_5954);
nand U11916 (N_11916,N_4378,N_4227);
xor U11917 (N_11917,N_2911,N_4436);
and U11918 (N_11918,N_2657,N_325);
or U11919 (N_11919,N_633,N_2373);
or U11920 (N_11920,N_3840,N_4854);
nor U11921 (N_11921,N_2830,N_5876);
nand U11922 (N_11922,N_1736,N_4526);
and U11923 (N_11923,N_1192,N_2559);
and U11924 (N_11924,N_4363,N_1936);
nor U11925 (N_11925,N_1172,N_1117);
nor U11926 (N_11926,N_2030,N_1473);
xor U11927 (N_11927,N_458,N_4832);
or U11928 (N_11928,N_4296,N_628);
xnor U11929 (N_11929,N_138,N_2394);
and U11930 (N_11930,N_2708,N_2604);
xnor U11931 (N_11931,N_24,N_227);
or U11932 (N_11932,N_1342,N_4691);
or U11933 (N_11933,N_3007,N_1129);
xor U11934 (N_11934,N_2029,N_3146);
or U11935 (N_11935,N_5754,N_1947);
and U11936 (N_11936,N_2940,N_3548);
nor U11937 (N_11937,N_2835,N_2216);
nor U11938 (N_11938,N_475,N_4676);
and U11939 (N_11939,N_792,N_2912);
or U11940 (N_11940,N_360,N_5524);
nand U11941 (N_11941,N_2686,N_4939);
nand U11942 (N_11942,N_1525,N_4678);
xnor U11943 (N_11943,N_5474,N_4817);
nor U11944 (N_11944,N_4117,N_3085);
xnor U11945 (N_11945,N_5696,N_2049);
nor U11946 (N_11946,N_2826,N_2233);
or U11947 (N_11947,N_3080,N_2126);
nand U11948 (N_11948,N_5243,N_2435);
or U11949 (N_11949,N_4170,N_1158);
or U11950 (N_11950,N_3943,N_531);
xor U11951 (N_11951,N_1166,N_4829);
or U11952 (N_11952,N_3232,N_1124);
nor U11953 (N_11953,N_828,N_1726);
nor U11954 (N_11954,N_4588,N_531);
nand U11955 (N_11955,N_5365,N_425);
nand U11956 (N_11956,N_299,N_1819);
nand U11957 (N_11957,N_1785,N_5224);
and U11958 (N_11958,N_4926,N_884);
xor U11959 (N_11959,N_2321,N_3991);
and U11960 (N_11960,N_4515,N_4532);
nand U11961 (N_11961,N_5089,N_4655);
or U11962 (N_11962,N_1367,N_2663);
xor U11963 (N_11963,N_294,N_5596);
and U11964 (N_11964,N_4959,N_915);
xor U11965 (N_11965,N_5026,N_4978);
xor U11966 (N_11966,N_858,N_3669);
nor U11967 (N_11967,N_1997,N_1960);
xnor U11968 (N_11968,N_221,N_3820);
nor U11969 (N_11969,N_3807,N_5727);
xnor U11970 (N_11970,N_2857,N_906);
and U11971 (N_11971,N_528,N_1556);
nor U11972 (N_11972,N_1948,N_867);
nand U11973 (N_11973,N_2854,N_2729);
or U11974 (N_11974,N_2884,N_432);
and U11975 (N_11975,N_2742,N_2945);
or U11976 (N_11976,N_1587,N_5910);
and U11977 (N_11977,N_2866,N_3133);
and U11978 (N_11978,N_2555,N_4315);
or U11979 (N_11979,N_3776,N_3487);
nand U11980 (N_11980,N_54,N_4041);
or U11981 (N_11981,N_4019,N_803);
or U11982 (N_11982,N_2023,N_5037);
nand U11983 (N_11983,N_2300,N_4165);
and U11984 (N_11984,N_3739,N_599);
nor U11985 (N_11985,N_3066,N_5494);
nor U11986 (N_11986,N_5887,N_2912);
nor U11987 (N_11987,N_2933,N_2509);
xnor U11988 (N_11988,N_5244,N_3979);
or U11989 (N_11989,N_3715,N_5861);
or U11990 (N_11990,N_2926,N_1927);
or U11991 (N_11991,N_2587,N_4418);
xor U11992 (N_11992,N_1874,N_4190);
and U11993 (N_11993,N_1961,N_1029);
and U11994 (N_11994,N_2576,N_603);
xnor U11995 (N_11995,N_4954,N_830);
nand U11996 (N_11996,N_5016,N_3479);
nor U11997 (N_11997,N_4555,N_4116);
xor U11998 (N_11998,N_1494,N_5836);
and U11999 (N_11999,N_5929,N_2088);
xnor U12000 (N_12000,N_6540,N_11459);
nand U12001 (N_12001,N_10955,N_10542);
nand U12002 (N_12002,N_10673,N_6041);
xnor U12003 (N_12003,N_10766,N_10048);
nand U12004 (N_12004,N_8418,N_8607);
or U12005 (N_12005,N_9078,N_8738);
xnor U12006 (N_12006,N_8626,N_7393);
xnor U12007 (N_12007,N_6498,N_6117);
and U12008 (N_12008,N_10055,N_11247);
nand U12009 (N_12009,N_9217,N_9375);
nand U12010 (N_12010,N_8494,N_7287);
nand U12011 (N_12011,N_9734,N_8481);
or U12012 (N_12012,N_10422,N_7415);
nand U12013 (N_12013,N_11258,N_6304);
xnor U12014 (N_12014,N_11624,N_11664);
xor U12015 (N_12015,N_8714,N_11505);
xor U12016 (N_12016,N_8147,N_11604);
xnor U12017 (N_12017,N_7298,N_11305);
or U12018 (N_12018,N_9194,N_6808);
and U12019 (N_12019,N_11701,N_8975);
and U12020 (N_12020,N_9663,N_7693);
nand U12021 (N_12021,N_9881,N_10167);
xnor U12022 (N_12022,N_9168,N_6620);
xnor U12023 (N_12023,N_7291,N_7252);
xnor U12024 (N_12024,N_10100,N_8369);
and U12025 (N_12025,N_11808,N_7228);
and U12026 (N_12026,N_8326,N_11140);
and U12027 (N_12027,N_10828,N_10540);
and U12028 (N_12028,N_7650,N_8917);
nand U12029 (N_12029,N_8403,N_6380);
xor U12030 (N_12030,N_11581,N_8094);
and U12031 (N_12031,N_9267,N_10792);
and U12032 (N_12032,N_8777,N_11519);
xnor U12033 (N_12033,N_8020,N_6306);
nor U12034 (N_12034,N_6678,N_9290);
nand U12035 (N_12035,N_7408,N_8669);
nand U12036 (N_12036,N_11399,N_11680);
nor U12037 (N_12037,N_8176,N_7741);
nand U12038 (N_12038,N_6581,N_7555);
nand U12039 (N_12039,N_9690,N_11048);
nand U12040 (N_12040,N_10757,N_8304);
or U12041 (N_12041,N_6630,N_6378);
and U12042 (N_12042,N_7307,N_10722);
xor U12043 (N_12043,N_11698,N_9334);
xnor U12044 (N_12044,N_7592,N_10341);
nand U12045 (N_12045,N_8531,N_10855);
and U12046 (N_12046,N_6456,N_11386);
or U12047 (N_12047,N_11997,N_7721);
xor U12048 (N_12048,N_6485,N_9356);
nand U12049 (N_12049,N_8128,N_7559);
and U12050 (N_12050,N_7691,N_10661);
nand U12051 (N_12051,N_8084,N_11354);
or U12052 (N_12052,N_9408,N_11525);
nor U12053 (N_12053,N_10162,N_9170);
xnor U12054 (N_12054,N_8796,N_7364);
xnor U12055 (N_12055,N_10275,N_10689);
xor U12056 (N_12056,N_11271,N_9232);
nor U12057 (N_12057,N_7867,N_10567);
nor U12058 (N_12058,N_8955,N_8654);
or U12059 (N_12059,N_6749,N_10186);
or U12060 (N_12060,N_10132,N_9101);
nor U12061 (N_12061,N_10406,N_8895);
xor U12062 (N_12062,N_7070,N_9965);
or U12063 (N_12063,N_7316,N_8981);
or U12064 (N_12064,N_11577,N_9973);
nor U12065 (N_12065,N_8676,N_9084);
nand U12066 (N_12066,N_7335,N_7714);
nor U12067 (N_12067,N_11380,N_10986);
and U12068 (N_12068,N_6008,N_10071);
and U12069 (N_12069,N_6431,N_6918);
and U12070 (N_12070,N_9887,N_9893);
or U12071 (N_12071,N_9717,N_6675);
nor U12072 (N_12072,N_6504,N_8642);
nand U12073 (N_12073,N_10089,N_11243);
and U12074 (N_12074,N_10631,N_8284);
nor U12075 (N_12075,N_10262,N_11544);
xnor U12076 (N_12076,N_8994,N_10934);
nand U12077 (N_12077,N_10664,N_6789);
nor U12078 (N_12078,N_8423,N_9668);
nor U12079 (N_12079,N_7088,N_9361);
and U12080 (N_12080,N_8733,N_10991);
xor U12081 (N_12081,N_7340,N_10650);
nand U12082 (N_12082,N_10534,N_9180);
and U12083 (N_12083,N_7068,N_9132);
or U12084 (N_12084,N_7853,N_6220);
and U12085 (N_12085,N_10491,N_7541);
xnor U12086 (N_12086,N_9343,N_8687);
nand U12087 (N_12087,N_6755,N_6059);
or U12088 (N_12088,N_11865,N_9975);
nor U12089 (N_12089,N_8258,N_6418);
nand U12090 (N_12090,N_11830,N_7821);
xor U12091 (N_12091,N_9289,N_11368);
xnor U12092 (N_12092,N_9569,N_11875);
nor U12093 (N_12093,N_10875,N_7229);
and U12094 (N_12094,N_8042,N_9857);
nand U12095 (N_12095,N_10470,N_11129);
and U12096 (N_12096,N_9910,N_9713);
or U12097 (N_12097,N_6164,N_10847);
nor U12098 (N_12098,N_7802,N_11475);
nand U12099 (N_12099,N_7005,N_7026);
nand U12100 (N_12100,N_9932,N_6539);
nor U12101 (N_12101,N_9622,N_11965);
xnor U12102 (N_12102,N_9620,N_10354);
nor U12103 (N_12103,N_11289,N_6005);
nand U12104 (N_12104,N_11576,N_8774);
nand U12105 (N_12105,N_9251,N_9712);
xor U12106 (N_12106,N_6238,N_7784);
and U12107 (N_12107,N_11104,N_8916);
and U12108 (N_12108,N_7869,N_7777);
nor U12109 (N_12109,N_7572,N_10874);
or U12110 (N_12110,N_6419,N_8978);
and U12111 (N_12111,N_11326,N_8844);
xor U12112 (N_12112,N_10723,N_8300);
and U12113 (N_12113,N_9417,N_9562);
nor U12114 (N_12114,N_11099,N_11801);
nor U12115 (N_12115,N_9803,N_8116);
nor U12116 (N_12116,N_6994,N_9039);
nor U12117 (N_12117,N_11187,N_6371);
and U12118 (N_12118,N_9166,N_7664);
nor U12119 (N_12119,N_6727,N_9397);
or U12120 (N_12120,N_6244,N_8689);
nor U12121 (N_12121,N_11824,N_6073);
and U12122 (N_12122,N_10392,N_11298);
and U12123 (N_12123,N_9777,N_6267);
nand U12124 (N_12124,N_8788,N_10767);
or U12125 (N_12125,N_7808,N_7654);
nand U12126 (N_12126,N_9792,N_6217);
nor U12127 (N_12127,N_10559,N_10786);
nand U12128 (N_12128,N_10046,N_7234);
and U12129 (N_12129,N_10806,N_7297);
or U12130 (N_12130,N_10479,N_7872);
and U12131 (N_12131,N_8853,N_11421);
xnor U12132 (N_12132,N_6021,N_9287);
nor U12133 (N_12133,N_9727,N_11778);
and U12134 (N_12134,N_11053,N_6616);
xnor U12135 (N_12135,N_8050,N_8396);
or U12136 (N_12136,N_6707,N_6200);
and U12137 (N_12137,N_8124,N_9344);
nand U12138 (N_12138,N_6828,N_9189);
or U12139 (N_12139,N_11898,N_7000);
xnor U12140 (N_12140,N_11699,N_8139);
and U12141 (N_12141,N_10781,N_8903);
nand U12142 (N_12142,N_11467,N_10105);
or U12143 (N_12143,N_11396,N_8108);
xor U12144 (N_12144,N_9383,N_10758);
or U12145 (N_12145,N_10982,N_9754);
or U12146 (N_12146,N_8239,N_9821);
nor U12147 (N_12147,N_10575,N_10395);
xnor U12148 (N_12148,N_8553,N_10798);
and U12149 (N_12149,N_10255,N_7757);
nand U12150 (N_12150,N_11920,N_7826);
and U12151 (N_12151,N_10173,N_7024);
nor U12152 (N_12152,N_8941,N_11630);
nor U12153 (N_12153,N_10373,N_7280);
or U12154 (N_12154,N_7686,N_6621);
xor U12155 (N_12155,N_6338,N_7161);
or U12156 (N_12156,N_9843,N_11737);
and U12157 (N_12157,N_8910,N_10908);
nor U12158 (N_12158,N_7842,N_7712);
or U12159 (N_12159,N_9260,N_6061);
and U12160 (N_12160,N_6113,N_11314);
and U12161 (N_12161,N_6915,N_11620);
nand U12162 (N_12162,N_7697,N_9427);
nand U12163 (N_12163,N_6078,N_7414);
xnor U12164 (N_12164,N_10620,N_8424);
nand U12165 (N_12165,N_8897,N_8806);
nand U12166 (N_12166,N_11647,N_8333);
xnor U12167 (N_12167,N_9323,N_9915);
and U12168 (N_12168,N_10456,N_9409);
nand U12169 (N_12169,N_11523,N_9658);
and U12170 (N_12170,N_7244,N_6387);
and U12171 (N_12171,N_8500,N_7497);
nand U12172 (N_12172,N_8133,N_10235);
nor U12173 (N_12173,N_6365,N_6770);
nand U12174 (N_12174,N_7300,N_11853);
and U12175 (N_12175,N_7780,N_10371);
xnor U12176 (N_12176,N_10247,N_9238);
or U12177 (N_12177,N_7695,N_6328);
nor U12178 (N_12178,N_10051,N_11278);
and U12179 (N_12179,N_8080,N_7602);
or U12180 (N_12180,N_7486,N_10180);
xor U12181 (N_12181,N_9228,N_8431);
xor U12182 (N_12182,N_6401,N_7806);
and U12183 (N_12183,N_6800,N_7525);
xnor U12184 (N_12184,N_9788,N_10599);
nand U12185 (N_12185,N_9675,N_9426);
nor U12186 (N_12186,N_8440,N_10049);
or U12187 (N_12187,N_11712,N_11330);
nor U12188 (N_12188,N_8259,N_7239);
or U12189 (N_12189,N_8739,N_9220);
nor U12190 (N_12190,N_11015,N_11975);
and U12191 (N_12191,N_9917,N_7450);
xnor U12192 (N_12192,N_7223,N_8013);
or U12193 (N_12193,N_10040,N_10230);
nor U12194 (N_12194,N_6051,N_7934);
nor U12195 (N_12195,N_10229,N_9859);
and U12196 (N_12196,N_7659,N_10367);
nor U12197 (N_12197,N_11339,N_9007);
nand U12198 (N_12198,N_10233,N_7220);
nand U12199 (N_12199,N_10912,N_6390);
nand U12200 (N_12200,N_10130,N_9762);
or U12201 (N_12201,N_11291,N_6774);
nand U12202 (N_12202,N_6657,N_8366);
or U12203 (N_12203,N_9799,N_6474);
or U12204 (N_12204,N_10648,N_6721);
or U12205 (N_12205,N_11121,N_11747);
and U12206 (N_12206,N_6705,N_6801);
nor U12207 (N_12207,N_7194,N_6744);
or U12208 (N_12208,N_10808,N_7775);
nand U12209 (N_12209,N_7539,N_6096);
nor U12210 (N_12210,N_10822,N_11041);
nand U12211 (N_12211,N_6559,N_8537);
xor U12212 (N_12212,N_8862,N_10091);
and U12213 (N_12213,N_7331,N_6099);
nand U12214 (N_12214,N_9879,N_9381);
and U12215 (N_12215,N_9738,N_6085);
and U12216 (N_12216,N_6946,N_6111);
xor U12217 (N_12217,N_11363,N_10950);
and U12218 (N_12218,N_11832,N_6564);
nand U12219 (N_12219,N_7455,N_9143);
xnor U12220 (N_12220,N_11275,N_9025);
nor U12221 (N_12221,N_9035,N_7681);
or U12222 (N_12222,N_11137,N_9532);
nand U12223 (N_12223,N_8538,N_9337);
xnor U12224 (N_12224,N_8245,N_11110);
nand U12225 (N_12225,N_10635,N_9233);
or U12226 (N_12226,N_8302,N_6364);
or U12227 (N_12227,N_10613,N_10602);
nand U12228 (N_12228,N_11014,N_8056);
or U12229 (N_12229,N_6221,N_7109);
and U12230 (N_12230,N_9031,N_10211);
nor U12231 (N_12231,N_7818,N_8331);
nand U12232 (N_12232,N_7571,N_9372);
xor U12233 (N_12233,N_10860,N_7781);
nor U12234 (N_12234,N_7150,N_10590);
or U12235 (N_12235,N_7803,N_7878);
xor U12236 (N_12236,N_11115,N_7608);
xor U12237 (N_12237,N_11654,N_8037);
nand U12238 (N_12238,N_6036,N_10878);
nor U12239 (N_12239,N_10183,N_10800);
nand U12240 (N_12240,N_10928,N_6553);
or U12241 (N_12241,N_9732,N_10363);
nand U12242 (N_12242,N_11311,N_10972);
nand U12243 (N_12243,N_7404,N_8857);
and U12244 (N_12244,N_8265,N_11955);
xnor U12245 (N_12245,N_10768,N_9850);
nand U12246 (N_12246,N_11583,N_10493);
nor U12247 (N_12247,N_11557,N_10434);
nor U12248 (N_12248,N_8047,N_7957);
and U12249 (N_12249,N_8623,N_6792);
xor U12250 (N_12250,N_6797,N_7547);
nand U12251 (N_12251,N_6053,N_7633);
or U12252 (N_12252,N_10699,N_8675);
and U12253 (N_12253,N_6140,N_11580);
xor U12254 (N_12254,N_10372,N_6382);
xnor U12255 (N_12255,N_8453,N_7827);
xnor U12256 (N_12256,N_11704,N_7049);
xnor U12257 (N_12257,N_8264,N_10345);
or U12258 (N_12258,N_7015,N_10578);
or U12259 (N_12259,N_11112,N_10539);
or U12260 (N_12260,N_8329,N_9662);
nand U12261 (N_12261,N_11681,N_11871);
nor U12262 (N_12262,N_9116,N_6854);
nand U12263 (N_12263,N_8564,N_10464);
or U12264 (N_12264,N_6628,N_9807);
and U12265 (N_12265,N_7709,N_10248);
nor U12266 (N_12266,N_10939,N_7983);
and U12267 (N_12267,N_10201,N_6100);
or U12268 (N_12268,N_8715,N_7584);
xor U12269 (N_12269,N_10576,N_9967);
xnor U12270 (N_12270,N_11161,N_7167);
and U12271 (N_12271,N_6398,N_8413);
nand U12272 (N_12272,N_6681,N_11987);
and U12273 (N_12273,N_7212,N_11001);
or U12274 (N_12274,N_6243,N_8855);
and U12275 (N_12275,N_11829,N_9244);
nand U12276 (N_12276,N_6237,N_10020);
and U12277 (N_12277,N_10283,N_6529);
or U12278 (N_12278,N_8439,N_8301);
xnor U12279 (N_12279,N_6700,N_6986);
and U12280 (N_12280,N_8604,N_10216);
nand U12281 (N_12281,N_6124,N_6092);
xnor U12282 (N_12282,N_10858,N_6460);
and U12283 (N_12283,N_7982,N_7427);
nor U12284 (N_12284,N_10155,N_9470);
xor U12285 (N_12285,N_6632,N_7158);
nand U12286 (N_12286,N_11274,N_8556);
nor U12287 (N_12287,N_8520,N_8241);
nor U12288 (N_12288,N_6031,N_9855);
nor U12289 (N_12289,N_9218,N_11558);
or U12290 (N_12290,N_9399,N_6511);
nor U12291 (N_12291,N_7852,N_9851);
and U12292 (N_12292,N_7887,N_10328);
nand U12293 (N_12293,N_7544,N_7516);
and U12294 (N_12294,N_8421,N_6533);
nand U12295 (N_12295,N_9638,N_10817);
or U12296 (N_12296,N_9618,N_8719);
xor U12297 (N_12297,N_6742,N_8129);
or U12298 (N_12298,N_9169,N_8711);
nand U12299 (N_12299,N_8804,N_9804);
xor U12300 (N_12300,N_6720,N_8352);
nor U12301 (N_12301,N_9537,N_10465);
or U12302 (N_12302,N_9506,N_11961);
nor U12303 (N_12303,N_7342,N_7357);
or U12304 (N_12304,N_6793,N_8647);
nand U12305 (N_12305,N_6670,N_6664);
xor U12306 (N_12306,N_6965,N_9311);
and U12307 (N_12307,N_7594,N_7046);
or U12308 (N_12308,N_8327,N_7372);
and U12309 (N_12309,N_11621,N_10690);
nand U12310 (N_12310,N_10962,N_9321);
and U12311 (N_12311,N_11530,N_10351);
nor U12312 (N_12312,N_10121,N_10831);
nand U12313 (N_12313,N_11803,N_7922);
nor U12314 (N_12314,N_6052,N_11455);
xor U12315 (N_12315,N_10555,N_6889);
xor U12316 (N_12316,N_7834,N_10067);
and U12317 (N_12317,N_9566,N_9403);
nand U12318 (N_12318,N_6831,N_10742);
nand U12319 (N_12319,N_9993,N_10510);
nand U12320 (N_12320,N_8203,N_7396);
nor U12321 (N_12321,N_8018,N_7155);
or U12322 (N_12322,N_9048,N_11249);
nand U12323 (N_12323,N_7771,N_11691);
or U12324 (N_12324,N_7743,N_9095);
or U12325 (N_12325,N_10148,N_6395);
nand U12326 (N_12326,N_7805,N_9500);
and U12327 (N_12327,N_7801,N_9045);
or U12328 (N_12328,N_9581,N_11083);
or U12329 (N_12329,N_6210,N_10625);
nor U12330 (N_12330,N_7487,N_6665);
or U12331 (N_12331,N_9933,N_11360);
xnor U12332 (N_12332,N_11619,N_6692);
nand U12333 (N_12333,N_7104,N_7875);
or U12334 (N_12334,N_7447,N_6483);
xor U12335 (N_12335,N_8314,N_10305);
nand U12336 (N_12336,N_8528,N_10423);
nand U12337 (N_12337,N_10407,N_8864);
nand U12338 (N_12338,N_8398,N_6601);
nand U12339 (N_12339,N_11128,N_8361);
nand U12340 (N_12340,N_10730,N_7341);
nand U12341 (N_12341,N_8513,N_7330);
and U12342 (N_12342,N_10017,N_11652);
nand U12343 (N_12343,N_11719,N_11253);
xnor U12344 (N_12344,N_11081,N_9086);
xor U12345 (N_12345,N_10488,N_8967);
nor U12346 (N_12346,N_10694,N_8816);
or U12347 (N_12347,N_11716,N_7689);
nor U12348 (N_12348,N_9496,N_7025);
or U12349 (N_12349,N_6453,N_10643);
xnor U12350 (N_12350,N_10866,N_11566);
or U12351 (N_12351,N_10789,N_8560);
nor U12352 (N_12352,N_7920,N_6989);
xnor U12353 (N_12353,N_10851,N_6050);
or U12354 (N_12354,N_11542,N_7997);
and U12355 (N_12355,N_9872,N_6772);
nor U12356 (N_12356,N_8803,N_6250);
and U12357 (N_12357,N_11711,N_6871);
xnor U12358 (N_12358,N_9960,N_9834);
nand U12359 (N_12359,N_9626,N_9655);
nand U12360 (N_12360,N_6876,N_11895);
or U12361 (N_12361,N_11184,N_8939);
and U12362 (N_12362,N_10289,N_7185);
nand U12363 (N_12363,N_10923,N_9840);
xnor U12364 (N_12364,N_9302,N_8943);
nand U12365 (N_12365,N_8089,N_6367);
nor U12366 (N_12366,N_6806,N_11886);
xor U12367 (N_12367,N_7529,N_11607);
nor U12368 (N_12368,N_7075,N_8613);
nor U12369 (N_12369,N_9012,N_10894);
or U12370 (N_12370,N_10770,N_11492);
nand U12371 (N_12371,N_6937,N_7910);
nor U12372 (N_12372,N_7765,N_7549);
xnor U12373 (N_12373,N_8652,N_11193);
and U12374 (N_12374,N_6852,N_9679);
or U12375 (N_12375,N_10992,N_8201);
xnor U12376 (N_12376,N_11199,N_11605);
or U12377 (N_12377,N_10966,N_8950);
nor U12378 (N_12378,N_6934,N_7640);
or U12379 (N_12379,N_8712,N_6415);
nor U12380 (N_12380,N_8610,N_8621);
nor U12381 (N_12381,N_9494,N_11606);
nor U12382 (N_12382,N_11248,N_11295);
xnor U12383 (N_12383,N_7948,N_10813);
xnor U12384 (N_12384,N_6291,N_8223);
nor U12385 (N_12385,N_7688,N_10172);
nor U12386 (N_12386,N_11230,N_10696);
xnor U12387 (N_12387,N_6642,N_6082);
xnor U12388 (N_12388,N_6935,N_11833);
and U12389 (N_12389,N_8492,N_10279);
nand U12390 (N_12390,N_9339,N_11097);
xor U12391 (N_12391,N_8743,N_10221);
xor U12392 (N_12392,N_8210,N_6607);
and U12393 (N_12393,N_8918,N_9136);
nor U12394 (N_12394,N_11792,N_7861);
and U12395 (N_12395,N_10317,N_7763);
or U12396 (N_12396,N_6216,N_11946);
xor U12397 (N_12397,N_7717,N_8160);
and U12398 (N_12398,N_11919,N_7864);
nand U12399 (N_12399,N_8106,N_10658);
or U12400 (N_12400,N_6068,N_6815);
xnor U12401 (N_12401,N_9241,N_6538);
and U12402 (N_12402,N_7774,N_9837);
or U12403 (N_12403,N_11316,N_9367);
nand U12404 (N_12404,N_9199,N_7125);
nor U12405 (N_12405,N_11046,N_11469);
or U12406 (N_12406,N_9684,N_7115);
xnor U12407 (N_12407,N_6207,N_8792);
or U12408 (N_12408,N_6039,N_11448);
and U12409 (N_12409,N_11934,N_6184);
or U12410 (N_12410,N_8673,N_6942);
nor U12411 (N_12411,N_10411,N_9695);
nor U12412 (N_12412,N_9032,N_6143);
xor U12413 (N_12413,N_7198,N_7116);
nand U12414 (N_12414,N_10885,N_8174);
or U12415 (N_12415,N_8581,N_7204);
xor U12416 (N_12416,N_8178,N_10915);
or U12417 (N_12417,N_7279,N_11706);
nand U12418 (N_12418,N_6583,N_9793);
nor U12419 (N_12419,N_11478,N_10557);
or U12420 (N_12420,N_11457,N_11256);
nor U12421 (N_12421,N_6163,N_9904);
nand U12422 (N_12422,N_7945,N_11036);
nor U12423 (N_12423,N_8249,N_11250);
nor U12424 (N_12424,N_8303,N_7747);
and U12425 (N_12425,N_7819,N_9573);
nand U12426 (N_12426,N_11513,N_6376);
and U12427 (N_12427,N_10708,N_8000);
and U12428 (N_12428,N_9276,N_8758);
nand U12429 (N_12429,N_11283,N_9196);
or U12430 (N_12430,N_8426,N_6669);
and U12431 (N_12431,N_6001,N_9480);
nor U12432 (N_12432,N_7295,N_11755);
nor U12433 (N_12433,N_11493,N_11645);
xor U12434 (N_12434,N_8725,N_8574);
xor U12435 (N_12435,N_8659,N_7030);
xor U12436 (N_12436,N_8121,N_10206);
nor U12437 (N_12437,N_6199,N_7169);
nand U12438 (N_12438,N_6762,N_8883);
nor U12439 (N_12439,N_9865,N_9471);
nand U12440 (N_12440,N_8888,N_8313);
nor U12441 (N_12441,N_8278,N_6997);
xnor U12442 (N_12442,N_10197,N_6107);
xor U12443 (N_12443,N_7646,N_10053);
or U12444 (N_12444,N_11391,N_8996);
or U12445 (N_12445,N_11464,N_10905);
and U12446 (N_12446,N_10104,N_6322);
or U12447 (N_12447,N_6780,N_9715);
xor U12448 (N_12448,N_9903,N_10124);
nor U12449 (N_12449,N_10118,N_10639);
or U12450 (N_12450,N_9280,N_9466);
nor U12451 (N_12451,N_8944,N_9605);
or U12452 (N_12452,N_8218,N_8963);
xor U12453 (N_12453,N_9130,N_9111);
xor U12454 (N_12454,N_9597,N_10628);
or U12455 (N_12455,N_10189,N_10429);
xnor U12456 (N_12456,N_6104,N_6270);
and U12457 (N_12457,N_11907,N_11150);
or U12458 (N_12458,N_8270,N_10850);
or U12459 (N_12459,N_7314,N_9414);
nor U12460 (N_12460,N_6834,N_7029);
nor U12461 (N_12461,N_11224,N_10794);
nor U12462 (N_12462,N_7038,N_8416);
nor U12463 (N_12463,N_11254,N_10942);
xnor U12464 (N_12464,N_6028,N_8100);
xnor U12465 (N_12465,N_6558,N_7459);
or U12466 (N_12466,N_9516,N_11034);
or U12467 (N_12467,N_10734,N_6475);
nand U12468 (N_12468,N_9949,N_8705);
nand U12469 (N_12469,N_7749,N_11126);
or U12470 (N_12470,N_11154,N_9393);
xor U12471 (N_12471,N_7092,N_8860);
xnor U12472 (N_12472,N_10772,N_10056);
nand U12473 (N_12473,N_7052,N_6286);
or U12474 (N_12474,N_8800,N_6927);
nand U12475 (N_12475,N_8901,N_11504);
nor U12476 (N_12476,N_11893,N_10277);
and U12477 (N_12477,N_9152,N_9273);
nor U12478 (N_12478,N_11731,N_6614);
xor U12479 (N_12479,N_9291,N_11425);
nor U12480 (N_12480,N_8510,N_7203);
nand U12481 (N_12481,N_10432,N_11892);
nor U12482 (N_12482,N_7352,N_11143);
nor U12483 (N_12483,N_7387,N_10519);
and U12484 (N_12484,N_7666,N_6305);
or U12485 (N_12485,N_8697,N_11553);
nand U12486 (N_12486,N_9721,N_6549);
nor U12487 (N_12487,N_10990,N_9345);
and U12488 (N_12488,N_8679,N_8049);
nor U12489 (N_12489,N_11214,N_7890);
xnor U12490 (N_12490,N_9058,N_8281);
nand U12491 (N_12491,N_6318,N_9833);
xor U12492 (N_12492,N_10701,N_9680);
xor U12493 (N_12493,N_7673,N_9292);
or U12494 (N_12494,N_11799,N_9546);
nand U12495 (N_12495,N_10615,N_7475);
nand U12496 (N_12496,N_9747,N_8987);
nand U12497 (N_12497,N_10083,N_11375);
or U12498 (N_12498,N_10738,N_10747);
nand U12499 (N_12499,N_6070,N_9875);
nor U12500 (N_12500,N_8957,N_11724);
and U12501 (N_12501,N_6423,N_6525);
or U12502 (N_12502,N_10603,N_10125);
xor U12503 (N_12503,N_9406,N_6582);
or U12504 (N_12504,N_11261,N_6303);
and U12505 (N_12505,N_6256,N_10359);
or U12506 (N_12506,N_6515,N_9431);
xnor U12507 (N_12507,N_9647,N_7967);
nand U12508 (N_12508,N_7443,N_7736);
nor U12509 (N_12509,N_7776,N_6491);
or U12510 (N_12510,N_9644,N_7242);
nor U12511 (N_12511,N_7611,N_7886);
and U12512 (N_12512,N_10930,N_9079);
nor U12513 (N_12513,N_9912,N_9866);
xor U12514 (N_12514,N_11656,N_9446);
nor U12515 (N_12515,N_9478,N_11173);
xnor U12516 (N_12516,N_7014,N_6747);
nor U12517 (N_12517,N_7752,N_10092);
nor U12518 (N_12518,N_9895,N_8933);
xnor U12519 (N_12519,N_10593,N_6197);
nand U12520 (N_12520,N_6905,N_8310);
or U12521 (N_12521,N_7502,N_9110);
nor U12522 (N_12522,N_11483,N_7665);
or U12523 (N_12523,N_7462,N_11913);
nor U12524 (N_12524,N_7449,N_8890);
nand U12525 (N_12525,N_7093,N_11093);
xor U12526 (N_12526,N_8651,N_8085);
and U12527 (N_12527,N_6178,N_10705);
or U12528 (N_12528,N_6847,N_6236);
and U12529 (N_12529,N_11013,N_7395);
nand U12530 (N_12530,N_8889,N_9508);
or U12531 (N_12531,N_11774,N_10011);
nand U12532 (N_12532,N_11348,N_6290);
or U12533 (N_12533,N_11287,N_10748);
and U12534 (N_12534,N_6473,N_8367);
nor U12535 (N_12535,N_8126,N_10944);
nor U12536 (N_12536,N_9034,N_11198);
or U12537 (N_12537,N_7748,N_8021);
and U12538 (N_12538,N_11125,N_9121);
nand U12539 (N_12539,N_10374,N_8098);
and U12540 (N_12540,N_6507,N_6417);
and U12541 (N_12541,N_10023,N_6147);
nand U12542 (N_12542,N_7837,N_7822);
and U12543 (N_12543,N_8199,N_6209);
xor U12544 (N_12544,N_7260,N_7386);
nor U12545 (N_12545,N_6817,N_9839);
or U12546 (N_12546,N_7519,N_7265);
and U12547 (N_12547,N_8388,N_8289);
and U12548 (N_12548,N_10417,N_11720);
nand U12549 (N_12549,N_9055,N_10804);
and U12550 (N_12550,N_8068,N_7456);
and U12551 (N_12551,N_9775,N_11301);
nor U12552 (N_12552,N_6366,N_8555);
or U12553 (N_12553,N_9051,N_8643);
xor U12554 (N_12554,N_8364,N_7192);
or U12555 (N_12555,N_11769,N_11263);
nor U12556 (N_12556,N_6856,N_10652);
and U12557 (N_12557,N_7345,N_7655);
nor U12558 (N_12558,N_11227,N_6201);
nor U12559 (N_12559,N_7467,N_6570);
and U12560 (N_12560,N_7699,N_7631);
or U12561 (N_12561,N_8923,N_11623);
and U12562 (N_12562,N_11178,N_6056);
or U12563 (N_12563,N_11461,N_8252);
or U12564 (N_12564,N_10541,N_6345);
nor U12565 (N_12565,N_8718,N_9202);
xnor U12566 (N_12566,N_10630,N_8519);
nor U12567 (N_12567,N_9000,N_10521);
or U12568 (N_12568,N_11402,N_7902);
xor U12569 (N_12569,N_7131,N_6796);
nor U12570 (N_12570,N_9610,N_7538);
nand U12571 (N_12571,N_9071,N_8575);
and U12572 (N_12572,N_8814,N_10916);
or U12573 (N_12573,N_10410,N_8149);
xor U12574 (N_12574,N_7968,N_11151);
or U12575 (N_12575,N_6406,N_8083);
or U12576 (N_12576,N_11246,N_11282);
and U12577 (N_12577,N_6898,N_9057);
or U12578 (N_12578,N_10498,N_10614);
nor U12579 (N_12579,N_7293,N_6866);
and U12580 (N_12580,N_10068,N_7055);
xor U12581 (N_12581,N_10644,N_11388);
or U12582 (N_12582,N_11175,N_11944);
xnor U12583 (N_12583,N_7593,N_9179);
nand U12584 (N_12584,N_11617,N_7246);
nand U12585 (N_12585,N_7129,N_9760);
and U12586 (N_12586,N_9200,N_8006);
xnor U12587 (N_12587,N_8605,N_10989);
nor U12588 (N_12588,N_8956,N_8843);
and U12589 (N_12589,N_11312,N_11191);
and U12590 (N_12590,N_7661,N_10334);
or U12591 (N_12591,N_11981,N_11255);
nand U12592 (N_12592,N_11346,N_10245);
xnor U12593 (N_12593,N_10054,N_10097);
or U12594 (N_12594,N_7960,N_6878);
or U12595 (N_12595,N_10709,N_10388);
and U12596 (N_12596,N_9783,N_11785);
or U12597 (N_12597,N_10700,N_9650);
nor U12598 (N_12598,N_6261,N_9380);
nand U12599 (N_12599,N_7453,N_8694);
or U12600 (N_12600,N_6729,N_9165);
and U12601 (N_12601,N_11649,N_9243);
and U12602 (N_12602,N_7779,N_8913);
nor U12603 (N_12603,N_7513,N_9832);
nor U12604 (N_12604,N_11891,N_10704);
nor U12605 (N_12605,N_10791,N_7740);
xnor U12606 (N_12606,N_9877,N_9972);
nor U12607 (N_12607,N_7301,N_6690);
nand U12608 (N_12608,N_9005,N_7172);
nand U12609 (N_12609,N_6067,N_7394);
or U12610 (N_12610,N_9968,N_6489);
or U12611 (N_12611,N_10030,N_6122);
and U12612 (N_12612,N_11176,N_11638);
nor U12613 (N_12613,N_6421,N_8569);
or U12614 (N_12614,N_8785,N_7281);
xnor U12615 (N_12615,N_11361,N_10670);
nand U12616 (N_12616,N_8095,N_6602);
nand U12617 (N_12617,N_9187,N_11479);
or U12618 (N_12618,N_7937,N_11527);
nor U12619 (N_12619,N_7445,N_6110);
and U12620 (N_12620,N_10202,N_10632);
nand U12621 (N_12621,N_9077,N_9861);
or U12622 (N_12622,N_9552,N_9673);
nand U12623 (N_12623,N_6374,N_8891);
and U12624 (N_12624,N_10945,N_11127);
or U12625 (N_12625,N_10910,N_11742);
xor U12626 (N_12626,N_10285,N_6463);
xor U12627 (N_12627,N_9479,N_6712);
nor U12628 (N_12628,N_11717,N_8311);
nor U12629 (N_12629,N_8161,N_7392);
or U12630 (N_12630,N_10663,N_11915);
or U12631 (N_12631,N_9534,N_7178);
or U12632 (N_12632,N_10318,N_11515);
nand U12633 (N_12633,N_11221,N_10320);
nor U12634 (N_12634,N_10610,N_8775);
nand U12635 (N_12635,N_10312,N_6551);
xor U12636 (N_12636,N_9296,N_11831);
and U12637 (N_12637,N_7984,N_9145);
and U12638 (N_12638,N_11304,N_8182);
nor U12639 (N_12639,N_7927,N_10047);
and U12640 (N_12640,N_10182,N_6953);
nor U12641 (N_12641,N_6868,N_9204);
xor U12642 (N_12642,N_7166,N_7701);
or U12643 (N_12643,N_10697,N_11463);
nor U12644 (N_12644,N_10188,N_10444);
or U12645 (N_12645,N_10356,N_11215);
nor U12646 (N_12646,N_8358,N_7508);
xnor U12647 (N_12647,N_7894,N_7254);
xnor U12648 (N_12648,N_8266,N_10041);
xor U12649 (N_12649,N_11456,N_8336);
and U12650 (N_12650,N_7011,N_9312);
or U12651 (N_12651,N_8059,N_11635);
nor U12652 (N_12652,N_8308,N_7458);
and U12653 (N_12653,N_6737,N_7570);
and U12654 (N_12654,N_9636,N_10270);
nand U12655 (N_12655,N_9578,N_10237);
nor U12656 (N_12656,N_11106,N_9744);
nand U12657 (N_12657,N_9587,N_9964);
nor U12658 (N_12658,N_11901,N_11300);
nand U12659 (N_12659,N_6974,N_8592);
nand U12660 (N_12660,N_6476,N_11334);
xor U12661 (N_12661,N_10379,N_9286);
or U12662 (N_12662,N_10967,N_10238);
nand U12663 (N_12663,N_11567,N_7174);
nand U12664 (N_12664,N_11024,N_6824);
nand U12665 (N_12665,N_7303,N_11411);
nor U12666 (N_12666,N_9856,N_7294);
nand U12667 (N_12667,N_11534,N_11069);
nor U12668 (N_12668,N_10840,N_6735);
nor U12669 (N_12669,N_6833,N_11959);
nor U12670 (N_12670,N_11903,N_9225);
xor U12671 (N_12671,N_6911,N_6676);
nor U12672 (N_12672,N_7403,N_10653);
and U12673 (N_12673,N_10760,N_7835);
and U12674 (N_12674,N_7463,N_8028);
and U12675 (N_12675,N_7737,N_10737);
and U12676 (N_12676,N_11922,N_8583);
nand U12677 (N_12677,N_9756,N_10115);
and U12678 (N_12678,N_7007,N_8925);
or U12679 (N_12679,N_6725,N_9319);
and U12680 (N_12680,N_8442,N_8382);
or U12681 (N_12681,N_10668,N_6751);
xnor U12682 (N_12682,N_6579,N_7258);
nor U12683 (N_12683,N_7542,N_11996);
nand U12684 (N_12684,N_9748,N_7530);
nand U12685 (N_12685,N_7457,N_11136);
nor U12686 (N_12686,N_7795,N_9019);
and U12687 (N_12687,N_8197,N_9213);
xor U12688 (N_12688,N_11625,N_6795);
nand U12689 (N_12689,N_6009,N_8238);
nand U12690 (N_12690,N_7344,N_9288);
xor U12691 (N_12691,N_10352,N_11760);
nor U12692 (N_12692,N_7195,N_11953);
and U12693 (N_12693,N_7788,N_9044);
and U12694 (N_12694,N_11307,N_6388);
or U12695 (N_12695,N_11209,N_7124);
nand U12696 (N_12696,N_6203,N_11631);
or U12697 (N_12697,N_11963,N_6279);
nand U12698 (N_12698,N_8187,N_10825);
nor U12699 (N_12699,N_11883,N_10545);
nor U12700 (N_12700,N_8912,N_6778);
xnor U12701 (N_12701,N_11657,N_6167);
xor U12702 (N_12702,N_10845,N_10340);
nor U12703 (N_12703,N_6212,N_8419);
xnor U12704 (N_12704,N_8344,N_11884);
nor U12705 (N_12705,N_8809,N_10269);
or U12706 (N_12706,N_6019,N_10301);
and U12707 (N_12707,N_9109,N_11537);
nand U12708 (N_12708,N_11038,N_10084);
xnor U12709 (N_12709,N_6166,N_9502);
nand U12710 (N_12710,N_10656,N_6230);
xor U12711 (N_12711,N_9752,N_9463);
nor U12712 (N_12712,N_7358,N_11403);
nor U12713 (N_12713,N_7596,N_6950);
nor U12714 (N_12714,N_7598,N_10087);
nand U12715 (N_12715,N_8219,N_8894);
nor U12716 (N_12716,N_6043,N_11333);
nor U12717 (N_12717,N_10232,N_7382);
and U12718 (N_12718,N_9353,N_9418);
and U12719 (N_12719,N_7435,N_6949);
or U12720 (N_12720,N_11614,N_8584);
or U12721 (N_12721,N_9693,N_8828);
or U12722 (N_12722,N_11434,N_10852);
xor U12723 (N_12723,N_7566,N_7157);
xnor U12724 (N_12724,N_9433,N_7895);
nor U12725 (N_12725,N_9621,N_11220);
and U12726 (N_12726,N_8122,N_6649);
xnor U12727 (N_12727,N_11378,N_10678);
and U12728 (N_12728,N_10166,N_10970);
nand U12729 (N_12729,N_7670,N_9664);
xor U12730 (N_12730,N_11814,N_8856);
nor U12731 (N_12731,N_11639,N_6312);
xor U12732 (N_12732,N_11618,N_11122);
nor U12733 (N_12733,N_11413,N_6677);
nand U12734 (N_12734,N_11075,N_9420);
xor U12735 (N_12735,N_10685,N_9089);
nor U12736 (N_12736,N_10389,N_9046);
nor U12737 (N_12737,N_8065,N_7306);
nor U12738 (N_12738,N_10775,N_6710);
or U12739 (N_12739,N_6813,N_8071);
and U12740 (N_12740,N_6807,N_8616);
and U12741 (N_12741,N_9284,N_9063);
nor U12742 (N_12742,N_8769,N_11881);
or U12743 (N_12743,N_6941,N_7552);
or U12744 (N_12744,N_9398,N_7089);
nand U12745 (N_12745,N_8051,N_11281);
or U12746 (N_12746,N_7050,N_9309);
nand U12747 (N_12747,N_8072,N_11372);
nand U12748 (N_12748,N_6763,N_10483);
or U12749 (N_12749,N_7409,N_8835);
and U12750 (N_12750,N_7001,N_9504);
xnor U12751 (N_12751,N_7421,N_8998);
xnor U12752 (N_12752,N_10025,N_9224);
and U12753 (N_12753,N_7272,N_10088);
nor U12754 (N_12754,N_6394,N_7815);
xnor U12755 (N_12755,N_10946,N_9127);
nor U12756 (N_12756,N_7081,N_8474);
xor U12757 (N_12757,N_10886,N_7145);
xnor U12758 (N_12758,N_11994,N_11167);
nand U12759 (N_12759,N_7928,N_11551);
nor U12760 (N_12760,N_6344,N_6098);
and U12761 (N_12761,N_6812,N_11673);
and U12762 (N_12762,N_6311,N_11783);
nor U12763 (N_12763,N_10589,N_6957);
nand U12764 (N_12764,N_9402,N_10228);
and U12765 (N_12765,N_10654,N_11357);
or U12766 (N_12766,N_11028,N_7630);
xnor U12767 (N_12767,N_10131,N_8069);
or U12768 (N_12768,N_9129,N_10679);
nor U12769 (N_12769,N_7959,N_11362);
nand U12770 (N_12770,N_11733,N_8293);
nor U12771 (N_12771,N_10622,N_9304);
nor U12772 (N_12772,N_10746,N_11650);
and U12773 (N_12773,N_6534,N_11728);
nor U12774 (N_12774,N_10531,N_10297);
or U12775 (N_12775,N_10261,N_11736);
and U12776 (N_12776,N_11590,N_10336);
xor U12777 (N_12777,N_8459,N_7273);
or U12778 (N_12778,N_9365,N_10347);
nand U12779 (N_12779,N_10588,N_9763);
xnor U12780 (N_12780,N_6150,N_9974);
nor U12781 (N_12781,N_11565,N_9645);
xor U12782 (N_12782,N_6186,N_7319);
nand U12783 (N_12783,N_7480,N_9210);
or U12784 (N_12784,N_6462,N_8376);
nor U12785 (N_12785,N_9898,N_8262);
or U12786 (N_12786,N_10583,N_10142);
or U12787 (N_12787,N_7099,N_9043);
and U12788 (N_12788,N_9040,N_8134);
or U12789 (N_12789,N_10739,N_8640);
and U12790 (N_12790,N_11392,N_11810);
nand U12791 (N_12791,N_9885,N_8638);
nor U12792 (N_12792,N_9531,N_9318);
nor U12793 (N_12793,N_10469,N_7027);
xor U12794 (N_12794,N_9771,N_6865);
and U12795 (N_12795,N_8807,N_6506);
and U12796 (N_12796,N_10997,N_6144);
nand U12797 (N_12797,N_7268,N_7434);
nor U12798 (N_12798,N_8732,N_8499);
and U12799 (N_12799,N_8660,N_7577);
xnor U12800 (N_12800,N_11152,N_11722);
and U12801 (N_12801,N_10196,N_6397);
nand U12802 (N_12802,N_9235,N_10494);
nor U12803 (N_12803,N_9015,N_6985);
and U12804 (N_12804,N_11259,N_9766);
nor U12805 (N_12805,N_6416,N_9259);
xnor U12806 (N_12806,N_11611,N_9689);
or U12807 (N_12807,N_7353,N_10412);
nand U12808 (N_12808,N_10543,N_10565);
nor U12809 (N_12809,N_7705,N_9347);
and U12810 (N_12810,N_8533,N_9720);
and U12811 (N_12811,N_8965,N_10451);
nand U12812 (N_12812,N_8798,N_8395);
nand U12813 (N_12813,N_7278,N_10138);
nand U12814 (N_12814,N_6245,N_10122);
xnor U12815 (N_12815,N_10585,N_6425);
nor U12816 (N_12816,N_11671,N_7755);
or U12817 (N_12817,N_9407,N_10787);
xor U12818 (N_12818,N_6386,N_11148);
or U12819 (N_12819,N_7008,N_6513);
and U12820 (N_12820,N_9444,N_9945);
or U12821 (N_12821,N_8778,N_8512);
xor U12822 (N_12822,N_10126,N_9172);
or U12823 (N_12823,N_9707,N_7493);
or U12824 (N_12824,N_7680,N_8750);
and U12825 (N_12825,N_10043,N_8480);
or U12826 (N_12826,N_6249,N_6340);
and U12827 (N_12827,N_7186,N_11909);
nand U12828 (N_12828,N_6010,N_9201);
or U12829 (N_12829,N_7035,N_11134);
nor U12830 (N_12830,N_7479,N_9894);
nand U12831 (N_12831,N_8668,N_11352);
nand U12832 (N_12832,N_7085,N_11843);
nor U12833 (N_12833,N_11770,N_8475);
nor U12834 (N_12834,N_11985,N_11569);
xor U12835 (N_12835,N_6923,N_9916);
and U12836 (N_12836,N_11047,N_8536);
and U12837 (N_12837,N_10712,N_6414);
nand U12838 (N_12838,N_7245,N_9382);
xor U12839 (N_12839,N_9049,N_10449);
or U12840 (N_12840,N_6637,N_10380);
or U12841 (N_12841,N_11071,N_6027);
and U12842 (N_12842,N_7903,N_11495);
and U12843 (N_12843,N_9666,N_7127);
xor U12844 (N_12844,N_6907,N_6713);
and U12845 (N_12845,N_11588,N_11856);
or U12846 (N_12846,N_8805,N_11313);
xor U12847 (N_12847,N_8818,N_8899);
nand U12848 (N_12848,N_8162,N_10338);
nor U12849 (N_12849,N_7782,N_9820);
or U12850 (N_12850,N_11613,N_9107);
nand U12851 (N_12851,N_10633,N_7692);
or U12852 (N_12852,N_11144,N_10755);
xnor U12853 (N_12853,N_6083,N_6136);
nor U12854 (N_12854,N_9404,N_9669);
nand U12855 (N_12855,N_8280,N_10448);
and U12856 (N_12856,N_6156,N_7484);
xor U12857 (N_12857,N_9724,N_10592);
and U12858 (N_12858,N_11443,N_8368);
xnor U12859 (N_12859,N_10820,N_6478);
or U12860 (N_12860,N_6530,N_10103);
or U12861 (N_12861,N_6004,N_10106);
or U12862 (N_12862,N_7647,N_10108);
or U12863 (N_12863,N_11767,N_8985);
and U12864 (N_12864,N_7995,N_11931);
xor U12865 (N_12865,N_10484,N_8271);
nor U12866 (N_12866,N_11947,N_8325);
or U12867 (N_12867,N_11488,N_7418);
and U12868 (N_12868,N_11286,N_8112);
or U12869 (N_12869,N_6784,N_11586);
xnor U12870 (N_12870,N_7133,N_7710);
xor U12871 (N_12871,N_8230,N_10052);
xor U12872 (N_12872,N_7607,N_6265);
or U12873 (N_12873,N_8982,N_7799);
or U12874 (N_12874,N_6919,N_9162);
or U12875 (N_12875,N_9052,N_8343);
nor U12876 (N_12876,N_10606,N_9108);
and U12877 (N_12877,N_11088,N_6999);
xor U12878 (N_12878,N_7994,N_9950);
nand U12879 (N_12879,N_11570,N_11223);
or U12880 (N_12880,N_10402,N_9460);
nand U12881 (N_12881,N_11820,N_8591);
nor U12882 (N_12882,N_9171,N_6955);
nor U12883 (N_12883,N_9701,N_10682);
xor U12884 (N_12884,N_10158,N_7476);
nand U12885 (N_12885,N_6223,N_11076);
or U12886 (N_12886,N_6643,N_9156);
nor U12887 (N_12887,N_6753,N_6264);
xnor U12888 (N_12888,N_7452,N_9795);
and U12889 (N_12889,N_6822,N_7940);
nand U12890 (N_12890,N_8620,N_10693);
xnor U12891 (N_12891,N_8786,N_11779);
or U12892 (N_12892,N_10873,N_6909);
and U12893 (N_12893,N_7856,N_7384);
nand U12894 (N_12894,N_11323,N_11482);
xor U12895 (N_12895,N_9002,N_8992);
xor U12896 (N_12896,N_8427,N_10940);
or U12897 (N_12897,N_9472,N_7399);
xor U12898 (N_12898,N_11244,N_11797);
xor U12899 (N_12899,N_6662,N_7610);
xor U12900 (N_12900,N_8866,N_11676);
nor U12901 (N_12901,N_10659,N_10313);
or U12902 (N_12902,N_7950,N_9927);
nor U12903 (N_12903,N_8283,N_10181);
nor U12904 (N_12904,N_8905,N_11758);
or U12905 (N_12905,N_6349,N_6277);
nand U12906 (N_12906,N_11707,N_11529);
and U12907 (N_12907,N_7231,N_10242);
and U12908 (N_12908,N_11859,N_10683);
and U12909 (N_12909,N_8256,N_9728);
or U12910 (N_12910,N_8167,N_7209);
and U12911 (N_12911,N_9011,N_10033);
nor U12912 (N_12912,N_11320,N_10662);
and U12913 (N_12913,N_6495,N_10191);
or U12914 (N_12914,N_10136,N_7140);
xor U12915 (N_12915,N_11775,N_6106);
or U12916 (N_12916,N_9849,N_8415);
nor U12917 (N_12917,N_6158,N_11860);
and U12918 (N_12918,N_6327,N_9359);
nand U12919 (N_12919,N_9739,N_10853);
or U12920 (N_12920,N_9796,N_10457);
nand U12921 (N_12921,N_10058,N_6299);
and U12922 (N_12922,N_8261,N_11389);
xor U12923 (N_12923,N_7296,N_8397);
xor U12924 (N_12924,N_6224,N_7898);
or U12925 (N_12925,N_10441,N_6208);
or U12926 (N_12926,N_8150,N_10556);
xnor U12927 (N_12927,N_6655,N_10477);
or U12928 (N_12928,N_11202,N_11751);
xnor U12929 (N_12929,N_7651,N_7876);
nand U12930 (N_12930,N_11358,N_6604);
or U12931 (N_12931,N_8665,N_6013);
xnor U12932 (N_12932,N_10520,N_11520);
nor U12933 (N_12933,N_11385,N_11878);
xnor U12934 (N_12934,N_10480,N_7080);
or U12935 (N_12935,N_10888,N_6862);
nor U12936 (N_12936,N_9369,N_6430);
nor U12937 (N_12937,N_10497,N_9743);
nor U12938 (N_12938,N_11022,N_9021);
nand U12939 (N_12939,N_6479,N_8909);
nand U12940 (N_12940,N_6947,N_8196);
and U12941 (N_12941,N_10061,N_10393);
or U12942 (N_12942,N_11718,N_7711);
and U12943 (N_12943,N_7332,N_9450);
xor U12944 (N_12944,N_7523,N_6017);
and U12945 (N_12945,N_10836,N_6181);
or U12946 (N_12946,N_11633,N_9640);
xnor U12947 (N_12947,N_9825,N_9203);
or U12948 (N_12948,N_11910,N_10869);
xor U12949 (N_12949,N_6899,N_10968);
nand U12950 (N_12950,N_10369,N_7580);
nor U12951 (N_12951,N_8635,N_10258);
nor U12952 (N_12952,N_10263,N_10117);
xnor U12953 (N_12953,N_6233,N_11827);
or U12954 (N_12954,N_9428,N_9711);
and U12955 (N_12955,N_8141,N_11252);
xnor U12956 (N_12956,N_11179,N_10293);
nand U12957 (N_12957,N_7051,N_10350);
or U12958 (N_12958,N_10762,N_6660);
nand U12959 (N_12959,N_7586,N_7674);
nand U12960 (N_12960,N_11477,N_8237);
and U12961 (N_12961,N_6672,N_10169);
nor U12962 (N_12962,N_10294,N_6773);
nor U12963 (N_12963,N_8337,N_9676);
nor U12964 (N_12964,N_9069,N_8111);
nand U12965 (N_12965,N_11296,N_11240);
nand U12966 (N_12966,N_7955,N_11874);
or U12967 (N_12967,N_10859,N_8079);
xnor U12968 (N_12968,N_9181,N_9816);
and U12969 (N_12969,N_9564,N_7087);
or U12970 (N_12970,N_11498,N_11438);
or U12971 (N_12971,N_9794,N_8852);
and U12972 (N_12972,N_10830,N_11939);
nor U12973 (N_12973,N_7488,N_9602);
or U12974 (N_12974,N_6917,N_6702);
or U12975 (N_12975,N_11738,N_7745);
nand U12976 (N_12976,N_11543,N_11982);
and U12977 (N_12977,N_10145,N_9691);
nor U12978 (N_12978,N_10260,N_9385);
and U12979 (N_12979,N_8737,N_8825);
or U12980 (N_12980,N_11436,N_11935);
xor U12981 (N_12981,N_10413,N_10719);
nor U12982 (N_12982,N_11908,N_8936);
nand U12983 (N_12983,N_8375,N_8653);
and U12984 (N_12984,N_10832,N_8168);
xor U12985 (N_12985,N_7311,N_7949);
nor U12986 (N_12986,N_9485,N_10774);
or U12987 (N_12987,N_10094,N_10133);
nor U12988 (N_12988,N_10360,N_7991);
or U12989 (N_12989,N_6827,N_6970);
nand U12990 (N_12990,N_6500,N_11957);
and U12991 (N_12991,N_11572,N_8231);
or U12992 (N_12992,N_8438,N_9882);
nand U12993 (N_12993,N_10081,N_10641);
nand U12994 (N_12994,N_11328,N_6225);
xor U12995 (N_12995,N_11726,N_10717);
and U12996 (N_12996,N_7017,N_7039);
nor U12997 (N_12997,N_7071,N_10007);
nor U12998 (N_12998,N_10642,N_6141);
and U12999 (N_12999,N_9831,N_11111);
xor U13000 (N_13000,N_7658,N_9360);
nand U13001 (N_13001,N_7054,N_8783);
and U13002 (N_13002,N_6587,N_9513);
nand U13003 (N_13003,N_9008,N_11309);
xor U13004 (N_13004,N_8630,N_6252);
and U13005 (N_13005,N_9930,N_9883);
and U13006 (N_13006,N_6169,N_10365);
nor U13007 (N_13007,N_6196,N_8027);
nand U13008 (N_13008,N_7320,N_8708);
and U13009 (N_13009,N_8054,N_9379);
and U13010 (N_13010,N_8444,N_7609);
or U13011 (N_13011,N_6906,N_6355);
or U13012 (N_13012,N_9298,N_10006);
xor U13013 (N_13013,N_11092,N_9105);
xnor U13014 (N_13014,N_11858,N_11232);
nor U13015 (N_13015,N_8041,N_8208);
nor U13016 (N_13016,N_9588,N_9456);
and U13017 (N_13017,N_11051,N_7569);
xnor U13018 (N_13018,N_11696,N_8873);
nand U13019 (N_13019,N_7832,N_7191);
nand U13020 (N_13020,N_8906,N_7160);
nand U13021 (N_13021,N_10016,N_10751);
xnor U13022 (N_13022,N_6447,N_9436);
nor U13023 (N_13023,N_11141,N_7760);
and U13024 (N_13024,N_11877,N_6274);
and U13025 (N_13025,N_6029,N_8067);
xor U13026 (N_13026,N_8646,N_11594);
and U13027 (N_13027,N_10208,N_8801);
nand U13028 (N_13028,N_6445,N_7582);
nor U13029 (N_13029,N_6154,N_6280);
xor U13030 (N_13030,N_10109,N_11342);
or U13031 (N_13031,N_11979,N_10909);
or U13032 (N_13032,N_7814,N_6925);
and U13033 (N_13033,N_6372,N_10645);
nor U13034 (N_13034,N_11462,N_11674);
and U13035 (N_13035,N_9190,N_9800);
nand U13036 (N_13036,N_11899,N_6362);
nand U13037 (N_13037,N_10922,N_6063);
xor U13038 (N_13038,N_8064,N_7964);
and U13039 (N_13039,N_6011,N_9614);
nor U13040 (N_13040,N_8062,N_9091);
or U13041 (N_13041,N_9947,N_10291);
xnor U13042 (N_13042,N_6968,N_10012);
xor U13043 (N_13043,N_6302,N_7823);
and U13044 (N_13044,N_10937,N_11672);
and U13045 (N_13045,N_8247,N_6076);
or U13046 (N_13046,N_11061,N_8441);
or U13047 (N_13047,N_11782,N_8496);
nor U13048 (N_13048,N_8931,N_7112);
and U13049 (N_13049,N_11552,N_9944);
or U13050 (N_13050,N_8577,N_9854);
xnor U13051 (N_13051,N_6895,N_7684);
nand U13052 (N_13052,N_7362,N_9841);
nor U13053 (N_13053,N_6138,N_7603);
nor U13054 (N_13054,N_7656,N_6168);
nand U13055 (N_13055,N_8974,N_7956);
and U13056 (N_13056,N_7614,N_8436);
or U13057 (N_13057,N_10924,N_8144);
xnor U13058 (N_13058,N_10014,N_9642);
nand U13059 (N_13059,N_7156,N_7590);
or U13060 (N_13060,N_9985,N_7628);
nand U13061 (N_13061,N_6329,N_10078);
nor U13062 (N_13062,N_9594,N_6552);
nor U13063 (N_13063,N_6932,N_11546);
nand U13064 (N_13064,N_9667,N_8276);
nand U13065 (N_13065,N_10153,N_10325);
nor U13066 (N_13066,N_10231,N_9250);
nor U13067 (N_13067,N_11587,N_10514);
and U13068 (N_13068,N_11969,N_11521);
xnor U13069 (N_13069,N_7930,N_9540);
nor U13070 (N_13070,N_9970,N_6396);
xnor U13071 (N_13071,N_6298,N_7064);
and U13072 (N_13072,N_6592,N_6651);
or U13073 (N_13073,N_9120,N_9245);
nor U13074 (N_13074,N_8504,N_6928);
xor U13075 (N_13075,N_11872,N_8295);
nor U13076 (N_13076,N_10735,N_7009);
nor U13077 (N_13077,N_7208,N_9567);
nor U13078 (N_13078,N_10066,N_11988);
and U13079 (N_13079,N_10549,N_7108);
xor U13080 (N_13080,N_6405,N_10740);
or U13081 (N_13081,N_8984,N_8472);
xor U13082 (N_13082,N_8684,N_11395);
nand U13083 (N_13083,N_6829,N_6636);
and U13084 (N_13084,N_9453,N_6971);
and U13085 (N_13085,N_7426,N_10881);
or U13086 (N_13086,N_11932,N_7840);
nand U13087 (N_13087,N_11522,N_11072);
and U13088 (N_13088,N_6555,N_9147);
and U13089 (N_13089,N_6128,N_8650);
nand U13090 (N_13090,N_10304,N_7269);
nor U13091 (N_13091,N_7739,N_8487);
xnor U13092 (N_13092,N_7059,N_7119);
nor U13093 (N_13093,N_8232,N_7499);
and U13094 (N_13094,N_6313,N_7365);
xnor U13095 (N_13095,N_10256,N_11427);
nor U13096 (N_13096,N_8549,N_7274);
nand U13097 (N_13097,N_8787,N_6701);
nor U13098 (N_13098,N_8473,N_10956);
and U13099 (N_13099,N_7347,N_9590);
or U13100 (N_13100,N_6436,N_6595);
nor U13101 (N_13101,N_7276,N_9176);
nor U13102 (N_13102,N_10876,N_10727);
xor U13103 (N_13103,N_8663,N_10698);
xor U13104 (N_13104,N_11539,N_11949);
xor U13105 (N_13105,N_11640,N_6650);
nor U13106 (N_13106,N_11692,N_6764);
and U13107 (N_13107,N_8506,N_11665);
xor U13108 (N_13108,N_10164,N_9753);
and U13109 (N_13109,N_11397,N_10079);
and U13110 (N_13110,N_9846,N_10948);
nand U13111 (N_13111,N_10240,N_9685);
or U13112 (N_13112,N_6734,N_6600);
xnor U13113 (N_13113,N_9038,N_6563);
nor U13114 (N_13114,N_9782,N_9346);
and U13115 (N_13115,N_10284,N_10788);
xnor U13116 (N_13116,N_7723,N_7932);
nor U13117 (N_13117,N_8991,N_7909);
or U13118 (N_13118,N_8961,N_10624);
xor U13119 (N_13119,N_9867,N_8972);
xnor U13120 (N_13120,N_8015,N_8664);
nand U13121 (N_13121,N_10298,N_8730);
xnor U13122 (N_13122,N_8032,N_7581);
nand U13123 (N_13123,N_11556,N_9612);
or U13124 (N_13124,N_11548,N_8859);
nor U13125 (N_13125,N_9373,N_7432);
or U13126 (N_13126,N_10637,N_8383);
nor U13127 (N_13127,N_6688,N_7766);
nor U13128 (N_13128,N_7369,N_11407);
and U13129 (N_13129,N_11070,N_9186);
xor U13130 (N_13130,N_6086,N_7889);
nand U13131 (N_13131,N_10752,N_11349);
nor U13132 (N_13132,N_10031,N_8847);
nand U13133 (N_13133,N_8544,N_7979);
nand U13134 (N_13134,N_9769,N_11849);
nand U13135 (N_13135,N_6709,N_6457);
or U13136 (N_13136,N_9599,N_6765);
nand U13137 (N_13137,N_8752,N_6428);
nand U13138 (N_13138,N_7883,N_11502);
nand U13139 (N_13139,N_8932,N_10797);
nand U13140 (N_13140,N_6739,N_8003);
xor U13141 (N_13141,N_8296,N_6874);
xor U13142 (N_13142,N_9491,N_8225);
or U13143 (N_13143,N_9490,N_7412);
nor U13144 (N_13144,N_7144,N_8606);
or U13145 (N_13145,N_6837,N_7880);
nor U13146 (N_13146,N_8175,N_8634);
nor U13147 (N_13147,N_11535,N_11584);
nand U13148 (N_13148,N_11452,N_8173);
xnor U13149 (N_13149,N_7768,N_8983);
xor U13150 (N_13150,N_9150,N_10801);
or U13151 (N_13151,N_10487,N_7522);
nor U13152 (N_13152,N_9637,N_11412);
xnor U13153 (N_13153,N_7971,N_7546);
xnor U13154 (N_13154,N_8841,N_10568);
and U13155 (N_13155,N_6673,N_9873);
and U13156 (N_13156,N_9757,N_6746);
nand U13157 (N_13157,N_7261,N_9081);
xnor U13158 (N_13158,N_7401,N_6920);
and U13159 (N_13159,N_6439,N_8125);
or U13160 (N_13160,N_10550,N_10343);
xor U13161 (N_13161,N_7987,N_8088);
and U13162 (N_13162,N_6057,N_7324);
and U13163 (N_13163,N_10251,N_7846);
xor U13164 (N_13164,N_9630,N_9016);
or U13165 (N_13165,N_10570,N_11978);
nand U13166 (N_13166,N_6861,N_11697);
nand U13167 (N_13167,N_10838,N_6605);
and U13168 (N_13168,N_8976,N_10795);
xnor U13169 (N_13169,N_10059,N_9223);
xor U13170 (N_13170,N_7371,N_6074);
xor U13171 (N_13171,N_8896,N_7521);
nand U13172 (N_13172,N_11918,N_11420);
and U13173 (N_13173,N_7010,N_8907);
and U13174 (N_13174,N_9262,N_7096);
nand U13175 (N_13175,N_7974,N_8279);
and U13176 (N_13176,N_10355,N_9149);
nand U13177 (N_13177,N_7134,N_8155);
nor U13178 (N_13178,N_10384,N_11045);
nor U13179 (N_13179,N_10461,N_6929);
nand U13180 (N_13180,N_10868,N_8568);
nor U13181 (N_13181,N_9990,N_8009);
nand U13182 (N_13182,N_6526,N_7811);
or U13183 (N_13183,N_8359,N_8746);
nand U13184 (N_13184,N_11485,N_11410);
xor U13185 (N_13185,N_8087,N_6336);
nand U13186 (N_13186,N_7700,N_8753);
or U13187 (N_13187,N_9657,N_9687);
nand U13188 (N_13188,N_10414,N_8587);
nor U13189 (N_13189,N_11332,N_11005);
xor U13190 (N_13190,N_10815,N_7496);
and U13191 (N_13191,N_7859,N_10471);
and U13192 (N_13192,N_6045,N_9696);
or U13193 (N_13193,N_8099,N_10366);
and U13194 (N_13194,N_10385,N_7004);
and U13195 (N_13195,N_11336,N_9708);
or U13196 (N_13196,N_7568,N_6403);
and U13197 (N_13197,N_8392,N_8834);
nor U13198 (N_13198,N_6914,N_6613);
and U13199 (N_13199,N_9677,N_8131);
or U13200 (N_13200,N_6146,N_11714);
nand U13201 (N_13201,N_7420,N_10307);
nor U13202 (N_13202,N_10731,N_10745);
xnor U13203 (N_13203,N_7943,N_8462);
and U13204 (N_13204,N_8482,N_8999);
or U13205 (N_13205,N_9278,N_11486);
nor U13206 (N_13206,N_6047,N_10060);
nor U13207 (N_13207,N_8552,N_11916);
nor U13208 (N_13208,N_10481,N_11353);
nor U13209 (N_13209,N_11771,N_8926);
or U13210 (N_13210,N_8316,N_8172);
xor U13211 (N_13211,N_11229,N_8153);
nor U13212 (N_13212,N_8390,N_8347);
nand U13213 (N_13213,N_8394,N_9389);
and U13214 (N_13214,N_7704,N_7619);
xor U13215 (N_13215,N_9611,N_6572);
or U13216 (N_13216,N_10478,N_6112);
or U13217 (N_13217,N_10370,N_8102);
xor U13218 (N_13218,N_6578,N_8380);
nand U13219 (N_13219,N_6731,N_9603);
and U13220 (N_13220,N_6227,N_11817);
xor U13221 (N_13221,N_6492,N_8721);
nand U13222 (N_13222,N_11204,N_6680);
nor U13223 (N_13223,N_10805,N_6253);
nand U13224 (N_13224,N_11279,N_6565);
or U13225 (N_13225,N_10707,N_8829);
or U13226 (N_13226,N_11484,N_6301);
xor U13227 (N_13227,N_11690,N_6897);
nor U13228 (N_13228,N_7012,N_11906);
nor U13229 (N_13229,N_7424,N_8221);
nor U13230 (N_13230,N_6556,N_6873);
nand U13231 (N_13231,N_6330,N_9686);
nand U13232 (N_13232,N_7110,N_11683);
or U13233 (N_13233,N_10045,N_8460);
or U13234 (N_13234,N_10926,N_9802);
and U13235 (N_13235,N_9570,N_8117);
or U13236 (N_13236,N_11764,N_11904);
xnor U13237 (N_13237,N_11977,N_11369);
nand U13238 (N_13238,N_11787,N_11554);
nand U13239 (N_13239,N_10903,N_9864);
nor U13240 (N_13240,N_8768,N_7073);
or U13241 (N_13241,N_7517,N_6435);
and U13242 (N_13242,N_6471,N_9559);
or U13243 (N_13243,N_7564,N_7151);
nor U13244 (N_13244,N_9890,N_9779);
nor U13245 (N_13245,N_7543,N_6251);
nor U13246 (N_13246,N_6443,N_7176);
xnor U13247 (N_13247,N_8946,N_7604);
nor U13248 (N_13248,N_9215,N_6410);
nand U13249 (N_13249,N_7491,N_9264);
and U13250 (N_13250,N_9988,N_10227);
nand U13251 (N_13251,N_11970,N_9525);
and U13252 (N_13252,N_9447,N_7676);
or U13253 (N_13253,N_11777,N_10949);
nor U13254 (N_13254,N_10833,N_7634);
or U13255 (N_13255,N_11382,N_8970);
nor U13256 (N_13256,N_9577,N_9682);
and U13257 (N_13257,N_10692,N_10779);
xnor U13258 (N_13258,N_11999,N_9362);
or U13259 (N_13259,N_8073,N_11643);
nand U13260 (N_13260,N_11976,N_10440);
nor U13261 (N_13261,N_8557,N_10824);
and U13262 (N_13262,N_6816,N_6361);
or U13263 (N_13263,N_11740,N_9761);
and U13264 (N_13264,N_8717,N_6509);
or U13265 (N_13265,N_6591,N_8461);
or U13266 (N_13266,N_6863,N_10496);
xor U13267 (N_13267,N_8093,N_11841);
and U13268 (N_13268,N_11265,N_8819);
and U13269 (N_13269,N_11500,N_9982);
nor U13270 (N_13270,N_7575,N_7255);
or U13271 (N_13271,N_9395,N_10249);
xor U13272 (N_13272,N_10616,N_10134);
nand U13273 (N_13273,N_10686,N_6294);
or U13274 (N_13274,N_11991,N_8007);
nand U13275 (N_13275,N_6465,N_11804);
nand U13276 (N_13276,N_6173,N_10785);
or U13277 (N_13277,N_7334,N_8114);
and U13278 (N_13278,N_8483,N_7339);
and U13279 (N_13279,N_7308,N_11888);
or U13280 (N_13280,N_6046,N_6791);
nor U13281 (N_13281,N_10515,N_6314);
xor U13282 (N_13282,N_11023,N_10680);
or U13283 (N_13283,N_9432,N_8002);
nand U13284 (N_13284,N_10368,N_6547);
xnor U13285 (N_13285,N_9575,N_8877);
xor U13286 (N_13286,N_7531,N_6619);
nand U13287 (N_13287,N_11035,N_8507);
nor U13288 (N_13288,N_9635,N_6836);
or U13289 (N_13289,N_11062,N_11659);
and U13290 (N_13290,N_11836,N_7152);
nand U13291 (N_13291,N_8070,N_9902);
and U13292 (N_13292,N_7288,N_9773);
and U13293 (N_13293,N_9421,N_10716);
and U13294 (N_13294,N_7707,N_8268);
xor U13295 (N_13295,N_11781,N_7214);
nor U13296 (N_13296,N_10288,N_11709);
xnor U13297 (N_13297,N_11472,N_9206);
nand U13298 (N_13298,N_7061,N_6821);
nor U13299 (N_13299,N_6566,N_8949);
xnor U13300 (N_13300,N_6393,N_11511);
and U13301 (N_13301,N_6859,N_10586);
xor U13302 (N_13302,N_8145,N_6072);
or U13303 (N_13303,N_7460,N_10880);
nand U13304 (N_13304,N_8846,N_8599);
xnor U13305 (N_13305,N_11776,N_7221);
nor U13306 (N_13306,N_6239,N_11648);
nand U13307 (N_13307,N_9639,N_9583);
xnor U13308 (N_13308,N_10582,N_10988);
nor U13309 (N_13309,N_11933,N_10364);
or U13310 (N_13310,N_10872,N_11923);
nor U13311 (N_13311,N_11589,N_8990);
nor U13312 (N_13312,N_6331,N_6023);
xor U13313 (N_13313,N_8875,N_10185);
nand U13314 (N_13314,N_7448,N_6258);
nor U13315 (N_13315,N_7153,N_11658);
xnor U13316 (N_13316,N_6926,N_10931);
nand U13317 (N_13317,N_11355,N_11880);
or U13318 (N_13318,N_7033,N_9411);
or U13319 (N_13319,N_6161,N_7642);
xnor U13320 (N_13320,N_11087,N_10349);
or U13321 (N_13321,N_10257,N_9989);
and U13322 (N_13322,N_8683,N_6903);
nor U13323 (N_13323,N_10907,N_9140);
xor U13324 (N_13324,N_6281,N_6219);
xor U13325 (N_13325,N_10400,N_11757);
or U13326 (N_13326,N_9117,N_9257);
and U13327 (N_13327,N_7841,N_8522);
or U13328 (N_13328,N_8422,N_8185);
nor U13329 (N_13329,N_6191,N_9412);
and U13330 (N_13330,N_8670,N_10399);
nor U13331 (N_13331,N_8485,N_8400);
xor U13332 (N_13332,N_8797,N_7163);
or U13333 (N_13333,N_8479,N_9492);
xor U13334 (N_13334,N_9335,N_6278);
and U13335 (N_13335,N_6069,N_7908);
and U13336 (N_13336,N_10947,N_11324);
and U13337 (N_13337,N_6379,N_6176);
and U13338 (N_13338,N_10102,N_11663);
xnor U13339 (N_13339,N_10149,N_11481);
nand U13340 (N_13340,N_11055,N_7407);
or U13341 (N_13341,N_11668,N_6933);
xor U13342 (N_13342,N_10063,N_8884);
and U13343 (N_13343,N_9193,N_7251);
nand U13344 (N_13344,N_7874,N_11700);
and U13345 (N_13345,N_9484,N_7390);
xor U13346 (N_13346,N_8541,N_7444);
or U13347 (N_13347,N_7809,N_9422);
or U13348 (N_13348,N_10580,N_10308);
or U13349 (N_13349,N_9310,N_9125);
or U13350 (N_13350,N_9758,N_10839);
xnor U13351 (N_13351,N_9455,N_11971);
xor U13352 (N_13352,N_6982,N_9295);
or U13353 (N_13353,N_10029,N_10893);
nor U13354 (N_13354,N_6995,N_11090);
xnor U13355 (N_13355,N_11146,N_8012);
xor U13356 (N_13356,N_6211,N_7118);
nand U13357 (N_13357,N_8404,N_11627);
and U13358 (N_13358,N_6308,N_11011);
nor U13359 (N_13359,N_10862,N_7213);
or U13360 (N_13360,N_10736,N_7113);
nand U13361 (N_13361,N_10376,N_10964);
or U13362 (N_13362,N_11517,N_7271);
nor U13363 (N_13363,N_6618,N_11964);
nand U13364 (N_13364,N_6826,N_8330);
xnor U13365 (N_13365,N_6629,N_11616);
nand U13366 (N_13366,N_7703,N_11794);
nand U13367 (N_13367,N_11404,N_10178);
or U13368 (N_13368,N_9263,N_6026);
nor U13369 (N_13369,N_6626,N_6133);
nor U13370 (N_13370,N_9817,N_10010);
or U13371 (N_13371,N_7132,N_6993);
xnor U13372 (N_13372,N_8622,N_9498);
nor U13373 (N_13373,N_9617,N_11563);
nand U13374 (N_13374,N_8342,N_6973);
xnor U13375 (N_13375,N_8110,N_6972);
or U13376 (N_13376,N_6769,N_10879);
or U13377 (N_13377,N_11102,N_6691);
or U13378 (N_13378,N_7355,N_8611);
or U13379 (N_13379,N_10170,N_7896);
and U13380 (N_13380,N_9073,N_7111);
xnor U13381 (N_13381,N_7492,N_10303);
nand U13382 (N_13382,N_7021,N_6840);
xnor U13383 (N_13383,N_11842,N_6732);
or U13384 (N_13384,N_11945,N_8602);
xor U13385 (N_13385,N_8408,N_6781);
nor U13386 (N_13386,N_6254,N_10563);
nor U13387 (N_13387,N_6639,N_9609);
and U13388 (N_13388,N_10454,N_11791);
or U13389 (N_13389,N_10861,N_6521);
and U13390 (N_13390,N_9835,N_6901);
or U13391 (N_13391,N_9997,N_7643);
or U13392 (N_13392,N_7413,N_10137);
or U13393 (N_13393,N_8324,N_11636);
xnor U13394 (N_13394,N_7873,N_9683);
nand U13395 (N_13395,N_7560,N_7731);
or U13396 (N_13396,N_7206,N_11601);
nand U13397 (N_13397,N_6562,N_9819);
nand U13398 (N_13398,N_11750,N_10687);
and U13399 (N_13399,N_10500,N_11226);
nand U13400 (N_13400,N_8779,N_6317);
nand U13401 (N_13401,N_8893,N_11063);
nand U13402 (N_13402,N_8734,N_7534);
or U13403 (N_13403,N_11509,N_6728);
nand U13404 (N_13404,N_7591,N_10936);
and U13405 (N_13405,N_11536,N_7899);
nor U13406 (N_13406,N_9454,N_9934);
and U13407 (N_13407,N_10763,N_9542);
or U13408 (N_13408,N_11120,N_6103);
xor U13409 (N_13409,N_11902,N_10093);
nor U13410 (N_13410,N_9791,N_11086);
xnor U13411 (N_13411,N_8678,N_10502);
nor U13412 (N_13412,N_7746,N_7230);
xnor U13413 (N_13413,N_9157,N_7146);
or U13414 (N_13414,N_7535,N_11746);
xor U13415 (N_13415,N_9275,N_10160);
or U13416 (N_13416,N_7207,N_10667);
and U13417 (N_13417,N_6014,N_6139);
and U13418 (N_13418,N_6357,N_9252);
or U13419 (N_13419,N_11124,N_9476);
xor U13420 (N_13420,N_11153,N_6759);
or U13421 (N_13421,N_7533,N_6598);
and U13422 (N_13422,N_11597,N_11667);
and U13423 (N_13423,N_9247,N_10299);
nor U13424 (N_13424,N_6975,N_6633);
or U13425 (N_13425,N_8820,N_6541);
or U13426 (N_13426,N_8876,N_9135);
nor U13427 (N_13427,N_6638,N_8254);
or U13428 (N_13428,N_8751,N_10703);
nor U13429 (N_13429,N_7286,N_10335);
nor U13430 (N_13430,N_6097,N_10536);
or U13431 (N_13431,N_11622,N_6016);
xnor U13432 (N_13432,N_6342,N_7877);
nand U13433 (N_13433,N_7130,N_6268);
nor U13434 (N_13434,N_6656,N_11424);
or U13435 (N_13435,N_9410,N_9452);
nor U13436 (N_13436,N_10143,N_11476);
nor U13437 (N_13437,N_7283,N_9188);
nor U13438 (N_13438,N_10396,N_7031);
nor U13439 (N_13439,N_9112,N_8973);
and U13440 (N_13440,N_7028,N_6434);
nor U13441 (N_13441,N_10547,N_7812);
xor U13442 (N_13442,N_7675,N_10526);
nand U13443 (N_13443,N_9208,N_11449);
and U13444 (N_13444,N_8542,N_8240);
or U13445 (N_13445,N_7338,N_6979);
nor U13446 (N_13446,N_9852,N_8195);
nand U13447 (N_13447,N_10226,N_11950);
nand U13448 (N_13448,N_11465,N_9884);
and U13449 (N_13449,N_7121,N_7944);
nand U13450 (N_13450,N_9745,N_11889);
nand U13451 (N_13451,N_9065,N_11468);
nand U13452 (N_13452,N_8170,N_10778);
nor U13453 (N_13453,N_7168,N_7224);
xnor U13454 (N_13454,N_10219,N_11608);
and U13455 (N_13455,N_11168,N_7257);
and U13456 (N_13456,N_9823,N_8593);
xnor U13457 (N_13457,N_7789,N_11007);
xnor U13458 (N_13458,N_7002,N_11754);
nor U13459 (N_13459,N_9390,N_8214);
nor U13460 (N_13460,N_6218,N_8934);
nand U13461 (N_13461,N_11662,N_11095);
nor U13462 (N_13462,N_11406,N_6429);
nand U13463 (N_13463,N_6064,N_11039);
nand U13464 (N_13464,N_6272,N_7256);
or U13465 (N_13465,N_9726,N_7720);
nand U13466 (N_13466,N_10253,N_9468);
nand U13467 (N_13467,N_10378,N_9207);
and U13468 (N_13468,N_7972,N_9138);
xor U13469 (N_13469,N_10070,N_9889);
xnor U13470 (N_13470,N_7181,N_8350);
nor U13471 (N_13471,N_11189,N_8306);
xnor U13472 (N_13472,N_11302,N_11164);
nand U13473 (N_13473,N_8795,N_8830);
or U13474 (N_13474,N_7735,N_8563);
xor U13475 (N_13475,N_11181,N_6922);
nor U13476 (N_13476,N_9075,N_10943);
nand U13477 (N_13477,N_10205,N_7756);
nand U13478 (N_13478,N_11828,N_10715);
and U13479 (N_13479,N_9306,N_9551);
or U13480 (N_13480,N_7374,N_8959);
nor U13481 (N_13481,N_7941,N_10473);
nand U13482 (N_13482,N_7713,N_6241);
or U13483 (N_13483,N_10187,N_11234);
nand U13484 (N_13484,N_7063,N_9474);
xor U13485 (N_13485,N_8498,N_7936);
nor U13486 (N_13486,N_6352,N_11562);
or U13487 (N_13487,N_7248,N_11693);
or U13488 (N_13488,N_7400,N_10139);
nand U13489 (N_13489,N_9047,N_9440);
xor U13490 (N_13490,N_7147,N_11065);
or U13491 (N_13491,N_11030,N_9465);
or U13492 (N_13492,N_8709,N_8921);
nor U13493 (N_13493,N_11646,N_9591);
nor U13494 (N_13494,N_8010,N_11310);
or U13495 (N_13495,N_6188,N_8486);
xnor U13496 (N_13496,N_8321,N_6155);
nor U13497 (N_13497,N_9272,N_6528);
or U13498 (N_13498,N_9174,N_7318);
or U13499 (N_13499,N_9178,N_11297);
nand U13500 (N_13500,N_11710,N_8060);
xor U13501 (N_13501,N_7605,N_6408);
and U13502 (N_13502,N_8038,N_10107);
nand U13503 (N_13503,N_8443,N_10439);
nor U13504 (N_13504,N_7285,N_6668);
nor U13505 (N_13505,N_7797,N_9723);
and U13506 (N_13506,N_8075,N_9694);
and U13507 (N_13507,N_9951,N_8180);
or U13508 (N_13508,N_6846,N_9548);
and U13509 (N_13509,N_8353,N_6560);
and U13510 (N_13510,N_11044,N_9749);
nor U13511 (N_13511,N_11768,N_10573);
xnor U13512 (N_13512,N_8244,N_6441);
nor U13513 (N_13513,N_9528,N_7952);
or U13514 (N_13514,N_11839,N_9308);
and U13515 (N_13515,N_7317,N_10601);
nand U13516 (N_13516,N_11057,N_8328);
nand U13517 (N_13517,N_10116,N_9842);
and U13518 (N_13518,N_9429,N_10082);
nor U13519 (N_13519,N_6424,N_10890);
nor U13520 (N_13520,N_11000,N_10960);
and U13521 (N_13521,N_7489,N_6262);
nor U13522 (N_13522,N_11031,N_10168);
xor U13523 (N_13523,N_9808,N_7041);
xor U13524 (N_13524,N_9173,N_11708);
xor U13525 (N_13525,N_9266,N_10241);
nor U13526 (N_13526,N_10175,N_6545);
xnor U13527 (N_13527,N_10489,N_10959);
and U13528 (N_13528,N_11943,N_7227);
nor U13529 (N_13529,N_6842,N_6115);
nor U13530 (N_13530,N_6830,N_10239);
xor U13531 (N_13531,N_11568,N_7990);
nor U13532 (N_13532,N_9853,N_9595);
and U13533 (N_13533,N_9459,N_9269);
nor U13534 (N_13534,N_8521,N_10681);
or U13535 (N_13535,N_11422,N_11806);
xnor U13536 (N_13536,N_6877,N_10598);
or U13537 (N_13537,N_11049,N_10431);
and U13538 (N_13538,N_9249,N_9122);
nand U13539 (N_13539,N_6916,N_8793);
nor U13540 (N_13540,N_7454,N_8495);
and U13541 (N_13541,N_10268,N_6646);
xor U13542 (N_13542,N_7978,N_9714);
or U13543 (N_13543,N_10485,N_6145);
nand U13544 (N_13544,N_9665,N_7668);
and U13545 (N_13545,N_8759,N_8566);
nand U13546 (N_13546,N_9100,N_8146);
or U13547 (N_13547,N_8850,N_6977);
and U13548 (N_13548,N_9719,N_10535);
nand U13549 (N_13549,N_9434,N_11489);
nor U13550 (N_13550,N_7078,N_7615);
nand U13551 (N_13551,N_9776,N_6350);
nor U13552 (N_13552,N_11876,N_9182);
and U13553 (N_13553,N_7926,N_11541);
nand U13554 (N_13554,N_9004,N_6231);
nand U13555 (N_13555,N_11384,N_10459);
and U13556 (N_13556,N_6931,N_8137);
nor U13557 (N_13557,N_11376,N_8234);
xnor U13558 (N_13558,N_8184,N_7696);
and U13559 (N_13559,N_6867,N_11813);
and U13560 (N_13560,N_6309,N_8183);
xnor U13561 (N_13561,N_7411,N_10537);
or U13562 (N_13562,N_6316,N_11043);
xor U13563 (N_13563,N_8579,N_6000);
and U13564 (N_13564,N_6573,N_10101);
nand U13565 (N_13565,N_8391,N_9589);
xor U13566 (N_13566,N_10999,N_7504);
and U13567 (N_13567,N_9317,N_8868);
and U13568 (N_13568,N_11117,N_11870);
xnor U13569 (N_13569,N_7100,N_10209);
or U13570 (N_13570,N_7325,N_8930);
and U13571 (N_13571,N_8780,N_11866);
or U13572 (N_13572,N_7750,N_9519);
xnor U13573 (N_13573,N_9598,N_11003);
xor U13574 (N_13574,N_10780,N_9764);
xnor U13575 (N_13575,N_9067,N_8202);
or U13576 (N_13576,N_7912,N_7120);
xor U13577 (N_13577,N_8467,N_10140);
nor U13578 (N_13578,N_10952,N_8189);
xor U13579 (N_13579,N_7637,N_9556);
xor U13580 (N_13580,N_6413,N_7193);
xnor U13581 (N_13581,N_8464,N_8101);
and U13582 (N_13582,N_6385,N_8432);
nor U13583 (N_13583,N_7817,N_6160);
or U13584 (N_13584,N_6809,N_8501);
or U13585 (N_13585,N_8948,N_9962);
xor U13586 (N_13586,N_8869,N_8736);
and U13587 (N_13587,N_6550,N_9625);
and U13588 (N_13588,N_7218,N_6296);
xor U13589 (N_13589,N_9443,N_11929);
and U13590 (N_13590,N_10516,N_6034);
nand U13591 (N_13591,N_7677,N_10383);
nor U13592 (N_13592,N_6467,N_11694);
xnor U13593 (N_13593,N_7023,N_9876);
and U13594 (N_13594,N_10314,N_9227);
nor U13595 (N_13595,N_9926,N_8617);
or U13596 (N_13596,N_11766,N_9330);
nand U13597 (N_13597,N_8854,N_9550);
and U13598 (N_13598,N_8724,N_11727);
and U13599 (N_13599,N_7657,N_9060);
nor U13600 (N_13600,N_7422,N_8120);
xor U13601 (N_13601,N_8754,N_8677);
or U13602 (N_13602,N_11366,N_10803);
nor U13603 (N_13603,N_11113,N_11322);
and U13604 (N_13604,N_7022,N_10309);
or U13605 (N_13605,N_10958,N_9526);
and U13606 (N_13606,N_8938,N_8839);
and U13607 (N_13607,N_8836,N_8096);
or U13608 (N_13608,N_7954,N_11374);
and U13609 (N_13609,N_10292,N_11869);
nand U13610 (N_13610,N_9209,N_8741);
nor U13611 (N_13611,N_7142,N_7527);
nand U13612 (N_13612,N_10995,N_6853);
and U13613 (N_13613,N_11526,N_6276);
and U13614 (N_13614,N_9545,N_7906);
and U13615 (N_13615,N_7336,N_11268);
nor U13616 (N_13616,N_6433,N_6324);
and U13617 (N_13617,N_7429,N_10193);
nor U13618 (N_13618,N_8543,N_7135);
or U13619 (N_13619,N_7148,N_7431);
xnor U13620 (N_13620,N_10273,N_8540);
nor U13621 (N_13621,N_6912,N_10210);
nand U13622 (N_13622,N_11180,N_9505);
nand U13623 (N_13623,N_6987,N_11393);
and U13624 (N_13624,N_11185,N_7617);
nor U13625 (N_13625,N_10329,N_11506);
xnor U13626 (N_13626,N_11862,N_7849);
nand U13627 (N_13627,N_10358,N_8035);
xor U13628 (N_13628,N_10404,N_9013);
nor U13629 (N_13629,N_6832,N_7095);
or U13630 (N_13630,N_7219,N_11266);
nand U13631 (N_13631,N_11835,N_6625);
and U13632 (N_13632,N_11423,N_7267);
and U13633 (N_13633,N_7327,N_6810);
nand U13634 (N_13634,N_8465,N_11789);
and U13635 (N_13635,N_11419,N_7751);
nand U13636 (N_13636,N_10501,N_9523);
or U13637 (N_13637,N_10021,N_8693);
nor U13638 (N_13638,N_10512,N_8360);
xnor U13639 (N_13639,N_10976,N_6908);
and U13640 (N_13640,N_11470,N_8823);
nand U13641 (N_13641,N_6961,N_9477);
nand U13642 (N_13642,N_8827,N_11591);
nand U13643 (N_13643,N_8188,N_11123);
nand U13644 (N_13644,N_6190,N_9845);
xnor U13645 (N_13645,N_7855,N_10897);
nor U13646 (N_13646,N_7143,N_11855);
or U13647 (N_13647,N_9939,N_9036);
or U13648 (N_13648,N_11725,N_6758);
nor U13649 (N_13649,N_10935,N_10250);
and U13650 (N_13650,N_10819,N_9118);
nor U13651 (N_13651,N_10039,N_6464);
nor U13652 (N_13652,N_10282,N_6568);
nand U13653 (N_13653,N_11429,N_8570);
or U13654 (N_13654,N_9142,N_9059);
and U13655 (N_13655,N_9299,N_9649);
nor U13656 (N_13656,N_8707,N_7103);
or U13657 (N_13657,N_8157,N_10150);
or U13658 (N_13658,N_7518,N_11318);
nor U13659 (N_13659,N_7551,N_8476);
xnor U13660 (N_13660,N_10706,N_11998);
nand U13661 (N_13661,N_6542,N_7217);
and U13662 (N_13662,N_9815,N_9924);
nor U13663 (N_13663,N_8103,N_7323);
xnor U13664 (N_13664,N_11114,N_7753);
nand U13665 (N_13665,N_9905,N_6090);
and U13666 (N_13666,N_9996,N_11993);
xnor U13667 (N_13667,N_7471,N_11203);
or U13668 (N_13668,N_8861,N_6938);
nor U13669 (N_13669,N_10829,N_7312);
and U13670 (N_13670,N_10669,N_7381);
nand U13671 (N_13671,N_10065,N_6756);
and U13672 (N_13672,N_6527,N_6246);
xnor U13673 (N_13673,N_7862,N_7238);
nor U13674 (N_13674,N_7321,N_8672);
and U13675 (N_13675,N_6089,N_7074);
and U13676 (N_13676,N_8692,N_8671);
nor U13677 (N_13677,N_10793,N_9652);
nor U13678 (N_13678,N_10128,N_8433);
nor U13679 (N_13679,N_9755,N_11564);
xnor U13680 (N_13680,N_6091,N_9113);
or U13681 (N_13681,N_10252,N_9042);
nor U13682 (N_13682,N_8667,N_6334);
or U13683 (N_13683,N_7865,N_6969);
or U13684 (N_13684,N_6580,N_9507);
or U13685 (N_13685,N_6939,N_10179);
xnor U13686 (N_13686,N_10711,N_8043);
nor U13687 (N_13687,N_10302,N_11454);
or U13688 (N_13688,N_11967,N_7556);
nand U13689 (N_13689,N_6594,N_10428);
xor U13690 (N_13690,N_9810,N_11426);
nand U13691 (N_13691,N_11276,N_8548);
and U13692 (N_13692,N_6232,N_11600);
or U13693 (N_13693,N_6032,N_8986);
nand U13694 (N_13694,N_9160,N_8551);
nand U13695 (N_13695,N_8004,N_8958);
nor U13696 (N_13696,N_11331,N_10938);
or U13697 (N_13697,N_11497,N_9377);
nor U13698 (N_13698,N_11447,N_7579);
and U13699 (N_13699,N_11990,N_11501);
nand U13700 (N_13700,N_9092,N_10278);
nand U13701 (N_13701,N_7505,N_11800);
nor U13702 (N_13702,N_6134,N_8235);
and U13703 (N_13703,N_11219,N_10194);
nor U13704 (N_13704,N_8039,N_6346);
xor U13705 (N_13705,N_6864,N_8597);
nand U13706 (N_13706,N_9563,N_11139);
xnor U13707 (N_13707,N_9464,N_6945);
and U13708 (N_13708,N_9270,N_11054);
and U13709 (N_13709,N_10377,N_11294);
nand U13710 (N_13710,N_9333,N_7907);
nand U13711 (N_13711,N_7086,N_9929);
and U13712 (N_13712,N_7913,N_8299);
nor U13713 (N_13713,N_6282,N_9327);
xnor U13714 (N_13714,N_9789,N_8250);
or U13715 (N_13715,N_7512,N_6777);
nor U13716 (N_13716,N_8322,N_11171);
and U13717 (N_13717,N_6400,N_10849);
nor U13718 (N_13718,N_9236,N_7199);
nor U13719 (N_13719,N_6875,N_8435);
or U13720 (N_13720,N_11131,N_11299);
and U13721 (N_13721,N_9518,N_6785);
and U13722 (N_13722,N_10472,N_10544);
xor U13723 (N_13723,N_8477,N_9848);
xnor U13724 (N_13724,N_7915,N_11684);
nor U13725 (N_13725,N_8696,N_10218);
or U13726 (N_13726,N_9037,N_10721);
nor U13727 (N_13727,N_6157,N_9586);
nor U13728 (N_13728,N_7315,N_9435);
nor U13729 (N_13729,N_11340,N_10154);
nand U13730 (N_13730,N_10425,N_10001);
nor U13731 (N_13731,N_10666,N_10814);
nor U13732 (N_13732,N_8815,N_9671);
xor U13733 (N_13733,N_6819,N_6466);
nand U13734 (N_13734,N_11531,N_10264);
and U13735 (N_13735,N_9822,N_10749);
xnor U13736 (N_13736,N_10353,N_8603);
nand U13737 (N_13737,N_6292,N_8319);
xor U13738 (N_13738,N_9509,N_6782);
and U13739 (N_13739,N_10146,N_8275);
or U13740 (N_13740,N_8430,N_11453);
nand U13741 (N_13741,N_9134,N_6482);
and U13742 (N_13742,N_6984,N_11966);
xor U13743 (N_13743,N_6776,N_6454);
nand U13744 (N_13744,N_10929,N_6240);
or U13745 (N_13745,N_8179,N_10802);
nand U13746 (N_13746,N_8190,N_9797);
nand U13747 (N_13747,N_7624,N_10917);
xnor U13748 (N_13748,N_8143,N_10394);
and U13749 (N_13749,N_7419,N_11809);
and U13750 (N_13750,N_9503,N_6363);
and U13751 (N_13751,N_10254,N_6631);
nor U13752 (N_13752,N_6487,N_10518);
and U13753 (N_13753,N_9818,N_9219);
nand U13754 (N_13754,N_10713,N_7045);
or U13755 (N_13755,N_10612,N_6879);
nand U13756 (N_13756,N_6347,N_6242);
nand U13757 (N_13757,N_8589,N_10906);
nand U13758 (N_13758,N_6733,N_9648);
nand U13759 (N_13759,N_7993,N_8565);
xnor U13760 (N_13760,N_10386,N_6696);
nand U13761 (N_13761,N_11503,N_7687);
or U13762 (N_13762,N_7398,N_8503);
or U13763 (N_13763,N_6893,N_11222);
and U13764 (N_13764,N_10993,N_9906);
xor U13765 (N_13765,N_8263,N_8105);
and U13766 (N_13766,N_10834,N_11236);
or U13767 (N_13767,N_10522,N_7406);
nor U13768 (N_13768,N_7744,N_9050);
nor U13769 (N_13769,N_8156,N_11201);
or U13770 (N_13770,N_6343,N_10112);
or U13771 (N_13771,N_7197,N_7425);
xor U13772 (N_13772,N_8320,N_11660);
nand U13773 (N_13773,N_10397,N_7200);
and U13774 (N_13774,N_11100,N_6172);
and U13775 (N_13775,N_8757,N_8842);
and U13776 (N_13776,N_8470,N_7938);
and U13777 (N_13777,N_11628,N_8135);
xnor U13778 (N_13778,N_11269,N_6814);
xnor U13779 (N_13779,N_8723,N_7524);
or U13780 (N_13780,N_6845,N_7929);
xnor U13781 (N_13781,N_7510,N_10790);
nand U13782 (N_13782,N_7897,N_10110);
nand U13783 (N_13783,N_7528,N_9416);
nor U13784 (N_13784,N_8578,N_8848);
nand U13785 (N_13785,N_9097,N_10724);
and U13786 (N_13786,N_6736,N_10640);
and U13787 (N_13787,N_11761,N_9539);
nand U13788 (N_13788,N_11356,N_11528);
or U13789 (N_13789,N_8887,N_11329);
nand U13790 (N_13790,N_7337,N_11431);
or U13791 (N_13791,N_6499,N_9786);
and U13792 (N_13792,N_8339,N_7225);
nor U13793 (N_13793,N_9226,N_9780);
nand U13794 (N_13794,N_9457,N_10574);
or U13795 (N_13795,N_6820,N_9396);
nand U13796 (N_13796,N_9331,N_11540);
or U13797 (N_13797,N_7553,N_8681);
or U13798 (N_13798,N_11197,N_7430);
nand U13799 (N_13799,N_10953,N_8833);
nor U13800 (N_13800,N_9030,N_11637);
and U13801 (N_13801,N_6182,N_6531);
xnor U13802 (N_13802,N_6384,N_6058);
nor U13803 (N_13803,N_6044,N_9512);
and U13804 (N_13804,N_10326,N_11942);
xor U13805 (N_13805,N_6718,N_10754);
and U13806 (N_13806,N_6040,N_6818);
nand U13807 (N_13807,N_7102,N_8066);
nand U13808 (N_13808,N_7638,N_10177);
nand U13809 (N_13809,N_11242,N_11073);
or U13810 (N_13810,N_7237,N_7933);
and U13811 (N_13811,N_10415,N_8163);
nand U13812 (N_13812,N_8040,N_7725);
nor U13813 (N_13813,N_11796,N_11021);
xor U13814 (N_13814,N_10776,N_9153);
nor U13815 (N_13815,N_11491,N_6584);
nand U13816 (N_13816,N_7882,N_6964);
xor U13817 (N_13817,N_9919,N_8628);
and U13818 (N_13818,N_6288,N_8658);
xor U13819 (N_13819,N_10821,N_8625);
xor U13820 (N_13820,N_8515,N_6838);
xnor U13821 (N_13821,N_9374,N_9329);
xnor U13822 (N_13822,N_10765,N_8904);
xnor U13823 (N_13823,N_10594,N_9956);
nand U13824 (N_13824,N_9787,N_11370);
xor U13825 (N_13825,N_7785,N_7215);
xnor U13826 (N_13826,N_7847,N_8762);
and U13827 (N_13827,N_9891,N_8879);
nor U13828 (N_13828,N_10156,N_11377);
and U13829 (N_13829,N_6335,N_11847);
nand U13830 (N_13830,N_9351,N_8118);
and U13831 (N_13831,N_8151,N_7299);
xnor U13832 (N_13832,N_6206,N_8892);
nor U13833 (N_13833,N_11661,N_8572);
nand U13834 (N_13834,N_7770,N_6635);
nor U13835 (N_13835,N_6645,N_7728);
xor U13836 (N_13836,N_6179,N_10099);
nand U13837 (N_13837,N_8632,N_8399);
xor U13838 (N_13838,N_10013,N_9197);
and U13839 (N_13839,N_6015,N_7813);
and U13840 (N_13840,N_7348,N_8726);
xnor U13841 (N_13841,N_8655,N_10098);
or U13842 (N_13842,N_8412,N_6590);
or U13843 (N_13843,N_9772,N_6603);
xor U13844 (N_13844,N_8286,N_11433);
or U13845 (N_13845,N_8995,N_7732);
or U13846 (N_13846,N_10438,N_9271);
xnor U13847 (N_13847,N_7716,N_6409);
xnor U13848 (N_13848,N_9216,N_11516);
xor U13849 (N_13849,N_8710,N_8911);
and U13850 (N_13850,N_9976,N_9584);
xor U13851 (N_13851,N_7916,N_6839);
or U13852 (N_13852,N_6693,N_7343);
and U13853 (N_13853,N_11816,N_10581);
xnor U13854 (N_13854,N_10391,N_6740);
or U13855 (N_13855,N_7625,N_7076);
nor U13856 (N_13856,N_11666,N_6886);
and U13857 (N_13857,N_9978,N_8484);
or U13858 (N_13858,N_6683,N_11818);
and U13859 (N_13859,N_10085,N_9928);
or U13860 (N_13860,N_6924,N_10846);
or U13861 (N_13861,N_7548,N_9838);
nor U13862 (N_13862,N_7442,N_10553);
nand U13863 (N_13863,N_10080,N_8997);
nand U13864 (N_13864,N_6171,N_9358);
nor U13865 (N_13865,N_9704,N_8385);
nor U13866 (N_13866,N_11306,N_11239);
or U13867 (N_13867,N_8511,N_8514);
and U13868 (N_13868,N_7117,N_7417);
or U13869 (N_13869,N_11026,N_7477);
and U13870 (N_13870,N_8227,N_8518);
or U13871 (N_13871,N_8123,N_10064);
xor U13872 (N_13872,N_8046,N_11571);
and U13873 (N_13873,N_7698,N_8393);
xnor U13874 (N_13874,N_11338,N_6888);
and U13875 (N_13875,N_6956,N_7969);
and U13876 (N_13876,N_7833,N_7892);
nand U13877 (N_13877,N_10152,N_6449);
nor U13878 (N_13878,N_7069,N_7249);
or U13879 (N_13879,N_7977,N_11514);
or U13880 (N_13880,N_6548,N_8968);
xor U13881 (N_13881,N_11857,N_11496);
or U13882 (N_13882,N_8747,N_8573);
xor U13883 (N_13883,N_11205,N_11451);
nand U13884 (N_13884,N_9338,N_6593);
nor U13885 (N_13885,N_10018,N_9958);
nor U13886 (N_13886,N_11142,N_9709);
or U13887 (N_13887,N_8115,N_9328);
nor U13888 (N_13888,N_7079,N_11593);
nand U13889 (N_13889,N_8154,N_10474);
xor U13890 (N_13890,N_6131,N_8340);
xor U13891 (N_13891,N_8539,N_8387);
xnor U13892 (N_13892,N_6717,N_7520);
nor U13893 (N_13893,N_6420,N_7870);
nand U13894 (N_13894,N_9940,N_9942);
and U13895 (N_13895,N_7558,N_7367);
nor U13896 (N_13896,N_10300,N_7136);
nand U13897 (N_13897,N_6353,N_11732);
nor U13898 (N_13898,N_11790,N_8298);
xor U13899 (N_13899,N_10032,N_7105);
xor U13900 (N_13900,N_6003,N_10163);
and U13901 (N_13901,N_10674,N_7201);
or U13902 (N_13902,N_11890,N_10629);
or U13903 (N_13903,N_8656,N_7077);
and U13904 (N_13904,N_10728,N_9613);
or U13905 (N_13905,N_11012,N_11705);
and U13906 (N_13906,N_9441,N_11960);
nor U13907 (N_13907,N_9368,N_9529);
or U13908 (N_13908,N_11138,N_7825);
nor U13909 (N_13909,N_6544,N_8688);
nor U13910 (N_13910,N_6502,N_6079);
xor U13911 (N_13911,N_9195,N_11042);
nand U13912 (N_13912,N_6659,N_8701);
xnor U13913 (N_13913,N_9971,N_9535);
nand U13914 (N_13914,N_11702,N_8478);
or U13915 (N_13915,N_8204,N_10324);
and U13916 (N_13916,N_7202,N_8641);
and U13917 (N_13917,N_10513,N_9576);
nor U13918 (N_13918,N_7800,N_7428);
or U13919 (N_13919,N_6494,N_10963);
or U13920 (N_13920,N_11629,N_7084);
and U13921 (N_13921,N_8881,N_11082);
nor U13922 (N_13922,N_6697,N_10467);
nor U13923 (N_13923,N_8052,N_10475);
xnor U13924 (N_13924,N_7094,N_11010);
nor U13925 (N_13925,N_8988,N_7481);
or U13926 (N_13926,N_11559,N_10490);
or U13927 (N_13927,N_10911,N_6512);
nand U13928 (N_13928,N_9722,N_10799);
nor U13929 (N_13929,N_6066,N_10015);
nand U13930 (N_13930,N_9438,N_10591);
xnor U13931 (N_13931,N_6611,N_9781);
nor U13932 (N_13932,N_7536,N_6967);
nor U13933 (N_13933,N_9538,N_9499);
nand U13934 (N_13934,N_6674,N_9706);
nor U13935 (N_13935,N_9458,N_10560);
nand U13936 (N_13936,N_8771,N_8288);
and U13937 (N_13937,N_8468,N_10812);
xor U13938 (N_13938,N_7175,N_6627);
and U13939 (N_13939,N_10977,N_9896);
nand U13940 (N_13940,N_11678,N_6273);
nand U13941 (N_13941,N_10684,N_11032);
or U13942 (N_13942,N_6648,N_9102);
or U13943 (N_13943,N_9580,N_9123);
or U13944 (N_13944,N_6743,N_6402);
or U13945 (N_13945,N_11756,N_7683);
xor U13946 (N_13946,N_7322,N_11602);
nor U13947 (N_13947,N_6963,N_6805);
xor U13948 (N_13948,N_11721,N_6617);
or U13949 (N_13949,N_9093,N_11812);
and U13950 (N_13950,N_6536,N_9300);
nor U13951 (N_13951,N_6951,N_8076);
nand U13952 (N_13952,N_6116,N_10259);
and U13953 (N_13953,N_8425,N_8927);
and U13954 (N_13954,N_10782,N_10996);
and U13955 (N_13955,N_9984,N_11861);
nand U13956 (N_13956,N_11212,N_8074);
nor U13957 (N_13957,N_7636,N_11344);
nand U13958 (N_13958,N_9068,N_8191);
or U13959 (N_13959,N_9277,N_8338);
nor U13960 (N_13960,N_7786,N_6894);
nand U13961 (N_13961,N_10090,N_8213);
nor U13962 (N_13962,N_8277,N_6459);
nand U13963 (N_13963,N_9901,N_10280);
nor U13964 (N_13964,N_9357,N_7988);
xnor U13965 (N_13965,N_11972,N_9899);
nor U13966 (N_13966,N_6446,N_11549);
xor U13967 (N_13967,N_9072,N_11008);
nand U13968 (N_13968,N_10729,N_11547);
nand U13969 (N_13969,N_8489,N_10174);
and U13970 (N_13970,N_6002,N_7433);
and U13971 (N_13971,N_9054,N_7662);
nor U13972 (N_13972,N_6348,N_7985);
nand U13973 (N_13973,N_6761,N_10453);
and U13974 (N_13974,N_10984,N_11798);
nor U13975 (N_13975,N_10604,N_7072);
nor U13976 (N_13976,N_6109,N_11211);
xnor U13977 (N_13977,N_6461,N_7981);
or U13978 (N_13978,N_6020,N_9514);
nand U13979 (N_13979,N_10424,N_8216);
and U13980 (N_13980,N_9340,N_8411);
xnor U13981 (N_13981,N_8417,N_10222);
nand U13982 (N_13982,N_10265,N_8871);
and U13983 (N_13983,N_10458,N_9469);
and U13984 (N_13984,N_8636,N_6326);
nand U13985 (N_13985,N_10843,N_11669);
and U13986 (N_13986,N_10037,N_10863);
nand U13987 (N_13987,N_11218,N_6679);
and U13988 (N_13988,N_11897,N_11555);
xor U13989 (N_13989,N_11319,N_9768);
or U13990 (N_13990,N_7845,N_10009);
xor U13991 (N_13991,N_6189,N_9628);
nand U13992 (N_13992,N_7998,N_10761);
and U13993 (N_13993,N_9938,N_7377);
xor U13994 (N_13994,N_7816,N_9770);
nand U13995 (N_13995,N_11441,N_9332);
or U13996 (N_13996,N_11303,N_7277);
nor U13997 (N_13997,N_9342,N_10072);
nor U13998 (N_13998,N_10971,N_9634);
and U13999 (N_13999,N_6177,N_10811);
and U14000 (N_14000,N_7062,N_8113);
and U14001 (N_14001,N_7866,N_7663);
nand U14002 (N_14002,N_11533,N_11163);
nor U14003 (N_14003,N_6841,N_11713);
nor U14004 (N_14004,N_7211,N_10323);
nand U14005 (N_14005,N_11238,N_10741);
and U14006 (N_14006,N_8735,N_6368);
nand U14007 (N_14007,N_11466,N_8686);
nand U14008 (N_14008,N_7798,N_10296);
nand U14009 (N_14009,N_9702,N_6194);
nor U14010 (N_14010,N_11414,N_11579);
xnor U14011 (N_14011,N_9868,N_7313);
nor U14012 (N_14012,N_7622,N_11208);
nor U14013 (N_14013,N_7262,N_6341);
nor U14014 (N_14014,N_10691,N_10190);
and U14015 (N_14015,N_10076,N_6654);
or U14016 (N_14016,N_8633,N_10319);
nand U14017 (N_14017,N_8608,N_7726);
nand U14018 (N_14018,N_11118,N_6844);
and U14019 (N_14019,N_11772,N_10636);
nand U14020 (N_14020,N_6698,N_8236);
nand U14021 (N_14021,N_6771,N_8001);
and U14022 (N_14022,N_8502,N_7483);
and U14023 (N_14023,N_9700,N_9961);
nor U14024 (N_14024,N_11398,N_7210);
nor U14025 (N_14025,N_9341,N_8055);
and U14026 (N_14026,N_10925,N_6321);
nor U14027 (N_14027,N_6065,N_9324);
and U14028 (N_14028,N_11315,N_6269);
nor U14029 (N_14029,N_9565,N_11474);
nand U14030 (N_14030,N_9378,N_6663);
nand U14031 (N_14031,N_11116,N_10171);
nand U14032 (N_14032,N_10675,N_9741);
nand U14033 (N_14033,N_6159,N_6518);
nand U14034 (N_14034,N_7375,N_6535);
nand U14035 (N_14035,N_8205,N_9146);
and U14036 (N_14036,N_9253,N_9660);
nor U14037 (N_14037,N_6135,N_8493);
and U14038 (N_14038,N_10509,N_6062);
and U14039 (N_14039,N_7360,N_6991);
nor U14040 (N_14040,N_6114,N_7884);
xnor U14041 (N_14041,N_10902,N_8645);
or U14042 (N_14042,N_8437,N_9751);
and U14043 (N_14043,N_9733,N_9255);
nand U14044 (N_14044,N_10276,N_10600);
and U14045 (N_14045,N_6976,N_11490);
and U14046 (N_14046,N_11009,N_9437);
nand U14047 (N_14047,N_11101,N_10151);
nor U14048 (N_14048,N_6033,N_6936);
and U14049 (N_14049,N_6323,N_10844);
xnor U14050 (N_14050,N_6585,N_9020);
and U14051 (N_14051,N_11327,N_8017);
nand U14052 (N_14052,N_11064,N_10038);
or U14053 (N_14053,N_11335,N_11401);
xor U14054 (N_14054,N_11079,N_10733);
and U14055 (N_14055,N_7767,N_8370);
nand U14056 (N_14056,N_9307,N_9656);
and U14057 (N_14057,N_6902,N_8713);
nor U14058 (N_14058,N_8022,N_9430);
xor U14059 (N_14059,N_8285,N_11609);
nor U14060 (N_14060,N_6121,N_9144);
nand U14061 (N_14061,N_10339,N_8586);
or U14062 (N_14062,N_7900,N_6850);
nand U14063 (N_14063,N_7639,N_8770);
nand U14064 (N_14064,N_7346,N_10331);
nor U14065 (N_14065,N_7935,N_8171);
nor U14066 (N_14066,N_11192,N_9765);
xor U14067 (N_14067,N_7563,N_6120);
nand U14068 (N_14068,N_7588,N_7366);
xnor U14069 (N_14069,N_8546,N_9515);
and U14070 (N_14070,N_9094,N_11610);
and U14071 (N_14071,N_7379,N_8317);
xnor U14072 (N_14072,N_7706,N_8119);
xor U14073 (N_14073,N_11262,N_6455);
and U14074 (N_14074,N_10246,N_9946);
nor U14075 (N_14075,N_9870,N_8935);
xor U14076 (N_14076,N_7376,N_7562);
xnor U14077 (N_14077,N_10114,N_11270);
or U14078 (N_14078,N_7473,N_10310);
or U14079 (N_14079,N_6884,N_6615);
nand U14080 (N_14080,N_11016,N_11937);
nand U14081 (N_14081,N_6126,N_7043);
xnor U14082 (N_14082,N_11940,N_9313);
xnor U14083 (N_14083,N_8242,N_8629);
or U14084 (N_14084,N_11911,N_11845);
nand U14085 (N_14085,N_11675,N_10732);
nand U14086 (N_14086,N_7180,N_6904);
xnor U14087 (N_14087,N_11442,N_8962);
xnor U14088 (N_14088,N_7730,N_9222);
and U14089 (N_14089,N_9350,N_7807);
nor U14090 (N_14090,N_7416,N_9062);
or U14091 (N_14091,N_10527,N_8228);
nor U14092 (N_14092,N_7514,N_8851);
or U14093 (N_14093,N_9497,N_8810);
nor U14094 (N_14094,N_10572,N_6037);
nand U14095 (N_14095,N_9099,N_11435);
xor U14096 (N_14096,N_9999,N_8033);
and U14097 (N_14097,N_9909,N_8097);
xnor U14098 (N_14098,N_6714,N_8136);
and U14099 (N_14099,N_9543,N_9631);
and U14100 (N_14100,N_6960,N_8784);
and U14101 (N_14101,N_7259,N_9085);
or U14102 (N_14102,N_7791,N_7247);
or U14103 (N_14103,N_10702,N_7470);
xnor U14104 (N_14104,N_8731,N_10161);
or U14105 (N_14105,N_10528,N_11574);
nand U14106 (N_14106,N_10192,N_11595);
or U14107 (N_14107,N_6983,N_10409);
nand U14108 (N_14108,N_11359,N_11573);
xor U14109 (N_14109,N_8446,N_8287);
nor U14110 (N_14110,N_9541,N_6283);
nand U14111 (N_14111,N_9511,N_11364);
or U14112 (N_14112,N_7839,N_9349);
nand U14113 (N_14113,N_11905,N_9133);
or U14114 (N_14114,N_11158,N_11260);
nand U14115 (N_14115,N_7183,N_6790);
nand U14116 (N_14116,N_8058,N_6170);
and U14117 (N_14117,N_8447,N_6699);
and U14118 (N_14118,N_6803,N_9325);
nor U14119 (N_14119,N_9106,N_6204);
nand U14120 (N_14120,N_11644,N_6229);
and U14121 (N_14121,N_8612,N_8166);
and U14122 (N_14122,N_7616,N_10203);
and U14123 (N_14123,N_8870,N_9980);
or U14124 (N_14124,N_9736,N_8838);
nor U14125 (N_14125,N_6094,N_11596);
nand U14126 (N_14126,N_10933,N_11924);
xor U14127 (N_14127,N_10854,N_6666);
nand U14128 (N_14128,N_6546,N_6356);
and U14129 (N_14129,N_9336,N_7719);
and U14130 (N_14130,N_6883,N_9074);
nor U14131 (N_14131,N_10486,N_11507);
and U14132 (N_14132,N_11653,N_8414);
xor U14133 (N_14133,N_9922,N_11288);
nand U14134 (N_14134,N_8727,N_6694);
or U14135 (N_14135,N_9305,N_11285);
nand U14136 (N_14136,N_9467,N_9729);
nand U14137 (N_14137,N_11343,N_9731);
nand U14138 (N_14138,N_7310,N_9242);
or U14139 (N_14139,N_7925,N_10044);
nor U14140 (N_14140,N_7578,N_9088);
xor U14141 (N_14141,N_9053,N_6333);
or U14142 (N_14142,N_7368,N_8649);
or U14143 (N_14143,N_6799,N_6944);
or U14144 (N_14144,N_6493,N_7141);
nor U14145 (N_14145,N_11612,N_10213);
nor U14146 (N_14146,N_7284,N_7205);
and U14147 (N_14147,N_11807,N_7918);
and U14148 (N_14148,N_6496,N_8497);
and U14149 (N_14149,N_9697,N_7060);
xor U14150 (N_14150,N_10517,N_9268);
nand U14151 (N_14151,N_6263,N_10220);
nand U14152 (N_14152,N_6523,N_9221);
and U14153 (N_14153,N_9812,N_8781);
nor U14154 (N_14154,N_11826,N_6307);
nor U14155 (N_14155,N_7359,N_9419);
or U14156 (N_14156,N_11293,N_9907);
nor U14157 (N_14157,N_11641,N_7097);
nor U14158 (N_14158,N_10022,N_11927);
or U14159 (N_14159,N_9141,N_7589);
and U14160 (N_14160,N_11284,N_7495);
xnor U14161 (N_14161,N_11166,N_9716);
and U14162 (N_14162,N_9554,N_8365);
xor U14163 (N_14163,N_9553,N_10617);
nor U14164 (N_14164,N_11900,N_6881);
nand U14165 (N_14165,N_6427,N_9596);
nand U14166 (N_14166,N_7989,N_6437);
and U14167 (N_14167,N_10306,N_9953);
xnor U14168 (N_14168,N_10387,N_6706);
and U14169 (N_14169,N_6373,N_9914);
nand U14170 (N_14170,N_8782,N_10274);
or U14171 (N_14171,N_8092,N_6954);
xnor U14172 (N_14172,N_8251,N_9616);
and U14173 (N_14173,N_11383,N_9568);
xor U14174 (N_14174,N_7734,N_7843);
nand U14175 (N_14175,N_9018,N_6757);
and U14176 (N_14176,N_8078,N_8452);
nand U14177 (N_14177,N_11730,N_7232);
nor U14178 (N_14178,N_10548,N_11068);
nand U14179 (N_14179,N_10816,N_11745);
xnor U14180 (N_14180,N_6988,N_11059);
and U14181 (N_14181,N_9869,N_11925);
nor U14182 (N_14182,N_11723,N_6205);
and U14183 (N_14183,N_8445,N_10004);
nor U14184 (N_14184,N_10921,N_11952);
or U14185 (N_14185,N_9858,N_6848);
or U14186 (N_14186,N_8159,N_6048);
and U14187 (N_14187,N_9921,N_6360);
xor U14188 (N_14188,N_10725,N_8217);
and U14189 (N_14189,N_6093,N_11715);
nand U14190 (N_14190,N_6682,N_11194);
and U14191 (N_14191,N_11560,N_8260);
or U14192 (N_14192,N_11040,N_10199);
nor U14193 (N_14193,N_11006,N_8207);
nor U14194 (N_14194,N_6458,N_9481);
xor U14195 (N_14195,N_7838,N_8885);
nand U14196 (N_14196,N_11351,N_7233);
or U14197 (N_14197,N_9627,N_10342);
or U14198 (N_14198,N_7501,N_7240);
nor U14199 (N_14199,N_7373,N_7942);
nor U14200 (N_14200,N_8937,N_7863);
nor U14201 (N_14201,N_7264,N_9425);
or U14202 (N_14202,N_9874,N_6569);
or U14203 (N_14203,N_6896,N_10994);
xnor U14204 (N_14204,N_8826,N_6175);
nor U14205 (N_14205,N_7042,N_6151);
and U14206 (N_14206,N_6381,N_7759);
or U14207 (N_14207,N_8448,N_7383);
nand U14208 (N_14208,N_10436,N_11844);
nor U14209 (N_14209,N_8253,N_6748);
xor U14210 (N_14210,N_7465,N_10215);
or U14211 (N_14211,N_6940,N_7171);
nor U14212 (N_14212,N_10532,N_6310);
nor U14213 (N_14213,N_7188,N_8517);
or U14214 (N_14214,N_11308,N_10000);
nor U14215 (N_14215,N_9527,N_9737);
and U14216 (N_14216,N_8627,N_7482);
or U14217 (N_14217,N_10571,N_9995);
nand U14218 (N_14218,N_8558,N_8169);
xnor U14219 (N_14219,N_6510,N_8193);
nand U14220 (N_14220,N_6887,N_6088);
nor U14221 (N_14221,N_6260,N_8132);
xnor U14222 (N_14222,N_11107,N_11815);
nand U14223 (N_14223,N_6255,N_11210);
xnor U14224 (N_14224,N_9376,N_8081);
xnor U14225 (N_14225,N_9354,N_8371);
or U14226 (N_14226,N_6823,N_6606);
xnor U14227 (N_14227,N_7649,N_7410);
and U14228 (N_14228,N_6557,N_6481);
and U14229 (N_14229,N_9790,N_8273);
nor U14230 (N_14230,N_8624,N_8766);
xor U14231 (N_14231,N_6383,N_7402);
or U14232 (N_14232,N_11105,N_8406);
nand U14233 (N_14233,N_7545,N_8695);
and U14234 (N_14234,N_8282,N_8571);
nand U14235 (N_14235,N_7464,N_7727);
xor U14236 (N_14236,N_8107,N_9185);
or U14237 (N_14237,N_8381,N_6183);
nor U14238 (N_14238,N_10028,N_9931);
and U14239 (N_14239,N_7629,N_8354);
and U14240 (N_14240,N_11802,N_11974);
nand U14241 (N_14241,N_6520,N_8609);
nor U14242 (N_14242,N_9829,N_6779);
nor U14243 (N_14243,N_11109,N_6319);
nand U14244 (N_14244,N_7623,N_10418);
and U14245 (N_14245,N_7905,N_7057);
nand U14246 (N_14246,N_8858,N_10435);
nor U14247 (N_14247,N_8142,N_6369);
xor U14248 (N_14248,N_8789,N_9624);
nand U14249 (N_14249,N_11879,N_9212);
nand U14250 (N_14250,N_9023,N_9862);
or U14251 (N_14251,N_6634,N_11585);
or U14252 (N_14252,N_9601,N_10207);
xnor U14253 (N_14253,N_8794,N_10271);
nand U14254 (N_14254,N_8200,N_11439);
nor U14255 (N_14255,N_8585,N_11251);
or U14256 (N_14256,N_10895,N_6035);
and U14257 (N_14257,N_9445,N_10827);
nor U14258 (N_14258,N_6287,N_9114);
nor U14259 (N_14259,N_7235,N_7498);
and U14260 (N_14260,N_9131,N_7758);
and U14261 (N_14261,N_11233,N_6332);
nor U14262 (N_14262,N_9530,N_10904);
nand U14263 (N_14263,N_11823,N_8874);
nor U14264 (N_14264,N_8524,N_7405);
xor U14265 (N_14265,N_8691,N_9813);
nand U14266 (N_14266,N_11984,N_7792);
nor U14267 (N_14267,N_11350,N_8812);
xnor U14268 (N_14268,N_10647,N_11394);
or U14269 (N_14269,N_9489,N_10120);
nand U14270 (N_14270,N_9205,N_6952);
or U14271 (N_14271,N_11096,N_11936);
nand U14272 (N_14272,N_8389,N_8813);
nor U14273 (N_14273,N_8534,N_9607);
and U14274 (N_14274,N_6284,N_6214);
nand U14275 (N_14275,N_10750,N_11458);
nor U14276 (N_14276,N_6766,N_11592);
and U14277 (N_14277,N_11642,N_10398);
nand U14278 (N_14278,N_10316,N_11850);
nor U14279 (N_14279,N_7349,N_11450);
nand U14280 (N_14280,N_7924,N_8821);
or U14281 (N_14281,N_8357,N_7351);
nor U14282 (N_14282,N_10330,N_10529);
xnor U14283 (N_14283,N_8530,N_8900);
or U14284 (N_14284,N_7266,N_7091);
and U14285 (N_14285,N_8772,N_11821);
xor U14286 (N_14286,N_10159,N_9897);
nor U14287 (N_14287,N_6438,N_7329);
nand U14288 (N_14288,N_10877,N_10784);
xor U14289 (N_14289,N_9536,N_7660);
and U14290 (N_14290,N_10981,N_9246);
nor U14291 (N_14291,N_9600,N_8952);
and U14292 (N_14292,N_7354,N_9056);
and U14293 (N_14293,N_8914,N_10605);
or U14294 (N_14294,N_7056,N_11440);
xor U14295 (N_14295,N_10665,N_11018);
nand U14296 (N_14296,N_6490,N_11020);
or U14297 (N_14297,N_8761,N_7438);
nor U14298 (N_14298,N_7016,N_11052);
and U14299 (N_14299,N_9986,N_6767);
xnor U14300 (N_14300,N_6671,N_7881);
and U14301 (N_14301,N_8516,N_6130);
and U14302 (N_14302,N_6561,N_10455);
or U14303 (N_14303,N_11852,N_8942);
or U14304 (N_14304,N_10941,N_11695);
and U14305 (N_14305,N_9705,N_9913);
xnor U14306 (N_14306,N_7515,N_10533);
and U14307 (N_14307,N_6149,N_10756);
and U14308 (N_14308,N_9303,N_9692);
nor U14309 (N_14309,N_11471,N_8229);
or U14310 (N_14310,N_6577,N_8401);
xnor U14311 (N_14311,N_9413,N_11598);
nor U14312 (N_14312,N_10419,N_6658);
xor U14313 (N_14313,N_7503,N_7250);
or U14314 (N_14314,N_8428,N_6966);
nor U14315 (N_14315,N_7644,N_7632);
nand U14316 (N_14316,N_9943,N_7829);
xnor U14317 (N_14317,N_7162,N_10646);
nor U14318 (N_14318,N_6129,N_11056);
and U14319 (N_14319,N_9164,N_9487);
and U14320 (N_14320,N_6300,N_7601);
xnor U14321 (N_14321,N_9809,N_10841);
and U14322 (N_14322,N_10566,N_7159);
nand U14323 (N_14323,N_7363,N_7292);
xor U14324 (N_14324,N_8243,N_11773);
and U14325 (N_14325,N_8702,N_11765);
or U14326 (N_14326,N_11603,N_10887);
and U14327 (N_14327,N_10677,N_6992);
nor U14328 (N_14328,N_7361,N_6450);
nor U14329 (N_14329,N_7810,N_9510);
xnor U14330 (N_14330,N_10987,N_10857);
nor U14331 (N_14331,N_6315,N_10401);
or U14332 (N_14332,N_8662,N_10626);
or U14333 (N_14333,N_6695,N_6858);
xor U14334 (N_14334,N_10882,N_8292);
nand U14335 (N_14335,N_7053,N_10649);
xor U14336 (N_14336,N_7671,N_11582);
xnor U14337 (N_14337,N_6647,N_10223);
nand U14338 (N_14338,N_9493,N_11257);
xnor U14339 (N_14339,N_11387,N_8063);
or U14340 (N_14340,N_10492,N_11753);
nor U14341 (N_14341,N_9230,N_7478);
or U14342 (N_14342,N_7540,N_10433);
or U14343 (N_14343,N_10695,N_9651);
or U14344 (N_14344,N_8849,N_10272);
nor U14345 (N_14345,N_6412,N_6375);
and U14346 (N_14346,N_10980,N_8755);
xnor U14347 (N_14347,N_11066,N_11188);
and U14348 (N_14348,N_8272,N_9557);
xnor U14349 (N_14349,N_8377,N_9424);
xnor U14350 (N_14350,N_7138,N_8831);
nand U14351 (N_14351,N_11108,N_8550);
nor U14352 (N_14352,N_6440,N_8024);
xnor U14353 (N_14353,N_11840,N_11085);
nand U14354 (N_14354,N_7653,N_8109);
nand U14355 (N_14355,N_11149,N_10427);
nand U14356 (N_14356,N_8882,N_7122);
or U14357 (N_14357,N_6042,N_11317);
or U14358 (N_14358,N_8561,N_7618);
and U14359 (N_14359,N_7500,N_11445);
nand U14360 (N_14360,N_11780,N_7423);
nor U14361 (N_14361,N_7573,N_11948);
and U14362 (N_14362,N_10157,N_7182);
nor U14363 (N_14363,N_8808,N_8335);
or U14364 (N_14364,N_7682,N_8822);
nand U14365 (N_14365,N_8920,N_9090);
nor U14366 (N_14366,N_7793,N_9871);
xnor U14367 (N_14367,N_11868,N_11159);
nor U14368 (N_14368,N_6783,N_6687);
nand U14369 (N_14369,N_7083,N_7170);
nor U14370 (N_14370,N_7606,N_10315);
nand U14371 (N_14371,N_6689,N_10856);
nand U14372 (N_14372,N_8527,N_8811);
or U14373 (N_14373,N_10287,N_10495);
nor U14374 (N_14374,N_10408,N_8315);
or U14375 (N_14375,N_6726,N_9606);
and U14376 (N_14376,N_9191,N_8728);
xnor U14377 (N_14377,N_6890,N_7963);
nor U14378 (N_14378,N_8576,N_8362);
nor U14379 (N_14379,N_10311,N_8165);
or U14380 (N_14380,N_11744,N_6038);
or U14381 (N_14381,N_10998,N_6609);
xnor U14382 (N_14382,N_10005,N_11409);
xor U14383 (N_14383,N_11078,N_10002);
or U14384 (N_14384,N_9148,N_9923);
xnor U14385 (N_14385,N_10463,N_8030);
and U14386 (N_14386,N_6007,N_11578);
xor U14387 (N_14387,N_10974,N_7494);
xor U14388 (N_14388,N_8700,N_10889);
nand U14389 (N_14389,N_8130,N_8799);
and U14390 (N_14390,N_8471,N_11968);
or U14391 (N_14391,N_7044,N_9558);
or U14392 (N_14392,N_6786,N_10332);
and U14393 (N_14393,N_10026,N_8346);
nand U14394 (N_14394,N_9643,N_11060);
xnor U14395 (N_14395,N_11228,N_8410);
xnor U14396 (N_14396,N_6885,N_8840);
and U14397 (N_14397,N_6358,N_7370);
nor U14398 (N_14398,N_10508,N_9767);
xor U14399 (N_14399,N_9725,N_7289);
and U14400 (N_14400,N_6652,N_10243);
nand U14401 (N_14401,N_10671,N_9811);
xor U14402 (N_14402,N_10123,N_6503);
nand U14403 (N_14403,N_8505,N_9391);
nor U14404 (N_14404,N_8186,N_11430);
nand U14405 (N_14405,N_8158,N_6125);
xnor U14406 (N_14406,N_10771,N_11838);
nor U14407 (N_14407,N_8601,N_9784);
xnor U14408 (N_14408,N_9495,N_8434);
or U14409 (N_14409,N_9759,N_9475);
xor U14410 (N_14410,N_9415,N_6185);
nor U14411 (N_14411,N_8405,N_6835);
xnor U14412 (N_14412,N_10564,N_9900);
nand U14413 (N_14413,N_8025,N_9234);
or U14414 (N_14414,N_7891,N_8596);
or U14415 (N_14415,N_9473,N_10129);
nor U14416 (N_14416,N_11050,N_7047);
nand U14417 (N_14417,N_11532,N_8767);
nor U14418 (N_14418,N_6202,N_8374);
and U14419 (N_14419,N_10530,N_6891);
and U14420 (N_14420,N_9730,N_8420);
xor U14421 (N_14421,N_11473,N_8164);
xnor U14422 (N_14422,N_9678,N_11954);
nor U14423 (N_14423,N_10008,N_6404);
and U14424 (N_14424,N_6622,N_10322);
or U14425 (N_14425,N_7048,N_10452);
or U14426 (N_14426,N_10003,N_9442);
and U14427 (N_14427,N_11273,N_9948);
or U14428 (N_14428,N_8192,N_10577);
and U14429 (N_14429,N_9082,N_11743);
nand U14430 (N_14430,N_10660,N_8508);
and U14431 (N_14431,N_7764,N_8523);
or U14432 (N_14432,N_9992,N_6448);
nand U14433 (N_14433,N_8290,N_10446);
nand U14434 (N_14434,N_9462,N_11235);
nand U14435 (N_14435,N_6589,N_10333);
or U14436 (N_14436,N_10499,N_6469);
nand U14437 (N_14437,N_8014,N_9935);
xnor U14438 (N_14438,N_9239,N_8966);
and U14439 (N_14439,N_10914,N_9742);
and U14440 (N_14440,N_10985,N_11004);
nor U14441 (N_14441,N_9010,N_8294);
xor U14442 (N_14442,N_11183,N_10074);
and U14443 (N_14443,N_6025,N_10979);
or U14444 (N_14444,N_10447,N_8898);
xor U14445 (N_14445,N_11207,N_9646);
or U14446 (N_14446,N_10957,N_8535);
xnor U14447 (N_14447,N_10818,N_6142);
xnor U14448 (N_14448,N_8323,N_7914);
xnor U14449 (N_14449,N_11956,N_9083);
or U14450 (N_14450,N_7574,N_11074);
and U14451 (N_14451,N_10609,N_7177);
nand U14452 (N_14452,N_8940,N_6703);
and U14453 (N_14453,N_6787,N_7975);
nor U14454 (N_14454,N_7787,N_11851);
or U14455 (N_14455,N_6608,N_7106);
or U14456 (N_14456,N_9632,N_11373);
or U14457 (N_14457,N_10551,N_8631);
nor U14458 (N_14458,N_6012,N_6162);
xor U14459 (N_14459,N_7733,N_9746);
nand U14460 (N_14460,N_8704,N_6213);
or U14461 (N_14461,N_9061,N_8274);
nor U14462 (N_14462,N_11216,N_9041);
nor U14463 (N_14463,N_10764,N_6981);
nor U14464 (N_14464,N_7020,N_7722);
nor U14465 (N_14465,N_7018,N_6127);
and U14466 (N_14466,N_11545,N_8547);
nor U14467 (N_14467,N_11980,N_9836);
xor U14468 (N_14468,N_9371,N_10826);
nor U14469 (N_14469,N_6996,N_7879);
nand U14470 (N_14470,N_6724,N_11973);
xnor U14471 (N_14471,N_7309,N_10867);
or U14472 (N_14472,N_11703,N_8802);
nand U14473 (N_14473,N_6486,N_8211);
nor U14474 (N_14474,N_6910,N_6153);
and U14475 (N_14475,N_8469,N_11615);
nor U14476 (N_14476,N_7032,N_9878);
and U14477 (N_14477,N_7597,N_9070);
or U14478 (N_14478,N_10975,N_6543);
and U14479 (N_14479,N_10346,N_11341);
nand U14480 (N_14480,N_11182,N_11160);
nand U14481 (N_14481,N_10558,N_6723);
xor U14482 (N_14482,N_11848,N_8332);
and U14483 (N_14483,N_8104,N_6775);
nand U14484 (N_14484,N_6174,N_6325);
and U14485 (N_14485,N_7561,N_7738);
and U14486 (N_14486,N_9254,N_7708);
or U14487 (N_14487,N_11983,N_11405);
nand U14488 (N_14488,N_10200,N_10445);
and U14489 (N_14489,N_10198,N_8598);
xnor U14490 (N_14490,N_8764,N_11575);
and U14491 (N_14491,N_9285,N_7290);
or U14492 (N_14492,N_10165,N_9547);
nor U14493 (N_14493,N_7965,N_6624);
xnor U14494 (N_14494,N_6484,N_7583);
nor U14495 (N_14495,N_6152,N_9022);
nand U14496 (N_14496,N_8053,N_7613);
nor U14497 (N_14497,N_9486,N_9214);
xnor U14498 (N_14498,N_8845,N_10961);
xnor U14499 (N_14499,N_6422,N_6022);
nor U14500 (N_14500,N_11873,N_8886);
and U14501 (N_14501,N_7037,N_9571);
nor U14502 (N_14502,N_10561,N_9735);
xor U14503 (N_14503,N_8177,N_9963);
nand U14504 (N_14504,N_10050,N_11417);
and U14505 (N_14505,N_10710,N_10466);
nor U14506 (N_14506,N_9137,N_9482);
and U14507 (N_14507,N_9801,N_6054);
nor U14508 (N_14508,N_8526,N_9672);
nor U14509 (N_14509,N_7992,N_7966);
and U14510 (N_14510,N_7090,N_9698);
nand U14511 (N_14511,N_9654,N_6337);
and U14512 (N_14512,N_10212,N_11930);
or U14513 (N_14513,N_9911,N_6913);
xor U14514 (N_14514,N_11670,N_7953);
nor U14515 (N_14515,N_8309,N_8989);
or U14516 (N_14516,N_10892,N_7196);
xnor U14517 (N_14517,N_6811,N_9674);
nor U14518 (N_14518,N_11157,N_9388);
or U14519 (N_14519,N_9281,N_9979);
or U14520 (N_14520,N_10918,N_11926);
nand U14521 (N_14521,N_7857,N_11321);
nand U14522 (N_14522,N_11186,N_10638);
xor U14523 (N_14523,N_7066,N_11524);
and U14524 (N_14524,N_9080,N_8748);
nor U14525 (N_14525,N_7844,N_6497);
nor U14526 (N_14526,N_8657,N_9006);
xor U14527 (N_14527,N_6320,N_10144);
or U14528 (N_14528,N_6049,N_10688);
xnor U14529 (N_14529,N_8077,N_9544);
xor U14530 (N_14530,N_6586,N_7126);
nor U14531 (N_14531,N_8019,N_10587);
nand U14532 (N_14532,N_6075,N_6105);
nand U14533 (N_14533,N_7067,N_8698);
nor U14534 (N_14534,N_11002,N_9699);
or U14535 (N_14535,N_6285,N_9163);
xor U14536 (N_14536,N_7678,N_8699);
xor U14537 (N_14537,N_10077,N_9555);
nor U14538 (N_14538,N_10569,N_7783);
and U14539 (N_14539,N_6118,N_10024);
or U14540 (N_14540,N_11682,N_8363);
nor U14541 (N_14541,N_8908,N_6686);
xor U14542 (N_14542,N_6248,N_9740);
nor U14543 (N_14543,N_9483,N_6575);
nand U14544 (N_14544,N_10954,N_9955);
and U14545 (N_14545,N_6990,N_8061);
or U14546 (N_14546,N_6505,N_10119);
nand U14547 (N_14547,N_9192,N_7599);
or U14548 (N_14548,N_11759,N_10281);
xor U14549 (N_14549,N_9615,N_9925);
nand U14550 (N_14550,N_6192,N_9623);
or U14551 (N_14551,N_8029,N_6377);
and U14552 (N_14552,N_7976,N_10969);
xor U14553 (N_14553,N_9104,N_8945);
nand U14554 (N_14554,N_6198,N_10777);
nor U14555 (N_14555,N_8562,N_7772);
xnor U14556 (N_14556,N_10596,N_6851);
xnor U14557 (N_14557,N_8525,N_11190);
or U14558 (N_14558,N_11325,N_8127);
or U14559 (N_14559,N_8267,N_11634);
xor U14560 (N_14560,N_10714,N_9824);
nor U14561 (N_14561,N_9064,N_7164);
xnor U14562 (N_14562,N_8407,N_6667);
nand U14563 (N_14563,N_9364,N_7451);
xor U14564 (N_14564,N_9977,N_8756);
nor U14565 (N_14565,N_9844,N_9521);
or U14566 (N_14566,N_11098,N_7385);
nor U14567 (N_14567,N_10420,N_11428);
or U14568 (N_14568,N_9258,N_7139);
xor U14569 (N_14569,N_11854,N_9366);
or U14570 (N_14570,N_11390,N_7669);
nand U14571 (N_14571,N_9952,N_6900);
xnor U14572 (N_14572,N_9326,N_7179);
or U14573 (N_14573,N_11938,N_11213);
nand U14574 (N_14574,N_10842,N_10442);
nor U14575 (N_14575,N_11225,N_11487);
nand U14576 (N_14576,N_8372,N_9151);
nor U14577 (N_14577,N_11067,N_6293);
nand U14578 (N_14578,N_11837,N_10214);
xnor U14579 (N_14579,N_6644,N_11365);
xor U14580 (N_14580,N_6472,N_9908);
nor U14581 (N_14581,N_9750,N_9998);
nand U14582 (N_14582,N_8615,N_10623);
or U14583 (N_14583,N_8450,N_8206);
and U14584 (N_14584,N_10870,N_6195);
or U14585 (N_14585,N_10357,N_11177);
nand U14586 (N_14586,N_6444,N_9653);
nor U14587 (N_14587,N_10460,N_7679);
and U14588 (N_14588,N_9451,N_11786);
nand U14589 (N_14589,N_6470,N_7871);
xnor U14590 (N_14590,N_9240,N_9681);
or U14591 (N_14591,N_7742,N_10069);
and U14592 (N_14592,N_10759,N_8082);
nand U14593 (N_14593,N_10783,N_9155);
nor U14594 (N_14594,N_9560,N_7923);
and U14595 (N_14595,N_6102,N_8318);
and U14596 (N_14596,N_10676,N_7820);
nor U14597 (N_14597,N_8005,N_7773);
and U14598 (N_14598,N_9294,N_9718);
nor U14599 (N_14599,N_6108,N_9969);
and U14600 (N_14600,N_7824,N_9983);
and U14601 (N_14601,N_6588,N_11264);
or U14602 (N_14602,N_8307,N_6235);
or U14603 (N_14603,N_10823,N_11735);
xor U14604 (N_14604,N_10430,N_6354);
xnor U14605 (N_14605,N_8373,N_8824);
or U14606 (N_14606,N_6860,N_6948);
xnor U14607 (N_14607,N_10450,N_7107);
nand U14608 (N_14608,N_7397,N_11237);
nor U14609 (N_14609,N_8922,N_11091);
nand U14610 (N_14610,N_8554,N_8008);
nand U14611 (N_14611,N_10184,N_10113);
xnor U14612 (N_14612,N_8269,N_9158);
xnor U14613 (N_14613,N_7850,N_8345);
xnor U14614 (N_14614,N_6006,N_10027);
nor U14615 (N_14615,N_10344,N_8233);
nor U14616 (N_14616,N_8614,N_8194);
and U14617 (N_14617,N_11749,N_9880);
or U14618 (N_14618,N_10651,N_8979);
and U14619 (N_14619,N_7253,N_8880);
nand U14620 (N_14620,N_6519,N_11894);
xnor U14621 (N_14621,N_6451,N_9028);
or U14622 (N_14622,N_9087,N_11480);
nor U14623 (N_14623,N_9608,N_10057);
or U14624 (N_14624,N_7904,N_7328);
and U14625 (N_14625,N_9322,N_10019);
nor U14626 (N_14626,N_6532,N_11914);
nand U14627 (N_14627,N_9394,N_11147);
xor U14628 (N_14628,N_10462,N_6978);
or U14629 (N_14629,N_9966,N_10608);
or U14630 (N_14630,N_11811,N_8451);
xor U14631 (N_14631,N_10796,N_8595);
or U14632 (N_14632,N_8817,N_10837);
or U14633 (N_14633,N_8867,N_10562);
and U14634 (N_14634,N_8902,N_11337);
nand U14635 (N_14635,N_11958,N_11887);
nand U14636 (N_14636,N_9619,N_11739);
xnor U14637 (N_14637,N_10225,N_10634);
nor U14638 (N_14638,N_8044,N_9184);
nor U14639 (N_14639,N_7804,N_7557);
and U14640 (N_14640,N_10983,N_6596);
or U14641 (N_14641,N_10348,N_8993);
or U14642 (N_14642,N_10607,N_9355);
or U14643 (N_14643,N_7490,N_7469);
nand U14644 (N_14644,N_8224,N_7302);
xnor U14645 (N_14645,N_9814,N_8919);
and U14646 (N_14646,N_6407,N_10773);
nand U14647 (N_14647,N_6684,N_8618);
xor U14648 (N_14648,N_8588,N_10405);
or U14649 (N_14649,N_11444,N_10900);
nand U14650 (N_14650,N_7222,N_7794);
and U14651 (N_14651,N_7036,N_8680);
and U14652 (N_14652,N_8291,N_8953);
nor U14653 (N_14653,N_8703,N_11896);
xnor U14654 (N_14654,N_9585,N_10267);
and U14655 (N_14655,N_11741,N_8355);
and U14656 (N_14656,N_8297,N_10726);
or U14657 (N_14657,N_7796,N_10523);
nand U14658 (N_14658,N_9488,N_9154);
and U14659 (N_14659,N_11882,N_10321);
nor U14660 (N_14660,N_7440,N_9863);
xor U14661 (N_14661,N_6760,N_9229);
and U14662 (N_14662,N_7226,N_11995);
nand U14663 (N_14663,N_10426,N_6704);
nand U14664 (N_14664,N_6612,N_7587);
and U14665 (N_14665,N_7999,N_9024);
xor U14666 (N_14666,N_11788,N_7946);
and U14667 (N_14667,N_6071,N_8212);
or U14668 (N_14668,N_6843,N_7082);
and U14669 (N_14669,N_7980,N_10579);
xnor U14670 (N_14670,N_8582,N_6745);
and U14671 (N_14671,N_6359,N_10135);
or U14672 (N_14672,N_8716,N_8045);
or U14673 (N_14673,N_6522,N_8964);
and U14674 (N_14674,N_11655,N_8409);
and U14675 (N_14675,N_9954,N_8580);
xor U14676 (N_14676,N_11145,N_9688);
nand U14677 (N_14677,N_7951,N_11292);
nand U14678 (N_14678,N_8458,N_8457);
or U14679 (N_14679,N_10204,N_9828);
nand U14680 (N_14680,N_10036,N_9128);
nand U14681 (N_14681,N_10552,N_7446);
nor U14682 (N_14682,N_11748,N_11689);
nand U14683 (N_14683,N_8969,N_9211);
or U14684 (N_14684,N_8865,N_11677);
nor U14685 (N_14685,N_9670,N_9959);
xnor U14686 (N_14686,N_11685,N_7350);
or U14687 (N_14687,N_9386,N_8929);
xor U14688 (N_14688,N_9888,N_10525);
or U14689 (N_14689,N_11418,N_7600);
and U14690 (N_14690,N_6711,N_9282);
or U14691 (N_14691,N_10920,N_7378);
xnor U14692 (N_14692,N_9957,N_10627);
or U14693 (N_14693,N_6653,N_11217);
nand U14694 (N_14694,N_8220,N_10034);
xnor U14695 (N_14695,N_7019,N_9886);
nor U14696 (N_14696,N_11135,N_7620);
nand U14697 (N_14697,N_8248,N_9119);
nor U14698 (N_14698,N_8682,N_7123);
xor U14699 (N_14699,N_10505,N_7537);
nand U14700 (N_14700,N_10871,N_7778);
nor U14701 (N_14701,N_10809,N_6018);
xor U14702 (N_14702,N_10744,N_7013);
nor U14703 (N_14703,N_9936,N_9124);
xnor U14704 (N_14704,N_6597,N_11921);
nand U14705 (N_14705,N_10266,N_6685);
or U14706 (N_14706,N_10597,N_7165);
or U14707 (N_14707,N_9392,N_11986);
and U14708 (N_14708,N_9937,N_11029);
or U14709 (N_14709,N_10234,N_9096);
xnor U14710 (N_14710,N_9703,N_11094);
xor U14711 (N_14711,N_10468,N_7860);
nand U14712 (N_14712,N_6411,N_7441);
and U14713 (N_14713,N_7507,N_11805);
xnor U14714 (N_14714,N_11174,N_7585);
xor U14715 (N_14715,N_10538,N_10621);
or U14716 (N_14716,N_10403,N_10127);
nand U14717 (N_14717,N_11156,N_11196);
nand U14718 (N_14718,N_9533,N_6567);
or U14719 (N_14719,N_10835,N_11989);
nor U14720 (N_14720,N_7511,N_7506);
xor U14721 (N_14721,N_11132,N_11432);
and U14722 (N_14722,N_11446,N_7567);
or U14723 (N_14723,N_10524,N_9574);
or U14724 (N_14724,N_11206,N_10657);
nand U14725 (N_14725,N_8356,N_10361);
and U14726 (N_14726,N_11155,N_7270);
and U14727 (N_14727,N_8878,N_8690);
nor U14728 (N_14728,N_10375,N_8449);
nand U14729 (N_14729,N_8215,N_6998);
nand U14730 (N_14730,N_9001,N_10095);
or U14731 (N_14731,N_7003,N_6930);
or U14732 (N_14732,N_6880,N_8832);
xor U14733 (N_14733,N_10236,N_8971);
nand U14734 (N_14734,N_9316,N_11734);
nor U14735 (N_14735,N_9991,N_9994);
and U14736 (N_14736,N_10743,N_11992);
nand U14737 (N_14737,N_11084,N_8351);
nand U14738 (N_14738,N_8637,N_9261);
xnor U14739 (N_14739,N_8246,N_8661);
or U14740 (N_14740,N_6392,N_11089);
xnor U14741 (N_14741,N_6215,N_11371);
nand U14742 (N_14742,N_7098,N_6623);
and U14743 (N_14743,N_11080,N_9387);
and U14744 (N_14744,N_6389,N_7626);
xor U14745 (N_14745,N_8463,N_10147);
nor U14746 (N_14746,N_9301,N_6081);
nand U14747 (N_14747,N_8454,N_7184);
or U14748 (N_14748,N_6708,N_9892);
xnor U14749 (N_14749,N_9126,N_10884);
or U14750 (N_14750,N_10042,N_6477);
xnor U14751 (N_14751,N_8198,N_11367);
or U14752 (N_14752,N_6468,N_7621);
nor U14753 (N_14753,N_9641,N_11499);
xor U14754 (N_14754,N_6297,N_10195);
or U14755 (N_14755,N_11510,N_10584);
and U14756 (N_14756,N_11494,N_10224);
xor U14757 (N_14757,N_9592,N_8488);
xnor U14758 (N_14758,N_7380,N_11599);
and U14759 (N_14759,N_10421,N_8545);
or U14760 (N_14760,N_11550,N_9661);
xor U14761 (N_14761,N_10899,N_9115);
nand U14762 (N_14762,N_6391,N_9027);
or U14763 (N_14763,N_8011,N_7645);
and U14764 (N_14764,N_8455,N_11885);
and U14765 (N_14765,N_7724,N_6722);
or U14766 (N_14766,N_7694,N_7532);
or U14767 (N_14767,N_6077,N_6501);
and U14768 (N_14768,N_10865,N_11017);
xor U14769 (N_14769,N_8749,N_11679);
xnor U14770 (N_14770,N_10390,N_11381);
nor U14771 (N_14771,N_8791,N_11172);
or U14772 (N_14772,N_9033,N_11133);
or U14773 (N_14773,N_11162,N_6193);
nand U14774 (N_14774,N_8872,N_7437);
nor U14775 (N_14775,N_10381,N_7919);
and U14776 (N_14776,N_11867,N_7391);
xnor U14777 (N_14777,N_7970,N_6980);
nor U14778 (N_14778,N_9279,N_9778);
xnor U14779 (N_14779,N_9604,N_8016);
nand U14780 (N_14780,N_7389,N_11752);
and U14781 (N_14781,N_7672,N_9579);
and U14782 (N_14782,N_11686,N_6554);
or U14783 (N_14783,N_6228,N_8928);
xnor U14784 (N_14784,N_8091,N_8140);
or U14785 (N_14785,N_10901,N_10506);
xor U14786 (N_14786,N_8257,N_8915);
and U14787 (N_14787,N_7939,N_10951);
or U14788 (N_14788,N_6857,N_11027);
nand U14789 (N_14789,N_8384,N_10062);
or U14790 (N_14790,N_9827,N_10416);
or U14791 (N_14791,N_9098,N_6180);
or U14792 (N_14792,N_8349,N_6370);
or U14793 (N_14793,N_6259,N_7472);
nor U14794 (N_14794,N_7715,N_11169);
or U14795 (N_14795,N_8181,N_9423);
nand U14796 (N_14796,N_10503,N_8255);
nor U14797 (N_14797,N_7388,N_8379);
and U14798 (N_14798,N_8348,N_10075);
nor U14799 (N_14799,N_6119,N_9175);
xor U14800 (N_14800,N_7304,N_7356);
and U14801 (N_14801,N_6752,N_11400);
and U14802 (N_14802,N_7718,N_7461);
nor U14803 (N_14803,N_7901,N_7436);
nor U14804 (N_14804,N_7762,N_8960);
and U14805 (N_14805,N_7961,N_8222);
and U14806 (N_14806,N_8760,N_7836);
nor U14807 (N_14807,N_10511,N_8057);
nand U14808 (N_14808,N_8036,N_10978);
or U14809 (N_14809,N_9549,N_8490);
and U14810 (N_14810,N_7996,N_6804);
or U14811 (N_14811,N_7885,N_9026);
xnor U14812 (N_14812,N_8863,N_8977);
nand U14813 (N_14813,N_9283,N_11784);
or U14814 (N_14814,N_6768,N_10932);
nor U14815 (N_14815,N_11508,N_11912);
or U14816 (N_14816,N_9461,N_6516);
and U14817 (N_14817,N_11626,N_6719);
xnor U14818 (N_14818,N_10898,N_8529);
xor U14819 (N_14819,N_9561,N_6524);
nand U14820 (N_14820,N_9076,N_6399);
or U14821 (N_14821,N_11962,N_11763);
nor U14822 (N_14822,N_10718,N_11025);
xor U14823 (N_14823,N_7305,N_7986);
nand U14824 (N_14824,N_11687,N_11231);
nand U14825 (N_14825,N_6480,N_11518);
nand U14826 (N_14826,N_6892,N_11165);
nor U14827 (N_14827,N_11241,N_8951);
and U14828 (N_14828,N_6275,N_7468);
and U14829 (N_14829,N_7474,N_10554);
and U14830 (N_14830,N_10035,N_6574);
xnor U14831 (N_14831,N_7275,N_9920);
and U14832 (N_14832,N_6289,N_6921);
or U14833 (N_14833,N_7187,N_7333);
nor U14834 (N_14834,N_6095,N_10217);
xor U14835 (N_14835,N_8639,N_9003);
nor U14836 (N_14836,N_6234,N_11077);
nand U14837 (N_14837,N_9593,N_7173);
and U14838 (N_14838,N_9348,N_9629);
nand U14839 (N_14839,N_11245,N_7888);
and U14840 (N_14840,N_6442,N_8765);
nor U14841 (N_14841,N_7868,N_11130);
xor U14842 (N_14842,N_7034,N_11280);
and U14843 (N_14843,N_9297,N_10286);
nand U14844 (N_14844,N_6222,N_7921);
nand U14845 (N_14845,N_10769,N_7962);
nor U14846 (N_14846,N_10443,N_8666);
and U14847 (N_14847,N_6351,N_7754);
nand U14848 (N_14848,N_11846,N_8312);
nand U14849 (N_14849,N_10618,N_10295);
or U14850 (N_14850,N_9582,N_9183);
and U14851 (N_14851,N_10672,N_9167);
nor U14852 (N_14852,N_6030,N_8305);
or U14853 (N_14853,N_6226,N_11416);
xor U14854 (N_14854,N_6869,N_6060);
nand U14855 (N_14855,N_8720,N_8048);
or U14856 (N_14856,N_7040,N_7149);
nand U14857 (N_14857,N_11834,N_9177);
xor U14858 (N_14858,N_7635,N_9401);
nor U14859 (N_14859,N_11538,N_6599);
nor U14860 (N_14860,N_9256,N_8745);
xor U14861 (N_14861,N_11119,N_6257);
and U14862 (N_14862,N_10073,N_11688);
or U14863 (N_14863,N_8226,N_6132);
nand U14864 (N_14864,N_6855,N_11795);
xor U14865 (N_14865,N_6641,N_8729);
or U14866 (N_14866,N_8790,N_8924);
xor U14867 (N_14867,N_6962,N_6750);
or U14868 (N_14868,N_11200,N_8334);
nor U14869 (N_14869,N_6825,N_11651);
nand U14870 (N_14870,N_11632,N_11941);
nor U14871 (N_14871,N_7958,N_7114);
and U14872 (N_14872,N_10611,N_9405);
or U14873 (N_14873,N_10482,N_10362);
and U14874 (N_14874,N_6452,N_8837);
nor U14875 (N_14875,N_8619,N_10913);
xnor U14876 (N_14876,N_8674,N_10141);
xnor U14877 (N_14877,N_6959,N_6055);
nand U14878 (N_14878,N_6958,N_11561);
or U14879 (N_14879,N_10507,N_7830);
and U14880 (N_14880,N_8644,N_10891);
and U14881 (N_14881,N_8026,N_7241);
xnor U14882 (N_14882,N_6517,N_6849);
nand U14883 (N_14883,N_7667,N_9805);
nand U14884 (N_14884,N_7509,N_9139);
and U14885 (N_14885,N_9860,N_6798);
nand U14886 (N_14886,N_10476,N_7485);
nand U14887 (N_14887,N_11170,N_11512);
nor U14888 (N_14888,N_8491,N_8152);
nor U14889 (N_14889,N_6537,N_7326);
nand U14890 (N_14890,N_10437,N_6870);
nor U14891 (N_14891,N_7526,N_8947);
or U14892 (N_14892,N_7690,N_6640);
nor U14893 (N_14893,N_10927,N_11037);
or U14894 (N_14894,N_9314,N_8402);
nand U14895 (N_14895,N_7565,N_7931);
nand U14896 (N_14896,N_7893,N_6080);
and U14897 (N_14897,N_6432,N_6514);
and U14898 (N_14898,N_9918,N_9826);
nand U14899 (N_14899,N_9161,N_10807);
nand U14900 (N_14900,N_11019,N_7282);
and U14901 (N_14901,N_9501,N_8763);
nor U14902 (N_14902,N_11058,N_8509);
or U14903 (N_14903,N_6610,N_8034);
nand U14904 (N_14904,N_9014,N_9517);
and U14905 (N_14905,N_9293,N_6715);
nand U14906 (N_14906,N_11347,N_10290);
nand U14907 (N_14907,N_8740,N_10504);
or U14908 (N_14908,N_7243,N_7917);
xnor U14909 (N_14909,N_11863,N_7006);
nand U14910 (N_14910,N_11272,N_9520);
xor U14911 (N_14911,N_7685,N_9231);
or U14912 (N_14912,N_7648,N_10864);
and U14913 (N_14913,N_7652,N_6576);
xor U14914 (N_14914,N_7831,N_7466);
or U14915 (N_14915,N_11928,N_6084);
or U14916 (N_14916,N_11345,N_11951);
or U14917 (N_14917,N_7851,N_7702);
and U14918 (N_14918,N_11290,N_8378);
xnor U14919 (N_14919,N_10595,N_6101);
nand U14920 (N_14920,N_9981,N_10086);
or U14921 (N_14921,N_9248,N_9009);
nor U14922 (N_14922,N_9439,N_6123);
or U14923 (N_14923,N_8138,N_8594);
nand U14924 (N_14924,N_9400,N_8532);
and U14925 (N_14925,N_6271,N_6802);
nor U14926 (N_14926,N_7554,N_9265);
xnor U14927 (N_14927,N_9524,N_8773);
or U14928 (N_14928,N_6794,N_6426);
or U14929 (N_14929,N_8744,N_7973);
nor U14930 (N_14930,N_10096,N_8954);
nand U14931 (N_14931,N_7101,N_9384);
nand U14932 (N_14932,N_7769,N_6165);
or U14933 (N_14933,N_9352,N_9029);
xor U14934 (N_14934,N_8386,N_8590);
and U14935 (N_14935,N_9710,N_9449);
nand U14936 (N_14936,N_7641,N_9320);
xor U14937 (N_14937,N_10176,N_9274);
nand U14938 (N_14938,N_6661,N_6882);
nand U14939 (N_14939,N_7729,N_11460);
and U14940 (N_14940,N_8466,N_7627);
xnor U14941 (N_14941,N_10720,N_7550);
nor U14942 (N_14942,N_10810,N_10753);
and U14943 (N_14943,N_7911,N_6295);
or U14944 (N_14944,N_10337,N_6024);
or U14945 (N_14945,N_7947,N_9774);
nor U14946 (N_14946,N_9448,N_11408);
nor U14947 (N_14947,N_8742,N_10244);
nor U14948 (N_14948,N_9017,N_8600);
or U14949 (N_14949,N_8456,N_6943);
or U14950 (N_14950,N_9987,N_10896);
nand U14951 (N_14951,N_6339,N_11267);
xnor U14952 (N_14952,N_10965,N_8090);
or U14953 (N_14953,N_11793,N_7190);
nand U14954 (N_14954,N_8648,N_6187);
xnor U14955 (N_14955,N_8567,N_7137);
and U14956 (N_14956,N_6087,N_9370);
nor U14957 (N_14957,N_6754,N_11379);
or U14958 (N_14958,N_8776,N_9847);
xor U14959 (N_14959,N_7263,N_9522);
nand U14960 (N_14960,N_11864,N_9633);
nor U14961 (N_14961,N_7848,N_11195);
xor U14962 (N_14962,N_9237,N_7858);
xor U14963 (N_14963,N_6872,N_9198);
and U14964 (N_14964,N_7236,N_7058);
xnor U14965 (N_14965,N_8685,N_10883);
and U14966 (N_14966,N_11103,N_8148);
or U14967 (N_14967,N_9830,N_11415);
nor U14968 (N_14968,N_9798,N_11917);
and U14969 (N_14969,N_6738,N_9572);
or U14970 (N_14970,N_11437,N_10619);
nor U14971 (N_14971,N_7154,N_6788);
nor U14972 (N_14972,N_7595,N_8086);
or U14973 (N_14973,N_7612,N_7128);
and U14974 (N_14974,N_8706,N_7439);
nand U14975 (N_14975,N_7790,N_9103);
or U14976 (N_14976,N_6137,N_11762);
or U14977 (N_14977,N_9785,N_11819);
nand U14978 (N_14978,N_9941,N_10848);
nand U14979 (N_14979,N_11277,N_6730);
xor U14980 (N_14980,N_6716,N_8722);
nand U14981 (N_14981,N_11033,N_6488);
or U14982 (N_14982,N_10327,N_7761);
or U14983 (N_14983,N_7576,N_6247);
nor U14984 (N_14984,N_9159,N_7065);
and U14985 (N_14985,N_8429,N_8209);
xor U14986 (N_14986,N_8341,N_8980);
and U14987 (N_14987,N_6148,N_8559);
or U14988 (N_14988,N_10111,N_7854);
nand U14989 (N_14989,N_6571,N_10655);
xnor U14990 (N_14990,N_11822,N_9066);
nand U14991 (N_14991,N_7216,N_11729);
or U14992 (N_14992,N_10973,N_7828);
and U14993 (N_14993,N_10382,N_8023);
nor U14994 (N_14994,N_6266,N_9659);
and U14995 (N_14995,N_9315,N_11825);
or U14996 (N_14996,N_6741,N_9363);
xnor U14997 (N_14997,N_10919,N_8031);
and U14998 (N_14998,N_9806,N_10546);
nor U14999 (N_14999,N_6508,N_7189);
xor U15000 (N_15000,N_11594,N_7946);
xor U15001 (N_15001,N_9802,N_11716);
nor U15002 (N_15002,N_9181,N_8454);
xor U15003 (N_15003,N_8849,N_7564);
xor U15004 (N_15004,N_7140,N_9481);
and U15005 (N_15005,N_11519,N_7020);
xnor U15006 (N_15006,N_11664,N_6020);
and U15007 (N_15007,N_8957,N_11142);
or U15008 (N_15008,N_10553,N_6963);
and U15009 (N_15009,N_10831,N_8768);
nor U15010 (N_15010,N_10424,N_8730);
and U15011 (N_15011,N_8584,N_10384);
and U15012 (N_15012,N_11183,N_11734);
nor U15013 (N_15013,N_6191,N_10171);
or U15014 (N_15014,N_8201,N_9726);
and U15015 (N_15015,N_6075,N_9812);
and U15016 (N_15016,N_6108,N_9455);
and U15017 (N_15017,N_7227,N_9512);
xnor U15018 (N_15018,N_6825,N_8697);
and U15019 (N_15019,N_8950,N_11421);
or U15020 (N_15020,N_6979,N_9576);
nor U15021 (N_15021,N_9211,N_9120);
nand U15022 (N_15022,N_9689,N_6256);
nor U15023 (N_15023,N_7658,N_8296);
xor U15024 (N_15024,N_11431,N_9142);
xor U15025 (N_15025,N_6908,N_9885);
or U15026 (N_15026,N_8925,N_6171);
nand U15027 (N_15027,N_8410,N_9059);
xor U15028 (N_15028,N_7984,N_8393);
nor U15029 (N_15029,N_8982,N_9869);
or U15030 (N_15030,N_10846,N_6337);
xnor U15031 (N_15031,N_10962,N_7608);
and U15032 (N_15032,N_11300,N_7688);
or U15033 (N_15033,N_8996,N_7361);
nor U15034 (N_15034,N_11145,N_9463);
nand U15035 (N_15035,N_10173,N_11402);
xnor U15036 (N_15036,N_10509,N_7299);
nand U15037 (N_15037,N_8589,N_7025);
nor U15038 (N_15038,N_6962,N_9581);
or U15039 (N_15039,N_7123,N_10717);
nor U15040 (N_15040,N_11440,N_9314);
and U15041 (N_15041,N_6207,N_6575);
or U15042 (N_15042,N_9211,N_10858);
or U15043 (N_15043,N_8873,N_9115);
or U15044 (N_15044,N_8885,N_10047);
xnor U15045 (N_15045,N_7742,N_7372);
xnor U15046 (N_15046,N_6034,N_8145);
xnor U15047 (N_15047,N_10865,N_7248);
nor U15048 (N_15048,N_8820,N_6596);
or U15049 (N_15049,N_11627,N_10544);
xnor U15050 (N_15050,N_8060,N_6532);
nand U15051 (N_15051,N_11343,N_9555);
xnor U15052 (N_15052,N_9824,N_7726);
nor U15053 (N_15053,N_7170,N_9719);
nor U15054 (N_15054,N_8457,N_10656);
nor U15055 (N_15055,N_6333,N_9602);
and U15056 (N_15056,N_7842,N_10561);
nand U15057 (N_15057,N_8112,N_8865);
or U15058 (N_15058,N_7760,N_10272);
nand U15059 (N_15059,N_11748,N_8356);
and U15060 (N_15060,N_6934,N_10173);
and U15061 (N_15061,N_10584,N_11760);
or U15062 (N_15062,N_6355,N_10906);
and U15063 (N_15063,N_7388,N_10167);
xnor U15064 (N_15064,N_6127,N_9613);
nand U15065 (N_15065,N_11139,N_9094);
and U15066 (N_15066,N_10365,N_9412);
or U15067 (N_15067,N_8769,N_8346);
nand U15068 (N_15068,N_7568,N_11638);
nor U15069 (N_15069,N_9525,N_10818);
and U15070 (N_15070,N_11004,N_9897);
nand U15071 (N_15071,N_10327,N_7613);
and U15072 (N_15072,N_11773,N_8867);
nor U15073 (N_15073,N_10180,N_11945);
nand U15074 (N_15074,N_6876,N_8439);
nor U15075 (N_15075,N_8079,N_6021);
and U15076 (N_15076,N_10088,N_11758);
nor U15077 (N_15077,N_8102,N_8773);
or U15078 (N_15078,N_10996,N_7677);
xor U15079 (N_15079,N_7496,N_10784);
or U15080 (N_15080,N_10968,N_9622);
nor U15081 (N_15081,N_7764,N_7027);
and U15082 (N_15082,N_11912,N_6738);
or U15083 (N_15083,N_9041,N_10180);
xor U15084 (N_15084,N_11523,N_9176);
nor U15085 (N_15085,N_6629,N_10963);
nor U15086 (N_15086,N_8717,N_10246);
xnor U15087 (N_15087,N_9328,N_6182);
nor U15088 (N_15088,N_6226,N_8087);
and U15089 (N_15089,N_8958,N_6456);
xnor U15090 (N_15090,N_8722,N_7439);
and U15091 (N_15091,N_11671,N_7627);
nor U15092 (N_15092,N_10272,N_8533);
and U15093 (N_15093,N_7077,N_7149);
or U15094 (N_15094,N_10182,N_9073);
nor U15095 (N_15095,N_8399,N_11614);
and U15096 (N_15096,N_6038,N_8070);
xnor U15097 (N_15097,N_7872,N_7707);
nor U15098 (N_15098,N_6559,N_9905);
nand U15099 (N_15099,N_11733,N_11250);
nor U15100 (N_15100,N_7265,N_9010);
nor U15101 (N_15101,N_6571,N_9766);
or U15102 (N_15102,N_9148,N_9979);
and U15103 (N_15103,N_7332,N_6069);
nor U15104 (N_15104,N_9149,N_6019);
or U15105 (N_15105,N_7580,N_9415);
nand U15106 (N_15106,N_6240,N_10896);
or U15107 (N_15107,N_10021,N_9457);
or U15108 (N_15108,N_8578,N_6005);
or U15109 (N_15109,N_11431,N_6369);
nand U15110 (N_15110,N_11197,N_11485);
nand U15111 (N_15111,N_7162,N_8959);
and U15112 (N_15112,N_8459,N_9732);
nand U15113 (N_15113,N_8073,N_8079);
nand U15114 (N_15114,N_11746,N_10407);
xor U15115 (N_15115,N_11539,N_11564);
and U15116 (N_15116,N_8110,N_8221);
nand U15117 (N_15117,N_10485,N_9003);
and U15118 (N_15118,N_10643,N_8309);
nor U15119 (N_15119,N_9623,N_8059);
nor U15120 (N_15120,N_8970,N_7678);
nand U15121 (N_15121,N_11273,N_8437);
or U15122 (N_15122,N_8056,N_6848);
xnor U15123 (N_15123,N_11281,N_8283);
nor U15124 (N_15124,N_8989,N_10956);
nand U15125 (N_15125,N_11217,N_10486);
nand U15126 (N_15126,N_8283,N_11092);
nor U15127 (N_15127,N_8721,N_11941);
nor U15128 (N_15128,N_6549,N_8386);
or U15129 (N_15129,N_6292,N_11794);
or U15130 (N_15130,N_11886,N_6492);
or U15131 (N_15131,N_11882,N_10999);
xor U15132 (N_15132,N_7703,N_6835);
nand U15133 (N_15133,N_7845,N_6297);
xnor U15134 (N_15134,N_11936,N_9569);
and U15135 (N_15135,N_9926,N_6290);
or U15136 (N_15136,N_7255,N_8764);
nor U15137 (N_15137,N_10607,N_9648);
nand U15138 (N_15138,N_8366,N_11067);
nand U15139 (N_15139,N_11842,N_11640);
xnor U15140 (N_15140,N_8506,N_9195);
and U15141 (N_15141,N_6127,N_7633);
nand U15142 (N_15142,N_8989,N_11780);
nor U15143 (N_15143,N_7792,N_9629);
nor U15144 (N_15144,N_7363,N_11750);
nand U15145 (N_15145,N_11451,N_7942);
xor U15146 (N_15146,N_8885,N_6647);
nor U15147 (N_15147,N_6014,N_9798);
nor U15148 (N_15148,N_10377,N_10688);
or U15149 (N_15149,N_6982,N_7471);
and U15150 (N_15150,N_9049,N_11288);
nor U15151 (N_15151,N_7517,N_11592);
xor U15152 (N_15152,N_6032,N_10271);
xor U15153 (N_15153,N_10703,N_8427);
nand U15154 (N_15154,N_9144,N_11294);
and U15155 (N_15155,N_11942,N_10313);
xor U15156 (N_15156,N_7304,N_10483);
nand U15157 (N_15157,N_8968,N_7882);
nor U15158 (N_15158,N_10479,N_9944);
or U15159 (N_15159,N_9262,N_9995);
and U15160 (N_15160,N_10488,N_10241);
xnor U15161 (N_15161,N_10743,N_9100);
and U15162 (N_15162,N_6756,N_6144);
or U15163 (N_15163,N_7910,N_10801);
or U15164 (N_15164,N_6021,N_10240);
xor U15165 (N_15165,N_9303,N_9098);
xnor U15166 (N_15166,N_11542,N_6281);
nor U15167 (N_15167,N_6011,N_10212);
nand U15168 (N_15168,N_7483,N_6204);
or U15169 (N_15169,N_8399,N_11096);
nor U15170 (N_15170,N_6118,N_7111);
or U15171 (N_15171,N_6693,N_8599);
nor U15172 (N_15172,N_8516,N_8771);
and U15173 (N_15173,N_7976,N_9718);
xor U15174 (N_15174,N_6095,N_7142);
or U15175 (N_15175,N_6358,N_8355);
or U15176 (N_15176,N_9629,N_9554);
or U15177 (N_15177,N_7847,N_8331);
nand U15178 (N_15178,N_6900,N_7415);
xor U15179 (N_15179,N_7502,N_9181);
and U15180 (N_15180,N_10485,N_11609);
and U15181 (N_15181,N_11251,N_7101);
and U15182 (N_15182,N_11764,N_11000);
or U15183 (N_15183,N_9402,N_7407);
nand U15184 (N_15184,N_6669,N_7735);
xor U15185 (N_15185,N_7384,N_10158);
and U15186 (N_15186,N_9736,N_8591);
xor U15187 (N_15187,N_9790,N_10130);
or U15188 (N_15188,N_10665,N_10224);
nor U15189 (N_15189,N_9552,N_7180);
or U15190 (N_15190,N_7858,N_10376);
nand U15191 (N_15191,N_9569,N_11279);
xor U15192 (N_15192,N_11351,N_7980);
or U15193 (N_15193,N_6274,N_10785);
nand U15194 (N_15194,N_9437,N_6654);
or U15195 (N_15195,N_11154,N_8609);
and U15196 (N_15196,N_10246,N_6566);
nand U15197 (N_15197,N_10965,N_11080);
xor U15198 (N_15198,N_8816,N_6939);
xnor U15199 (N_15199,N_11646,N_6098);
or U15200 (N_15200,N_7815,N_11656);
xor U15201 (N_15201,N_7453,N_11114);
xor U15202 (N_15202,N_8484,N_11641);
nand U15203 (N_15203,N_11923,N_8859);
xnor U15204 (N_15204,N_10303,N_6832);
nand U15205 (N_15205,N_11133,N_9516);
nand U15206 (N_15206,N_7264,N_10255);
nor U15207 (N_15207,N_6515,N_9942);
nor U15208 (N_15208,N_8227,N_8056);
and U15209 (N_15209,N_11688,N_10623);
or U15210 (N_15210,N_7082,N_8325);
and U15211 (N_15211,N_11658,N_7836);
and U15212 (N_15212,N_9164,N_8597);
or U15213 (N_15213,N_6688,N_6305);
nor U15214 (N_15214,N_8099,N_9598);
nor U15215 (N_15215,N_9527,N_10433);
or U15216 (N_15216,N_6161,N_9312);
nor U15217 (N_15217,N_9928,N_7671);
nor U15218 (N_15218,N_7639,N_6683);
or U15219 (N_15219,N_6655,N_6426);
or U15220 (N_15220,N_11889,N_10581);
xnor U15221 (N_15221,N_10189,N_9017);
xor U15222 (N_15222,N_9982,N_10419);
nand U15223 (N_15223,N_8406,N_11955);
nand U15224 (N_15224,N_7129,N_7804);
and U15225 (N_15225,N_7085,N_9630);
xor U15226 (N_15226,N_8140,N_8823);
and U15227 (N_15227,N_11763,N_9031);
and U15228 (N_15228,N_7034,N_8286);
and U15229 (N_15229,N_9540,N_7290);
or U15230 (N_15230,N_6489,N_7259);
nor U15231 (N_15231,N_8983,N_7155);
or U15232 (N_15232,N_6115,N_9251);
and U15233 (N_15233,N_9703,N_10152);
or U15234 (N_15234,N_11491,N_11511);
or U15235 (N_15235,N_8490,N_10258);
and U15236 (N_15236,N_10958,N_10688);
and U15237 (N_15237,N_11618,N_9784);
nor U15238 (N_15238,N_9621,N_6185);
or U15239 (N_15239,N_10328,N_7087);
nand U15240 (N_15240,N_10238,N_11110);
xnor U15241 (N_15241,N_9010,N_6700);
xnor U15242 (N_15242,N_10849,N_9513);
and U15243 (N_15243,N_9372,N_11483);
and U15244 (N_15244,N_9256,N_11294);
nand U15245 (N_15245,N_10850,N_11377);
or U15246 (N_15246,N_11119,N_7955);
nand U15247 (N_15247,N_7475,N_7502);
and U15248 (N_15248,N_6681,N_7550);
and U15249 (N_15249,N_11649,N_8345);
or U15250 (N_15250,N_6057,N_11945);
nor U15251 (N_15251,N_9582,N_11903);
nand U15252 (N_15252,N_6992,N_9208);
nor U15253 (N_15253,N_7487,N_9067);
nand U15254 (N_15254,N_11131,N_7109);
nand U15255 (N_15255,N_7777,N_10107);
and U15256 (N_15256,N_8133,N_9102);
nand U15257 (N_15257,N_11005,N_7587);
nand U15258 (N_15258,N_7110,N_6999);
nor U15259 (N_15259,N_10786,N_11790);
nor U15260 (N_15260,N_8243,N_9971);
or U15261 (N_15261,N_11520,N_9088);
nor U15262 (N_15262,N_8875,N_8905);
or U15263 (N_15263,N_7682,N_7188);
nand U15264 (N_15264,N_8791,N_10773);
xnor U15265 (N_15265,N_9852,N_8279);
nor U15266 (N_15266,N_6877,N_7499);
and U15267 (N_15267,N_10059,N_10518);
nand U15268 (N_15268,N_7130,N_7251);
nand U15269 (N_15269,N_9407,N_7741);
nand U15270 (N_15270,N_6934,N_10060);
and U15271 (N_15271,N_7308,N_6705);
nand U15272 (N_15272,N_11205,N_11569);
nand U15273 (N_15273,N_9528,N_6802);
or U15274 (N_15274,N_7733,N_10559);
nor U15275 (N_15275,N_11951,N_8539);
and U15276 (N_15276,N_11018,N_9475);
nor U15277 (N_15277,N_7168,N_7801);
xor U15278 (N_15278,N_9244,N_9038);
or U15279 (N_15279,N_6213,N_9627);
xor U15280 (N_15280,N_9565,N_9173);
or U15281 (N_15281,N_9134,N_11663);
nand U15282 (N_15282,N_8304,N_11594);
xnor U15283 (N_15283,N_7912,N_7171);
and U15284 (N_15284,N_6481,N_11142);
nand U15285 (N_15285,N_6734,N_10078);
nand U15286 (N_15286,N_11206,N_10310);
xnor U15287 (N_15287,N_7132,N_6174);
and U15288 (N_15288,N_7401,N_9846);
nand U15289 (N_15289,N_7853,N_6215);
xor U15290 (N_15290,N_7227,N_7780);
and U15291 (N_15291,N_7330,N_8912);
nor U15292 (N_15292,N_10536,N_11771);
and U15293 (N_15293,N_8009,N_11091);
nor U15294 (N_15294,N_6089,N_6955);
and U15295 (N_15295,N_10693,N_8052);
or U15296 (N_15296,N_8931,N_7708);
and U15297 (N_15297,N_7874,N_10797);
and U15298 (N_15298,N_10715,N_6773);
nand U15299 (N_15299,N_9100,N_8671);
nand U15300 (N_15300,N_8169,N_7205);
nor U15301 (N_15301,N_9459,N_6520);
and U15302 (N_15302,N_9153,N_11720);
or U15303 (N_15303,N_9048,N_10544);
xnor U15304 (N_15304,N_10687,N_6406);
nand U15305 (N_15305,N_10828,N_7099);
or U15306 (N_15306,N_11615,N_7170);
nor U15307 (N_15307,N_9110,N_11628);
or U15308 (N_15308,N_9500,N_8818);
nor U15309 (N_15309,N_9579,N_10668);
and U15310 (N_15310,N_6447,N_7036);
nor U15311 (N_15311,N_9357,N_7835);
or U15312 (N_15312,N_9455,N_8447);
nand U15313 (N_15313,N_10597,N_11783);
nor U15314 (N_15314,N_11613,N_7075);
nor U15315 (N_15315,N_10360,N_8382);
and U15316 (N_15316,N_6322,N_11921);
nand U15317 (N_15317,N_7229,N_9438);
or U15318 (N_15318,N_8226,N_8153);
nor U15319 (N_15319,N_8306,N_8831);
xor U15320 (N_15320,N_9431,N_10138);
and U15321 (N_15321,N_11764,N_10120);
or U15322 (N_15322,N_10335,N_8522);
nand U15323 (N_15323,N_9296,N_8214);
or U15324 (N_15324,N_11240,N_8205);
nand U15325 (N_15325,N_7683,N_7452);
or U15326 (N_15326,N_7243,N_7901);
nand U15327 (N_15327,N_10446,N_6519);
or U15328 (N_15328,N_9663,N_6242);
xnor U15329 (N_15329,N_8694,N_8638);
and U15330 (N_15330,N_11275,N_7417);
or U15331 (N_15331,N_11176,N_8545);
and U15332 (N_15332,N_10686,N_7989);
and U15333 (N_15333,N_11132,N_9851);
or U15334 (N_15334,N_9676,N_6067);
nand U15335 (N_15335,N_7002,N_11663);
xnor U15336 (N_15336,N_11408,N_8470);
and U15337 (N_15337,N_7534,N_9460);
or U15338 (N_15338,N_9388,N_11661);
and U15339 (N_15339,N_8518,N_9530);
nand U15340 (N_15340,N_11428,N_6577);
or U15341 (N_15341,N_10816,N_8038);
nand U15342 (N_15342,N_8093,N_8894);
xor U15343 (N_15343,N_6611,N_11673);
nor U15344 (N_15344,N_8011,N_7100);
or U15345 (N_15345,N_7375,N_6862);
nor U15346 (N_15346,N_7544,N_9612);
or U15347 (N_15347,N_6622,N_9156);
and U15348 (N_15348,N_9396,N_10774);
nand U15349 (N_15349,N_10936,N_9264);
nand U15350 (N_15350,N_11177,N_7087);
xnor U15351 (N_15351,N_8345,N_7187);
and U15352 (N_15352,N_10018,N_8216);
xor U15353 (N_15353,N_10227,N_10197);
and U15354 (N_15354,N_8458,N_7331);
or U15355 (N_15355,N_7640,N_10649);
nor U15356 (N_15356,N_7516,N_7882);
and U15357 (N_15357,N_9662,N_9101);
nand U15358 (N_15358,N_7602,N_6587);
nor U15359 (N_15359,N_10395,N_11782);
xnor U15360 (N_15360,N_9175,N_6231);
nand U15361 (N_15361,N_10505,N_8444);
and U15362 (N_15362,N_8388,N_8421);
nor U15363 (N_15363,N_8063,N_6669);
and U15364 (N_15364,N_11527,N_8968);
xnor U15365 (N_15365,N_8711,N_7250);
xnor U15366 (N_15366,N_11697,N_10449);
or U15367 (N_15367,N_6201,N_10835);
or U15368 (N_15368,N_8329,N_9870);
xnor U15369 (N_15369,N_8750,N_9810);
and U15370 (N_15370,N_9559,N_7911);
and U15371 (N_15371,N_9478,N_6055);
nor U15372 (N_15372,N_8698,N_6080);
nor U15373 (N_15373,N_9255,N_9342);
or U15374 (N_15374,N_8737,N_9846);
xnor U15375 (N_15375,N_9606,N_7886);
or U15376 (N_15376,N_9728,N_11311);
nor U15377 (N_15377,N_7841,N_6030);
nor U15378 (N_15378,N_10634,N_10395);
nor U15379 (N_15379,N_11825,N_6444);
or U15380 (N_15380,N_10433,N_7118);
nor U15381 (N_15381,N_6246,N_10454);
nand U15382 (N_15382,N_7573,N_8113);
and U15383 (N_15383,N_7867,N_9800);
nand U15384 (N_15384,N_11340,N_11727);
xor U15385 (N_15385,N_8921,N_10020);
nor U15386 (N_15386,N_10985,N_10870);
and U15387 (N_15387,N_11813,N_9191);
xor U15388 (N_15388,N_7860,N_9964);
xor U15389 (N_15389,N_10136,N_10222);
xor U15390 (N_15390,N_8105,N_11844);
or U15391 (N_15391,N_8547,N_10033);
nand U15392 (N_15392,N_7298,N_7826);
and U15393 (N_15393,N_7555,N_10560);
nand U15394 (N_15394,N_8801,N_9828);
and U15395 (N_15395,N_8673,N_10375);
nand U15396 (N_15396,N_8445,N_6064);
xnor U15397 (N_15397,N_9745,N_6214);
and U15398 (N_15398,N_9036,N_11409);
or U15399 (N_15399,N_9110,N_7144);
or U15400 (N_15400,N_10949,N_7546);
nor U15401 (N_15401,N_8045,N_10215);
nand U15402 (N_15402,N_6353,N_8810);
nor U15403 (N_15403,N_11231,N_9184);
xnor U15404 (N_15404,N_6677,N_6876);
xor U15405 (N_15405,N_6527,N_10831);
and U15406 (N_15406,N_8655,N_7518);
or U15407 (N_15407,N_11376,N_11869);
xor U15408 (N_15408,N_9675,N_6872);
and U15409 (N_15409,N_9259,N_8135);
xnor U15410 (N_15410,N_11884,N_10939);
nor U15411 (N_15411,N_7597,N_11788);
xnor U15412 (N_15412,N_9069,N_8675);
nor U15413 (N_15413,N_6750,N_11149);
xnor U15414 (N_15414,N_8750,N_9179);
xnor U15415 (N_15415,N_9660,N_9613);
nor U15416 (N_15416,N_11544,N_11709);
xnor U15417 (N_15417,N_9463,N_10483);
and U15418 (N_15418,N_8680,N_11317);
nand U15419 (N_15419,N_6793,N_7717);
or U15420 (N_15420,N_7302,N_8978);
nand U15421 (N_15421,N_11710,N_10122);
and U15422 (N_15422,N_6738,N_6304);
xor U15423 (N_15423,N_8414,N_10388);
xor U15424 (N_15424,N_6504,N_10318);
nand U15425 (N_15425,N_10606,N_7962);
and U15426 (N_15426,N_6382,N_8506);
and U15427 (N_15427,N_8130,N_7500);
nand U15428 (N_15428,N_11942,N_6521);
or U15429 (N_15429,N_10260,N_9459);
and U15430 (N_15430,N_6612,N_9965);
and U15431 (N_15431,N_6781,N_10709);
or U15432 (N_15432,N_11208,N_7947);
or U15433 (N_15433,N_8883,N_11817);
and U15434 (N_15434,N_9076,N_11916);
or U15435 (N_15435,N_7398,N_9715);
or U15436 (N_15436,N_6585,N_6922);
nor U15437 (N_15437,N_8951,N_9305);
or U15438 (N_15438,N_8539,N_7628);
nand U15439 (N_15439,N_8923,N_7724);
and U15440 (N_15440,N_6583,N_9333);
xor U15441 (N_15441,N_11278,N_6092);
or U15442 (N_15442,N_9789,N_7044);
nor U15443 (N_15443,N_7354,N_10401);
and U15444 (N_15444,N_7450,N_11037);
and U15445 (N_15445,N_7503,N_11943);
nor U15446 (N_15446,N_9879,N_9019);
or U15447 (N_15447,N_10758,N_8713);
xnor U15448 (N_15448,N_7501,N_9380);
or U15449 (N_15449,N_9524,N_9778);
nor U15450 (N_15450,N_10705,N_6888);
nor U15451 (N_15451,N_11692,N_11061);
nor U15452 (N_15452,N_7228,N_7154);
nor U15453 (N_15453,N_7981,N_11391);
and U15454 (N_15454,N_6451,N_6408);
and U15455 (N_15455,N_6857,N_8602);
nand U15456 (N_15456,N_9556,N_9125);
or U15457 (N_15457,N_7819,N_6894);
and U15458 (N_15458,N_9094,N_9241);
nor U15459 (N_15459,N_11924,N_6447);
xor U15460 (N_15460,N_6924,N_6876);
nor U15461 (N_15461,N_10438,N_8917);
or U15462 (N_15462,N_6807,N_8562);
nor U15463 (N_15463,N_8846,N_10633);
and U15464 (N_15464,N_9998,N_8656);
and U15465 (N_15465,N_6322,N_10391);
nand U15466 (N_15466,N_9251,N_8867);
nand U15467 (N_15467,N_10638,N_8262);
nor U15468 (N_15468,N_7568,N_9658);
nand U15469 (N_15469,N_6251,N_6038);
nor U15470 (N_15470,N_6424,N_6849);
nand U15471 (N_15471,N_11893,N_10168);
nor U15472 (N_15472,N_6542,N_6162);
or U15473 (N_15473,N_10088,N_11188);
xor U15474 (N_15474,N_6009,N_9444);
xor U15475 (N_15475,N_7024,N_6588);
xor U15476 (N_15476,N_10132,N_10654);
nor U15477 (N_15477,N_7387,N_7886);
xnor U15478 (N_15478,N_6441,N_8427);
xor U15479 (N_15479,N_10139,N_10841);
xnor U15480 (N_15480,N_6301,N_9677);
nor U15481 (N_15481,N_11774,N_7981);
nand U15482 (N_15482,N_11859,N_6235);
xnor U15483 (N_15483,N_10028,N_6357);
nand U15484 (N_15484,N_9421,N_8621);
or U15485 (N_15485,N_8537,N_10762);
nor U15486 (N_15486,N_11933,N_10117);
nor U15487 (N_15487,N_6470,N_10437);
and U15488 (N_15488,N_10751,N_6607);
nand U15489 (N_15489,N_8132,N_11839);
xor U15490 (N_15490,N_11075,N_11139);
or U15491 (N_15491,N_7550,N_10157);
nand U15492 (N_15492,N_8181,N_8239);
xnor U15493 (N_15493,N_7980,N_10029);
nor U15494 (N_15494,N_11654,N_7172);
nand U15495 (N_15495,N_8725,N_9555);
and U15496 (N_15496,N_6757,N_6241);
or U15497 (N_15497,N_10287,N_10664);
nand U15498 (N_15498,N_7686,N_6812);
and U15499 (N_15499,N_9588,N_8824);
and U15500 (N_15500,N_11863,N_10548);
nor U15501 (N_15501,N_9638,N_6363);
nand U15502 (N_15502,N_7254,N_7293);
or U15503 (N_15503,N_8198,N_7892);
nand U15504 (N_15504,N_6925,N_6955);
xnor U15505 (N_15505,N_10518,N_6841);
or U15506 (N_15506,N_9044,N_8039);
nor U15507 (N_15507,N_7187,N_8150);
xor U15508 (N_15508,N_11226,N_6344);
and U15509 (N_15509,N_10602,N_10211);
or U15510 (N_15510,N_9605,N_10667);
nand U15511 (N_15511,N_6878,N_11673);
or U15512 (N_15512,N_7145,N_6992);
and U15513 (N_15513,N_8197,N_9814);
and U15514 (N_15514,N_11667,N_10546);
nand U15515 (N_15515,N_10403,N_11233);
xnor U15516 (N_15516,N_11584,N_8039);
or U15517 (N_15517,N_8827,N_8512);
xnor U15518 (N_15518,N_6495,N_10319);
xnor U15519 (N_15519,N_6687,N_10488);
nor U15520 (N_15520,N_10467,N_11540);
or U15521 (N_15521,N_7486,N_7212);
nor U15522 (N_15522,N_7176,N_7347);
and U15523 (N_15523,N_8439,N_6372);
and U15524 (N_15524,N_11760,N_11067);
nor U15525 (N_15525,N_9281,N_6107);
and U15526 (N_15526,N_10089,N_6062);
and U15527 (N_15527,N_6017,N_7705);
or U15528 (N_15528,N_10295,N_11298);
xor U15529 (N_15529,N_11605,N_10445);
nor U15530 (N_15530,N_10066,N_8713);
nor U15531 (N_15531,N_8784,N_9713);
nand U15532 (N_15532,N_7438,N_6829);
nand U15533 (N_15533,N_10942,N_10450);
or U15534 (N_15534,N_6105,N_10985);
nand U15535 (N_15535,N_10632,N_11290);
nor U15536 (N_15536,N_9361,N_8828);
or U15537 (N_15537,N_6957,N_11625);
nor U15538 (N_15538,N_7376,N_9102);
nand U15539 (N_15539,N_9320,N_9577);
xor U15540 (N_15540,N_6505,N_6773);
or U15541 (N_15541,N_6273,N_11402);
and U15542 (N_15542,N_9178,N_8023);
nor U15543 (N_15543,N_6073,N_6046);
xor U15544 (N_15544,N_8029,N_11790);
or U15545 (N_15545,N_9029,N_11932);
nor U15546 (N_15546,N_7026,N_8339);
or U15547 (N_15547,N_8898,N_10161);
or U15548 (N_15548,N_8019,N_9385);
xnor U15549 (N_15549,N_8559,N_6206);
and U15550 (N_15550,N_9036,N_9207);
nor U15551 (N_15551,N_10679,N_11319);
and U15552 (N_15552,N_8922,N_10262);
or U15553 (N_15553,N_11090,N_7173);
nor U15554 (N_15554,N_11586,N_10671);
nor U15555 (N_15555,N_9718,N_9404);
nor U15556 (N_15556,N_9077,N_6889);
xnor U15557 (N_15557,N_7626,N_10715);
or U15558 (N_15558,N_8064,N_10923);
xnor U15559 (N_15559,N_7329,N_9451);
nand U15560 (N_15560,N_9845,N_11152);
or U15561 (N_15561,N_6116,N_11216);
nor U15562 (N_15562,N_6581,N_8207);
nor U15563 (N_15563,N_10916,N_9951);
nor U15564 (N_15564,N_7878,N_10030);
nand U15565 (N_15565,N_7238,N_10890);
xor U15566 (N_15566,N_8311,N_6882);
nand U15567 (N_15567,N_7075,N_11843);
nor U15568 (N_15568,N_6029,N_9683);
nand U15569 (N_15569,N_11641,N_7540);
and U15570 (N_15570,N_11382,N_8071);
nand U15571 (N_15571,N_9604,N_11606);
xnor U15572 (N_15572,N_6402,N_11869);
nor U15573 (N_15573,N_9739,N_11072);
and U15574 (N_15574,N_7195,N_11783);
nand U15575 (N_15575,N_7823,N_8277);
xor U15576 (N_15576,N_11229,N_6293);
nor U15577 (N_15577,N_7151,N_8827);
nor U15578 (N_15578,N_8743,N_7518);
nor U15579 (N_15579,N_6856,N_10723);
and U15580 (N_15580,N_8168,N_10269);
xor U15581 (N_15581,N_6360,N_10190);
and U15582 (N_15582,N_11065,N_11200);
and U15583 (N_15583,N_8405,N_9295);
nand U15584 (N_15584,N_6498,N_6245);
and U15585 (N_15585,N_6780,N_11208);
or U15586 (N_15586,N_7712,N_10181);
or U15587 (N_15587,N_6139,N_7417);
and U15588 (N_15588,N_6249,N_6878);
nor U15589 (N_15589,N_9353,N_9339);
xnor U15590 (N_15590,N_7221,N_8649);
nor U15591 (N_15591,N_7971,N_11469);
xnor U15592 (N_15592,N_9193,N_6951);
nand U15593 (N_15593,N_11221,N_6468);
and U15594 (N_15594,N_9945,N_10189);
nand U15595 (N_15595,N_11410,N_10141);
nor U15596 (N_15596,N_6962,N_10405);
xnor U15597 (N_15597,N_7165,N_11106);
or U15598 (N_15598,N_9907,N_7200);
xnor U15599 (N_15599,N_10754,N_9997);
xor U15600 (N_15600,N_11574,N_11307);
and U15601 (N_15601,N_7777,N_11700);
xor U15602 (N_15602,N_11791,N_6145);
nor U15603 (N_15603,N_7281,N_7717);
and U15604 (N_15604,N_7216,N_10003);
nor U15605 (N_15605,N_7004,N_7403);
xnor U15606 (N_15606,N_8855,N_9655);
or U15607 (N_15607,N_7707,N_8053);
nand U15608 (N_15608,N_6140,N_6876);
or U15609 (N_15609,N_11514,N_9738);
or U15610 (N_15610,N_7983,N_6940);
nand U15611 (N_15611,N_7918,N_9423);
and U15612 (N_15612,N_7965,N_9114);
or U15613 (N_15613,N_10337,N_7348);
and U15614 (N_15614,N_11160,N_9295);
xnor U15615 (N_15615,N_7369,N_9883);
nand U15616 (N_15616,N_11472,N_10593);
nand U15617 (N_15617,N_8550,N_7613);
and U15618 (N_15618,N_11791,N_10829);
and U15619 (N_15619,N_8765,N_11542);
and U15620 (N_15620,N_9709,N_6304);
or U15621 (N_15621,N_8977,N_8535);
nor U15622 (N_15622,N_11537,N_6667);
nor U15623 (N_15623,N_9937,N_9838);
nor U15624 (N_15624,N_9500,N_6115);
nand U15625 (N_15625,N_11569,N_9929);
and U15626 (N_15626,N_6592,N_7269);
xor U15627 (N_15627,N_8483,N_8406);
and U15628 (N_15628,N_6359,N_8911);
and U15629 (N_15629,N_11813,N_6243);
nand U15630 (N_15630,N_9673,N_6531);
xnor U15631 (N_15631,N_9275,N_8986);
and U15632 (N_15632,N_7387,N_11816);
or U15633 (N_15633,N_10665,N_10142);
nor U15634 (N_15634,N_7949,N_6187);
and U15635 (N_15635,N_9642,N_7072);
nand U15636 (N_15636,N_6548,N_8243);
nor U15637 (N_15637,N_9987,N_11320);
or U15638 (N_15638,N_7343,N_7757);
nor U15639 (N_15639,N_8389,N_7955);
nand U15640 (N_15640,N_10116,N_9868);
and U15641 (N_15641,N_9702,N_10640);
nor U15642 (N_15642,N_11238,N_10726);
and U15643 (N_15643,N_7942,N_10766);
or U15644 (N_15644,N_6345,N_7926);
nand U15645 (N_15645,N_10805,N_10887);
nand U15646 (N_15646,N_7411,N_7021);
and U15647 (N_15647,N_7202,N_10801);
and U15648 (N_15648,N_7739,N_9728);
nand U15649 (N_15649,N_7385,N_7163);
nor U15650 (N_15650,N_9421,N_8652);
or U15651 (N_15651,N_8064,N_7327);
xor U15652 (N_15652,N_7327,N_10185);
xnor U15653 (N_15653,N_10817,N_10618);
or U15654 (N_15654,N_7745,N_7049);
xor U15655 (N_15655,N_10249,N_8321);
and U15656 (N_15656,N_7585,N_11799);
or U15657 (N_15657,N_6205,N_11715);
nand U15658 (N_15658,N_7421,N_11030);
nand U15659 (N_15659,N_7197,N_7661);
nand U15660 (N_15660,N_7104,N_8443);
or U15661 (N_15661,N_7603,N_6057);
and U15662 (N_15662,N_6751,N_6642);
and U15663 (N_15663,N_7122,N_7349);
xnor U15664 (N_15664,N_8060,N_11995);
xnor U15665 (N_15665,N_7556,N_7945);
nor U15666 (N_15666,N_10832,N_8414);
and U15667 (N_15667,N_10714,N_11672);
xor U15668 (N_15668,N_9563,N_10716);
or U15669 (N_15669,N_9297,N_8390);
nand U15670 (N_15670,N_10395,N_10764);
and U15671 (N_15671,N_10176,N_6986);
nand U15672 (N_15672,N_8412,N_8896);
xor U15673 (N_15673,N_6831,N_9945);
nand U15674 (N_15674,N_9660,N_7690);
or U15675 (N_15675,N_7348,N_7651);
xor U15676 (N_15676,N_10767,N_8537);
xor U15677 (N_15677,N_11227,N_10232);
nand U15678 (N_15678,N_8220,N_11377);
nand U15679 (N_15679,N_11426,N_11192);
and U15680 (N_15680,N_10552,N_8116);
nor U15681 (N_15681,N_6994,N_11737);
and U15682 (N_15682,N_10897,N_9048);
nand U15683 (N_15683,N_9742,N_7939);
xor U15684 (N_15684,N_8422,N_11547);
nand U15685 (N_15685,N_7306,N_9299);
or U15686 (N_15686,N_8601,N_6296);
and U15687 (N_15687,N_11713,N_8052);
and U15688 (N_15688,N_8066,N_11103);
nand U15689 (N_15689,N_11592,N_8129);
nand U15690 (N_15690,N_10143,N_6537);
or U15691 (N_15691,N_11322,N_11455);
nand U15692 (N_15692,N_10826,N_6974);
nand U15693 (N_15693,N_10907,N_10797);
or U15694 (N_15694,N_11146,N_6387);
or U15695 (N_15695,N_11779,N_9457);
nand U15696 (N_15696,N_9873,N_11642);
and U15697 (N_15697,N_9037,N_11652);
and U15698 (N_15698,N_11239,N_6877);
xor U15699 (N_15699,N_6685,N_10218);
or U15700 (N_15700,N_9918,N_9603);
and U15701 (N_15701,N_8447,N_6243);
nand U15702 (N_15702,N_7641,N_7962);
or U15703 (N_15703,N_8142,N_7030);
xnor U15704 (N_15704,N_9785,N_10224);
xnor U15705 (N_15705,N_6200,N_7519);
nor U15706 (N_15706,N_9589,N_6153);
nor U15707 (N_15707,N_7981,N_11434);
or U15708 (N_15708,N_8813,N_7906);
nand U15709 (N_15709,N_11785,N_10466);
or U15710 (N_15710,N_6222,N_11831);
nand U15711 (N_15711,N_6782,N_10016);
or U15712 (N_15712,N_9718,N_9489);
or U15713 (N_15713,N_11502,N_6231);
or U15714 (N_15714,N_8163,N_7797);
and U15715 (N_15715,N_9531,N_8203);
and U15716 (N_15716,N_9754,N_6551);
and U15717 (N_15717,N_8921,N_6269);
nand U15718 (N_15718,N_9100,N_6486);
or U15719 (N_15719,N_11951,N_7573);
nand U15720 (N_15720,N_7694,N_10085);
or U15721 (N_15721,N_11139,N_8813);
nand U15722 (N_15722,N_9239,N_8180);
or U15723 (N_15723,N_9242,N_6945);
nor U15724 (N_15724,N_11244,N_10533);
nor U15725 (N_15725,N_7022,N_8521);
nor U15726 (N_15726,N_6675,N_8122);
nand U15727 (N_15727,N_9931,N_6377);
or U15728 (N_15728,N_6648,N_7327);
and U15729 (N_15729,N_7808,N_10314);
xnor U15730 (N_15730,N_9891,N_9467);
xor U15731 (N_15731,N_11305,N_10807);
and U15732 (N_15732,N_7520,N_8350);
or U15733 (N_15733,N_10157,N_8585);
xor U15734 (N_15734,N_11289,N_8167);
xnor U15735 (N_15735,N_10228,N_11056);
and U15736 (N_15736,N_7864,N_10993);
nand U15737 (N_15737,N_9164,N_9878);
or U15738 (N_15738,N_11243,N_7694);
or U15739 (N_15739,N_8057,N_11846);
xor U15740 (N_15740,N_11397,N_7302);
and U15741 (N_15741,N_11379,N_8208);
or U15742 (N_15742,N_7720,N_6141);
nand U15743 (N_15743,N_9429,N_6821);
nor U15744 (N_15744,N_6808,N_7298);
nor U15745 (N_15745,N_9425,N_7298);
nand U15746 (N_15746,N_11794,N_9089);
xnor U15747 (N_15747,N_11744,N_6475);
nor U15748 (N_15748,N_8265,N_7662);
and U15749 (N_15749,N_7141,N_11503);
nand U15750 (N_15750,N_11926,N_7655);
or U15751 (N_15751,N_7389,N_6800);
and U15752 (N_15752,N_9740,N_11940);
nor U15753 (N_15753,N_6809,N_10734);
and U15754 (N_15754,N_8000,N_6447);
or U15755 (N_15755,N_6209,N_8321);
nor U15756 (N_15756,N_9810,N_9375);
xnor U15757 (N_15757,N_7544,N_6363);
and U15758 (N_15758,N_9157,N_11281);
or U15759 (N_15759,N_9863,N_10936);
or U15760 (N_15760,N_10700,N_10509);
and U15761 (N_15761,N_11921,N_9259);
nor U15762 (N_15762,N_10290,N_11777);
and U15763 (N_15763,N_11589,N_7435);
nor U15764 (N_15764,N_9487,N_6361);
nor U15765 (N_15765,N_7434,N_11888);
xnor U15766 (N_15766,N_8562,N_11847);
nor U15767 (N_15767,N_11014,N_6774);
or U15768 (N_15768,N_9477,N_6752);
xor U15769 (N_15769,N_9666,N_11680);
nand U15770 (N_15770,N_9721,N_6638);
or U15771 (N_15771,N_7604,N_6065);
xor U15772 (N_15772,N_11215,N_8683);
nor U15773 (N_15773,N_9574,N_11218);
nor U15774 (N_15774,N_6980,N_8538);
nor U15775 (N_15775,N_10349,N_10260);
or U15776 (N_15776,N_11929,N_6229);
nor U15777 (N_15777,N_11159,N_8710);
xnor U15778 (N_15778,N_8902,N_11256);
nand U15779 (N_15779,N_11627,N_8057);
nand U15780 (N_15780,N_6286,N_8145);
and U15781 (N_15781,N_8356,N_11230);
or U15782 (N_15782,N_6023,N_10209);
nand U15783 (N_15783,N_6300,N_7584);
or U15784 (N_15784,N_6340,N_6785);
nand U15785 (N_15785,N_6198,N_10822);
and U15786 (N_15786,N_10966,N_6750);
nand U15787 (N_15787,N_8108,N_6891);
xor U15788 (N_15788,N_11673,N_10612);
or U15789 (N_15789,N_9518,N_11868);
nor U15790 (N_15790,N_6746,N_10797);
nand U15791 (N_15791,N_7915,N_6267);
nor U15792 (N_15792,N_7182,N_8229);
nand U15793 (N_15793,N_8616,N_8193);
and U15794 (N_15794,N_8088,N_10577);
or U15795 (N_15795,N_10733,N_9331);
and U15796 (N_15796,N_9602,N_11838);
nor U15797 (N_15797,N_8741,N_7314);
nor U15798 (N_15798,N_10210,N_8881);
or U15799 (N_15799,N_10936,N_6030);
xnor U15800 (N_15800,N_7470,N_9164);
nand U15801 (N_15801,N_7310,N_11799);
or U15802 (N_15802,N_6308,N_6073);
nand U15803 (N_15803,N_8828,N_10896);
nor U15804 (N_15804,N_6595,N_6958);
and U15805 (N_15805,N_9114,N_9382);
nand U15806 (N_15806,N_10889,N_11532);
nor U15807 (N_15807,N_10442,N_7866);
and U15808 (N_15808,N_7736,N_7655);
nor U15809 (N_15809,N_6705,N_11114);
and U15810 (N_15810,N_9327,N_8915);
nand U15811 (N_15811,N_8471,N_7375);
nor U15812 (N_15812,N_7253,N_7164);
xnor U15813 (N_15813,N_11326,N_6965);
xor U15814 (N_15814,N_7057,N_8012);
nor U15815 (N_15815,N_9952,N_7828);
nand U15816 (N_15816,N_11169,N_8219);
nand U15817 (N_15817,N_11827,N_9911);
nand U15818 (N_15818,N_9730,N_8013);
and U15819 (N_15819,N_11680,N_6177);
and U15820 (N_15820,N_8970,N_9971);
and U15821 (N_15821,N_7676,N_9127);
and U15822 (N_15822,N_8307,N_10286);
nand U15823 (N_15823,N_8739,N_6434);
nor U15824 (N_15824,N_6557,N_10990);
nor U15825 (N_15825,N_7155,N_9454);
and U15826 (N_15826,N_6410,N_10077);
xnor U15827 (N_15827,N_7774,N_7422);
and U15828 (N_15828,N_8614,N_11975);
or U15829 (N_15829,N_6033,N_8684);
nor U15830 (N_15830,N_9290,N_6515);
or U15831 (N_15831,N_9257,N_8630);
and U15832 (N_15832,N_11804,N_6442);
and U15833 (N_15833,N_7936,N_10163);
xor U15834 (N_15834,N_9860,N_8988);
nand U15835 (N_15835,N_6334,N_8874);
nand U15836 (N_15836,N_8927,N_10520);
nand U15837 (N_15837,N_10754,N_9202);
or U15838 (N_15838,N_9554,N_7819);
or U15839 (N_15839,N_11312,N_8354);
or U15840 (N_15840,N_7094,N_9620);
and U15841 (N_15841,N_7473,N_11453);
and U15842 (N_15842,N_11143,N_8996);
nor U15843 (N_15843,N_8678,N_10953);
and U15844 (N_15844,N_11486,N_6237);
or U15845 (N_15845,N_8928,N_7270);
nand U15846 (N_15846,N_11955,N_11047);
or U15847 (N_15847,N_11676,N_7518);
nor U15848 (N_15848,N_9916,N_10217);
and U15849 (N_15849,N_6247,N_6294);
or U15850 (N_15850,N_6979,N_8187);
xor U15851 (N_15851,N_6604,N_6390);
nor U15852 (N_15852,N_8076,N_10833);
and U15853 (N_15853,N_11080,N_10003);
xor U15854 (N_15854,N_9912,N_7544);
nor U15855 (N_15855,N_10131,N_9004);
nand U15856 (N_15856,N_6098,N_7104);
xor U15857 (N_15857,N_11916,N_9881);
and U15858 (N_15858,N_10099,N_7983);
nor U15859 (N_15859,N_10511,N_8444);
nand U15860 (N_15860,N_7728,N_8228);
nor U15861 (N_15861,N_7146,N_7865);
nand U15862 (N_15862,N_10728,N_8670);
nand U15863 (N_15863,N_10974,N_9535);
and U15864 (N_15864,N_11991,N_9645);
and U15865 (N_15865,N_11422,N_10826);
and U15866 (N_15866,N_8786,N_9353);
or U15867 (N_15867,N_8357,N_9397);
nor U15868 (N_15868,N_8560,N_11445);
nand U15869 (N_15869,N_10815,N_9328);
or U15870 (N_15870,N_7937,N_10927);
nor U15871 (N_15871,N_7866,N_10013);
nor U15872 (N_15872,N_7702,N_8930);
nor U15873 (N_15873,N_6204,N_8910);
nand U15874 (N_15874,N_7689,N_7308);
and U15875 (N_15875,N_7891,N_11927);
nand U15876 (N_15876,N_7962,N_10476);
or U15877 (N_15877,N_11891,N_6657);
and U15878 (N_15878,N_9547,N_6445);
nand U15879 (N_15879,N_10362,N_6892);
xnor U15880 (N_15880,N_10221,N_11661);
and U15881 (N_15881,N_11451,N_8320);
nand U15882 (N_15882,N_8930,N_10712);
nand U15883 (N_15883,N_9219,N_8241);
and U15884 (N_15884,N_10666,N_6186);
nand U15885 (N_15885,N_9309,N_6536);
nand U15886 (N_15886,N_8395,N_10398);
nor U15887 (N_15887,N_11234,N_10943);
nor U15888 (N_15888,N_10729,N_10889);
or U15889 (N_15889,N_6845,N_6698);
or U15890 (N_15890,N_7855,N_8477);
nor U15891 (N_15891,N_11317,N_10444);
nand U15892 (N_15892,N_10046,N_8815);
and U15893 (N_15893,N_8281,N_11626);
nand U15894 (N_15894,N_7400,N_10267);
nand U15895 (N_15895,N_11980,N_7425);
and U15896 (N_15896,N_9918,N_9988);
nor U15897 (N_15897,N_9019,N_11118);
and U15898 (N_15898,N_6416,N_9640);
xnor U15899 (N_15899,N_8108,N_8992);
nor U15900 (N_15900,N_7996,N_9931);
or U15901 (N_15901,N_11815,N_7668);
nand U15902 (N_15902,N_11662,N_8962);
and U15903 (N_15903,N_6908,N_9112);
and U15904 (N_15904,N_6358,N_9845);
and U15905 (N_15905,N_6600,N_10721);
or U15906 (N_15906,N_9161,N_9374);
or U15907 (N_15907,N_9629,N_9391);
and U15908 (N_15908,N_7076,N_8395);
and U15909 (N_15909,N_9107,N_8623);
or U15910 (N_15910,N_8793,N_6193);
and U15911 (N_15911,N_8969,N_11980);
or U15912 (N_15912,N_6029,N_7681);
nand U15913 (N_15913,N_11932,N_8669);
nand U15914 (N_15914,N_9649,N_6796);
xor U15915 (N_15915,N_11192,N_10791);
or U15916 (N_15916,N_6043,N_11076);
and U15917 (N_15917,N_8136,N_6659);
nand U15918 (N_15918,N_7900,N_10391);
nor U15919 (N_15919,N_8428,N_8292);
or U15920 (N_15920,N_11501,N_9310);
nor U15921 (N_15921,N_7510,N_7414);
nor U15922 (N_15922,N_6187,N_7054);
and U15923 (N_15923,N_11949,N_11388);
or U15924 (N_15924,N_10836,N_8570);
xor U15925 (N_15925,N_9056,N_6955);
and U15926 (N_15926,N_9554,N_9971);
or U15927 (N_15927,N_7921,N_9294);
and U15928 (N_15928,N_8473,N_8045);
nand U15929 (N_15929,N_9426,N_7725);
or U15930 (N_15930,N_8348,N_6540);
and U15931 (N_15931,N_8698,N_6950);
or U15932 (N_15932,N_7428,N_6009);
and U15933 (N_15933,N_11804,N_10079);
or U15934 (N_15934,N_10821,N_10357);
xnor U15935 (N_15935,N_11489,N_7008);
or U15936 (N_15936,N_10614,N_10359);
or U15937 (N_15937,N_7992,N_6416);
or U15938 (N_15938,N_7863,N_7861);
xor U15939 (N_15939,N_11141,N_6663);
nor U15940 (N_15940,N_7648,N_7369);
xor U15941 (N_15941,N_9875,N_7140);
nor U15942 (N_15942,N_7591,N_11872);
nor U15943 (N_15943,N_6258,N_11179);
or U15944 (N_15944,N_6814,N_9431);
and U15945 (N_15945,N_11641,N_7594);
nor U15946 (N_15946,N_7715,N_9399);
nor U15947 (N_15947,N_8425,N_6718);
and U15948 (N_15948,N_10044,N_9126);
xnor U15949 (N_15949,N_10609,N_10592);
xor U15950 (N_15950,N_8477,N_9860);
nor U15951 (N_15951,N_10631,N_6632);
xor U15952 (N_15952,N_8928,N_7428);
nand U15953 (N_15953,N_6325,N_7797);
nand U15954 (N_15954,N_11509,N_10641);
and U15955 (N_15955,N_9803,N_6139);
and U15956 (N_15956,N_9582,N_7367);
nor U15957 (N_15957,N_10031,N_7002);
xor U15958 (N_15958,N_8516,N_6942);
nor U15959 (N_15959,N_6889,N_6312);
and U15960 (N_15960,N_6981,N_6174);
nand U15961 (N_15961,N_7032,N_11712);
nor U15962 (N_15962,N_11135,N_9431);
nor U15963 (N_15963,N_11192,N_11270);
nor U15964 (N_15964,N_11877,N_9938);
nor U15965 (N_15965,N_9484,N_10010);
xor U15966 (N_15966,N_8703,N_6771);
nor U15967 (N_15967,N_9506,N_6638);
nor U15968 (N_15968,N_10956,N_6123);
or U15969 (N_15969,N_7757,N_10855);
nor U15970 (N_15970,N_10336,N_9271);
nor U15971 (N_15971,N_10545,N_9492);
nand U15972 (N_15972,N_6262,N_10619);
nor U15973 (N_15973,N_11786,N_11198);
or U15974 (N_15974,N_6600,N_7176);
or U15975 (N_15975,N_9114,N_8789);
xor U15976 (N_15976,N_6718,N_11651);
nand U15977 (N_15977,N_11346,N_9843);
nor U15978 (N_15978,N_10833,N_7486);
and U15979 (N_15979,N_10545,N_10709);
nor U15980 (N_15980,N_11207,N_11721);
nor U15981 (N_15981,N_10400,N_8848);
and U15982 (N_15982,N_7089,N_10362);
and U15983 (N_15983,N_7472,N_11982);
or U15984 (N_15984,N_8185,N_8908);
xor U15985 (N_15985,N_7769,N_10938);
and U15986 (N_15986,N_11198,N_11610);
nand U15987 (N_15987,N_11890,N_6514);
nand U15988 (N_15988,N_10681,N_10814);
xnor U15989 (N_15989,N_11625,N_9587);
and U15990 (N_15990,N_9479,N_7918);
nor U15991 (N_15991,N_9517,N_9296);
nand U15992 (N_15992,N_6246,N_9341);
nand U15993 (N_15993,N_6023,N_9067);
and U15994 (N_15994,N_8900,N_8578);
or U15995 (N_15995,N_8291,N_8714);
nand U15996 (N_15996,N_11755,N_7995);
xnor U15997 (N_15997,N_10787,N_8611);
and U15998 (N_15998,N_8535,N_7761);
and U15999 (N_15999,N_6516,N_11825);
nand U16000 (N_16000,N_9438,N_11697);
and U16001 (N_16001,N_11120,N_7092);
nand U16002 (N_16002,N_7456,N_9551);
nor U16003 (N_16003,N_6992,N_11404);
and U16004 (N_16004,N_9036,N_11471);
and U16005 (N_16005,N_7878,N_10514);
or U16006 (N_16006,N_8636,N_6351);
xor U16007 (N_16007,N_7620,N_11465);
nand U16008 (N_16008,N_9207,N_10204);
and U16009 (N_16009,N_9273,N_10891);
nand U16010 (N_16010,N_11620,N_10132);
and U16011 (N_16011,N_8690,N_6329);
xnor U16012 (N_16012,N_11624,N_10909);
and U16013 (N_16013,N_9230,N_8089);
and U16014 (N_16014,N_6383,N_10140);
and U16015 (N_16015,N_10587,N_6737);
or U16016 (N_16016,N_8394,N_10481);
or U16017 (N_16017,N_11135,N_8794);
nand U16018 (N_16018,N_11173,N_8988);
nand U16019 (N_16019,N_8862,N_9758);
and U16020 (N_16020,N_7219,N_9103);
xor U16021 (N_16021,N_11257,N_11881);
or U16022 (N_16022,N_6847,N_11914);
or U16023 (N_16023,N_8577,N_6066);
nand U16024 (N_16024,N_11788,N_9915);
xor U16025 (N_16025,N_7392,N_10407);
nand U16026 (N_16026,N_11402,N_7890);
and U16027 (N_16027,N_8321,N_6944);
and U16028 (N_16028,N_8493,N_6823);
nor U16029 (N_16029,N_8300,N_9910);
or U16030 (N_16030,N_7335,N_6065);
nand U16031 (N_16031,N_9943,N_7114);
xor U16032 (N_16032,N_9290,N_7509);
xor U16033 (N_16033,N_9815,N_6201);
xor U16034 (N_16034,N_11217,N_10923);
xnor U16035 (N_16035,N_11776,N_7126);
nand U16036 (N_16036,N_6120,N_8470);
nor U16037 (N_16037,N_11644,N_9671);
or U16038 (N_16038,N_10254,N_9541);
nor U16039 (N_16039,N_11402,N_8887);
nand U16040 (N_16040,N_11614,N_10725);
xnor U16041 (N_16041,N_9016,N_9386);
or U16042 (N_16042,N_10772,N_7963);
or U16043 (N_16043,N_6689,N_7962);
and U16044 (N_16044,N_11676,N_8934);
nor U16045 (N_16045,N_8219,N_11364);
xor U16046 (N_16046,N_9070,N_10938);
nor U16047 (N_16047,N_8664,N_9132);
or U16048 (N_16048,N_9462,N_10420);
xor U16049 (N_16049,N_7771,N_8238);
nand U16050 (N_16050,N_7923,N_8800);
or U16051 (N_16051,N_6595,N_8318);
and U16052 (N_16052,N_7972,N_7960);
xor U16053 (N_16053,N_10647,N_7529);
nand U16054 (N_16054,N_8227,N_8050);
and U16055 (N_16055,N_7852,N_9119);
or U16056 (N_16056,N_10454,N_6125);
and U16057 (N_16057,N_10654,N_8089);
and U16058 (N_16058,N_8973,N_10811);
nor U16059 (N_16059,N_6027,N_7601);
xor U16060 (N_16060,N_11378,N_11024);
nor U16061 (N_16061,N_10981,N_6409);
nand U16062 (N_16062,N_11792,N_11537);
nor U16063 (N_16063,N_6354,N_10876);
nor U16064 (N_16064,N_8262,N_8025);
xor U16065 (N_16065,N_10338,N_10792);
nor U16066 (N_16066,N_11518,N_10855);
and U16067 (N_16067,N_8346,N_10465);
nand U16068 (N_16068,N_10486,N_8039);
xnor U16069 (N_16069,N_7635,N_9608);
nor U16070 (N_16070,N_11909,N_8126);
nand U16071 (N_16071,N_7761,N_7438);
or U16072 (N_16072,N_7550,N_7432);
nand U16073 (N_16073,N_11312,N_10865);
xor U16074 (N_16074,N_11853,N_7856);
or U16075 (N_16075,N_7612,N_8623);
nor U16076 (N_16076,N_7225,N_8204);
xor U16077 (N_16077,N_7790,N_11217);
nand U16078 (N_16078,N_9679,N_10047);
nand U16079 (N_16079,N_7879,N_7528);
and U16080 (N_16080,N_8041,N_8033);
nor U16081 (N_16081,N_8114,N_8433);
or U16082 (N_16082,N_11614,N_9035);
nand U16083 (N_16083,N_9074,N_6635);
or U16084 (N_16084,N_9294,N_10931);
nand U16085 (N_16085,N_6347,N_6105);
nand U16086 (N_16086,N_7103,N_6893);
nor U16087 (N_16087,N_6528,N_6659);
nor U16088 (N_16088,N_8857,N_6142);
xnor U16089 (N_16089,N_10770,N_9696);
nor U16090 (N_16090,N_10651,N_11248);
nor U16091 (N_16091,N_6258,N_8057);
and U16092 (N_16092,N_6550,N_7312);
or U16093 (N_16093,N_11158,N_9682);
nand U16094 (N_16094,N_6614,N_10789);
and U16095 (N_16095,N_11630,N_8504);
xnor U16096 (N_16096,N_10355,N_10771);
xor U16097 (N_16097,N_7313,N_8113);
nand U16098 (N_16098,N_6397,N_9276);
nand U16099 (N_16099,N_6945,N_9608);
xnor U16100 (N_16100,N_10819,N_6215);
nor U16101 (N_16101,N_7444,N_10807);
nand U16102 (N_16102,N_8851,N_10307);
nor U16103 (N_16103,N_11075,N_11123);
nor U16104 (N_16104,N_9020,N_7676);
nor U16105 (N_16105,N_8641,N_6199);
nand U16106 (N_16106,N_9234,N_6463);
nor U16107 (N_16107,N_10135,N_11120);
nand U16108 (N_16108,N_8647,N_6011);
and U16109 (N_16109,N_7226,N_8570);
or U16110 (N_16110,N_7463,N_8558);
xor U16111 (N_16111,N_10600,N_11737);
and U16112 (N_16112,N_8942,N_8059);
and U16113 (N_16113,N_8420,N_9160);
xor U16114 (N_16114,N_10642,N_9240);
or U16115 (N_16115,N_9419,N_9884);
and U16116 (N_16116,N_10168,N_7314);
and U16117 (N_16117,N_11569,N_11694);
nor U16118 (N_16118,N_9329,N_10043);
and U16119 (N_16119,N_11269,N_8664);
xnor U16120 (N_16120,N_6590,N_10145);
nand U16121 (N_16121,N_7541,N_8031);
xor U16122 (N_16122,N_11427,N_11819);
nor U16123 (N_16123,N_6542,N_6675);
xnor U16124 (N_16124,N_10896,N_11293);
nor U16125 (N_16125,N_7774,N_8605);
and U16126 (N_16126,N_7802,N_6928);
nor U16127 (N_16127,N_10303,N_8680);
or U16128 (N_16128,N_11074,N_9204);
or U16129 (N_16129,N_7851,N_11277);
nand U16130 (N_16130,N_7847,N_8676);
and U16131 (N_16131,N_10889,N_9539);
and U16132 (N_16132,N_9405,N_10108);
nand U16133 (N_16133,N_6081,N_9973);
xor U16134 (N_16134,N_6281,N_6020);
or U16135 (N_16135,N_11160,N_11516);
nor U16136 (N_16136,N_6262,N_6508);
xnor U16137 (N_16137,N_10949,N_11284);
xor U16138 (N_16138,N_7746,N_9453);
xor U16139 (N_16139,N_7105,N_7359);
nand U16140 (N_16140,N_7988,N_9641);
nand U16141 (N_16141,N_9713,N_8742);
nor U16142 (N_16142,N_7160,N_10353);
nor U16143 (N_16143,N_8934,N_11055);
and U16144 (N_16144,N_7286,N_9519);
nor U16145 (N_16145,N_8471,N_11205);
and U16146 (N_16146,N_10627,N_8693);
nand U16147 (N_16147,N_6642,N_10456);
nor U16148 (N_16148,N_6409,N_9910);
nand U16149 (N_16149,N_6080,N_11042);
and U16150 (N_16150,N_9955,N_10801);
nand U16151 (N_16151,N_6655,N_10883);
or U16152 (N_16152,N_11075,N_7453);
nor U16153 (N_16153,N_10575,N_9212);
nand U16154 (N_16154,N_6797,N_7196);
nor U16155 (N_16155,N_11371,N_7860);
nor U16156 (N_16156,N_10748,N_7249);
and U16157 (N_16157,N_9316,N_9065);
or U16158 (N_16158,N_10824,N_8319);
or U16159 (N_16159,N_11746,N_10453);
or U16160 (N_16160,N_6088,N_10433);
or U16161 (N_16161,N_10015,N_6628);
or U16162 (N_16162,N_8572,N_6396);
xor U16163 (N_16163,N_11821,N_11651);
or U16164 (N_16164,N_7872,N_10141);
nand U16165 (N_16165,N_7657,N_10483);
xor U16166 (N_16166,N_10399,N_7034);
nor U16167 (N_16167,N_8481,N_11714);
nor U16168 (N_16168,N_11655,N_6567);
or U16169 (N_16169,N_10649,N_9251);
and U16170 (N_16170,N_10066,N_6423);
nand U16171 (N_16171,N_9750,N_9389);
and U16172 (N_16172,N_6569,N_10666);
or U16173 (N_16173,N_8755,N_7956);
and U16174 (N_16174,N_10584,N_7178);
and U16175 (N_16175,N_11723,N_7584);
xor U16176 (N_16176,N_7470,N_7361);
or U16177 (N_16177,N_6198,N_7831);
or U16178 (N_16178,N_6500,N_6663);
or U16179 (N_16179,N_11466,N_6520);
and U16180 (N_16180,N_8054,N_6355);
and U16181 (N_16181,N_6625,N_6350);
nor U16182 (N_16182,N_7871,N_7493);
or U16183 (N_16183,N_11151,N_7840);
nand U16184 (N_16184,N_6792,N_9335);
nand U16185 (N_16185,N_7793,N_7801);
nand U16186 (N_16186,N_8833,N_9065);
xnor U16187 (N_16187,N_10872,N_9393);
or U16188 (N_16188,N_11026,N_9409);
xnor U16189 (N_16189,N_8657,N_11563);
and U16190 (N_16190,N_6602,N_9597);
xor U16191 (N_16191,N_9036,N_9441);
nor U16192 (N_16192,N_11444,N_7298);
or U16193 (N_16193,N_10307,N_8655);
xor U16194 (N_16194,N_11573,N_8504);
or U16195 (N_16195,N_11195,N_9207);
xnor U16196 (N_16196,N_10594,N_9145);
and U16197 (N_16197,N_8334,N_10954);
nor U16198 (N_16198,N_7681,N_10908);
and U16199 (N_16199,N_9915,N_9743);
xor U16200 (N_16200,N_11762,N_9902);
xor U16201 (N_16201,N_11859,N_6523);
nand U16202 (N_16202,N_10842,N_11280);
nand U16203 (N_16203,N_7959,N_9059);
or U16204 (N_16204,N_11714,N_7565);
or U16205 (N_16205,N_7501,N_10884);
and U16206 (N_16206,N_8279,N_7171);
nand U16207 (N_16207,N_6511,N_10876);
xor U16208 (N_16208,N_6357,N_8994);
nand U16209 (N_16209,N_6748,N_7824);
xor U16210 (N_16210,N_11119,N_9764);
xnor U16211 (N_16211,N_7724,N_7363);
nor U16212 (N_16212,N_8378,N_10150);
nand U16213 (N_16213,N_6594,N_7007);
xnor U16214 (N_16214,N_9406,N_9788);
nand U16215 (N_16215,N_9256,N_8818);
or U16216 (N_16216,N_10127,N_11098);
nor U16217 (N_16217,N_9507,N_8061);
nor U16218 (N_16218,N_10527,N_8656);
or U16219 (N_16219,N_9291,N_11565);
nor U16220 (N_16220,N_6944,N_11684);
nor U16221 (N_16221,N_8334,N_11984);
and U16222 (N_16222,N_9849,N_6356);
xnor U16223 (N_16223,N_9820,N_10448);
and U16224 (N_16224,N_11183,N_9708);
or U16225 (N_16225,N_9514,N_10828);
nor U16226 (N_16226,N_9954,N_7658);
nor U16227 (N_16227,N_8735,N_7448);
and U16228 (N_16228,N_7000,N_11807);
or U16229 (N_16229,N_11983,N_8121);
xnor U16230 (N_16230,N_9933,N_8442);
or U16231 (N_16231,N_11556,N_10161);
and U16232 (N_16232,N_6697,N_11698);
and U16233 (N_16233,N_8373,N_8577);
nor U16234 (N_16234,N_9709,N_11694);
and U16235 (N_16235,N_7075,N_11794);
and U16236 (N_16236,N_7363,N_7500);
and U16237 (N_16237,N_10865,N_9012);
nor U16238 (N_16238,N_11078,N_10490);
or U16239 (N_16239,N_7759,N_10896);
xor U16240 (N_16240,N_10471,N_8446);
and U16241 (N_16241,N_6602,N_10554);
nor U16242 (N_16242,N_7095,N_8129);
or U16243 (N_16243,N_7392,N_11837);
or U16244 (N_16244,N_6526,N_7452);
and U16245 (N_16245,N_10575,N_7233);
nand U16246 (N_16246,N_8698,N_10443);
nor U16247 (N_16247,N_9395,N_10640);
or U16248 (N_16248,N_7594,N_10342);
nand U16249 (N_16249,N_6425,N_11085);
or U16250 (N_16250,N_9426,N_10951);
or U16251 (N_16251,N_6563,N_11061);
or U16252 (N_16252,N_9593,N_7019);
xor U16253 (N_16253,N_6170,N_7058);
xor U16254 (N_16254,N_9552,N_11259);
or U16255 (N_16255,N_6087,N_11670);
nor U16256 (N_16256,N_8194,N_6465);
xnor U16257 (N_16257,N_6214,N_6501);
or U16258 (N_16258,N_10140,N_7116);
nor U16259 (N_16259,N_9980,N_9672);
xor U16260 (N_16260,N_6841,N_6412);
xor U16261 (N_16261,N_7081,N_9797);
xor U16262 (N_16262,N_10842,N_9947);
and U16263 (N_16263,N_9510,N_11916);
or U16264 (N_16264,N_8813,N_9853);
xor U16265 (N_16265,N_6273,N_6138);
nand U16266 (N_16266,N_6847,N_9095);
and U16267 (N_16267,N_8569,N_8303);
nand U16268 (N_16268,N_10953,N_11538);
and U16269 (N_16269,N_9771,N_7386);
xor U16270 (N_16270,N_10200,N_6040);
nor U16271 (N_16271,N_7612,N_7436);
and U16272 (N_16272,N_9130,N_10314);
xnor U16273 (N_16273,N_7876,N_9003);
nand U16274 (N_16274,N_7084,N_6347);
or U16275 (N_16275,N_10023,N_11768);
and U16276 (N_16276,N_8880,N_6458);
nor U16277 (N_16277,N_9039,N_7231);
xor U16278 (N_16278,N_9731,N_8968);
xnor U16279 (N_16279,N_6996,N_8291);
nand U16280 (N_16280,N_8468,N_11436);
nor U16281 (N_16281,N_7804,N_7090);
nand U16282 (N_16282,N_11931,N_10658);
and U16283 (N_16283,N_9478,N_7872);
or U16284 (N_16284,N_11189,N_11087);
nor U16285 (N_16285,N_9279,N_6786);
nor U16286 (N_16286,N_10070,N_7489);
or U16287 (N_16287,N_7169,N_11677);
and U16288 (N_16288,N_8029,N_6306);
nor U16289 (N_16289,N_10795,N_6160);
xor U16290 (N_16290,N_7276,N_8515);
nor U16291 (N_16291,N_6058,N_8610);
nand U16292 (N_16292,N_6845,N_9855);
nor U16293 (N_16293,N_8914,N_7564);
and U16294 (N_16294,N_10585,N_8642);
nand U16295 (N_16295,N_11166,N_9597);
or U16296 (N_16296,N_8018,N_7835);
or U16297 (N_16297,N_8815,N_10345);
or U16298 (N_16298,N_8478,N_8669);
nor U16299 (N_16299,N_10499,N_8130);
nand U16300 (N_16300,N_11640,N_10636);
nand U16301 (N_16301,N_6939,N_6216);
xnor U16302 (N_16302,N_10825,N_8071);
and U16303 (N_16303,N_7094,N_11451);
nand U16304 (N_16304,N_11382,N_8668);
and U16305 (N_16305,N_7688,N_7069);
xnor U16306 (N_16306,N_8720,N_10502);
nor U16307 (N_16307,N_10880,N_11262);
nor U16308 (N_16308,N_10706,N_7702);
and U16309 (N_16309,N_8859,N_9090);
xor U16310 (N_16310,N_7797,N_10663);
and U16311 (N_16311,N_11836,N_8994);
xnor U16312 (N_16312,N_6899,N_6712);
xor U16313 (N_16313,N_8982,N_8152);
and U16314 (N_16314,N_6128,N_8678);
or U16315 (N_16315,N_8460,N_11996);
or U16316 (N_16316,N_11791,N_6337);
nor U16317 (N_16317,N_9108,N_7972);
xnor U16318 (N_16318,N_6725,N_6473);
nand U16319 (N_16319,N_9498,N_6292);
and U16320 (N_16320,N_11175,N_6252);
and U16321 (N_16321,N_6644,N_8761);
or U16322 (N_16322,N_10878,N_8620);
xor U16323 (N_16323,N_7298,N_8150);
and U16324 (N_16324,N_11691,N_6019);
xnor U16325 (N_16325,N_8468,N_11772);
nor U16326 (N_16326,N_10875,N_10731);
nand U16327 (N_16327,N_7007,N_11161);
or U16328 (N_16328,N_6901,N_8693);
and U16329 (N_16329,N_10251,N_6386);
nor U16330 (N_16330,N_11639,N_6367);
or U16331 (N_16331,N_11108,N_6319);
or U16332 (N_16332,N_9116,N_10919);
xor U16333 (N_16333,N_11160,N_8952);
xnor U16334 (N_16334,N_9328,N_6817);
and U16335 (N_16335,N_6437,N_11530);
nor U16336 (N_16336,N_7221,N_9386);
xor U16337 (N_16337,N_8181,N_7346);
and U16338 (N_16338,N_6279,N_11007);
nand U16339 (N_16339,N_6111,N_7453);
xnor U16340 (N_16340,N_10546,N_11774);
nor U16341 (N_16341,N_8188,N_6459);
xor U16342 (N_16342,N_7128,N_8940);
or U16343 (N_16343,N_7989,N_6028);
and U16344 (N_16344,N_10125,N_8113);
or U16345 (N_16345,N_8804,N_10113);
nor U16346 (N_16346,N_11869,N_10616);
and U16347 (N_16347,N_7069,N_7406);
and U16348 (N_16348,N_8571,N_7461);
or U16349 (N_16349,N_6847,N_6705);
nor U16350 (N_16350,N_9534,N_11141);
or U16351 (N_16351,N_10023,N_7906);
or U16352 (N_16352,N_9741,N_8444);
nand U16353 (N_16353,N_9356,N_7482);
xor U16354 (N_16354,N_11198,N_7710);
xnor U16355 (N_16355,N_9890,N_8252);
and U16356 (N_16356,N_6225,N_9087);
xnor U16357 (N_16357,N_11567,N_7480);
or U16358 (N_16358,N_10878,N_10057);
and U16359 (N_16359,N_10044,N_6295);
xor U16360 (N_16360,N_11977,N_7887);
or U16361 (N_16361,N_9412,N_8149);
or U16362 (N_16362,N_6283,N_11731);
and U16363 (N_16363,N_7050,N_11856);
or U16364 (N_16364,N_6435,N_10359);
xor U16365 (N_16365,N_10412,N_6218);
nand U16366 (N_16366,N_6985,N_6021);
and U16367 (N_16367,N_7153,N_11311);
and U16368 (N_16368,N_6347,N_8860);
xnor U16369 (N_16369,N_7139,N_10636);
nor U16370 (N_16370,N_6104,N_6500);
and U16371 (N_16371,N_10971,N_6895);
and U16372 (N_16372,N_7636,N_10350);
nand U16373 (N_16373,N_11756,N_8572);
or U16374 (N_16374,N_11078,N_7069);
xor U16375 (N_16375,N_8655,N_6544);
nand U16376 (N_16376,N_10587,N_7096);
xnor U16377 (N_16377,N_10817,N_11199);
nor U16378 (N_16378,N_9032,N_11783);
and U16379 (N_16379,N_7799,N_11035);
nor U16380 (N_16380,N_8034,N_8403);
nor U16381 (N_16381,N_6062,N_8684);
or U16382 (N_16382,N_9933,N_8082);
and U16383 (N_16383,N_6983,N_7828);
nor U16384 (N_16384,N_11443,N_11737);
nand U16385 (N_16385,N_10259,N_10960);
and U16386 (N_16386,N_9195,N_7066);
nand U16387 (N_16387,N_8965,N_6844);
or U16388 (N_16388,N_11198,N_7224);
nor U16389 (N_16389,N_6045,N_11537);
nand U16390 (N_16390,N_10479,N_9708);
or U16391 (N_16391,N_8645,N_9247);
xor U16392 (N_16392,N_7267,N_10566);
and U16393 (N_16393,N_9191,N_9957);
xnor U16394 (N_16394,N_10230,N_11409);
nor U16395 (N_16395,N_7933,N_9623);
and U16396 (N_16396,N_6253,N_11232);
nor U16397 (N_16397,N_11526,N_7467);
nand U16398 (N_16398,N_8713,N_8376);
and U16399 (N_16399,N_9621,N_7722);
xor U16400 (N_16400,N_10546,N_10281);
or U16401 (N_16401,N_6293,N_6798);
and U16402 (N_16402,N_9702,N_9798);
and U16403 (N_16403,N_10866,N_11476);
nor U16404 (N_16404,N_7401,N_6317);
or U16405 (N_16405,N_9504,N_11668);
and U16406 (N_16406,N_11453,N_8860);
and U16407 (N_16407,N_6756,N_11877);
nor U16408 (N_16408,N_7071,N_6023);
and U16409 (N_16409,N_10488,N_10029);
xnor U16410 (N_16410,N_9146,N_7719);
or U16411 (N_16411,N_10572,N_6341);
xor U16412 (N_16412,N_9773,N_7999);
xor U16413 (N_16413,N_8880,N_7442);
or U16414 (N_16414,N_7822,N_6818);
and U16415 (N_16415,N_11396,N_9203);
and U16416 (N_16416,N_6347,N_11097);
or U16417 (N_16417,N_8175,N_8070);
nand U16418 (N_16418,N_9154,N_11934);
nor U16419 (N_16419,N_11624,N_11566);
nand U16420 (N_16420,N_6609,N_7314);
nand U16421 (N_16421,N_11023,N_6526);
nor U16422 (N_16422,N_11117,N_11313);
xnor U16423 (N_16423,N_10681,N_7259);
xor U16424 (N_16424,N_6261,N_6723);
or U16425 (N_16425,N_8346,N_9577);
or U16426 (N_16426,N_6769,N_6654);
and U16427 (N_16427,N_11510,N_10104);
or U16428 (N_16428,N_11942,N_8197);
nand U16429 (N_16429,N_11139,N_10794);
or U16430 (N_16430,N_11140,N_6194);
nor U16431 (N_16431,N_6402,N_6885);
or U16432 (N_16432,N_11530,N_11192);
and U16433 (N_16433,N_10523,N_10702);
xnor U16434 (N_16434,N_6024,N_9045);
or U16435 (N_16435,N_6449,N_9286);
and U16436 (N_16436,N_6434,N_6855);
and U16437 (N_16437,N_8483,N_8032);
and U16438 (N_16438,N_6428,N_6498);
xor U16439 (N_16439,N_10549,N_9759);
and U16440 (N_16440,N_9587,N_8922);
nor U16441 (N_16441,N_7936,N_10716);
or U16442 (N_16442,N_10879,N_10984);
xnor U16443 (N_16443,N_8573,N_9785);
nor U16444 (N_16444,N_11705,N_10202);
nand U16445 (N_16445,N_10652,N_7898);
xnor U16446 (N_16446,N_8687,N_8233);
nor U16447 (N_16447,N_7700,N_11327);
and U16448 (N_16448,N_10712,N_8513);
nand U16449 (N_16449,N_8756,N_10038);
xnor U16450 (N_16450,N_6332,N_9913);
nand U16451 (N_16451,N_10133,N_8802);
nand U16452 (N_16452,N_7074,N_6575);
nor U16453 (N_16453,N_8385,N_7274);
and U16454 (N_16454,N_7029,N_11898);
or U16455 (N_16455,N_11843,N_10040);
nand U16456 (N_16456,N_7515,N_6110);
xor U16457 (N_16457,N_8732,N_7650);
or U16458 (N_16458,N_9920,N_6626);
and U16459 (N_16459,N_7551,N_6715);
and U16460 (N_16460,N_7996,N_7590);
nor U16461 (N_16461,N_7665,N_11831);
or U16462 (N_16462,N_7621,N_11123);
nor U16463 (N_16463,N_11763,N_10121);
xor U16464 (N_16464,N_7756,N_11478);
xnor U16465 (N_16465,N_8755,N_7200);
or U16466 (N_16466,N_9330,N_10535);
and U16467 (N_16467,N_9889,N_10032);
nor U16468 (N_16468,N_11171,N_7720);
nand U16469 (N_16469,N_8860,N_7536);
nor U16470 (N_16470,N_7344,N_10831);
or U16471 (N_16471,N_6198,N_9939);
nand U16472 (N_16472,N_6166,N_11877);
nand U16473 (N_16473,N_10740,N_11597);
and U16474 (N_16474,N_8191,N_7222);
xor U16475 (N_16475,N_9880,N_10422);
or U16476 (N_16476,N_11132,N_7011);
and U16477 (N_16477,N_8294,N_7942);
or U16478 (N_16478,N_7154,N_9641);
or U16479 (N_16479,N_6382,N_8931);
xnor U16480 (N_16480,N_11763,N_9346);
or U16481 (N_16481,N_7923,N_8611);
or U16482 (N_16482,N_10308,N_6844);
nor U16483 (N_16483,N_7891,N_7468);
xor U16484 (N_16484,N_11851,N_6824);
nand U16485 (N_16485,N_9678,N_10011);
or U16486 (N_16486,N_10456,N_6741);
xor U16487 (N_16487,N_9940,N_10688);
xor U16488 (N_16488,N_8286,N_11315);
nand U16489 (N_16489,N_11204,N_8538);
nor U16490 (N_16490,N_7056,N_8104);
nor U16491 (N_16491,N_8405,N_8718);
nor U16492 (N_16492,N_11894,N_8833);
xnor U16493 (N_16493,N_9851,N_9070);
nor U16494 (N_16494,N_6521,N_8905);
and U16495 (N_16495,N_8890,N_9965);
nor U16496 (N_16496,N_6788,N_6771);
or U16497 (N_16497,N_7935,N_7162);
nor U16498 (N_16498,N_7247,N_8821);
nor U16499 (N_16499,N_6780,N_7565);
or U16500 (N_16500,N_6202,N_10643);
and U16501 (N_16501,N_9619,N_8495);
and U16502 (N_16502,N_7351,N_9139);
nand U16503 (N_16503,N_8794,N_10475);
or U16504 (N_16504,N_7690,N_6264);
or U16505 (N_16505,N_7593,N_9454);
and U16506 (N_16506,N_8004,N_9645);
nor U16507 (N_16507,N_6405,N_11878);
and U16508 (N_16508,N_10555,N_11448);
or U16509 (N_16509,N_10736,N_8096);
nand U16510 (N_16510,N_11847,N_11306);
or U16511 (N_16511,N_11294,N_6639);
and U16512 (N_16512,N_10555,N_10080);
nor U16513 (N_16513,N_11331,N_9142);
nor U16514 (N_16514,N_9502,N_8162);
xor U16515 (N_16515,N_9347,N_8933);
and U16516 (N_16516,N_11652,N_11314);
nor U16517 (N_16517,N_6255,N_11628);
and U16518 (N_16518,N_11855,N_10320);
nor U16519 (N_16519,N_8708,N_8241);
and U16520 (N_16520,N_11608,N_8137);
and U16521 (N_16521,N_7642,N_6576);
and U16522 (N_16522,N_11201,N_8673);
or U16523 (N_16523,N_9082,N_8471);
nand U16524 (N_16524,N_7282,N_7542);
nand U16525 (N_16525,N_8024,N_9615);
nor U16526 (N_16526,N_8440,N_8020);
and U16527 (N_16527,N_10434,N_8604);
xnor U16528 (N_16528,N_11536,N_11156);
and U16529 (N_16529,N_10253,N_10769);
nand U16530 (N_16530,N_10699,N_6649);
nor U16531 (N_16531,N_11358,N_7310);
and U16532 (N_16532,N_8444,N_11295);
and U16533 (N_16533,N_9383,N_6027);
nand U16534 (N_16534,N_6716,N_9076);
or U16535 (N_16535,N_11737,N_6097);
nand U16536 (N_16536,N_8207,N_7004);
nor U16537 (N_16537,N_11979,N_6557);
and U16538 (N_16538,N_7074,N_6585);
nor U16539 (N_16539,N_7283,N_10213);
nand U16540 (N_16540,N_7376,N_7018);
xnor U16541 (N_16541,N_10809,N_10278);
nor U16542 (N_16542,N_8373,N_10617);
and U16543 (N_16543,N_10303,N_7387);
and U16544 (N_16544,N_10009,N_8106);
nand U16545 (N_16545,N_11796,N_9986);
nor U16546 (N_16546,N_9932,N_6326);
xnor U16547 (N_16547,N_8027,N_10543);
and U16548 (N_16548,N_11021,N_11865);
xor U16549 (N_16549,N_7420,N_9537);
xnor U16550 (N_16550,N_9116,N_11267);
nand U16551 (N_16551,N_11656,N_9639);
xnor U16552 (N_16552,N_11046,N_7738);
xor U16553 (N_16553,N_8618,N_8839);
nand U16554 (N_16554,N_7620,N_6248);
and U16555 (N_16555,N_8338,N_9183);
xnor U16556 (N_16556,N_6807,N_8608);
and U16557 (N_16557,N_9338,N_7947);
xnor U16558 (N_16558,N_7814,N_7190);
and U16559 (N_16559,N_9444,N_11522);
or U16560 (N_16560,N_10199,N_10637);
or U16561 (N_16561,N_10425,N_9841);
or U16562 (N_16562,N_6263,N_10504);
xnor U16563 (N_16563,N_8614,N_9624);
and U16564 (N_16564,N_9936,N_10176);
xnor U16565 (N_16565,N_8370,N_6996);
xnor U16566 (N_16566,N_9025,N_9390);
nand U16567 (N_16567,N_8732,N_6736);
xor U16568 (N_16568,N_6717,N_10896);
xor U16569 (N_16569,N_7927,N_10465);
nor U16570 (N_16570,N_8790,N_7911);
or U16571 (N_16571,N_8291,N_7459);
and U16572 (N_16572,N_8279,N_8198);
or U16573 (N_16573,N_10966,N_6321);
or U16574 (N_16574,N_11054,N_11688);
and U16575 (N_16575,N_10309,N_10848);
or U16576 (N_16576,N_9878,N_7943);
or U16577 (N_16577,N_11562,N_9467);
or U16578 (N_16578,N_9028,N_8935);
nand U16579 (N_16579,N_10278,N_7883);
nand U16580 (N_16580,N_7541,N_9437);
nand U16581 (N_16581,N_9026,N_6884);
nor U16582 (N_16582,N_9858,N_9624);
and U16583 (N_16583,N_9333,N_11190);
nor U16584 (N_16584,N_11509,N_8506);
nand U16585 (N_16585,N_8687,N_6292);
nand U16586 (N_16586,N_11104,N_10194);
and U16587 (N_16587,N_6936,N_10463);
nor U16588 (N_16588,N_9090,N_10294);
nand U16589 (N_16589,N_9712,N_11090);
or U16590 (N_16590,N_10641,N_6825);
nor U16591 (N_16591,N_7429,N_9430);
xor U16592 (N_16592,N_7510,N_7943);
nor U16593 (N_16593,N_9432,N_6166);
and U16594 (N_16594,N_10502,N_10483);
nor U16595 (N_16595,N_10318,N_7907);
nand U16596 (N_16596,N_9591,N_6269);
nand U16597 (N_16597,N_11488,N_9992);
xnor U16598 (N_16598,N_11439,N_7400);
xnor U16599 (N_16599,N_9126,N_8135);
xor U16600 (N_16600,N_10177,N_9455);
nor U16601 (N_16601,N_7903,N_8537);
nor U16602 (N_16602,N_6538,N_8086);
and U16603 (N_16603,N_8265,N_11949);
nor U16604 (N_16604,N_9309,N_11805);
nand U16605 (N_16605,N_6384,N_8743);
xnor U16606 (N_16606,N_8468,N_9916);
nor U16607 (N_16607,N_6885,N_10205);
or U16608 (N_16608,N_6213,N_10431);
or U16609 (N_16609,N_8579,N_6529);
or U16610 (N_16610,N_11511,N_7609);
and U16611 (N_16611,N_6971,N_11288);
nor U16612 (N_16612,N_9154,N_11774);
xor U16613 (N_16613,N_9576,N_8594);
nor U16614 (N_16614,N_6802,N_9974);
or U16615 (N_16615,N_7976,N_6384);
or U16616 (N_16616,N_6152,N_7057);
and U16617 (N_16617,N_10763,N_9571);
or U16618 (N_16618,N_7631,N_6314);
xnor U16619 (N_16619,N_6500,N_6464);
xnor U16620 (N_16620,N_6105,N_10369);
or U16621 (N_16621,N_10728,N_6575);
or U16622 (N_16622,N_10830,N_11812);
and U16623 (N_16623,N_7528,N_10489);
nor U16624 (N_16624,N_10768,N_6856);
nor U16625 (N_16625,N_6515,N_7723);
nand U16626 (N_16626,N_6331,N_7962);
and U16627 (N_16627,N_8815,N_8998);
nand U16628 (N_16628,N_7952,N_8221);
xnor U16629 (N_16629,N_6497,N_7202);
xnor U16630 (N_16630,N_11026,N_11322);
xor U16631 (N_16631,N_9279,N_7925);
nor U16632 (N_16632,N_6203,N_6364);
and U16633 (N_16633,N_7259,N_6059);
or U16634 (N_16634,N_6961,N_9079);
nand U16635 (N_16635,N_8079,N_9972);
and U16636 (N_16636,N_8765,N_6660);
nand U16637 (N_16637,N_10536,N_11895);
or U16638 (N_16638,N_7022,N_9029);
nor U16639 (N_16639,N_7931,N_11703);
or U16640 (N_16640,N_8817,N_9875);
nand U16641 (N_16641,N_10009,N_10173);
xnor U16642 (N_16642,N_11697,N_7322);
xnor U16643 (N_16643,N_10272,N_10538);
nand U16644 (N_16644,N_11645,N_10705);
and U16645 (N_16645,N_8485,N_8080);
nor U16646 (N_16646,N_8878,N_6973);
xnor U16647 (N_16647,N_10218,N_8476);
xor U16648 (N_16648,N_11332,N_8085);
nand U16649 (N_16649,N_7150,N_6825);
nand U16650 (N_16650,N_6729,N_10652);
nor U16651 (N_16651,N_11703,N_10419);
nand U16652 (N_16652,N_7537,N_9120);
xnor U16653 (N_16653,N_10239,N_6161);
xnor U16654 (N_16654,N_9549,N_9316);
nand U16655 (N_16655,N_6289,N_6575);
and U16656 (N_16656,N_8900,N_10864);
or U16657 (N_16657,N_7807,N_11925);
or U16658 (N_16658,N_10455,N_11137);
nor U16659 (N_16659,N_7477,N_6484);
nand U16660 (N_16660,N_7591,N_11627);
or U16661 (N_16661,N_9052,N_8334);
or U16662 (N_16662,N_8376,N_7563);
xor U16663 (N_16663,N_9467,N_8995);
xor U16664 (N_16664,N_7525,N_9981);
or U16665 (N_16665,N_10728,N_6669);
nor U16666 (N_16666,N_10451,N_6538);
nand U16667 (N_16667,N_7266,N_7609);
and U16668 (N_16668,N_10168,N_7447);
nor U16669 (N_16669,N_9556,N_10640);
nor U16670 (N_16670,N_7446,N_10816);
or U16671 (N_16671,N_9092,N_11474);
or U16672 (N_16672,N_9622,N_10457);
nor U16673 (N_16673,N_10106,N_10065);
xnor U16674 (N_16674,N_9082,N_6573);
xnor U16675 (N_16675,N_7563,N_11835);
xnor U16676 (N_16676,N_11843,N_10237);
nand U16677 (N_16677,N_6379,N_7935);
and U16678 (N_16678,N_7480,N_8024);
xnor U16679 (N_16679,N_10241,N_9305);
nand U16680 (N_16680,N_7552,N_11682);
nand U16681 (N_16681,N_11157,N_11339);
nor U16682 (N_16682,N_11922,N_6558);
and U16683 (N_16683,N_7131,N_6147);
nor U16684 (N_16684,N_6755,N_8351);
nand U16685 (N_16685,N_10647,N_6943);
nor U16686 (N_16686,N_10429,N_11195);
and U16687 (N_16687,N_6515,N_6405);
or U16688 (N_16688,N_7733,N_11210);
nor U16689 (N_16689,N_10817,N_10279);
and U16690 (N_16690,N_6706,N_8774);
nand U16691 (N_16691,N_6680,N_11613);
nand U16692 (N_16692,N_10770,N_8276);
xor U16693 (N_16693,N_10705,N_10421);
nor U16694 (N_16694,N_6408,N_10840);
nand U16695 (N_16695,N_9543,N_6798);
xor U16696 (N_16696,N_6433,N_11587);
xnor U16697 (N_16697,N_7904,N_8550);
or U16698 (N_16698,N_9417,N_11739);
xnor U16699 (N_16699,N_8517,N_9854);
nand U16700 (N_16700,N_7134,N_11227);
nand U16701 (N_16701,N_9894,N_6541);
nand U16702 (N_16702,N_10944,N_8826);
nor U16703 (N_16703,N_10497,N_11813);
xnor U16704 (N_16704,N_8699,N_8131);
xnor U16705 (N_16705,N_6739,N_7463);
nor U16706 (N_16706,N_11932,N_6586);
nor U16707 (N_16707,N_11853,N_6281);
and U16708 (N_16708,N_11913,N_10320);
nor U16709 (N_16709,N_11088,N_8185);
or U16710 (N_16710,N_9443,N_8716);
or U16711 (N_16711,N_7396,N_8683);
or U16712 (N_16712,N_9196,N_9013);
and U16713 (N_16713,N_8829,N_8124);
nor U16714 (N_16714,N_9917,N_8160);
and U16715 (N_16715,N_10574,N_10615);
nand U16716 (N_16716,N_7108,N_9716);
xnor U16717 (N_16717,N_10657,N_7589);
xor U16718 (N_16718,N_10937,N_6726);
or U16719 (N_16719,N_10927,N_8407);
or U16720 (N_16720,N_11828,N_7052);
nor U16721 (N_16721,N_11938,N_7361);
nor U16722 (N_16722,N_6169,N_9317);
and U16723 (N_16723,N_9218,N_9983);
or U16724 (N_16724,N_10189,N_6606);
or U16725 (N_16725,N_7020,N_6790);
xor U16726 (N_16726,N_11370,N_6683);
and U16727 (N_16727,N_6237,N_8672);
xnor U16728 (N_16728,N_9710,N_10746);
and U16729 (N_16729,N_9603,N_10226);
xor U16730 (N_16730,N_8350,N_7845);
or U16731 (N_16731,N_11886,N_9831);
nor U16732 (N_16732,N_11614,N_11974);
or U16733 (N_16733,N_6216,N_6625);
and U16734 (N_16734,N_7461,N_7561);
nand U16735 (N_16735,N_10335,N_6714);
or U16736 (N_16736,N_7790,N_8820);
or U16737 (N_16737,N_7480,N_8868);
nand U16738 (N_16738,N_10633,N_6539);
and U16739 (N_16739,N_11990,N_9662);
nor U16740 (N_16740,N_10792,N_8624);
nand U16741 (N_16741,N_10452,N_6372);
xnor U16742 (N_16742,N_11941,N_11718);
nor U16743 (N_16743,N_7889,N_8329);
nor U16744 (N_16744,N_11220,N_10399);
and U16745 (N_16745,N_7844,N_9507);
or U16746 (N_16746,N_9392,N_10016);
nor U16747 (N_16747,N_7859,N_6026);
xor U16748 (N_16748,N_6944,N_11871);
and U16749 (N_16749,N_6891,N_7943);
and U16750 (N_16750,N_8366,N_6732);
nand U16751 (N_16751,N_9170,N_7267);
nor U16752 (N_16752,N_10489,N_10298);
nor U16753 (N_16753,N_6287,N_6527);
nor U16754 (N_16754,N_10788,N_7770);
xor U16755 (N_16755,N_11001,N_8887);
and U16756 (N_16756,N_8128,N_11040);
or U16757 (N_16757,N_11480,N_10264);
xor U16758 (N_16758,N_11000,N_9284);
xnor U16759 (N_16759,N_6115,N_11477);
nor U16760 (N_16760,N_10082,N_10190);
and U16761 (N_16761,N_7744,N_6528);
nand U16762 (N_16762,N_6154,N_8164);
or U16763 (N_16763,N_6345,N_9401);
nor U16764 (N_16764,N_8532,N_10815);
nand U16765 (N_16765,N_11985,N_6199);
nor U16766 (N_16766,N_8055,N_11245);
nand U16767 (N_16767,N_9353,N_10918);
xor U16768 (N_16768,N_6867,N_11904);
nor U16769 (N_16769,N_9680,N_10542);
nand U16770 (N_16770,N_10628,N_6169);
nand U16771 (N_16771,N_8712,N_9832);
nor U16772 (N_16772,N_8524,N_7133);
and U16773 (N_16773,N_10114,N_11976);
or U16774 (N_16774,N_9124,N_11105);
nor U16775 (N_16775,N_9051,N_7845);
or U16776 (N_16776,N_7286,N_10386);
or U16777 (N_16777,N_7341,N_11622);
nand U16778 (N_16778,N_10271,N_9778);
nor U16779 (N_16779,N_8634,N_9323);
nor U16780 (N_16780,N_9927,N_10163);
xor U16781 (N_16781,N_11001,N_9761);
xnor U16782 (N_16782,N_10006,N_6864);
nand U16783 (N_16783,N_8396,N_11261);
or U16784 (N_16784,N_6532,N_11166);
or U16785 (N_16785,N_7108,N_10707);
xor U16786 (N_16786,N_6018,N_7401);
or U16787 (N_16787,N_6260,N_10503);
or U16788 (N_16788,N_11506,N_6734);
nand U16789 (N_16789,N_8045,N_9973);
nor U16790 (N_16790,N_6774,N_7226);
and U16791 (N_16791,N_6032,N_10945);
xor U16792 (N_16792,N_6958,N_6742);
xnor U16793 (N_16793,N_6083,N_7372);
xor U16794 (N_16794,N_9577,N_7639);
nor U16795 (N_16795,N_6359,N_6910);
nand U16796 (N_16796,N_6376,N_6176);
nor U16797 (N_16797,N_6081,N_11975);
or U16798 (N_16798,N_8254,N_6936);
xnor U16799 (N_16799,N_10213,N_9631);
nor U16800 (N_16800,N_8471,N_10151);
nor U16801 (N_16801,N_11178,N_6270);
xnor U16802 (N_16802,N_8403,N_6027);
nor U16803 (N_16803,N_9396,N_10874);
xnor U16804 (N_16804,N_8334,N_10109);
nor U16805 (N_16805,N_6034,N_8741);
nor U16806 (N_16806,N_8104,N_6847);
or U16807 (N_16807,N_7325,N_11222);
or U16808 (N_16808,N_8403,N_7228);
xnor U16809 (N_16809,N_7191,N_11584);
nor U16810 (N_16810,N_6965,N_6264);
or U16811 (N_16811,N_11315,N_8005);
and U16812 (N_16812,N_6116,N_6373);
and U16813 (N_16813,N_9138,N_7864);
or U16814 (N_16814,N_9895,N_9260);
nand U16815 (N_16815,N_10024,N_7947);
nor U16816 (N_16816,N_10355,N_9382);
nand U16817 (N_16817,N_7633,N_6635);
nand U16818 (N_16818,N_11933,N_8531);
xor U16819 (N_16819,N_7183,N_8237);
xor U16820 (N_16820,N_6731,N_7947);
xnor U16821 (N_16821,N_10526,N_11859);
or U16822 (N_16822,N_10728,N_11095);
nor U16823 (N_16823,N_11121,N_9117);
nor U16824 (N_16824,N_6866,N_7573);
or U16825 (N_16825,N_6395,N_8837);
nor U16826 (N_16826,N_11259,N_7807);
xor U16827 (N_16827,N_10951,N_11487);
nor U16828 (N_16828,N_8445,N_10391);
xnor U16829 (N_16829,N_8365,N_7472);
or U16830 (N_16830,N_11513,N_10131);
and U16831 (N_16831,N_6092,N_8415);
nor U16832 (N_16832,N_8863,N_6496);
or U16833 (N_16833,N_10262,N_9025);
nor U16834 (N_16834,N_6893,N_10929);
xor U16835 (N_16835,N_10631,N_10924);
and U16836 (N_16836,N_9520,N_8645);
xnor U16837 (N_16837,N_7629,N_10126);
nor U16838 (N_16838,N_6524,N_9786);
and U16839 (N_16839,N_10856,N_11692);
nand U16840 (N_16840,N_7722,N_9163);
xnor U16841 (N_16841,N_7326,N_10715);
and U16842 (N_16842,N_6976,N_8736);
and U16843 (N_16843,N_9541,N_8674);
or U16844 (N_16844,N_9831,N_11903);
nand U16845 (N_16845,N_7528,N_7189);
xor U16846 (N_16846,N_11169,N_9642);
and U16847 (N_16847,N_9884,N_6622);
nor U16848 (N_16848,N_9310,N_7170);
nor U16849 (N_16849,N_8734,N_7350);
and U16850 (N_16850,N_6723,N_7836);
nand U16851 (N_16851,N_7263,N_11565);
or U16852 (N_16852,N_6244,N_11928);
nor U16853 (N_16853,N_6136,N_8639);
and U16854 (N_16854,N_9015,N_7642);
or U16855 (N_16855,N_10390,N_9570);
xnor U16856 (N_16856,N_11951,N_9702);
or U16857 (N_16857,N_9775,N_7781);
and U16858 (N_16858,N_9398,N_10704);
nor U16859 (N_16859,N_10341,N_9060);
xnor U16860 (N_16860,N_7203,N_8566);
xor U16861 (N_16861,N_8434,N_10209);
xnor U16862 (N_16862,N_9289,N_7437);
and U16863 (N_16863,N_11277,N_11953);
or U16864 (N_16864,N_9976,N_9211);
nor U16865 (N_16865,N_6150,N_9035);
and U16866 (N_16866,N_7644,N_8391);
nor U16867 (N_16867,N_10910,N_9399);
and U16868 (N_16868,N_11824,N_8820);
xor U16869 (N_16869,N_6026,N_9953);
nor U16870 (N_16870,N_8709,N_9947);
and U16871 (N_16871,N_6045,N_6475);
or U16872 (N_16872,N_9828,N_9433);
or U16873 (N_16873,N_11145,N_9204);
or U16874 (N_16874,N_6738,N_9487);
nor U16875 (N_16875,N_11739,N_10673);
xnor U16876 (N_16876,N_7288,N_10537);
xor U16877 (N_16877,N_10158,N_11608);
or U16878 (N_16878,N_11661,N_6829);
or U16879 (N_16879,N_8982,N_9261);
or U16880 (N_16880,N_7037,N_9041);
or U16881 (N_16881,N_9574,N_10311);
nand U16882 (N_16882,N_6465,N_11147);
xor U16883 (N_16883,N_8801,N_11439);
or U16884 (N_16884,N_7322,N_6450);
nor U16885 (N_16885,N_6159,N_10978);
nor U16886 (N_16886,N_10954,N_9241);
nand U16887 (N_16887,N_7800,N_8916);
or U16888 (N_16888,N_9448,N_9276);
and U16889 (N_16889,N_9844,N_7850);
and U16890 (N_16890,N_11820,N_8163);
and U16891 (N_16891,N_9549,N_8348);
nor U16892 (N_16892,N_8994,N_11591);
or U16893 (N_16893,N_10765,N_9879);
nor U16894 (N_16894,N_7259,N_6832);
or U16895 (N_16895,N_6671,N_8654);
and U16896 (N_16896,N_11749,N_11856);
xor U16897 (N_16897,N_10841,N_6039);
or U16898 (N_16898,N_6620,N_9470);
nor U16899 (N_16899,N_7081,N_6989);
xnor U16900 (N_16900,N_10075,N_9229);
xor U16901 (N_16901,N_6865,N_10331);
or U16902 (N_16902,N_6563,N_9577);
or U16903 (N_16903,N_6828,N_11592);
xnor U16904 (N_16904,N_8650,N_9493);
xor U16905 (N_16905,N_10556,N_8410);
or U16906 (N_16906,N_9298,N_8850);
or U16907 (N_16907,N_10499,N_10700);
nor U16908 (N_16908,N_6473,N_8549);
and U16909 (N_16909,N_11267,N_11296);
and U16910 (N_16910,N_10136,N_7050);
or U16911 (N_16911,N_10376,N_6701);
and U16912 (N_16912,N_9895,N_9351);
nand U16913 (N_16913,N_7475,N_8641);
xor U16914 (N_16914,N_8353,N_6086);
xor U16915 (N_16915,N_8211,N_7737);
or U16916 (N_16916,N_11136,N_7126);
and U16917 (N_16917,N_7531,N_6189);
and U16918 (N_16918,N_9592,N_10446);
xnor U16919 (N_16919,N_8169,N_6255);
or U16920 (N_16920,N_8531,N_8258);
nand U16921 (N_16921,N_10970,N_8590);
nand U16922 (N_16922,N_9855,N_6106);
and U16923 (N_16923,N_8364,N_9431);
nand U16924 (N_16924,N_8132,N_10177);
and U16925 (N_16925,N_9688,N_6027);
nand U16926 (N_16926,N_10709,N_11141);
nor U16927 (N_16927,N_11328,N_11372);
and U16928 (N_16928,N_6942,N_8125);
nand U16929 (N_16929,N_9340,N_11253);
and U16930 (N_16930,N_8551,N_9813);
or U16931 (N_16931,N_8047,N_9250);
and U16932 (N_16932,N_8945,N_7486);
nor U16933 (N_16933,N_11710,N_9823);
and U16934 (N_16934,N_10777,N_6877);
or U16935 (N_16935,N_9097,N_10892);
nand U16936 (N_16936,N_9681,N_7286);
xor U16937 (N_16937,N_7260,N_6946);
and U16938 (N_16938,N_8135,N_10435);
xor U16939 (N_16939,N_7173,N_6847);
xnor U16940 (N_16940,N_6740,N_6977);
and U16941 (N_16941,N_7257,N_6761);
or U16942 (N_16942,N_6093,N_7889);
and U16943 (N_16943,N_10538,N_7365);
nand U16944 (N_16944,N_7674,N_6737);
nor U16945 (N_16945,N_9485,N_8858);
nor U16946 (N_16946,N_7619,N_7761);
and U16947 (N_16947,N_6876,N_6999);
nand U16948 (N_16948,N_10781,N_9069);
or U16949 (N_16949,N_11305,N_8981);
xor U16950 (N_16950,N_7041,N_7219);
nand U16951 (N_16951,N_8468,N_6772);
nor U16952 (N_16952,N_10543,N_9857);
or U16953 (N_16953,N_9737,N_7966);
and U16954 (N_16954,N_10975,N_11924);
and U16955 (N_16955,N_6623,N_9637);
nor U16956 (N_16956,N_11405,N_7353);
and U16957 (N_16957,N_11680,N_6540);
nand U16958 (N_16958,N_10756,N_9401);
nor U16959 (N_16959,N_11538,N_7682);
or U16960 (N_16960,N_8667,N_9218);
and U16961 (N_16961,N_11945,N_9091);
or U16962 (N_16962,N_8596,N_11413);
nor U16963 (N_16963,N_9116,N_6036);
nor U16964 (N_16964,N_9602,N_8085);
nor U16965 (N_16965,N_7428,N_11328);
nand U16966 (N_16966,N_7667,N_9543);
xor U16967 (N_16967,N_8398,N_8927);
and U16968 (N_16968,N_8453,N_10209);
or U16969 (N_16969,N_11124,N_9162);
and U16970 (N_16970,N_8940,N_8585);
nand U16971 (N_16971,N_6542,N_11916);
or U16972 (N_16972,N_9962,N_6632);
or U16973 (N_16973,N_10626,N_7219);
or U16974 (N_16974,N_6829,N_11325);
nor U16975 (N_16975,N_10807,N_6506);
and U16976 (N_16976,N_6777,N_9688);
xor U16977 (N_16977,N_7678,N_7552);
xnor U16978 (N_16978,N_6421,N_6184);
or U16979 (N_16979,N_8523,N_7324);
xnor U16980 (N_16980,N_11723,N_6082);
xnor U16981 (N_16981,N_7748,N_9131);
nor U16982 (N_16982,N_8371,N_7341);
or U16983 (N_16983,N_7735,N_7906);
or U16984 (N_16984,N_7328,N_10102);
xor U16985 (N_16985,N_7357,N_6340);
and U16986 (N_16986,N_8912,N_9719);
and U16987 (N_16987,N_8793,N_11279);
and U16988 (N_16988,N_7370,N_7441);
nor U16989 (N_16989,N_11810,N_10268);
or U16990 (N_16990,N_9916,N_8813);
nor U16991 (N_16991,N_10703,N_8394);
and U16992 (N_16992,N_8909,N_10890);
xor U16993 (N_16993,N_11784,N_8007);
nand U16994 (N_16994,N_6016,N_9955);
xnor U16995 (N_16995,N_9168,N_10068);
and U16996 (N_16996,N_8515,N_8692);
nand U16997 (N_16997,N_8418,N_11793);
and U16998 (N_16998,N_9157,N_9920);
nand U16999 (N_16999,N_11406,N_9708);
nand U17000 (N_17000,N_7099,N_8804);
xor U17001 (N_17001,N_7721,N_11439);
xnor U17002 (N_17002,N_9616,N_6906);
and U17003 (N_17003,N_10552,N_10488);
nand U17004 (N_17004,N_11036,N_7973);
or U17005 (N_17005,N_6265,N_7586);
nand U17006 (N_17006,N_6236,N_11432);
nor U17007 (N_17007,N_9677,N_8033);
and U17008 (N_17008,N_10952,N_7628);
xor U17009 (N_17009,N_8938,N_10360);
and U17010 (N_17010,N_7490,N_7932);
and U17011 (N_17011,N_9023,N_7906);
and U17012 (N_17012,N_6548,N_10025);
or U17013 (N_17013,N_8300,N_10010);
and U17014 (N_17014,N_8618,N_8511);
xnor U17015 (N_17015,N_6890,N_8022);
nand U17016 (N_17016,N_9477,N_8307);
and U17017 (N_17017,N_9968,N_7559);
nor U17018 (N_17018,N_10564,N_10654);
xnor U17019 (N_17019,N_7058,N_10312);
xor U17020 (N_17020,N_8222,N_9773);
xor U17021 (N_17021,N_6952,N_8003);
xnor U17022 (N_17022,N_9676,N_9535);
xnor U17023 (N_17023,N_9871,N_11779);
xor U17024 (N_17024,N_7906,N_10063);
or U17025 (N_17025,N_8236,N_6738);
xnor U17026 (N_17026,N_10195,N_9417);
and U17027 (N_17027,N_6682,N_10138);
xor U17028 (N_17028,N_6071,N_8033);
or U17029 (N_17029,N_6374,N_8398);
xnor U17030 (N_17030,N_7704,N_11851);
or U17031 (N_17031,N_6518,N_8045);
nor U17032 (N_17032,N_7372,N_11124);
and U17033 (N_17033,N_10822,N_11697);
nor U17034 (N_17034,N_10678,N_10980);
nand U17035 (N_17035,N_10458,N_6758);
or U17036 (N_17036,N_8385,N_10517);
xor U17037 (N_17037,N_10055,N_9148);
nand U17038 (N_17038,N_10857,N_11948);
nor U17039 (N_17039,N_7041,N_10943);
xnor U17040 (N_17040,N_8881,N_6630);
or U17041 (N_17041,N_11618,N_9857);
and U17042 (N_17042,N_9515,N_6923);
nor U17043 (N_17043,N_6496,N_7789);
xor U17044 (N_17044,N_7734,N_11885);
and U17045 (N_17045,N_11584,N_11519);
and U17046 (N_17046,N_8930,N_7660);
nand U17047 (N_17047,N_11423,N_10518);
or U17048 (N_17048,N_11667,N_10678);
nor U17049 (N_17049,N_9333,N_6996);
xnor U17050 (N_17050,N_7067,N_6813);
and U17051 (N_17051,N_10631,N_9517);
nand U17052 (N_17052,N_10314,N_7250);
nand U17053 (N_17053,N_11268,N_11348);
or U17054 (N_17054,N_6604,N_9398);
nand U17055 (N_17055,N_8473,N_7861);
or U17056 (N_17056,N_11838,N_9981);
nand U17057 (N_17057,N_10082,N_9103);
or U17058 (N_17058,N_10480,N_9290);
and U17059 (N_17059,N_9150,N_7559);
nand U17060 (N_17060,N_6026,N_11325);
nor U17061 (N_17061,N_11945,N_6347);
xor U17062 (N_17062,N_7811,N_8337);
and U17063 (N_17063,N_8883,N_7077);
and U17064 (N_17064,N_8290,N_7665);
or U17065 (N_17065,N_10047,N_7953);
xnor U17066 (N_17066,N_6547,N_7490);
xnor U17067 (N_17067,N_9590,N_11521);
nor U17068 (N_17068,N_6709,N_7769);
xor U17069 (N_17069,N_7764,N_10046);
and U17070 (N_17070,N_8388,N_6461);
nor U17071 (N_17071,N_7312,N_7531);
nor U17072 (N_17072,N_10126,N_7391);
xor U17073 (N_17073,N_10510,N_10422);
nor U17074 (N_17074,N_6262,N_11712);
nand U17075 (N_17075,N_6838,N_6146);
nor U17076 (N_17076,N_9054,N_7240);
or U17077 (N_17077,N_10240,N_8859);
and U17078 (N_17078,N_8573,N_9821);
nor U17079 (N_17079,N_9061,N_10758);
nor U17080 (N_17080,N_6230,N_11694);
nand U17081 (N_17081,N_8026,N_6026);
nand U17082 (N_17082,N_6759,N_7286);
and U17083 (N_17083,N_8317,N_8484);
xnor U17084 (N_17084,N_6754,N_6721);
xor U17085 (N_17085,N_8753,N_11278);
nor U17086 (N_17086,N_6688,N_10689);
nand U17087 (N_17087,N_6065,N_6026);
nor U17088 (N_17088,N_8208,N_8650);
or U17089 (N_17089,N_10944,N_6385);
nand U17090 (N_17090,N_10988,N_11698);
and U17091 (N_17091,N_6009,N_8858);
and U17092 (N_17092,N_11547,N_9397);
nor U17093 (N_17093,N_9915,N_6909);
xor U17094 (N_17094,N_11482,N_10636);
nor U17095 (N_17095,N_7129,N_9009);
or U17096 (N_17096,N_11728,N_6068);
and U17097 (N_17097,N_9991,N_8319);
xnor U17098 (N_17098,N_8804,N_9471);
nor U17099 (N_17099,N_6372,N_9161);
nand U17100 (N_17100,N_9346,N_11516);
or U17101 (N_17101,N_8267,N_6975);
and U17102 (N_17102,N_8444,N_8601);
nand U17103 (N_17103,N_7738,N_11244);
nor U17104 (N_17104,N_9550,N_6950);
xnor U17105 (N_17105,N_10038,N_7921);
and U17106 (N_17106,N_7591,N_8536);
and U17107 (N_17107,N_10613,N_8250);
xnor U17108 (N_17108,N_7261,N_7528);
or U17109 (N_17109,N_8119,N_11149);
xnor U17110 (N_17110,N_7191,N_11040);
or U17111 (N_17111,N_6080,N_9114);
or U17112 (N_17112,N_6922,N_7098);
or U17113 (N_17113,N_7667,N_9525);
or U17114 (N_17114,N_11516,N_11278);
xor U17115 (N_17115,N_11353,N_7870);
nand U17116 (N_17116,N_9755,N_7041);
or U17117 (N_17117,N_10812,N_11646);
nand U17118 (N_17118,N_11631,N_8242);
nor U17119 (N_17119,N_9083,N_11546);
and U17120 (N_17120,N_11276,N_10830);
xor U17121 (N_17121,N_11335,N_8696);
or U17122 (N_17122,N_6037,N_6268);
nor U17123 (N_17123,N_7053,N_10719);
nand U17124 (N_17124,N_11935,N_11030);
and U17125 (N_17125,N_8552,N_6269);
nand U17126 (N_17126,N_11847,N_11327);
and U17127 (N_17127,N_8058,N_10908);
nor U17128 (N_17128,N_10291,N_8425);
nor U17129 (N_17129,N_7518,N_6173);
xnor U17130 (N_17130,N_6094,N_9843);
nand U17131 (N_17131,N_8376,N_10644);
nand U17132 (N_17132,N_7877,N_11677);
or U17133 (N_17133,N_6986,N_10951);
nand U17134 (N_17134,N_9902,N_11021);
nand U17135 (N_17135,N_9281,N_7965);
nand U17136 (N_17136,N_7123,N_6260);
xnor U17137 (N_17137,N_6994,N_11696);
nor U17138 (N_17138,N_10357,N_10981);
xnor U17139 (N_17139,N_8901,N_10051);
xnor U17140 (N_17140,N_11794,N_8918);
nand U17141 (N_17141,N_7167,N_9066);
nand U17142 (N_17142,N_10463,N_6170);
and U17143 (N_17143,N_9634,N_11252);
nand U17144 (N_17144,N_7351,N_8775);
nand U17145 (N_17145,N_8382,N_11492);
nor U17146 (N_17146,N_10380,N_9750);
and U17147 (N_17147,N_11959,N_11459);
xnor U17148 (N_17148,N_11661,N_7927);
nor U17149 (N_17149,N_7115,N_8595);
xor U17150 (N_17150,N_11355,N_9450);
xor U17151 (N_17151,N_10391,N_11102);
nor U17152 (N_17152,N_8306,N_8304);
or U17153 (N_17153,N_11361,N_11334);
xor U17154 (N_17154,N_11937,N_10536);
or U17155 (N_17155,N_9799,N_6217);
nand U17156 (N_17156,N_7474,N_10938);
xnor U17157 (N_17157,N_7156,N_9599);
xnor U17158 (N_17158,N_8113,N_8283);
xor U17159 (N_17159,N_11475,N_8425);
and U17160 (N_17160,N_11548,N_8139);
nand U17161 (N_17161,N_6890,N_11687);
nor U17162 (N_17162,N_10867,N_11627);
and U17163 (N_17163,N_6131,N_7090);
or U17164 (N_17164,N_10266,N_8233);
xnor U17165 (N_17165,N_11240,N_11860);
or U17166 (N_17166,N_6220,N_9349);
nor U17167 (N_17167,N_9228,N_6693);
and U17168 (N_17168,N_7807,N_7614);
xnor U17169 (N_17169,N_11006,N_10937);
nor U17170 (N_17170,N_8233,N_9237);
nand U17171 (N_17171,N_7503,N_8335);
nor U17172 (N_17172,N_8704,N_10037);
xnor U17173 (N_17173,N_8607,N_7463);
xnor U17174 (N_17174,N_11381,N_8216);
and U17175 (N_17175,N_6724,N_8146);
or U17176 (N_17176,N_10910,N_8024);
nand U17177 (N_17177,N_6436,N_8023);
or U17178 (N_17178,N_8475,N_11878);
nand U17179 (N_17179,N_6925,N_10176);
or U17180 (N_17180,N_11110,N_11505);
nor U17181 (N_17181,N_8816,N_10771);
nor U17182 (N_17182,N_10152,N_6563);
or U17183 (N_17183,N_8186,N_11360);
nor U17184 (N_17184,N_9674,N_7519);
and U17185 (N_17185,N_8661,N_10000);
nand U17186 (N_17186,N_10353,N_11756);
xor U17187 (N_17187,N_9272,N_6071);
or U17188 (N_17188,N_6249,N_9360);
nor U17189 (N_17189,N_8133,N_10898);
xor U17190 (N_17190,N_10287,N_7336);
nand U17191 (N_17191,N_7304,N_10030);
or U17192 (N_17192,N_8137,N_8122);
nor U17193 (N_17193,N_8834,N_10876);
or U17194 (N_17194,N_7212,N_6984);
nor U17195 (N_17195,N_6522,N_7639);
or U17196 (N_17196,N_11820,N_8805);
nor U17197 (N_17197,N_8712,N_9300);
nor U17198 (N_17198,N_7013,N_11296);
xor U17199 (N_17199,N_8879,N_8905);
and U17200 (N_17200,N_8368,N_8032);
and U17201 (N_17201,N_8847,N_6007);
xor U17202 (N_17202,N_9358,N_9001);
xnor U17203 (N_17203,N_6542,N_8474);
and U17204 (N_17204,N_6913,N_10033);
and U17205 (N_17205,N_11327,N_9332);
nor U17206 (N_17206,N_8807,N_6263);
and U17207 (N_17207,N_11956,N_7012);
or U17208 (N_17208,N_10012,N_11292);
or U17209 (N_17209,N_9326,N_11426);
nor U17210 (N_17210,N_10069,N_8199);
nand U17211 (N_17211,N_10178,N_7534);
nand U17212 (N_17212,N_8771,N_11663);
xnor U17213 (N_17213,N_11074,N_6648);
and U17214 (N_17214,N_11739,N_7726);
xnor U17215 (N_17215,N_7192,N_10871);
xor U17216 (N_17216,N_7157,N_11274);
or U17217 (N_17217,N_6584,N_9964);
xnor U17218 (N_17218,N_10621,N_7655);
and U17219 (N_17219,N_6027,N_11813);
nand U17220 (N_17220,N_11635,N_7740);
nand U17221 (N_17221,N_9648,N_7827);
xnor U17222 (N_17222,N_9429,N_7917);
nand U17223 (N_17223,N_8973,N_8751);
nand U17224 (N_17224,N_8957,N_9411);
xnor U17225 (N_17225,N_9848,N_6195);
xnor U17226 (N_17226,N_8902,N_8251);
nor U17227 (N_17227,N_11119,N_11140);
and U17228 (N_17228,N_6986,N_8249);
or U17229 (N_17229,N_10387,N_10392);
xor U17230 (N_17230,N_9548,N_6609);
and U17231 (N_17231,N_10882,N_10814);
and U17232 (N_17232,N_8509,N_9727);
and U17233 (N_17233,N_9652,N_11070);
xor U17234 (N_17234,N_7266,N_11638);
or U17235 (N_17235,N_10293,N_9675);
nor U17236 (N_17236,N_11248,N_7051);
or U17237 (N_17237,N_10464,N_6866);
and U17238 (N_17238,N_11814,N_10907);
and U17239 (N_17239,N_7495,N_10157);
nand U17240 (N_17240,N_8185,N_9422);
xor U17241 (N_17241,N_6141,N_9227);
xnor U17242 (N_17242,N_9273,N_10403);
nor U17243 (N_17243,N_10275,N_6855);
nor U17244 (N_17244,N_7313,N_11825);
nand U17245 (N_17245,N_10055,N_7911);
or U17246 (N_17246,N_8948,N_9948);
and U17247 (N_17247,N_6009,N_10065);
and U17248 (N_17248,N_6289,N_6751);
and U17249 (N_17249,N_7278,N_10705);
nand U17250 (N_17250,N_10590,N_7578);
or U17251 (N_17251,N_9770,N_10200);
nand U17252 (N_17252,N_7468,N_10533);
and U17253 (N_17253,N_10847,N_10554);
nor U17254 (N_17254,N_6206,N_10437);
nor U17255 (N_17255,N_7266,N_10055);
or U17256 (N_17256,N_8412,N_8813);
and U17257 (N_17257,N_8513,N_11354);
or U17258 (N_17258,N_11253,N_11963);
and U17259 (N_17259,N_8569,N_10773);
nor U17260 (N_17260,N_10512,N_9983);
nand U17261 (N_17261,N_10451,N_10485);
and U17262 (N_17262,N_6736,N_9064);
nand U17263 (N_17263,N_8971,N_10518);
nand U17264 (N_17264,N_6126,N_10990);
nand U17265 (N_17265,N_7007,N_8025);
nor U17266 (N_17266,N_7654,N_7390);
nor U17267 (N_17267,N_8733,N_6677);
nand U17268 (N_17268,N_6887,N_11165);
nor U17269 (N_17269,N_9547,N_7885);
or U17270 (N_17270,N_10625,N_7633);
nor U17271 (N_17271,N_11337,N_9041);
nand U17272 (N_17272,N_11905,N_11889);
and U17273 (N_17273,N_10020,N_8714);
nand U17274 (N_17274,N_9620,N_11248);
nand U17275 (N_17275,N_11548,N_9461);
xor U17276 (N_17276,N_11215,N_11923);
and U17277 (N_17277,N_7780,N_9609);
and U17278 (N_17278,N_7392,N_8003);
nor U17279 (N_17279,N_11351,N_7710);
nand U17280 (N_17280,N_9867,N_11929);
xor U17281 (N_17281,N_8975,N_8389);
nor U17282 (N_17282,N_7212,N_7866);
nand U17283 (N_17283,N_10526,N_7009);
and U17284 (N_17284,N_10262,N_7438);
nand U17285 (N_17285,N_10340,N_6569);
and U17286 (N_17286,N_6753,N_10640);
nand U17287 (N_17287,N_10220,N_11212);
nand U17288 (N_17288,N_8335,N_9521);
nor U17289 (N_17289,N_10000,N_6680);
xnor U17290 (N_17290,N_7706,N_7499);
and U17291 (N_17291,N_9745,N_6231);
xor U17292 (N_17292,N_10426,N_8704);
and U17293 (N_17293,N_6581,N_9795);
nand U17294 (N_17294,N_7016,N_9999);
nor U17295 (N_17295,N_10795,N_9626);
nor U17296 (N_17296,N_8998,N_7139);
nor U17297 (N_17297,N_10227,N_8459);
nand U17298 (N_17298,N_11460,N_9972);
and U17299 (N_17299,N_6047,N_10435);
or U17300 (N_17300,N_8412,N_9457);
nor U17301 (N_17301,N_9600,N_7372);
and U17302 (N_17302,N_10296,N_8516);
or U17303 (N_17303,N_9134,N_7037);
and U17304 (N_17304,N_9184,N_6463);
nand U17305 (N_17305,N_10376,N_7473);
and U17306 (N_17306,N_8541,N_7611);
or U17307 (N_17307,N_7699,N_7567);
nand U17308 (N_17308,N_7278,N_7172);
or U17309 (N_17309,N_8489,N_7228);
nand U17310 (N_17310,N_11720,N_10964);
nor U17311 (N_17311,N_7556,N_10556);
nand U17312 (N_17312,N_9171,N_8861);
and U17313 (N_17313,N_10278,N_11663);
and U17314 (N_17314,N_6900,N_7114);
and U17315 (N_17315,N_9896,N_10213);
and U17316 (N_17316,N_6691,N_8601);
and U17317 (N_17317,N_8263,N_7784);
and U17318 (N_17318,N_6344,N_6556);
xnor U17319 (N_17319,N_10045,N_7065);
or U17320 (N_17320,N_8351,N_8298);
nor U17321 (N_17321,N_8486,N_10263);
xor U17322 (N_17322,N_10196,N_6077);
and U17323 (N_17323,N_6552,N_6511);
and U17324 (N_17324,N_8199,N_8338);
and U17325 (N_17325,N_8399,N_10928);
xnor U17326 (N_17326,N_9133,N_6618);
and U17327 (N_17327,N_7306,N_9412);
or U17328 (N_17328,N_8090,N_7408);
or U17329 (N_17329,N_7143,N_10277);
nor U17330 (N_17330,N_10134,N_11952);
xnor U17331 (N_17331,N_10563,N_9681);
and U17332 (N_17332,N_7791,N_7649);
xor U17333 (N_17333,N_9800,N_10676);
and U17334 (N_17334,N_9262,N_8893);
or U17335 (N_17335,N_11450,N_10515);
or U17336 (N_17336,N_8447,N_6163);
or U17337 (N_17337,N_8345,N_7522);
or U17338 (N_17338,N_11617,N_9387);
nand U17339 (N_17339,N_6935,N_9897);
or U17340 (N_17340,N_6388,N_10183);
xor U17341 (N_17341,N_9600,N_8398);
or U17342 (N_17342,N_10624,N_10486);
xor U17343 (N_17343,N_9985,N_9614);
nor U17344 (N_17344,N_10190,N_8949);
xnor U17345 (N_17345,N_10312,N_11700);
and U17346 (N_17346,N_6153,N_6235);
xnor U17347 (N_17347,N_9331,N_11112);
xor U17348 (N_17348,N_8803,N_9107);
nor U17349 (N_17349,N_8250,N_11671);
nor U17350 (N_17350,N_10148,N_11110);
and U17351 (N_17351,N_6865,N_9379);
nand U17352 (N_17352,N_7521,N_9412);
nand U17353 (N_17353,N_6293,N_10449);
nand U17354 (N_17354,N_11034,N_8697);
xor U17355 (N_17355,N_11298,N_11956);
nand U17356 (N_17356,N_7641,N_9070);
or U17357 (N_17357,N_9438,N_8885);
and U17358 (N_17358,N_11355,N_7953);
nor U17359 (N_17359,N_8427,N_6158);
nand U17360 (N_17360,N_10366,N_9799);
nor U17361 (N_17361,N_7687,N_9984);
xor U17362 (N_17362,N_11000,N_11034);
xnor U17363 (N_17363,N_8065,N_8433);
or U17364 (N_17364,N_10357,N_9610);
or U17365 (N_17365,N_9783,N_9760);
nand U17366 (N_17366,N_6907,N_7428);
nand U17367 (N_17367,N_6412,N_8720);
nand U17368 (N_17368,N_7276,N_8168);
nand U17369 (N_17369,N_7112,N_9071);
nand U17370 (N_17370,N_10477,N_11922);
nand U17371 (N_17371,N_8565,N_11818);
or U17372 (N_17372,N_11735,N_7517);
or U17373 (N_17373,N_11779,N_11525);
nor U17374 (N_17374,N_11072,N_9251);
nand U17375 (N_17375,N_6639,N_9044);
nand U17376 (N_17376,N_8666,N_8742);
and U17377 (N_17377,N_7794,N_8846);
or U17378 (N_17378,N_6265,N_8862);
xor U17379 (N_17379,N_7928,N_6366);
or U17380 (N_17380,N_6995,N_10326);
nor U17381 (N_17381,N_11924,N_6705);
and U17382 (N_17382,N_8572,N_8146);
nor U17383 (N_17383,N_7185,N_8912);
nor U17384 (N_17384,N_7702,N_8440);
nand U17385 (N_17385,N_9587,N_10816);
nand U17386 (N_17386,N_9783,N_8198);
nor U17387 (N_17387,N_10089,N_9051);
or U17388 (N_17388,N_6581,N_9427);
xnor U17389 (N_17389,N_6124,N_10801);
nand U17390 (N_17390,N_7013,N_8683);
nor U17391 (N_17391,N_11556,N_10107);
nand U17392 (N_17392,N_7653,N_6290);
nand U17393 (N_17393,N_7123,N_6346);
nor U17394 (N_17394,N_10019,N_7739);
nand U17395 (N_17395,N_10224,N_9247);
or U17396 (N_17396,N_7347,N_6528);
or U17397 (N_17397,N_11881,N_8418);
nand U17398 (N_17398,N_6444,N_8725);
nor U17399 (N_17399,N_11637,N_6542);
or U17400 (N_17400,N_11638,N_10003);
nor U17401 (N_17401,N_8580,N_11708);
nand U17402 (N_17402,N_7883,N_9924);
nor U17403 (N_17403,N_11331,N_11941);
nand U17404 (N_17404,N_7477,N_11384);
xnor U17405 (N_17405,N_10167,N_6665);
and U17406 (N_17406,N_7065,N_7052);
xnor U17407 (N_17407,N_10517,N_8210);
nor U17408 (N_17408,N_9218,N_6436);
xnor U17409 (N_17409,N_6312,N_10195);
and U17410 (N_17410,N_11547,N_10843);
and U17411 (N_17411,N_8322,N_6461);
nor U17412 (N_17412,N_7465,N_7418);
xor U17413 (N_17413,N_6701,N_9596);
and U17414 (N_17414,N_10820,N_9254);
nor U17415 (N_17415,N_8462,N_10275);
xor U17416 (N_17416,N_9431,N_11579);
xor U17417 (N_17417,N_7511,N_11547);
or U17418 (N_17418,N_6409,N_9956);
nand U17419 (N_17419,N_6626,N_6792);
or U17420 (N_17420,N_11957,N_10458);
nor U17421 (N_17421,N_7738,N_8964);
nand U17422 (N_17422,N_8751,N_9790);
and U17423 (N_17423,N_9600,N_7318);
nor U17424 (N_17424,N_7048,N_7785);
nand U17425 (N_17425,N_8236,N_11394);
and U17426 (N_17426,N_8722,N_6653);
and U17427 (N_17427,N_6566,N_10827);
and U17428 (N_17428,N_10488,N_10621);
or U17429 (N_17429,N_9777,N_10358);
nand U17430 (N_17430,N_8928,N_11778);
nor U17431 (N_17431,N_6203,N_11291);
nand U17432 (N_17432,N_11150,N_8469);
and U17433 (N_17433,N_10962,N_11954);
nand U17434 (N_17434,N_11697,N_6423);
nor U17435 (N_17435,N_9947,N_8227);
or U17436 (N_17436,N_7246,N_10740);
xnor U17437 (N_17437,N_9751,N_7680);
or U17438 (N_17438,N_11308,N_8166);
nor U17439 (N_17439,N_9113,N_11321);
or U17440 (N_17440,N_9985,N_7629);
and U17441 (N_17441,N_8681,N_11702);
nand U17442 (N_17442,N_10543,N_11259);
xnor U17443 (N_17443,N_6877,N_9184);
or U17444 (N_17444,N_8137,N_7638);
nor U17445 (N_17445,N_7051,N_8793);
nand U17446 (N_17446,N_6766,N_7761);
and U17447 (N_17447,N_11603,N_8995);
xnor U17448 (N_17448,N_9391,N_9404);
nor U17449 (N_17449,N_11178,N_7758);
and U17450 (N_17450,N_6360,N_6835);
xnor U17451 (N_17451,N_8524,N_9000);
nand U17452 (N_17452,N_8231,N_7877);
and U17453 (N_17453,N_8586,N_6366);
nand U17454 (N_17454,N_8035,N_10946);
and U17455 (N_17455,N_9620,N_8660);
and U17456 (N_17456,N_7768,N_8300);
xor U17457 (N_17457,N_8419,N_9988);
and U17458 (N_17458,N_8950,N_11408);
or U17459 (N_17459,N_7154,N_9995);
and U17460 (N_17460,N_9466,N_11786);
or U17461 (N_17461,N_9911,N_6984);
nand U17462 (N_17462,N_9770,N_11444);
nor U17463 (N_17463,N_10574,N_10881);
and U17464 (N_17464,N_7201,N_6340);
or U17465 (N_17465,N_10527,N_9538);
xor U17466 (N_17466,N_9139,N_11588);
and U17467 (N_17467,N_11748,N_11225);
nor U17468 (N_17468,N_7752,N_10737);
xor U17469 (N_17469,N_9085,N_7918);
and U17470 (N_17470,N_8144,N_6501);
or U17471 (N_17471,N_9137,N_11091);
or U17472 (N_17472,N_6551,N_8385);
or U17473 (N_17473,N_9231,N_9187);
or U17474 (N_17474,N_9641,N_9963);
xnor U17475 (N_17475,N_11350,N_6883);
xnor U17476 (N_17476,N_8058,N_7789);
nand U17477 (N_17477,N_8569,N_7015);
or U17478 (N_17478,N_10130,N_9995);
and U17479 (N_17479,N_9799,N_9843);
nor U17480 (N_17480,N_6475,N_10409);
nand U17481 (N_17481,N_8134,N_10348);
nand U17482 (N_17482,N_8769,N_7784);
nand U17483 (N_17483,N_8720,N_11376);
nand U17484 (N_17484,N_8830,N_7867);
and U17485 (N_17485,N_10124,N_7354);
nand U17486 (N_17486,N_11305,N_8572);
and U17487 (N_17487,N_11910,N_6573);
xor U17488 (N_17488,N_10181,N_11485);
and U17489 (N_17489,N_10744,N_11361);
nand U17490 (N_17490,N_7947,N_11444);
and U17491 (N_17491,N_7915,N_6150);
or U17492 (N_17492,N_10345,N_6314);
nor U17493 (N_17493,N_8880,N_7489);
xor U17494 (N_17494,N_11709,N_7820);
xor U17495 (N_17495,N_11911,N_6454);
nand U17496 (N_17496,N_7076,N_6777);
and U17497 (N_17497,N_8384,N_7665);
and U17498 (N_17498,N_6870,N_9817);
and U17499 (N_17499,N_9903,N_9509);
nand U17500 (N_17500,N_6132,N_7410);
or U17501 (N_17501,N_11094,N_11780);
nand U17502 (N_17502,N_11116,N_8824);
nor U17503 (N_17503,N_8432,N_6741);
nand U17504 (N_17504,N_6701,N_8425);
xnor U17505 (N_17505,N_9018,N_6425);
or U17506 (N_17506,N_8547,N_9751);
nand U17507 (N_17507,N_6273,N_10723);
and U17508 (N_17508,N_9723,N_8607);
xnor U17509 (N_17509,N_8770,N_11840);
nor U17510 (N_17510,N_9240,N_11386);
or U17511 (N_17511,N_9479,N_10951);
or U17512 (N_17512,N_10359,N_9000);
and U17513 (N_17513,N_10223,N_6857);
xnor U17514 (N_17514,N_6433,N_7683);
xor U17515 (N_17515,N_8936,N_11670);
nand U17516 (N_17516,N_6493,N_6372);
nand U17517 (N_17517,N_9642,N_7174);
nand U17518 (N_17518,N_8313,N_10248);
nand U17519 (N_17519,N_9903,N_6192);
or U17520 (N_17520,N_9591,N_8418);
or U17521 (N_17521,N_6787,N_9237);
nand U17522 (N_17522,N_7674,N_8378);
nand U17523 (N_17523,N_7615,N_9891);
or U17524 (N_17524,N_9267,N_9858);
nor U17525 (N_17525,N_11813,N_11234);
and U17526 (N_17526,N_6826,N_7059);
xnor U17527 (N_17527,N_8147,N_11415);
xnor U17528 (N_17528,N_7690,N_8179);
and U17529 (N_17529,N_6774,N_10928);
or U17530 (N_17530,N_9853,N_11824);
xnor U17531 (N_17531,N_10065,N_8296);
or U17532 (N_17532,N_7596,N_9362);
nor U17533 (N_17533,N_6959,N_10583);
or U17534 (N_17534,N_8301,N_8048);
or U17535 (N_17535,N_6260,N_10421);
nand U17536 (N_17536,N_10959,N_10320);
xnor U17537 (N_17537,N_9303,N_10769);
or U17538 (N_17538,N_10683,N_6597);
nor U17539 (N_17539,N_8244,N_8694);
and U17540 (N_17540,N_11888,N_10302);
nor U17541 (N_17541,N_11796,N_9277);
xor U17542 (N_17542,N_10551,N_10897);
or U17543 (N_17543,N_6962,N_7789);
nor U17544 (N_17544,N_6309,N_8217);
nor U17545 (N_17545,N_6311,N_11790);
nor U17546 (N_17546,N_9501,N_7664);
nand U17547 (N_17547,N_11462,N_9798);
nand U17548 (N_17548,N_10644,N_7758);
nor U17549 (N_17549,N_7489,N_6334);
nand U17550 (N_17550,N_9320,N_11876);
xnor U17551 (N_17551,N_10975,N_11818);
or U17552 (N_17552,N_11385,N_6643);
nand U17553 (N_17553,N_6542,N_11472);
and U17554 (N_17554,N_11578,N_7319);
xnor U17555 (N_17555,N_6321,N_9739);
xnor U17556 (N_17556,N_9507,N_11144);
or U17557 (N_17557,N_6378,N_8352);
and U17558 (N_17558,N_6462,N_9835);
xnor U17559 (N_17559,N_7442,N_10325);
nand U17560 (N_17560,N_9186,N_7224);
xor U17561 (N_17561,N_6204,N_7260);
and U17562 (N_17562,N_8519,N_8833);
xnor U17563 (N_17563,N_11075,N_6047);
xnor U17564 (N_17564,N_7665,N_11730);
or U17565 (N_17565,N_11659,N_8732);
xnor U17566 (N_17566,N_6167,N_10029);
nand U17567 (N_17567,N_11929,N_10576);
or U17568 (N_17568,N_11641,N_11247);
xor U17569 (N_17569,N_9064,N_7020);
xnor U17570 (N_17570,N_10495,N_10773);
and U17571 (N_17571,N_11007,N_9227);
nor U17572 (N_17572,N_9235,N_6730);
and U17573 (N_17573,N_6076,N_6959);
or U17574 (N_17574,N_9182,N_11591);
nor U17575 (N_17575,N_11188,N_6050);
or U17576 (N_17576,N_6379,N_11716);
nand U17577 (N_17577,N_11296,N_10646);
nor U17578 (N_17578,N_6805,N_7925);
or U17579 (N_17579,N_8307,N_7330);
and U17580 (N_17580,N_10086,N_9855);
or U17581 (N_17581,N_9938,N_9215);
and U17582 (N_17582,N_6494,N_7002);
and U17583 (N_17583,N_8427,N_11409);
nor U17584 (N_17584,N_11301,N_6941);
or U17585 (N_17585,N_7995,N_6013);
nor U17586 (N_17586,N_11085,N_7566);
nor U17587 (N_17587,N_8637,N_10847);
xnor U17588 (N_17588,N_8958,N_9273);
or U17589 (N_17589,N_6450,N_11353);
nor U17590 (N_17590,N_11088,N_11239);
or U17591 (N_17591,N_6096,N_6605);
or U17592 (N_17592,N_11781,N_6257);
xnor U17593 (N_17593,N_8157,N_7190);
or U17594 (N_17594,N_10366,N_10351);
nor U17595 (N_17595,N_8831,N_10557);
nand U17596 (N_17596,N_11267,N_7913);
nor U17597 (N_17597,N_6838,N_7875);
xor U17598 (N_17598,N_10081,N_10229);
nand U17599 (N_17599,N_6214,N_10345);
xor U17600 (N_17600,N_9933,N_11681);
or U17601 (N_17601,N_8655,N_6789);
nand U17602 (N_17602,N_7110,N_9391);
or U17603 (N_17603,N_7395,N_6797);
nand U17604 (N_17604,N_7016,N_6682);
xor U17605 (N_17605,N_8781,N_10349);
xnor U17606 (N_17606,N_9062,N_10156);
and U17607 (N_17607,N_9510,N_8231);
nand U17608 (N_17608,N_11169,N_10127);
xnor U17609 (N_17609,N_8633,N_6360);
nor U17610 (N_17610,N_9961,N_6785);
or U17611 (N_17611,N_6386,N_7316);
and U17612 (N_17612,N_10748,N_6481);
nor U17613 (N_17613,N_11274,N_6591);
xnor U17614 (N_17614,N_6227,N_10184);
nand U17615 (N_17615,N_9510,N_6150);
nor U17616 (N_17616,N_7935,N_10773);
nor U17617 (N_17617,N_7835,N_9504);
nand U17618 (N_17618,N_6158,N_7969);
nand U17619 (N_17619,N_6545,N_6923);
nor U17620 (N_17620,N_8789,N_8537);
xor U17621 (N_17621,N_6053,N_8953);
and U17622 (N_17622,N_8606,N_11263);
nand U17623 (N_17623,N_6320,N_6391);
and U17624 (N_17624,N_10810,N_11518);
and U17625 (N_17625,N_10302,N_11543);
or U17626 (N_17626,N_8726,N_9322);
or U17627 (N_17627,N_7558,N_10831);
nor U17628 (N_17628,N_6023,N_7969);
nor U17629 (N_17629,N_7020,N_7260);
xor U17630 (N_17630,N_7780,N_11394);
nor U17631 (N_17631,N_7778,N_10094);
xor U17632 (N_17632,N_10954,N_10923);
and U17633 (N_17633,N_9146,N_8266);
or U17634 (N_17634,N_10323,N_6301);
nand U17635 (N_17635,N_9220,N_8349);
nor U17636 (N_17636,N_10713,N_7311);
xor U17637 (N_17637,N_7874,N_7841);
and U17638 (N_17638,N_6227,N_9239);
nor U17639 (N_17639,N_9146,N_10961);
nand U17640 (N_17640,N_10926,N_11320);
or U17641 (N_17641,N_8555,N_6241);
nand U17642 (N_17642,N_7208,N_8435);
nor U17643 (N_17643,N_7358,N_6838);
nand U17644 (N_17644,N_11252,N_6186);
xor U17645 (N_17645,N_6786,N_9090);
or U17646 (N_17646,N_9694,N_6820);
xnor U17647 (N_17647,N_9984,N_9348);
and U17648 (N_17648,N_11693,N_8232);
and U17649 (N_17649,N_8791,N_10550);
nand U17650 (N_17650,N_8143,N_6937);
nand U17651 (N_17651,N_11145,N_8659);
or U17652 (N_17652,N_8215,N_8256);
nor U17653 (N_17653,N_11591,N_9897);
or U17654 (N_17654,N_9776,N_11416);
xor U17655 (N_17655,N_10907,N_7491);
or U17656 (N_17656,N_8524,N_11009);
or U17657 (N_17657,N_10502,N_10746);
nand U17658 (N_17658,N_11742,N_11065);
or U17659 (N_17659,N_8917,N_6482);
or U17660 (N_17660,N_10129,N_10598);
or U17661 (N_17661,N_11703,N_11961);
xnor U17662 (N_17662,N_9421,N_9774);
and U17663 (N_17663,N_8059,N_6130);
and U17664 (N_17664,N_8567,N_9353);
xnor U17665 (N_17665,N_11819,N_9408);
xnor U17666 (N_17666,N_7736,N_9043);
nand U17667 (N_17667,N_10305,N_8444);
xnor U17668 (N_17668,N_7790,N_7266);
and U17669 (N_17669,N_8423,N_10912);
nand U17670 (N_17670,N_11383,N_6695);
nor U17671 (N_17671,N_10874,N_6165);
nor U17672 (N_17672,N_11100,N_9443);
xnor U17673 (N_17673,N_8047,N_6105);
and U17674 (N_17674,N_11457,N_8840);
or U17675 (N_17675,N_7108,N_7211);
or U17676 (N_17676,N_7368,N_8955);
nand U17677 (N_17677,N_6456,N_10233);
and U17678 (N_17678,N_9337,N_9420);
and U17679 (N_17679,N_8671,N_6662);
nor U17680 (N_17680,N_9400,N_11512);
nand U17681 (N_17681,N_7216,N_11006);
nor U17682 (N_17682,N_8320,N_11207);
or U17683 (N_17683,N_8031,N_9291);
and U17684 (N_17684,N_8567,N_10788);
and U17685 (N_17685,N_9666,N_11095);
nand U17686 (N_17686,N_11505,N_7614);
xor U17687 (N_17687,N_11227,N_9538);
or U17688 (N_17688,N_7015,N_10475);
or U17689 (N_17689,N_7552,N_10138);
xnor U17690 (N_17690,N_7084,N_7330);
nand U17691 (N_17691,N_11851,N_7116);
and U17692 (N_17692,N_11857,N_9159);
and U17693 (N_17693,N_6544,N_9099);
nor U17694 (N_17694,N_10550,N_10149);
and U17695 (N_17695,N_9010,N_11505);
nor U17696 (N_17696,N_8050,N_9201);
and U17697 (N_17697,N_8957,N_7403);
nand U17698 (N_17698,N_7567,N_11002);
nor U17699 (N_17699,N_8610,N_6501);
and U17700 (N_17700,N_6747,N_8838);
or U17701 (N_17701,N_7292,N_7720);
xor U17702 (N_17702,N_7091,N_7792);
nand U17703 (N_17703,N_11657,N_11132);
or U17704 (N_17704,N_11441,N_8379);
nand U17705 (N_17705,N_8471,N_10323);
and U17706 (N_17706,N_8626,N_6381);
or U17707 (N_17707,N_11370,N_11991);
xnor U17708 (N_17708,N_9415,N_11679);
nand U17709 (N_17709,N_9998,N_6732);
xnor U17710 (N_17710,N_11404,N_8517);
nor U17711 (N_17711,N_11715,N_10821);
nand U17712 (N_17712,N_6638,N_11693);
xnor U17713 (N_17713,N_9899,N_8428);
xor U17714 (N_17714,N_9744,N_6802);
nor U17715 (N_17715,N_7374,N_9567);
and U17716 (N_17716,N_7205,N_6310);
xnor U17717 (N_17717,N_11100,N_6991);
and U17718 (N_17718,N_6835,N_9580);
xor U17719 (N_17719,N_9584,N_10548);
or U17720 (N_17720,N_9116,N_8295);
or U17721 (N_17721,N_10055,N_10794);
and U17722 (N_17722,N_7738,N_6859);
nand U17723 (N_17723,N_9638,N_11405);
xor U17724 (N_17724,N_10669,N_9716);
or U17725 (N_17725,N_7165,N_6876);
or U17726 (N_17726,N_8506,N_11074);
nand U17727 (N_17727,N_8582,N_11865);
xor U17728 (N_17728,N_9984,N_6862);
nor U17729 (N_17729,N_11677,N_6438);
nand U17730 (N_17730,N_6317,N_9829);
nand U17731 (N_17731,N_7846,N_11513);
nand U17732 (N_17732,N_11585,N_6579);
nor U17733 (N_17733,N_10778,N_9489);
xor U17734 (N_17734,N_7018,N_9661);
nand U17735 (N_17735,N_6262,N_6476);
nor U17736 (N_17736,N_10474,N_9364);
or U17737 (N_17737,N_8595,N_10232);
nand U17738 (N_17738,N_6295,N_10899);
nor U17739 (N_17739,N_10353,N_7088);
nor U17740 (N_17740,N_10273,N_6421);
xnor U17741 (N_17741,N_9663,N_10279);
or U17742 (N_17742,N_10734,N_7262);
and U17743 (N_17743,N_8050,N_6203);
or U17744 (N_17744,N_8532,N_7159);
xor U17745 (N_17745,N_8540,N_6064);
and U17746 (N_17746,N_9969,N_7928);
nand U17747 (N_17747,N_7165,N_9266);
xnor U17748 (N_17748,N_9758,N_11264);
nand U17749 (N_17749,N_8570,N_7470);
xnor U17750 (N_17750,N_10212,N_7724);
xnor U17751 (N_17751,N_11740,N_6435);
nor U17752 (N_17752,N_6189,N_11357);
xnor U17753 (N_17753,N_8631,N_9133);
nor U17754 (N_17754,N_8619,N_9454);
nor U17755 (N_17755,N_10104,N_10047);
xor U17756 (N_17756,N_8814,N_11750);
xor U17757 (N_17757,N_11770,N_7361);
nor U17758 (N_17758,N_9592,N_6661);
and U17759 (N_17759,N_11891,N_9641);
and U17760 (N_17760,N_9957,N_8956);
nor U17761 (N_17761,N_11835,N_11260);
nand U17762 (N_17762,N_6192,N_6722);
and U17763 (N_17763,N_8412,N_8268);
and U17764 (N_17764,N_10820,N_6196);
nand U17765 (N_17765,N_7576,N_9101);
nand U17766 (N_17766,N_8820,N_9182);
or U17767 (N_17767,N_8590,N_6294);
and U17768 (N_17768,N_10815,N_7070);
xor U17769 (N_17769,N_9676,N_9482);
nor U17770 (N_17770,N_6759,N_7739);
or U17771 (N_17771,N_6783,N_7933);
and U17772 (N_17772,N_8368,N_7540);
and U17773 (N_17773,N_9248,N_8962);
or U17774 (N_17774,N_8086,N_8115);
and U17775 (N_17775,N_9175,N_9152);
nor U17776 (N_17776,N_11807,N_11671);
and U17777 (N_17777,N_11106,N_11042);
or U17778 (N_17778,N_6444,N_7266);
nor U17779 (N_17779,N_6815,N_8829);
nand U17780 (N_17780,N_9054,N_10643);
or U17781 (N_17781,N_6503,N_11881);
or U17782 (N_17782,N_10104,N_9591);
nand U17783 (N_17783,N_7711,N_10617);
xnor U17784 (N_17784,N_11445,N_7310);
nor U17785 (N_17785,N_9632,N_8337);
and U17786 (N_17786,N_10624,N_10520);
or U17787 (N_17787,N_11250,N_10927);
and U17788 (N_17788,N_10768,N_10446);
xor U17789 (N_17789,N_11945,N_6283);
or U17790 (N_17790,N_8416,N_10544);
nand U17791 (N_17791,N_8211,N_6427);
nor U17792 (N_17792,N_7836,N_7192);
xnor U17793 (N_17793,N_9554,N_9827);
and U17794 (N_17794,N_8596,N_7613);
or U17795 (N_17795,N_11191,N_7316);
and U17796 (N_17796,N_11769,N_8865);
or U17797 (N_17797,N_6179,N_7693);
or U17798 (N_17798,N_6782,N_11807);
and U17799 (N_17799,N_6148,N_11768);
and U17800 (N_17800,N_6863,N_6160);
or U17801 (N_17801,N_8705,N_8361);
and U17802 (N_17802,N_11074,N_9154);
and U17803 (N_17803,N_8369,N_7172);
nor U17804 (N_17804,N_9397,N_8226);
or U17805 (N_17805,N_9220,N_11006);
and U17806 (N_17806,N_8199,N_7983);
or U17807 (N_17807,N_9060,N_8947);
and U17808 (N_17808,N_10389,N_6649);
or U17809 (N_17809,N_10508,N_11224);
xor U17810 (N_17810,N_7130,N_11877);
and U17811 (N_17811,N_11025,N_6106);
nor U17812 (N_17812,N_8178,N_6462);
or U17813 (N_17813,N_6686,N_11488);
nor U17814 (N_17814,N_7144,N_10066);
or U17815 (N_17815,N_8229,N_10293);
and U17816 (N_17816,N_9180,N_8270);
and U17817 (N_17817,N_9905,N_7048);
xnor U17818 (N_17818,N_9383,N_8055);
or U17819 (N_17819,N_11170,N_6064);
nand U17820 (N_17820,N_8563,N_8954);
nor U17821 (N_17821,N_8230,N_10866);
or U17822 (N_17822,N_10387,N_9679);
or U17823 (N_17823,N_6351,N_6017);
nand U17824 (N_17824,N_10395,N_11881);
nand U17825 (N_17825,N_9650,N_8013);
nor U17826 (N_17826,N_10074,N_6403);
or U17827 (N_17827,N_8496,N_7505);
xor U17828 (N_17828,N_8591,N_8977);
and U17829 (N_17829,N_11230,N_10683);
nand U17830 (N_17830,N_9270,N_9755);
and U17831 (N_17831,N_8546,N_8091);
xor U17832 (N_17832,N_6053,N_7097);
or U17833 (N_17833,N_8899,N_10047);
xor U17834 (N_17834,N_8735,N_9985);
nor U17835 (N_17835,N_6599,N_6805);
nand U17836 (N_17836,N_8052,N_7973);
and U17837 (N_17837,N_9890,N_7882);
xnor U17838 (N_17838,N_7657,N_6117);
and U17839 (N_17839,N_9724,N_7908);
nand U17840 (N_17840,N_6883,N_8095);
xnor U17841 (N_17841,N_8704,N_11093);
or U17842 (N_17842,N_8686,N_8293);
nand U17843 (N_17843,N_10580,N_10367);
nor U17844 (N_17844,N_9865,N_9268);
xor U17845 (N_17845,N_8681,N_6103);
nor U17846 (N_17846,N_7089,N_6491);
nand U17847 (N_17847,N_6041,N_7117);
nor U17848 (N_17848,N_7920,N_8504);
and U17849 (N_17849,N_6840,N_11041);
and U17850 (N_17850,N_7471,N_7859);
and U17851 (N_17851,N_10813,N_10197);
xor U17852 (N_17852,N_8981,N_7475);
nor U17853 (N_17853,N_8280,N_10855);
xor U17854 (N_17854,N_9828,N_9569);
nor U17855 (N_17855,N_8339,N_7395);
xnor U17856 (N_17856,N_9581,N_6128);
nor U17857 (N_17857,N_7764,N_6789);
or U17858 (N_17858,N_8421,N_6844);
and U17859 (N_17859,N_9046,N_8851);
or U17860 (N_17860,N_9300,N_8512);
nand U17861 (N_17861,N_8171,N_11168);
xnor U17862 (N_17862,N_10462,N_8139);
xor U17863 (N_17863,N_11116,N_10709);
nand U17864 (N_17864,N_8815,N_9897);
and U17865 (N_17865,N_7174,N_8891);
xnor U17866 (N_17866,N_11789,N_9413);
nand U17867 (N_17867,N_10729,N_7381);
and U17868 (N_17868,N_8155,N_8442);
and U17869 (N_17869,N_11051,N_7873);
or U17870 (N_17870,N_11217,N_11966);
xor U17871 (N_17871,N_7711,N_8113);
or U17872 (N_17872,N_11516,N_10248);
and U17873 (N_17873,N_11445,N_10622);
xor U17874 (N_17874,N_8108,N_7417);
nor U17875 (N_17875,N_6239,N_6055);
nor U17876 (N_17876,N_11229,N_7573);
or U17877 (N_17877,N_9668,N_10514);
and U17878 (N_17878,N_11794,N_7463);
or U17879 (N_17879,N_11665,N_11977);
nand U17880 (N_17880,N_10543,N_9931);
or U17881 (N_17881,N_9636,N_8554);
and U17882 (N_17882,N_10935,N_8539);
nor U17883 (N_17883,N_6754,N_9992);
or U17884 (N_17884,N_11409,N_8357);
xnor U17885 (N_17885,N_11673,N_8783);
nand U17886 (N_17886,N_7905,N_10335);
xor U17887 (N_17887,N_7064,N_10686);
xor U17888 (N_17888,N_9351,N_6962);
xor U17889 (N_17889,N_7076,N_9497);
nand U17890 (N_17890,N_9319,N_6708);
nor U17891 (N_17891,N_8705,N_7417);
nand U17892 (N_17892,N_8761,N_7297);
nor U17893 (N_17893,N_8411,N_6145);
xnor U17894 (N_17894,N_11603,N_10303);
or U17895 (N_17895,N_6732,N_7391);
or U17896 (N_17896,N_7912,N_7888);
xor U17897 (N_17897,N_8459,N_8155);
nor U17898 (N_17898,N_8364,N_10796);
xor U17899 (N_17899,N_10935,N_8425);
or U17900 (N_17900,N_8826,N_8216);
nor U17901 (N_17901,N_7177,N_6619);
nor U17902 (N_17902,N_8210,N_11995);
xnor U17903 (N_17903,N_7788,N_8465);
nor U17904 (N_17904,N_6815,N_7692);
xnor U17905 (N_17905,N_6974,N_6414);
nand U17906 (N_17906,N_10122,N_6202);
nor U17907 (N_17907,N_9948,N_6719);
or U17908 (N_17908,N_7680,N_11359);
or U17909 (N_17909,N_9792,N_8741);
nor U17910 (N_17910,N_6921,N_11435);
nor U17911 (N_17911,N_6922,N_11218);
nor U17912 (N_17912,N_6499,N_11329);
or U17913 (N_17913,N_8031,N_8268);
nand U17914 (N_17914,N_11532,N_6406);
and U17915 (N_17915,N_11919,N_6198);
nand U17916 (N_17916,N_9161,N_10364);
xnor U17917 (N_17917,N_11656,N_6555);
and U17918 (N_17918,N_9355,N_7105);
nand U17919 (N_17919,N_7712,N_11466);
nand U17920 (N_17920,N_6607,N_9212);
or U17921 (N_17921,N_11171,N_10027);
xor U17922 (N_17922,N_7977,N_8032);
nand U17923 (N_17923,N_8391,N_8304);
and U17924 (N_17924,N_7828,N_11889);
and U17925 (N_17925,N_8728,N_10088);
nor U17926 (N_17926,N_11820,N_7823);
xor U17927 (N_17927,N_11765,N_7011);
or U17928 (N_17928,N_6907,N_9648);
nand U17929 (N_17929,N_10850,N_6884);
or U17930 (N_17930,N_11431,N_10970);
and U17931 (N_17931,N_11891,N_6103);
or U17932 (N_17932,N_7209,N_6836);
xor U17933 (N_17933,N_6881,N_7671);
nand U17934 (N_17934,N_6882,N_7907);
or U17935 (N_17935,N_6961,N_9088);
nor U17936 (N_17936,N_7995,N_9223);
or U17937 (N_17937,N_8729,N_8403);
or U17938 (N_17938,N_6723,N_8450);
nand U17939 (N_17939,N_7417,N_9920);
nor U17940 (N_17940,N_8936,N_9011);
nor U17941 (N_17941,N_6817,N_7708);
nand U17942 (N_17942,N_9368,N_7700);
and U17943 (N_17943,N_6987,N_8953);
nand U17944 (N_17944,N_7729,N_10653);
and U17945 (N_17945,N_7436,N_11954);
xnor U17946 (N_17946,N_7628,N_10887);
xor U17947 (N_17947,N_10695,N_6449);
or U17948 (N_17948,N_7198,N_11274);
xnor U17949 (N_17949,N_11224,N_8386);
nor U17950 (N_17950,N_10734,N_9402);
nand U17951 (N_17951,N_8421,N_7003);
and U17952 (N_17952,N_6570,N_6207);
xnor U17953 (N_17953,N_9371,N_7862);
and U17954 (N_17954,N_10943,N_11422);
nor U17955 (N_17955,N_9500,N_9490);
nor U17956 (N_17956,N_11418,N_8436);
nand U17957 (N_17957,N_7612,N_8222);
and U17958 (N_17958,N_9825,N_7917);
and U17959 (N_17959,N_11065,N_8576);
nor U17960 (N_17960,N_8901,N_8588);
nor U17961 (N_17961,N_6230,N_6758);
nand U17962 (N_17962,N_10127,N_11857);
or U17963 (N_17963,N_7085,N_8788);
xor U17964 (N_17964,N_7938,N_11086);
or U17965 (N_17965,N_10289,N_7156);
nor U17966 (N_17966,N_6326,N_8370);
nand U17967 (N_17967,N_9193,N_7911);
nor U17968 (N_17968,N_6154,N_7223);
nand U17969 (N_17969,N_7787,N_8016);
nand U17970 (N_17970,N_9839,N_10003);
nand U17971 (N_17971,N_9831,N_8193);
and U17972 (N_17972,N_6833,N_10597);
nand U17973 (N_17973,N_11057,N_10085);
nand U17974 (N_17974,N_6269,N_8619);
nand U17975 (N_17975,N_8500,N_8990);
xor U17976 (N_17976,N_7546,N_6515);
nand U17977 (N_17977,N_9681,N_9425);
nor U17978 (N_17978,N_6402,N_8470);
and U17979 (N_17979,N_9599,N_6626);
or U17980 (N_17980,N_7708,N_8018);
nand U17981 (N_17981,N_11203,N_6093);
xor U17982 (N_17982,N_11591,N_10221);
xnor U17983 (N_17983,N_9035,N_8777);
nand U17984 (N_17984,N_9439,N_9400);
or U17985 (N_17985,N_10721,N_6939);
and U17986 (N_17986,N_9096,N_7872);
nand U17987 (N_17987,N_7111,N_11988);
xnor U17988 (N_17988,N_9429,N_8356);
nand U17989 (N_17989,N_8936,N_11616);
nand U17990 (N_17990,N_11375,N_8801);
nand U17991 (N_17991,N_6639,N_8930);
nand U17992 (N_17992,N_8171,N_9490);
or U17993 (N_17993,N_10049,N_7552);
nand U17994 (N_17994,N_9981,N_9134);
xor U17995 (N_17995,N_6310,N_10836);
or U17996 (N_17996,N_11882,N_9985);
or U17997 (N_17997,N_9799,N_7983);
and U17998 (N_17998,N_6205,N_9625);
and U17999 (N_17999,N_9422,N_7918);
nand U18000 (N_18000,N_14306,N_14988);
xor U18001 (N_18001,N_17776,N_16624);
and U18002 (N_18002,N_14882,N_15947);
or U18003 (N_18003,N_14608,N_15301);
nand U18004 (N_18004,N_17654,N_16657);
and U18005 (N_18005,N_15487,N_14137);
xnor U18006 (N_18006,N_17923,N_17289);
nand U18007 (N_18007,N_16201,N_12024);
and U18008 (N_18008,N_13535,N_16332);
xor U18009 (N_18009,N_13215,N_17881);
nor U18010 (N_18010,N_17630,N_14980);
nand U18011 (N_18011,N_13401,N_13434);
nand U18012 (N_18012,N_13039,N_15883);
and U18013 (N_18013,N_16252,N_12645);
nand U18014 (N_18014,N_13157,N_13399);
and U18015 (N_18015,N_14849,N_17047);
nor U18016 (N_18016,N_16777,N_12956);
nand U18017 (N_18017,N_14714,N_17804);
nand U18018 (N_18018,N_15967,N_15779);
and U18019 (N_18019,N_13185,N_17502);
xnor U18020 (N_18020,N_15662,N_13885);
or U18021 (N_18021,N_14694,N_17615);
xnor U18022 (N_18022,N_12705,N_13833);
xor U18023 (N_18023,N_16858,N_13330);
xnor U18024 (N_18024,N_14405,N_13411);
and U18025 (N_18025,N_13000,N_15655);
xor U18026 (N_18026,N_14266,N_14625);
xnor U18027 (N_18027,N_17256,N_13934);
nand U18028 (N_18028,N_15636,N_16779);
nand U18029 (N_18029,N_12595,N_12665);
nand U18030 (N_18030,N_14635,N_13114);
or U18031 (N_18031,N_13072,N_16143);
xnor U18032 (N_18032,N_13458,N_14052);
nand U18033 (N_18033,N_12409,N_12265);
and U18034 (N_18034,N_13881,N_16012);
nand U18035 (N_18035,N_17141,N_15252);
nand U18036 (N_18036,N_16043,N_16129);
and U18037 (N_18037,N_12742,N_12385);
nand U18038 (N_18038,N_17532,N_15019);
nor U18039 (N_18039,N_15821,N_16786);
nand U18040 (N_18040,N_17833,N_17544);
and U18041 (N_18041,N_16602,N_17810);
xor U18042 (N_18042,N_16381,N_13971);
xor U18043 (N_18043,N_14834,N_17943);
nor U18044 (N_18044,N_13802,N_15095);
xor U18045 (N_18045,N_12816,N_13266);
or U18046 (N_18046,N_12515,N_15932);
or U18047 (N_18047,N_12890,N_15812);
and U18048 (N_18048,N_17004,N_15331);
nand U18049 (N_18049,N_15530,N_16555);
or U18050 (N_18050,N_14931,N_13619);
nor U18051 (N_18051,N_13291,N_14339);
or U18052 (N_18052,N_14343,N_12969);
nor U18053 (N_18053,N_17262,N_15341);
nand U18054 (N_18054,N_16476,N_17494);
nor U18055 (N_18055,N_12843,N_14921);
xor U18056 (N_18056,N_13969,N_13181);
nand U18057 (N_18057,N_16666,N_16000);
or U18058 (N_18058,N_15234,N_16185);
or U18059 (N_18059,N_16656,N_12579);
and U18060 (N_18060,N_16312,N_13436);
nand U18061 (N_18061,N_17671,N_14582);
xnor U18062 (N_18062,N_15075,N_15406);
and U18063 (N_18063,N_14830,N_14402);
xor U18064 (N_18064,N_15783,N_12247);
xor U18065 (N_18065,N_17665,N_14518);
or U18066 (N_18066,N_14406,N_14575);
and U18067 (N_18067,N_13255,N_15585);
and U18068 (N_18068,N_16058,N_15877);
nor U18069 (N_18069,N_15300,N_14043);
nor U18070 (N_18070,N_17296,N_12818);
and U18071 (N_18071,N_16735,N_12797);
and U18072 (N_18072,N_13310,N_12317);
nor U18073 (N_18073,N_15933,N_15140);
nand U18074 (N_18074,N_17829,N_13653);
xor U18075 (N_18075,N_17041,N_15448);
nand U18076 (N_18076,N_14507,N_16340);
nor U18077 (N_18077,N_14887,N_13496);
and U18078 (N_18078,N_13263,N_15759);
xor U18079 (N_18079,N_13205,N_15880);
xor U18080 (N_18080,N_15789,N_13575);
nor U18081 (N_18081,N_15419,N_15318);
xor U18082 (N_18082,N_13128,N_16292);
nor U18083 (N_18083,N_13849,N_12751);
nor U18084 (N_18084,N_14421,N_15244);
xor U18085 (N_18085,N_12625,N_15383);
nand U18086 (N_18086,N_14163,N_12292);
and U18087 (N_18087,N_12219,N_17099);
xnor U18088 (N_18088,N_15981,N_15553);
or U18089 (N_18089,N_13447,N_17164);
xor U18090 (N_18090,N_16342,N_12239);
nand U18091 (N_18091,N_17990,N_16220);
nor U18092 (N_18092,N_15510,N_13736);
or U18093 (N_18093,N_13369,N_16133);
or U18094 (N_18094,N_12055,N_16648);
xnor U18095 (N_18095,N_13970,N_15389);
nor U18096 (N_18096,N_12868,N_15181);
nand U18097 (N_18097,N_12531,N_16331);
or U18098 (N_18098,N_15692,N_15698);
or U18099 (N_18099,N_14065,N_13499);
or U18100 (N_18100,N_17126,N_13754);
nor U18101 (N_18101,N_12025,N_12944);
xnor U18102 (N_18102,N_12837,N_14783);
nand U18103 (N_18103,N_17799,N_15020);
or U18104 (N_18104,N_16447,N_14764);
or U18105 (N_18105,N_17701,N_16053);
nand U18106 (N_18106,N_16251,N_16887);
and U18107 (N_18107,N_14657,N_17343);
or U18108 (N_18108,N_12841,N_17015);
or U18109 (N_18109,N_16830,N_16927);
or U18110 (N_18110,N_12270,N_13835);
nor U18111 (N_18111,N_15513,N_17127);
nor U18112 (N_18112,N_14915,N_15342);
and U18113 (N_18113,N_14804,N_16788);
and U18114 (N_18114,N_14621,N_14674);
and U18115 (N_18115,N_17095,N_14152);
nor U18116 (N_18116,N_12507,N_13875);
nand U18117 (N_18117,N_15423,N_16209);
or U18118 (N_18118,N_13895,N_17619);
or U18119 (N_18119,N_14205,N_13916);
or U18120 (N_18120,N_13356,N_12176);
and U18121 (N_18121,N_17559,N_12570);
xnor U18122 (N_18122,N_14789,N_16806);
nor U18123 (N_18123,N_17321,N_16967);
and U18124 (N_18124,N_13946,N_12585);
and U18125 (N_18125,N_12903,N_16695);
nand U18126 (N_18126,N_17857,N_15519);
or U18127 (N_18127,N_16245,N_17310);
and U18128 (N_18128,N_17794,N_17113);
nand U18129 (N_18129,N_14226,N_12527);
nand U18130 (N_18130,N_17979,N_13697);
and U18131 (N_18131,N_12351,N_15505);
and U18132 (N_18132,N_15474,N_17678);
xor U18133 (N_18133,N_12202,N_17094);
nand U18134 (N_18134,N_15078,N_16552);
nor U18135 (N_18135,N_17846,N_14824);
nor U18136 (N_18136,N_15337,N_13710);
nand U18137 (N_18137,N_13329,N_15567);
and U18138 (N_18138,N_16075,N_13410);
and U18139 (N_18139,N_14530,N_13592);
xnor U18140 (N_18140,N_13957,N_13612);
and U18141 (N_18141,N_15617,N_15669);
and U18142 (N_18142,N_12426,N_15228);
and U18143 (N_18143,N_14650,N_14842);
or U18144 (N_18144,N_14470,N_17854);
xor U18145 (N_18145,N_12183,N_13096);
or U18146 (N_18146,N_13995,N_15881);
nand U18147 (N_18147,N_13374,N_17426);
nand U18148 (N_18148,N_17398,N_13509);
or U18149 (N_18149,N_16671,N_12454);
nor U18150 (N_18150,N_13587,N_15499);
nand U18151 (N_18151,N_17009,N_13122);
nor U18152 (N_18152,N_15674,N_15472);
xor U18153 (N_18153,N_16847,N_17153);
nor U18154 (N_18154,N_17301,N_16029);
xor U18155 (N_18155,N_14498,N_17664);
nor U18156 (N_18156,N_14062,N_12557);
and U18157 (N_18157,N_13088,N_17805);
and U18158 (N_18158,N_12178,N_13649);
nor U18159 (N_18159,N_16509,N_14550);
nand U18160 (N_18160,N_15230,N_13209);
nor U18161 (N_18161,N_12869,N_13170);
nand U18162 (N_18162,N_12282,N_16047);
nor U18163 (N_18163,N_17403,N_15801);
and U18164 (N_18164,N_12235,N_13270);
xnor U18165 (N_18165,N_14893,N_16274);
nor U18166 (N_18166,N_14861,N_13467);
nor U18167 (N_18167,N_12614,N_16931);
nand U18168 (N_18168,N_15564,N_12408);
nor U18169 (N_18169,N_17516,N_17602);
nor U18170 (N_18170,N_12510,N_12330);
xor U18171 (N_18171,N_13904,N_15722);
xor U18172 (N_18172,N_15885,N_15670);
and U18173 (N_18173,N_14543,N_15964);
xnor U18174 (N_18174,N_17035,N_13493);
or U18175 (N_18175,N_13968,N_17467);
nor U18176 (N_18176,N_12143,N_12702);
nor U18177 (N_18177,N_15046,N_15882);
and U18178 (N_18178,N_16427,N_14314);
or U18179 (N_18179,N_17731,N_13917);
xnor U18180 (N_18180,N_12878,N_17937);
nor U18181 (N_18181,N_16780,N_14353);
or U18182 (N_18182,N_15468,N_12714);
nand U18183 (N_18183,N_15540,N_13191);
nand U18184 (N_18184,N_16463,N_15130);
and U18185 (N_18185,N_13562,N_12783);
nand U18186 (N_18186,N_13817,N_16156);
nor U18187 (N_18187,N_14207,N_12602);
nor U18188 (N_18188,N_12785,N_13857);
nand U18189 (N_18189,N_16782,N_14193);
xor U18190 (N_18190,N_13732,N_17878);
or U18191 (N_18191,N_17220,N_13613);
nor U18192 (N_18192,N_13139,N_15041);
xnor U18193 (N_18193,N_13309,N_17484);
and U18194 (N_18194,N_15570,N_15476);
nand U18195 (N_18195,N_13184,N_16392);
nor U18196 (N_18196,N_13452,N_15339);
nand U18197 (N_18197,N_14217,N_14559);
xnor U18198 (N_18198,N_13507,N_17160);
and U18199 (N_18199,N_12889,N_13197);
nor U18200 (N_18200,N_17292,N_13002);
or U18201 (N_18201,N_14671,N_15489);
nor U18202 (N_18202,N_12638,N_15725);
nand U18203 (N_18203,N_15566,N_14091);
xnor U18204 (N_18204,N_14620,N_13664);
nor U18205 (N_18205,N_14110,N_17775);
and U18206 (N_18206,N_12000,N_13961);
nor U18207 (N_18207,N_17003,N_16679);
nand U18208 (N_18208,N_17255,N_17211);
and U18209 (N_18209,N_13034,N_16686);
and U18210 (N_18210,N_13005,N_16682);
nand U18211 (N_18211,N_14715,N_13015);
nand U18212 (N_18212,N_13195,N_15271);
nor U18213 (N_18213,N_14593,N_16890);
xnor U18214 (N_18214,N_14135,N_14221);
or U18215 (N_18215,N_14612,N_13728);
nor U18216 (N_18216,N_14547,N_12499);
or U18217 (N_18217,N_15755,N_13520);
or U18218 (N_18218,N_15637,N_16396);
or U18219 (N_18219,N_13094,N_15621);
and U18220 (N_18220,N_17515,N_16365);
and U18221 (N_18221,N_15833,N_13077);
nor U18222 (N_18222,N_12363,N_13229);
or U18223 (N_18223,N_15641,N_17563);
nor U18224 (N_18224,N_14422,N_15913);
or U18225 (N_18225,N_16601,N_12787);
and U18226 (N_18226,N_12489,N_17493);
nand U18227 (N_18227,N_13823,N_17155);
nor U18228 (N_18228,N_17750,N_12471);
or U18229 (N_18229,N_13661,N_16044);
nand U18230 (N_18230,N_13379,N_12850);
or U18231 (N_18231,N_17722,N_16275);
nor U18232 (N_18232,N_13611,N_15622);
nand U18233 (N_18233,N_16878,N_13407);
and U18234 (N_18234,N_16165,N_12600);
or U18235 (N_18235,N_13668,N_17176);
xor U18236 (N_18236,N_17920,N_16369);
nor U18237 (N_18237,N_17295,N_16234);
nand U18238 (N_18238,N_13757,N_15296);
and U18239 (N_18239,N_14943,N_13759);
nand U18240 (N_18240,N_14648,N_13599);
and U18241 (N_18241,N_15183,N_13589);
nor U18242 (N_18242,N_16716,N_15104);
or U18243 (N_18243,N_15950,N_16320);
or U18244 (N_18244,N_14642,N_15646);
xor U18245 (N_18245,N_15490,N_17019);
or U18246 (N_18246,N_17699,N_14699);
and U18247 (N_18247,N_17062,N_14799);
nor U18248 (N_18248,N_13361,N_14377);
nand U18249 (N_18249,N_16457,N_14454);
nand U18250 (N_18250,N_16354,N_14555);
or U18251 (N_18251,N_13483,N_14145);
nand U18252 (N_18252,N_17567,N_12684);
or U18253 (N_18253,N_12578,N_16981);
nor U18254 (N_18254,N_13800,N_16805);
or U18255 (N_18255,N_13083,N_16709);
and U18256 (N_18256,N_12214,N_16142);
or U18257 (N_18257,N_16702,N_16266);
xnor U18258 (N_18258,N_16092,N_17243);
or U18259 (N_18259,N_12781,N_15015);
or U18260 (N_18260,N_13519,N_15809);
and U18261 (N_18261,N_15189,N_17347);
and U18262 (N_18262,N_14428,N_16464);
nor U18263 (N_18263,N_15278,N_14430);
and U18264 (N_18264,N_16431,N_15410);
nor U18265 (N_18265,N_14576,N_13280);
or U18266 (N_18266,N_15713,N_12768);
xor U18267 (N_18267,N_17632,N_16579);
nor U18268 (N_18268,N_14203,N_14060);
or U18269 (N_18269,N_16647,N_13024);
nand U18270 (N_18270,N_16995,N_13773);
nor U18271 (N_18271,N_13684,N_17133);
and U18272 (N_18272,N_17589,N_12793);
nor U18273 (N_18273,N_12070,N_12554);
or U18274 (N_18274,N_13156,N_12607);
nor U18275 (N_18275,N_12336,N_15853);
nor U18276 (N_18276,N_17717,N_16717);
nor U18277 (N_18277,N_15627,N_13045);
or U18278 (N_18278,N_16045,N_13030);
or U18279 (N_18279,N_16963,N_17235);
xnor U18280 (N_18280,N_14464,N_17709);
nand U18281 (N_18281,N_15257,N_15691);
or U18282 (N_18282,N_16619,N_16934);
nand U18283 (N_18283,N_17065,N_13975);
xnor U18284 (N_18284,N_17172,N_17887);
xor U18285 (N_18285,N_12367,N_17088);
and U18286 (N_18286,N_12035,N_15065);
nand U18287 (N_18287,N_17459,N_12014);
and U18288 (N_18288,N_16242,N_14218);
nor U18289 (N_18289,N_12445,N_12998);
xnor U18290 (N_18290,N_13941,N_17600);
or U18291 (N_18291,N_15576,N_12713);
nor U18292 (N_18292,N_15224,N_16147);
nand U18293 (N_18293,N_14199,N_13689);
xor U18294 (N_18294,N_14118,N_15836);
nand U18295 (N_18295,N_17784,N_15386);
and U18296 (N_18296,N_17227,N_13782);
xor U18297 (N_18297,N_15162,N_12318);
xnor U18298 (N_18298,N_15479,N_15477);
or U18299 (N_18299,N_13672,N_12370);
and U18300 (N_18300,N_16168,N_14668);
nand U18301 (N_18301,N_14165,N_15437);
and U18302 (N_18302,N_12468,N_14971);
xnor U18303 (N_18303,N_16363,N_12011);
nand U18304 (N_18304,N_16290,N_13796);
or U18305 (N_18305,N_15592,N_12240);
and U18306 (N_18306,N_15105,N_13299);
nor U18307 (N_18307,N_15049,N_14248);
xnor U18308 (N_18308,N_13593,N_12474);
nand U18309 (N_18309,N_13490,N_12572);
nand U18310 (N_18310,N_14829,N_13443);
nand U18311 (N_18311,N_17638,N_16529);
nor U18312 (N_18312,N_12970,N_12854);
nor U18313 (N_18313,N_17861,N_17434);
nor U18314 (N_18314,N_16672,N_13918);
xor U18315 (N_18315,N_12676,N_17033);
nand U18316 (N_18316,N_12865,N_14926);
and U18317 (N_18317,N_17233,N_15732);
xor U18318 (N_18318,N_15748,N_12796);
nor U18319 (N_18319,N_16102,N_13186);
xnor U18320 (N_18320,N_16958,N_12126);
nor U18321 (N_18321,N_12509,N_14275);
nand U18322 (N_18322,N_14795,N_12194);
nor U18323 (N_18323,N_14775,N_15220);
xor U18324 (N_18324,N_12144,N_14153);
nor U18325 (N_18325,N_17852,N_16177);
xor U18326 (N_18326,N_14144,N_17476);
xor U18327 (N_18327,N_14952,N_15741);
or U18328 (N_18328,N_12091,N_15599);
xnor U18329 (N_18329,N_13175,N_12184);
xor U18330 (N_18330,N_13964,N_14227);
nor U18331 (N_18331,N_14182,N_14189);
and U18332 (N_18332,N_14916,N_13258);
xor U18333 (N_18333,N_14756,N_16336);
or U18334 (N_18334,N_14810,N_12932);
xor U18335 (N_18335,N_12897,N_16341);
and U18336 (N_18336,N_17478,N_14607);
nand U18337 (N_18337,N_16415,N_13897);
nor U18338 (N_18338,N_14667,N_15360);
xnor U18339 (N_18339,N_17596,N_12166);
xnor U18340 (N_18340,N_17116,N_15822);
and U18341 (N_18341,N_14661,N_15209);
nand U18342 (N_18342,N_13297,N_16364);
or U18343 (N_18343,N_15335,N_13498);
and U18344 (N_18344,N_17734,N_13482);
or U18345 (N_18345,N_15849,N_12963);
xor U18346 (N_18346,N_15940,N_13358);
and U18347 (N_18347,N_17159,N_14776);
xor U18348 (N_18348,N_15525,N_14603);
xnor U18349 (N_18349,N_12789,N_13870);
and U18350 (N_18350,N_15290,N_12441);
or U18351 (N_18351,N_14438,N_12672);
nand U18352 (N_18352,N_15664,N_13264);
xnor U18353 (N_18353,N_14706,N_17844);
and U18354 (N_18354,N_13014,N_17504);
nor U18355 (N_18355,N_12013,N_14214);
nand U18356 (N_18356,N_13880,N_14341);
nor U18357 (N_18357,N_12028,N_13505);
nand U18358 (N_18358,N_16605,N_14286);
xor U18359 (N_18359,N_16550,N_15488);
or U18360 (N_18360,N_16018,N_13237);
and U18361 (N_18361,N_16783,N_17533);
nor U18362 (N_18362,N_14005,N_13283);
xor U18363 (N_18363,N_17171,N_15526);
nand U18364 (N_18364,N_17093,N_13285);
xnor U18365 (N_18365,N_14449,N_17963);
and U18366 (N_18366,N_17877,N_15000);
or U18367 (N_18367,N_12007,N_12726);
nand U18368 (N_18368,N_13900,N_13388);
or U18369 (N_18369,N_17071,N_13752);
nand U18370 (N_18370,N_15557,N_16905);
nand U18371 (N_18371,N_16808,N_14492);
nor U18372 (N_18372,N_14914,N_13814);
nor U18373 (N_18373,N_16920,N_15215);
and U18374 (N_18374,N_16733,N_17674);
or U18375 (N_18375,N_13856,N_15361);
nand U18376 (N_18376,N_16329,N_16257);
nand U18377 (N_18377,N_14981,N_15862);
or U18378 (N_18378,N_12494,N_16346);
nand U18379 (N_18379,N_16028,N_17306);
or U18380 (N_18380,N_12398,N_12165);
and U18381 (N_18381,N_12634,N_12817);
and U18382 (N_18382,N_12110,N_16060);
xor U18383 (N_18383,N_12983,N_13337);
nor U18384 (N_18384,N_12978,N_14619);
or U18385 (N_18385,N_13805,N_14491);
nand U18386 (N_18386,N_17328,N_17320);
xor U18387 (N_18387,N_13949,N_14857);
nand U18388 (N_18388,N_15577,N_13394);
nor U18389 (N_18389,N_16070,N_14401);
and U18390 (N_18390,N_15098,N_12838);
nand U18391 (N_18391,N_13019,N_17834);
nor U18392 (N_18392,N_14445,N_16310);
xor U18393 (N_18393,N_14379,N_15050);
xor U18394 (N_18394,N_12986,N_15515);
or U18395 (N_18395,N_13546,N_16395);
xnor U18396 (N_18396,N_16673,N_13303);
or U18397 (N_18397,N_12756,N_13769);
and U18398 (N_18398,N_15618,N_13178);
nor U18399 (N_18399,N_17636,N_13472);
or U18400 (N_18400,N_16994,N_16240);
nand U18401 (N_18401,N_17265,N_12737);
xor U18402 (N_18402,N_14179,N_13985);
xnor U18403 (N_18403,N_12874,N_17926);
nand U18404 (N_18404,N_13539,N_15204);
and U18405 (N_18405,N_12264,N_14664);
xnor U18406 (N_18406,N_17901,N_17361);
and U18407 (N_18407,N_17442,N_14574);
or U18408 (N_18408,N_17336,N_16712);
xnor U18409 (N_18409,N_14411,N_16787);
xor U18410 (N_18410,N_15369,N_14848);
or U18411 (N_18411,N_15970,N_14124);
xnor U18412 (N_18412,N_17914,N_15185);
xnor U18413 (N_18413,N_12338,N_15260);
xor U18414 (N_18414,N_17726,N_15355);
nand U18415 (N_18415,N_14742,N_12922);
nor U18416 (N_18416,N_17054,N_17154);
or U18417 (N_18417,N_12609,N_12618);
xnor U18418 (N_18418,N_17245,N_16781);
or U18419 (N_18419,N_15959,N_17349);
and U18420 (N_18420,N_12241,N_16596);
xnor U18421 (N_18421,N_15834,N_12008);
xnor U18422 (N_18422,N_14302,N_17766);
and U18423 (N_18423,N_16929,N_12608);
nor U18424 (N_18424,N_16056,N_14689);
and U18425 (N_18425,N_14488,N_13163);
and U18426 (N_18426,N_16635,N_16193);
nand U18427 (N_18427,N_13313,N_16703);
nand U18428 (N_18428,N_13105,N_16035);
and U18429 (N_18429,N_15819,N_16385);
xnor U18430 (N_18430,N_15989,N_16155);
or U18431 (N_18431,N_15718,N_14333);
or U18432 (N_18432,N_17606,N_13688);
and U18433 (N_18433,N_12112,N_13565);
xnor U18434 (N_18434,N_14298,N_12439);
or U18435 (N_18435,N_16451,N_16059);
or U18436 (N_18436,N_17711,N_15009);
xnor U18437 (N_18437,N_16520,N_17823);
xnor U18438 (N_18438,N_13798,N_14838);
nor U18439 (N_18439,N_14708,N_16816);
xor U18440 (N_18440,N_14898,N_17572);
or U18441 (N_18441,N_16390,N_14447);
or U18442 (N_18442,N_13396,N_15986);
nor U18443 (N_18443,N_15974,N_17807);
or U18444 (N_18444,N_13883,N_14054);
nand U18445 (N_18445,N_16950,N_16940);
and U18446 (N_18446,N_12775,N_13616);
xor U18447 (N_18447,N_14245,N_15594);
and U18448 (N_18448,N_17365,N_15973);
nor U18449 (N_18449,N_16636,N_14517);
or U18450 (N_18450,N_17389,N_15711);
xnor U18451 (N_18451,N_17221,N_14251);
xnor U18452 (N_18452,N_15914,N_14023);
and U18453 (N_18453,N_16306,N_15710);
or U18454 (N_18454,N_14811,N_16253);
xnor U18455 (N_18455,N_15716,N_17897);
and U18456 (N_18456,N_13465,N_12772);
nor U18457 (N_18457,N_13470,N_14076);
xor U18458 (N_18458,N_14698,N_16430);
or U18459 (N_18459,N_13775,N_12347);
xnor U18460 (N_18460,N_17645,N_17800);
or U18461 (N_18461,N_17457,N_15679);
nand U18462 (N_18462,N_14277,N_12244);
or U18463 (N_18463,N_12044,N_16281);
nand U18464 (N_18464,N_12048,N_15044);
xor U18465 (N_18465,N_13084,N_14812);
nor U18466 (N_18466,N_16842,N_15056);
and U18467 (N_18467,N_14386,N_17820);
nor U18468 (N_18468,N_15299,N_14317);
nand U18469 (N_18469,N_17974,N_14335);
nand U18470 (N_18470,N_16652,N_16353);
nand U18471 (N_18471,N_12552,N_17982);
nor U18472 (N_18472,N_14900,N_13333);
nor U18473 (N_18473,N_13536,N_16025);
nor U18474 (N_18474,N_15689,N_12694);
and U18475 (N_18475,N_17465,N_13842);
nand U18476 (N_18476,N_14691,N_17779);
or U18477 (N_18477,N_12231,N_16206);
nand U18478 (N_18478,N_13043,N_13846);
nor U18479 (N_18479,N_15038,N_15208);
nand U18480 (N_18480,N_12733,N_13044);
nor U18481 (N_18481,N_17754,N_16538);
xor U18482 (N_18482,N_15280,N_17613);
and U18483 (N_18483,N_16162,N_12950);
and U18484 (N_18484,N_17101,N_12719);
nor U18485 (N_18485,N_14733,N_12378);
or U18486 (N_18486,N_12092,N_12763);
nor U18487 (N_18487,N_15830,N_13892);
or U18488 (N_18488,N_16492,N_15658);
nand U18489 (N_18489,N_16874,N_17186);
nor U18490 (N_18490,N_17299,N_13323);
or U18491 (N_18491,N_16852,N_14647);
nor U18492 (N_18492,N_13065,N_14390);
or U18493 (N_18493,N_14604,N_15303);
xor U18494 (N_18494,N_16272,N_17228);
xnor U18495 (N_18495,N_13687,N_14224);
xor U18496 (N_18496,N_16465,N_13335);
nor U18497 (N_18497,N_15133,N_17952);
and U18498 (N_18498,N_15701,N_15961);
nand U18499 (N_18499,N_16986,N_13972);
xnor U18500 (N_18500,N_13614,N_14676);
or U18501 (N_18501,N_15866,N_17191);
and U18502 (N_18502,N_16384,N_13305);
xnor U18503 (N_18503,N_15551,N_17752);
xnor U18504 (N_18504,N_15651,N_16333);
or U18505 (N_18505,N_17657,N_17614);
nor U18506 (N_18506,N_17860,N_15835);
and U18507 (N_18507,N_17813,N_17557);
xnor U18508 (N_18508,N_13722,N_13481);
xor U18509 (N_18509,N_13319,N_13491);
and U18510 (N_18510,N_16584,N_17385);
nor U18511 (N_18511,N_15432,N_16042);
xor U18512 (N_18512,N_15756,N_17382);
and U18513 (N_18513,N_12542,N_12761);
nor U18514 (N_18514,N_15659,N_17826);
or U18515 (N_18515,N_15219,N_16848);
nand U18516 (N_18516,N_14802,N_12260);
nor U18517 (N_18517,N_15022,N_12917);
or U18518 (N_18518,N_12227,N_16135);
xor U18519 (N_18519,N_16032,N_17649);
and U18520 (N_18520,N_14305,N_13888);
and U18521 (N_18521,N_17662,N_14174);
or U18522 (N_18522,N_16719,N_17634);
xnor U18523 (N_18523,N_14629,N_14992);
nand U18524 (N_18524,N_13473,N_16639);
or U18525 (N_18525,N_12780,N_12636);
or U18526 (N_18526,N_16822,N_14382);
and U18527 (N_18527,N_17950,N_13763);
and U18528 (N_18528,N_17639,N_13431);
or U18529 (N_18529,N_17659,N_14618);
or U18530 (N_18530,N_16813,N_13439);
and U18531 (N_18531,N_13279,N_14954);
xor U18532 (N_18532,N_17378,N_12858);
nand U18533 (N_18533,N_12920,N_13268);
xor U18534 (N_18534,N_14164,N_16244);
and U18535 (N_18535,N_15843,N_12650);
xnor U18536 (N_18536,N_12943,N_14679);
nand U18537 (N_18537,N_12724,N_17415);
xnor U18538 (N_18538,N_12071,N_16738);
or U18539 (N_18539,N_14064,N_16641);
and U18540 (N_18540,N_17055,N_12957);
or U18541 (N_18541,N_12171,N_17747);
nand U18542 (N_18542,N_15198,N_14768);
nand U18543 (N_18543,N_14999,N_16117);
and U18544 (N_18544,N_16741,N_17682);
and U18545 (N_18545,N_15889,N_15307);
or U18546 (N_18546,N_14587,N_16105);
nand U18547 (N_18547,N_15416,N_14461);
nor U18548 (N_18548,N_14777,N_17072);
xnor U18549 (N_18549,N_14038,N_12682);
and U18550 (N_18550,N_12271,N_17733);
nor U18551 (N_18551,N_16984,N_17135);
nand U18552 (N_18552,N_16284,N_13445);
and U18553 (N_18553,N_17485,N_14007);
or U18554 (N_18554,N_12953,N_17771);
or U18555 (N_18555,N_14741,N_17407);
xnor U18556 (N_18556,N_12623,N_17564);
xor U18557 (N_18557,N_17705,N_17609);
or U18558 (N_18558,N_14458,N_16642);
and U18559 (N_18559,N_14310,N_12925);
or U18560 (N_18560,N_16659,N_13100);
nand U18561 (N_18561,N_12755,N_13741);
nand U18562 (N_18562,N_17446,N_15815);
or U18563 (N_18563,N_13809,N_14410);
or U18564 (N_18564,N_13937,N_17819);
nand U18565 (N_18565,N_12644,N_16864);
xor U18566 (N_18566,N_13675,N_14089);
xnor U18567 (N_18567,N_14511,N_15575);
nand U18568 (N_18568,N_12397,N_16344);
or U18569 (N_18569,N_17370,N_13988);
and U18570 (N_18570,N_14823,N_15733);
xnor U18571 (N_18571,N_16139,N_15820);
nor U18572 (N_18572,N_15899,N_17134);
nand U18573 (N_18573,N_14677,N_16500);
and U18574 (N_18574,N_17364,N_14116);
nand U18575 (N_18575,N_16687,N_16432);
nand U18576 (N_18576,N_14173,N_12629);
nand U18577 (N_18577,N_15745,N_12182);
and U18578 (N_18578,N_16291,N_16740);
and U18579 (N_18579,N_12405,N_13116);
xor U18580 (N_18580,N_12043,N_14787);
and U18581 (N_18581,N_13729,N_17917);
or U18582 (N_18582,N_13646,N_17984);
nand U18583 (N_18583,N_13570,N_15518);
nand U18584 (N_18584,N_16853,N_15322);
or U18585 (N_18585,N_16397,N_12667);
nor U18586 (N_18586,N_12569,N_17886);
nand U18587 (N_18587,N_15966,N_17008);
or U18588 (N_18588,N_16744,N_16126);
nand U18589 (N_18589,N_16566,N_14327);
and U18590 (N_18590,N_13076,N_14102);
nand U18591 (N_18591,N_16479,N_17744);
nand U18592 (N_18592,N_14985,N_14580);
and U18593 (N_18593,N_12281,N_16737);
nor U18594 (N_18594,N_12040,N_17791);
and U18595 (N_18595,N_14143,N_16704);
and U18596 (N_18596,N_17879,N_12162);
nor U18597 (N_18597,N_17972,N_17646);
nand U18598 (N_18598,N_16543,N_16153);
or U18599 (N_18599,N_14961,N_13497);
and U18600 (N_18600,N_13207,N_15178);
xnor U18601 (N_18601,N_13657,N_12460);
and U18602 (N_18602,N_17396,N_15844);
nor U18603 (N_18603,N_13256,N_14496);
nor U18604 (N_18604,N_14026,N_17331);
or U18605 (N_18605,N_16881,N_15426);
and U18606 (N_18606,N_12310,N_13223);
or U18607 (N_18607,N_14726,N_12919);
nor U18608 (N_18608,N_15740,N_17402);
nand U18609 (N_18609,N_15729,N_13325);
xnor U18610 (N_18610,N_16522,N_13444);
or U18611 (N_18611,N_12999,N_13787);
xnor U18612 (N_18612,N_13525,N_14426);
and U18613 (N_18613,N_12597,N_14093);
xor U18614 (N_18614,N_16953,N_13954);
xor U18615 (N_18615,N_14015,N_12221);
nor U18616 (N_18616,N_17685,N_17346);
nand U18617 (N_18617,N_12729,N_12149);
nand U18618 (N_18618,N_17416,N_12267);
xnor U18619 (N_18619,N_14241,N_15420);
or U18620 (N_18620,N_13795,N_16960);
xor U18621 (N_18621,N_16693,N_17540);
or U18622 (N_18622,N_12615,N_12565);
or U18623 (N_18623,N_12019,N_13837);
and U18624 (N_18624,N_16891,N_13087);
nor U18625 (N_18625,N_15758,N_12864);
and U18626 (N_18626,N_14098,N_17795);
nand U18627 (N_18627,N_16987,N_13669);
and U18628 (N_18628,N_13561,N_12464);
nor U18629 (N_18629,N_15926,N_12004);
and U18630 (N_18630,N_17537,N_13878);
and U18631 (N_18631,N_17721,N_17332);
xnor U18632 (N_18632,N_16263,N_17286);
nor U18633 (N_18633,N_17529,N_14594);
nor U18634 (N_18634,N_13022,N_16754);
and U18635 (N_18635,N_15528,N_14424);
or U18636 (N_18636,N_12798,N_17908);
nand U18637 (N_18637,N_17114,N_16828);
nand U18638 (N_18638,N_14039,N_12076);
nand U18639 (N_18639,N_12435,N_12975);
xor U18640 (N_18640,N_16404,N_16884);
nor U18641 (N_18641,N_15643,N_12147);
and U18642 (N_18642,N_16594,N_12757);
nor U18643 (N_18643,N_13306,N_14311);
or U18644 (N_18644,N_14905,N_12513);
nor U18645 (N_18645,N_12586,N_14325);
xor U18646 (N_18646,N_13772,N_13425);
or U18647 (N_18647,N_15186,N_14397);
and U18648 (N_18648,N_15352,N_15172);
nor U18649 (N_18649,N_13110,N_14254);
and U18650 (N_18650,N_17411,N_12977);
or U18651 (N_18651,N_12229,N_12770);
and U18652 (N_18652,N_17915,N_14818);
nand U18653 (N_18653,N_15400,N_12877);
nand U18654 (N_18654,N_15869,N_15737);
xnor U18655 (N_18655,N_13569,N_16907);
xnor U18656 (N_18656,N_15868,N_15359);
nor U18657 (N_18657,N_12412,N_12300);
nand U18658 (N_18658,N_15870,N_14280);
and U18659 (N_18659,N_13981,N_17097);
and U18660 (N_18660,N_15304,N_17092);
xnor U18661 (N_18661,N_16785,N_12328);
and U18662 (N_18662,N_16918,N_14184);
or U18663 (N_18663,N_15043,N_15905);
xor U18664 (N_18664,N_12191,N_16407);
nor U18665 (N_18665,N_15522,N_16225);
nand U18666 (N_18666,N_17166,N_12010);
or U18667 (N_18667,N_14913,N_17394);
nor U18668 (N_18668,N_13321,N_16328);
nand U18669 (N_18669,N_15106,N_13694);
nor U18670 (N_18670,N_14436,N_14378);
or U18671 (N_18671,N_15221,N_12590);
nand U18672 (N_18672,N_14821,N_12819);
xor U18673 (N_18673,N_13595,N_17831);
or U18674 (N_18674,N_14150,N_13013);
and U18675 (N_18675,N_14729,N_17787);
xnor U18676 (N_18676,N_15247,N_13028);
nand U18677 (N_18677,N_12290,N_12658);
xnor U18678 (N_18678,N_17903,N_16489);
xnor U18679 (N_18679,N_16423,N_15937);
and U18680 (N_18680,N_13709,N_15010);
and U18681 (N_18681,N_12414,N_17932);
and U18682 (N_18682,N_15457,N_13318);
nor U18683 (N_18683,N_17375,N_12674);
nor U18684 (N_18684,N_17719,N_16661);
nand U18685 (N_18685,N_14942,N_16658);
xnor U18686 (N_18686,N_14746,N_17951);
xnor U18687 (N_18687,N_12895,N_16157);
xor U18688 (N_18688,N_12508,N_16241);
or U18689 (N_18689,N_13199,N_16869);
and U18690 (N_18690,N_12769,N_15102);
or U18691 (N_18691,N_13225,N_17156);
xor U18692 (N_18692,N_13699,N_14965);
or U18693 (N_18693,N_17973,N_16149);
nand U18694 (N_18694,N_14216,N_15357);
nor U18695 (N_18695,N_15925,N_13126);
or U18696 (N_18696,N_13398,N_14223);
xnor U18697 (N_18697,N_13075,N_12334);
xnor U18698 (N_18698,N_16954,N_12862);
nand U18699 (N_18699,N_14732,N_14499);
nand U18700 (N_18700,N_13086,N_13609);
nor U18701 (N_18701,N_13241,N_13945);
nand U18702 (N_18702,N_13278,N_14984);
and U18703 (N_18703,N_13326,N_15305);
and U18704 (N_18704,N_15538,N_13492);
nor U18705 (N_18705,N_12547,N_13416);
nand U18706 (N_18706,N_14602,N_12666);
or U18707 (N_18707,N_14238,N_16007);
nor U18708 (N_18708,N_16236,N_17969);
and U18709 (N_18709,N_14903,N_13488);
nand U18710 (N_18710,N_16836,N_16065);
or U18711 (N_18711,N_17257,N_12706);
and U18712 (N_18712,N_16375,N_17277);
or U18713 (N_18713,N_12163,N_16085);
nand U18714 (N_18714,N_13747,N_16237);
and U18715 (N_18715,N_12718,N_17362);
xor U18716 (N_18716,N_14538,N_15609);
nor U18717 (N_18717,N_16979,N_12437);
xnor U18718 (N_18718,N_13288,N_12086);
nand U18719 (N_18719,N_17832,N_12581);
and U18720 (N_18720,N_15648,N_14852);
or U18721 (N_18721,N_16628,N_17736);
and U18722 (N_18722,N_13915,N_13006);
nor U18723 (N_18723,N_15534,N_15680);
and U18724 (N_18724,N_12872,N_17444);
xnor U18725 (N_18725,N_17311,N_16454);
or U18726 (N_18726,N_17716,N_12945);
or U18727 (N_18727,N_12613,N_12987);
nor U18728 (N_18728,N_17936,N_16623);
nand U18729 (N_18729,N_13284,N_13239);
xor U18730 (N_18730,N_17070,N_12278);
nand U18731 (N_18731,N_17971,N_17570);
nor U18732 (N_18732,N_13963,N_13054);
or U18733 (N_18733,N_16039,N_12469);
nand U18734 (N_18734,N_12685,N_13638);
and U18735 (N_18735,N_12324,N_13777);
xnor U18736 (N_18736,N_13538,N_15580);
or U18737 (N_18737,N_13140,N_17770);
and U18738 (N_18738,N_14563,N_14565);
nand U18739 (N_18739,N_12993,N_14571);
nand U18740 (N_18740,N_17273,N_15370);
nand U18741 (N_18741,N_12635,N_17059);
nor U18742 (N_18742,N_12536,N_13652);
or U18743 (N_18743,N_17430,N_14740);
and U18744 (N_18744,N_16293,N_15442);
or U18745 (N_18745,N_16399,N_12285);
xor U18746 (N_18746,N_16902,N_17425);
and U18747 (N_18747,N_13879,N_14101);
and U18748 (N_18748,N_14730,N_15971);
or U18749 (N_18749,N_12381,N_16899);
nor U18750 (N_18750,N_12699,N_15638);
or U18751 (N_18751,N_16760,N_12931);
and U18752 (N_18752,N_14973,N_15571);
nand U18753 (N_18753,N_16189,N_15326);
and U18754 (N_18754,N_13269,N_16387);
nor U18755 (N_18755,N_13951,N_13456);
and U18756 (N_18756,N_16608,N_16956);
and U18757 (N_18757,N_17241,N_12394);
nor U18758 (N_18758,N_17507,N_13676);
nor U18759 (N_18759,N_16524,N_12611);
xnor U18760 (N_18760,N_17593,N_15639);
nor U18761 (N_18761,N_13926,N_16736);
nor U18762 (N_18762,N_13294,N_13068);
xnor U18763 (N_18763,N_16685,N_12177);
xnor U18764 (N_18764,N_12927,N_15957);
and U18765 (N_18765,N_13053,N_12490);
nand U18766 (N_18766,N_17641,N_15997);
or U18767 (N_18767,N_12882,N_17527);
xor U18768 (N_18768,N_17456,N_14720);
nand U18769 (N_18769,N_13011,N_17472);
nor U18770 (N_18770,N_12924,N_14590);
nor U18771 (N_18771,N_13755,N_12384);
xor U18772 (N_18772,N_12103,N_14844);
xor U18773 (N_18773,N_14990,N_14112);
nand U18774 (N_18774,N_14955,N_13786);
nor U18775 (N_18775,N_15226,N_13441);
xnor U18776 (N_18776,N_15417,N_15552);
nand U18777 (N_18777,N_16893,N_14681);
nor U18778 (N_18778,N_12037,N_13989);
xnor U18779 (N_18779,N_15760,N_15332);
xor U18780 (N_18780,N_12734,N_17212);
and U18781 (N_18781,N_16103,N_17843);
and U18782 (N_18782,N_17218,N_13610);
nor U18783 (N_18783,N_15317,N_16928);
nor U18784 (N_18784,N_14859,N_16141);
and U18785 (N_18785,N_17522,N_17152);
nor U18786 (N_18786,N_13414,N_15144);
and U18787 (N_18787,N_15207,N_17414);
nand U18788 (N_18788,N_14253,N_17006);
nor U18789 (N_18789,N_14285,N_15806);
and U18790 (N_18790,N_13745,N_13151);
or U18791 (N_18791,N_16212,N_12051);
and U18792 (N_18792,N_13847,N_17392);
and U18793 (N_18793,N_16807,N_14704);
nor U18794 (N_18794,N_14331,N_13923);
and U18795 (N_18795,N_15404,N_13298);
xnor U18796 (N_18796,N_16882,N_12169);
nand U18797 (N_18797,N_17957,N_12111);
xor U18798 (N_18798,N_17975,N_13596);
or U18799 (N_18799,N_15403,N_16254);
xnor U18800 (N_18800,N_16617,N_17201);
nor U18801 (N_18801,N_16398,N_12411);
nor U18802 (N_18802,N_13751,N_17748);
and U18803 (N_18803,N_12263,N_14573);
nor U18804 (N_18804,N_14960,N_13104);
and U18805 (N_18805,N_14349,N_16698);
xor U18806 (N_18806,N_15962,N_12252);
xnor U18807 (N_18807,N_12428,N_13047);
nor U18808 (N_18808,N_16812,N_15995);
xor U18809 (N_18809,N_13936,N_15793);
and U18810 (N_18810,N_14516,N_12821);
nor U18811 (N_18811,N_15120,N_12544);
nand U18812 (N_18812,N_15464,N_13138);
xor U18813 (N_18813,N_15874,N_14968);
nor U18814 (N_18814,N_12773,N_14465);
and U18815 (N_18815,N_16502,N_15568);
xor U18816 (N_18816,N_15851,N_16799);
or U18817 (N_18817,N_13166,N_16964);
or U18818 (N_18818,N_13603,N_13750);
or U18819 (N_18819,N_15248,N_17209);
xor U18820 (N_18820,N_13655,N_14639);
or U18821 (N_18821,N_17232,N_14373);
nor U18822 (N_18822,N_14813,N_15895);
xor U18823 (N_18823,N_17895,N_14068);
xor U18824 (N_18824,N_12288,N_15011);
nand U18825 (N_18825,N_15969,N_12820);
nor U18826 (N_18826,N_16957,N_17983);
nor U18827 (N_18827,N_14272,N_12795);
nand U18828 (N_18828,N_14393,N_14294);
and U18829 (N_18829,N_15478,N_16137);
or U18830 (N_18830,N_17231,N_16924);
xnor U18831 (N_18831,N_17991,N_13403);
nor U18832 (N_18832,N_15256,N_15589);
nand U18833 (N_18833,N_15194,N_12245);
xnor U18834 (N_18834,N_13556,N_12502);
and U18835 (N_18835,N_17715,N_12480);
xor U18836 (N_18836,N_13591,N_15717);
nor U18837 (N_18837,N_17994,N_14974);
nor U18838 (N_18838,N_16680,N_14147);
nor U18839 (N_18839,N_14528,N_13203);
nor U18840 (N_18840,N_12457,N_16930);
nor U18841 (N_18841,N_12201,N_12871);
or U18842 (N_18842,N_16776,N_15356);
and U18843 (N_18843,N_17539,N_17839);
nand U18844 (N_18844,N_17675,N_17528);
or U18845 (N_18845,N_14088,N_15539);
nor U18846 (N_18846,N_15018,N_12211);
xor U18847 (N_18847,N_14148,N_17139);
nand U18848 (N_18848,N_14997,N_15797);
nor U18849 (N_18849,N_17302,N_12514);
or U18850 (N_18850,N_14917,N_13449);
xor U18851 (N_18851,N_16484,N_13877);
xnor U18852 (N_18852,N_14745,N_12012);
nor U18853 (N_18853,N_13377,N_13423);
nor U18854 (N_18854,N_12023,N_14552);
and U18855 (N_18855,N_13690,N_15544);
nor U18856 (N_18856,N_17550,N_16831);
nand U18857 (N_18857,N_15601,N_15847);
xor U18858 (N_18858,N_16949,N_14387);
nand U18859 (N_18859,N_15956,N_14047);
nor U18860 (N_18860,N_16160,N_15082);
nand U18861 (N_18861,N_12778,N_13544);
and U18862 (N_18862,N_14190,N_14982);
or U18863 (N_18863,N_14504,N_14268);
nor U18864 (N_18864,N_17574,N_13070);
or U18865 (N_18865,N_17552,N_12958);
nand U18866 (N_18866,N_17254,N_17656);
nand U18867 (N_18867,N_16469,N_16562);
nor U18868 (N_18868,N_15379,N_16194);
xor U18869 (N_18869,N_14713,N_16181);
nand U18870 (N_18870,N_14967,N_12511);
nor U18871 (N_18871,N_15624,N_12901);
xor U18872 (N_18872,N_17690,N_12475);
nor U18873 (N_18873,N_15161,N_13987);
and U18874 (N_18874,N_13023,N_12422);
or U18875 (N_18875,N_13531,N_17086);
or U18876 (N_18876,N_16403,N_17806);
nand U18877 (N_18877,N_17048,N_12485);
or U18878 (N_18878,N_15512,N_16071);
nand U18879 (N_18879,N_13744,N_12621);
and U18880 (N_18880,N_13380,N_13580);
and U18881 (N_18881,N_17612,N_12735);
nand U18882 (N_18882,N_16980,N_17585);
or U18883 (N_18883,N_16714,N_16824);
xor U18884 (N_18884,N_15193,N_15469);
or U18885 (N_18885,N_12348,N_12332);
or U18886 (N_18886,N_16273,N_15795);
nand U18887 (N_18887,N_15273,N_12960);
xnor U18888 (N_18888,N_17452,N_16798);
xnor U18889 (N_18889,N_12289,N_17828);
and U18890 (N_18890,N_15855,N_14222);
nand U18891 (N_18891,N_13502,N_14288);
nand U18892 (N_18892,N_14067,N_15588);
nor U18893 (N_18893,N_12242,N_17742);
and U18894 (N_18894,N_15714,N_13632);
or U18895 (N_18895,N_16198,N_15131);
or U18896 (N_18896,N_12036,N_14107);
or U18897 (N_18897,N_14198,N_16358);
nand U18898 (N_18898,N_16114,N_14856);
and U18899 (N_18899,N_15562,N_13240);
nand U18900 (N_18900,N_17872,N_14463);
nand U18901 (N_18901,N_13807,N_16211);
nand U18902 (N_18902,N_14510,N_15507);
or U18903 (N_18903,N_16900,N_12391);
or U18904 (N_18904,N_14876,N_17815);
nor U18905 (N_18905,N_17366,N_17500);
nor U18906 (N_18906,N_13395,N_12443);
and U18907 (N_18907,N_16446,N_17495);
nor U18908 (N_18908,N_13667,N_13927);
nand U18909 (N_18909,N_17558,N_14928);
xnor U18910 (N_18910,N_14053,N_14041);
and U18911 (N_18911,N_13248,N_16443);
nor U18912 (N_18912,N_16146,N_17226);
xnor U18913 (N_18913,N_14886,N_17698);
nand U18914 (N_18914,N_13349,N_15249);
nand U18915 (N_18915,N_16978,N_16743);
or U18916 (N_18916,N_14494,N_13397);
or U18917 (N_18917,N_12750,N_14175);
nand U18918 (N_18918,N_12933,N_12605);
nand U18919 (N_18919,N_13063,N_13633);
nand U18920 (N_18920,N_14794,N_16116);
nand U18921 (N_18921,N_17693,N_12743);
and U18922 (N_18922,N_15503,N_12701);
xnor U18923 (N_18923,N_12880,N_15565);
nor U18924 (N_18924,N_12712,N_13994);
nand U18925 (N_18925,N_16553,N_12361);
and U18926 (N_18926,N_17145,N_13521);
or U18927 (N_18927,N_15362,N_13990);
or U18928 (N_18928,N_13242,N_13357);
xor U18929 (N_18929,N_17487,N_14927);
or U18930 (N_18930,N_16976,N_16402);
nand U18931 (N_18931,N_15996,N_14252);
and U18932 (N_18932,N_13617,N_16593);
nor U18933 (N_18933,N_16879,N_12825);
xor U18934 (N_18934,N_17263,N_17356);
or U18935 (N_18935,N_17439,N_17317);
nand U18936 (N_18936,N_17595,N_12866);
or U18937 (N_18937,N_16287,N_15771);
nor U18938 (N_18938,N_13686,N_13246);
nor U18939 (N_18939,N_13737,N_17110);
nor U18940 (N_18940,N_15259,N_16926);
or U18941 (N_18941,N_12307,N_17464);
or U18942 (N_18942,N_17569,N_14570);
nand U18943 (N_18943,N_15030,N_17285);
or U18944 (N_18944,N_17125,N_17236);
nand U18945 (N_18945,N_14236,N_14388);
or U18946 (N_18946,N_12344,N_15536);
nand U18947 (N_18947,N_17945,N_15919);
nor U18948 (N_18948,N_13429,N_14443);
xor U18949 (N_18949,N_15064,N_16033);
nand U18950 (N_18950,N_13236,N_15832);
xor U18951 (N_18951,N_16343,N_14865);
xnor U18952 (N_18952,N_12857,N_14711);
nor U18953 (N_18953,N_15275,N_17506);
xor U18954 (N_18954,N_14279,N_12135);
and U18955 (N_18955,N_15032,N_15039);
xnor U18956 (N_18956,N_12914,N_16910);
nand U18957 (N_18957,N_17509,N_16046);
and U18958 (N_18958,N_16199,N_17728);
and U18959 (N_18959,N_17988,N_15447);
nand U18960 (N_18960,N_17024,N_14450);
nor U18961 (N_18961,N_17921,N_17314);
nand U18962 (N_18962,N_17371,N_14264);
and U18963 (N_18963,N_13523,N_16021);
nor U18964 (N_18964,N_12973,N_15393);
nor U18965 (N_18965,N_17038,N_12298);
xor U18966 (N_18966,N_13517,N_17941);
nor U18967 (N_18967,N_16439,N_14581);
nand U18968 (N_18968,N_15395,N_13484);
nor U18969 (N_18969,N_17391,N_16386);
and U18970 (N_18970,N_13064,N_13471);
or U18971 (N_18971,N_12368,N_15254);
or U18972 (N_18972,N_14213,N_15608);
xnor U18973 (N_18973,N_14322,N_17083);
xnor U18974 (N_18974,N_17610,N_16561);
nand U18975 (N_18975,N_17293,N_14762);
nand U18976 (N_18976,N_16123,N_14791);
or U18977 (N_18977,N_13412,N_13332);
or U18978 (N_18978,N_12096,N_15412);
nor U18979 (N_18979,N_13659,N_15149);
nor U18980 (N_18980,N_13974,N_12686);
or U18981 (N_18981,N_16372,N_14295);
and U18982 (N_18982,N_16170,N_12584);
nor U18983 (N_18983,N_14319,N_17591);
nand U18984 (N_18984,N_15385,N_15205);
nor U18985 (N_18985,N_12366,N_14493);
nor U18986 (N_18986,N_17707,N_13808);
nand U18987 (N_18987,N_16091,N_15293);
nand U18988 (N_18988,N_15243,N_15233);
nor U18989 (N_18989,N_16080,N_12967);
or U18990 (N_18990,N_16894,N_16218);
nand U18991 (N_18991,N_17562,N_12192);
or U18992 (N_18992,N_16510,N_17117);
nor U18993 (N_18993,N_14209,N_13393);
nand U18994 (N_18994,N_17651,N_15901);
nor U18995 (N_18995,N_17195,N_16690);
nand U18996 (N_18996,N_13315,N_13046);
or U18997 (N_18997,N_12913,N_15554);
nand U18998 (N_18998,N_17175,N_12847);
nand U18999 (N_18999,N_15481,N_17179);
and U19000 (N_19000,N_13274,N_13487);
nand U19001 (N_19001,N_14284,N_16217);
nor U19002 (N_19002,N_16360,N_12279);
nor U19003 (N_19003,N_14953,N_14276);
and U19004 (N_19004,N_13822,N_16675);
or U19005 (N_19005,N_16655,N_14585);
xnor U19006 (N_19006,N_15936,N_12466);
nand U19007 (N_19007,N_14853,N_17298);
nand U19008 (N_19008,N_16511,N_15814);
nor U19009 (N_19009,N_17925,N_14300);
and U19010 (N_19010,N_17115,N_17989);
nand U19011 (N_19011,N_16013,N_14316);
or U19012 (N_19012,N_12208,N_16722);
xor U19013 (N_19013,N_14949,N_13813);
nand U19014 (N_19014,N_14993,N_16968);
nand U19015 (N_19015,N_17599,N_14500);
or U19016 (N_19016,N_16497,N_17801);
nor U19017 (N_19017,N_16633,N_17964);
or U19018 (N_19018,N_17002,N_17348);
nor U19019 (N_19019,N_15738,N_13124);
and U19020 (N_19020,N_16904,N_12079);
nor U19021 (N_19021,N_15040,N_12254);
nand U19022 (N_19022,N_15825,N_16077);
and U19023 (N_19023,N_17626,N_15892);
and U19024 (N_19024,N_17387,N_17835);
nand U19025 (N_19025,N_13433,N_12379);
nor U19026 (N_19026,N_14389,N_13408);
nor U19027 (N_19027,N_13766,N_16580);
nand U19028 (N_19028,N_12121,N_15502);
and U19029 (N_19029,N_17308,N_13148);
or U19030 (N_19030,N_12054,N_16750);
nor U19031 (N_19031,N_16606,N_13810);
or U19032 (N_19032,N_12548,N_12387);
nor U19033 (N_19033,N_17448,N_12131);
nor U19034 (N_19034,N_13906,N_13495);
and U19035 (N_19035,N_17453,N_12098);
nand U19036 (N_19036,N_17229,N_16911);
and U19037 (N_19037,N_13437,N_13553);
xor U19038 (N_19038,N_12687,N_12938);
xor U19039 (N_19039,N_12939,N_13327);
and U19040 (N_19040,N_14767,N_13639);
nand U19041 (N_19041,N_17420,N_17124);
or U19042 (N_19042,N_14033,N_17667);
xor U19043 (N_19043,N_15380,N_16279);
nand U19044 (N_19044,N_17350,N_17825);
and U19045 (N_19045,N_13913,N_17997);
nor U19046 (N_19046,N_12497,N_12168);
nand U19047 (N_19047,N_15066,N_15724);
nor U19048 (N_19048,N_15640,N_16537);
xor U19049 (N_19049,N_14375,N_13254);
nand U19050 (N_19050,N_17761,N_14234);
nand U19051 (N_19051,N_15676,N_16663);
nand U19052 (N_19052,N_17249,N_13049);
xnor U19053 (N_19053,N_15791,N_15645);
nand U19054 (N_19054,N_12164,N_12088);
nand U19055 (N_19055,N_12042,N_12782);
nand U19056 (N_19056,N_16650,N_17774);
xnor U19057 (N_19057,N_14601,N_12350);
nand U19058 (N_19058,N_13224,N_12139);
or U19059 (N_19059,N_17724,N_15785);
or U19060 (N_19060,N_17616,N_17429);
and U19061 (N_19061,N_12093,N_17954);
and U19062 (N_19062,N_17778,N_16868);
or U19063 (N_19063,N_14854,N_17661);
or U19064 (N_19064,N_14082,N_12991);
xnor U19065 (N_19065,N_12749,N_15993);
nand U19066 (N_19066,N_16764,N_13730);
nor U19067 (N_19067,N_13602,N_13943);
or U19068 (N_19068,N_17995,N_17618);
xor U19069 (N_19069,N_13942,N_15747);
nand U19070 (N_19070,N_13723,N_17655);
and U19071 (N_19071,N_15826,N_12459);
nand U19072 (N_19072,N_16164,N_17898);
nor U19073 (N_19073,N_15212,N_17323);
nand U19074 (N_19074,N_15127,N_13486);
nor U19075 (N_19075,N_12032,N_17140);
or U19076 (N_19076,N_15327,N_12389);
nor U19077 (N_19077,N_17802,N_13211);
nand U19078 (N_19078,N_15320,N_15225);
or U19079 (N_19079,N_14467,N_16379);
nand U19080 (N_19080,N_17803,N_16031);
nor U19081 (N_19081,N_16866,N_14956);
or U19082 (N_19082,N_12345,N_13784);
nor U19083 (N_19083,N_16122,N_15190);
nor U19084 (N_19084,N_14119,N_13574);
or U19085 (N_19085,N_14123,N_17548);
or U19086 (N_19086,N_16265,N_14030);
xnor U19087 (N_19087,N_16528,N_14380);
nor U19088 (N_19088,N_15980,N_17594);
and U19089 (N_19089,N_14659,N_12180);
nor U19090 (N_19090,N_12301,N_12077);
and U19091 (N_19091,N_14354,N_13476);
and U19092 (N_19092,N_15218,N_14263);
and U19093 (N_19093,N_15520,N_16773);
or U19094 (N_19094,N_12337,N_13829);
nand U19095 (N_19095,N_17104,N_17981);
or U19096 (N_19096,N_16849,N_13150);
nor U19097 (N_19097,N_14548,N_14369);
or U19098 (N_19098,N_13438,N_14462);
xnor U19099 (N_19099,N_13060,N_13642);
nand U19100 (N_19100,N_17479,N_17143);
nand U19101 (N_19101,N_14645,N_15865);
nor U19102 (N_19102,N_13113,N_14701);
xor U19103 (N_19103,N_17809,N_16505);
or U19104 (N_19104,N_17422,N_16725);
and U19105 (N_19105,N_16335,N_12894);
nor U19106 (N_19106,N_17633,N_12722);
and U19107 (N_19107,N_15549,N_13212);
xor U19108 (N_19108,N_15772,N_16258);
xor U19109 (N_19109,N_17944,N_16626);
or U19110 (N_19110,N_15726,N_13307);
nor U19111 (N_19111,N_15232,N_17329);
nand U19112 (N_19112,N_15097,N_12574);
and U19113 (N_19113,N_13360,N_16898);
xnor U19114 (N_19114,N_15311,N_12114);
and U19115 (N_19115,N_16491,N_15695);
nand U19116 (N_19116,N_14977,N_12393);
nor U19117 (N_19117,N_15827,N_15348);
and U19118 (N_19118,N_15061,N_16532);
nand U19119 (N_19119,N_12601,N_15103);
or U19120 (N_19120,N_12205,N_16079);
nand U19121 (N_19121,N_12424,N_16228);
nand U19122 (N_19122,N_16371,N_16621);
or U19123 (N_19123,N_12266,N_13713);
or U19124 (N_19124,N_14941,N_13365);
nand U19125 (N_19125,N_16880,N_13980);
or U19126 (N_19126,N_17797,N_13914);
nand U19127 (N_19127,N_14815,N_15292);
xor U19128 (N_19128,N_12233,N_17894);
xor U19129 (N_19129,N_12662,N_17782);
or U19130 (N_19130,N_17132,N_15787);
nand U19131 (N_19131,N_12179,N_17473);
and U19132 (N_19132,N_15171,N_14700);
nor U19133 (N_19133,N_14692,N_12851);
or U19134 (N_19134,N_13073,N_12315);
nor U19135 (N_19135,N_12910,N_17085);
and U19136 (N_19136,N_12646,N_14414);
and U19137 (N_19137,N_15656,N_13362);
xnor U19138 (N_19138,N_14763,N_13158);
and U19139 (N_19139,N_16232,N_17341);
or U19140 (N_19140,N_15917,N_17290);
or U19141 (N_19141,N_14873,N_13815);
nand U19142 (N_19142,N_15313,N_16144);
xnor U19143 (N_19143,N_14337,N_14807);
nand U19144 (N_19144,N_16547,N_16355);
and U19145 (N_19145,N_13993,N_16700);
and U19146 (N_19146,N_13426,N_15616);
xnor U19147 (N_19147,N_13890,N_12203);
nand U19148 (N_19148,N_17666,N_12525);
or U19149 (N_19149,N_14356,N_12900);
nand U19150 (N_19150,N_15285,N_16804);
xor U19151 (N_19151,N_16932,N_14399);
nand U19152 (N_19152,N_14889,N_16231);
nor U19153 (N_19153,N_17150,N_12683);
nor U19154 (N_19154,N_15096,N_14437);
nand U19155 (N_19155,N_12730,N_17217);
nand U19156 (N_19156,N_14611,N_16833);
or U19157 (N_19157,N_14201,N_17334);
and U19158 (N_19158,N_14727,N_16896);
xor U19159 (N_19159,N_16669,N_15441);
xnor U19160 (N_19160,N_15845,N_16724);
nand U19161 (N_19161,N_12884,N_17207);
or U19162 (N_19162,N_17746,N_13091);
or U19163 (N_19163,N_12606,N_16651);
nor U19164 (N_19164,N_14957,N_15734);
nor U19165 (N_19165,N_12392,N_14899);
and U19166 (N_19166,N_17049,N_17653);
xor U19167 (N_19167,N_14055,N_15911);
nand U19168 (N_19168,N_17868,N_14210);
nand U19169 (N_19169,N_16434,N_17935);
xor U19170 (N_19170,N_13677,N_14723);
or U19171 (N_19171,N_16972,N_12997);
xor U19172 (N_19172,N_12966,N_15761);
nand U19173 (N_19173,N_14395,N_12108);
nand U19174 (N_19174,N_15650,N_13781);
nor U19175 (N_19175,N_15527,N_13386);
and U19176 (N_19176,N_14615,N_13791);
nor U19177 (N_19177,N_12115,N_17130);
nor U19178 (N_19178,N_13261,N_13738);
xnor U19179 (N_19179,N_15268,N_16756);
and U19180 (N_19180,N_14440,N_16084);
and U19181 (N_19181,N_12085,N_16101);
or U19182 (N_19182,N_15721,N_12799);
xnor U19183 (N_19183,N_17729,N_17607);
xor U19184 (N_19184,N_17676,N_15069);
xnor U19185 (N_19185,N_15114,N_16394);
nor U19186 (N_19186,N_13103,N_14800);
nand U19187 (N_19187,N_15720,N_13127);
nand U19188 (N_19188,N_14779,N_17210);
or U19189 (N_19189,N_13080,N_15878);
and U19190 (N_19190,N_15694,N_13637);
or U19191 (N_19191,N_12286,N_17788);
xnor U19192 (N_19192,N_15840,N_13375);
xor U19193 (N_19193,N_15297,N_12275);
xnor U19194 (N_19194,N_13273,N_16416);
xor U19195 (N_19195,N_12711,N_13402);
nor U19196 (N_19196,N_17066,N_17381);
and U19197 (N_19197,N_12971,N_12656);
nor U19198 (N_19198,N_14120,N_17068);
and U19199 (N_19199,N_14564,N_14600);
and U19200 (N_19200,N_16490,N_17924);
nor U19201 (N_19201,N_13295,N_14019);
or U19202 (N_19202,N_17460,N_15439);
xnor U19203 (N_19203,N_12598,N_12752);
and U19204 (N_19204,N_13625,N_14096);
or U19205 (N_19205,N_15431,N_14951);
and U19206 (N_19206,N_14308,N_16026);
nand U19207 (N_19207,N_15697,N_12476);
and U19208 (N_19208,N_16723,N_17027);
or U19209 (N_19209,N_17075,N_15523);
and U19210 (N_19210,N_13955,N_17058);
nor U19211 (N_19211,N_15282,N_14239);
nand U19212 (N_19212,N_17732,N_15462);
nand U19213 (N_19213,N_14016,N_16453);
and U19214 (N_19214,N_17102,N_13025);
xor U19215 (N_19215,N_16951,N_17953);
xnor U19216 (N_19216,N_14297,N_12200);
nor U19217 (N_19217,N_14318,N_12295);
nor U19218 (N_19218,N_13581,N_13226);
xor U19219 (N_19219,N_15117,N_14863);
xnor U19220 (N_19220,N_16989,N_15988);
nand U19221 (N_19221,N_13344,N_15908);
and U19222 (N_19222,N_15059,N_13924);
and U19223 (N_19223,N_17106,N_16513);
nand U19224 (N_19224,N_17089,N_12371);
nor U19225 (N_19225,N_17021,N_12416);
and U19226 (N_19226,N_12860,N_16865);
xor U19227 (N_19227,N_15378,N_14484);
and U19228 (N_19228,N_14056,N_12172);
or U19229 (N_19229,N_17413,N_16426);
xor U19230 (N_19230,N_15199,N_15353);
xor U19231 (N_19231,N_17224,N_16020);
or U19232 (N_19232,N_12765,N_13758);
nand U19233 (N_19233,N_15281,N_14346);
and U19234 (N_19234,N_13940,N_15168);
and U19235 (N_19235,N_12062,N_15242);
nand U19236 (N_19236,N_13244,N_16036);
nand U19237 (N_19237,N_16006,N_13983);
xor U19238 (N_19238,N_12762,N_17326);
and U19239 (N_19239,N_13334,N_14912);
xnor U19240 (N_19240,N_17313,N_17162);
nor U19241 (N_19241,N_14293,N_17783);
or U19242 (N_19242,N_12580,N_12717);
nor U19243 (N_19243,N_13803,N_13041);
nand U19244 (N_19244,N_12881,N_12523);
nand U19245 (N_19245,N_13245,N_13190);
or U19246 (N_19246,N_13771,N_17372);
nand U19247 (N_19247,N_14374,N_13997);
and U19248 (N_19248,N_13317,N_15690);
nor U19249 (N_19249,N_12431,N_17962);
nand U19250 (N_19250,N_16670,N_13886);
nor U19251 (N_19251,N_14925,N_13705);
nand U19252 (N_19252,N_17488,N_17841);
xnor U19253 (N_19253,N_13541,N_15517);
nor U19254 (N_19254,N_16393,N_16747);
and U19255 (N_19255,N_12589,N_17684);
or U19256 (N_19256,N_17694,N_12815);
and U19257 (N_19257,N_13442,N_14008);
nand U19258 (N_19258,N_14798,N_17324);
or U19259 (N_19259,N_16745,N_14031);
nand U19260 (N_19260,N_15846,N_12410);
xnor U19261 (N_19261,N_17177,N_16775);
nand U19262 (N_19262,N_14797,N_12642);
and U19263 (N_19263,N_16708,N_16758);
and U19264 (N_19264,N_17428,N_17621);
xnor U19265 (N_19265,N_15354,N_16134);
or U19266 (N_19266,N_12453,N_15455);
and U19267 (N_19267,N_16405,N_13979);
or U19268 (N_19268,N_15985,N_14177);
nand U19269 (N_19269,N_17628,N_13061);
xnor U19270 (N_19270,N_13704,N_14180);
and U19271 (N_19271,N_17692,N_17629);
xor U19272 (N_19272,N_12374,N_13389);
nor U19273 (N_19273,N_12487,N_14598);
or U19274 (N_19274,N_14012,N_15893);
and U19275 (N_19275,N_15165,N_15073);
and U19276 (N_19276,N_14592,N_13167);
or U19277 (N_19277,N_12876,N_14324);
and U19278 (N_19278,N_17122,N_13952);
nand U19279 (N_19279,N_17498,N_15723);
and U19280 (N_19280,N_16856,N_14313);
nor U19281 (N_19281,N_16169,N_16731);
nand U19282 (N_19282,N_12856,N_15633);
and U19283 (N_19283,N_12806,N_16288);
nand U19284 (N_19284,N_13066,N_13693);
nand U19285 (N_19285,N_16271,N_14935);
nand U19286 (N_19286,N_17773,N_17808);
nand U19287 (N_19287,N_14696,N_14365);
xor U19288 (N_19288,N_13912,N_17269);
nor U19289 (N_19289,N_16285,N_14540);
nor U19290 (N_19290,N_13761,N_17798);
and U19291 (N_19291,N_17073,N_13925);
and U19292 (N_19292,N_17151,N_13050);
nand U19293 (N_19293,N_13123,N_15047);
nor U19294 (N_19294,N_14892,N_15173);
or U19295 (N_19295,N_17436,N_17142);
nor U19296 (N_19296,N_16598,N_12097);
nand U19297 (N_19297,N_12359,N_14188);
nand U19298 (N_19298,N_15912,N_16452);
xor U19299 (N_19299,N_14534,N_17789);
nor U19300 (N_19300,N_15707,N_14250);
nor U19301 (N_19301,N_17642,N_14194);
or U19302 (N_19302,N_16094,N_16697);
and U19303 (N_19303,N_15237,N_13155);
nand U19304 (N_19304,N_12715,N_16378);
nor U19305 (N_19305,N_13540,N_14274);
nand U19306 (N_19306,N_13874,N_17510);
nand U19307 (N_19307,N_12936,N_16886);
or U19308 (N_19308,N_15533,N_12261);
or U19309 (N_19309,N_13033,N_13510);
and U19310 (N_19310,N_15333,N_15660);
nand U19311 (N_19311,N_13042,N_15894);
xor U19312 (N_19312,N_14850,N_13131);
xnor U19313 (N_19313,N_14649,N_15495);
xor U19314 (N_19314,N_17644,N_15902);
nand U19315 (N_19315,N_12448,N_14754);
nor U19316 (N_19316,N_14501,N_12912);
nand U19317 (N_19317,N_14103,N_12677);
nor U19318 (N_19318,N_17173,N_13275);
nand U19319 (N_19319,N_14185,N_16121);
or U19320 (N_19320,N_14660,N_16068);
nand U19321 (N_19321,N_16644,N_17827);
or U19322 (N_19322,N_13780,N_17816);
xor U19323 (N_19323,N_12655,N_17695);
nand U19324 (N_19324,N_15121,N_12786);
xor U19325 (N_19325,N_14790,N_15497);
nand U19326 (N_19326,N_15414,N_12905);
nor U19327 (N_19327,N_13764,N_15712);
nand U19328 (N_19328,N_14827,N_17242);
xnor U19329 (N_19329,N_12668,N_17545);
xnor U19330 (N_19330,N_14719,N_17930);
or U19331 (N_19331,N_12125,N_14459);
nor U19332 (N_19332,N_17005,N_14930);
nor U19333 (N_19333,N_12376,N_16990);
or U19334 (N_19334,N_12708,N_13188);
nor U19335 (N_19335,N_15752,N_14906);
and U19336 (N_19336,N_14666,N_13461);
or U19337 (N_19337,N_14478,N_12306);
nand U19338 (N_19338,N_14532,N_12784);
or U19339 (N_19339,N_15486,N_13898);
or U19340 (N_19340,N_12916,N_17696);
or U19341 (N_19341,N_16778,N_15547);
xnor U19342 (N_19342,N_14028,N_16889);
and U19343 (N_19343,N_12732,N_14705);
or U19344 (N_19344,N_15261,N_17561);
nor U19345 (N_19345,N_17704,N_17584);
nor U19346 (N_19346,N_13085,N_16933);
and U19347 (N_19347,N_13630,N_12404);
or U19348 (N_19348,N_15093,N_14235);
xor U19349 (N_19349,N_16516,N_16406);
and U19350 (N_19350,N_15842,N_13806);
xor U19351 (N_19351,N_12535,N_12174);
or U19352 (N_19352,N_13198,N_14195);
or U19353 (N_19353,N_15463,N_17845);
or U19354 (N_19354,N_14159,N_15798);
nor U19355 (N_19355,N_12524,N_14141);
or U19356 (N_19356,N_15351,N_12528);
or U19357 (N_19357,N_12311,N_12220);
and U19358 (N_19358,N_15610,N_13790);
or U19359 (N_19359,N_17553,N_17076);
xnor U19360 (N_19360,N_13355,N_13867);
and U19361 (N_19361,N_13792,N_12020);
nand U19362 (N_19362,N_12175,N_14665);
nor U19363 (N_19363,N_14229,N_12520);
and U19364 (N_19364,N_15975,N_17198);
nor U19365 (N_19365,N_14609,N_15605);
or U19366 (N_19366,N_13142,N_15916);
nand U19367 (N_19367,N_16389,N_16326);
or U19368 (N_19368,N_13605,N_13965);
and U19369 (N_19369,N_14628,N_14412);
or U19370 (N_19370,N_13626,N_16303);
or U19371 (N_19371,N_13598,N_13577);
or U19372 (N_19372,N_12209,N_12099);
nand U19373 (N_19373,N_14237,N_16696);
xor U19374 (N_19374,N_15573,N_15910);
and U19375 (N_19375,N_13161,N_17968);
nand U19376 (N_19376,N_12959,N_13132);
or U19377 (N_19377,N_12940,N_16321);
xor U19378 (N_19378,N_17174,N_15808);
and U19379 (N_19379,N_12447,N_15267);
nand U19380 (N_19380,N_17309,N_13930);
nor U19381 (N_19381,N_17672,N_12664);
xnor U19382 (N_19382,N_15742,N_14489);
nand U19383 (N_19383,N_16531,N_14273);
xnor U19384 (N_19384,N_17751,N_13721);
and U19385 (N_19385,N_12128,N_15569);
xnor U19386 (N_19386,N_17590,N_12303);
nor U19387 (N_19387,N_16936,N_14323);
xor U19388 (N_19388,N_14524,N_15058);
or U19389 (N_19389,N_15574,N_15100);
or U19390 (N_19390,N_13435,N_13250);
nand U19391 (N_19391,N_15931,N_13055);
and U19392 (N_19392,N_15336,N_13262);
nor U19393 (N_19393,N_16349,N_12058);
or U19394 (N_19394,N_12481,N_13622);
nand U19395 (N_19395,N_17438,N_16061);
xor U19396 (N_19396,N_16435,N_14215);
xor U19397 (N_19397,N_12828,N_17441);
xnor U19398 (N_19398,N_16573,N_14752);
or U19399 (N_19399,N_15316,N_13217);
nand U19400 (N_19400,N_12673,N_16462);
nor U19401 (N_19401,N_15739,N_14364);
or U19402 (N_19402,N_14072,N_15315);
nand U19403 (N_19403,N_12305,N_16380);
and U19404 (N_19404,N_16983,N_14553);
nand U19405 (N_19405,N_16027,N_13543);
or U19406 (N_19406,N_12549,N_13051);
nor U19407 (N_19407,N_14816,N_14011);
nor U19408 (N_19408,N_12084,N_16734);
nor U19409 (N_19409,N_14161,N_12388);
xor U19410 (N_19410,N_14170,N_13671);
nor U19411 (N_19411,N_15141,N_15657);
xnor U19412 (N_19412,N_16262,N_16248);
and U19413 (N_19413,N_15607,N_13932);
nand U19414 (N_19414,N_13584,N_17688);
or U19415 (N_19415,N_15581,N_12521);
xor U19416 (N_19416,N_17822,N_13685);
xnor U19417 (N_19417,N_13785,N_16370);
xnor U19418 (N_19418,N_15377,N_12587);
xnor U19419 (N_19419,N_16485,N_14683);
and U19420 (N_19420,N_17551,N_12996);
or U19421 (N_19421,N_14420,N_17635);
or U19422 (N_19422,N_17870,N_12863);
and U19423 (N_19423,N_15083,N_17069);
xnor U19424 (N_19424,N_16563,N_15155);
xnor U19425 (N_19425,N_13868,N_12794);
nor U19426 (N_19426,N_17474,N_14452);
or U19427 (N_19427,N_16567,N_13801);
or U19428 (N_19428,N_12132,N_17481);
nand U19429 (N_19429,N_12731,N_16259);
nand U19430 (N_19430,N_16839,N_16710);
nand U19431 (N_19431,N_15347,N_16797);
xnor U19432 (N_19432,N_12222,N_17196);
xnor U19433 (N_19433,N_17786,N_13382);
nor U19434 (N_19434,N_13788,N_13698);
nand U19435 (N_19435,N_15661,N_17148);
nor U19436 (N_19436,N_17910,N_13464);
nor U19437 (N_19437,N_15828,N_12810);
xnor U19438 (N_19438,N_17279,N_13478);
and U19439 (N_19439,N_15111,N_15424);
nor U19440 (N_19440,N_15308,N_12505);
and U19441 (N_19441,N_16186,N_12562);
nor U19442 (N_19442,N_12824,N_14117);
or U19443 (N_19443,N_17996,N_12988);
or U19444 (N_19444,N_17890,N_13727);
nand U19445 (N_19445,N_14206,N_13853);
nor U19446 (N_19446,N_13322,N_15663);
xor U19447 (N_19447,N_16440,N_13511);
xor U19448 (N_19448,N_16350,N_12026);
nand U19449 (N_19449,N_15026,N_14441);
nor U19450 (N_19450,N_17282,N_15145);
and U19451 (N_19451,N_15206,N_15115);
and U19452 (N_19452,N_16726,N_14747);
or U19453 (N_19453,N_16860,N_13119);
or U19454 (N_19454,N_12158,N_17358);
or U19455 (N_19455,N_13107,N_12228);
or U19456 (N_19456,N_13568,N_15492);
or U19457 (N_19457,N_16749,N_16857);
nand U19458 (N_19458,N_17185,N_12961);
or U19459 (N_19459,N_14843,N_15159);
nand U19460 (N_19460,N_15556,N_13343);
nor U19461 (N_19461,N_13316,N_15366);
and U19462 (N_19462,N_16100,N_15654);
xnor U19463 (N_19463,N_16826,N_14572);
nor U19464 (N_19464,N_12758,N_14000);
xor U19465 (N_19465,N_14391,N_17966);
and U19466 (N_19466,N_13422,N_13420);
and U19467 (N_19467,N_15231,N_17549);
or U19468 (N_19468,N_13919,N_17393);
or U19469 (N_19469,N_17999,N_16246);
xnor U19470 (N_19470,N_17397,N_17377);
nand U19471 (N_19471,N_17395,N_14508);
xor U19472 (N_19472,N_14057,N_15358);
and U19473 (N_19473,N_16587,N_14772);
and U19474 (N_19474,N_14315,N_14077);
xor U19475 (N_19475,N_13716,N_13999);
and U19476 (N_19476,N_17181,N_16362);
xnor U19477 (N_19477,N_16088,N_14472);
xor U19478 (N_19478,N_12308,N_16591);
or U19479 (N_19479,N_15596,N_14724);
nor U19480 (N_19480,N_16223,N_15746);
nor U19481 (N_19481,N_17060,N_13089);
xor U19482 (N_19482,N_14413,N_17376);
or U19483 (N_19483,N_14613,N_12748);
xnor U19484 (N_19484,N_17624,N_15077);
xor U19485 (N_19485,N_17520,N_17743);
nor U19486 (N_19486,N_15991,N_14805);
and U19487 (N_19487,N_14782,N_16796);
and U19488 (N_19488,N_12995,N_15005);
and U19489 (N_19489,N_16111,N_15668);
nor U19490 (N_19490,N_17103,N_13756);
or U19491 (N_19491,N_14875,N_13474);
or U19492 (N_19492,N_14652,N_14579);
xor U19493 (N_19493,N_13187,N_17909);
nor U19494 (N_19494,N_13228,N_12450);
xnor U19495 (N_19495,N_16270,N_14267);
nor U19496 (N_19496,N_15425,N_15164);
xor U19497 (N_19497,N_16173,N_15384);
and U19498 (N_19498,N_14920,N_14950);
and U19499 (N_19499,N_17769,N_14158);
xor U19500 (N_19500,N_16145,N_14765);
and U19501 (N_19501,N_17888,N_13608);
nor U19502 (N_19502,N_15623,N_13272);
nor U19503 (N_19503,N_15631,N_16519);
nor U19504 (N_19504,N_12362,N_12541);
and U19505 (N_19505,N_17026,N_17566);
or U19506 (N_19506,N_12212,N_13615);
xor U19507 (N_19507,N_15415,N_16125);
xnor U19508 (N_19508,N_12704,N_16851);
nor U19509 (N_19509,N_16466,N_13290);
nor U19510 (N_19510,N_16827,N_14169);
nand U19511 (N_19511,N_12067,N_16938);
nand U19512 (N_19512,N_12826,N_13016);
and U19513 (N_19513,N_16916,N_14819);
nor U19514 (N_19514,N_12626,N_16062);
and U19515 (N_19515,N_15350,N_12045);
xnor U19516 (N_19516,N_12831,N_16643);
nand U19517 (N_19517,N_12577,N_16496);
nand U19518 (N_19518,N_16475,N_12974);
or U19519 (N_19519,N_14136,N_12942);
xor U19520 (N_19520,N_15025,N_13726);
nand U19521 (N_19521,N_12571,N_12199);
or U19522 (N_19522,N_12822,N_15147);
nand U19523 (N_19523,N_16720,N_12506);
nand U19524 (N_19524,N_16589,N_14140);
nor U19525 (N_19525,N_14166,N_12477);
nand U19526 (N_19526,N_14269,N_15496);
nand U19527 (N_19527,N_12941,N_12329);
nand U19528 (N_19528,N_14157,N_12697);
and U19529 (N_19529,N_16239,N_15965);
nand U19530 (N_19530,N_17044,N_12083);
nand U19531 (N_19531,N_17505,N_17889);
or U19532 (N_19532,N_17283,N_12652);
and U19533 (N_19533,N_17344,N_15473);
and U19534 (N_19534,N_12413,N_14634);
nand U19535 (N_19535,N_12284,N_15590);
xnor U19536 (N_19536,N_15388,N_17184);
or U19537 (N_19537,N_14425,N_13739);
or U19538 (N_19538,N_15928,N_14523);
nor U19539 (N_19539,N_16301,N_16455);
nor U19540 (N_19540,N_16993,N_13056);
nor U19541 (N_19541,N_16684,N_17580);
and U19542 (N_19542,N_14351,N_13982);
nand U19543 (N_19543,N_13760,N_12709);
xnor U19544 (N_19544,N_15930,N_15545);
xor U19545 (N_19545,N_14947,N_14901);
and U19546 (N_19546,N_17543,N_13921);
and U19547 (N_19547,N_13962,N_15649);
and U19548 (N_19548,N_14208,N_16161);
nor U19549 (N_19549,N_17518,N_17812);
xnor U19550 (N_19550,N_15227,N_13134);
or U19551 (N_19551,N_17576,N_16939);
and U19552 (N_19552,N_14338,N_16247);
or U19553 (N_19553,N_16008,N_15440);
nand U19554 (N_19554,N_16067,N_16313);
and U19555 (N_19555,N_16914,N_12047);
xnor U19556 (N_19556,N_13147,N_17270);
xor U19557 (N_19557,N_12236,N_15770);
xor U19558 (N_19558,N_12057,N_16197);
or U19559 (N_19559,N_13840,N_17078);
or U19560 (N_19560,N_14111,N_16037);
xor U19561 (N_19561,N_14670,N_12063);
xnor U19562 (N_19562,N_17739,N_17355);
and U19563 (N_19563,N_12339,N_17708);
xnor U19564 (N_19564,N_12801,N_12660);
or U19565 (N_19565,N_17949,N_17555);
nor U19566 (N_19566,N_13276,N_14439);
nand U19567 (N_19567,N_12105,N_16441);
nand U19568 (N_19568,N_17904,N_14021);
and U19569 (N_19569,N_16742,N_16770);
xor U19570 (N_19570,N_16467,N_15774);
xor U19571 (N_19571,N_15682,N_13421);
xor U19572 (N_19572,N_12215,N_12478);
and U19573 (N_19573,N_15434,N_17884);
xor U19574 (N_19574,N_16233,N_13302);
nor U19575 (N_19575,N_16992,N_14987);
nand U19576 (N_19576,N_15644,N_12273);
nand U19577 (N_19577,N_15888,N_14870);
and U19578 (N_19578,N_14329,N_14839);
or U19579 (N_19579,N_15788,N_14864);
or U19580 (N_19580,N_14408,N_14092);
nand U19581 (N_19581,N_13725,N_12560);
nor U19582 (N_19582,N_12498,N_17271);
or U19583 (N_19583,N_14562,N_12619);
nand U19584 (N_19584,N_17725,N_13783);
nor U19585 (N_19585,N_14910,N_12451);
or U19586 (N_19586,N_15286,N_12226);
nor U19587 (N_19587,N_16104,N_13947);
xor U19588 (N_19588,N_16424,N_17760);
xnor U19589 (N_19589,N_17455,N_15433);
nand U19590 (N_19590,N_16318,N_12563);
and U19591 (N_19591,N_16536,N_15365);
nand U19592 (N_19592,N_13529,N_15861);
or U19593 (N_19593,N_16998,N_17082);
nand U19594 (N_19594,N_13135,N_12456);
xnor U19595 (N_19595,N_14219,N_16112);
nand U19596 (N_19596,N_12333,N_16662);
and U19597 (N_19597,N_17755,N_13662);
xor U19598 (N_19598,N_15436,N_14781);
xor U19599 (N_19599,N_15709,N_12679);
xnor U19600 (N_19600,N_13460,N_17764);
nand U19601 (N_19601,N_12224,N_17131);
or U19602 (N_19602,N_15200,N_14330);
nor U19603 (N_19603,N_17297,N_15036);
or U19604 (N_19604,N_16572,N_13348);
and U19605 (N_19605,N_17039,N_17447);
nand U19606 (N_19606,N_13029,N_14128);
nand U19607 (N_19607,N_13090,N_14678);
nand U19608 (N_19608,N_17896,N_14130);
nor U19609 (N_19609,N_14036,N_12546);
xor U19610 (N_19610,N_14983,N_14744);
or U19611 (N_19611,N_14243,N_15775);
and U19612 (N_19612,N_13165,N_15953);
or U19613 (N_19613,N_13102,N_15854);
and U19614 (N_19614,N_15754,N_16727);
nand U19615 (N_19615,N_15521,N_12452);
nor U19616 (N_19616,N_14233,N_17683);
and U19617 (N_19617,N_16883,N_14846);
and U19618 (N_19618,N_16338,N_13986);
or U19619 (N_19619,N_14368,N_14121);
and U19620 (N_19620,N_14937,N_14114);
nand U19621 (N_19621,N_14071,N_17121);
nand U19622 (N_19622,N_15831,N_15399);
or U19623 (N_19623,N_12918,N_16115);
and U19624 (N_19624,N_14881,N_14867);
or U19625 (N_19625,N_14178,N_16542);
or U19626 (N_19626,N_17938,N_17859);
or U19627 (N_19627,N_15735,N_15291);
xor U19628 (N_19628,N_13367,N_14376);
xor U19629 (N_19629,N_15968,N_15482);
nand U19630 (N_19630,N_14663,N_14907);
and U19631 (N_19631,N_14037,N_16412);
or U19632 (N_19632,N_15153,N_15762);
nor U19633 (N_19633,N_17492,N_16461);
xnor U19634 (N_19634,N_16610,N_17234);
nand U19635 (N_19635,N_16213,N_14069);
or U19636 (N_19636,N_14287,N_12540);
nand U19637 (N_19637,N_14475,N_17036);
nor U19638 (N_19638,N_16140,N_17637);
nand U19639 (N_19639,N_12739,N_15188);
nand U19640 (N_19640,N_15027,N_17530);
nand U19641 (N_19641,N_14154,N_15466);
nor U19642 (N_19642,N_14321,N_16677);
nand U19643 (N_19643,N_14247,N_12710);
or U19644 (N_19644,N_16996,N_16159);
or U19645 (N_19645,N_14271,N_14825);
or U19646 (N_19646,N_12915,N_13387);
and U19647 (N_19647,N_16269,N_15647);
nor U19648 (N_19648,N_14936,N_13901);
nand U19649 (N_19649,N_13059,N_13865);
xnor U19650 (N_19650,N_16646,N_13673);
nand U19651 (N_19651,N_15051,N_13027);
and U19652 (N_19652,N_12186,N_14945);
and U19653 (N_19653,N_12101,N_14860);
and U19654 (N_19654,N_14710,N_13152);
or U19655 (N_19655,N_13300,N_14686);
and U19656 (N_19656,N_13504,N_16837);
and U19657 (N_19657,N_15004,N_14520);
nor U19658 (N_19658,N_14918,N_15598);
xnor U19659 (N_19659,N_15766,N_16674);
nor U19660 (N_19660,N_14042,N_13922);
nand U19661 (N_19661,N_12449,N_14132);
nand U19662 (N_19662,N_13012,N_15702);
xnor U19663 (N_19663,N_12599,N_13871);
and U19664 (N_19664,N_14972,N_13074);
or U19665 (N_19665,N_12346,N_15392);
nor U19666 (N_19666,N_14595,N_12002);
nand U19667 (N_19667,N_16766,N_17568);
nor U19668 (N_19668,N_12001,N_16002);
xor U19669 (N_19669,N_17351,N_17405);
xnor U19670 (N_19670,N_13406,N_16005);
nand U19671 (N_19671,N_14167,N_15509);
nand U19672 (N_19672,N_14948,N_14084);
xor U19673 (N_19673,N_17817,N_14029);
and U19674 (N_19674,N_14513,N_12146);
nor U19675 (N_19675,N_12150,N_14868);
xor U19676 (N_19676,N_13082,N_12046);
or U19677 (N_19677,N_17360,N_12985);
nor U19678 (N_19678,N_16592,N_14605);
or U19679 (N_19679,N_17267,N_14583);
xor U19680 (N_19680,N_12848,N_15875);
nand U19681 (N_19681,N_16614,N_17677);
nor U19682 (N_19682,N_15578,N_17608);
and U19683 (N_19683,N_12754,N_16925);
or U19684 (N_19684,N_17623,N_17556);
or U19685 (N_19685,N_12526,N_16459);
nand U19686 (N_19686,N_16004,N_14578);
or U19687 (N_19687,N_16600,N_12262);
xnor U19688 (N_19688,N_14168,N_13956);
xnor U19689 (N_19689,N_16627,N_12207);
nor U19690 (N_19690,N_16977,N_16559);
and U19691 (N_19691,N_13804,N_13370);
nand U19692 (N_19692,N_13635,N_13700);
and U19693 (N_19693,N_17777,N_13111);
xnor U19694 (N_19694,N_13067,N_17919);
nor U19695 (N_19695,N_12792,N_17052);
xnor U19696 (N_19696,N_13182,N_17390);
and U19697 (N_19697,N_17955,N_13169);
xor U19698 (N_19698,N_17074,N_14400);
nor U19699 (N_19699,N_14542,N_16055);
xor U19700 (N_19700,N_14196,N_12314);
nor U19701 (N_19701,N_17582,N_14392);
and U19702 (N_19702,N_12250,N_15454);
nand U19703 (N_19703,N_14010,N_15560);
or U19704 (N_19704,N_14480,N_17288);
xnor U19705 (N_19705,N_14644,N_17601);
nor U19706 (N_19706,N_15274,N_13929);
nand U19707 (N_19707,N_17625,N_14808);
and U19708 (N_19708,N_17617,N_14242);
nor U19709 (N_19709,N_12444,N_16630);
xnor U19710 (N_19710,N_12736,N_16472);
and U19711 (N_19711,N_15070,N_13354);
xor U19712 (N_19712,N_16540,N_13692);
xor U19713 (N_19713,N_15859,N_14403);
nor U19714 (N_19714,N_14998,N_17927);
or U19715 (N_19715,N_13928,N_12159);
and U19716 (N_19716,N_16751,N_17010);
or U19717 (N_19717,N_15310,N_16961);
xnor U19718 (N_19718,N_13141,N_17258);
nor U19719 (N_19719,N_15107,N_16556);
nor U19720 (N_19720,N_17111,N_16568);
and U19721 (N_19721,N_15753,N_16945);
nor U19722 (N_19722,N_16631,N_14656);
xor U19723 (N_19723,N_13740,N_17340);
or U19724 (N_19724,N_15394,N_14304);
xnor U19725 (N_19725,N_15251,N_13213);
or U19726 (N_19726,N_13733,N_14142);
xor U19727 (N_19727,N_17592,N_16825);
nand U19728 (N_19728,N_16692,N_14817);
and U19729 (N_19729,N_12979,N_14278);
nand U19730 (N_19730,N_16581,N_12415);
or U19731 (N_19731,N_13515,N_16337);
nor U19732 (N_19732,N_16534,N_16767);
nand U19733 (N_19733,N_12113,N_14512);
nor U19734 (N_19734,N_14778,N_14097);
xor U19735 (N_19735,N_13020,N_14638);
or U19736 (N_19736,N_16935,N_14567);
nor U19737 (N_19737,N_16645,N_12365);
xnor U19738 (N_19738,N_14962,N_16622);
and U19739 (N_19739,N_13566,N_14904);
xor U19740 (N_19740,N_16632,N_15728);
xnor U19741 (N_19741,N_15012,N_17718);
nand U19742 (N_19742,N_16113,N_16870);
or U19743 (N_19743,N_17604,N_14073);
xnor U19744 (N_19744,N_12463,N_17333);
nand U19745 (N_19745,N_15014,N_16527);
xor U19746 (N_19746,N_14641,N_13463);
or U19747 (N_19747,N_17374,N_15508);
nand U19748 (N_19748,N_15094,N_15535);
and U19749 (N_19749,N_12257,N_15016);
or U19750 (N_19750,N_15074,N_12759);
nand U19751 (N_19751,N_13862,N_15241);
or U19752 (N_19752,N_15154,N_16014);
and U19753 (N_19753,N_16203,N_16413);
xnor U19754 (N_19754,N_14880,N_17029);
xnor U19755 (N_19755,N_12935,N_15086);
nand U19756 (N_19756,N_14929,N_17727);
nor U19757 (N_19757,N_14890,N_14616);
nor U19758 (N_19758,N_15461,N_13308);
nor U19759 (N_19759,N_12087,N_12433);
xnor U19760 (N_19760,N_14139,N_12420);
and U19761 (N_19761,N_16583,N_14786);
nand U19762 (N_19762,N_16444,N_12326);
and U19763 (N_19763,N_17906,N_16753);
nor U19764 (N_19764,N_15555,N_14334);
nand U19765 (N_19765,N_16437,N_14125);
and U19766 (N_19766,N_17902,N_16118);
and U19767 (N_19767,N_13891,N_12018);
or U19768 (N_19768,N_16128,N_16474);
nor U19769 (N_19769,N_13572,N_15909);
nand U19770 (N_19770,N_13618,N_15216);
and U19771 (N_19771,N_14788,N_13889);
nand U19772 (N_19772,N_12050,N_13691);
nand U19773 (N_19773,N_12727,N_17535);
xor U19774 (N_19774,N_14034,N_15794);
and U19775 (N_19775,N_16003,N_17081);
and U19776 (N_19776,N_15563,N_17523);
or U19777 (N_19777,N_14630,N_13524);
nor U19778 (N_19778,N_12561,N_17266);
nand U19779 (N_19779,N_13252,N_16367);
and U19780 (N_19780,N_14418,N_13887);
and U19781 (N_19781,N_13627,N_15632);
nor U19782 (N_19782,N_13206,N_17780);
xnor U19783 (N_19783,N_15704,N_15876);
nor U19784 (N_19784,N_15346,N_17466);
nor U19785 (N_19785,N_12356,N_15451);
nor U19786 (N_19786,N_15625,N_16871);
or U19787 (N_19787,N_16083,N_16654);
nand U19788 (N_19788,N_12947,N_13843);
nand U19789 (N_19789,N_16515,N_15289);
nand U19790 (N_19790,N_17410,N_16975);
nor U19791 (N_19791,N_14606,N_12188);
and U19792 (N_19792,N_17408,N_16701);
or U19793 (N_19793,N_16410,N_12926);
nand U19794 (N_19794,N_13550,N_15898);
or U19795 (N_19795,N_14753,N_16207);
xor U19796 (N_19796,N_17998,N_15174);
xnor U19797 (N_19797,N_17758,N_17067);
nand U19798 (N_19798,N_14289,N_17893);
nor U19799 (N_19799,N_17640,N_16603);
nand U19800 (N_19800,N_13179,N_15824);
xor U19801 (N_19801,N_12283,N_16917);
nand U19802 (N_19802,N_12833,N_17445);
nand U19803 (N_19803,N_15169,N_12482);
nor U19804 (N_19804,N_12896,N_14695);
or U19805 (N_19805,N_17239,N_12573);
xnor U19806 (N_19806,N_12403,N_16625);
nand U19807 (N_19807,N_14366,N_15184);
nor U19808 (N_19808,N_14884,N_17276);
or U19809 (N_19809,N_12145,N_14133);
nand U19810 (N_19810,N_17546,N_12321);
xnor U19811 (N_19811,N_17305,N_14569);
or U19812 (N_19812,N_14685,N_14200);
and U19813 (N_19813,N_13415,N_15867);
or U19814 (N_19814,N_16921,N_17208);
nand U19815 (N_19815,N_13324,N_12360);
and U19816 (N_19816,N_13227,N_15166);
nor U19817 (N_19817,N_17322,N_15177);
nand U19818 (N_19818,N_13506,N_15072);
xnor U19819 (N_19819,N_14535,N_14086);
or U19820 (N_19820,N_14774,N_12299);
xnor U19821 (N_19821,N_15684,N_14637);
and U19822 (N_19822,N_14544,N_14106);
xnor U19823 (N_19823,N_14558,N_16098);
xor U19824 (N_19824,N_15757,N_15700);
and U19825 (N_19825,N_15927,N_17946);
nor U19826 (N_19826,N_15334,N_13400);
xor U19827 (N_19827,N_13368,N_16985);
nand U19828 (N_19828,N_16238,N_16689);
nor U19829 (N_19829,N_14969,N_15450);
and U19830 (N_19830,N_16001,N_16322);
nand U19831 (N_19831,N_12981,N_17230);
xor U19832 (N_19832,N_14770,N_14466);
or U19833 (N_19833,N_16876,N_12078);
nand U19834 (N_19834,N_12072,N_13117);
nand U19835 (N_19835,N_14522,N_17180);
xor U19836 (N_19836,N_13631,N_12551);
or U19837 (N_19837,N_13552,N_16863);
and U19838 (N_19838,N_12320,N_16728);
nor U19839 (N_19839,N_16095,N_14113);
or U19840 (N_19840,N_13257,N_14551);
and U19841 (N_19841,N_15401,N_15924);
or U19842 (N_19842,N_17579,N_15438);
and U19843 (N_19843,N_14627,N_12671);
or U19844 (N_19844,N_16541,N_16034);
nor U19845 (N_19845,N_15841,N_13168);
xor U19846 (N_19846,N_14095,N_13902);
xnor U19847 (N_19847,N_13858,N_16087);
nand U19848 (N_19848,N_16493,N_12873);
nand U19849 (N_19849,N_14320,N_12845);
nor U19850 (N_19850,N_14866,N_13670);
and U19851 (N_19851,N_13489,N_17443);
and U19852 (N_19852,N_14002,N_13701);
xor U19853 (N_19853,N_13742,N_14290);
xor U19854 (N_19854,N_17193,N_14874);
and U19855 (N_19855,N_12327,N_12788);
nor U19856 (N_19856,N_17129,N_16052);
xnor U19857 (N_19857,N_12811,N_13682);
or U19858 (N_19858,N_14171,N_16268);
or U19859 (N_19859,N_16942,N_13350);
xor U19860 (N_19860,N_13479,N_12738);
or U19861 (N_19861,N_16276,N_15678);
nand U19862 (N_19862,N_16219,N_13149);
nand U19863 (N_19863,N_15730,N_16982);
and U19864 (N_19864,N_13081,N_17987);
or U19865 (N_19865,N_12022,N_13154);
or U19866 (N_19866,N_16609,N_14862);
xnor U19867 (N_19867,N_14728,N_15119);
and U19868 (N_19868,N_17658,N_14361);
xor U19869 (N_19869,N_17554,N_12255);
xor U19870 (N_19870,N_14658,N_15480);
and U19871 (N_19871,N_16729,N_15201);
or U19872 (N_19872,N_14536,N_13905);
xor U19873 (N_19873,N_13260,N_17100);
nand U19874 (N_19874,N_13717,N_13336);
and U19875 (N_19875,N_16969,N_15864);
or U19876 (N_19876,N_12225,N_14456);
and U19877 (N_19877,N_17652,N_13036);
and U19878 (N_19878,N_15699,N_15396);
or U19879 (N_19879,N_12904,N_13106);
nor U19880 (N_19880,N_17401,N_16311);
and U19881 (N_19881,N_14448,N_12421);
xnor U19882 (N_19882,N_15021,N_14151);
or U19883 (N_19883,N_13579,N_13749);
or U19884 (N_19884,N_17976,N_14623);
and U19885 (N_19885,N_12104,N_13277);
or U19886 (N_19886,N_15805,N_16297);
xor U19887 (N_19887,N_14291,N_14855);
nand U19888 (N_19888,N_17312,N_13678);
xor U19889 (N_19889,N_16649,N_17307);
nand U19890 (N_19890,N_13378,N_17703);
nand U19891 (N_19891,N_14924,N_14455);
and U19892 (N_19892,N_16495,N_13409);
nor U19893 (N_19893,N_15405,N_16514);
xnor U19894 (N_19894,N_17811,N_12982);
nor U19895 (N_19895,N_15686,N_17578);
nor U19896 (N_19896,N_13876,N_13253);
and U19897 (N_19897,N_13219,N_12690);
nor U19898 (N_19898,N_14682,N_12657);
or U19899 (N_19899,N_15561,N_12631);
nand U19900 (N_19900,N_15387,N_17790);
nand U19901 (N_19901,N_15089,N_17012);
nor U19902 (N_19902,N_16763,N_12277);
nor U19903 (N_19903,N_13606,N_15108);
xnor U19904 (N_19904,N_17874,N_13896);
or U19905 (N_19905,N_17291,N_12643);
nor U19906 (N_19906,N_13032,N_12396);
xor U19907 (N_19907,N_17673,N_16388);
nand U19908 (N_19908,N_15769,N_12632);
nand U19909 (N_19909,N_13851,N_17225);
and U19910 (N_19910,N_12566,N_13628);
nand U19911 (N_19911,N_12134,N_13666);
or U19912 (N_19912,N_13462,N_12968);
nor U19913 (N_19913,N_17663,N_14959);
nor U19914 (N_19914,N_12867,N_16224);
and U19915 (N_19915,N_15897,N_14027);
nand U19916 (N_19916,N_13767,N_13998);
nor U19917 (N_19917,N_12467,N_12946);
or U19918 (N_19918,N_17118,N_16325);
xnor U19919 (N_19919,N_17359,N_15977);
or U19920 (N_19920,N_16076,N_13656);
nand U19921 (N_19921,N_14736,N_15767);
nand U19922 (N_19922,N_17948,N_14643);
nor U19923 (N_19923,N_15642,N_14191);
or U19924 (N_19924,N_12238,N_16611);
xor U19925 (N_19925,N_13457,N_13991);
nor U19926 (N_19926,N_13417,N_16226);
or U19927 (N_19927,N_12522,N_15949);
xnor U19928 (N_19928,N_16877,N_17223);
xor U19929 (N_19929,N_13548,N_13620);
or U19930 (N_19930,N_14045,N_12839);
and U19931 (N_19931,N_16178,N_16732);
nand U19932 (N_19932,N_13040,N_16518);
and U19933 (N_19933,N_17105,N_17240);
nor U19934 (N_19934,N_12596,N_16304);
or U19935 (N_19935,N_12929,N_13658);
or U19936 (N_19936,N_14471,N_16667);
or U19937 (N_19937,N_12316,N_13557);
or U19938 (N_19938,N_17993,N_15449);
nand U19939 (N_19939,N_12556,N_15132);
nor U19940 (N_19940,N_13651,N_16578);
and U19941 (N_19941,N_16892,N_16944);
and U19942 (N_19942,N_12304,N_15653);
nor U19943 (N_19943,N_13312,N_12342);
and U19944 (N_19944,N_13118,N_16300);
or U19945 (N_19945,N_13774,N_14596);
and U19946 (N_19946,N_13143,N_14384);
nand U19947 (N_19947,N_16150,N_14722);
and U19948 (N_19948,N_15850,N_13418);
and U19949 (N_19949,N_16179,N_12061);
xor U19950 (N_19950,N_17079,N_13271);
and U19951 (N_19951,N_17367,N_12102);
and U19952 (N_19952,N_12382,N_17486);
nand U19953 (N_19953,N_16607,N_16832);
or U19954 (N_19954,N_13172,N_14894);
nand U19955 (N_19955,N_17194,N_15493);
and U19956 (N_19956,N_17253,N_13718);
and U19957 (N_19957,N_14537,N_13281);
xnor U19958 (N_19958,N_13789,N_12764);
xor U19959 (N_19959,N_13978,N_14506);
and U19960 (N_19960,N_14826,N_14599);
xor U19961 (N_19961,N_12624,N_16821);
nand U19962 (N_19962,N_17650,N_13018);
nand U19963 (N_19963,N_15002,N_16120);
nor U19964 (N_19964,N_17931,N_12603);
xnor U19965 (N_19965,N_17960,N_14495);
and U19966 (N_19966,N_17824,N_13567);
xor U19967 (N_19967,N_12648,N_16166);
or U19968 (N_19968,N_12503,N_14431);
nand U19969 (N_19969,N_17197,N_12155);
xnor U19970 (N_19970,N_16264,N_16041);
xnor U19971 (N_19971,N_16368,N_12419);
nor U19972 (N_19972,N_16713,N_15501);
and U19973 (N_19973,N_15063,N_13180);
and U19974 (N_19974,N_15559,N_16174);
nor U19975 (N_19975,N_12015,N_15211);
nand U19976 (N_19976,N_13301,N_12073);
nor U19977 (N_19977,N_15634,N_17689);
nand U19978 (N_19978,N_17513,N_13092);
or U19979 (N_19979,N_15890,N_12039);
xor U19980 (N_19980,N_15491,N_13818);
nand U19981 (N_19981,N_14885,N_15781);
xor U19982 (N_19982,N_13654,N_16498);
xnor U19983 (N_19983,N_13894,N_13831);
xnor U19984 (N_19984,N_15418,N_15176);
nand U19985 (N_19985,N_17483,N_14759);
nor U19986 (N_19986,N_14094,N_15099);
nor U19987 (N_19987,N_12297,N_15743);
nand U19988 (N_19988,N_13017,N_13545);
or U19989 (N_19989,N_15652,N_16009);
xnor U19990 (N_19990,N_17037,N_16521);
and U19991 (N_19991,N_14244,N_12707);
or U19992 (N_19992,N_13428,N_13004);
nand U19993 (N_19993,N_12852,N_17264);
nor U19994 (N_19994,N_16182,N_12532);
and U19995 (N_19995,N_17875,N_14090);
nand U19996 (N_19996,N_14061,N_15306);
or U19997 (N_19997,N_15023,N_12170);
or U19998 (N_19998,N_13826,N_14858);
or U19999 (N_19999,N_14944,N_17409);
xnor U20000 (N_20000,N_13707,N_15800);
and U20001 (N_20001,N_16897,N_13838);
xor U20002 (N_20002,N_12814,N_13232);
nand U20003 (N_20003,N_12809,N_17189);
or U20004 (N_20004,N_16629,N_15587);
xnor U20005 (N_20005,N_15896,N_13208);
nand U20006 (N_20006,N_14081,N_17319);
nand U20007 (N_20007,N_16222,N_17165);
xnor U20008 (N_20008,N_16535,N_14785);
xor U20009 (N_20009,N_14879,N_12776);
xor U20010 (N_20010,N_12518,N_15148);
or U20011 (N_20011,N_15671,N_15804);
and U20012 (N_20012,N_14332,N_13218);
or U20013 (N_20013,N_15765,N_17051);
nor U20014 (N_20014,N_14083,N_16200);
and U20015 (N_20015,N_17146,N_17252);
nor U20016 (N_20016,N_14326,N_17337);
nor U20017 (N_20017,N_15460,N_14979);
nand U20018 (N_20018,N_15467,N_13293);
nor U20019 (N_20019,N_12016,N_13578);
xor U20020 (N_20020,N_14282,N_13600);
and U20021 (N_20021,N_16487,N_15920);
xor U20022 (N_20022,N_16214,N_15279);
nor U20023 (N_20023,N_17905,N_17017);
or U20024 (N_20024,N_17958,N_17710);
and U20025 (N_20025,N_16769,N_17373);
nor U20026 (N_20026,N_15283,N_12617);
nor U20027 (N_20027,N_17281,N_12675);
nand U20028 (N_20028,N_17090,N_15817);
nand U20029 (N_20029,N_14396,N_15272);
or U20030 (N_20030,N_15749,N_13503);
nor U20031 (N_20031,N_16221,N_17785);
nor U20032 (N_20032,N_15092,N_15524);
and U20033 (N_20033,N_16688,N_16793);
nor U20034 (N_20034,N_14624,N_16791);
or U20035 (N_20035,N_12157,N_15612);
xor U20036 (N_20036,N_14105,N_17187);
nor U20037 (N_20037,N_13607,N_17598);
or U20038 (N_20038,N_15764,N_16829);
and U20039 (N_20039,N_14566,N_13372);
and U20040 (N_20040,N_17577,N_17338);
xnor U20041 (N_20041,N_14372,N_13062);
or U20042 (N_20042,N_13448,N_16570);
and U20043 (N_20043,N_15763,N_15340);
and U20044 (N_20044,N_17163,N_13238);
xor U20045 (N_20045,N_12870,N_17182);
and U20046 (N_20046,N_13174,N_13996);
nand U20047 (N_20047,N_14932,N_16309);
xor U20048 (N_20048,N_16205,N_12053);
and U20049 (N_20049,N_14479,N_16295);
xor U20050 (N_20050,N_12698,N_12358);
xnor U20051 (N_20051,N_13644,N_12681);
xor U20052 (N_20052,N_15673,N_16577);
xor U20053 (N_20053,N_16048,N_14568);
xnor U20054 (N_20054,N_16973,N_14891);
and U20055 (N_20055,N_12545,N_16838);
xor U20056 (N_20056,N_16676,N_16422);
xor U20057 (N_20057,N_15052,N_17246);
or U20058 (N_20058,N_14675,N_14476);
or U20059 (N_20059,N_14126,N_15514);
and U20060 (N_20060,N_17458,N_13196);
xor U20061 (N_20061,N_12031,N_13230);
xnor U20062 (N_20062,N_17471,N_15872);
xor U20063 (N_20063,N_16294,N_14966);
nand U20064 (N_20064,N_17001,N_13451);
or U20065 (N_20065,N_13645,N_17712);
and U20066 (N_20066,N_14473,N_13432);
nand U20067 (N_20067,N_15790,N_16530);
and U20068 (N_20068,N_12992,N_16974);
and U20069 (N_20069,N_17842,N_17980);
nor U20070 (N_20070,N_16545,N_12249);
xor U20071 (N_20071,N_14022,N_12343);
nor U20072 (N_20072,N_15963,N_15091);
or U20073 (N_20073,N_12100,N_16952);
xor U20074 (N_20074,N_12296,N_17648);
nor U20075 (N_20075,N_15626,N_14546);
nor U20076 (N_20076,N_13663,N_15323);
xnor U20077 (N_20077,N_14589,N_15295);
and U20078 (N_20078,N_13037,N_13547);
or U20079 (N_20079,N_15407,N_12891);
nor U20080 (N_20080,N_13459,N_16681);
and U20081 (N_20081,N_13872,N_16066);
xor U20082 (N_20082,N_13660,N_12117);
and U20083 (N_20083,N_16327,N_14509);
nand U20084 (N_20084,N_17851,N_17213);
or U20085 (N_20085,N_12984,N_14451);
xnor U20086 (N_20086,N_15780,N_16906);
or U20087 (N_20087,N_13973,N_12232);
nor U20088 (N_20088,N_16595,N_12516);
or U20089 (N_20089,N_15591,N_17581);
or U20090 (N_20090,N_15006,N_14078);
and U20091 (N_20091,N_12659,N_15443);
nand U20092 (N_20092,N_15294,N_16759);
nand U20093 (N_20093,N_15085,N_12774);
nand U20094 (N_20094,N_13339,N_16525);
xor U20095 (N_20095,N_13711,N_12616);
and U20096 (N_20096,N_13347,N_15321);
or U20097 (N_20097,N_16414,N_15045);
nor U20098 (N_20098,N_14355,N_13861);
nand U20099 (N_20099,N_14561,N_14262);
or U20100 (N_20100,N_16748,N_14514);
or U20101 (N_20101,N_16795,N_15034);
nand U20102 (N_20102,N_14841,N_15548);
and U20103 (N_20103,N_16941,N_12620);
or U20104 (N_20104,N_13058,N_13555);
nand U20105 (N_20105,N_13799,N_13371);
nand U20106 (N_20106,N_14490,N_14202);
or U20107 (N_20107,N_13893,N_12156);
or U20108 (N_20108,N_12041,N_12610);
or U20109 (N_20109,N_17042,N_14059);
xnor U20110 (N_20110,N_12976,N_14994);
xnor U20111 (N_20111,N_14721,N_14554);
and U20112 (N_20112,N_17203,N_17749);
xor U20113 (N_20113,N_14847,N_15196);
xnor U20114 (N_20114,N_15954,N_14383);
xnor U20115 (N_20115,N_12118,N_15054);
or U20116 (N_20116,N_17922,N_16478);
nor U20117 (N_20117,N_13683,N_12377);
and U20118 (N_20118,N_15731,N_12495);
nor U20119 (N_20119,N_15446,N_12331);
nand U20120 (N_20120,N_15373,N_12291);
xor U20121 (N_20121,N_12539,N_17541);
nand U20122 (N_20122,N_15222,N_13811);
and U20123 (N_20123,N_17034,N_12140);
nand U20124 (N_20124,N_16947,N_13977);
nor U20125 (N_20125,N_15619,N_16250);
and U20126 (N_20126,N_14134,N_13164);
xnor U20127 (N_20127,N_12148,N_17011);
xor U20128 (N_20128,N_15250,N_17339);
nor U20129 (N_20129,N_13026,N_14655);
nor U20130 (N_20130,N_12349,N_15053);
nor U20131 (N_20131,N_13588,N_16943);
and U20132 (N_20132,N_17503,N_17796);
xnor U20133 (N_20133,N_14761,N_12120);
nand U20134 (N_20134,N_15060,N_16377);
xor U20135 (N_20135,N_12800,N_13243);
nand U20136 (N_20136,N_14482,N_17916);
and U20137 (N_20137,N_15179,N_13863);
xnor U20138 (N_20138,N_16481,N_17511);
nor U20139 (N_20139,N_14883,N_15214);
nand U20140 (N_20140,N_16305,N_17547);
nor U20141 (N_20141,N_12181,N_12364);
nor U20142 (N_20142,N_17053,N_14212);
and U20143 (N_20143,N_13719,N_17040);
xor U20144 (N_20144,N_16074,N_13960);
nor U20145 (N_20145,N_14614,N_17108);
or U20146 (N_20146,N_12380,N_17412);
xor U20147 (N_20147,N_16180,N_12760);
or U20148 (N_20148,N_16908,N_12033);
or U20149 (N_20149,N_15124,N_16330);
nand U20150 (N_20150,N_14350,N_17985);
nand U20151 (N_20151,N_12080,N_14474);
and U20152 (N_20152,N_14486,N_16959);
xor U20153 (N_20153,N_16283,N_15693);
or U20154 (N_20154,N_14964,N_16762);
or U20155 (N_20155,N_17192,N_13583);
and U20156 (N_20156,N_12069,N_15773);
nand U20157 (N_20157,N_17170,N_16183);
or U20158 (N_20158,N_16718,N_14230);
nand U20159 (N_20159,N_13959,N_12122);
nor U20160 (N_20160,N_13259,N_12567);
nor U20161 (N_20161,N_14398,N_14131);
and U20162 (N_20162,N_17490,N_16366);
and U20163 (N_20163,N_16429,N_14453);
xor U20164 (N_20164,N_17470,N_17023);
nand U20165 (N_20165,N_12253,N_12888);
or U20166 (N_20166,N_12892,N_12994);
nor U20167 (N_20167,N_13133,N_15344);
xnor U20168 (N_20168,N_16840,N_16835);
nand U20169 (N_20169,N_17587,N_12689);
xnor U20170 (N_20170,N_14345,N_17524);
nor U20171 (N_20171,N_17781,N_17691);
and U20172 (N_20172,N_13604,N_15452);
and U20173 (N_20173,N_14183,N_17482);
nor U20174 (N_20174,N_15688,N_17611);
nand U20175 (N_20175,N_14358,N_12465);
nand U20176 (N_20176,N_12630,N_13527);
or U20177 (N_20177,N_16923,N_14146);
nand U20178 (N_20178,N_14160,N_16425);
nor U20179 (N_20179,N_17885,N_14385);
or U20180 (N_20180,N_13908,N_12534);
xor U20181 (N_20181,N_17316,N_12898);
nor U20182 (N_20182,N_17475,N_15391);
nand U20183 (N_20183,N_15602,N_13419);
nand U20184 (N_20184,N_14265,N_12538);
nor U20185 (N_20185,N_17517,N_13931);
or U20186 (N_20186,N_17565,N_12006);
nand U20187 (N_20187,N_12425,N_13821);
xor U20188 (N_20188,N_16955,N_16599);
nor U20189 (N_20189,N_12234,N_13859);
xnor U20190 (N_20190,N_16286,N_16420);
nand U20191 (N_20191,N_15736,N_15118);
and U20192 (N_20192,N_13384,N_16010);
nor U20193 (N_20193,N_13816,N_14556);
nor U20194 (N_20194,N_12335,N_14281);
and U20195 (N_20195,N_14688,N_13404);
xnor U20196 (N_20196,N_15465,N_17031);
xor U20197 (N_20197,N_17251,N_16308);
nand U20198 (N_20198,N_13624,N_15915);
xor U20199 (N_20199,N_16400,N_14703);
xor U20200 (N_20200,N_13331,N_13125);
nand U20201 (N_20201,N_15349,N_16417);
and U20202 (N_20202,N_15003,N_15192);
and U20203 (N_20203,N_17112,N_13724);
nor U20204 (N_20204,N_12223,N_15500);
nand U20205 (N_20205,N_16458,N_14460);
and U20206 (N_20206,N_14240,N_16850);
and U20207 (N_20207,N_13559,N_12907);
or U20208 (N_20208,N_15037,N_16683);
nor U20209 (N_20209,N_15839,N_12720);
xor U20210 (N_20210,N_14809,N_13146);
and U20211 (N_20211,N_15125,N_16110);
nand U20212 (N_20212,N_12309,N_13183);
or U20213 (N_20213,N_14840,N_14100);
and U20214 (N_20214,N_15459,N_13153);
and U20215 (N_20215,N_12246,N_16017);
xor U20216 (N_20216,N_12160,N_12030);
nand U20217 (N_20217,N_13910,N_13909);
nor U20218 (N_20218,N_12803,N_14577);
or U20219 (N_20219,N_13214,N_15429);
or U20220 (N_20220,N_13953,N_13468);
nor U20221 (N_20221,N_13162,N_17793);
and U20222 (N_20222,N_17575,N_16948);
xor U20223 (N_20223,N_15858,N_15860);
nor U20224 (N_20224,N_13537,N_12353);
and U20225 (N_20225,N_14481,N_15444);
and U20226 (N_20226,N_13748,N_13827);
or U20227 (N_20227,N_12564,N_15620);
xnor U20228 (N_20228,N_15258,N_16792);
nor U20229 (N_20229,N_15708,N_14357);
nor U20230 (N_20230,N_12746,N_14780);
nand U20231 (N_20231,N_17838,N_16548);
or U20232 (N_20232,N_14261,N_13765);
nand U20233 (N_20233,N_17178,N_12855);
nor U20234 (N_20234,N_16317,N_16549);
and U20235 (N_20235,N_14040,N_13585);
and U20236 (N_20236,N_15586,N_16409);
nand U20237 (N_20237,N_14340,N_16315);
nand U20238 (N_20238,N_16569,N_12123);
and U20239 (N_20239,N_17244,N_17850);
and U20240 (N_20240,N_14483,N_12357);
nand U20241 (N_20241,N_14299,N_16844);
or U20242 (N_20242,N_16705,N_17597);
nor U20243 (N_20243,N_14309,N_13852);
xnor U20244 (N_20244,N_13516,N_16093);
xor U20245 (N_20245,N_16480,N_16158);
or U20246 (N_20246,N_12823,N_15972);
nor U20247 (N_20247,N_15813,N_13292);
and U20248 (N_20248,N_13345,N_16319);
nand U20249 (N_20249,N_12805,N_14001);
nand U20250 (N_20250,N_14149,N_17462);
or U20251 (N_20251,N_15884,N_12325);
xor U20252 (N_20252,N_14995,N_16361);
nand U20253 (N_20253,N_17491,N_17499);
or U20254 (N_20254,N_12280,N_15667);
nor U20255 (N_20255,N_17199,N_12790);
nor U20256 (N_20256,N_12691,N_12034);
or U20257 (N_20257,N_14978,N_14731);
and U20258 (N_20258,N_17961,N_17848);
xor U20259 (N_20259,N_16582,N_14636);
xor U20260 (N_20260,N_12455,N_14672);
or U20261 (N_20261,N_15666,N_14836);
nand U20262 (N_20262,N_14938,N_16784);
nor U20263 (N_20263,N_14526,N_16765);
xor U20264 (N_20264,N_17538,N_15485);
or U20265 (N_20265,N_17583,N_15411);
or U20266 (N_20266,N_14503,N_17865);
or U20267 (N_20267,N_12753,N_12029);
xnor U20268 (N_20268,N_16356,N_14869);
nor U20269 (N_20269,N_16057,N_17534);
nor U20270 (N_20270,N_15134,N_15270);
xnor U20271 (N_20271,N_14970,N_16620);
nand U20272 (N_20272,N_15593,N_13078);
nor U20273 (N_20273,N_13112,N_15029);
nand U20274 (N_20274,N_15223,N_15312);
nor U20275 (N_20275,N_17098,N_12906);
nand U20276 (N_20276,N_16664,N_15484);
nand U20277 (N_20277,N_17419,N_14588);
xnor U20278 (N_20278,N_13352,N_17043);
xor U20279 (N_20279,N_14750,N_13558);
nor U20280 (N_20280,N_14423,N_17369);
and U20281 (N_20281,N_14032,N_12500);
or U20282 (N_20282,N_13145,N_14303);
and U20283 (N_20283,N_12056,N_14404);
nand U20284 (N_20284,N_13144,N_17168);
xor U20285 (N_20285,N_15309,N_13564);
and U20286 (N_20286,N_17294,N_17022);
xor U20287 (N_20287,N_16069,N_12640);
xor U20288 (N_20288,N_13528,N_13251);
or U20289 (N_20289,N_14129,N_15615);
nor U20290 (N_20290,N_16820,N_16401);
nor U20291 (N_20291,N_16138,N_17433);
and U20292 (N_20292,N_15681,N_17091);
and U20293 (N_20293,N_17818,N_13714);
xnor U20294 (N_20294,N_17670,N_16721);
nand U20295 (N_20295,N_12312,N_13825);
xnor U20296 (N_20296,N_12779,N_16494);
nand U20297 (N_20297,N_15110,N_12390);
nand U20298 (N_20298,N_12151,N_12747);
xnor U20299 (N_20299,N_15471,N_13176);
xnor U20300 (N_20300,N_17489,N_13551);
xor U20301 (N_20301,N_13193,N_13935);
nand U20302 (N_20302,N_16470,N_14631);
or U20303 (N_20303,N_14773,N_17354);
or U20304 (N_20304,N_16482,N_15998);
xor U20305 (N_20305,N_13731,N_15938);
or U20306 (N_20306,N_14828,N_17454);
or U20307 (N_20307,N_15857,N_12276);
xnor U20308 (N_20308,N_15511,N_17025);
nor U20309 (N_20309,N_15024,N_14312);
nand U20310 (N_20310,N_15838,N_14307);
and U20311 (N_20311,N_14690,N_16539);
or U20312 (N_20312,N_12302,N_12533);
xnor U20313 (N_20313,N_12899,N_16971);
xnor U20314 (N_20314,N_14359,N_14653);
nand U20315 (N_20315,N_14020,N_15343);
or U20316 (N_20316,N_13834,N_16167);
and U20317 (N_20317,N_12119,N_17206);
nand U20318 (N_20318,N_12909,N_15048);
nand U20319 (N_20319,N_12248,N_12074);
and U20320 (N_20320,N_15088,N_16334);
or U20321 (N_20321,N_15368,N_13099);
nor U20322 (N_20322,N_15175,N_16546);
or U20323 (N_20323,N_12592,N_17863);
nor U20324 (N_20324,N_13920,N_14342);
or U20325 (N_20325,N_12550,N_16618);
nand U20326 (N_20326,N_13681,N_12152);
and U20327 (N_20327,N_15084,N_15891);
and U20328 (N_20328,N_16506,N_15613);
nor U20329 (N_20329,N_12129,N_17869);
nand U20330 (N_20330,N_17300,N_12827);
or U20331 (N_20331,N_15146,N_13003);
or U20332 (N_20332,N_16374,N_12355);
nand U20333 (N_20333,N_12089,N_12021);
xnor U20334 (N_20334,N_16099,N_12807);
nand U20335 (N_20335,N_14716,N_14908);
nand U20336 (N_20336,N_12090,N_12512);
nor U20337 (N_20337,N_13351,N_15579);
xor U20338 (N_20338,N_17432,N_16640);
xor U20339 (N_20339,N_12372,N_16229);
or U20340 (N_20340,N_13231,N_14751);
nor U20341 (N_20341,N_12434,N_16859);
nor U20342 (N_20342,N_16351,N_13079);
or U20343 (N_20343,N_16638,N_16818);
nor U20344 (N_20344,N_16023,N_15182);
nand U20345 (N_20345,N_13830,N_12383);
nand U20346 (N_20346,N_15873,N_16557);
nor U20347 (N_20347,N_12829,N_17451);
nand U20348 (N_20348,N_17353,N_16196);
xor U20349 (N_20349,N_13636,N_14085);
and U20350 (N_20350,N_17202,N_15904);
or U20351 (N_20351,N_17918,N_13597);
nor U20352 (N_20352,N_14766,N_14370);
xnor U20353 (N_20353,N_14749,N_17929);
nor U20354 (N_20354,N_13984,N_12438);
xnor U20355 (N_20355,N_16867,N_16210);
nand U20356 (N_20356,N_17250,N_12294);
xnor U20357 (N_20357,N_14934,N_12432);
nand U20358 (N_20358,N_16991,N_16774);
nor U20359 (N_20359,N_16558,N_16090);
and U20360 (N_20360,N_15079,N_14796);
and U20361 (N_20361,N_12322,N_15402);
or U20362 (N_20362,N_12206,N_15603);
nand U20363 (N_20363,N_13159,N_14877);
xnor U20364 (N_20364,N_16192,N_17730);
nor U20365 (N_20365,N_14360,N_12375);
nand U20366 (N_20366,N_15113,N_15157);
nand U20367 (N_20367,N_16501,N_12352);
and U20368 (N_20368,N_13413,N_15363);
nand U20369 (N_20369,N_16106,N_16574);
xnor U20370 (N_20370,N_17849,N_17144);
and U20371 (N_20371,N_16054,N_17287);
xor U20372 (N_20372,N_15803,N_17247);
or U20373 (N_20373,N_14079,N_14831);
or U20374 (N_20374,N_13576,N_16216);
xnor U20375 (N_20375,N_15076,N_12185);
xnor U20376 (N_20376,N_16050,N_12728);
xnor U20377 (N_20377,N_16997,N_14632);
or U20378 (N_20378,N_17188,N_12210);
xnor U20379 (N_20379,N_16862,N_13069);
nor U20380 (N_20380,N_17867,N_12116);
nand U20381 (N_20381,N_12402,N_15374);
and U20382 (N_20382,N_17046,N_16267);
or U20383 (N_20383,N_16885,N_14584);
or U20384 (N_20384,N_12853,N_15529);
xor U20385 (N_20385,N_14622,N_17687);
nor U20386 (N_20386,N_14044,N_16691);
nor U20387 (N_20387,N_16913,N_17384);
nand U20388 (N_20388,N_17219,N_15163);
xor U20389 (N_20389,N_16966,N_17627);
nand U20390 (N_20390,N_17573,N_12075);
nand U20391 (N_20391,N_13216,N_15203);
or U20392 (N_20392,N_17158,N_14549);
xor U20393 (N_20393,N_12517,N_13621);
xor U20394 (N_20394,N_14232,N_12190);
or U20395 (N_20395,N_16597,N_12095);
xnor U20396 (N_20396,N_16188,N_13177);
xnor U20397 (N_20397,N_16072,N_13903);
xnor U20398 (N_20398,N_14996,N_15246);
or U20399 (N_20399,N_16854,N_13746);
xor U20400 (N_20400,N_14211,N_16019);
or U20401 (N_20401,N_13794,N_17107);
nand U20402 (N_20402,N_16289,N_15033);
nor U20403 (N_20403,N_17404,N_15284);
and U20404 (N_20404,N_13848,N_15786);
nand U20405 (N_20405,N_14626,N_16299);
nor U20406 (N_20406,N_14976,N_13121);
or U20407 (N_20407,N_17477,N_17061);
nor U20408 (N_20408,N_16127,N_17928);
nand U20409 (N_20409,N_13381,N_13590);
nor U20410 (N_20410,N_15952,N_15992);
or U20411 (N_20411,N_15537,N_17268);
xnor U20412 (N_20412,N_13383,N_12791);
and U20413 (N_20413,N_17417,N_17977);
and U20414 (N_20414,N_16803,N_17840);
xor U20415 (N_20415,N_13832,N_14702);
nand U20416 (N_20416,N_13201,N_12354);
nor U20417 (N_20417,N_17435,N_15210);
or U20418 (N_20418,N_16433,N_16483);
nand U20419 (N_20419,N_15090,N_16707);
nor U20420 (N_20420,N_14533,N_17007);
or U20421 (N_20421,N_13353,N_16660);
xor U20422 (N_20422,N_14709,N_15398);
and U20423 (N_20423,N_13009,N_13768);
or U20424 (N_20424,N_16801,N_17259);
xor U20425 (N_20425,N_13532,N_12641);
nand U20426 (N_20426,N_15558,N_17706);
nand U20427 (N_20427,N_15253,N_17304);
or U20428 (N_20428,N_14718,N_12972);
nor U20429 (N_20429,N_17303,N_16845);
or U20430 (N_20430,N_17335,N_14803);
xnor U20431 (N_20431,N_12937,N_15062);
xor U20432 (N_20432,N_17057,N_17970);
and U20433 (N_20433,N_12399,N_12313);
or U20434 (N_20434,N_15900,N_15236);
or U20435 (N_20435,N_12908,N_14231);
xnor U20436 (N_20436,N_12725,N_15376);
and U20437 (N_20437,N_13530,N_14429);
and U20438 (N_20438,N_13390,N_16348);
and U20439 (N_20439,N_16339,N_15422);
xnor U20440 (N_20440,N_16030,N_13735);
nand U20441 (N_20441,N_16278,N_15135);
and U20442 (N_20442,N_14381,N_14417);
or U20443 (N_20443,N_13907,N_17480);
and U20444 (N_20444,N_15240,N_14014);
xor U20445 (N_20445,N_15768,N_17427);
nor U20446 (N_20446,N_16665,N_17669);
or U20447 (N_20447,N_17900,N_14519);
nand U20448 (N_20448,N_13948,N_16445);
nor U20449 (N_20449,N_16249,N_12189);
xor U20450 (N_20450,N_12923,N_12576);
and U20451 (N_20451,N_16503,N_12766);
or U20452 (N_20452,N_12196,N_14525);
nor U20453 (N_20453,N_16438,N_15017);
and U20454 (N_20454,N_14793,N_16064);
or U20455 (N_20455,N_12558,N_15138);
and U20456 (N_20456,N_13494,N_17871);
nand U20457 (N_20457,N_13475,N_15371);
and U20458 (N_20458,N_15421,N_17363);
xnor U20459 (N_20459,N_14301,N_14541);
and U20460 (N_20460,N_16460,N_13501);
or U20461 (N_20461,N_15408,N_15629);
xnor U20462 (N_20462,N_14127,N_17756);
nand U20463 (N_20463,N_16323,N_12486);
and U20464 (N_20464,N_14878,N_16049);
xor U20465 (N_20465,N_12703,N_15028);
nor U20466 (N_20466,N_14249,N_15187);
nor U20467 (N_20467,N_16739,N_16136);
xnor U20468 (N_20468,N_15013,N_15483);
xnor U20469 (N_20469,N_15167,N_16051);
nand U20470 (N_20470,N_13314,N_12721);
xor U20471 (N_20471,N_12949,N_13560);
or U20472 (N_20472,N_14155,N_13286);
nor U20473 (N_20473,N_17327,N_12272);
nand U20474 (N_20474,N_16421,N_14049);
or U20475 (N_20475,N_14487,N_17643);
nor U20476 (N_20476,N_17461,N_14760);
or U20477 (N_20477,N_13466,N_12989);
nand U20478 (N_20478,N_15498,N_16843);
and U20479 (N_20479,N_16888,N_12407);
and U20480 (N_20480,N_13234,N_17318);
nor U20481 (N_20481,N_12027,N_13359);
nand U20482 (N_20482,N_17018,N_17753);
nor U20483 (N_20483,N_14156,N_17855);
nor U20484 (N_20484,N_13267,N_15600);
or U20485 (N_20485,N_17315,N_17056);
xnor U20486 (N_20486,N_12886,N_12663);
xnor U20487 (N_20487,N_17215,N_12138);
nand U20488 (N_20488,N_15504,N_14923);
xor U20489 (N_20489,N_17525,N_13287);
xnor U20490 (N_20490,N_17431,N_12173);
nand U20491 (N_20491,N_17205,N_14529);
nor U20492 (N_20492,N_17109,N_13373);
nand U20493 (N_20493,N_17120,N_17222);
nand U20494 (N_20494,N_15143,N_12948);
or U20495 (N_20495,N_17137,N_15583);
or U20496 (N_20496,N_14246,N_13533);
or U20497 (N_20497,N_17388,N_17080);
or U20498 (N_20498,N_15823,N_16383);
nand U20499 (N_20499,N_13424,N_15277);
nand U20500 (N_20500,N_12582,N_15799);
nor U20501 (N_20501,N_12458,N_15319);
and U20502 (N_20502,N_13514,N_14009);
or U20503 (N_20503,N_16172,N_17907);
xnor U20504 (N_20504,N_13634,N_15364);
or U20505 (N_20505,N_16119,N_17757);
nand U20506 (N_20506,N_16965,N_14181);
or U20507 (N_20507,N_14347,N_13247);
and U20508 (N_20508,N_13304,N_16215);
and U20509 (N_20509,N_15982,N_12479);
xnor U20510 (N_20510,N_16314,N_14225);
or U20511 (N_20511,N_17345,N_12406);
nor U20512 (N_20512,N_14792,N_12049);
or U20513 (N_20513,N_14204,N_16357);
and U20514 (N_20514,N_17496,N_14801);
nor U20515 (N_20515,N_12649,N_12038);
xor U20516 (N_20516,N_14435,N_16038);
or U20517 (N_20517,N_15635,N_16912);
or U20518 (N_20518,N_15976,N_15263);
or U20519 (N_20519,N_13770,N_12427);
nand U20520 (N_20520,N_12423,N_13743);
nand U20521 (N_20521,N_16533,N_17912);
or U20522 (N_20522,N_12472,N_12902);
and U20523 (N_20523,N_16477,N_15245);
xor U20524 (N_20524,N_14025,N_14006);
or U20525 (N_20525,N_15287,N_15675);
nor U20526 (N_20526,N_17965,N_12243);
nand U20527 (N_20527,N_16616,N_14896);
or U20528 (N_20528,N_13508,N_17768);
and U20529 (N_20529,N_15943,N_14515);
or U20530 (N_20530,N_12218,N_17668);
and U20531 (N_20531,N_13854,N_17357);
xnor U20532 (N_20532,N_16752,N_15719);
nand U20533 (N_20533,N_17123,N_16089);
nor U20534 (N_20534,N_17016,N_12647);
nor U20535 (N_20535,N_15978,N_16260);
nor U20536 (N_20536,N_12928,N_16152);
nand U20537 (N_20537,N_13392,N_16024);
nand U20538 (N_20538,N_12633,N_17449);
and U20539 (N_20539,N_13136,N_12256);
or U20540 (N_20540,N_17020,N_13884);
and U20541 (N_20541,N_13643,N_12879);
nand U20542 (N_20542,N_13571,N_13549);
xnor U20543 (N_20543,N_17714,N_15922);
xnor U20544 (N_20544,N_16895,N_15217);
xor U20545 (N_20545,N_13097,N_13812);
nand U20546 (N_20546,N_12962,N_16903);
or U20547 (N_20547,N_13071,N_12543);
nor U20548 (N_20548,N_16382,N_16715);
and U20549 (N_20549,N_13031,N_17497);
and U20550 (N_20550,N_15470,N_15727);
nor U20551 (N_20551,N_13120,N_16755);
xnor U20552 (N_20552,N_12341,N_16757);
xor U20553 (N_20553,N_12268,N_12952);
and U20554 (N_20554,N_14192,N_15903);
nor U20555 (N_20555,N_16919,N_16846);
nor U20556 (N_20556,N_15150,N_14646);
nor U20557 (N_20557,N_12005,N_15031);
xor U20558 (N_20558,N_12930,N_16873);
nor U20559 (N_20559,N_16124,N_12653);
and U20560 (N_20560,N_16815,N_14485);
nand U20561 (N_20561,N_16771,N_17605);
xnor U20562 (N_20562,N_14743,N_17386);
or U20563 (N_20563,N_12593,N_14074);
nor U20564 (N_20564,N_13647,N_14531);
or U20565 (N_20565,N_13328,N_12193);
or U20566 (N_20566,N_13629,N_17836);
nand U20567 (N_20567,N_15935,N_14922);
or U20568 (N_20568,N_17275,N_12483);
xnor U20569 (N_20569,N_17959,N_17214);
nor U20570 (N_20570,N_15595,N_17571);
nand U20571 (N_20571,N_15604,N_15802);
and U20572 (N_20572,N_15606,N_14017);
or U20573 (N_20573,N_14633,N_15067);
or U20574 (N_20574,N_12693,N_17762);
nor U20575 (N_20575,N_14066,N_17862);
nor U20576 (N_20576,N_14735,N_12504);
nor U20577 (N_20577,N_16419,N_16428);
and U20578 (N_20578,N_14363,N_15934);
and U20579 (N_20579,N_13778,N_17713);
nor U20580 (N_20580,N_14662,N_15035);
nor U20581 (N_20581,N_12052,N_13346);
xor U20582 (N_20582,N_13776,N_17647);
or U20583 (N_20583,N_12418,N_13010);
and U20584 (N_20584,N_12553,N_15456);
nor U20585 (N_20585,N_17631,N_13430);
nor U20586 (N_20586,N_12060,N_16107);
or U20587 (N_20587,N_13265,N_15008);
nand U20588 (N_20588,N_16915,N_12696);
xnor U20589 (N_20589,N_15848,N_16999);
or U20590 (N_20590,N_16901,N_12835);
xnor U20591 (N_20591,N_13385,N_13522);
nor U20592 (N_20592,N_15375,N_13793);
nand U20593 (N_20593,N_12153,N_15427);
and U20594 (N_20594,N_16699,N_17084);
and U20595 (N_20595,N_15907,N_16800);
and U20596 (N_20596,N_16909,N_15829);
xnor U20597 (N_20597,N_14806,N_15871);
and U20598 (N_20598,N_12692,N_15923);
or U20599 (N_20599,N_17933,N_14697);
and U20600 (N_20600,N_12875,N_14024);
nor U20601 (N_20601,N_17149,N_16376);
and U20602 (N_20602,N_16564,N_15597);
and U20603 (N_20603,N_14651,N_13048);
nand U20604 (N_20604,N_13696,N_17864);
nand U20605 (N_20605,N_15265,N_15262);
and U20606 (N_20606,N_17368,N_13958);
or U20607 (N_20607,N_15126,N_17847);
nor U20608 (N_20608,N_12217,N_15068);
xnor U20609 (N_20609,N_13734,N_16615);
xor U20610 (N_20610,N_16576,N_14122);
and U20611 (N_20611,N_14946,N_12980);
and U20612 (N_20612,N_13841,N_12395);
or U20613 (N_20613,N_14457,N_13021);
or U20614 (N_20614,N_13512,N_17237);
xnor U20615 (N_20615,N_14739,N_15941);
and U20616 (N_20616,N_14939,N_14468);
nand U20617 (N_20617,N_13204,N_12430);
xnor U20618 (N_20618,N_17421,N_17013);
xnor U20619 (N_20619,N_15750,N_14259);
and U20620 (N_20620,N_12141,N_14680);
nor U20621 (N_20621,N_12462,N_17284);
or U20622 (N_20622,N_14197,N_14769);
xnor U20623 (N_20623,N_13220,N_14717);
and U20624 (N_20624,N_16109,N_14004);
or U20625 (N_20625,N_17759,N_17450);
or U20626 (N_20626,N_17992,N_13405);
or U20627 (N_20627,N_13366,N_16590);
xor U20628 (N_20628,N_15381,N_14758);
and U20629 (N_20629,N_12323,N_14109);
and U20630 (N_20630,N_14895,N_15057);
xor U20631 (N_20631,N_12583,N_16507);
and U20632 (N_20632,N_13762,N_12059);
nor U20633 (N_20633,N_12716,N_13469);
nand U20634 (N_20634,N_14755,N_12530);
nor U20635 (N_20635,N_12401,N_13296);
or U20636 (N_20636,N_13526,N_15001);
nor U20637 (N_20637,N_16988,N_15705);
nand U20638 (N_20638,N_16612,N_15715);
nand U20639 (N_20639,N_14087,N_16359);
and U20640 (N_20640,N_12911,N_16296);
nor U20641 (N_20641,N_15112,N_16586);
and U20642 (N_20642,N_15863,N_16132);
nor U20643 (N_20643,N_15960,N_14617);
nor U20644 (N_20644,N_12107,N_16486);
and U20645 (N_20645,N_12849,N_12319);
and U20646 (N_20646,N_17723,N_13282);
nand U20647 (N_20647,N_16450,N_14693);
and U20648 (N_20648,N_12846,N_14162);
nor U20649 (N_20649,N_16471,N_16148);
or U20650 (N_20650,N_16227,N_14051);
and U20651 (N_20651,N_17342,N_12830);
nand U20652 (N_20652,N_15946,N_14003);
nand U20653 (N_20653,N_13249,N_13194);
nand U20654 (N_20654,N_13650,N_16184);
nand U20655 (N_20655,N_17508,N_12496);
nor U20656 (N_20656,N_12628,N_17380);
xor U20657 (N_20657,N_17735,N_17680);
and U20658 (N_20658,N_15264,N_13753);
and U20659 (N_20659,N_17913,N_13446);
nand U20660 (N_20660,N_13855,N_15266);
and U20661 (N_20661,N_15382,N_12400);
or U20662 (N_20662,N_14427,N_17512);
and U20663 (N_20663,N_17014,N_13601);
nor U20664 (N_20664,N_13342,N_16011);
or U20665 (N_20665,N_17045,N_14725);
or U20666 (N_20666,N_12842,N_15906);
or U20667 (N_20667,N_12142,N_12559);
nor U20668 (N_20668,N_16324,N_15288);
nand U20669 (N_20669,N_16204,N_16456);
nor U20670 (N_20670,N_14336,N_17087);
nor U20671 (N_20671,N_16097,N_14888);
and U20672 (N_20672,N_16946,N_17911);
xnor U20673 (N_20673,N_15958,N_15532);
nor U20674 (N_20674,N_12639,N_14058);
nor U20675 (N_20675,N_17030,N_14963);
and U20676 (N_20676,N_17167,N_15614);
nand U20677 (N_20677,N_14035,N_14909);
and U20678 (N_20678,N_13202,N_12009);
and U20679 (N_20679,N_16512,N_16411);
nor U20680 (N_20680,N_16544,N_14415);
xor U20681 (N_20681,N_17873,N_12287);
nor U20682 (N_20682,N_15458,N_16768);
xor U20683 (N_20683,N_15235,N_12198);
or U20684 (N_20684,N_16255,N_17077);
xnor U20685 (N_20685,N_17536,N_14497);
and U20686 (N_20686,N_13235,N_13882);
nor U20687 (N_20687,N_16861,N_17330);
or U20688 (N_20688,N_17956,N_14344);
xor U20689 (N_20689,N_17000,N_14940);
xor U20690 (N_20690,N_15818,N_12802);
nand U20691 (N_20691,N_15951,N_12990);
nand U20692 (N_20692,N_16488,N_17526);
nand U20693 (N_20693,N_16473,N_15229);
nand U20694 (N_20694,N_15550,N_16922);
nor U20695 (N_20695,N_12568,N_17468);
nor U20696 (N_20696,N_15372,N_14080);
nand U20697 (N_20697,N_17858,N_17032);
nand U20698 (N_20698,N_13391,N_12127);
xor U20699 (N_20699,N_15687,N_12501);
xor U20700 (N_20700,N_17876,N_17064);
nor U20701 (N_20701,N_12859,N_12161);
and U20702 (N_20702,N_13582,N_16151);
and U20703 (N_20703,N_17260,N_17406);
or U20704 (N_20704,N_15390,N_16408);
xnor U20705 (N_20705,N_12369,N_12082);
or U20706 (N_20706,N_15543,N_16588);
xor U20707 (N_20707,N_17423,N_13869);
nand U20708 (N_20708,N_13115,N_12167);
and U20709 (N_20709,N_16819,N_16711);
or U20710 (N_20710,N_15630,N_14902);
and U20711 (N_20711,N_16256,N_16761);
and U20712 (N_20712,N_12661,N_12771);
nor U20713 (N_20713,N_17740,N_17169);
nand U20714 (N_20714,N_12484,N_13007);
xor U20715 (N_20715,N_17424,N_16634);
or U20716 (N_20716,N_12834,N_14851);
or U20717 (N_20717,N_14919,N_12493);
or U20718 (N_20718,N_14654,N_14099);
or U20719 (N_20719,N_13680,N_13866);
nand U20720 (N_20720,N_14527,N_13938);
nor U20721 (N_20721,N_15345,N_12678);
and U20722 (N_20722,N_17899,N_15939);
nand U20723 (N_20723,N_17096,N_13453);
xor U20724 (N_20724,N_14434,N_16345);
nand U20725 (N_20725,N_14597,N_12861);
nor U20726 (N_20726,N_15239,N_12373);
xnor U20727 (N_20727,N_12340,N_17765);
nor U20728 (N_20728,N_13455,N_15984);
or U20729 (N_20729,N_14046,N_15665);
nand U20730 (N_20730,N_12591,N_14409);
and U20731 (N_20731,N_14833,N_15516);
and U20732 (N_20732,N_13850,N_15330);
nand U20733 (N_20733,N_13563,N_15409);
nand U20734 (N_20734,N_14748,N_17866);
nor U20735 (N_20735,N_16108,N_16195);
nand U20736 (N_20736,N_12529,N_13137);
or U20737 (N_20737,N_14013,N_14684);
nor U20738 (N_20738,N_15776,N_12519);
xor U20739 (N_20739,N_15921,N_15156);
and U20740 (N_20740,N_17737,N_14442);
xor U20741 (N_20741,N_15887,N_15129);
xnor U20742 (N_20742,N_12840,N_14018);
nand U20743 (N_20743,N_12537,N_12440);
and U20744 (N_20744,N_12745,N_16202);
nand U20745 (N_20745,N_17437,N_14707);
and U20746 (N_20746,N_17767,N_15197);
xor U20747 (N_20747,N_13702,N_17469);
or U20748 (N_20748,N_16834,N_15990);
or U20749 (N_20749,N_12259,N_12204);
nor U20750 (N_20750,N_17947,N_13779);
or U20751 (N_20751,N_15180,N_14260);
nor U20752 (N_20752,N_16073,N_12216);
and U20753 (N_20753,N_13836,N_16468);
and U20754 (N_20754,N_12258,N_12492);
nand U20755 (N_20755,N_17200,N_13860);
xor U20756 (N_20756,N_14444,N_17136);
xor U20757 (N_20757,N_17891,N_14557);
nor U20758 (N_20758,N_16449,N_15531);
nand U20759 (N_20759,N_15983,N_14586);
and U20760 (N_20760,N_13586,N_14820);
and U20761 (N_20761,N_12893,N_14986);
or U20762 (N_20762,N_16015,N_12627);
nor U20763 (N_20763,N_12446,N_13500);
nor U20764 (N_20764,N_14832,N_14991);
and U20765 (N_20765,N_15683,N_14371);
and U20766 (N_20766,N_12417,N_16789);
nand U20767 (N_20767,N_12442,N_14737);
nor U20768 (N_20768,N_16794,N_15942);
nand U20769 (N_20769,N_17934,N_12813);
xnor U20770 (N_20770,N_12832,N_16436);
or U20771 (N_20771,N_16694,N_13450);
xnor U20772 (N_20772,N_13933,N_12588);
nor U20773 (N_20773,N_15329,N_13706);
or U20774 (N_20774,N_16171,N_13341);
and U20775 (N_20775,N_16517,N_15999);
or U20776 (N_20776,N_14610,N_12594);
nor U20777 (N_20777,N_12488,N_12429);
or U20778 (N_20778,N_13966,N_16730);
or U20779 (N_20779,N_16554,N_16508);
nor U20780 (N_20780,N_16063,N_14845);
or U20781 (N_20781,N_17501,N_15541);
nor U20782 (N_20782,N_16163,N_13720);
or U20783 (N_20783,N_17853,N_15191);
or U20784 (N_20784,N_15136,N_16347);
or U20785 (N_20785,N_17697,N_15152);
nand U20786 (N_20786,N_16316,N_12109);
xor U20787 (N_20787,N_12386,N_14446);
nand U20788 (N_20788,N_12133,N_14837);
xnor U20789 (N_20789,N_17986,N_16208);
or U20790 (N_20790,N_15948,N_12964);
and U20791 (N_20791,N_15582,N_13440);
or U20792 (N_20792,N_13864,N_15255);
or U20793 (N_20793,N_13001,N_12804);
and U20794 (N_20794,N_12883,N_13008);
nand U20795 (N_20795,N_15879,N_13708);
or U20796 (N_20796,N_17814,N_15784);
or U20797 (N_20797,N_17837,N_12934);
or U20798 (N_20798,N_12237,N_15852);
and U20799 (N_20799,N_12921,N_16523);
or U20800 (N_20800,N_14545,N_12230);
or U20801 (N_20801,N_13992,N_13480);
nor U20802 (N_20802,N_15109,N_17352);
xnor U20803 (N_20803,N_12293,N_17883);
nand U20804 (N_20804,N_16790,N_17238);
or U20805 (N_20805,N_13129,N_17119);
and U20806 (N_20806,N_15276,N_13233);
nand U20807 (N_20807,N_15158,N_13093);
and U20808 (N_20808,N_16841,N_16096);
xnor U20809 (N_20809,N_12130,N_17531);
nand U20810 (N_20810,N_14138,N_14673);
and U20811 (N_20811,N_12461,N_16373);
nand U20812 (N_20812,N_14348,N_16937);
nor U20813 (N_20813,N_12068,N_14283);
nor U20814 (N_20814,N_16154,N_17519);
xor U20815 (N_20815,N_15778,N_17939);
nor U20816 (N_20816,N_15994,N_17028);
nand U20817 (N_20817,N_14352,N_12154);
and U20818 (N_20818,N_14176,N_15929);
or U20819 (N_20819,N_14228,N_14757);
nand U20820 (N_20820,N_16078,N_13967);
nand U20821 (N_20821,N_16746,N_17880);
nand U20822 (N_20822,N_17521,N_13109);
nor U20823 (N_20823,N_13679,N_15042);
and U20824 (N_20824,N_16175,N_13222);
or U20825 (N_20825,N_17892,N_13189);
xor U20826 (N_20826,N_13819,N_12844);
and U20827 (N_20827,N_13542,N_14063);
nor U20828 (N_20828,N_13641,N_14771);
nand U20829 (N_20829,N_13594,N_15796);
or U20830 (N_20830,N_14328,N_12723);
nand U20831 (N_20831,N_13320,N_14734);
nor U20832 (N_20832,N_15139,N_14505);
xor U20833 (N_20833,N_13824,N_15328);
and U20834 (N_20834,N_14669,N_15397);
xor U20835 (N_20835,N_16814,N_17821);
and U20836 (N_20836,N_15703,N_17399);
nor U20837 (N_20837,N_16086,N_14367);
xor U20838 (N_20838,N_13376,N_14362);
and U20839 (N_20839,N_12017,N_17190);
xnor U20840 (N_20840,N_12137,N_13844);
nand U20841 (N_20841,N_16176,N_15314);
or U20842 (N_20842,N_15080,N_15435);
nand U20843 (N_20843,N_13828,N_15628);
nor U20844 (N_20844,N_12436,N_16604);
or U20845 (N_20845,N_17161,N_17603);
nor U20846 (N_20846,N_17702,N_13820);
or U20847 (N_20847,N_15160,N_15071);
nand U20848 (N_20848,N_12836,N_17681);
or U20849 (N_20849,N_13057,N_14871);
or U20850 (N_20850,N_17216,N_15428);
xor U20851 (N_20851,N_13098,N_13518);
xor U20852 (N_20852,N_16082,N_12744);
or U20853 (N_20853,N_15810,N_15979);
and U20854 (N_20854,N_16653,N_14075);
xnor U20855 (N_20855,N_12767,N_16499);
nand U20856 (N_20856,N_17440,N_12094);
and U20857 (N_20857,N_15672,N_17720);
and U20858 (N_20858,N_12680,N_15298);
and U20859 (N_20859,N_13715,N_13095);
nand U20860 (N_20860,N_17063,N_17940);
nand U20861 (N_20861,N_17942,N_14048);
nand U20862 (N_20862,N_16391,N_12066);
or U20863 (N_20863,N_14407,N_16872);
or U20864 (N_20864,N_16637,N_16282);
nand U20865 (N_20865,N_13171,N_16810);
and U20866 (N_20866,N_16817,N_16668);
nand U20867 (N_20867,N_12473,N_14255);
nor U20868 (N_20868,N_14432,N_12555);
nand U20869 (N_20869,N_15475,N_16678);
xnor U20870 (N_20870,N_12812,N_12637);
nor U20871 (N_20871,N_14872,N_17679);
and U20872 (N_20872,N_14220,N_13340);
nand U20873 (N_20873,N_17157,N_13674);
xnor U20874 (N_20874,N_13573,N_14296);
and U20875 (N_20875,N_15987,N_17792);
or U20876 (N_20876,N_13289,N_13623);
or U20877 (N_20877,N_15170,N_12654);
nand U20878 (N_20878,N_17745,N_13363);
or U20879 (N_20879,N_15546,N_17400);
nand U20880 (N_20880,N_16875,N_15751);
nand U20881 (N_20881,N_12195,N_17882);
nor U20882 (N_20882,N_14911,N_16131);
nor U20883 (N_20883,N_17248,N_16823);
or U20884 (N_20884,N_15494,N_13200);
nand U20885 (N_20885,N_14070,N_12670);
nand U20886 (N_20886,N_15572,N_12700);
nor U20887 (N_20887,N_17741,N_16571);
nand U20888 (N_20888,N_15792,N_12955);
nor U20889 (N_20889,N_12951,N_16277);
xor U20890 (N_20890,N_13101,N_16307);
xnor U20891 (N_20891,N_16352,N_15142);
and U20892 (N_20892,N_16230,N_17272);
xor U20893 (N_20893,N_12003,N_13108);
and U20894 (N_20894,N_16243,N_16560);
nand U20895 (N_20895,N_14477,N_15856);
xor U20896 (N_20896,N_12251,N_14784);
and U20897 (N_20897,N_15706,N_14050);
and U20898 (N_20898,N_13950,N_13038);
nand U20899 (N_20899,N_16575,N_14104);
nor U20900 (N_20900,N_15302,N_14433);
or U20901 (N_20901,N_12622,N_14897);
or U20902 (N_20902,N_13035,N_17967);
or U20903 (N_20903,N_14822,N_14270);
xor U20904 (N_20904,N_12741,N_14257);
and U20905 (N_20905,N_13703,N_15413);
nand U20906 (N_20906,N_17204,N_13485);
nand U20907 (N_20907,N_12885,N_15202);
nor U20908 (N_20908,N_15584,N_16585);
xnor U20909 (N_20909,N_12491,N_17700);
nor U20910 (N_20910,N_13477,N_15213);
and U20911 (N_20911,N_13052,N_16504);
and U20912 (N_20912,N_17560,N_15122);
nor U20913 (N_20913,N_15338,N_14738);
nor U20914 (N_20914,N_14712,N_16191);
or U20915 (N_20915,N_15238,N_16811);
xor U20916 (N_20916,N_15101,N_12965);
xnor U20917 (N_20917,N_15807,N_12064);
or U20918 (N_20918,N_12604,N_15269);
or U20919 (N_20919,N_13665,N_17856);
xnor U20920 (N_20920,N_12612,N_12124);
xor U20921 (N_20921,N_14469,N_15453);
nand U20922 (N_20922,N_12187,N_17763);
and U20923 (N_20923,N_16565,N_17325);
nand U20924 (N_20924,N_17542,N_15123);
and U20925 (N_20925,N_15886,N_15007);
nand U20926 (N_20926,N_14419,N_13695);
xnor U20927 (N_20927,N_15816,N_12269);
nor U20928 (N_20928,N_16772,N_17660);
or U20929 (N_20929,N_15955,N_15611);
nand U20930 (N_20930,N_17379,N_13534);
nand U20931 (N_20931,N_12081,N_15081);
nor U20932 (N_20932,N_12808,N_16040);
nand U20933 (N_20933,N_17686,N_12065);
and U20934 (N_20934,N_17280,N_16855);
and U20935 (N_20935,N_16081,N_14560);
and U20936 (N_20936,N_15506,N_13839);
nor U20937 (N_20937,N_15430,N_16802);
nor U20938 (N_20938,N_15777,N_15677);
or U20939 (N_20939,N_14256,N_13554);
nand U20940 (N_20940,N_12470,N_17138);
and U20941 (N_20941,N_13130,N_13944);
nand U20942 (N_20942,N_13911,N_13976);
nor U20943 (N_20943,N_17514,N_13712);
or U20944 (N_20944,N_12688,N_13797);
nor U20945 (N_20945,N_15151,N_16280);
xnor U20946 (N_20946,N_14958,N_15325);
and U20947 (N_20947,N_14591,N_16235);
or U20948 (N_20948,N_17383,N_14502);
nand U20949 (N_20949,N_14521,N_12575);
xor U20950 (N_20950,N_13640,N_16418);
and U20951 (N_20951,N_13221,N_14292);
or U20952 (N_20952,N_12197,N_16613);
nor U20953 (N_20953,N_17050,N_17274);
nand U20954 (N_20954,N_13364,N_15744);
and U20955 (N_20955,N_13873,N_17772);
xor U20956 (N_20956,N_15918,N_15128);
or U20957 (N_20957,N_15055,N_15944);
and U20958 (N_20958,N_16962,N_15137);
nand U20959 (N_20959,N_17738,N_14187);
xnor U20960 (N_20960,N_16970,N_15087);
nand U20961 (N_20961,N_15945,N_13939);
or U20962 (N_20962,N_14989,N_13311);
xnor U20963 (N_20963,N_16187,N_13173);
nand U20964 (N_20964,N_16261,N_16706);
or U20965 (N_20965,N_14975,N_14258);
and U20966 (N_20966,N_16016,N_14115);
nor U20967 (N_20967,N_13513,N_17463);
xor U20968 (N_20968,N_16526,N_16130);
nor U20969 (N_20969,N_15782,N_13210);
and U20970 (N_20970,N_16448,N_14640);
or U20971 (N_20971,N_13427,N_17183);
nand U20972 (N_20972,N_14108,N_16809);
or U20973 (N_20973,N_17588,N_17418);
and U20974 (N_20974,N_16190,N_14835);
and U20975 (N_20975,N_13192,N_17128);
or U20976 (N_20976,N_17147,N_15367);
or U20977 (N_20977,N_13899,N_15542);
nor U20978 (N_20978,N_13160,N_12136);
nor U20979 (N_20979,N_12954,N_14186);
nand U20980 (N_20980,N_16022,N_15324);
and U20981 (N_20981,N_14416,N_15685);
xor U20982 (N_20982,N_12740,N_17278);
nand U20983 (N_20983,N_17978,N_12777);
nand U20984 (N_20984,N_15116,N_17261);
and U20985 (N_20985,N_16302,N_15837);
and U20986 (N_20986,N_15195,N_12669);
nor U20987 (N_20987,N_17622,N_17830);
or U20988 (N_20988,N_13338,N_14539);
xor U20989 (N_20989,N_12213,N_13648);
xor U20990 (N_20990,N_12651,N_14394);
or U20991 (N_20991,N_14814,N_16551);
and U20992 (N_20992,N_15811,N_15445);
nor U20993 (N_20993,N_12887,N_14933);
nor U20994 (N_20994,N_14172,N_12106);
xnor U20995 (N_20995,N_16442,N_15696);
nor U20996 (N_20996,N_17620,N_14687);
xnor U20997 (N_20997,N_13454,N_17586);
or U20998 (N_20998,N_13845,N_16298);
nand U20999 (N_20999,N_12274,N_12695);
xnor U21000 (N_21000,N_17080,N_13959);
and U21001 (N_21001,N_13546,N_17027);
or U21002 (N_21002,N_13641,N_14790);
and U21003 (N_21003,N_12760,N_14933);
and U21004 (N_21004,N_16570,N_13359);
nor U21005 (N_21005,N_15089,N_13723);
or U21006 (N_21006,N_17506,N_14425);
nand U21007 (N_21007,N_13105,N_14453);
or U21008 (N_21008,N_15784,N_13292);
nor U21009 (N_21009,N_17235,N_16721);
xor U21010 (N_21010,N_16017,N_16173);
xnor U21011 (N_21011,N_14200,N_14962);
and U21012 (N_21012,N_16599,N_13077);
nand U21013 (N_21013,N_13149,N_13224);
nand U21014 (N_21014,N_17609,N_16989);
nor U21015 (N_21015,N_16680,N_15549);
nor U21016 (N_21016,N_12419,N_15487);
or U21017 (N_21017,N_14381,N_13586);
nor U21018 (N_21018,N_13845,N_15353);
xnor U21019 (N_21019,N_14197,N_13229);
nand U21020 (N_21020,N_15848,N_16608);
and U21021 (N_21021,N_16669,N_17597);
and U21022 (N_21022,N_15878,N_17555);
nand U21023 (N_21023,N_17663,N_17425);
xor U21024 (N_21024,N_16679,N_13354);
nor U21025 (N_21025,N_14943,N_15111);
and U21026 (N_21026,N_13403,N_13299);
nor U21027 (N_21027,N_16204,N_14800);
xor U21028 (N_21028,N_17305,N_12528);
nor U21029 (N_21029,N_14879,N_14695);
or U21030 (N_21030,N_13657,N_14790);
xnor U21031 (N_21031,N_13612,N_14309);
nand U21032 (N_21032,N_17478,N_14186);
or U21033 (N_21033,N_16078,N_14190);
xnor U21034 (N_21034,N_12449,N_16426);
or U21035 (N_21035,N_14014,N_12190);
nor U21036 (N_21036,N_17614,N_15628);
nor U21037 (N_21037,N_13758,N_17433);
xor U21038 (N_21038,N_13952,N_15192);
and U21039 (N_21039,N_17326,N_12102);
nand U21040 (N_21040,N_17542,N_14813);
and U21041 (N_21041,N_16006,N_14266);
nor U21042 (N_21042,N_17376,N_17902);
nand U21043 (N_21043,N_14117,N_13786);
and U21044 (N_21044,N_15285,N_13437);
and U21045 (N_21045,N_15024,N_14047);
and U21046 (N_21046,N_15597,N_16617);
and U21047 (N_21047,N_14322,N_13319);
nor U21048 (N_21048,N_16819,N_14040);
nor U21049 (N_21049,N_13415,N_14385);
and U21050 (N_21050,N_15940,N_15540);
or U21051 (N_21051,N_13092,N_17746);
or U21052 (N_21052,N_12239,N_14795);
and U21053 (N_21053,N_16938,N_14387);
xnor U21054 (N_21054,N_14014,N_15326);
and U21055 (N_21055,N_12801,N_14561);
nor U21056 (N_21056,N_16847,N_13072);
nand U21057 (N_21057,N_13196,N_13732);
or U21058 (N_21058,N_12588,N_12639);
nand U21059 (N_21059,N_14438,N_14100);
and U21060 (N_21060,N_12216,N_12979);
xor U21061 (N_21061,N_16005,N_14730);
and U21062 (N_21062,N_15132,N_12407);
or U21063 (N_21063,N_15017,N_17320);
xor U21064 (N_21064,N_14761,N_13478);
nor U21065 (N_21065,N_14107,N_12884);
nor U21066 (N_21066,N_16134,N_14882);
nand U21067 (N_21067,N_16303,N_17268);
and U21068 (N_21068,N_17953,N_12591);
nand U21069 (N_21069,N_12544,N_12001);
nor U21070 (N_21070,N_17161,N_15722);
nand U21071 (N_21071,N_13774,N_13956);
or U21072 (N_21072,N_12124,N_15572);
nor U21073 (N_21073,N_14634,N_14748);
xor U21074 (N_21074,N_15656,N_12180);
or U21075 (N_21075,N_13036,N_14123);
xnor U21076 (N_21076,N_13370,N_13969);
or U21077 (N_21077,N_16626,N_12093);
or U21078 (N_21078,N_14720,N_14396);
nand U21079 (N_21079,N_16841,N_16778);
and U21080 (N_21080,N_14361,N_16342);
xnor U21081 (N_21081,N_17060,N_12354);
xnor U21082 (N_21082,N_15643,N_15936);
nor U21083 (N_21083,N_16432,N_15055);
or U21084 (N_21084,N_13177,N_16334);
nand U21085 (N_21085,N_15239,N_15085);
or U21086 (N_21086,N_17426,N_14666);
nand U21087 (N_21087,N_17495,N_12108);
or U21088 (N_21088,N_14737,N_16987);
nand U21089 (N_21089,N_14575,N_15820);
xor U21090 (N_21090,N_14889,N_14200);
xnor U21091 (N_21091,N_17262,N_13947);
and U21092 (N_21092,N_12798,N_16387);
xnor U21093 (N_21093,N_14884,N_13941);
and U21094 (N_21094,N_17103,N_12774);
and U21095 (N_21095,N_15363,N_15858);
nand U21096 (N_21096,N_17928,N_15852);
nand U21097 (N_21097,N_15845,N_14433);
and U21098 (N_21098,N_17852,N_14624);
or U21099 (N_21099,N_15862,N_17653);
xnor U21100 (N_21100,N_12934,N_12385);
xnor U21101 (N_21101,N_14848,N_15396);
nand U21102 (N_21102,N_16146,N_17950);
nand U21103 (N_21103,N_13032,N_13247);
nand U21104 (N_21104,N_15199,N_12880);
nand U21105 (N_21105,N_17230,N_13116);
nand U21106 (N_21106,N_17077,N_16412);
and U21107 (N_21107,N_12036,N_16297);
or U21108 (N_21108,N_17590,N_12772);
nor U21109 (N_21109,N_14480,N_12781);
nand U21110 (N_21110,N_16309,N_16292);
xor U21111 (N_21111,N_12776,N_16000);
or U21112 (N_21112,N_14508,N_17166);
or U21113 (N_21113,N_16593,N_12455);
and U21114 (N_21114,N_13556,N_16738);
and U21115 (N_21115,N_12795,N_14850);
nand U21116 (N_21116,N_15361,N_17397);
xnor U21117 (N_21117,N_13384,N_17214);
or U21118 (N_21118,N_13715,N_12686);
nor U21119 (N_21119,N_16102,N_16384);
or U21120 (N_21120,N_15620,N_12941);
xor U21121 (N_21121,N_14781,N_12958);
and U21122 (N_21122,N_15436,N_15955);
nor U21123 (N_21123,N_13217,N_12727);
xnor U21124 (N_21124,N_15926,N_14792);
xnor U21125 (N_21125,N_12360,N_13133);
xor U21126 (N_21126,N_14816,N_16011);
nor U21127 (N_21127,N_14619,N_16732);
xnor U21128 (N_21128,N_17145,N_12320);
and U21129 (N_21129,N_17684,N_17380);
xor U21130 (N_21130,N_12457,N_15293);
xor U21131 (N_21131,N_14126,N_12331);
and U21132 (N_21132,N_13010,N_12072);
nand U21133 (N_21133,N_13474,N_17462);
nor U21134 (N_21134,N_14235,N_13618);
nor U21135 (N_21135,N_16320,N_17747);
nor U21136 (N_21136,N_14912,N_13222);
xnor U21137 (N_21137,N_16733,N_12738);
and U21138 (N_21138,N_12471,N_16168);
nor U21139 (N_21139,N_12098,N_16009);
or U21140 (N_21140,N_12444,N_12071);
nand U21141 (N_21141,N_16966,N_16540);
or U21142 (N_21142,N_17562,N_15009);
nor U21143 (N_21143,N_16360,N_14279);
or U21144 (N_21144,N_17457,N_12008);
or U21145 (N_21145,N_13401,N_17762);
nor U21146 (N_21146,N_17075,N_14631);
nor U21147 (N_21147,N_16494,N_16183);
nor U21148 (N_21148,N_16537,N_15745);
xor U21149 (N_21149,N_15245,N_13254);
and U21150 (N_21150,N_17568,N_15292);
xor U21151 (N_21151,N_17606,N_12740);
xor U21152 (N_21152,N_14630,N_12800);
and U21153 (N_21153,N_15904,N_17413);
nand U21154 (N_21154,N_16420,N_16384);
and U21155 (N_21155,N_17931,N_13367);
or U21156 (N_21156,N_12258,N_16042);
xor U21157 (N_21157,N_13385,N_14843);
nor U21158 (N_21158,N_16706,N_16211);
xor U21159 (N_21159,N_14015,N_17337);
xnor U21160 (N_21160,N_14035,N_15990);
and U21161 (N_21161,N_12858,N_14684);
and U21162 (N_21162,N_17997,N_14151);
or U21163 (N_21163,N_12515,N_15208);
nand U21164 (N_21164,N_12748,N_13910);
nor U21165 (N_21165,N_12490,N_14880);
and U21166 (N_21166,N_15371,N_15294);
nand U21167 (N_21167,N_17368,N_17301);
nor U21168 (N_21168,N_12021,N_13243);
or U21169 (N_21169,N_16975,N_15830);
or U21170 (N_21170,N_17567,N_15551);
or U21171 (N_21171,N_12298,N_17145);
nor U21172 (N_21172,N_14444,N_15334);
and U21173 (N_21173,N_13819,N_16981);
nand U21174 (N_21174,N_13333,N_13883);
nor U21175 (N_21175,N_14408,N_14380);
or U21176 (N_21176,N_16444,N_15755);
or U21177 (N_21177,N_13623,N_15012);
nand U21178 (N_21178,N_14153,N_13611);
nor U21179 (N_21179,N_12596,N_13727);
nand U21180 (N_21180,N_12519,N_14206);
xor U21181 (N_21181,N_15199,N_17549);
or U21182 (N_21182,N_14412,N_15635);
and U21183 (N_21183,N_13569,N_13507);
nor U21184 (N_21184,N_17623,N_13425);
xnor U21185 (N_21185,N_14640,N_13650);
nor U21186 (N_21186,N_13607,N_12323);
nor U21187 (N_21187,N_13392,N_14633);
xnor U21188 (N_21188,N_12361,N_14843);
nand U21189 (N_21189,N_15669,N_15560);
or U21190 (N_21190,N_15723,N_17591);
nor U21191 (N_21191,N_13378,N_12379);
nand U21192 (N_21192,N_16682,N_16066);
nand U21193 (N_21193,N_14249,N_16159);
or U21194 (N_21194,N_15144,N_17153);
xor U21195 (N_21195,N_17829,N_16951);
xor U21196 (N_21196,N_12286,N_13504);
nor U21197 (N_21197,N_16612,N_13927);
or U21198 (N_21198,N_14057,N_14666);
or U21199 (N_21199,N_16003,N_16069);
xnor U21200 (N_21200,N_13317,N_16970);
and U21201 (N_21201,N_17850,N_13621);
nor U21202 (N_21202,N_12462,N_12276);
xor U21203 (N_21203,N_15424,N_17656);
xor U21204 (N_21204,N_12737,N_13377);
and U21205 (N_21205,N_17227,N_13822);
and U21206 (N_21206,N_15373,N_16769);
nor U21207 (N_21207,N_15887,N_13132);
and U21208 (N_21208,N_17280,N_16239);
and U21209 (N_21209,N_16487,N_17661);
xor U21210 (N_21210,N_13968,N_16951);
and U21211 (N_21211,N_13663,N_16577);
nor U21212 (N_21212,N_13824,N_16255);
and U21213 (N_21213,N_14676,N_16031);
or U21214 (N_21214,N_14952,N_17327);
xor U21215 (N_21215,N_17339,N_14616);
nand U21216 (N_21216,N_16286,N_16870);
xnor U21217 (N_21217,N_14027,N_16029);
or U21218 (N_21218,N_16522,N_12104);
xor U21219 (N_21219,N_13001,N_16745);
nand U21220 (N_21220,N_13299,N_16733);
nand U21221 (N_21221,N_15460,N_17305);
nand U21222 (N_21222,N_16553,N_15748);
and U21223 (N_21223,N_15545,N_12441);
xnor U21224 (N_21224,N_15949,N_16806);
nand U21225 (N_21225,N_15829,N_16614);
nand U21226 (N_21226,N_15539,N_14928);
xor U21227 (N_21227,N_17407,N_13637);
xnor U21228 (N_21228,N_17463,N_12129);
nand U21229 (N_21229,N_15636,N_15962);
and U21230 (N_21230,N_17279,N_13888);
xor U21231 (N_21231,N_13209,N_13506);
nor U21232 (N_21232,N_17182,N_12203);
nand U21233 (N_21233,N_15753,N_15166);
and U21234 (N_21234,N_13311,N_14935);
or U21235 (N_21235,N_14430,N_13229);
nand U21236 (N_21236,N_17146,N_14590);
xor U21237 (N_21237,N_16933,N_15641);
and U21238 (N_21238,N_17183,N_12379);
nand U21239 (N_21239,N_13191,N_13031);
nor U21240 (N_21240,N_17673,N_12463);
nand U21241 (N_21241,N_17051,N_17122);
xor U21242 (N_21242,N_17139,N_16308);
xor U21243 (N_21243,N_13086,N_13931);
nor U21244 (N_21244,N_15364,N_15691);
xor U21245 (N_21245,N_14097,N_17599);
nor U21246 (N_21246,N_17780,N_15409);
nand U21247 (N_21247,N_17026,N_12025);
or U21248 (N_21248,N_15838,N_12112);
or U21249 (N_21249,N_13563,N_17831);
or U21250 (N_21250,N_13614,N_15441);
and U21251 (N_21251,N_16621,N_17953);
and U21252 (N_21252,N_17673,N_15810);
nand U21253 (N_21253,N_14541,N_15949);
and U21254 (N_21254,N_13388,N_17545);
and U21255 (N_21255,N_13019,N_12411);
or U21256 (N_21256,N_17183,N_14112);
nor U21257 (N_21257,N_14529,N_13669);
nand U21258 (N_21258,N_14601,N_16490);
xnor U21259 (N_21259,N_13678,N_14591);
xnor U21260 (N_21260,N_15296,N_17306);
or U21261 (N_21261,N_14873,N_14731);
nor U21262 (N_21262,N_12684,N_13175);
and U21263 (N_21263,N_15479,N_15306);
and U21264 (N_21264,N_17518,N_12084);
nand U21265 (N_21265,N_17514,N_15896);
or U21266 (N_21266,N_13152,N_17476);
xnor U21267 (N_21267,N_17532,N_14322);
and U21268 (N_21268,N_15325,N_15481);
nand U21269 (N_21269,N_17055,N_12981);
and U21270 (N_21270,N_15907,N_12412);
nand U21271 (N_21271,N_13111,N_13509);
or U21272 (N_21272,N_14986,N_17356);
xor U21273 (N_21273,N_17700,N_16231);
nand U21274 (N_21274,N_14838,N_15809);
and U21275 (N_21275,N_15135,N_16057);
xnor U21276 (N_21276,N_13755,N_13199);
nand U21277 (N_21277,N_17145,N_14317);
nor U21278 (N_21278,N_13344,N_12589);
and U21279 (N_21279,N_17874,N_15439);
nor U21280 (N_21280,N_12936,N_14700);
or U21281 (N_21281,N_12837,N_14689);
and U21282 (N_21282,N_17069,N_12419);
nor U21283 (N_21283,N_12799,N_16940);
or U21284 (N_21284,N_13260,N_13372);
and U21285 (N_21285,N_17690,N_13669);
nand U21286 (N_21286,N_14594,N_14583);
nor U21287 (N_21287,N_17873,N_12942);
and U21288 (N_21288,N_13087,N_12176);
or U21289 (N_21289,N_12552,N_13334);
nor U21290 (N_21290,N_13903,N_15903);
or U21291 (N_21291,N_13552,N_16573);
nand U21292 (N_21292,N_12939,N_13242);
and U21293 (N_21293,N_17549,N_15606);
nor U21294 (N_21294,N_15888,N_13214);
nor U21295 (N_21295,N_17840,N_17914);
or U21296 (N_21296,N_13536,N_16187);
xor U21297 (N_21297,N_17340,N_16975);
nand U21298 (N_21298,N_16548,N_14702);
nand U21299 (N_21299,N_12658,N_17170);
nor U21300 (N_21300,N_14171,N_12354);
or U21301 (N_21301,N_16819,N_17302);
xnor U21302 (N_21302,N_13181,N_14629);
nor U21303 (N_21303,N_17931,N_12827);
nor U21304 (N_21304,N_13069,N_17200);
and U21305 (N_21305,N_15565,N_15951);
or U21306 (N_21306,N_17449,N_16876);
xor U21307 (N_21307,N_12356,N_15604);
nand U21308 (N_21308,N_13292,N_15433);
or U21309 (N_21309,N_16872,N_14059);
and U21310 (N_21310,N_15630,N_16134);
nor U21311 (N_21311,N_16733,N_16611);
nor U21312 (N_21312,N_16375,N_17901);
or U21313 (N_21313,N_15765,N_13032);
and U21314 (N_21314,N_13715,N_16084);
xor U21315 (N_21315,N_17436,N_16605);
or U21316 (N_21316,N_16019,N_13611);
nor U21317 (N_21317,N_14644,N_13681);
nand U21318 (N_21318,N_14181,N_17442);
xnor U21319 (N_21319,N_13928,N_15399);
xnor U21320 (N_21320,N_16023,N_15173);
xnor U21321 (N_21321,N_12349,N_13985);
nor U21322 (N_21322,N_12043,N_12545);
nand U21323 (N_21323,N_15995,N_17343);
and U21324 (N_21324,N_16604,N_14137);
nor U21325 (N_21325,N_14800,N_14962);
nor U21326 (N_21326,N_13655,N_15891);
xnor U21327 (N_21327,N_13325,N_17108);
nand U21328 (N_21328,N_17367,N_15529);
and U21329 (N_21329,N_15218,N_16965);
nand U21330 (N_21330,N_17355,N_15030);
nand U21331 (N_21331,N_14229,N_15256);
and U21332 (N_21332,N_14703,N_17861);
and U21333 (N_21333,N_14970,N_16717);
or U21334 (N_21334,N_13063,N_16527);
nand U21335 (N_21335,N_12190,N_16347);
nor U21336 (N_21336,N_12537,N_13867);
nand U21337 (N_21337,N_15523,N_16875);
xor U21338 (N_21338,N_13702,N_13514);
or U21339 (N_21339,N_15059,N_16645);
nand U21340 (N_21340,N_13498,N_17246);
xnor U21341 (N_21341,N_14932,N_15642);
xor U21342 (N_21342,N_13468,N_14340);
xor U21343 (N_21343,N_13933,N_14017);
or U21344 (N_21344,N_15889,N_17929);
xnor U21345 (N_21345,N_12940,N_13012);
nand U21346 (N_21346,N_13136,N_17276);
nor U21347 (N_21347,N_17006,N_15176);
nand U21348 (N_21348,N_16261,N_17035);
or U21349 (N_21349,N_16719,N_17717);
xnor U21350 (N_21350,N_15772,N_17019);
or U21351 (N_21351,N_14748,N_12434);
xnor U21352 (N_21352,N_14484,N_16341);
and U21353 (N_21353,N_15967,N_14039);
nand U21354 (N_21354,N_15157,N_12213);
or U21355 (N_21355,N_16480,N_16817);
nand U21356 (N_21356,N_12140,N_12838);
xor U21357 (N_21357,N_16323,N_13193);
or U21358 (N_21358,N_15663,N_15951);
xor U21359 (N_21359,N_14028,N_14462);
xor U21360 (N_21360,N_15080,N_17731);
nand U21361 (N_21361,N_14708,N_16227);
and U21362 (N_21362,N_13910,N_16957);
and U21363 (N_21363,N_12553,N_15562);
or U21364 (N_21364,N_13804,N_16068);
nand U21365 (N_21365,N_17069,N_16709);
and U21366 (N_21366,N_14680,N_17594);
nor U21367 (N_21367,N_14377,N_17344);
and U21368 (N_21368,N_17172,N_16735);
nor U21369 (N_21369,N_12985,N_13192);
xor U21370 (N_21370,N_17200,N_14667);
xnor U21371 (N_21371,N_12514,N_14937);
and U21372 (N_21372,N_16572,N_15162);
xor U21373 (N_21373,N_17760,N_17874);
and U21374 (N_21374,N_17985,N_12360);
and U21375 (N_21375,N_12022,N_13374);
nand U21376 (N_21376,N_16123,N_14915);
xor U21377 (N_21377,N_16964,N_14281);
or U21378 (N_21378,N_12781,N_16449);
nor U21379 (N_21379,N_16752,N_13094);
xor U21380 (N_21380,N_14307,N_12767);
nand U21381 (N_21381,N_14682,N_12825);
or U21382 (N_21382,N_13538,N_13119);
nand U21383 (N_21383,N_14779,N_14727);
and U21384 (N_21384,N_14074,N_14359);
xor U21385 (N_21385,N_17282,N_14605);
nor U21386 (N_21386,N_14119,N_12617);
nor U21387 (N_21387,N_15004,N_15297);
nand U21388 (N_21388,N_14097,N_15074);
xnor U21389 (N_21389,N_17274,N_15516);
nand U21390 (N_21390,N_17278,N_13563);
xor U21391 (N_21391,N_12904,N_17257);
nand U21392 (N_21392,N_12666,N_12752);
nand U21393 (N_21393,N_14567,N_17950);
nand U21394 (N_21394,N_16777,N_17024);
xor U21395 (N_21395,N_13836,N_14350);
xor U21396 (N_21396,N_16012,N_13747);
and U21397 (N_21397,N_16916,N_14503);
nor U21398 (N_21398,N_14024,N_15892);
nor U21399 (N_21399,N_16557,N_17477);
xor U21400 (N_21400,N_13737,N_13442);
and U21401 (N_21401,N_14229,N_17031);
and U21402 (N_21402,N_16937,N_16753);
nor U21403 (N_21403,N_13186,N_17169);
xor U21404 (N_21404,N_15218,N_12535);
xor U21405 (N_21405,N_15310,N_17030);
xnor U21406 (N_21406,N_13058,N_15783);
or U21407 (N_21407,N_14440,N_15902);
and U21408 (N_21408,N_16334,N_17291);
xnor U21409 (N_21409,N_12441,N_12185);
nand U21410 (N_21410,N_12290,N_13841);
xor U21411 (N_21411,N_13967,N_13554);
xor U21412 (N_21412,N_15762,N_17015);
and U21413 (N_21413,N_14533,N_17135);
and U21414 (N_21414,N_16766,N_14341);
xnor U21415 (N_21415,N_12841,N_17534);
nor U21416 (N_21416,N_16966,N_17178);
nor U21417 (N_21417,N_14256,N_12004);
or U21418 (N_21418,N_16995,N_13467);
nand U21419 (N_21419,N_17116,N_12375);
nor U21420 (N_21420,N_15147,N_15985);
nand U21421 (N_21421,N_12836,N_12657);
and U21422 (N_21422,N_17534,N_13408);
or U21423 (N_21423,N_12329,N_13202);
or U21424 (N_21424,N_12144,N_12315);
nor U21425 (N_21425,N_15978,N_15960);
xnor U21426 (N_21426,N_12545,N_12729);
nor U21427 (N_21427,N_15063,N_16409);
or U21428 (N_21428,N_16600,N_15687);
and U21429 (N_21429,N_14328,N_17276);
and U21430 (N_21430,N_13483,N_13164);
and U21431 (N_21431,N_14240,N_12253);
nor U21432 (N_21432,N_13132,N_14642);
and U21433 (N_21433,N_14398,N_13924);
or U21434 (N_21434,N_17550,N_17463);
nand U21435 (N_21435,N_17238,N_17403);
nor U21436 (N_21436,N_13053,N_12320);
nor U21437 (N_21437,N_17184,N_12335);
xnor U21438 (N_21438,N_16750,N_15560);
nor U21439 (N_21439,N_17095,N_16686);
nor U21440 (N_21440,N_12133,N_17725);
nand U21441 (N_21441,N_12952,N_15536);
or U21442 (N_21442,N_13474,N_17409);
nand U21443 (N_21443,N_14377,N_17463);
nor U21444 (N_21444,N_16945,N_16959);
or U21445 (N_21445,N_13835,N_13642);
xnor U21446 (N_21446,N_13263,N_15419);
nand U21447 (N_21447,N_12620,N_15405);
and U21448 (N_21448,N_17497,N_14215);
nor U21449 (N_21449,N_16916,N_12778);
xor U21450 (N_21450,N_13425,N_17997);
xnor U21451 (N_21451,N_15299,N_16528);
xor U21452 (N_21452,N_14694,N_12714);
or U21453 (N_21453,N_13075,N_15210);
or U21454 (N_21454,N_13862,N_15265);
nand U21455 (N_21455,N_13169,N_16741);
or U21456 (N_21456,N_15913,N_16955);
and U21457 (N_21457,N_14214,N_13027);
or U21458 (N_21458,N_12710,N_15861);
or U21459 (N_21459,N_13725,N_16079);
xnor U21460 (N_21460,N_13106,N_14564);
xor U21461 (N_21461,N_15261,N_12153);
or U21462 (N_21462,N_14738,N_12738);
nand U21463 (N_21463,N_17873,N_16452);
xor U21464 (N_21464,N_16090,N_15930);
or U21465 (N_21465,N_17813,N_13786);
or U21466 (N_21466,N_16136,N_14707);
nand U21467 (N_21467,N_15703,N_13270);
xnor U21468 (N_21468,N_16505,N_14423);
xnor U21469 (N_21469,N_17432,N_16797);
nor U21470 (N_21470,N_15037,N_17001);
xor U21471 (N_21471,N_15963,N_13832);
or U21472 (N_21472,N_15949,N_15023);
or U21473 (N_21473,N_14980,N_12330);
nor U21474 (N_21474,N_14164,N_16823);
nand U21475 (N_21475,N_15159,N_12156);
nand U21476 (N_21476,N_17908,N_14863);
nand U21477 (N_21477,N_12525,N_12897);
xnor U21478 (N_21478,N_13872,N_14053);
xor U21479 (N_21479,N_17432,N_16206);
nor U21480 (N_21480,N_17378,N_17537);
nor U21481 (N_21481,N_16968,N_12506);
nand U21482 (N_21482,N_17160,N_17550);
and U21483 (N_21483,N_17880,N_12318);
and U21484 (N_21484,N_12937,N_14404);
xor U21485 (N_21485,N_12503,N_14902);
nand U21486 (N_21486,N_14361,N_14860);
and U21487 (N_21487,N_17677,N_17407);
nand U21488 (N_21488,N_16654,N_12724);
or U21489 (N_21489,N_12603,N_13099);
nor U21490 (N_21490,N_15004,N_14186);
xor U21491 (N_21491,N_14805,N_14189);
xnor U21492 (N_21492,N_17598,N_16336);
nor U21493 (N_21493,N_12791,N_13284);
or U21494 (N_21494,N_17529,N_17587);
or U21495 (N_21495,N_15232,N_14738);
or U21496 (N_21496,N_15653,N_12593);
nand U21497 (N_21497,N_14797,N_15456);
or U21498 (N_21498,N_14432,N_14402);
nand U21499 (N_21499,N_14216,N_14068);
and U21500 (N_21500,N_12418,N_12621);
and U21501 (N_21501,N_14178,N_17489);
nand U21502 (N_21502,N_13098,N_15586);
nor U21503 (N_21503,N_15227,N_13328);
or U21504 (N_21504,N_16303,N_17186);
or U21505 (N_21505,N_17820,N_17628);
nor U21506 (N_21506,N_14260,N_17935);
or U21507 (N_21507,N_15680,N_14632);
xor U21508 (N_21508,N_13131,N_12330);
or U21509 (N_21509,N_12897,N_16563);
nor U21510 (N_21510,N_17985,N_12209);
or U21511 (N_21511,N_16775,N_13310);
or U21512 (N_21512,N_17697,N_17609);
xor U21513 (N_21513,N_14517,N_14969);
or U21514 (N_21514,N_14034,N_17538);
and U21515 (N_21515,N_16663,N_15920);
nand U21516 (N_21516,N_14151,N_12971);
nor U21517 (N_21517,N_16307,N_16752);
nor U21518 (N_21518,N_17505,N_12264);
or U21519 (N_21519,N_12969,N_12542);
and U21520 (N_21520,N_17850,N_17340);
and U21521 (N_21521,N_16338,N_14104);
and U21522 (N_21522,N_14832,N_13152);
nand U21523 (N_21523,N_15224,N_14918);
xor U21524 (N_21524,N_17965,N_17746);
or U21525 (N_21525,N_14326,N_15586);
nor U21526 (N_21526,N_12865,N_15432);
nand U21527 (N_21527,N_15261,N_13075);
xnor U21528 (N_21528,N_12951,N_17079);
nand U21529 (N_21529,N_13778,N_15764);
nor U21530 (N_21530,N_15616,N_14833);
nand U21531 (N_21531,N_13766,N_15495);
or U21532 (N_21532,N_14070,N_16894);
nor U21533 (N_21533,N_13897,N_17545);
nor U21534 (N_21534,N_12739,N_17112);
nand U21535 (N_21535,N_14313,N_12876);
or U21536 (N_21536,N_14954,N_14211);
xor U21537 (N_21537,N_13585,N_16719);
nand U21538 (N_21538,N_15002,N_16988);
nor U21539 (N_21539,N_14569,N_14874);
nor U21540 (N_21540,N_13988,N_13712);
xor U21541 (N_21541,N_14523,N_17304);
or U21542 (N_21542,N_13606,N_12000);
and U21543 (N_21543,N_15844,N_14177);
nand U21544 (N_21544,N_15359,N_16390);
xnor U21545 (N_21545,N_17521,N_13774);
nor U21546 (N_21546,N_17394,N_15489);
nand U21547 (N_21547,N_12986,N_17218);
nand U21548 (N_21548,N_13803,N_15400);
nor U21549 (N_21549,N_17492,N_12674);
and U21550 (N_21550,N_14778,N_15727);
nand U21551 (N_21551,N_17547,N_16931);
xor U21552 (N_21552,N_16875,N_17289);
nor U21553 (N_21553,N_12671,N_17926);
xor U21554 (N_21554,N_13814,N_13721);
nand U21555 (N_21555,N_17978,N_12711);
and U21556 (N_21556,N_17638,N_15097);
or U21557 (N_21557,N_14377,N_13932);
nand U21558 (N_21558,N_17386,N_12243);
xor U21559 (N_21559,N_15913,N_15303);
and U21560 (N_21560,N_17580,N_15856);
or U21561 (N_21561,N_17467,N_15057);
nand U21562 (N_21562,N_16669,N_13570);
and U21563 (N_21563,N_13981,N_17333);
and U21564 (N_21564,N_15579,N_17742);
nand U21565 (N_21565,N_14775,N_15259);
nand U21566 (N_21566,N_15440,N_16727);
xnor U21567 (N_21567,N_17196,N_16335);
or U21568 (N_21568,N_15458,N_14853);
xor U21569 (N_21569,N_16506,N_12184);
nand U21570 (N_21570,N_15688,N_13529);
nor U21571 (N_21571,N_17343,N_16235);
nor U21572 (N_21572,N_15678,N_12362);
xor U21573 (N_21573,N_14065,N_14491);
xnor U21574 (N_21574,N_17724,N_16522);
nor U21575 (N_21575,N_12714,N_15507);
or U21576 (N_21576,N_13502,N_15223);
nor U21577 (N_21577,N_14063,N_15374);
nand U21578 (N_21578,N_15198,N_13854);
or U21579 (N_21579,N_12334,N_13589);
nand U21580 (N_21580,N_17863,N_13602);
nor U21581 (N_21581,N_15423,N_12362);
nor U21582 (N_21582,N_13072,N_15229);
and U21583 (N_21583,N_12635,N_16187);
and U21584 (N_21584,N_12302,N_15871);
nand U21585 (N_21585,N_13720,N_14309);
nor U21586 (N_21586,N_16986,N_12222);
and U21587 (N_21587,N_17322,N_12402);
or U21588 (N_21588,N_13863,N_12034);
and U21589 (N_21589,N_15038,N_16250);
nor U21590 (N_21590,N_17203,N_12887);
nand U21591 (N_21591,N_13520,N_16711);
nor U21592 (N_21592,N_13495,N_13182);
and U21593 (N_21593,N_17036,N_14157);
and U21594 (N_21594,N_15334,N_13195);
and U21595 (N_21595,N_16970,N_12560);
nor U21596 (N_21596,N_12667,N_16030);
nand U21597 (N_21597,N_16989,N_15260);
and U21598 (N_21598,N_13118,N_14974);
nor U21599 (N_21599,N_15508,N_13319);
nand U21600 (N_21600,N_13023,N_12812);
nor U21601 (N_21601,N_15628,N_16191);
nand U21602 (N_21602,N_15077,N_16337);
nor U21603 (N_21603,N_16220,N_14855);
and U21604 (N_21604,N_15728,N_12318);
or U21605 (N_21605,N_13432,N_17062);
xnor U21606 (N_21606,N_14612,N_16023);
xor U21607 (N_21607,N_14424,N_13335);
and U21608 (N_21608,N_14238,N_13452);
nor U21609 (N_21609,N_12347,N_14670);
nand U21610 (N_21610,N_16700,N_16885);
nor U21611 (N_21611,N_16583,N_12224);
and U21612 (N_21612,N_13499,N_14303);
nand U21613 (N_21613,N_15919,N_14525);
nor U21614 (N_21614,N_17854,N_16301);
and U21615 (N_21615,N_13773,N_14563);
xnor U21616 (N_21616,N_15267,N_17169);
and U21617 (N_21617,N_14253,N_13368);
nor U21618 (N_21618,N_17091,N_12274);
and U21619 (N_21619,N_16078,N_17990);
nand U21620 (N_21620,N_14166,N_13009);
xnor U21621 (N_21621,N_12336,N_13231);
xor U21622 (N_21622,N_16936,N_12024);
or U21623 (N_21623,N_15822,N_12145);
and U21624 (N_21624,N_16545,N_13119);
nor U21625 (N_21625,N_13686,N_15190);
nor U21626 (N_21626,N_17313,N_17386);
nand U21627 (N_21627,N_12536,N_15298);
nor U21628 (N_21628,N_15066,N_12590);
nor U21629 (N_21629,N_13623,N_17488);
nand U21630 (N_21630,N_14236,N_12537);
xor U21631 (N_21631,N_15596,N_15966);
nor U21632 (N_21632,N_16666,N_15729);
or U21633 (N_21633,N_14311,N_15405);
xnor U21634 (N_21634,N_15403,N_15976);
xnor U21635 (N_21635,N_13199,N_16326);
nand U21636 (N_21636,N_12174,N_14712);
and U21637 (N_21637,N_12010,N_12048);
and U21638 (N_21638,N_15238,N_17968);
xnor U21639 (N_21639,N_14865,N_17134);
xor U21640 (N_21640,N_13799,N_14006);
or U21641 (N_21641,N_15471,N_17528);
nand U21642 (N_21642,N_17079,N_13958);
nand U21643 (N_21643,N_14651,N_12715);
xor U21644 (N_21644,N_13373,N_17864);
or U21645 (N_21645,N_12858,N_14629);
xor U21646 (N_21646,N_16628,N_12497);
xnor U21647 (N_21647,N_16442,N_15043);
and U21648 (N_21648,N_13496,N_12566);
nor U21649 (N_21649,N_15720,N_12227);
or U21650 (N_21650,N_16289,N_14693);
nor U21651 (N_21651,N_14243,N_14408);
nor U21652 (N_21652,N_14333,N_16288);
or U21653 (N_21653,N_13158,N_17196);
xor U21654 (N_21654,N_14208,N_13861);
or U21655 (N_21655,N_16926,N_14154);
or U21656 (N_21656,N_16382,N_13113);
or U21657 (N_21657,N_14849,N_13877);
xnor U21658 (N_21658,N_13160,N_14030);
and U21659 (N_21659,N_12070,N_12541);
nor U21660 (N_21660,N_13798,N_15888);
nand U21661 (N_21661,N_16306,N_13987);
xnor U21662 (N_21662,N_16196,N_15479);
or U21663 (N_21663,N_15854,N_17195);
nor U21664 (N_21664,N_15545,N_13704);
nand U21665 (N_21665,N_13783,N_15371);
xnor U21666 (N_21666,N_12972,N_15768);
or U21667 (N_21667,N_15498,N_15096);
nand U21668 (N_21668,N_13528,N_14328);
or U21669 (N_21669,N_16110,N_17945);
xnor U21670 (N_21670,N_16711,N_15973);
xor U21671 (N_21671,N_13290,N_13520);
nor U21672 (N_21672,N_17707,N_15865);
nor U21673 (N_21673,N_12767,N_13890);
and U21674 (N_21674,N_12617,N_14080);
nand U21675 (N_21675,N_15064,N_15541);
or U21676 (N_21676,N_14115,N_17763);
xor U21677 (N_21677,N_16772,N_13419);
xnor U21678 (N_21678,N_17935,N_14732);
or U21679 (N_21679,N_16313,N_16630);
xnor U21680 (N_21680,N_17789,N_14159);
or U21681 (N_21681,N_15741,N_13617);
nor U21682 (N_21682,N_17642,N_13712);
nor U21683 (N_21683,N_13318,N_15714);
nor U21684 (N_21684,N_17752,N_15759);
nand U21685 (N_21685,N_15968,N_13637);
nand U21686 (N_21686,N_15590,N_15210);
or U21687 (N_21687,N_13587,N_15915);
nand U21688 (N_21688,N_14085,N_15429);
xnor U21689 (N_21689,N_13435,N_13893);
nand U21690 (N_21690,N_14637,N_13265);
or U21691 (N_21691,N_15323,N_15593);
or U21692 (N_21692,N_16592,N_13647);
nand U21693 (N_21693,N_16155,N_13307);
nor U21694 (N_21694,N_15190,N_12078);
and U21695 (N_21695,N_16578,N_15239);
xor U21696 (N_21696,N_16062,N_17325);
xor U21697 (N_21697,N_17924,N_13238);
nor U21698 (N_21698,N_13816,N_13336);
nor U21699 (N_21699,N_17016,N_16359);
xor U21700 (N_21700,N_15214,N_14919);
nand U21701 (N_21701,N_16033,N_12091);
xor U21702 (N_21702,N_16567,N_17420);
or U21703 (N_21703,N_14618,N_16587);
or U21704 (N_21704,N_15259,N_15311);
nor U21705 (N_21705,N_13100,N_17321);
xnor U21706 (N_21706,N_17584,N_12173);
and U21707 (N_21707,N_17739,N_15159);
nor U21708 (N_21708,N_17707,N_15139);
nand U21709 (N_21709,N_17683,N_13309);
or U21710 (N_21710,N_12305,N_17459);
or U21711 (N_21711,N_13546,N_12077);
nor U21712 (N_21712,N_17216,N_15784);
nand U21713 (N_21713,N_14482,N_13192);
xnor U21714 (N_21714,N_16263,N_16554);
nor U21715 (N_21715,N_17395,N_17628);
nand U21716 (N_21716,N_14613,N_17252);
xor U21717 (N_21717,N_14559,N_13270);
or U21718 (N_21718,N_16102,N_17359);
or U21719 (N_21719,N_15405,N_13294);
xor U21720 (N_21720,N_14678,N_15982);
or U21721 (N_21721,N_15077,N_15629);
nand U21722 (N_21722,N_13993,N_13334);
and U21723 (N_21723,N_13332,N_14016);
xnor U21724 (N_21724,N_14534,N_15544);
nor U21725 (N_21725,N_17333,N_12279);
or U21726 (N_21726,N_16162,N_12393);
xor U21727 (N_21727,N_12810,N_16985);
or U21728 (N_21728,N_12481,N_13118);
or U21729 (N_21729,N_17312,N_15156);
xnor U21730 (N_21730,N_12148,N_12172);
nand U21731 (N_21731,N_12866,N_13825);
xnor U21732 (N_21732,N_13191,N_17112);
and U21733 (N_21733,N_17699,N_17659);
or U21734 (N_21734,N_12248,N_16977);
nor U21735 (N_21735,N_16758,N_15807);
and U21736 (N_21736,N_13318,N_17570);
nor U21737 (N_21737,N_17763,N_17542);
nand U21738 (N_21738,N_12479,N_16108);
xor U21739 (N_21739,N_16478,N_12299);
xnor U21740 (N_21740,N_13824,N_17257);
or U21741 (N_21741,N_17758,N_17888);
or U21742 (N_21742,N_13152,N_16806);
and U21743 (N_21743,N_13019,N_17663);
and U21744 (N_21744,N_14985,N_12459);
xnor U21745 (N_21745,N_17500,N_15141);
nor U21746 (N_21746,N_15492,N_17330);
and U21747 (N_21747,N_15674,N_16414);
nand U21748 (N_21748,N_12854,N_15336);
xor U21749 (N_21749,N_12167,N_15250);
nand U21750 (N_21750,N_12193,N_14675);
or U21751 (N_21751,N_17667,N_12961);
and U21752 (N_21752,N_16971,N_12100);
xnor U21753 (N_21753,N_17493,N_16608);
or U21754 (N_21754,N_14099,N_14901);
nor U21755 (N_21755,N_14973,N_13216);
nor U21756 (N_21756,N_17351,N_15750);
nand U21757 (N_21757,N_17605,N_15691);
and U21758 (N_21758,N_15350,N_12008);
and U21759 (N_21759,N_15751,N_16320);
nor U21760 (N_21760,N_14685,N_17567);
nor U21761 (N_21761,N_15943,N_13631);
nor U21762 (N_21762,N_14681,N_14885);
and U21763 (N_21763,N_14442,N_15490);
nand U21764 (N_21764,N_13818,N_12078);
and U21765 (N_21765,N_12194,N_16994);
nand U21766 (N_21766,N_13758,N_12704);
xnor U21767 (N_21767,N_15437,N_12211);
nand U21768 (N_21768,N_14066,N_12598);
xnor U21769 (N_21769,N_14900,N_16122);
nor U21770 (N_21770,N_12997,N_12531);
or U21771 (N_21771,N_15167,N_12048);
nor U21772 (N_21772,N_13264,N_17299);
nand U21773 (N_21773,N_13160,N_17584);
nor U21774 (N_21774,N_14471,N_14685);
nor U21775 (N_21775,N_12563,N_15083);
and U21776 (N_21776,N_13325,N_15722);
or U21777 (N_21777,N_14912,N_15275);
nand U21778 (N_21778,N_16909,N_16521);
and U21779 (N_21779,N_16093,N_17494);
or U21780 (N_21780,N_13511,N_16797);
or U21781 (N_21781,N_16241,N_13706);
and U21782 (N_21782,N_15500,N_12742);
nor U21783 (N_21783,N_17897,N_17640);
nor U21784 (N_21784,N_13719,N_17668);
xnor U21785 (N_21785,N_13183,N_14864);
or U21786 (N_21786,N_12192,N_16088);
and U21787 (N_21787,N_13458,N_17779);
nand U21788 (N_21788,N_16960,N_14689);
nor U21789 (N_21789,N_14583,N_17147);
xnor U21790 (N_21790,N_13137,N_16951);
nand U21791 (N_21791,N_14698,N_17663);
xor U21792 (N_21792,N_12328,N_17915);
xnor U21793 (N_21793,N_15778,N_13213);
or U21794 (N_21794,N_17580,N_16733);
or U21795 (N_21795,N_16080,N_13371);
nand U21796 (N_21796,N_12952,N_13652);
and U21797 (N_21797,N_14536,N_13087);
xor U21798 (N_21798,N_14813,N_12244);
or U21799 (N_21799,N_16243,N_13789);
or U21800 (N_21800,N_16634,N_12913);
xnor U21801 (N_21801,N_17054,N_12434);
and U21802 (N_21802,N_16166,N_16035);
xnor U21803 (N_21803,N_14194,N_17563);
xnor U21804 (N_21804,N_13242,N_16457);
or U21805 (N_21805,N_12309,N_17421);
nand U21806 (N_21806,N_17446,N_16939);
nor U21807 (N_21807,N_14717,N_15908);
xor U21808 (N_21808,N_17434,N_15864);
and U21809 (N_21809,N_14033,N_17357);
nand U21810 (N_21810,N_17185,N_14424);
and U21811 (N_21811,N_15887,N_15998);
xnor U21812 (N_21812,N_12043,N_16836);
xnor U21813 (N_21813,N_13447,N_16493);
xnor U21814 (N_21814,N_12004,N_12309);
nor U21815 (N_21815,N_13709,N_13146);
or U21816 (N_21816,N_16044,N_16763);
nand U21817 (N_21817,N_14978,N_14475);
or U21818 (N_21818,N_12974,N_15843);
or U21819 (N_21819,N_16344,N_12673);
xnor U21820 (N_21820,N_12038,N_15875);
nor U21821 (N_21821,N_16664,N_12258);
nand U21822 (N_21822,N_16631,N_16069);
xnor U21823 (N_21823,N_16482,N_16500);
nand U21824 (N_21824,N_16819,N_12638);
or U21825 (N_21825,N_16797,N_15527);
xnor U21826 (N_21826,N_14323,N_14383);
xnor U21827 (N_21827,N_13298,N_14897);
nand U21828 (N_21828,N_15195,N_14422);
nor U21829 (N_21829,N_17409,N_17672);
and U21830 (N_21830,N_12146,N_14200);
xor U21831 (N_21831,N_15962,N_14607);
nor U21832 (N_21832,N_14729,N_15119);
and U21833 (N_21833,N_16820,N_15339);
nand U21834 (N_21834,N_15582,N_13070);
nand U21835 (N_21835,N_17824,N_15296);
xor U21836 (N_21836,N_13943,N_14473);
xnor U21837 (N_21837,N_16039,N_16996);
xor U21838 (N_21838,N_16143,N_16550);
and U21839 (N_21839,N_17765,N_15823);
xor U21840 (N_21840,N_13405,N_15492);
xnor U21841 (N_21841,N_12560,N_13908);
nand U21842 (N_21842,N_16964,N_13261);
or U21843 (N_21843,N_17557,N_14204);
nand U21844 (N_21844,N_17498,N_13619);
and U21845 (N_21845,N_15375,N_17313);
xnor U21846 (N_21846,N_17221,N_15677);
xor U21847 (N_21847,N_16774,N_12452);
xor U21848 (N_21848,N_13597,N_13409);
nand U21849 (N_21849,N_16846,N_17018);
nand U21850 (N_21850,N_15297,N_14509);
and U21851 (N_21851,N_12275,N_14510);
or U21852 (N_21852,N_14074,N_15775);
xnor U21853 (N_21853,N_15066,N_13990);
or U21854 (N_21854,N_17873,N_12831);
nand U21855 (N_21855,N_13659,N_14988);
and U21856 (N_21856,N_14346,N_12693);
or U21857 (N_21857,N_12511,N_12604);
nand U21858 (N_21858,N_13443,N_12369);
nor U21859 (N_21859,N_14466,N_13853);
and U21860 (N_21860,N_15009,N_13104);
nor U21861 (N_21861,N_14955,N_17941);
nor U21862 (N_21862,N_12524,N_14662);
and U21863 (N_21863,N_15439,N_17333);
nand U21864 (N_21864,N_17807,N_13871);
nand U21865 (N_21865,N_13272,N_12591);
nor U21866 (N_21866,N_15015,N_15610);
xor U21867 (N_21867,N_15953,N_12689);
xor U21868 (N_21868,N_13621,N_13187);
xnor U21869 (N_21869,N_17199,N_15702);
nand U21870 (N_21870,N_14068,N_13502);
xor U21871 (N_21871,N_13048,N_17541);
nor U21872 (N_21872,N_15773,N_16005);
or U21873 (N_21873,N_14174,N_15323);
xnor U21874 (N_21874,N_14600,N_15402);
or U21875 (N_21875,N_16767,N_15569);
and U21876 (N_21876,N_15452,N_12809);
xnor U21877 (N_21877,N_17020,N_15815);
xnor U21878 (N_21878,N_12719,N_15681);
nor U21879 (N_21879,N_13456,N_16878);
nand U21880 (N_21880,N_15155,N_12063);
and U21881 (N_21881,N_14886,N_13442);
nor U21882 (N_21882,N_13301,N_12465);
and U21883 (N_21883,N_13109,N_15404);
and U21884 (N_21884,N_16045,N_12827);
and U21885 (N_21885,N_14361,N_13587);
xnor U21886 (N_21886,N_12403,N_14847);
nor U21887 (N_21887,N_15288,N_14162);
nand U21888 (N_21888,N_13690,N_17525);
nor U21889 (N_21889,N_15603,N_14336);
xor U21890 (N_21890,N_17071,N_13940);
xor U21891 (N_21891,N_15804,N_16100);
nand U21892 (N_21892,N_15098,N_16591);
nor U21893 (N_21893,N_14711,N_15421);
or U21894 (N_21894,N_14050,N_14830);
xnor U21895 (N_21895,N_12495,N_16089);
xnor U21896 (N_21896,N_14759,N_15440);
or U21897 (N_21897,N_14505,N_17754);
or U21898 (N_21898,N_13697,N_16227);
or U21899 (N_21899,N_13280,N_16812);
xor U21900 (N_21900,N_15480,N_17562);
nand U21901 (N_21901,N_16970,N_13946);
nand U21902 (N_21902,N_16220,N_13120);
nor U21903 (N_21903,N_17877,N_15576);
and U21904 (N_21904,N_13695,N_16375);
xor U21905 (N_21905,N_15900,N_13409);
and U21906 (N_21906,N_12280,N_15404);
or U21907 (N_21907,N_17072,N_14309);
and U21908 (N_21908,N_17976,N_15578);
and U21909 (N_21909,N_13356,N_17802);
nand U21910 (N_21910,N_17999,N_13263);
or U21911 (N_21911,N_15602,N_14102);
nand U21912 (N_21912,N_13677,N_16098);
and U21913 (N_21913,N_14792,N_12565);
or U21914 (N_21914,N_12808,N_12079);
or U21915 (N_21915,N_15152,N_12113);
nor U21916 (N_21916,N_16328,N_16090);
and U21917 (N_21917,N_12415,N_12090);
and U21918 (N_21918,N_15716,N_15061);
nor U21919 (N_21919,N_15506,N_16418);
nand U21920 (N_21920,N_15839,N_15008);
or U21921 (N_21921,N_12380,N_15015);
or U21922 (N_21922,N_13096,N_16425);
or U21923 (N_21923,N_12749,N_12947);
and U21924 (N_21924,N_12966,N_12088);
and U21925 (N_21925,N_14333,N_13489);
nor U21926 (N_21926,N_16029,N_17364);
nor U21927 (N_21927,N_14210,N_15867);
or U21928 (N_21928,N_12386,N_15915);
and U21929 (N_21929,N_15320,N_15715);
nor U21930 (N_21930,N_17564,N_15009);
or U21931 (N_21931,N_15043,N_15243);
or U21932 (N_21932,N_17573,N_15177);
nand U21933 (N_21933,N_17380,N_14671);
and U21934 (N_21934,N_14452,N_14584);
nor U21935 (N_21935,N_14231,N_13309);
and U21936 (N_21936,N_17629,N_15003);
nor U21937 (N_21937,N_12697,N_17636);
xor U21938 (N_21938,N_14435,N_16314);
nor U21939 (N_21939,N_12938,N_14942);
and U21940 (N_21940,N_15445,N_13417);
xnor U21941 (N_21941,N_17277,N_16606);
and U21942 (N_21942,N_13560,N_16761);
or U21943 (N_21943,N_12380,N_14496);
nand U21944 (N_21944,N_14615,N_16337);
nand U21945 (N_21945,N_15771,N_16481);
nand U21946 (N_21946,N_15894,N_13626);
and U21947 (N_21947,N_14070,N_12146);
nand U21948 (N_21948,N_14464,N_12428);
nand U21949 (N_21949,N_14597,N_13524);
nor U21950 (N_21950,N_14664,N_14099);
xor U21951 (N_21951,N_13745,N_13808);
xor U21952 (N_21952,N_16451,N_17799);
nor U21953 (N_21953,N_15927,N_15235);
nor U21954 (N_21954,N_12591,N_13355);
and U21955 (N_21955,N_16501,N_17928);
and U21956 (N_21956,N_14082,N_12215);
or U21957 (N_21957,N_17005,N_16734);
and U21958 (N_21958,N_17325,N_15118);
nor U21959 (N_21959,N_14811,N_16987);
nor U21960 (N_21960,N_14767,N_17281);
xor U21961 (N_21961,N_12164,N_14479);
xnor U21962 (N_21962,N_12372,N_15574);
nand U21963 (N_21963,N_13821,N_12728);
and U21964 (N_21964,N_17427,N_13542);
nor U21965 (N_21965,N_15842,N_17521);
and U21966 (N_21966,N_16286,N_17497);
xnor U21967 (N_21967,N_13755,N_14092);
xnor U21968 (N_21968,N_16360,N_14007);
or U21969 (N_21969,N_13367,N_16388);
and U21970 (N_21970,N_12623,N_14305);
nand U21971 (N_21971,N_16655,N_17959);
xor U21972 (N_21972,N_13216,N_15625);
nor U21973 (N_21973,N_16791,N_13720);
or U21974 (N_21974,N_16050,N_17580);
and U21975 (N_21975,N_17894,N_17322);
nor U21976 (N_21976,N_14343,N_15688);
and U21977 (N_21977,N_15047,N_17377);
and U21978 (N_21978,N_15422,N_12127);
nand U21979 (N_21979,N_12752,N_12028);
and U21980 (N_21980,N_14492,N_15915);
nor U21981 (N_21981,N_12841,N_13067);
xnor U21982 (N_21982,N_17651,N_15010);
nor U21983 (N_21983,N_16988,N_13814);
nor U21984 (N_21984,N_14221,N_13851);
or U21985 (N_21985,N_16794,N_16304);
nand U21986 (N_21986,N_14543,N_15574);
or U21987 (N_21987,N_15188,N_13736);
xnor U21988 (N_21988,N_13767,N_15611);
nor U21989 (N_21989,N_16679,N_17917);
nand U21990 (N_21990,N_13591,N_14374);
nor U21991 (N_21991,N_15746,N_16453);
xor U21992 (N_21992,N_15648,N_14527);
nor U21993 (N_21993,N_16487,N_14271);
and U21994 (N_21994,N_16715,N_17091);
xor U21995 (N_21995,N_13277,N_13043);
nand U21996 (N_21996,N_14654,N_15989);
and U21997 (N_21997,N_14948,N_14541);
nor U21998 (N_21998,N_12010,N_16857);
and U21999 (N_21999,N_17008,N_12197);
or U22000 (N_22000,N_17056,N_12103);
and U22001 (N_22001,N_14979,N_12998);
and U22002 (N_22002,N_12118,N_14240);
nor U22003 (N_22003,N_15183,N_12963);
and U22004 (N_22004,N_16465,N_17158);
nand U22005 (N_22005,N_12343,N_16448);
nand U22006 (N_22006,N_12234,N_13703);
and U22007 (N_22007,N_13199,N_17649);
or U22008 (N_22008,N_15604,N_12670);
or U22009 (N_22009,N_14448,N_15057);
or U22010 (N_22010,N_14350,N_14351);
or U22011 (N_22011,N_12290,N_15130);
or U22012 (N_22012,N_13140,N_14250);
and U22013 (N_22013,N_14818,N_16311);
xor U22014 (N_22014,N_13922,N_15421);
and U22015 (N_22015,N_17922,N_15094);
nor U22016 (N_22016,N_17466,N_16771);
and U22017 (N_22017,N_12507,N_13374);
and U22018 (N_22018,N_15887,N_13345);
xnor U22019 (N_22019,N_15063,N_15512);
or U22020 (N_22020,N_14074,N_16188);
xor U22021 (N_22021,N_14086,N_15729);
and U22022 (N_22022,N_17844,N_12306);
nor U22023 (N_22023,N_15259,N_13832);
xnor U22024 (N_22024,N_17455,N_17331);
nand U22025 (N_22025,N_13083,N_14762);
nand U22026 (N_22026,N_12332,N_12706);
xor U22027 (N_22027,N_14261,N_12020);
nor U22028 (N_22028,N_16904,N_15654);
or U22029 (N_22029,N_17190,N_16831);
xor U22030 (N_22030,N_12106,N_17528);
xor U22031 (N_22031,N_12840,N_13028);
and U22032 (N_22032,N_17915,N_12187);
or U22033 (N_22033,N_16184,N_13251);
or U22034 (N_22034,N_15413,N_16755);
xnor U22035 (N_22035,N_15684,N_15631);
nand U22036 (N_22036,N_12883,N_16962);
or U22037 (N_22037,N_16496,N_12219);
or U22038 (N_22038,N_16936,N_14267);
and U22039 (N_22039,N_17755,N_14332);
nor U22040 (N_22040,N_15894,N_14507);
nor U22041 (N_22041,N_14065,N_15926);
nand U22042 (N_22042,N_12242,N_12012);
or U22043 (N_22043,N_16273,N_17221);
nor U22044 (N_22044,N_13587,N_12724);
or U22045 (N_22045,N_17384,N_16267);
and U22046 (N_22046,N_15530,N_16175);
or U22047 (N_22047,N_15978,N_15015);
xor U22048 (N_22048,N_12664,N_15471);
xor U22049 (N_22049,N_14126,N_12163);
nor U22050 (N_22050,N_16940,N_16610);
nand U22051 (N_22051,N_13068,N_16557);
nor U22052 (N_22052,N_17671,N_16132);
and U22053 (N_22053,N_14669,N_14079);
or U22054 (N_22054,N_17384,N_14502);
and U22055 (N_22055,N_13685,N_13499);
and U22056 (N_22056,N_16785,N_14142);
or U22057 (N_22057,N_15982,N_13154);
or U22058 (N_22058,N_14949,N_12787);
and U22059 (N_22059,N_13234,N_14358);
nand U22060 (N_22060,N_13800,N_16916);
xor U22061 (N_22061,N_17109,N_16128);
nor U22062 (N_22062,N_15645,N_14050);
xnor U22063 (N_22063,N_16735,N_16634);
xor U22064 (N_22064,N_17671,N_12560);
nand U22065 (N_22065,N_16382,N_16429);
and U22066 (N_22066,N_15512,N_13975);
nor U22067 (N_22067,N_15375,N_12550);
xnor U22068 (N_22068,N_13692,N_16122);
nand U22069 (N_22069,N_16937,N_14395);
nand U22070 (N_22070,N_16119,N_15260);
and U22071 (N_22071,N_13376,N_15666);
or U22072 (N_22072,N_13670,N_15156);
nor U22073 (N_22073,N_17494,N_17539);
xnor U22074 (N_22074,N_16941,N_16006);
nand U22075 (N_22075,N_16188,N_17230);
nand U22076 (N_22076,N_13953,N_17798);
or U22077 (N_22077,N_14280,N_16348);
nand U22078 (N_22078,N_16567,N_12314);
and U22079 (N_22079,N_13201,N_16944);
nand U22080 (N_22080,N_17746,N_15356);
xor U22081 (N_22081,N_16714,N_17511);
or U22082 (N_22082,N_15061,N_12061);
nor U22083 (N_22083,N_14186,N_13218);
xnor U22084 (N_22084,N_17467,N_15561);
xor U22085 (N_22085,N_16254,N_15176);
and U22086 (N_22086,N_17557,N_12133);
and U22087 (N_22087,N_12807,N_17752);
nor U22088 (N_22088,N_16724,N_16006);
or U22089 (N_22089,N_13275,N_16685);
nor U22090 (N_22090,N_15704,N_14388);
and U22091 (N_22091,N_15939,N_15764);
nor U22092 (N_22092,N_16965,N_13173);
nor U22093 (N_22093,N_14121,N_16114);
or U22094 (N_22094,N_14662,N_12664);
nand U22095 (N_22095,N_12425,N_14137);
xor U22096 (N_22096,N_12153,N_16003);
xnor U22097 (N_22097,N_14682,N_14530);
nand U22098 (N_22098,N_13879,N_17678);
nand U22099 (N_22099,N_12754,N_14553);
nand U22100 (N_22100,N_12590,N_17752);
and U22101 (N_22101,N_15628,N_16974);
xnor U22102 (N_22102,N_17168,N_17715);
nand U22103 (N_22103,N_13368,N_14921);
xor U22104 (N_22104,N_13723,N_12017);
xnor U22105 (N_22105,N_17466,N_12649);
xnor U22106 (N_22106,N_12119,N_16104);
nand U22107 (N_22107,N_17864,N_14370);
and U22108 (N_22108,N_13854,N_17563);
nor U22109 (N_22109,N_16085,N_14163);
xor U22110 (N_22110,N_16633,N_16574);
xnor U22111 (N_22111,N_17532,N_13348);
xnor U22112 (N_22112,N_14970,N_12381);
or U22113 (N_22113,N_17726,N_15582);
or U22114 (N_22114,N_13683,N_13409);
and U22115 (N_22115,N_16569,N_17346);
nor U22116 (N_22116,N_14747,N_14397);
and U22117 (N_22117,N_15496,N_12161);
nor U22118 (N_22118,N_12601,N_14692);
and U22119 (N_22119,N_15767,N_16400);
xnor U22120 (N_22120,N_17912,N_12440);
nand U22121 (N_22121,N_12422,N_17080);
nand U22122 (N_22122,N_15235,N_17097);
nor U22123 (N_22123,N_13287,N_15691);
or U22124 (N_22124,N_13891,N_16084);
and U22125 (N_22125,N_17233,N_14745);
or U22126 (N_22126,N_13435,N_16475);
and U22127 (N_22127,N_12480,N_17254);
nor U22128 (N_22128,N_17600,N_14172);
or U22129 (N_22129,N_15184,N_17842);
nor U22130 (N_22130,N_13961,N_16478);
nand U22131 (N_22131,N_12254,N_12749);
or U22132 (N_22132,N_13723,N_15354);
nand U22133 (N_22133,N_12365,N_13103);
and U22134 (N_22134,N_16796,N_16918);
nand U22135 (N_22135,N_15306,N_13978);
and U22136 (N_22136,N_17999,N_16295);
xnor U22137 (N_22137,N_17536,N_14039);
xor U22138 (N_22138,N_12239,N_13010);
or U22139 (N_22139,N_16250,N_17129);
or U22140 (N_22140,N_13254,N_15894);
xor U22141 (N_22141,N_17637,N_12490);
and U22142 (N_22142,N_17655,N_12508);
or U22143 (N_22143,N_12754,N_17202);
and U22144 (N_22144,N_12283,N_17219);
nand U22145 (N_22145,N_17553,N_16541);
and U22146 (N_22146,N_13735,N_12726);
xnor U22147 (N_22147,N_15473,N_16268);
and U22148 (N_22148,N_17629,N_12630);
nand U22149 (N_22149,N_17280,N_15873);
nor U22150 (N_22150,N_16190,N_12234);
nand U22151 (N_22151,N_15853,N_12378);
nor U22152 (N_22152,N_14620,N_16074);
xor U22153 (N_22153,N_16241,N_16002);
xor U22154 (N_22154,N_16975,N_14845);
xnor U22155 (N_22155,N_16449,N_13940);
nor U22156 (N_22156,N_15121,N_16840);
and U22157 (N_22157,N_13122,N_12314);
and U22158 (N_22158,N_13255,N_13395);
and U22159 (N_22159,N_17817,N_13200);
xnor U22160 (N_22160,N_17958,N_14246);
and U22161 (N_22161,N_13832,N_14533);
xor U22162 (N_22162,N_17367,N_12184);
or U22163 (N_22163,N_17309,N_13373);
nor U22164 (N_22164,N_15458,N_16553);
xor U22165 (N_22165,N_14059,N_16384);
and U22166 (N_22166,N_17150,N_14890);
nand U22167 (N_22167,N_12087,N_12596);
xnor U22168 (N_22168,N_14281,N_15838);
nor U22169 (N_22169,N_16399,N_16496);
or U22170 (N_22170,N_14805,N_16907);
nand U22171 (N_22171,N_15227,N_16452);
nor U22172 (N_22172,N_17953,N_14066);
nand U22173 (N_22173,N_17614,N_14829);
xor U22174 (N_22174,N_17868,N_15091);
nor U22175 (N_22175,N_17340,N_16175);
or U22176 (N_22176,N_12678,N_17253);
or U22177 (N_22177,N_17106,N_17448);
nand U22178 (N_22178,N_12297,N_13779);
nand U22179 (N_22179,N_15693,N_13279);
or U22180 (N_22180,N_12860,N_15993);
nand U22181 (N_22181,N_13238,N_16890);
xnor U22182 (N_22182,N_13438,N_12432);
or U22183 (N_22183,N_14021,N_15155);
xor U22184 (N_22184,N_14233,N_15245);
xor U22185 (N_22185,N_16180,N_14526);
nor U22186 (N_22186,N_12800,N_14656);
nor U22187 (N_22187,N_12478,N_13657);
nand U22188 (N_22188,N_12284,N_17865);
or U22189 (N_22189,N_12256,N_17906);
or U22190 (N_22190,N_16166,N_16099);
xor U22191 (N_22191,N_12482,N_13123);
nand U22192 (N_22192,N_12273,N_16401);
nand U22193 (N_22193,N_14259,N_13685);
xor U22194 (N_22194,N_17778,N_14100);
nor U22195 (N_22195,N_15854,N_12955);
xnor U22196 (N_22196,N_16476,N_15155);
or U22197 (N_22197,N_13746,N_14194);
and U22198 (N_22198,N_12362,N_14805);
or U22199 (N_22199,N_12413,N_13587);
xor U22200 (N_22200,N_17356,N_16855);
or U22201 (N_22201,N_12006,N_16408);
or U22202 (N_22202,N_12583,N_17049);
nor U22203 (N_22203,N_12481,N_12807);
xor U22204 (N_22204,N_14126,N_13834);
nor U22205 (N_22205,N_17404,N_13051);
and U22206 (N_22206,N_12588,N_17636);
xor U22207 (N_22207,N_12728,N_16410);
nor U22208 (N_22208,N_17539,N_14175);
and U22209 (N_22209,N_13213,N_12221);
nand U22210 (N_22210,N_13505,N_17626);
or U22211 (N_22211,N_16086,N_16540);
xor U22212 (N_22212,N_12650,N_17803);
nand U22213 (N_22213,N_15699,N_16977);
and U22214 (N_22214,N_15471,N_16834);
nand U22215 (N_22215,N_15056,N_16782);
xor U22216 (N_22216,N_16258,N_17117);
and U22217 (N_22217,N_15001,N_13753);
nor U22218 (N_22218,N_15976,N_17454);
or U22219 (N_22219,N_15092,N_12722);
nand U22220 (N_22220,N_14747,N_16282);
or U22221 (N_22221,N_15270,N_17736);
nor U22222 (N_22222,N_16880,N_14380);
xor U22223 (N_22223,N_17447,N_12536);
and U22224 (N_22224,N_14785,N_16652);
nand U22225 (N_22225,N_13366,N_13572);
nor U22226 (N_22226,N_14286,N_12104);
xor U22227 (N_22227,N_17670,N_17547);
nor U22228 (N_22228,N_14087,N_13276);
nor U22229 (N_22229,N_16875,N_13620);
xor U22230 (N_22230,N_16315,N_16222);
nor U22231 (N_22231,N_12066,N_14463);
or U22232 (N_22232,N_14347,N_12782);
or U22233 (N_22233,N_13425,N_14612);
or U22234 (N_22234,N_17824,N_12855);
or U22235 (N_22235,N_12200,N_17920);
or U22236 (N_22236,N_12237,N_15338);
xor U22237 (N_22237,N_16158,N_16575);
and U22238 (N_22238,N_15257,N_17627);
nand U22239 (N_22239,N_12503,N_14287);
and U22240 (N_22240,N_14044,N_13285);
xor U22241 (N_22241,N_16598,N_13345);
xnor U22242 (N_22242,N_16465,N_14107);
or U22243 (N_22243,N_14180,N_17726);
and U22244 (N_22244,N_15711,N_14732);
or U22245 (N_22245,N_12601,N_12903);
nand U22246 (N_22246,N_17958,N_14733);
nand U22247 (N_22247,N_16003,N_15939);
nor U22248 (N_22248,N_17535,N_12423);
xnor U22249 (N_22249,N_12730,N_16933);
xnor U22250 (N_22250,N_16165,N_12046);
nand U22251 (N_22251,N_13743,N_16405);
nor U22252 (N_22252,N_12183,N_15753);
nand U22253 (N_22253,N_16062,N_16359);
nand U22254 (N_22254,N_14649,N_17527);
xnor U22255 (N_22255,N_14018,N_13672);
and U22256 (N_22256,N_12297,N_16966);
nor U22257 (N_22257,N_13433,N_15061);
xor U22258 (N_22258,N_12153,N_14881);
xor U22259 (N_22259,N_16893,N_12600);
or U22260 (N_22260,N_15445,N_15705);
nor U22261 (N_22261,N_14321,N_13301);
and U22262 (N_22262,N_13351,N_15926);
or U22263 (N_22263,N_15891,N_15107);
and U22264 (N_22264,N_13910,N_16959);
or U22265 (N_22265,N_14652,N_17674);
xnor U22266 (N_22266,N_14348,N_15811);
nand U22267 (N_22267,N_17843,N_17844);
and U22268 (N_22268,N_13129,N_12578);
or U22269 (N_22269,N_14792,N_17551);
xor U22270 (N_22270,N_13510,N_15099);
or U22271 (N_22271,N_16714,N_16612);
nor U22272 (N_22272,N_16071,N_16951);
nor U22273 (N_22273,N_17181,N_12304);
xnor U22274 (N_22274,N_15939,N_16831);
nor U22275 (N_22275,N_16230,N_14669);
nand U22276 (N_22276,N_14240,N_13079);
nor U22277 (N_22277,N_12133,N_16047);
nor U22278 (N_22278,N_15175,N_15593);
nand U22279 (N_22279,N_12336,N_14562);
nor U22280 (N_22280,N_12986,N_12288);
nand U22281 (N_22281,N_12527,N_15747);
nor U22282 (N_22282,N_12272,N_12602);
nor U22283 (N_22283,N_12890,N_17265);
xor U22284 (N_22284,N_16148,N_13818);
nand U22285 (N_22285,N_16562,N_14118);
nor U22286 (N_22286,N_16725,N_12852);
nand U22287 (N_22287,N_14808,N_12590);
nor U22288 (N_22288,N_15576,N_17529);
and U22289 (N_22289,N_15093,N_13555);
or U22290 (N_22290,N_12568,N_17271);
nor U22291 (N_22291,N_16774,N_16102);
nor U22292 (N_22292,N_15885,N_12260);
nand U22293 (N_22293,N_14996,N_12079);
or U22294 (N_22294,N_14295,N_15414);
or U22295 (N_22295,N_16458,N_16820);
nor U22296 (N_22296,N_17419,N_16524);
and U22297 (N_22297,N_17836,N_14832);
or U22298 (N_22298,N_12745,N_13913);
nor U22299 (N_22299,N_16932,N_14474);
xor U22300 (N_22300,N_15331,N_13966);
nor U22301 (N_22301,N_16934,N_16758);
nand U22302 (N_22302,N_14390,N_16251);
and U22303 (N_22303,N_13500,N_13414);
nor U22304 (N_22304,N_17009,N_16890);
xnor U22305 (N_22305,N_17274,N_12165);
nand U22306 (N_22306,N_16912,N_12966);
xnor U22307 (N_22307,N_17136,N_17320);
and U22308 (N_22308,N_16720,N_17909);
or U22309 (N_22309,N_17475,N_17176);
and U22310 (N_22310,N_16656,N_17357);
and U22311 (N_22311,N_17197,N_15820);
or U22312 (N_22312,N_13054,N_14700);
and U22313 (N_22313,N_16591,N_14336);
nand U22314 (N_22314,N_17918,N_14150);
xnor U22315 (N_22315,N_17399,N_15900);
and U22316 (N_22316,N_13054,N_15763);
or U22317 (N_22317,N_14091,N_16701);
or U22318 (N_22318,N_16447,N_12330);
nand U22319 (N_22319,N_12139,N_12634);
or U22320 (N_22320,N_15978,N_14947);
nand U22321 (N_22321,N_14057,N_12665);
nor U22322 (N_22322,N_17652,N_14891);
xnor U22323 (N_22323,N_14431,N_15523);
nor U22324 (N_22324,N_12226,N_12867);
nand U22325 (N_22325,N_16685,N_15890);
and U22326 (N_22326,N_16636,N_16558);
nand U22327 (N_22327,N_13836,N_13360);
or U22328 (N_22328,N_14154,N_16966);
nand U22329 (N_22329,N_16783,N_13293);
nor U22330 (N_22330,N_13229,N_14199);
and U22331 (N_22331,N_15220,N_14387);
nand U22332 (N_22332,N_15395,N_16227);
xnor U22333 (N_22333,N_12864,N_15099);
nor U22334 (N_22334,N_15151,N_12544);
and U22335 (N_22335,N_14294,N_16697);
nor U22336 (N_22336,N_13160,N_13690);
or U22337 (N_22337,N_13616,N_13778);
xnor U22338 (N_22338,N_16783,N_13181);
or U22339 (N_22339,N_16244,N_14016);
xor U22340 (N_22340,N_13791,N_17315);
nor U22341 (N_22341,N_12900,N_17231);
and U22342 (N_22342,N_14559,N_15821);
nand U22343 (N_22343,N_16825,N_14872);
nand U22344 (N_22344,N_13274,N_16777);
nand U22345 (N_22345,N_17659,N_12010);
xor U22346 (N_22346,N_15926,N_14929);
nor U22347 (N_22347,N_15750,N_13317);
or U22348 (N_22348,N_12558,N_12846);
xor U22349 (N_22349,N_13112,N_12274);
nand U22350 (N_22350,N_15924,N_15196);
nor U22351 (N_22351,N_14861,N_15529);
nor U22352 (N_22352,N_12997,N_16755);
xnor U22353 (N_22353,N_12120,N_15899);
and U22354 (N_22354,N_17266,N_12603);
xor U22355 (N_22355,N_14195,N_16717);
or U22356 (N_22356,N_15538,N_13199);
and U22357 (N_22357,N_12960,N_13257);
or U22358 (N_22358,N_17891,N_15711);
nor U22359 (N_22359,N_15808,N_15908);
xnor U22360 (N_22360,N_13733,N_15209);
xnor U22361 (N_22361,N_17884,N_16168);
xor U22362 (N_22362,N_13267,N_15304);
xor U22363 (N_22363,N_17613,N_12460);
xnor U22364 (N_22364,N_14754,N_15291);
and U22365 (N_22365,N_15765,N_15972);
and U22366 (N_22366,N_12034,N_16626);
nor U22367 (N_22367,N_14238,N_15248);
nand U22368 (N_22368,N_13338,N_12301);
xnor U22369 (N_22369,N_13703,N_15710);
nor U22370 (N_22370,N_13796,N_17972);
xor U22371 (N_22371,N_14844,N_14265);
and U22372 (N_22372,N_15920,N_14394);
nor U22373 (N_22373,N_14604,N_12870);
nand U22374 (N_22374,N_13387,N_16187);
nor U22375 (N_22375,N_15853,N_13476);
xnor U22376 (N_22376,N_16177,N_16130);
nand U22377 (N_22377,N_16140,N_16677);
xnor U22378 (N_22378,N_17632,N_14228);
and U22379 (N_22379,N_17319,N_17284);
or U22380 (N_22380,N_14666,N_17774);
or U22381 (N_22381,N_13869,N_12170);
xor U22382 (N_22382,N_12956,N_15260);
nand U22383 (N_22383,N_12260,N_15689);
and U22384 (N_22384,N_15263,N_16010);
or U22385 (N_22385,N_17888,N_14488);
nor U22386 (N_22386,N_17712,N_14475);
and U22387 (N_22387,N_12509,N_16538);
and U22388 (N_22388,N_15032,N_12499);
and U22389 (N_22389,N_13694,N_17529);
xnor U22390 (N_22390,N_15517,N_14979);
nor U22391 (N_22391,N_16829,N_12717);
xnor U22392 (N_22392,N_17935,N_17622);
xor U22393 (N_22393,N_15392,N_14557);
or U22394 (N_22394,N_15531,N_14541);
nor U22395 (N_22395,N_17769,N_14503);
nor U22396 (N_22396,N_12699,N_12719);
xor U22397 (N_22397,N_17200,N_17989);
nor U22398 (N_22398,N_15801,N_15925);
xor U22399 (N_22399,N_13254,N_14052);
nor U22400 (N_22400,N_12999,N_13379);
and U22401 (N_22401,N_15030,N_15182);
nor U22402 (N_22402,N_12903,N_12481);
or U22403 (N_22403,N_13705,N_13992);
nand U22404 (N_22404,N_17738,N_16329);
or U22405 (N_22405,N_14577,N_14920);
xnor U22406 (N_22406,N_13075,N_12350);
or U22407 (N_22407,N_15053,N_14498);
nand U22408 (N_22408,N_12111,N_12907);
or U22409 (N_22409,N_12449,N_13646);
or U22410 (N_22410,N_15040,N_12859);
or U22411 (N_22411,N_14936,N_14855);
and U22412 (N_22412,N_14030,N_16250);
xnor U22413 (N_22413,N_14446,N_13363);
or U22414 (N_22414,N_12160,N_14665);
xnor U22415 (N_22415,N_16853,N_17070);
xor U22416 (N_22416,N_12770,N_13185);
or U22417 (N_22417,N_13617,N_15672);
nor U22418 (N_22418,N_16035,N_17029);
or U22419 (N_22419,N_15301,N_17185);
and U22420 (N_22420,N_16314,N_14350);
and U22421 (N_22421,N_15566,N_15801);
xnor U22422 (N_22422,N_12056,N_12631);
or U22423 (N_22423,N_17325,N_14458);
or U22424 (N_22424,N_14750,N_16060);
nand U22425 (N_22425,N_12173,N_13634);
nand U22426 (N_22426,N_16478,N_12138);
or U22427 (N_22427,N_17317,N_12585);
and U22428 (N_22428,N_13048,N_13203);
nand U22429 (N_22429,N_15786,N_15085);
nor U22430 (N_22430,N_16509,N_15247);
or U22431 (N_22431,N_15544,N_14905);
nand U22432 (N_22432,N_14478,N_16371);
or U22433 (N_22433,N_16316,N_14180);
xor U22434 (N_22434,N_17534,N_14644);
xnor U22435 (N_22435,N_16120,N_14435);
xnor U22436 (N_22436,N_17318,N_15193);
xor U22437 (N_22437,N_16464,N_16085);
nor U22438 (N_22438,N_15754,N_16733);
nand U22439 (N_22439,N_17515,N_17533);
and U22440 (N_22440,N_15538,N_12062);
nor U22441 (N_22441,N_17808,N_14871);
nor U22442 (N_22442,N_15642,N_13373);
or U22443 (N_22443,N_14873,N_13132);
nand U22444 (N_22444,N_17443,N_13159);
or U22445 (N_22445,N_16405,N_16570);
nand U22446 (N_22446,N_12784,N_15363);
nand U22447 (N_22447,N_12283,N_15032);
nand U22448 (N_22448,N_14678,N_16738);
or U22449 (N_22449,N_16127,N_17329);
or U22450 (N_22450,N_17325,N_13993);
and U22451 (N_22451,N_15051,N_12881);
nor U22452 (N_22452,N_15174,N_15158);
xor U22453 (N_22453,N_16972,N_16356);
xnor U22454 (N_22454,N_16306,N_13706);
nand U22455 (N_22455,N_13301,N_15605);
xnor U22456 (N_22456,N_14685,N_17537);
nand U22457 (N_22457,N_15563,N_12283);
or U22458 (N_22458,N_15495,N_12820);
or U22459 (N_22459,N_13394,N_17125);
nor U22460 (N_22460,N_14910,N_17653);
nand U22461 (N_22461,N_16814,N_16790);
nand U22462 (N_22462,N_15763,N_17298);
nor U22463 (N_22463,N_17582,N_17111);
nor U22464 (N_22464,N_14495,N_13904);
nor U22465 (N_22465,N_16091,N_16847);
nor U22466 (N_22466,N_14102,N_17674);
or U22467 (N_22467,N_17497,N_12249);
xor U22468 (N_22468,N_17972,N_17010);
nor U22469 (N_22469,N_14424,N_17715);
or U22470 (N_22470,N_13537,N_17848);
xor U22471 (N_22471,N_13599,N_16879);
or U22472 (N_22472,N_12894,N_12656);
nand U22473 (N_22473,N_16144,N_13012);
or U22474 (N_22474,N_16933,N_15089);
xor U22475 (N_22475,N_13286,N_14449);
xor U22476 (N_22476,N_16373,N_13102);
and U22477 (N_22477,N_15636,N_17184);
nand U22478 (N_22478,N_12663,N_15140);
nand U22479 (N_22479,N_17725,N_16334);
or U22480 (N_22480,N_17318,N_17219);
nor U22481 (N_22481,N_15819,N_14965);
xor U22482 (N_22482,N_16966,N_12935);
nand U22483 (N_22483,N_16016,N_12835);
nand U22484 (N_22484,N_13789,N_15112);
nor U22485 (N_22485,N_14378,N_12162);
xor U22486 (N_22486,N_15505,N_16487);
or U22487 (N_22487,N_12544,N_12669);
or U22488 (N_22488,N_16453,N_12708);
and U22489 (N_22489,N_17427,N_14518);
and U22490 (N_22490,N_15639,N_15333);
nand U22491 (N_22491,N_17540,N_15338);
nor U22492 (N_22492,N_12110,N_12361);
and U22493 (N_22493,N_14038,N_12912);
xor U22494 (N_22494,N_17696,N_13988);
or U22495 (N_22495,N_13966,N_12336);
and U22496 (N_22496,N_17340,N_15619);
nand U22497 (N_22497,N_16350,N_13088);
nand U22498 (N_22498,N_15937,N_15011);
or U22499 (N_22499,N_17099,N_17049);
xor U22500 (N_22500,N_16989,N_16614);
nand U22501 (N_22501,N_16105,N_17790);
and U22502 (N_22502,N_15697,N_13666);
nor U22503 (N_22503,N_15709,N_12247);
nor U22504 (N_22504,N_15514,N_13869);
or U22505 (N_22505,N_17560,N_17202);
xor U22506 (N_22506,N_14246,N_16567);
nor U22507 (N_22507,N_15498,N_14118);
or U22508 (N_22508,N_14797,N_16701);
xor U22509 (N_22509,N_15865,N_14533);
xor U22510 (N_22510,N_16052,N_17105);
or U22511 (N_22511,N_15802,N_17688);
nor U22512 (N_22512,N_13828,N_17099);
or U22513 (N_22513,N_16099,N_16052);
or U22514 (N_22514,N_17071,N_17055);
nor U22515 (N_22515,N_13643,N_13653);
xnor U22516 (N_22516,N_17834,N_16113);
and U22517 (N_22517,N_17261,N_12938);
nand U22518 (N_22518,N_17461,N_16901);
nor U22519 (N_22519,N_15965,N_13166);
xnor U22520 (N_22520,N_16169,N_17708);
nor U22521 (N_22521,N_16437,N_15024);
and U22522 (N_22522,N_13077,N_12553);
nand U22523 (N_22523,N_17386,N_16947);
nor U22524 (N_22524,N_14440,N_14794);
or U22525 (N_22525,N_12567,N_17218);
nor U22526 (N_22526,N_13105,N_14350);
nand U22527 (N_22527,N_17720,N_14097);
xnor U22528 (N_22528,N_12561,N_15274);
and U22529 (N_22529,N_15548,N_14587);
and U22530 (N_22530,N_14393,N_17184);
and U22531 (N_22531,N_16704,N_17846);
and U22532 (N_22532,N_16606,N_16617);
or U22533 (N_22533,N_15393,N_14468);
and U22534 (N_22534,N_13020,N_16696);
nand U22535 (N_22535,N_12604,N_15423);
nand U22536 (N_22536,N_16610,N_13131);
and U22537 (N_22537,N_12229,N_14784);
nand U22538 (N_22538,N_15001,N_14511);
and U22539 (N_22539,N_14342,N_16187);
or U22540 (N_22540,N_13773,N_15409);
nand U22541 (N_22541,N_16762,N_16454);
nand U22542 (N_22542,N_17769,N_15597);
nor U22543 (N_22543,N_15523,N_13813);
nor U22544 (N_22544,N_17120,N_17565);
nor U22545 (N_22545,N_17599,N_15228);
nor U22546 (N_22546,N_17981,N_15181);
xor U22547 (N_22547,N_13664,N_16575);
nand U22548 (N_22548,N_16151,N_17064);
nor U22549 (N_22549,N_14228,N_13262);
nor U22550 (N_22550,N_14529,N_16795);
and U22551 (N_22551,N_13687,N_13207);
nor U22552 (N_22552,N_13471,N_17574);
xor U22553 (N_22553,N_14883,N_14179);
or U22554 (N_22554,N_12957,N_15270);
nor U22555 (N_22555,N_12655,N_16651);
nor U22556 (N_22556,N_14513,N_13329);
xor U22557 (N_22557,N_12956,N_15590);
or U22558 (N_22558,N_12085,N_14198);
and U22559 (N_22559,N_16199,N_17226);
nor U22560 (N_22560,N_16780,N_13183);
nor U22561 (N_22561,N_16166,N_17558);
or U22562 (N_22562,N_12199,N_17688);
xnor U22563 (N_22563,N_13528,N_12555);
nand U22564 (N_22564,N_16977,N_14129);
or U22565 (N_22565,N_12077,N_12000);
nand U22566 (N_22566,N_12401,N_13795);
xnor U22567 (N_22567,N_12370,N_13048);
and U22568 (N_22568,N_16342,N_16642);
nor U22569 (N_22569,N_12126,N_17200);
or U22570 (N_22570,N_13358,N_12534);
and U22571 (N_22571,N_16369,N_16777);
nand U22572 (N_22572,N_15752,N_16487);
nor U22573 (N_22573,N_14178,N_16194);
or U22574 (N_22574,N_12757,N_17087);
or U22575 (N_22575,N_13061,N_13648);
and U22576 (N_22576,N_15941,N_12166);
nand U22577 (N_22577,N_12961,N_16850);
and U22578 (N_22578,N_14123,N_13148);
nor U22579 (N_22579,N_15240,N_14517);
xor U22580 (N_22580,N_13757,N_17208);
xor U22581 (N_22581,N_15265,N_16647);
or U22582 (N_22582,N_17309,N_16375);
xnor U22583 (N_22583,N_15455,N_14850);
or U22584 (N_22584,N_16877,N_14239);
or U22585 (N_22585,N_16069,N_15190);
xor U22586 (N_22586,N_16980,N_12248);
xnor U22587 (N_22587,N_13984,N_13108);
or U22588 (N_22588,N_15460,N_14522);
nand U22589 (N_22589,N_17734,N_15754);
nor U22590 (N_22590,N_17578,N_13700);
nor U22591 (N_22591,N_16090,N_13335);
xor U22592 (N_22592,N_15269,N_15437);
or U22593 (N_22593,N_15117,N_14543);
nand U22594 (N_22594,N_15965,N_16140);
xnor U22595 (N_22595,N_13774,N_14854);
nor U22596 (N_22596,N_12370,N_15669);
nor U22597 (N_22597,N_14241,N_16208);
nor U22598 (N_22598,N_17896,N_13521);
nand U22599 (N_22599,N_12406,N_16980);
nand U22600 (N_22600,N_14744,N_17255);
or U22601 (N_22601,N_12808,N_15597);
or U22602 (N_22602,N_12679,N_14963);
or U22603 (N_22603,N_16371,N_14672);
xnor U22604 (N_22604,N_15079,N_16190);
nand U22605 (N_22605,N_13602,N_12318);
nand U22606 (N_22606,N_17466,N_12750);
nand U22607 (N_22607,N_12370,N_16558);
or U22608 (N_22608,N_13102,N_13973);
nor U22609 (N_22609,N_15769,N_14125);
or U22610 (N_22610,N_16803,N_16760);
nor U22611 (N_22611,N_16996,N_17092);
xnor U22612 (N_22612,N_12656,N_14760);
xor U22613 (N_22613,N_12491,N_16793);
or U22614 (N_22614,N_17160,N_17009);
or U22615 (N_22615,N_13184,N_13475);
nor U22616 (N_22616,N_14755,N_15687);
nand U22617 (N_22617,N_15937,N_15892);
and U22618 (N_22618,N_13304,N_14225);
and U22619 (N_22619,N_15730,N_15312);
or U22620 (N_22620,N_15134,N_13146);
nor U22621 (N_22621,N_17709,N_15566);
or U22622 (N_22622,N_15322,N_13140);
xor U22623 (N_22623,N_14328,N_16470);
and U22624 (N_22624,N_15252,N_17642);
or U22625 (N_22625,N_17008,N_16031);
nor U22626 (N_22626,N_17114,N_12612);
and U22627 (N_22627,N_17932,N_17386);
xnor U22628 (N_22628,N_17885,N_17083);
nand U22629 (N_22629,N_16835,N_16642);
nor U22630 (N_22630,N_14745,N_17047);
nor U22631 (N_22631,N_14797,N_16670);
nand U22632 (N_22632,N_14819,N_12820);
or U22633 (N_22633,N_12593,N_13634);
or U22634 (N_22634,N_12978,N_15916);
nand U22635 (N_22635,N_12629,N_12646);
or U22636 (N_22636,N_14486,N_15675);
and U22637 (N_22637,N_15588,N_13532);
xnor U22638 (N_22638,N_13953,N_13766);
and U22639 (N_22639,N_17250,N_17203);
nand U22640 (N_22640,N_17955,N_16610);
nor U22641 (N_22641,N_12865,N_12821);
or U22642 (N_22642,N_14826,N_16853);
nor U22643 (N_22643,N_12814,N_13178);
nor U22644 (N_22644,N_12004,N_13238);
nand U22645 (N_22645,N_13269,N_16258);
or U22646 (N_22646,N_14642,N_13782);
or U22647 (N_22647,N_13524,N_16937);
nor U22648 (N_22648,N_13072,N_16220);
nand U22649 (N_22649,N_17703,N_12160);
and U22650 (N_22650,N_12142,N_14018);
or U22651 (N_22651,N_16419,N_16113);
or U22652 (N_22652,N_16742,N_17448);
or U22653 (N_22653,N_13928,N_15997);
or U22654 (N_22654,N_13573,N_14734);
nor U22655 (N_22655,N_17279,N_12535);
and U22656 (N_22656,N_14391,N_17798);
or U22657 (N_22657,N_13992,N_14720);
nand U22658 (N_22658,N_17274,N_12320);
nand U22659 (N_22659,N_14964,N_12711);
nor U22660 (N_22660,N_16188,N_16117);
nand U22661 (N_22661,N_15340,N_12398);
nor U22662 (N_22662,N_14740,N_16466);
and U22663 (N_22663,N_13337,N_13365);
and U22664 (N_22664,N_17612,N_14630);
nor U22665 (N_22665,N_16654,N_13481);
nand U22666 (N_22666,N_17961,N_15563);
xnor U22667 (N_22667,N_13828,N_17060);
and U22668 (N_22668,N_15596,N_16782);
nor U22669 (N_22669,N_17246,N_14308);
or U22670 (N_22670,N_16391,N_13351);
nand U22671 (N_22671,N_13753,N_12301);
xor U22672 (N_22672,N_15795,N_12834);
xor U22673 (N_22673,N_15429,N_12215);
nand U22674 (N_22674,N_14990,N_12382);
and U22675 (N_22675,N_13282,N_12663);
nor U22676 (N_22676,N_13058,N_13887);
xnor U22677 (N_22677,N_13057,N_16244);
nor U22678 (N_22678,N_16960,N_13763);
xor U22679 (N_22679,N_17934,N_14349);
xor U22680 (N_22680,N_14628,N_13913);
nor U22681 (N_22681,N_13987,N_12552);
nand U22682 (N_22682,N_16332,N_16392);
xnor U22683 (N_22683,N_14108,N_12089);
nor U22684 (N_22684,N_17802,N_16750);
or U22685 (N_22685,N_17218,N_12140);
and U22686 (N_22686,N_17505,N_15845);
nand U22687 (N_22687,N_16502,N_17089);
and U22688 (N_22688,N_15208,N_16804);
nor U22689 (N_22689,N_16663,N_17687);
or U22690 (N_22690,N_13132,N_14085);
nor U22691 (N_22691,N_15682,N_17988);
nor U22692 (N_22692,N_12481,N_12716);
xor U22693 (N_22693,N_16956,N_14562);
or U22694 (N_22694,N_12420,N_17019);
nand U22695 (N_22695,N_15849,N_15879);
or U22696 (N_22696,N_13478,N_15828);
nor U22697 (N_22697,N_13019,N_15489);
nor U22698 (N_22698,N_16884,N_15776);
and U22699 (N_22699,N_12388,N_12726);
xnor U22700 (N_22700,N_13504,N_13987);
xor U22701 (N_22701,N_14506,N_15531);
xnor U22702 (N_22702,N_16909,N_15661);
nand U22703 (N_22703,N_12162,N_17344);
nand U22704 (N_22704,N_15767,N_17027);
and U22705 (N_22705,N_14018,N_15891);
and U22706 (N_22706,N_12512,N_15005);
xnor U22707 (N_22707,N_16655,N_13665);
xor U22708 (N_22708,N_17525,N_17111);
or U22709 (N_22709,N_13449,N_15433);
and U22710 (N_22710,N_17081,N_12264);
nor U22711 (N_22711,N_12050,N_15367);
or U22712 (N_22712,N_17421,N_16022);
nor U22713 (N_22713,N_17216,N_14016);
and U22714 (N_22714,N_17497,N_14483);
xor U22715 (N_22715,N_16989,N_14990);
nor U22716 (N_22716,N_14188,N_12596);
or U22717 (N_22717,N_16418,N_17419);
xnor U22718 (N_22718,N_17990,N_12268);
nand U22719 (N_22719,N_17656,N_16824);
nor U22720 (N_22720,N_14737,N_13840);
xnor U22721 (N_22721,N_13395,N_15203);
and U22722 (N_22722,N_15321,N_12632);
and U22723 (N_22723,N_16527,N_14729);
or U22724 (N_22724,N_12450,N_14260);
or U22725 (N_22725,N_17489,N_15317);
and U22726 (N_22726,N_17994,N_17233);
xor U22727 (N_22727,N_13593,N_15245);
nand U22728 (N_22728,N_13062,N_13707);
and U22729 (N_22729,N_13925,N_17737);
xnor U22730 (N_22730,N_13527,N_15186);
and U22731 (N_22731,N_14970,N_17504);
nand U22732 (N_22732,N_13435,N_15574);
xnor U22733 (N_22733,N_13271,N_16197);
and U22734 (N_22734,N_12705,N_12161);
xnor U22735 (N_22735,N_12262,N_14365);
xor U22736 (N_22736,N_13014,N_17767);
and U22737 (N_22737,N_16396,N_15262);
nor U22738 (N_22738,N_15250,N_14182);
or U22739 (N_22739,N_12582,N_12389);
nand U22740 (N_22740,N_14162,N_17274);
xor U22741 (N_22741,N_14200,N_14444);
xnor U22742 (N_22742,N_13558,N_12573);
nor U22743 (N_22743,N_12657,N_12096);
and U22744 (N_22744,N_12779,N_15629);
nand U22745 (N_22745,N_16591,N_14568);
nor U22746 (N_22746,N_14756,N_16023);
xor U22747 (N_22747,N_14853,N_12630);
nand U22748 (N_22748,N_14092,N_13686);
and U22749 (N_22749,N_16639,N_17650);
and U22750 (N_22750,N_15723,N_16740);
and U22751 (N_22751,N_14673,N_16880);
xor U22752 (N_22752,N_15569,N_16770);
and U22753 (N_22753,N_12371,N_13600);
nor U22754 (N_22754,N_13780,N_17807);
and U22755 (N_22755,N_12269,N_14336);
nor U22756 (N_22756,N_17168,N_14197);
or U22757 (N_22757,N_14790,N_13234);
nand U22758 (N_22758,N_14989,N_14707);
xor U22759 (N_22759,N_13524,N_16141);
nand U22760 (N_22760,N_13566,N_16459);
and U22761 (N_22761,N_12370,N_15997);
nor U22762 (N_22762,N_16300,N_13675);
xor U22763 (N_22763,N_13231,N_13889);
or U22764 (N_22764,N_16470,N_16954);
nand U22765 (N_22765,N_14450,N_15639);
xor U22766 (N_22766,N_16137,N_15175);
nand U22767 (N_22767,N_13887,N_15285);
nand U22768 (N_22768,N_17151,N_12042);
and U22769 (N_22769,N_14127,N_13024);
and U22770 (N_22770,N_16814,N_16394);
xor U22771 (N_22771,N_13293,N_17818);
nand U22772 (N_22772,N_14318,N_12675);
xnor U22773 (N_22773,N_17394,N_14713);
xor U22774 (N_22774,N_13213,N_12213);
nor U22775 (N_22775,N_13364,N_16147);
xor U22776 (N_22776,N_13297,N_17687);
nor U22777 (N_22777,N_17864,N_16274);
or U22778 (N_22778,N_17955,N_14820);
xnor U22779 (N_22779,N_13091,N_15355);
and U22780 (N_22780,N_16634,N_14233);
nor U22781 (N_22781,N_15889,N_15832);
or U22782 (N_22782,N_16614,N_16538);
nand U22783 (N_22783,N_15365,N_13531);
nand U22784 (N_22784,N_17364,N_16680);
and U22785 (N_22785,N_14747,N_14954);
nand U22786 (N_22786,N_17605,N_17506);
xnor U22787 (N_22787,N_12394,N_14374);
nor U22788 (N_22788,N_12656,N_15969);
nor U22789 (N_22789,N_14612,N_16136);
and U22790 (N_22790,N_15690,N_13261);
nand U22791 (N_22791,N_14588,N_16714);
and U22792 (N_22792,N_17553,N_17815);
nor U22793 (N_22793,N_16980,N_17501);
nand U22794 (N_22794,N_17458,N_16333);
and U22795 (N_22795,N_13701,N_16883);
and U22796 (N_22796,N_15022,N_14552);
nand U22797 (N_22797,N_16444,N_17775);
or U22798 (N_22798,N_12141,N_13620);
and U22799 (N_22799,N_17597,N_15670);
or U22800 (N_22800,N_16596,N_16563);
or U22801 (N_22801,N_14070,N_13014);
and U22802 (N_22802,N_16083,N_12540);
nor U22803 (N_22803,N_13515,N_16891);
nor U22804 (N_22804,N_12428,N_17820);
and U22805 (N_22805,N_13588,N_16545);
and U22806 (N_22806,N_14177,N_13296);
or U22807 (N_22807,N_12212,N_12383);
nor U22808 (N_22808,N_16707,N_12400);
and U22809 (N_22809,N_16096,N_12084);
nor U22810 (N_22810,N_16043,N_13129);
nand U22811 (N_22811,N_16652,N_16323);
nand U22812 (N_22812,N_14365,N_16128);
nand U22813 (N_22813,N_17647,N_14538);
nor U22814 (N_22814,N_16555,N_12325);
nand U22815 (N_22815,N_16949,N_15566);
nor U22816 (N_22816,N_15499,N_12363);
nor U22817 (N_22817,N_12189,N_15286);
or U22818 (N_22818,N_16546,N_15671);
or U22819 (N_22819,N_14855,N_12990);
nand U22820 (N_22820,N_12509,N_12075);
or U22821 (N_22821,N_13539,N_17629);
xnor U22822 (N_22822,N_17643,N_12339);
xor U22823 (N_22823,N_13794,N_15589);
and U22824 (N_22824,N_13052,N_14221);
and U22825 (N_22825,N_16812,N_15520);
nor U22826 (N_22826,N_16438,N_13012);
or U22827 (N_22827,N_16074,N_14751);
and U22828 (N_22828,N_15205,N_17075);
and U22829 (N_22829,N_17358,N_12831);
and U22830 (N_22830,N_13789,N_13258);
nor U22831 (N_22831,N_16927,N_14374);
xnor U22832 (N_22832,N_17812,N_13323);
xor U22833 (N_22833,N_14153,N_12398);
or U22834 (N_22834,N_12910,N_12354);
nor U22835 (N_22835,N_12609,N_16726);
nor U22836 (N_22836,N_13581,N_12044);
nand U22837 (N_22837,N_14665,N_17173);
xnor U22838 (N_22838,N_17891,N_17755);
nor U22839 (N_22839,N_15342,N_16227);
nand U22840 (N_22840,N_15406,N_13009);
nand U22841 (N_22841,N_15022,N_12160);
or U22842 (N_22842,N_16506,N_15035);
nand U22843 (N_22843,N_12946,N_17964);
xnor U22844 (N_22844,N_14141,N_14941);
xor U22845 (N_22845,N_15894,N_16157);
nand U22846 (N_22846,N_13687,N_15845);
xnor U22847 (N_22847,N_14207,N_12835);
or U22848 (N_22848,N_16863,N_16612);
nand U22849 (N_22849,N_15405,N_12456);
xor U22850 (N_22850,N_12179,N_12970);
nor U22851 (N_22851,N_16421,N_15034);
and U22852 (N_22852,N_15909,N_16899);
or U22853 (N_22853,N_17469,N_13553);
nor U22854 (N_22854,N_15048,N_13305);
xor U22855 (N_22855,N_13737,N_17163);
and U22856 (N_22856,N_16389,N_16760);
nand U22857 (N_22857,N_16017,N_16056);
nand U22858 (N_22858,N_12836,N_17952);
nand U22859 (N_22859,N_17872,N_13667);
and U22860 (N_22860,N_13791,N_17917);
nor U22861 (N_22861,N_13437,N_16267);
nor U22862 (N_22862,N_12892,N_12453);
xor U22863 (N_22863,N_16443,N_17427);
or U22864 (N_22864,N_16438,N_17461);
xnor U22865 (N_22865,N_17035,N_14029);
or U22866 (N_22866,N_13398,N_14123);
nand U22867 (N_22867,N_16865,N_17287);
or U22868 (N_22868,N_16720,N_16036);
xnor U22869 (N_22869,N_15081,N_13816);
xor U22870 (N_22870,N_13005,N_16264);
or U22871 (N_22871,N_14902,N_16959);
and U22872 (N_22872,N_13645,N_17047);
nor U22873 (N_22873,N_14310,N_15538);
nand U22874 (N_22874,N_12626,N_14942);
nor U22875 (N_22875,N_13020,N_12308);
nor U22876 (N_22876,N_15622,N_17870);
and U22877 (N_22877,N_17764,N_12419);
and U22878 (N_22878,N_16489,N_13655);
and U22879 (N_22879,N_17658,N_16819);
nor U22880 (N_22880,N_12151,N_17146);
and U22881 (N_22881,N_16156,N_15870);
nor U22882 (N_22882,N_13375,N_17167);
nor U22883 (N_22883,N_16932,N_14917);
xor U22884 (N_22884,N_16029,N_13046);
nor U22885 (N_22885,N_15786,N_12099);
nor U22886 (N_22886,N_12230,N_16549);
and U22887 (N_22887,N_15147,N_14337);
or U22888 (N_22888,N_14542,N_17670);
nor U22889 (N_22889,N_14301,N_15697);
and U22890 (N_22890,N_17156,N_17396);
nor U22891 (N_22891,N_14316,N_15153);
and U22892 (N_22892,N_14489,N_17603);
or U22893 (N_22893,N_16375,N_12413);
xnor U22894 (N_22894,N_16022,N_15069);
and U22895 (N_22895,N_13997,N_15379);
nand U22896 (N_22896,N_13283,N_16950);
nor U22897 (N_22897,N_17325,N_12215);
nand U22898 (N_22898,N_14537,N_14805);
nand U22899 (N_22899,N_15737,N_16127);
or U22900 (N_22900,N_17224,N_17107);
or U22901 (N_22901,N_12466,N_13752);
nand U22902 (N_22902,N_16156,N_14975);
xnor U22903 (N_22903,N_12820,N_15717);
and U22904 (N_22904,N_12302,N_17279);
nor U22905 (N_22905,N_14160,N_16331);
and U22906 (N_22906,N_12135,N_16354);
and U22907 (N_22907,N_14405,N_15648);
xor U22908 (N_22908,N_16750,N_17894);
xnor U22909 (N_22909,N_13288,N_14713);
xnor U22910 (N_22910,N_14261,N_14647);
nor U22911 (N_22911,N_12053,N_13816);
or U22912 (N_22912,N_12847,N_15066);
nand U22913 (N_22913,N_13661,N_15907);
nand U22914 (N_22914,N_13724,N_16369);
or U22915 (N_22915,N_17760,N_15173);
nor U22916 (N_22916,N_17308,N_16845);
or U22917 (N_22917,N_14988,N_13312);
nand U22918 (N_22918,N_17113,N_16317);
xor U22919 (N_22919,N_16654,N_16082);
nor U22920 (N_22920,N_15562,N_15790);
nor U22921 (N_22921,N_14696,N_14524);
and U22922 (N_22922,N_14702,N_13151);
nor U22923 (N_22923,N_16153,N_15515);
xnor U22924 (N_22924,N_15295,N_16506);
or U22925 (N_22925,N_14379,N_13453);
and U22926 (N_22926,N_16349,N_14559);
or U22927 (N_22927,N_12142,N_16450);
nor U22928 (N_22928,N_16774,N_17585);
xnor U22929 (N_22929,N_17030,N_12508);
nand U22930 (N_22930,N_16601,N_16980);
or U22931 (N_22931,N_12073,N_15526);
nor U22932 (N_22932,N_13804,N_13926);
or U22933 (N_22933,N_12559,N_13132);
nand U22934 (N_22934,N_17582,N_17730);
and U22935 (N_22935,N_16400,N_14093);
xor U22936 (N_22936,N_12344,N_15782);
or U22937 (N_22937,N_17601,N_17901);
nand U22938 (N_22938,N_12308,N_12352);
or U22939 (N_22939,N_14021,N_15551);
nand U22940 (N_22940,N_16710,N_14109);
nor U22941 (N_22941,N_13181,N_17746);
nor U22942 (N_22942,N_12460,N_14380);
and U22943 (N_22943,N_12418,N_16917);
or U22944 (N_22944,N_16427,N_12051);
xor U22945 (N_22945,N_16927,N_15802);
and U22946 (N_22946,N_13510,N_17530);
or U22947 (N_22947,N_13910,N_13506);
nand U22948 (N_22948,N_15390,N_16069);
xor U22949 (N_22949,N_12583,N_13979);
nand U22950 (N_22950,N_14612,N_15800);
nand U22951 (N_22951,N_12245,N_17866);
and U22952 (N_22952,N_17638,N_13987);
xor U22953 (N_22953,N_12765,N_17969);
nand U22954 (N_22954,N_14815,N_13053);
and U22955 (N_22955,N_16822,N_15909);
nor U22956 (N_22956,N_14285,N_14576);
nor U22957 (N_22957,N_16418,N_14814);
nand U22958 (N_22958,N_12569,N_17002);
nand U22959 (N_22959,N_16278,N_12408);
or U22960 (N_22960,N_17513,N_12988);
nand U22961 (N_22961,N_13913,N_12184);
and U22962 (N_22962,N_17297,N_15932);
and U22963 (N_22963,N_13556,N_15387);
nor U22964 (N_22964,N_15989,N_15377);
nor U22965 (N_22965,N_15376,N_16365);
and U22966 (N_22966,N_14444,N_17889);
or U22967 (N_22967,N_13393,N_16239);
nor U22968 (N_22968,N_14314,N_15479);
nand U22969 (N_22969,N_13902,N_16671);
nor U22970 (N_22970,N_17476,N_12012);
and U22971 (N_22971,N_15456,N_16492);
nand U22972 (N_22972,N_17865,N_15841);
nor U22973 (N_22973,N_13756,N_17695);
xnor U22974 (N_22974,N_12098,N_15349);
nand U22975 (N_22975,N_15338,N_17367);
nand U22976 (N_22976,N_17618,N_12974);
nor U22977 (N_22977,N_15351,N_16368);
nor U22978 (N_22978,N_16703,N_14506);
or U22979 (N_22979,N_16445,N_14144);
xnor U22980 (N_22980,N_17624,N_14008);
or U22981 (N_22981,N_15061,N_13393);
or U22982 (N_22982,N_14080,N_12886);
or U22983 (N_22983,N_14796,N_17609);
xnor U22984 (N_22984,N_14303,N_14195);
and U22985 (N_22985,N_16906,N_17253);
or U22986 (N_22986,N_14936,N_16150);
and U22987 (N_22987,N_16395,N_17662);
xnor U22988 (N_22988,N_14563,N_15734);
or U22989 (N_22989,N_16237,N_12574);
or U22990 (N_22990,N_17758,N_17631);
or U22991 (N_22991,N_16020,N_13828);
nor U22992 (N_22992,N_13740,N_13007);
xnor U22993 (N_22993,N_14956,N_13812);
xnor U22994 (N_22994,N_16953,N_12473);
xnor U22995 (N_22995,N_15994,N_13854);
nand U22996 (N_22996,N_14832,N_12646);
or U22997 (N_22997,N_16211,N_15360);
and U22998 (N_22998,N_15539,N_13836);
xor U22999 (N_22999,N_15381,N_12676);
or U23000 (N_23000,N_16870,N_16033);
nor U23001 (N_23001,N_17231,N_17260);
nand U23002 (N_23002,N_13147,N_16732);
xor U23003 (N_23003,N_14261,N_15153);
nor U23004 (N_23004,N_15573,N_12990);
or U23005 (N_23005,N_15712,N_13331);
xor U23006 (N_23006,N_14740,N_15920);
or U23007 (N_23007,N_14709,N_15860);
nand U23008 (N_23008,N_13373,N_15759);
or U23009 (N_23009,N_16704,N_12271);
nand U23010 (N_23010,N_17090,N_17607);
or U23011 (N_23011,N_16651,N_15002);
xor U23012 (N_23012,N_14517,N_17721);
xnor U23013 (N_23013,N_14866,N_17133);
nand U23014 (N_23014,N_15624,N_14493);
and U23015 (N_23015,N_13643,N_16539);
and U23016 (N_23016,N_14203,N_16494);
xnor U23017 (N_23017,N_13279,N_14726);
xor U23018 (N_23018,N_15536,N_13582);
nor U23019 (N_23019,N_15647,N_13232);
nor U23020 (N_23020,N_13233,N_16257);
and U23021 (N_23021,N_12901,N_16734);
nor U23022 (N_23022,N_13769,N_17960);
nor U23023 (N_23023,N_12161,N_14140);
nor U23024 (N_23024,N_17849,N_14992);
nand U23025 (N_23025,N_12111,N_14936);
nor U23026 (N_23026,N_15230,N_14477);
and U23027 (N_23027,N_12723,N_17642);
xnor U23028 (N_23028,N_13330,N_12830);
xnor U23029 (N_23029,N_13959,N_15909);
nor U23030 (N_23030,N_16370,N_17315);
xnor U23031 (N_23031,N_15295,N_13402);
and U23032 (N_23032,N_15974,N_12974);
or U23033 (N_23033,N_17326,N_14647);
nor U23034 (N_23034,N_15087,N_17430);
nor U23035 (N_23035,N_13354,N_12146);
nand U23036 (N_23036,N_13287,N_15414);
nor U23037 (N_23037,N_16930,N_16378);
or U23038 (N_23038,N_17984,N_14737);
nor U23039 (N_23039,N_14424,N_12261);
and U23040 (N_23040,N_13440,N_15054);
nor U23041 (N_23041,N_12198,N_17946);
or U23042 (N_23042,N_15219,N_16188);
nand U23043 (N_23043,N_13709,N_16429);
and U23044 (N_23044,N_16807,N_15825);
nand U23045 (N_23045,N_13211,N_17571);
or U23046 (N_23046,N_12816,N_17421);
or U23047 (N_23047,N_15507,N_17136);
nand U23048 (N_23048,N_14275,N_12578);
or U23049 (N_23049,N_12661,N_15125);
or U23050 (N_23050,N_12889,N_15519);
nand U23051 (N_23051,N_12578,N_12357);
or U23052 (N_23052,N_12675,N_17093);
xnor U23053 (N_23053,N_12875,N_16134);
or U23054 (N_23054,N_14088,N_13684);
or U23055 (N_23055,N_12155,N_17145);
or U23056 (N_23056,N_15870,N_17851);
nand U23057 (N_23057,N_13391,N_14940);
xnor U23058 (N_23058,N_17171,N_14232);
xnor U23059 (N_23059,N_12867,N_15107);
and U23060 (N_23060,N_14208,N_13225);
nand U23061 (N_23061,N_12738,N_12768);
nand U23062 (N_23062,N_14576,N_17576);
and U23063 (N_23063,N_17258,N_12361);
nand U23064 (N_23064,N_14739,N_14826);
nand U23065 (N_23065,N_15592,N_16662);
xnor U23066 (N_23066,N_15534,N_12100);
or U23067 (N_23067,N_17046,N_13723);
nand U23068 (N_23068,N_12137,N_17505);
and U23069 (N_23069,N_12054,N_14073);
xor U23070 (N_23070,N_12215,N_17017);
nand U23071 (N_23071,N_14787,N_17232);
xnor U23072 (N_23072,N_16339,N_12401);
and U23073 (N_23073,N_13447,N_14491);
xnor U23074 (N_23074,N_17772,N_14327);
nor U23075 (N_23075,N_14215,N_16944);
nand U23076 (N_23076,N_13951,N_17913);
xnor U23077 (N_23077,N_13299,N_16468);
nand U23078 (N_23078,N_15040,N_15414);
xor U23079 (N_23079,N_15464,N_14727);
or U23080 (N_23080,N_16779,N_14203);
and U23081 (N_23081,N_15987,N_17545);
or U23082 (N_23082,N_12135,N_13313);
and U23083 (N_23083,N_14058,N_12588);
or U23084 (N_23084,N_17480,N_16655);
xor U23085 (N_23085,N_16121,N_17060);
nand U23086 (N_23086,N_14867,N_15789);
and U23087 (N_23087,N_12403,N_13257);
and U23088 (N_23088,N_17601,N_13498);
xor U23089 (N_23089,N_17437,N_14877);
or U23090 (N_23090,N_17679,N_14783);
xor U23091 (N_23091,N_14156,N_13915);
or U23092 (N_23092,N_17706,N_16490);
or U23093 (N_23093,N_17749,N_17763);
nand U23094 (N_23094,N_12567,N_17988);
nor U23095 (N_23095,N_13984,N_12530);
xor U23096 (N_23096,N_14430,N_16937);
nor U23097 (N_23097,N_14953,N_14358);
nor U23098 (N_23098,N_16624,N_13642);
and U23099 (N_23099,N_13297,N_14587);
nor U23100 (N_23100,N_16362,N_17608);
or U23101 (N_23101,N_16698,N_13217);
nand U23102 (N_23102,N_14549,N_15950);
xor U23103 (N_23103,N_13158,N_13389);
xnor U23104 (N_23104,N_13271,N_13064);
nand U23105 (N_23105,N_14737,N_12893);
xor U23106 (N_23106,N_16316,N_12988);
and U23107 (N_23107,N_12568,N_15366);
nand U23108 (N_23108,N_17642,N_14289);
or U23109 (N_23109,N_13648,N_12685);
nand U23110 (N_23110,N_16369,N_15739);
and U23111 (N_23111,N_16103,N_15292);
and U23112 (N_23112,N_14593,N_14870);
nand U23113 (N_23113,N_16415,N_16515);
nor U23114 (N_23114,N_16097,N_13597);
nor U23115 (N_23115,N_17613,N_13085);
and U23116 (N_23116,N_12774,N_15962);
and U23117 (N_23117,N_12636,N_12929);
or U23118 (N_23118,N_17894,N_12002);
xnor U23119 (N_23119,N_13759,N_14547);
and U23120 (N_23120,N_14492,N_13283);
nor U23121 (N_23121,N_17599,N_12049);
xnor U23122 (N_23122,N_12855,N_13106);
or U23123 (N_23123,N_16122,N_14516);
xor U23124 (N_23124,N_13204,N_12067);
nor U23125 (N_23125,N_12065,N_16883);
and U23126 (N_23126,N_17581,N_15754);
and U23127 (N_23127,N_15550,N_14665);
or U23128 (N_23128,N_16067,N_12768);
nand U23129 (N_23129,N_13644,N_14854);
nor U23130 (N_23130,N_15732,N_16553);
nand U23131 (N_23131,N_14597,N_17016);
or U23132 (N_23132,N_17484,N_16011);
nand U23133 (N_23133,N_16826,N_14701);
nand U23134 (N_23134,N_14881,N_13331);
and U23135 (N_23135,N_12430,N_15453);
and U23136 (N_23136,N_13032,N_12945);
nor U23137 (N_23137,N_12013,N_16761);
nor U23138 (N_23138,N_15036,N_17739);
xnor U23139 (N_23139,N_15579,N_13056);
nor U23140 (N_23140,N_14237,N_15095);
nand U23141 (N_23141,N_16330,N_12580);
nand U23142 (N_23142,N_15272,N_12547);
nor U23143 (N_23143,N_13043,N_13073);
nor U23144 (N_23144,N_17980,N_16557);
nor U23145 (N_23145,N_13341,N_16584);
nand U23146 (N_23146,N_14253,N_16716);
xnor U23147 (N_23147,N_13162,N_15479);
nor U23148 (N_23148,N_13114,N_14674);
or U23149 (N_23149,N_15029,N_12922);
nor U23150 (N_23150,N_14033,N_12928);
nand U23151 (N_23151,N_12179,N_14279);
xor U23152 (N_23152,N_15208,N_14287);
nor U23153 (N_23153,N_15526,N_13481);
or U23154 (N_23154,N_16660,N_16037);
or U23155 (N_23155,N_14381,N_13162);
xnor U23156 (N_23156,N_15123,N_17854);
or U23157 (N_23157,N_13078,N_15280);
xor U23158 (N_23158,N_12192,N_15749);
or U23159 (N_23159,N_15674,N_16569);
xor U23160 (N_23160,N_12667,N_17533);
and U23161 (N_23161,N_12706,N_15186);
xor U23162 (N_23162,N_13506,N_17874);
xor U23163 (N_23163,N_16095,N_14083);
nor U23164 (N_23164,N_15995,N_17989);
and U23165 (N_23165,N_16831,N_14745);
and U23166 (N_23166,N_15196,N_14209);
and U23167 (N_23167,N_13068,N_15046);
xor U23168 (N_23168,N_15141,N_14301);
and U23169 (N_23169,N_14810,N_15787);
xor U23170 (N_23170,N_15207,N_13536);
nand U23171 (N_23171,N_16747,N_14074);
nor U23172 (N_23172,N_17898,N_17299);
and U23173 (N_23173,N_12617,N_14174);
xor U23174 (N_23174,N_17454,N_15487);
or U23175 (N_23175,N_13363,N_12126);
nand U23176 (N_23176,N_17157,N_14656);
nand U23177 (N_23177,N_14527,N_13183);
xor U23178 (N_23178,N_17016,N_15019);
and U23179 (N_23179,N_17202,N_13763);
or U23180 (N_23180,N_15386,N_14933);
and U23181 (N_23181,N_14703,N_12131);
xor U23182 (N_23182,N_15836,N_14222);
and U23183 (N_23183,N_13966,N_15961);
nor U23184 (N_23184,N_15659,N_13222);
nor U23185 (N_23185,N_13520,N_16151);
or U23186 (N_23186,N_14907,N_14847);
or U23187 (N_23187,N_17962,N_16307);
xnor U23188 (N_23188,N_13876,N_17510);
or U23189 (N_23189,N_16337,N_17233);
and U23190 (N_23190,N_14845,N_15331);
nor U23191 (N_23191,N_16119,N_12987);
nor U23192 (N_23192,N_17867,N_16422);
xor U23193 (N_23193,N_17804,N_15650);
xor U23194 (N_23194,N_16826,N_16299);
nand U23195 (N_23195,N_16755,N_15421);
and U23196 (N_23196,N_12015,N_14760);
nand U23197 (N_23197,N_15596,N_16239);
nand U23198 (N_23198,N_15445,N_12838);
and U23199 (N_23199,N_14974,N_16206);
or U23200 (N_23200,N_17155,N_12248);
and U23201 (N_23201,N_14459,N_15286);
xor U23202 (N_23202,N_13834,N_16506);
nor U23203 (N_23203,N_16953,N_14804);
and U23204 (N_23204,N_13997,N_17367);
or U23205 (N_23205,N_16127,N_15351);
and U23206 (N_23206,N_13075,N_14710);
or U23207 (N_23207,N_16789,N_17974);
or U23208 (N_23208,N_14994,N_12529);
nor U23209 (N_23209,N_13252,N_13813);
nor U23210 (N_23210,N_13040,N_13764);
nand U23211 (N_23211,N_16555,N_14546);
and U23212 (N_23212,N_16828,N_14072);
or U23213 (N_23213,N_13061,N_14351);
and U23214 (N_23214,N_12394,N_13032);
or U23215 (N_23215,N_15530,N_15839);
nor U23216 (N_23216,N_14064,N_15898);
nand U23217 (N_23217,N_14309,N_16392);
nand U23218 (N_23218,N_12661,N_15081);
and U23219 (N_23219,N_12614,N_14230);
nor U23220 (N_23220,N_16402,N_15941);
or U23221 (N_23221,N_13184,N_12187);
or U23222 (N_23222,N_14253,N_14101);
nor U23223 (N_23223,N_13586,N_16501);
or U23224 (N_23224,N_16770,N_15018);
nand U23225 (N_23225,N_16991,N_16023);
nor U23226 (N_23226,N_14665,N_13391);
xor U23227 (N_23227,N_14798,N_16962);
and U23228 (N_23228,N_15824,N_15693);
nand U23229 (N_23229,N_15762,N_14643);
nand U23230 (N_23230,N_14857,N_16587);
and U23231 (N_23231,N_17244,N_13272);
and U23232 (N_23232,N_16240,N_17101);
or U23233 (N_23233,N_16294,N_16680);
xnor U23234 (N_23234,N_15482,N_12461);
xnor U23235 (N_23235,N_16932,N_15243);
nand U23236 (N_23236,N_17173,N_12948);
nand U23237 (N_23237,N_16021,N_14764);
xor U23238 (N_23238,N_15890,N_15844);
or U23239 (N_23239,N_16438,N_16144);
and U23240 (N_23240,N_17414,N_13069);
nand U23241 (N_23241,N_12319,N_17754);
nand U23242 (N_23242,N_16674,N_16275);
xor U23243 (N_23243,N_17997,N_14010);
nor U23244 (N_23244,N_15565,N_17911);
or U23245 (N_23245,N_17627,N_14020);
and U23246 (N_23246,N_13718,N_12930);
nor U23247 (N_23247,N_12292,N_15903);
nand U23248 (N_23248,N_13254,N_12100);
and U23249 (N_23249,N_14768,N_12569);
nand U23250 (N_23250,N_15989,N_13375);
nor U23251 (N_23251,N_16929,N_15769);
xnor U23252 (N_23252,N_13643,N_16016);
or U23253 (N_23253,N_17543,N_14078);
nand U23254 (N_23254,N_13484,N_17513);
xnor U23255 (N_23255,N_14104,N_13932);
nor U23256 (N_23256,N_12252,N_14270);
nand U23257 (N_23257,N_12023,N_13991);
nor U23258 (N_23258,N_14919,N_16192);
nor U23259 (N_23259,N_15427,N_13876);
nand U23260 (N_23260,N_14470,N_13504);
or U23261 (N_23261,N_17780,N_15185);
nor U23262 (N_23262,N_13147,N_13813);
nand U23263 (N_23263,N_13506,N_14815);
or U23264 (N_23264,N_14215,N_14198);
nor U23265 (N_23265,N_16643,N_17033);
or U23266 (N_23266,N_14818,N_12814);
nand U23267 (N_23267,N_12973,N_15962);
xnor U23268 (N_23268,N_16394,N_13845);
xor U23269 (N_23269,N_15756,N_14571);
and U23270 (N_23270,N_14664,N_16786);
or U23271 (N_23271,N_17474,N_13610);
nor U23272 (N_23272,N_15781,N_16037);
and U23273 (N_23273,N_17378,N_14407);
xnor U23274 (N_23274,N_12264,N_15075);
xor U23275 (N_23275,N_14856,N_15394);
nor U23276 (N_23276,N_17991,N_14894);
xnor U23277 (N_23277,N_16904,N_16897);
nand U23278 (N_23278,N_15455,N_15356);
or U23279 (N_23279,N_17806,N_14619);
xnor U23280 (N_23280,N_13345,N_16585);
or U23281 (N_23281,N_13959,N_13302);
xor U23282 (N_23282,N_12804,N_17002);
nor U23283 (N_23283,N_15182,N_16982);
xnor U23284 (N_23284,N_14423,N_14481);
and U23285 (N_23285,N_13963,N_14128);
or U23286 (N_23286,N_12040,N_12234);
or U23287 (N_23287,N_16100,N_12098);
and U23288 (N_23288,N_17709,N_16688);
xor U23289 (N_23289,N_16726,N_15898);
nor U23290 (N_23290,N_14280,N_16011);
and U23291 (N_23291,N_14072,N_13201);
or U23292 (N_23292,N_17936,N_16484);
nand U23293 (N_23293,N_14309,N_13383);
xor U23294 (N_23294,N_12543,N_13541);
and U23295 (N_23295,N_12483,N_14923);
or U23296 (N_23296,N_12298,N_17248);
xnor U23297 (N_23297,N_16131,N_15266);
nor U23298 (N_23298,N_16497,N_15626);
xnor U23299 (N_23299,N_17873,N_14087);
xnor U23300 (N_23300,N_15708,N_13198);
nor U23301 (N_23301,N_16922,N_17360);
and U23302 (N_23302,N_16321,N_13391);
nand U23303 (N_23303,N_14875,N_16671);
nand U23304 (N_23304,N_17807,N_15047);
or U23305 (N_23305,N_14601,N_16851);
or U23306 (N_23306,N_13185,N_15383);
or U23307 (N_23307,N_12467,N_14068);
or U23308 (N_23308,N_17398,N_16824);
xor U23309 (N_23309,N_14103,N_17935);
xor U23310 (N_23310,N_12150,N_16054);
nand U23311 (N_23311,N_15510,N_14716);
xor U23312 (N_23312,N_13422,N_15976);
nor U23313 (N_23313,N_17993,N_15272);
xnor U23314 (N_23314,N_13551,N_14995);
nor U23315 (N_23315,N_15192,N_13968);
nand U23316 (N_23316,N_14162,N_14988);
nor U23317 (N_23317,N_13308,N_17474);
xnor U23318 (N_23318,N_13350,N_12539);
xor U23319 (N_23319,N_15382,N_16933);
nand U23320 (N_23320,N_13601,N_16209);
and U23321 (N_23321,N_12657,N_15830);
xnor U23322 (N_23322,N_15585,N_17606);
xor U23323 (N_23323,N_12396,N_16661);
or U23324 (N_23324,N_14317,N_16232);
and U23325 (N_23325,N_13061,N_12458);
xor U23326 (N_23326,N_15565,N_14541);
nor U23327 (N_23327,N_15630,N_13020);
nand U23328 (N_23328,N_12939,N_17574);
or U23329 (N_23329,N_14457,N_16437);
nand U23330 (N_23330,N_12358,N_17460);
nand U23331 (N_23331,N_12280,N_15479);
nor U23332 (N_23332,N_17347,N_15444);
and U23333 (N_23333,N_12967,N_16413);
and U23334 (N_23334,N_16452,N_13854);
xnor U23335 (N_23335,N_15083,N_14942);
nand U23336 (N_23336,N_13116,N_12029);
or U23337 (N_23337,N_14859,N_16276);
and U23338 (N_23338,N_12273,N_16999);
and U23339 (N_23339,N_15843,N_12118);
nor U23340 (N_23340,N_17813,N_14931);
xor U23341 (N_23341,N_16974,N_17819);
and U23342 (N_23342,N_15630,N_17022);
nor U23343 (N_23343,N_17859,N_16446);
nor U23344 (N_23344,N_17196,N_16676);
nor U23345 (N_23345,N_16495,N_12221);
nand U23346 (N_23346,N_13535,N_13155);
nor U23347 (N_23347,N_14069,N_14043);
nand U23348 (N_23348,N_14270,N_14904);
and U23349 (N_23349,N_17838,N_13973);
nor U23350 (N_23350,N_15194,N_17261);
or U23351 (N_23351,N_14809,N_13841);
xor U23352 (N_23352,N_16154,N_14527);
nand U23353 (N_23353,N_14070,N_17452);
nor U23354 (N_23354,N_17166,N_16433);
nand U23355 (N_23355,N_12766,N_15176);
and U23356 (N_23356,N_13433,N_15993);
xnor U23357 (N_23357,N_13447,N_16129);
nor U23358 (N_23358,N_15857,N_12553);
or U23359 (N_23359,N_17049,N_13311);
xnor U23360 (N_23360,N_13462,N_14926);
or U23361 (N_23361,N_16862,N_12732);
or U23362 (N_23362,N_12909,N_14306);
nand U23363 (N_23363,N_16574,N_14890);
nor U23364 (N_23364,N_17734,N_13583);
nor U23365 (N_23365,N_14274,N_12247);
nand U23366 (N_23366,N_17511,N_16761);
xnor U23367 (N_23367,N_15932,N_16497);
nor U23368 (N_23368,N_17603,N_12874);
xnor U23369 (N_23369,N_13455,N_16064);
and U23370 (N_23370,N_14689,N_17148);
xnor U23371 (N_23371,N_15036,N_15050);
and U23372 (N_23372,N_15264,N_13375);
nand U23373 (N_23373,N_12473,N_13554);
or U23374 (N_23374,N_17067,N_17495);
or U23375 (N_23375,N_13757,N_15108);
xor U23376 (N_23376,N_13597,N_15667);
and U23377 (N_23377,N_15394,N_17677);
nor U23378 (N_23378,N_17863,N_13108);
and U23379 (N_23379,N_15324,N_16484);
nor U23380 (N_23380,N_12401,N_14608);
nand U23381 (N_23381,N_13492,N_13662);
xnor U23382 (N_23382,N_12643,N_17195);
and U23383 (N_23383,N_16751,N_17219);
or U23384 (N_23384,N_14289,N_12645);
nor U23385 (N_23385,N_15473,N_15288);
nand U23386 (N_23386,N_14754,N_15944);
or U23387 (N_23387,N_13177,N_12937);
nand U23388 (N_23388,N_17778,N_17091);
xnor U23389 (N_23389,N_14309,N_16639);
xnor U23390 (N_23390,N_13996,N_12124);
nor U23391 (N_23391,N_14494,N_13936);
or U23392 (N_23392,N_17610,N_12682);
or U23393 (N_23393,N_15145,N_16413);
xnor U23394 (N_23394,N_15817,N_17742);
nand U23395 (N_23395,N_12427,N_15457);
nand U23396 (N_23396,N_15800,N_15773);
or U23397 (N_23397,N_14304,N_14345);
or U23398 (N_23398,N_17653,N_12295);
and U23399 (N_23399,N_15431,N_16911);
nor U23400 (N_23400,N_12462,N_16612);
nor U23401 (N_23401,N_12782,N_14720);
xnor U23402 (N_23402,N_14088,N_15599);
xor U23403 (N_23403,N_13442,N_15116);
or U23404 (N_23404,N_12198,N_17456);
nand U23405 (N_23405,N_13725,N_14544);
or U23406 (N_23406,N_13971,N_15556);
xnor U23407 (N_23407,N_17195,N_12566);
nor U23408 (N_23408,N_16698,N_14053);
and U23409 (N_23409,N_16454,N_13236);
nor U23410 (N_23410,N_12582,N_13903);
nor U23411 (N_23411,N_12607,N_16016);
nor U23412 (N_23412,N_14377,N_14495);
xnor U23413 (N_23413,N_14466,N_17174);
xor U23414 (N_23414,N_15072,N_17289);
nand U23415 (N_23415,N_16352,N_15201);
nand U23416 (N_23416,N_14729,N_14711);
or U23417 (N_23417,N_15399,N_17683);
or U23418 (N_23418,N_15349,N_16479);
or U23419 (N_23419,N_13152,N_17224);
and U23420 (N_23420,N_16701,N_16576);
nor U23421 (N_23421,N_17880,N_13880);
nor U23422 (N_23422,N_17696,N_14370);
nor U23423 (N_23423,N_16719,N_12547);
or U23424 (N_23424,N_17992,N_14584);
nand U23425 (N_23425,N_15522,N_17259);
or U23426 (N_23426,N_14747,N_14528);
nand U23427 (N_23427,N_12328,N_16677);
xnor U23428 (N_23428,N_13027,N_15132);
and U23429 (N_23429,N_13638,N_14873);
or U23430 (N_23430,N_14212,N_14677);
nor U23431 (N_23431,N_14160,N_13257);
nor U23432 (N_23432,N_12558,N_14696);
nand U23433 (N_23433,N_15621,N_14888);
xor U23434 (N_23434,N_13828,N_13943);
nand U23435 (N_23435,N_17695,N_12473);
xor U23436 (N_23436,N_12957,N_16730);
and U23437 (N_23437,N_13608,N_15377);
nand U23438 (N_23438,N_12629,N_13410);
or U23439 (N_23439,N_17246,N_17627);
xor U23440 (N_23440,N_15980,N_16970);
nand U23441 (N_23441,N_14117,N_14297);
xor U23442 (N_23442,N_12971,N_14407);
and U23443 (N_23443,N_16370,N_14513);
and U23444 (N_23444,N_15456,N_15492);
or U23445 (N_23445,N_15347,N_17842);
and U23446 (N_23446,N_12690,N_16578);
nor U23447 (N_23447,N_13873,N_17337);
or U23448 (N_23448,N_14316,N_16247);
nor U23449 (N_23449,N_14375,N_13977);
or U23450 (N_23450,N_15642,N_13115);
or U23451 (N_23451,N_17967,N_17956);
nor U23452 (N_23452,N_14239,N_17104);
nand U23453 (N_23453,N_13166,N_15511);
or U23454 (N_23454,N_15902,N_13723);
nor U23455 (N_23455,N_17772,N_15518);
and U23456 (N_23456,N_16527,N_13745);
or U23457 (N_23457,N_14891,N_17739);
or U23458 (N_23458,N_15083,N_14073);
nor U23459 (N_23459,N_13492,N_15264);
nand U23460 (N_23460,N_12526,N_14179);
or U23461 (N_23461,N_15019,N_13777);
or U23462 (N_23462,N_13359,N_13101);
and U23463 (N_23463,N_14530,N_17252);
nand U23464 (N_23464,N_14205,N_12217);
and U23465 (N_23465,N_12694,N_15239);
xor U23466 (N_23466,N_12470,N_12111);
xnor U23467 (N_23467,N_13507,N_14257);
and U23468 (N_23468,N_15431,N_16368);
and U23469 (N_23469,N_12310,N_12991);
nor U23470 (N_23470,N_15190,N_13241);
nand U23471 (N_23471,N_16482,N_13587);
nand U23472 (N_23472,N_17509,N_16778);
nor U23473 (N_23473,N_13569,N_15477);
and U23474 (N_23474,N_15555,N_13993);
and U23475 (N_23475,N_17901,N_15529);
or U23476 (N_23476,N_12736,N_15871);
nor U23477 (N_23477,N_15488,N_14516);
xnor U23478 (N_23478,N_15141,N_15775);
and U23479 (N_23479,N_12911,N_14011);
and U23480 (N_23480,N_13461,N_15644);
or U23481 (N_23481,N_15707,N_12354);
or U23482 (N_23482,N_14497,N_12693);
nor U23483 (N_23483,N_14330,N_13724);
nor U23484 (N_23484,N_13830,N_17718);
or U23485 (N_23485,N_16801,N_12518);
nor U23486 (N_23486,N_16540,N_17397);
nand U23487 (N_23487,N_14925,N_16170);
nand U23488 (N_23488,N_13575,N_12276);
and U23489 (N_23489,N_13932,N_15888);
nand U23490 (N_23490,N_15487,N_13379);
and U23491 (N_23491,N_12241,N_17299);
or U23492 (N_23492,N_14690,N_14834);
and U23493 (N_23493,N_14560,N_17124);
or U23494 (N_23494,N_15284,N_14981);
xor U23495 (N_23495,N_16696,N_17801);
nor U23496 (N_23496,N_12797,N_12880);
nand U23497 (N_23497,N_12730,N_14405);
and U23498 (N_23498,N_12360,N_12116);
or U23499 (N_23499,N_13470,N_12600);
nor U23500 (N_23500,N_13937,N_15038);
and U23501 (N_23501,N_12482,N_14112);
nor U23502 (N_23502,N_15817,N_13116);
xnor U23503 (N_23503,N_17943,N_17673);
xnor U23504 (N_23504,N_16067,N_17822);
and U23505 (N_23505,N_13872,N_17681);
or U23506 (N_23506,N_15075,N_17375);
xnor U23507 (N_23507,N_16308,N_15360);
nor U23508 (N_23508,N_15528,N_17977);
nand U23509 (N_23509,N_17707,N_16164);
nor U23510 (N_23510,N_16255,N_13370);
nand U23511 (N_23511,N_17713,N_13398);
and U23512 (N_23512,N_15582,N_16302);
nand U23513 (N_23513,N_13039,N_12790);
nor U23514 (N_23514,N_12352,N_17096);
nor U23515 (N_23515,N_16482,N_17329);
nand U23516 (N_23516,N_13670,N_13097);
or U23517 (N_23517,N_12446,N_16473);
xnor U23518 (N_23518,N_17255,N_13172);
nand U23519 (N_23519,N_12631,N_13335);
nand U23520 (N_23520,N_14763,N_12655);
nand U23521 (N_23521,N_14895,N_15660);
nor U23522 (N_23522,N_14916,N_16783);
nand U23523 (N_23523,N_12408,N_15943);
xnor U23524 (N_23524,N_16866,N_14385);
or U23525 (N_23525,N_17165,N_16218);
or U23526 (N_23526,N_14912,N_15458);
or U23527 (N_23527,N_12756,N_15444);
or U23528 (N_23528,N_15626,N_14647);
xor U23529 (N_23529,N_14546,N_14452);
xor U23530 (N_23530,N_15059,N_16661);
or U23531 (N_23531,N_13678,N_14151);
xnor U23532 (N_23532,N_12399,N_12676);
nand U23533 (N_23533,N_16445,N_15956);
and U23534 (N_23534,N_13854,N_14979);
xor U23535 (N_23535,N_13777,N_17060);
nor U23536 (N_23536,N_15300,N_13101);
nor U23537 (N_23537,N_12679,N_16556);
and U23538 (N_23538,N_12442,N_15893);
nand U23539 (N_23539,N_15195,N_14463);
nand U23540 (N_23540,N_17511,N_13545);
and U23541 (N_23541,N_13242,N_17517);
or U23542 (N_23542,N_17855,N_14849);
nor U23543 (N_23543,N_14644,N_17005);
or U23544 (N_23544,N_17596,N_17840);
nor U23545 (N_23545,N_16591,N_15553);
and U23546 (N_23546,N_12629,N_17342);
nand U23547 (N_23547,N_13464,N_16723);
nor U23548 (N_23548,N_17863,N_14840);
nand U23549 (N_23549,N_15422,N_15279);
or U23550 (N_23550,N_12790,N_15020);
xnor U23551 (N_23551,N_15495,N_12270);
and U23552 (N_23552,N_14129,N_15705);
nand U23553 (N_23553,N_15903,N_15629);
or U23554 (N_23554,N_14207,N_16605);
or U23555 (N_23555,N_16230,N_16515);
xor U23556 (N_23556,N_15408,N_15807);
or U23557 (N_23557,N_16493,N_14254);
or U23558 (N_23558,N_12299,N_12880);
and U23559 (N_23559,N_14820,N_12653);
or U23560 (N_23560,N_13238,N_13441);
and U23561 (N_23561,N_12098,N_17498);
or U23562 (N_23562,N_13662,N_13454);
nor U23563 (N_23563,N_17273,N_15946);
and U23564 (N_23564,N_16445,N_17340);
or U23565 (N_23565,N_17691,N_17698);
and U23566 (N_23566,N_15020,N_14249);
nor U23567 (N_23567,N_16622,N_14634);
nand U23568 (N_23568,N_17763,N_14666);
nand U23569 (N_23569,N_16440,N_14333);
or U23570 (N_23570,N_17796,N_15897);
nor U23571 (N_23571,N_12380,N_15252);
nor U23572 (N_23572,N_17403,N_16002);
nor U23573 (N_23573,N_14730,N_15378);
xor U23574 (N_23574,N_12415,N_16104);
nor U23575 (N_23575,N_16933,N_17329);
and U23576 (N_23576,N_16511,N_14295);
xnor U23577 (N_23577,N_13915,N_14733);
or U23578 (N_23578,N_13819,N_13211);
nand U23579 (N_23579,N_17464,N_14332);
or U23580 (N_23580,N_14389,N_12862);
and U23581 (N_23581,N_14179,N_15447);
nand U23582 (N_23582,N_13633,N_15054);
nor U23583 (N_23583,N_15784,N_16735);
or U23584 (N_23584,N_17457,N_15254);
and U23585 (N_23585,N_16408,N_12451);
and U23586 (N_23586,N_13880,N_16160);
nor U23587 (N_23587,N_15916,N_17736);
xnor U23588 (N_23588,N_12126,N_16927);
nand U23589 (N_23589,N_15273,N_14415);
nand U23590 (N_23590,N_17547,N_13638);
xnor U23591 (N_23591,N_15316,N_16273);
nand U23592 (N_23592,N_14691,N_15375);
nand U23593 (N_23593,N_14705,N_16551);
nand U23594 (N_23594,N_15869,N_12536);
nor U23595 (N_23595,N_14288,N_15709);
nor U23596 (N_23596,N_15884,N_15523);
nor U23597 (N_23597,N_15644,N_14232);
nand U23598 (N_23598,N_12641,N_17782);
nand U23599 (N_23599,N_14902,N_12800);
nor U23600 (N_23600,N_12047,N_16076);
and U23601 (N_23601,N_12433,N_15993);
and U23602 (N_23602,N_15946,N_14874);
or U23603 (N_23603,N_17720,N_16555);
nand U23604 (N_23604,N_16120,N_13835);
and U23605 (N_23605,N_12134,N_14361);
nand U23606 (N_23606,N_16258,N_13145);
nor U23607 (N_23607,N_16435,N_12196);
nand U23608 (N_23608,N_17120,N_13438);
nand U23609 (N_23609,N_15980,N_13076);
or U23610 (N_23610,N_15824,N_12934);
nor U23611 (N_23611,N_13852,N_13766);
or U23612 (N_23612,N_15247,N_16069);
nor U23613 (N_23613,N_17731,N_15246);
or U23614 (N_23614,N_14753,N_15268);
nand U23615 (N_23615,N_17288,N_12795);
nor U23616 (N_23616,N_14101,N_13262);
xor U23617 (N_23617,N_12186,N_16719);
nand U23618 (N_23618,N_12686,N_16834);
or U23619 (N_23619,N_12797,N_16382);
xor U23620 (N_23620,N_15034,N_16879);
or U23621 (N_23621,N_17353,N_17620);
and U23622 (N_23622,N_17972,N_14959);
xor U23623 (N_23623,N_16383,N_13648);
nor U23624 (N_23624,N_16590,N_15604);
nor U23625 (N_23625,N_16876,N_12006);
or U23626 (N_23626,N_17786,N_16184);
or U23627 (N_23627,N_12845,N_16185);
xor U23628 (N_23628,N_14662,N_17512);
or U23629 (N_23629,N_17735,N_12458);
and U23630 (N_23630,N_16624,N_17200);
and U23631 (N_23631,N_16406,N_15476);
nand U23632 (N_23632,N_15907,N_16815);
or U23633 (N_23633,N_14840,N_16745);
nor U23634 (N_23634,N_13014,N_16857);
nand U23635 (N_23635,N_12716,N_13204);
nor U23636 (N_23636,N_12131,N_16612);
xnor U23637 (N_23637,N_15216,N_13769);
or U23638 (N_23638,N_15211,N_12410);
and U23639 (N_23639,N_12911,N_12959);
and U23640 (N_23640,N_14050,N_16410);
or U23641 (N_23641,N_15155,N_17259);
or U23642 (N_23642,N_13367,N_12464);
or U23643 (N_23643,N_17396,N_14741);
or U23644 (N_23644,N_12653,N_17426);
nor U23645 (N_23645,N_14596,N_12787);
or U23646 (N_23646,N_14027,N_13927);
xnor U23647 (N_23647,N_15156,N_15532);
nand U23648 (N_23648,N_14928,N_17083);
or U23649 (N_23649,N_17657,N_16685);
and U23650 (N_23650,N_17306,N_13897);
nor U23651 (N_23651,N_13885,N_14569);
nor U23652 (N_23652,N_17070,N_16707);
nor U23653 (N_23653,N_13241,N_17404);
xor U23654 (N_23654,N_16665,N_17633);
xor U23655 (N_23655,N_17534,N_15204);
or U23656 (N_23656,N_12587,N_14339);
or U23657 (N_23657,N_15903,N_15580);
nand U23658 (N_23658,N_15730,N_15906);
nor U23659 (N_23659,N_14747,N_17188);
and U23660 (N_23660,N_12233,N_15802);
nor U23661 (N_23661,N_15249,N_14593);
xor U23662 (N_23662,N_12413,N_15226);
xor U23663 (N_23663,N_15181,N_13126);
and U23664 (N_23664,N_17646,N_16187);
nor U23665 (N_23665,N_13106,N_12905);
xnor U23666 (N_23666,N_15190,N_12738);
xnor U23667 (N_23667,N_14660,N_16188);
or U23668 (N_23668,N_15324,N_14024);
nand U23669 (N_23669,N_12294,N_14791);
and U23670 (N_23670,N_15586,N_14786);
nand U23671 (N_23671,N_16819,N_16326);
nand U23672 (N_23672,N_12290,N_13583);
and U23673 (N_23673,N_16117,N_14897);
or U23674 (N_23674,N_13056,N_13238);
xor U23675 (N_23675,N_14110,N_12249);
xnor U23676 (N_23676,N_16636,N_12582);
or U23677 (N_23677,N_12672,N_15260);
xnor U23678 (N_23678,N_15787,N_12201);
and U23679 (N_23679,N_17296,N_13607);
or U23680 (N_23680,N_14665,N_13638);
and U23681 (N_23681,N_17727,N_16136);
nand U23682 (N_23682,N_13458,N_16794);
nand U23683 (N_23683,N_17822,N_15491);
nand U23684 (N_23684,N_15069,N_14204);
or U23685 (N_23685,N_15965,N_15867);
or U23686 (N_23686,N_16574,N_16657);
nand U23687 (N_23687,N_16545,N_17782);
nor U23688 (N_23688,N_12264,N_14912);
nand U23689 (N_23689,N_16183,N_15010);
nand U23690 (N_23690,N_14939,N_15769);
nor U23691 (N_23691,N_15287,N_12548);
nand U23692 (N_23692,N_15016,N_13195);
nand U23693 (N_23693,N_12204,N_14620);
or U23694 (N_23694,N_16496,N_13894);
xnor U23695 (N_23695,N_17971,N_16171);
xnor U23696 (N_23696,N_14898,N_17871);
nor U23697 (N_23697,N_13891,N_17225);
xnor U23698 (N_23698,N_16861,N_12325);
or U23699 (N_23699,N_14770,N_17428);
nand U23700 (N_23700,N_13762,N_12716);
or U23701 (N_23701,N_15803,N_13432);
nor U23702 (N_23702,N_15937,N_12056);
or U23703 (N_23703,N_14796,N_15195);
nor U23704 (N_23704,N_16576,N_14255);
and U23705 (N_23705,N_13536,N_16655);
xnor U23706 (N_23706,N_15036,N_13274);
and U23707 (N_23707,N_15294,N_14504);
nor U23708 (N_23708,N_12600,N_16136);
nor U23709 (N_23709,N_17752,N_13874);
nand U23710 (N_23710,N_12572,N_14015);
nand U23711 (N_23711,N_12096,N_17679);
xnor U23712 (N_23712,N_12116,N_17381);
nand U23713 (N_23713,N_12845,N_16745);
xor U23714 (N_23714,N_13765,N_12336);
xor U23715 (N_23715,N_17618,N_17415);
or U23716 (N_23716,N_12446,N_13703);
and U23717 (N_23717,N_16269,N_15630);
or U23718 (N_23718,N_13066,N_15836);
nand U23719 (N_23719,N_13966,N_13208);
nand U23720 (N_23720,N_17280,N_13630);
and U23721 (N_23721,N_17567,N_13239);
nand U23722 (N_23722,N_12082,N_13600);
nand U23723 (N_23723,N_12859,N_13421);
or U23724 (N_23724,N_12639,N_13635);
nor U23725 (N_23725,N_16896,N_14890);
nor U23726 (N_23726,N_13469,N_14513);
nand U23727 (N_23727,N_14468,N_15983);
nor U23728 (N_23728,N_12766,N_13300);
nand U23729 (N_23729,N_14388,N_17345);
nand U23730 (N_23730,N_15603,N_15324);
nor U23731 (N_23731,N_16538,N_14878);
nor U23732 (N_23732,N_13469,N_13732);
or U23733 (N_23733,N_13062,N_14513);
or U23734 (N_23734,N_13048,N_14902);
nor U23735 (N_23735,N_17873,N_12636);
and U23736 (N_23736,N_16417,N_12543);
xnor U23737 (N_23737,N_14553,N_17761);
nor U23738 (N_23738,N_17740,N_13111);
or U23739 (N_23739,N_13713,N_12019);
and U23740 (N_23740,N_13718,N_17688);
xor U23741 (N_23741,N_15381,N_16669);
and U23742 (N_23742,N_17825,N_15529);
xnor U23743 (N_23743,N_14594,N_15322);
nand U23744 (N_23744,N_14987,N_15529);
nand U23745 (N_23745,N_16542,N_13513);
nand U23746 (N_23746,N_16431,N_14306);
nor U23747 (N_23747,N_16323,N_13216);
xor U23748 (N_23748,N_13519,N_12772);
xnor U23749 (N_23749,N_17116,N_13970);
nand U23750 (N_23750,N_13758,N_13003);
nor U23751 (N_23751,N_14460,N_12536);
nor U23752 (N_23752,N_13342,N_13195);
or U23753 (N_23753,N_12385,N_17543);
nand U23754 (N_23754,N_15948,N_14851);
or U23755 (N_23755,N_12369,N_17917);
and U23756 (N_23756,N_13722,N_14698);
and U23757 (N_23757,N_13317,N_15421);
and U23758 (N_23758,N_15611,N_17994);
nor U23759 (N_23759,N_16774,N_12611);
or U23760 (N_23760,N_14231,N_16904);
xnor U23761 (N_23761,N_16348,N_14819);
nand U23762 (N_23762,N_17589,N_13024);
nand U23763 (N_23763,N_16037,N_12737);
and U23764 (N_23764,N_12742,N_12689);
nor U23765 (N_23765,N_17021,N_12503);
nor U23766 (N_23766,N_15513,N_15876);
nand U23767 (N_23767,N_12043,N_13451);
or U23768 (N_23768,N_12694,N_15471);
and U23769 (N_23769,N_13495,N_15955);
nand U23770 (N_23770,N_15789,N_16223);
or U23771 (N_23771,N_15861,N_16601);
xnor U23772 (N_23772,N_15139,N_13159);
and U23773 (N_23773,N_12604,N_16099);
nand U23774 (N_23774,N_17687,N_16783);
or U23775 (N_23775,N_16493,N_12535);
nor U23776 (N_23776,N_12449,N_14467);
nand U23777 (N_23777,N_16791,N_13201);
nor U23778 (N_23778,N_16745,N_16437);
nand U23779 (N_23779,N_15166,N_15502);
nand U23780 (N_23780,N_17045,N_15729);
nor U23781 (N_23781,N_17149,N_13847);
xnor U23782 (N_23782,N_12798,N_15800);
nand U23783 (N_23783,N_14206,N_13768);
xnor U23784 (N_23784,N_17067,N_16653);
nand U23785 (N_23785,N_13274,N_15691);
nand U23786 (N_23786,N_17490,N_17234);
xor U23787 (N_23787,N_15446,N_14391);
and U23788 (N_23788,N_15365,N_14699);
and U23789 (N_23789,N_14208,N_16139);
or U23790 (N_23790,N_12692,N_16388);
or U23791 (N_23791,N_16754,N_16145);
nor U23792 (N_23792,N_15203,N_12682);
nor U23793 (N_23793,N_15604,N_12428);
nor U23794 (N_23794,N_12492,N_12347);
and U23795 (N_23795,N_13755,N_13118);
or U23796 (N_23796,N_12360,N_14822);
and U23797 (N_23797,N_13371,N_17682);
nand U23798 (N_23798,N_14984,N_12326);
nand U23799 (N_23799,N_13312,N_15865);
nand U23800 (N_23800,N_13454,N_13466);
nor U23801 (N_23801,N_17075,N_13147);
or U23802 (N_23802,N_13111,N_12069);
nor U23803 (N_23803,N_13618,N_13437);
nand U23804 (N_23804,N_15652,N_15907);
or U23805 (N_23805,N_13759,N_13421);
nand U23806 (N_23806,N_12442,N_12782);
nor U23807 (N_23807,N_16161,N_12834);
or U23808 (N_23808,N_16263,N_14139);
nor U23809 (N_23809,N_15185,N_14626);
xor U23810 (N_23810,N_12979,N_13735);
nand U23811 (N_23811,N_16067,N_16592);
or U23812 (N_23812,N_12987,N_15296);
xor U23813 (N_23813,N_15962,N_17062);
and U23814 (N_23814,N_17174,N_12197);
nand U23815 (N_23815,N_17336,N_17129);
and U23816 (N_23816,N_15196,N_14593);
xnor U23817 (N_23817,N_17601,N_15969);
xor U23818 (N_23818,N_12638,N_14547);
nand U23819 (N_23819,N_16036,N_13497);
nand U23820 (N_23820,N_16141,N_16181);
xor U23821 (N_23821,N_14443,N_12001);
and U23822 (N_23822,N_16444,N_16849);
nor U23823 (N_23823,N_12261,N_14071);
nand U23824 (N_23824,N_17092,N_12845);
or U23825 (N_23825,N_16771,N_12139);
or U23826 (N_23826,N_17436,N_12669);
and U23827 (N_23827,N_12680,N_13777);
or U23828 (N_23828,N_14512,N_15762);
xnor U23829 (N_23829,N_16116,N_17217);
nand U23830 (N_23830,N_17120,N_17445);
nor U23831 (N_23831,N_15213,N_16034);
nand U23832 (N_23832,N_16585,N_15113);
or U23833 (N_23833,N_16979,N_16662);
nor U23834 (N_23834,N_12191,N_17492);
and U23835 (N_23835,N_12174,N_16781);
or U23836 (N_23836,N_12060,N_14754);
nor U23837 (N_23837,N_14610,N_14483);
and U23838 (N_23838,N_14777,N_16477);
nand U23839 (N_23839,N_14460,N_16662);
or U23840 (N_23840,N_15766,N_12811);
xor U23841 (N_23841,N_17500,N_15080);
nor U23842 (N_23842,N_12057,N_14054);
xor U23843 (N_23843,N_12985,N_15510);
nor U23844 (N_23844,N_14222,N_17852);
and U23845 (N_23845,N_17635,N_14156);
and U23846 (N_23846,N_15434,N_17746);
nand U23847 (N_23847,N_16030,N_14370);
nand U23848 (N_23848,N_16040,N_13378);
or U23849 (N_23849,N_13049,N_17181);
nand U23850 (N_23850,N_15699,N_13042);
or U23851 (N_23851,N_13540,N_16794);
and U23852 (N_23852,N_15555,N_14189);
or U23853 (N_23853,N_16048,N_14034);
nand U23854 (N_23854,N_12593,N_14402);
or U23855 (N_23855,N_14644,N_16615);
or U23856 (N_23856,N_16063,N_14521);
nor U23857 (N_23857,N_12852,N_15395);
or U23858 (N_23858,N_14872,N_16715);
nand U23859 (N_23859,N_17525,N_13433);
or U23860 (N_23860,N_12556,N_12304);
xor U23861 (N_23861,N_17672,N_17772);
nand U23862 (N_23862,N_12398,N_13114);
nor U23863 (N_23863,N_16389,N_17924);
xnor U23864 (N_23864,N_14483,N_12320);
or U23865 (N_23865,N_15463,N_15441);
and U23866 (N_23866,N_15114,N_14701);
or U23867 (N_23867,N_15985,N_14418);
xnor U23868 (N_23868,N_16724,N_12454);
xor U23869 (N_23869,N_15357,N_12171);
xor U23870 (N_23870,N_12387,N_13353);
and U23871 (N_23871,N_15795,N_12470);
nor U23872 (N_23872,N_14603,N_16088);
and U23873 (N_23873,N_15752,N_12591);
nor U23874 (N_23874,N_14172,N_16094);
and U23875 (N_23875,N_13911,N_12444);
xor U23876 (N_23876,N_17889,N_13833);
xor U23877 (N_23877,N_14848,N_16252);
nor U23878 (N_23878,N_16148,N_16430);
nor U23879 (N_23879,N_13124,N_17130);
nand U23880 (N_23880,N_16737,N_13629);
or U23881 (N_23881,N_15330,N_12676);
or U23882 (N_23882,N_17010,N_14223);
nor U23883 (N_23883,N_16106,N_15019);
and U23884 (N_23884,N_16440,N_12164);
or U23885 (N_23885,N_17569,N_17575);
and U23886 (N_23886,N_17751,N_12226);
nand U23887 (N_23887,N_16484,N_17609);
and U23888 (N_23888,N_12656,N_13710);
and U23889 (N_23889,N_15578,N_14437);
or U23890 (N_23890,N_15221,N_16486);
nor U23891 (N_23891,N_14690,N_13683);
nand U23892 (N_23892,N_17942,N_13674);
nand U23893 (N_23893,N_16787,N_15652);
nor U23894 (N_23894,N_13258,N_16342);
nand U23895 (N_23895,N_15631,N_13926);
or U23896 (N_23896,N_12861,N_13509);
nand U23897 (N_23897,N_16695,N_12111);
xnor U23898 (N_23898,N_16985,N_17535);
xnor U23899 (N_23899,N_17077,N_13886);
and U23900 (N_23900,N_12855,N_15250);
nor U23901 (N_23901,N_17308,N_15924);
or U23902 (N_23902,N_12773,N_13512);
nand U23903 (N_23903,N_14053,N_16363);
and U23904 (N_23904,N_12173,N_17418);
and U23905 (N_23905,N_16978,N_15607);
nor U23906 (N_23906,N_17924,N_13830);
and U23907 (N_23907,N_13464,N_17104);
nor U23908 (N_23908,N_17530,N_12441);
nand U23909 (N_23909,N_14879,N_14003);
nand U23910 (N_23910,N_15378,N_12593);
xor U23911 (N_23911,N_17684,N_13871);
and U23912 (N_23912,N_17768,N_15187);
xnor U23913 (N_23913,N_13480,N_13823);
xor U23914 (N_23914,N_12205,N_12796);
and U23915 (N_23915,N_16639,N_14759);
or U23916 (N_23916,N_12742,N_12767);
or U23917 (N_23917,N_14325,N_16388);
nand U23918 (N_23918,N_14591,N_13799);
or U23919 (N_23919,N_17499,N_17752);
or U23920 (N_23920,N_15293,N_14812);
and U23921 (N_23921,N_16356,N_17375);
xnor U23922 (N_23922,N_17882,N_14852);
xnor U23923 (N_23923,N_17797,N_15023);
and U23924 (N_23924,N_16297,N_16505);
xor U23925 (N_23925,N_16894,N_12239);
nor U23926 (N_23926,N_17596,N_14800);
nor U23927 (N_23927,N_17294,N_16366);
and U23928 (N_23928,N_14263,N_17326);
and U23929 (N_23929,N_14176,N_16085);
nor U23930 (N_23930,N_13383,N_14734);
and U23931 (N_23931,N_17130,N_15670);
xnor U23932 (N_23932,N_12997,N_16994);
and U23933 (N_23933,N_12537,N_16487);
and U23934 (N_23934,N_12721,N_12124);
xnor U23935 (N_23935,N_12753,N_14353);
and U23936 (N_23936,N_12128,N_12650);
nor U23937 (N_23937,N_15057,N_12749);
nor U23938 (N_23938,N_12170,N_14868);
xor U23939 (N_23939,N_17141,N_16207);
xnor U23940 (N_23940,N_16421,N_13100);
or U23941 (N_23941,N_13446,N_14724);
nand U23942 (N_23942,N_12629,N_14734);
xnor U23943 (N_23943,N_16200,N_14878);
nor U23944 (N_23944,N_12318,N_15933);
xor U23945 (N_23945,N_16864,N_16429);
nor U23946 (N_23946,N_12799,N_16186);
or U23947 (N_23947,N_15054,N_17682);
or U23948 (N_23948,N_12282,N_14399);
nor U23949 (N_23949,N_12774,N_16058);
nand U23950 (N_23950,N_12189,N_16208);
xor U23951 (N_23951,N_13755,N_17984);
xor U23952 (N_23952,N_16878,N_16125);
and U23953 (N_23953,N_15619,N_17217);
xor U23954 (N_23954,N_17663,N_16677);
and U23955 (N_23955,N_14016,N_15203);
xnor U23956 (N_23956,N_17983,N_12322);
xor U23957 (N_23957,N_17221,N_13806);
nand U23958 (N_23958,N_15985,N_12106);
nand U23959 (N_23959,N_17569,N_12816);
nor U23960 (N_23960,N_17348,N_13528);
nand U23961 (N_23961,N_17234,N_15300);
or U23962 (N_23962,N_13107,N_13737);
or U23963 (N_23963,N_17845,N_15655);
nor U23964 (N_23964,N_13249,N_12903);
nor U23965 (N_23965,N_16999,N_14676);
nor U23966 (N_23966,N_15138,N_16108);
xor U23967 (N_23967,N_14933,N_12931);
nor U23968 (N_23968,N_17963,N_14492);
nand U23969 (N_23969,N_15930,N_17448);
and U23970 (N_23970,N_12139,N_13702);
xnor U23971 (N_23971,N_16097,N_15501);
xnor U23972 (N_23972,N_14132,N_15070);
and U23973 (N_23973,N_14978,N_17676);
xor U23974 (N_23974,N_13742,N_15806);
or U23975 (N_23975,N_12697,N_13670);
nor U23976 (N_23976,N_13342,N_17949);
xnor U23977 (N_23977,N_13109,N_13739);
nor U23978 (N_23978,N_17811,N_12234);
nor U23979 (N_23979,N_12309,N_15210);
and U23980 (N_23980,N_14966,N_15199);
nand U23981 (N_23981,N_15169,N_14943);
and U23982 (N_23982,N_15676,N_14977);
nor U23983 (N_23983,N_16290,N_15814);
nor U23984 (N_23984,N_12069,N_13427);
xnor U23985 (N_23985,N_14064,N_16372);
or U23986 (N_23986,N_14812,N_15982);
and U23987 (N_23987,N_16106,N_12818);
nor U23988 (N_23988,N_14510,N_15931);
xor U23989 (N_23989,N_12273,N_12685);
and U23990 (N_23990,N_13329,N_16107);
xor U23991 (N_23991,N_16339,N_14173);
nand U23992 (N_23992,N_17020,N_12385);
and U23993 (N_23993,N_12468,N_15257);
or U23994 (N_23994,N_13695,N_16276);
xor U23995 (N_23995,N_16240,N_12978);
or U23996 (N_23996,N_12804,N_14053);
nand U23997 (N_23997,N_17631,N_12818);
or U23998 (N_23998,N_12053,N_12849);
and U23999 (N_23999,N_17339,N_16455);
nor U24000 (N_24000,N_18061,N_23551);
or U24001 (N_24001,N_22164,N_22355);
nand U24002 (N_24002,N_18723,N_22056);
nand U24003 (N_24003,N_23356,N_23616);
nand U24004 (N_24004,N_22444,N_19337);
nand U24005 (N_24005,N_18388,N_19457);
or U24006 (N_24006,N_21557,N_20193);
or U24007 (N_24007,N_19490,N_21509);
or U24008 (N_24008,N_20346,N_22065);
nor U24009 (N_24009,N_22887,N_20101);
nor U24010 (N_24010,N_22769,N_21853);
and U24011 (N_24011,N_21751,N_23598);
xor U24012 (N_24012,N_19630,N_23798);
and U24013 (N_24013,N_21474,N_18341);
nor U24014 (N_24014,N_22699,N_19240);
and U24015 (N_24015,N_22920,N_21738);
or U24016 (N_24016,N_20648,N_20722);
or U24017 (N_24017,N_23420,N_21426);
nand U24018 (N_24018,N_20117,N_21952);
nand U24019 (N_24019,N_21116,N_18133);
xor U24020 (N_24020,N_19577,N_20561);
nand U24021 (N_24021,N_22380,N_22679);
and U24022 (N_24022,N_22029,N_21461);
nor U24023 (N_24023,N_20814,N_23107);
or U24024 (N_24024,N_19592,N_20979);
or U24025 (N_24025,N_20058,N_19778);
or U24026 (N_24026,N_22815,N_21196);
xor U24027 (N_24027,N_20332,N_22497);
or U24028 (N_24028,N_20761,N_20160);
nand U24029 (N_24029,N_23458,N_19154);
nor U24030 (N_24030,N_23821,N_22194);
xor U24031 (N_24031,N_23627,N_19176);
and U24032 (N_24032,N_18486,N_20831);
nor U24033 (N_24033,N_22795,N_20137);
nor U24034 (N_24034,N_20339,N_23635);
nand U24035 (N_24035,N_22547,N_21482);
and U24036 (N_24036,N_21489,N_20978);
xor U24037 (N_24037,N_21723,N_18897);
xor U24038 (N_24038,N_22425,N_18577);
nor U24039 (N_24039,N_20866,N_21925);
or U24040 (N_24040,N_19836,N_21264);
or U24041 (N_24041,N_23118,N_19053);
xor U24042 (N_24042,N_18040,N_20037);
nand U24043 (N_24043,N_18609,N_21206);
nand U24044 (N_24044,N_23923,N_23871);
nor U24045 (N_24045,N_18914,N_20508);
and U24046 (N_24046,N_18640,N_20183);
xor U24047 (N_24047,N_18627,N_20249);
or U24048 (N_24048,N_18999,N_19487);
nor U24049 (N_24049,N_19178,N_20119);
nand U24050 (N_24050,N_18860,N_23605);
or U24051 (N_24051,N_21939,N_19159);
xor U24052 (N_24052,N_22918,N_21987);
xor U24053 (N_24053,N_22138,N_18413);
or U24054 (N_24054,N_20057,N_22664);
or U24055 (N_24055,N_20710,N_19584);
xor U24056 (N_24056,N_22202,N_21997);
nor U24057 (N_24057,N_18219,N_22381);
and U24058 (N_24058,N_18479,N_23610);
xnor U24059 (N_24059,N_23588,N_18262);
xor U24060 (N_24060,N_20076,N_18283);
xor U24061 (N_24061,N_20447,N_20727);
or U24062 (N_24062,N_18801,N_20837);
or U24063 (N_24063,N_19792,N_23590);
nand U24064 (N_24064,N_21859,N_21917);
or U24065 (N_24065,N_19498,N_20389);
or U24066 (N_24066,N_21831,N_20211);
xnor U24067 (N_24067,N_23484,N_22790);
or U24068 (N_24068,N_20194,N_22717);
xor U24069 (N_24069,N_23796,N_19274);
xor U24070 (N_24070,N_19064,N_23761);
xnor U24071 (N_24071,N_21942,N_20421);
xnor U24072 (N_24072,N_18037,N_23989);
and U24073 (N_24073,N_21096,N_18724);
nand U24074 (N_24074,N_19122,N_20751);
and U24075 (N_24075,N_23323,N_18543);
nor U24076 (N_24076,N_20683,N_20056);
nand U24077 (N_24077,N_21944,N_19935);
xnor U24078 (N_24078,N_23535,N_20155);
xor U24079 (N_24079,N_19761,N_19162);
or U24080 (N_24080,N_22373,N_18440);
or U24081 (N_24081,N_19619,N_20207);
and U24082 (N_24082,N_18195,N_18359);
nand U24083 (N_24083,N_19010,N_22148);
nor U24084 (N_24084,N_21608,N_22615);
xor U24085 (N_24085,N_19067,N_18296);
or U24086 (N_24086,N_18209,N_19206);
nor U24087 (N_24087,N_21636,N_20904);
nand U24088 (N_24088,N_21869,N_22191);
xor U24089 (N_24089,N_20908,N_18474);
nand U24090 (N_24090,N_22124,N_22299);
or U24091 (N_24091,N_19462,N_23060);
nor U24092 (N_24092,N_19124,N_19934);
and U24093 (N_24093,N_20413,N_22938);
or U24094 (N_24094,N_23999,N_21329);
xnor U24095 (N_24095,N_19833,N_23864);
xnor U24096 (N_24096,N_18302,N_23565);
nand U24097 (N_24097,N_22489,N_21356);
xor U24098 (N_24098,N_22017,N_22341);
xor U24099 (N_24099,N_22290,N_20475);
or U24100 (N_24100,N_19597,N_21178);
nand U24101 (N_24101,N_22180,N_19629);
nor U24102 (N_24102,N_20450,N_22632);
and U24103 (N_24103,N_19397,N_21388);
nand U24104 (N_24104,N_18258,N_23813);
or U24105 (N_24105,N_18533,N_20747);
xor U24106 (N_24106,N_18395,N_22586);
nor U24107 (N_24107,N_18631,N_19327);
and U24108 (N_24108,N_23106,N_23500);
xnor U24109 (N_24109,N_20457,N_20403);
nor U24110 (N_24110,N_19252,N_23325);
xnor U24111 (N_24111,N_19062,N_20542);
nor U24112 (N_24112,N_23329,N_23430);
or U24113 (N_24113,N_19423,N_21275);
nand U24114 (N_24114,N_22889,N_20750);
xor U24115 (N_24115,N_18214,N_21445);
and U24116 (N_24116,N_20243,N_18957);
nor U24117 (N_24117,N_18535,N_21501);
nor U24118 (N_24118,N_19198,N_22727);
nand U24119 (N_24119,N_22430,N_22197);
and U24120 (N_24120,N_20601,N_23976);
nor U24121 (N_24121,N_18970,N_23443);
nand U24122 (N_24122,N_21247,N_23874);
nor U24123 (N_24123,N_21915,N_22096);
or U24124 (N_24124,N_21435,N_19455);
nor U24125 (N_24125,N_21644,N_18152);
xor U24126 (N_24126,N_19434,N_23956);
nand U24127 (N_24127,N_19098,N_22859);
and U24128 (N_24128,N_19039,N_22480);
and U24129 (N_24129,N_20417,N_21778);
nor U24130 (N_24130,N_20643,N_19142);
xnor U24131 (N_24131,N_22808,N_18688);
or U24132 (N_24132,N_23052,N_19869);
nand U24133 (N_24133,N_18514,N_18298);
and U24134 (N_24134,N_19486,N_22090);
xnor U24135 (N_24135,N_18008,N_18216);
xnor U24136 (N_24136,N_21397,N_20340);
xor U24137 (N_24137,N_23068,N_19231);
nor U24138 (N_24138,N_21232,N_22143);
or U24139 (N_24139,N_21009,N_19196);
nor U24140 (N_24140,N_22289,N_19849);
xnor U24141 (N_24141,N_19071,N_21121);
nand U24142 (N_24142,N_21289,N_19601);
or U24143 (N_24143,N_20479,N_22357);
or U24144 (N_24144,N_19336,N_21606);
and U24145 (N_24145,N_21671,N_23340);
nor U24146 (N_24146,N_19741,N_18944);
or U24147 (N_24147,N_20480,N_21787);
nand U24148 (N_24148,N_19326,N_23379);
nor U24149 (N_24149,N_20506,N_23926);
and U24150 (N_24150,N_18975,N_19082);
and U24151 (N_24151,N_21662,N_20846);
or U24152 (N_24152,N_23130,N_19729);
or U24153 (N_24153,N_22418,N_19179);
nand U24154 (N_24154,N_18929,N_22944);
nand U24155 (N_24155,N_20008,N_20014);
or U24156 (N_24156,N_23488,N_22494);
xor U24157 (N_24157,N_21286,N_18843);
xor U24158 (N_24158,N_18115,N_20826);
and U24159 (N_24159,N_22121,N_20865);
xor U24160 (N_24160,N_18267,N_18222);
and U24161 (N_24161,N_22565,N_23811);
xor U24162 (N_24162,N_23364,N_22453);
or U24163 (N_24163,N_22222,N_19727);
and U24164 (N_24164,N_20314,N_18541);
or U24165 (N_24165,N_18727,N_21358);
or U24166 (N_24166,N_22362,N_20595);
nor U24167 (N_24167,N_23229,N_19746);
nand U24168 (N_24168,N_23782,N_22916);
nor U24169 (N_24169,N_19234,N_21188);
nand U24170 (N_24170,N_19535,N_20639);
nand U24171 (N_24171,N_18123,N_21423);
nor U24172 (N_24172,N_19784,N_22467);
nand U24173 (N_24173,N_19607,N_22348);
nand U24174 (N_24174,N_23353,N_21607);
nand U24175 (N_24175,N_20344,N_22957);
and U24176 (N_24176,N_19004,N_20034);
and U24177 (N_24177,N_18063,N_23254);
nor U24178 (N_24178,N_21699,N_22496);
nand U24179 (N_24179,N_23581,N_23680);
or U24180 (N_24180,N_20424,N_21821);
or U24181 (N_24181,N_22302,N_21255);
xor U24182 (N_24182,N_18854,N_20536);
nor U24183 (N_24183,N_21702,N_18278);
and U24184 (N_24184,N_23165,N_22922);
and U24185 (N_24185,N_23149,N_21514);
nor U24186 (N_24186,N_18781,N_18891);
and U24187 (N_24187,N_21389,N_22747);
or U24188 (N_24188,N_18044,N_23925);
nor U24189 (N_24189,N_21937,N_23460);
nor U24190 (N_24190,N_19165,N_23421);
or U24191 (N_24191,N_18976,N_22612);
and U24192 (N_24192,N_23791,N_18839);
nand U24193 (N_24193,N_18177,N_20633);
xnor U24194 (N_24194,N_20329,N_20199);
nor U24195 (N_24195,N_19675,N_21768);
and U24196 (N_24196,N_20774,N_23313);
and U24197 (N_24197,N_23843,N_20619);
xor U24198 (N_24198,N_23144,N_20516);
xnor U24199 (N_24199,N_21830,N_19238);
or U24200 (N_24200,N_22602,N_21626);
or U24201 (N_24201,N_18339,N_23508);
or U24202 (N_24202,N_20621,N_19436);
or U24203 (N_24203,N_18587,N_18469);
or U24204 (N_24204,N_22195,N_23018);
or U24205 (N_24205,N_19489,N_21954);
xnor U24206 (N_24206,N_23301,N_21318);
nor U24207 (N_24207,N_20540,N_23092);
or U24208 (N_24208,N_18538,N_18311);
nor U24209 (N_24209,N_20290,N_18441);
nand U24210 (N_24210,N_19323,N_21039);
nor U24211 (N_24211,N_22970,N_19959);
nand U24212 (N_24212,N_22101,N_23260);
xor U24213 (N_24213,N_23034,N_20238);
or U24214 (N_24214,N_23775,N_22371);
and U24215 (N_24215,N_23636,N_18504);
and U24216 (N_24216,N_20848,N_21585);
nand U24217 (N_24217,N_23647,N_19576);
xnor U24218 (N_24218,N_19172,N_22935);
or U24219 (N_24219,N_21680,N_18299);
xnor U24220 (N_24220,N_22074,N_22926);
or U24221 (N_24221,N_21355,N_19202);
or U24222 (N_24222,N_19979,N_19406);
or U24223 (N_24223,N_19856,N_19570);
nand U24224 (N_24224,N_18066,N_23187);
xnor U24225 (N_24225,N_18360,N_21016);
nor U24226 (N_24226,N_19351,N_22883);
nor U24227 (N_24227,N_18210,N_21569);
nand U24228 (N_24228,N_22345,N_22134);
and U24229 (N_24229,N_21470,N_22842);
xnor U24230 (N_24230,N_18842,N_19542);
and U24231 (N_24231,N_22219,N_19461);
nand U24232 (N_24232,N_19954,N_20179);
and U24233 (N_24233,N_20994,N_20266);
and U24234 (N_24234,N_21105,N_23041);
xor U24235 (N_24235,N_19285,N_18110);
nor U24236 (N_24236,N_22482,N_22158);
nor U24237 (N_24237,N_18900,N_18480);
xor U24238 (N_24238,N_19350,N_20330);
xor U24239 (N_24239,N_23897,N_21238);
or U24240 (N_24240,N_22526,N_18766);
nand U24241 (N_24241,N_22420,N_21635);
xnor U24242 (N_24242,N_22989,N_20322);
nor U24243 (N_24243,N_18191,N_22672);
xor U24244 (N_24244,N_21234,N_19250);
xnor U24245 (N_24245,N_23157,N_20033);
or U24246 (N_24246,N_19025,N_22503);
nand U24247 (N_24247,N_21604,N_23634);
and U24248 (N_24248,N_22917,N_20018);
nor U24249 (N_24249,N_22083,N_18620);
and U24250 (N_24250,N_19569,N_19107);
nand U24251 (N_24251,N_22495,N_22667);
and U24252 (N_24252,N_23218,N_18990);
nand U24253 (N_24253,N_18899,N_18259);
and U24254 (N_24254,N_21120,N_21686);
and U24255 (N_24255,N_22486,N_21624);
xnor U24256 (N_24256,N_18977,N_19665);
xnor U24257 (N_24257,N_21008,N_21602);
and U24258 (N_24258,N_21341,N_22811);
xor U24259 (N_24259,N_20736,N_20562);
and U24260 (N_24260,N_20154,N_23583);
nor U24261 (N_24261,N_19735,N_23790);
xor U24262 (N_24262,N_18372,N_20684);
nand U24263 (N_24263,N_20597,N_23110);
nand U24264 (N_24264,N_19043,N_21259);
nor U24265 (N_24265,N_19783,N_22548);
nand U24266 (N_24266,N_20105,N_21776);
nor U24267 (N_24267,N_22974,N_18104);
nand U24268 (N_24268,N_19550,N_18552);
nor U24269 (N_24269,N_20434,N_19505);
or U24270 (N_24270,N_18266,N_18599);
or U24271 (N_24271,N_18771,N_23071);
and U24272 (N_24272,N_18462,N_18374);
nor U24273 (N_24273,N_22846,N_18633);
nor U24274 (N_24274,N_21309,N_21066);
and U24275 (N_24275,N_18429,N_20061);
nand U24276 (N_24276,N_19687,N_23405);
nor U24277 (N_24277,N_19603,N_19716);
xor U24278 (N_24278,N_18128,N_21674);
and U24279 (N_24279,N_20307,N_19278);
or U24280 (N_24280,N_18434,N_20660);
nand U24281 (N_24281,N_19771,N_23475);
nor U24282 (N_24282,N_19248,N_20564);
or U24283 (N_24283,N_21003,N_18755);
nand U24284 (N_24284,N_19808,N_21529);
xnor U24285 (N_24285,N_21148,N_23227);
nor U24286 (N_24286,N_20163,N_20212);
nand U24287 (N_24287,N_22648,N_19546);
and U24288 (N_24288,N_20527,N_22446);
and U24289 (N_24289,N_20796,N_23518);
or U24290 (N_24290,N_19690,N_22443);
nand U24291 (N_24291,N_21215,N_22350);
nand U24292 (N_24292,N_21442,N_18164);
or U24293 (N_24293,N_18320,N_23755);
xnor U24294 (N_24294,N_19964,N_22744);
nand U24295 (N_24295,N_22235,N_21448);
or U24296 (N_24296,N_21861,N_22913);
nor U24297 (N_24297,N_18795,N_23006);
or U24298 (N_24298,N_20252,N_20869);
or U24299 (N_24299,N_18686,N_19681);
xor U24300 (N_24300,N_18827,N_18074);
nand U24301 (N_24301,N_23764,N_21620);
xor U24302 (N_24302,N_23346,N_20777);
or U24303 (N_24303,N_18098,N_23174);
or U24304 (N_24304,N_20513,N_21172);
nor U24305 (N_24305,N_18287,N_19863);
or U24306 (N_24306,N_21160,N_18786);
nand U24307 (N_24307,N_20334,N_21263);
nor U24308 (N_24308,N_22270,N_19637);
nor U24309 (N_24309,N_22410,N_22988);
nor U24310 (N_24310,N_20626,N_22563);
or U24311 (N_24311,N_23357,N_18606);
and U24312 (N_24312,N_21927,N_19089);
nor U24313 (N_24313,N_19867,N_19268);
and U24314 (N_24314,N_23817,N_19017);
or U24315 (N_24315,N_20204,N_21319);
nor U24316 (N_24316,N_20721,N_20559);
nor U24317 (N_24317,N_23131,N_18992);
xor U24318 (N_24318,N_23861,N_23961);
and U24319 (N_24319,N_23244,N_18377);
nand U24320 (N_24320,N_22269,N_22059);
nand U24321 (N_24321,N_23614,N_22654);
nor U24322 (N_24322,N_19348,N_21849);
nor U24323 (N_24323,N_18549,N_20939);
and U24324 (N_24324,N_21325,N_20235);
nor U24325 (N_24325,N_18347,N_23902);
nand U24326 (N_24326,N_21536,N_19270);
nor U24327 (N_24327,N_23362,N_21531);
xnor U24328 (N_24328,N_18271,N_22661);
nor U24329 (N_24329,N_22841,N_23432);
and U24330 (N_24330,N_20821,N_22868);
and U24331 (N_24331,N_20827,N_18525);
nor U24332 (N_24332,N_18850,N_21578);
or U24333 (N_24333,N_18231,N_18519);
nor U24334 (N_24334,N_23368,N_22668);
nor U24335 (N_24335,N_20894,N_22187);
nor U24336 (N_24336,N_20872,N_21854);
or U24337 (N_24337,N_21025,N_23517);
nor U24338 (N_24338,N_18171,N_21735);
nor U24339 (N_24339,N_20967,N_22995);
nand U24340 (N_24340,N_21223,N_18861);
nor U24341 (N_24341,N_22839,N_21185);
nor U24342 (N_24342,N_23162,N_23249);
or U24343 (N_24343,N_21486,N_21783);
nor U24344 (N_24344,N_23274,N_18314);
or U24345 (N_24345,N_22624,N_22538);
nor U24346 (N_24346,N_19084,N_21230);
xnor U24347 (N_24347,N_20004,N_23954);
and U24348 (N_24348,N_18695,N_18404);
xnor U24349 (N_24349,N_20700,N_19038);
nand U24350 (N_24350,N_23893,N_20893);
nand U24351 (N_24351,N_22799,N_22904);
and U24352 (N_24352,N_20589,N_22646);
xnor U24353 (N_24353,N_23669,N_18728);
xor U24354 (N_24354,N_22070,N_23258);
or U24355 (N_24355,N_21946,N_19352);
and U24356 (N_24356,N_23880,N_19511);
xnor U24357 (N_24357,N_21288,N_18812);
nand U24358 (N_24358,N_21848,N_23077);
and U24359 (N_24359,N_19517,N_23461);
nor U24360 (N_24360,N_19157,N_23792);
nand U24361 (N_24361,N_23418,N_23648);
xnor U24362 (N_24362,N_23054,N_23373);
and U24363 (N_24363,N_19247,N_23711);
or U24364 (N_24364,N_22570,N_23177);
nand U24365 (N_24365,N_18465,N_21011);
nor U24366 (N_24366,N_18075,N_22261);
nor U24367 (N_24367,N_20682,N_22292);
nand U24368 (N_24368,N_18580,N_21453);
nand U24369 (N_24369,N_23851,N_19042);
or U24370 (N_24370,N_22971,N_21819);
and U24371 (N_24371,N_22166,N_18141);
xor U24372 (N_24372,N_21334,N_20962);
and U24373 (N_24373,N_19627,N_19086);
and U24374 (N_24374,N_20184,N_19918);
nor U24375 (N_24375,N_23169,N_21069);
or U24376 (N_24376,N_21119,N_20368);
nor U24377 (N_24377,N_22750,N_21451);
nor U24378 (N_24378,N_22759,N_21256);
xnor U24379 (N_24379,N_20729,N_19655);
xor U24380 (N_24380,N_22590,N_22878);
nand U24381 (N_24381,N_18651,N_18604);
nor U24382 (N_24382,N_22849,N_23526);
nor U24383 (N_24383,N_22892,N_19593);
xnor U24384 (N_24384,N_18150,N_18634);
nor U24385 (N_24385,N_22524,N_19823);
nor U24386 (N_24386,N_23264,N_23221);
xor U24387 (N_24387,N_21558,N_20398);
nand U24388 (N_24388,N_19521,N_21568);
or U24389 (N_24389,N_23644,N_21432);
xor U24390 (N_24390,N_21335,N_22004);
or U24391 (N_24391,N_22338,N_20707);
or U24392 (N_24392,N_23028,N_18522);
or U24393 (N_24393,N_20711,N_21043);
or U24394 (N_24394,N_21454,N_22905);
or U24395 (N_24395,N_21026,N_19925);
and U24396 (N_24396,N_18826,N_20049);
nor U24397 (N_24397,N_19923,N_19605);
or U24398 (N_24398,N_18904,N_23347);
nor U24399 (N_24399,N_19600,N_19555);
and U24400 (N_24400,N_18358,N_21712);
nand U24401 (N_24401,N_20704,N_18931);
and U24402 (N_24402,N_19775,N_21641);
nor U24403 (N_24403,N_23516,N_18124);
or U24404 (N_24404,N_19649,N_22356);
xor U24405 (N_24405,N_21610,N_21634);
nand U24406 (N_24406,N_18199,N_21818);
nor U24407 (N_24407,N_21065,N_19420);
or U24408 (N_24408,N_23543,N_22850);
xnor U24409 (N_24409,N_19415,N_18007);
nand U24410 (N_24410,N_20969,N_20845);
xnor U24411 (N_24411,N_21802,N_22399);
nor U24412 (N_24412,N_23993,N_19661);
nand U24413 (N_24413,N_22386,N_22689);
or U24414 (N_24414,N_21551,N_18276);
or U24415 (N_24415,N_21421,N_22738);
nor U24416 (N_24416,N_23429,N_18601);
nand U24417 (N_24417,N_23238,N_18249);
xnor U24418 (N_24418,N_19456,N_22579);
nand U24419 (N_24419,N_21840,N_23867);
and U24420 (N_24420,N_23291,N_20582);
xnor U24421 (N_24421,N_19890,N_23309);
or U24422 (N_24422,N_20524,N_20571);
nand U24423 (N_24423,N_22775,N_20782);
or U24424 (N_24424,N_18593,N_20487);
xor U24425 (N_24425,N_18491,N_21244);
xnor U24426 (N_24426,N_22510,N_18153);
nand U24427 (N_24427,N_21328,N_20820);
xnor U24428 (N_24428,N_20658,N_20239);
nor U24429 (N_24429,N_22990,N_20818);
nor U24430 (N_24430,N_20118,N_20987);
and U24431 (N_24431,N_19552,N_18273);
and U24432 (N_24432,N_21863,N_22315);
and U24433 (N_24433,N_18521,N_21817);
nand U24434 (N_24434,N_21571,N_20566);
and U24435 (N_24435,N_19108,N_21138);
xnor U24436 (N_24436,N_19512,N_23360);
nor U24437 (N_24437,N_22394,N_18706);
nor U24438 (N_24438,N_23538,N_22851);
and U24439 (N_24439,N_23850,N_22968);
or U24440 (N_24440,N_23170,N_23048);
xnor U24441 (N_24441,N_19894,N_21855);
xor U24442 (N_24442,N_20986,N_18117);
xor U24443 (N_24443,N_22768,N_21431);
or U24444 (N_24444,N_23126,N_22165);
xnor U24445 (N_24445,N_23513,N_22071);
and U24446 (N_24446,N_20795,N_22823);
and U24447 (N_24447,N_20862,N_18647);
nor U24448 (N_24448,N_23878,N_22871);
xnor U24449 (N_24449,N_20731,N_19791);
or U24450 (N_24450,N_22599,N_23779);
nand U24451 (N_24451,N_20678,N_23793);
or U24452 (N_24452,N_20580,N_22320);
or U24453 (N_24453,N_20147,N_21732);
or U24454 (N_24454,N_18031,N_21382);
or U24455 (N_24455,N_21458,N_22644);
xor U24456 (N_24456,N_18707,N_23289);
nand U24457 (N_24457,N_20488,N_18607);
xor U24458 (N_24458,N_23494,N_19214);
xnor U24459 (N_24459,N_21570,N_18770);
and U24460 (N_24460,N_19479,N_19114);
nor U24461 (N_24461,N_22899,N_19658);
nand U24462 (N_24462,N_22885,N_22925);
xor U24463 (N_24463,N_20276,N_23259);
or U24464 (N_24464,N_23603,N_19344);
and U24465 (N_24465,N_21941,N_22332);
and U24466 (N_24466,N_22103,N_20832);
nand U24467 (N_24467,N_21627,N_20654);
xor U24468 (N_24468,N_19779,N_20455);
xor U24469 (N_24469,N_23904,N_19169);
or U24470 (N_24470,N_19300,N_19001);
nor U24471 (N_24471,N_23102,N_22147);
or U24472 (N_24472,N_19093,N_22118);
xnor U24473 (N_24473,N_20937,N_23702);
nand U24474 (N_24474,N_19547,N_18645);
nor U24475 (N_24475,N_19732,N_20882);
nor U24476 (N_24476,N_22791,N_18758);
nor U24477 (N_24477,N_22940,N_21416);
nand U24478 (N_24478,N_23969,N_23771);
or U24479 (N_24479,N_18819,N_21218);
or U24480 (N_24480,N_19029,N_22647);
and U24481 (N_24481,N_20006,N_18715);
xnor U24482 (N_24482,N_23802,N_18917);
and U24483 (N_24483,N_19312,N_20446);
nor U24484 (N_24484,N_20040,N_21933);
xnor U24485 (N_24485,N_22142,N_22972);
nand U24486 (N_24486,N_18922,N_21015);
or U24487 (N_24487,N_23220,N_19738);
xnor U24488 (N_24488,N_18878,N_23774);
nor U24489 (N_24489,N_21575,N_19320);
nor U24490 (N_24490,N_18814,N_20743);
nand U24491 (N_24491,N_20860,N_21455);
xnor U24492 (N_24492,N_18749,N_22020);
nor U24493 (N_24493,N_23160,N_21704);
and U24494 (N_24494,N_20936,N_23288);
and U24495 (N_24495,N_23182,N_23416);
xnor U24496 (N_24496,N_21851,N_20030);
xnor U24497 (N_24497,N_22608,N_22778);
nand U24498 (N_24498,N_21067,N_19538);
xor U24499 (N_24499,N_22033,N_19019);
and U24500 (N_24500,N_23367,N_23942);
nor U24501 (N_24501,N_21708,N_18083);
or U24502 (N_24502,N_21823,N_22464);
or U24503 (N_24503,N_18516,N_20718);
xor U24504 (N_24504,N_18557,N_20975);
nor U24505 (N_24505,N_19910,N_22330);
and U24506 (N_24506,N_18090,N_22955);
xnor U24507 (N_24507,N_20778,N_23837);
xnor U24508 (N_24508,N_20054,N_19800);
xnor U24509 (N_24509,N_21826,N_20444);
or U24510 (N_24510,N_18559,N_21369);
xor U24511 (N_24511,N_19310,N_22244);
and U24512 (N_24512,N_22604,N_21904);
xnor U24513 (N_24513,N_20174,N_20573);
and U24514 (N_24514,N_21112,N_21886);
xor U24515 (N_24515,N_21332,N_18051);
and U24516 (N_24516,N_21093,N_22500);
nand U24517 (N_24517,N_22863,N_22785);
and U24518 (N_24518,N_23065,N_18334);
nor U24519 (N_24519,N_19328,N_18336);
xnor U24520 (N_24520,N_22130,N_23814);
nand U24521 (N_24521,N_22911,N_18963);
xnor U24522 (N_24522,N_21961,N_18730);
nor U24523 (N_24523,N_18229,N_19692);
xnor U24524 (N_24524,N_20520,N_22383);
nor U24525 (N_24525,N_19693,N_22535);
and U24526 (N_24526,N_21834,N_22757);
and U24527 (N_24527,N_22631,N_22681);
nand U24528 (N_24528,N_20310,N_20521);
nor U24529 (N_24529,N_18608,N_23763);
or U24530 (N_24530,N_23045,N_20753);
xor U24531 (N_24531,N_23673,N_23132);
nor U24532 (N_24532,N_23098,N_22694);
and U24533 (N_24533,N_19287,N_23011);
nor U24534 (N_24534,N_21175,N_19701);
nor U24535 (N_24535,N_18280,N_19070);
and U24536 (N_24536,N_23281,N_21616);
xnor U24537 (N_24537,N_19610,N_23846);
nor U24538 (N_24538,N_18473,N_20726);
xnor U24539 (N_24539,N_22076,N_23228);
nand U24540 (N_24540,N_20000,N_18077);
or U24541 (N_24541,N_21074,N_21343);
xor U24542 (N_24542,N_23671,N_22377);
xor U24543 (N_24543,N_22445,N_22660);
or U24544 (N_24544,N_21920,N_19500);
and U24545 (N_24545,N_18499,N_19551);
or U24546 (N_24546,N_21748,N_21829);
xnor U24547 (N_24547,N_19301,N_20496);
or U24548 (N_24548,N_19708,N_21806);
or U24549 (N_24549,N_23570,N_18823);
or U24550 (N_24550,N_21901,N_21685);
or U24551 (N_24551,N_22736,N_21078);
xnor U24552 (N_24552,N_21354,N_19030);
nor U24553 (N_24553,N_20280,N_20180);
xor U24554 (N_24554,N_23501,N_19548);
xnor U24555 (N_24555,N_20623,N_21365);
nor U24556 (N_24556,N_21556,N_22218);
and U24557 (N_24557,N_20690,N_22898);
or U24558 (N_24558,N_21740,N_21642);
xnor U24559 (N_24559,N_22369,N_19504);
or U24560 (N_24560,N_19912,N_20287);
nor U24561 (N_24561,N_21714,N_21598);
nand U24562 (N_24562,N_18029,N_21505);
or U24563 (N_24563,N_18912,N_19740);
or U24564 (N_24564,N_22561,N_19286);
nand U24565 (N_24565,N_23426,N_21579);
and U24566 (N_24566,N_18632,N_23713);
nand U24567 (N_24567,N_18673,N_22550);
nand U24568 (N_24568,N_18996,N_21133);
nand U24569 (N_24569,N_22806,N_19494);
or U24570 (N_24570,N_22587,N_21940);
or U24571 (N_24571,N_20679,N_20531);
nor U24572 (N_24572,N_20348,N_22440);
xnor U24573 (N_24573,N_19385,N_18241);
or U24574 (N_24574,N_19844,N_22172);
nor U24575 (N_24575,N_23971,N_19468);
nand U24576 (N_24576,N_19798,N_18524);
and U24577 (N_24577,N_21197,N_19145);
xor U24578 (N_24578,N_22400,N_23109);
xnor U24579 (N_24579,N_20545,N_20672);
xor U24580 (N_24580,N_19119,N_21528);
or U24581 (N_24581,N_22848,N_20491);
nor U24582 (N_24582,N_18591,N_19789);
xor U24583 (N_24583,N_21368,N_21587);
nor U24584 (N_24584,N_19702,N_19956);
xor U24585 (N_24585,N_23696,N_20022);
nor U24586 (N_24586,N_22122,N_18765);
or U24587 (N_24587,N_23964,N_21593);
or U24588 (N_24588,N_23600,N_18409);
and U24589 (N_24589,N_19390,N_19191);
nand U24590 (N_24590,N_20220,N_18338);
nand U24591 (N_24591,N_20069,N_20171);
xnor U24592 (N_24592,N_21733,N_21401);
nand U24593 (N_24593,N_21656,N_20955);
and U24594 (N_24594,N_23502,N_20089);
xor U24595 (N_24595,N_23284,N_18700);
xor U24596 (N_24596,N_19762,N_22678);
and U24597 (N_24597,N_22513,N_18274);
or U24598 (N_24598,N_23267,N_18178);
xnor U24599 (N_24599,N_23395,N_22937);
or U24600 (N_24600,N_18845,N_20576);
and U24601 (N_24601,N_19453,N_23746);
and U24602 (N_24602,N_19367,N_18513);
xor U24603 (N_24603,N_18445,N_21480);
and U24604 (N_24604,N_19854,N_20925);
or U24605 (N_24605,N_22233,N_22150);
xor U24606 (N_24606,N_20349,N_19813);
or U24607 (N_24607,N_19141,N_19897);
nor U24608 (N_24608,N_23021,N_20100);
and U24609 (N_24609,N_21418,N_22465);
xnor U24610 (N_24610,N_19049,N_19369);
nor U24611 (N_24611,N_20624,N_19467);
and U24612 (N_24612,N_22653,N_22705);
and U24613 (N_24613,N_23935,N_18109);
nand U24614 (N_24614,N_21136,N_18628);
nor U24615 (N_24615,N_23730,N_19678);
xnor U24616 (N_24616,N_18163,N_19233);
xnor U24617 (N_24617,N_19188,N_21669);
and U24618 (N_24618,N_18004,N_20094);
or U24619 (N_24619,N_23370,N_23737);
nor U24620 (N_24620,N_18517,N_22516);
or U24621 (N_24621,N_20382,N_21775);
and U24622 (N_24622,N_20553,N_19616);
xor U24623 (N_24623,N_22555,N_19837);
nand U24624 (N_24624,N_18255,N_19501);
and U24625 (N_24625,N_21673,N_19138);
and U24626 (N_24626,N_22016,N_23654);
nand U24627 (N_24627,N_20459,N_23148);
and U24628 (N_24628,N_18385,N_20665);
or U24629 (N_24629,N_20294,N_22025);
nor U24630 (N_24630,N_22962,N_18100);
nor U24631 (N_24631,N_21801,N_22886);
or U24632 (N_24632,N_21311,N_19485);
nor U24633 (N_24633,N_21844,N_20471);
xnor U24634 (N_24634,N_19862,N_19939);
or U24635 (N_24635,N_20701,N_19646);
and U24636 (N_24636,N_20523,N_18671);
or U24637 (N_24637,N_23085,N_21950);
and U24638 (N_24638,N_21449,N_20271);
and U24639 (N_24639,N_22406,N_21565);
xnor U24640 (N_24640,N_21314,N_22894);
nand U24641 (N_24641,N_22404,N_20592);
xor U24642 (N_24642,N_21895,N_23093);
nor U24643 (N_24643,N_22789,N_20360);
or U24644 (N_24644,N_23579,N_21315);
xnor U24645 (N_24645,N_22977,N_20799);
or U24646 (N_24646,N_18942,N_21367);
nor U24647 (N_24647,N_20112,N_18295);
and U24648 (N_24648,N_23991,N_21099);
and U24649 (N_24649,N_21777,N_19674);
nand U24650 (N_24650,N_23542,N_20328);
or U24651 (N_24651,N_20972,N_23747);
or U24652 (N_24652,N_21691,N_22651);
xnor U24653 (N_24653,N_22488,N_21773);
xnor U24654 (N_24654,N_22682,N_19944);
nand U24655 (N_24655,N_19158,N_20614);
nand U24656 (N_24656,N_19725,N_18583);
nand U24657 (N_24657,N_19356,N_22463);
xnor U24658 (N_24658,N_22127,N_20405);
or U24659 (N_24659,N_23273,N_19335);
and U24660 (N_24660,N_19744,N_21681);
xnor U24661 (N_24661,N_19933,N_21645);
nor U24662 (N_24662,N_23949,N_21980);
nand U24663 (N_24663,N_23789,N_23236);
or U24664 (N_24664,N_20149,N_19292);
nor U24665 (N_24665,N_19832,N_23180);
and U24666 (N_24666,N_21767,N_21323);
xnor U24667 (N_24667,N_18256,N_21171);
and U24668 (N_24668,N_22755,N_19773);
or U24669 (N_24669,N_19458,N_23431);
and U24670 (N_24670,N_19684,N_18760);
or U24671 (N_24671,N_21468,N_23096);
or U24672 (N_24672,N_21996,N_22415);
nand U24673 (N_24673,N_20312,N_23597);
and U24674 (N_24674,N_21731,N_22567);
nand U24675 (N_24675,N_18646,N_20724);
xnor U24676 (N_24676,N_19193,N_23975);
nor U24677 (N_24677,N_22558,N_21243);
nand U24678 (N_24678,N_22021,N_22961);
or U24679 (N_24679,N_22766,N_20847);
or U24680 (N_24680,N_23623,N_19513);
and U24681 (N_24681,N_23599,N_22546);
and U24682 (N_24682,N_19186,N_18641);
and U24683 (N_24683,N_20541,N_20416);
nand U24684 (N_24684,N_19414,N_19332);
nand U24685 (N_24685,N_20250,N_22929);
nor U24686 (N_24686,N_20086,N_23743);
or U24687 (N_24687,N_18348,N_22984);
and U24688 (N_24688,N_18089,N_20139);
nor U24689 (N_24689,N_23912,N_22728);
nand U24690 (N_24690,N_18272,N_19571);
nor U24691 (N_24691,N_19146,N_20669);
or U24692 (N_24692,N_19722,N_19893);
nand U24693 (N_24693,N_22853,N_23984);
nand U24694 (N_24694,N_23142,N_19116);
or U24695 (N_24695,N_20422,N_20044);
nand U24696 (N_24696,N_22649,N_18757);
nor U24697 (N_24697,N_21338,N_19282);
and U24698 (N_24698,N_23459,N_18805);
nand U24699 (N_24699,N_20336,N_23171);
nand U24700 (N_24700,N_20984,N_20189);
or U24701 (N_24701,N_23499,N_21377);
xnor U24702 (N_24702,N_23722,N_20232);
xor U24703 (N_24703,N_22047,N_23216);
nand U24704 (N_24704,N_20958,N_18612);
and U24705 (N_24705,N_21688,N_18742);
nor U24706 (N_24706,N_22264,N_21652);
and U24707 (N_24707,N_22478,N_22451);
nor U24708 (N_24708,N_18159,N_20699);
nor U24709 (N_24709,N_21502,N_23914);
nor U24710 (N_24710,N_20608,N_20657);
xnor U24711 (N_24711,N_18353,N_19032);
nand U24712 (N_24712,N_23831,N_22748);
nand U24713 (N_24713,N_22030,N_23498);
nand U24714 (N_24714,N_23064,N_21890);
nor U24715 (N_24715,N_23013,N_21824);
nor U24716 (N_24716,N_19572,N_18431);
nand U24717 (N_24717,N_19679,N_20478);
and U24718 (N_24718,N_20995,N_23652);
or U24719 (N_24719,N_19958,N_19983);
nor U24720 (N_24720,N_21566,N_20321);
or U24721 (N_24721,N_20507,N_18866);
or U24722 (N_24722,N_20203,N_21202);
nand U24723 (N_24723,N_20656,N_20485);
nand U24724 (N_24724,N_19000,N_18855);
xor U24725 (N_24725,N_20855,N_19936);
and U24726 (N_24726,N_19363,N_23534);
nor U24727 (N_24727,N_21438,N_22284);
xnor U24728 (N_24728,N_22407,N_20708);
nor U24729 (N_24729,N_22114,N_18481);
and U24730 (N_24730,N_20002,N_23891);
xnor U24731 (N_24731,N_23847,N_18660);
xor U24732 (N_24732,N_19509,N_22434);
and U24733 (N_24733,N_18078,N_18656);
nand U24734 (N_24734,N_19794,N_18568);
xnor U24735 (N_24735,N_18122,N_23787);
or U24736 (N_24736,N_22636,N_19845);
nand U24737 (N_24737,N_20948,N_21153);
nand U24738 (N_24738,N_23137,N_21182);
and U24739 (N_24739,N_19705,N_21525);
xor U24740 (N_24740,N_21333,N_23253);
nand U24741 (N_24741,N_18894,N_18851);
xor U24742 (N_24742,N_19528,N_19885);
or U24743 (N_24743,N_23877,N_18279);
nand U24744 (N_24744,N_21719,N_19612);
nand U24745 (N_24745,N_22829,N_19088);
nor U24746 (N_24746,N_23198,N_21663);
nand U24747 (N_24747,N_20610,N_20090);
and U24748 (N_24748,N_22007,N_20104);
nor U24749 (N_24749,N_21270,N_18903);
nand U24750 (N_24750,N_19560,N_18927);
and U24751 (N_24751,N_19776,N_18102);
xnor U24752 (N_24752,N_22462,N_20912);
nand U24753 (N_24753,N_19633,N_19626);
nor U24754 (N_24754,N_18328,N_21532);
nor U24755 (N_24755,N_22994,N_18149);
nor U24756 (N_24756,N_21743,N_20247);
xnor U24757 (N_24757,N_18945,N_21664);
nand U24758 (N_24758,N_21109,N_20025);
xor U24759 (N_24759,N_23910,N_21956);
or U24760 (N_24760,N_20286,N_19520);
or U24761 (N_24761,N_20558,N_18598);
nor U24762 (N_24762,N_18011,N_20469);
nand U24763 (N_24763,N_18869,N_23608);
and U24764 (N_24764,N_22723,N_18959);
or U24765 (N_24765,N_23113,N_19408);
or U24766 (N_24766,N_19686,N_23478);
nand U24767 (N_24767,N_21059,N_21543);
xnor U24768 (N_24768,N_18307,N_23403);
xnor U24769 (N_24769,N_21928,N_21476);
and U24770 (N_24770,N_22712,N_18908);
nand U24771 (N_24771,N_19156,N_20663);
nand U24772 (N_24772,N_21352,N_22754);
nand U24773 (N_24773,N_19412,N_22876);
xnor U24774 (N_24774,N_18972,N_22870);
or U24775 (N_24775,N_21413,N_22600);
nand U24776 (N_24776,N_23855,N_20638);
or U24777 (N_24777,N_23797,N_22964);
or U24778 (N_24778,N_18412,N_20709);
nand U24779 (N_24779,N_18834,N_19594);
or U24780 (N_24780,N_18166,N_18183);
and U24781 (N_24781,N_22864,N_19785);
nor U24782 (N_24782,N_18971,N_18173);
and U24783 (N_24783,N_22137,N_20785);
xor U24784 (N_24784,N_18863,N_19527);
or U24785 (N_24785,N_22975,N_20135);
or U24786 (N_24786,N_18458,N_21484);
xnor U24787 (N_24787,N_23397,N_18346);
nand U24788 (N_24788,N_18979,N_19200);
xnor U24789 (N_24789,N_22098,N_18138);
xor U24790 (N_24790,N_18547,N_19452);
nor U24791 (N_24791,N_23677,N_19628);
or U24792 (N_24792,N_20099,N_23750);
or U24793 (N_24793,N_19596,N_18046);
nor U24794 (N_24794,N_18788,N_18733);
xor U24795 (N_24795,N_21144,N_19739);
nand U24796 (N_24796,N_20363,N_22693);
and U24797 (N_24797,N_23869,N_22327);
nand U24798 (N_24798,N_19843,N_20935);
xnor U24799 (N_24799,N_20953,N_22306);
or U24800 (N_24800,N_21675,N_21013);
and U24801 (N_24801,N_19653,N_18678);
or U24802 (N_24802,N_19999,N_18662);
or U24803 (N_24803,N_19115,N_20063);
or U24804 (N_24804,N_21971,N_23477);
xor U24805 (N_24805,N_18364,N_23901);
nand U24806 (N_24806,N_18918,N_19241);
nand U24807 (N_24807,N_18416,N_19841);
and U24808 (N_24808,N_18493,N_23799);
xnor U24809 (N_24809,N_23528,N_22200);
nand U24810 (N_24810,N_18808,N_21152);
or U24811 (N_24811,N_21140,N_23525);
nor U24812 (N_24812,N_21183,N_18862);
nand U24813 (N_24813,N_18915,N_21117);
nand U24814 (N_24814,N_23633,N_21228);
xor U24815 (N_24815,N_23252,N_21524);
xor U24816 (N_24816,N_23401,N_20460);
nand U24817 (N_24817,N_18201,N_22131);
and U24818 (N_24818,N_23222,N_22701);
and U24819 (N_24819,N_22135,N_18966);
or U24820 (N_24820,N_20532,N_20224);
nand U24821 (N_24821,N_18816,N_20065);
or U24822 (N_24822,N_18876,N_23121);
or U24823 (N_24823,N_21870,N_22243);
nand U24824 (N_24824,N_20915,N_20631);
or U24825 (N_24825,N_19256,N_23794);
xnor U24826 (N_24826,N_23400,N_20952);
xnor U24827 (N_24827,N_18013,N_23858);
nand U24828 (N_24828,N_21345,N_22210);
nand U24829 (N_24829,N_23996,N_20877);
or U24830 (N_24830,N_22674,N_20001);
and U24831 (N_24831,N_18731,N_22735);
nand U24832 (N_24832,N_20053,N_19916);
xor U24833 (N_24833,N_22797,N_18433);
nand U24834 (N_24834,N_18571,N_20629);
nor U24835 (N_24835,N_18676,N_23752);
nand U24836 (N_24836,N_18560,N_21544);
or U24837 (N_24837,N_23906,N_22436);
nand U24838 (N_24838,N_22773,N_22454);
and U24839 (N_24839,N_19275,N_21722);
nor U24840 (N_24840,N_18033,N_22487);
or U24841 (N_24841,N_19997,N_23153);
nand U24842 (N_24842,N_19382,N_19360);
nor U24843 (N_24843,N_18774,N_21494);
or U24844 (N_24844,N_23047,N_19222);
and U24845 (N_24845,N_19008,N_20841);
and U24846 (N_24846,N_20773,N_18653);
and U24847 (N_24847,N_19166,N_21676);
xnor U24848 (N_24848,N_23974,N_19907);
nand U24849 (N_24849,N_19950,N_18950);
xor U24850 (N_24850,N_23262,N_18297);
nor U24851 (N_24851,N_19216,N_19267);
xor U24852 (N_24852,N_20583,N_22520);
nand U24853 (N_24853,N_23832,N_20501);
or U24854 (N_24854,N_23510,N_21161);
and U24855 (N_24855,N_18094,N_20586);
xnor U24856 (N_24856,N_19720,N_20461);
and U24857 (N_24857,N_20585,N_22043);
nand U24858 (N_24858,N_18370,N_22080);
or U24859 (N_24859,N_21597,N_18107);
and U24860 (N_24860,N_19297,N_18323);
nor U24861 (N_24861,N_22449,N_22733);
xor U24862 (N_24862,N_21005,N_19793);
nor U24863 (N_24863,N_23734,N_21101);
and U24864 (N_24864,N_21955,N_18463);
nor U24865 (N_24865,N_22522,N_23297);
xor U24866 (N_24866,N_18248,N_21293);
xnor U24867 (N_24867,N_23039,N_19664);
nand U24868 (N_24868,N_19239,N_23385);
nand U24869 (N_24869,N_23161,N_23445);
and U24870 (N_24870,N_22034,N_19758);
or U24871 (N_24871,N_23191,N_21415);
nor U24872 (N_24872,N_23492,N_21020);
xnor U24873 (N_24873,N_21530,N_23410);
or U24874 (N_24874,N_19949,N_20871);
and U24875 (N_24875,N_19113,N_19445);
nor U24876 (N_24876,N_18603,N_23592);
and U24877 (N_24877,N_21770,N_22676);
or U24878 (N_24878,N_23626,N_20429);
and U24879 (N_24879,N_19957,N_20108);
nand U24880 (N_24880,N_21727,N_21868);
nor U24881 (N_24881,N_18285,N_21647);
nor U24882 (N_24882,N_23960,N_22256);
nor U24883 (N_24883,N_23757,N_22333);
xnor U24884 (N_24884,N_19711,N_21812);
nor U24885 (N_24885,N_23331,N_23208);
and U24886 (N_24886,N_18344,N_19148);
nand U24887 (N_24887,N_20511,N_22063);
or U24888 (N_24888,N_18384,N_18746);
xor U24889 (N_24889,N_21595,N_19243);
and U24890 (N_24890,N_19905,N_18451);
xor U24891 (N_24891,N_20256,N_18125);
and U24892 (N_24892,N_19481,N_20644);
nand U24893 (N_24893,N_22086,N_21986);
xnor U24894 (N_24894,N_19755,N_18470);
and U24895 (N_24895,N_19026,N_21307);
or U24896 (N_24896,N_22403,N_19081);
or U24897 (N_24897,N_22157,N_22069);
nor U24898 (N_24898,N_19715,N_20892);
and U24899 (N_24899,N_18382,N_23759);
nand U24900 (N_24900,N_19334,N_18309);
nand U24901 (N_24901,N_21024,N_22673);
xnor U24902 (N_24902,N_22387,N_21887);
or U24903 (N_24903,N_18196,N_19212);
and U24904 (N_24904,N_21405,N_21874);
nor U24905 (N_24905,N_21810,N_22123);
nor U24906 (N_24906,N_19754,N_20950);
nand U24907 (N_24907,N_19266,N_23352);
xnor U24908 (N_24908,N_18072,N_22433);
or U24909 (N_24909,N_18084,N_18887);
or U24910 (N_24910,N_20324,N_19132);
and U24911 (N_24911,N_23613,N_19491);
nor U24912 (N_24912,N_20842,N_23008);
or U24913 (N_24913,N_18847,N_20395);
or U24914 (N_24914,N_20142,N_23235);
nand U24915 (N_24915,N_20843,N_21761);
xor U24916 (N_24916,N_19695,N_22814);
xnor U24917 (N_24917,N_23803,N_18162);
or U24918 (N_24918,N_18430,N_22732);
nor U24919 (N_24919,N_21774,N_20677);
nand U24920 (N_24920,N_20924,N_21184);
xor U24921 (N_24921,N_22050,N_22731);
or U24922 (N_24922,N_21118,N_20440);
or U24923 (N_24923,N_23540,N_20265);
nand U24924 (N_24924,N_19488,N_19790);
xor U24925 (N_24925,N_20024,N_22238);
or U24926 (N_24926,N_18447,N_23094);
nand U24927 (N_24927,N_19037,N_19683);
or U24928 (N_24928,N_23932,N_18319);
xor U24929 (N_24929,N_20676,N_20738);
nand U24930 (N_24930,N_22708,N_18215);
and U24931 (N_24931,N_19309,N_19254);
or U24932 (N_24932,N_23727,N_22714);
and U24933 (N_24933,N_20362,N_23084);
or U24934 (N_24934,N_20436,N_18087);
or U24935 (N_24935,N_18650,N_21370);
xnor U24936 (N_24936,N_20430,N_20803);
nor U24937 (N_24937,N_20169,N_21785);
nor U24938 (N_24938,N_22344,N_21298);
nand U24939 (N_24939,N_18349,N_20674);
and U24940 (N_24940,N_18459,N_19745);
or U24941 (N_24941,N_20214,N_22417);
nand U24942 (N_24942,N_22052,N_19318);
or U24943 (N_24943,N_19036,N_23469);
xor U24944 (N_24944,N_18738,N_21277);
nor U24945 (N_24945,N_21924,N_20156);
and U24946 (N_24946,N_18000,N_18403);
nor U24947 (N_24947,N_23541,N_18674);
or U24948 (N_24948,N_21771,N_21504);
or U24949 (N_24949,N_21301,N_18485);
or U24950 (N_24950,N_21304,N_21222);
or U24951 (N_24951,N_23462,N_19974);
nor U24952 (N_24952,N_20233,N_23195);
and U24953 (N_24953,N_21520,N_21717);
nor U24954 (N_24954,N_19807,N_23655);
or U24955 (N_24955,N_18811,N_23602);
nand U24956 (N_24956,N_21252,N_21495);
xor U24957 (N_24957,N_20071,N_23452);
xnor U24958 (N_24958,N_22361,N_23396);
nor U24959 (N_24959,N_21670,N_18437);
and U24960 (N_24960,N_22439,N_19449);
xnor U24961 (N_24961,N_20739,N_20765);
nor U24962 (N_24962,N_22336,N_20850);
nor U24963 (N_24963,N_21657,N_20901);
and U24964 (N_24964,N_19237,N_21380);
nor U24965 (N_24965,N_18873,N_23256);
and U24966 (N_24966,N_18322,N_20667);
xor U24967 (N_24967,N_19225,N_19209);
nor U24968 (N_24968,N_21167,N_23196);
or U24969 (N_24969,N_21926,N_21693);
xnor U24970 (N_24970,N_20066,N_19694);
or U24971 (N_24971,N_21856,N_20477);
and U24972 (N_24972,N_21629,N_20081);
nand U24973 (N_24973,N_20996,N_19210);
xnor U24974 (N_24974,N_20415,N_19853);
xnor U24975 (N_24975,N_19872,N_20113);
xor U24976 (N_24976,N_23665,N_20769);
xnor U24977 (N_24977,N_23887,N_18635);
and U24978 (N_24978,N_19103,N_23807);
nand U24979 (N_24979,N_19358,N_22949);
xnor U24980 (N_24980,N_22553,N_23230);
xnor U24981 (N_24981,N_20505,N_20555);
nor U24982 (N_24982,N_19565,N_19476);
nand U24983 (N_24983,N_21385,N_18895);
nor U24984 (N_24984,N_23990,N_21150);
nor U24985 (N_24985,N_18408,N_23027);
nor U24986 (N_24986,N_18703,N_23316);
xnor U24987 (N_24987,N_19073,N_22777);
nand U24988 (N_24988,N_20019,N_19662);
and U24989 (N_24989,N_23795,N_21056);
and U24990 (N_24990,N_18567,N_22562);
xnor U24991 (N_24991,N_18363,N_23172);
nor U24992 (N_24992,N_21631,N_18802);
nor U24993 (N_24993,N_19938,N_22483);
nor U24994 (N_24994,N_22826,N_18930);
nand U24995 (N_24995,N_21051,N_19127);
xor U24996 (N_24996,N_21752,N_18672);
and U24997 (N_24997,N_19850,N_21427);
nor U24998 (N_24998,N_19035,N_19472);
nand U24999 (N_24999,N_23892,N_19322);
nand U25000 (N_25000,N_22902,N_20274);
xnor U25001 (N_25001,N_20900,N_21533);
or U25002 (N_25002,N_21795,N_20092);
xnor U25003 (N_25003,N_23183,N_22120);
nand U25004 (N_25004,N_19180,N_18157);
and U25005 (N_25005,N_21383,N_19522);
nand U25006 (N_25006,N_19112,N_18569);
and U25007 (N_25007,N_19881,N_19102);
or U25008 (N_25008,N_20880,N_20988);
nor U25009 (N_25009,N_20273,N_18367);
nor U25010 (N_25010,N_21998,N_22328);
or U25011 (N_25011,N_20284,N_19273);
and U25012 (N_25012,N_21224,N_22573);
nand U25013 (N_25013,N_18060,N_21021);
or U25014 (N_25014,N_20451,N_22266);
nor U25015 (N_25015,N_23242,N_22584);
or U25016 (N_25016,N_23037,N_18753);
xnor U25017 (N_25017,N_21033,N_22305);
nor U25018 (N_25018,N_20035,N_19747);
and U25019 (N_25019,N_20309,N_22657);
or U25020 (N_25020,N_21281,N_21825);
and U25021 (N_25021,N_21651,N_22634);
nor U25022 (N_25022,N_19982,N_22448);
and U25023 (N_25023,N_21273,N_18986);
and U25024 (N_25024,N_21091,N_19953);
and U25025 (N_25025,N_23186,N_23023);
and U25026 (N_25026,N_18584,N_22756);
and U25027 (N_25027,N_23857,N_23943);
nor U25028 (N_25028,N_23726,N_21879);
or U25029 (N_25029,N_19995,N_20418);
xnor U25030 (N_25030,N_20812,N_22471);
nor U25031 (N_25031,N_22626,N_22834);
or U25032 (N_25032,N_23456,N_19543);
or U25033 (N_25033,N_20551,N_19556);
nor U25034 (N_25034,N_20993,N_20130);
nand U25035 (N_25035,N_20257,N_21331);
and U25036 (N_25036,N_18234,N_20366);
nand U25037 (N_25037,N_22873,N_20680);
or U25038 (N_25038,N_20133,N_18217);
and U25039 (N_25039,N_21209,N_20062);
xnor U25040 (N_25040,N_19228,N_23555);
and U25041 (N_25041,N_20167,N_23883);
and U25042 (N_25042,N_23338,N_21507);
xnor U25043 (N_25043,N_19892,N_19861);
nand U25044 (N_25044,N_22236,N_23839);
xnor U25045 (N_25045,N_20182,N_19688);
nor U25046 (N_25046,N_22543,N_20941);
and U25047 (N_25047,N_22285,N_21177);
or U25048 (N_25048,N_18190,N_22959);
or U25049 (N_25049,N_21892,N_22659);
and U25050 (N_25050,N_21703,N_19417);
xnor U25051 (N_25051,N_18244,N_20752);
nor U25052 (N_25052,N_20313,N_18366);
or U25053 (N_25053,N_20762,N_18419);
nor U25054 (N_25054,N_21061,N_18467);
nand U25055 (N_25055,N_20494,N_20693);
nand U25056 (N_25056,N_18417,N_19575);
xor U25057 (N_25057,N_23896,N_19333);
and U25058 (N_25058,N_19183,N_19640);
xor U25059 (N_25059,N_18888,N_21866);
or U25060 (N_25060,N_23742,N_22335);
or U25061 (N_25061,N_19359,N_20043);
nor U25062 (N_25062,N_21724,N_21794);
or U25063 (N_25063,N_23650,N_18204);
xor U25064 (N_25064,N_22979,N_22620);
or U25065 (N_25065,N_23578,N_23411);
nor U25066 (N_25066,N_20578,N_21363);
xnor U25067 (N_25067,N_19343,N_23417);
nor U25068 (N_25068,N_19561,N_18565);
xnor U25069 (N_25069,N_23576,N_19377);
nand U25070 (N_25070,N_19051,N_23318);
or U25071 (N_25071,N_21408,N_22912);
nor U25072 (N_25072,N_18994,N_21984);
nand U25073 (N_25073,N_21027,N_20045);
nor U25074 (N_25074,N_22254,N_20807);
nand U25075 (N_25075,N_22276,N_18902);
nand U25076 (N_25076,N_23561,N_18085);
and U25077 (N_25077,N_19516,N_23970);
nor U25078 (N_25078,N_23785,N_21554);
nand U25079 (N_25079,N_21537,N_19591);
xor U25080 (N_25080,N_19615,N_19579);
nand U25081 (N_25081,N_19803,N_18865);
nand U25082 (N_25082,N_19652,N_20687);
xnor U25083 (N_25083,N_21220,N_22993);
nand U25084 (N_25084,N_23681,N_22616);
nor U25085 (N_25085,N_20162,N_23736);
and U25086 (N_25086,N_22384,N_18780);
xor U25087 (N_25087,N_20789,N_18511);
nor U25088 (N_25088,N_19345,N_18424);
nand U25089 (N_25089,N_19588,N_22275);
and U25090 (N_25090,N_22452,N_21113);
xnor U25091 (N_25091,N_22239,N_18235);
nand U25092 (N_25092,N_19710,N_22211);
or U25093 (N_25093,N_19518,N_20931);
or U25094 (N_25094,N_23381,N_21217);
and U25095 (N_25095,N_18946,N_19659);
or U25096 (N_25096,N_18211,N_23948);
nor U25097 (N_25097,N_20437,N_21267);
nand U25098 (N_25098,N_18722,N_20126);
nand U25099 (N_25099,N_20150,N_19041);
nand U25100 (N_25100,N_19418,N_22536);
and U25101 (N_25101,N_18003,N_19224);
and U25102 (N_25102,N_20628,N_18617);
or U25103 (N_25103,N_23097,N_20352);
or U25104 (N_25104,N_23886,N_23472);
nor U25105 (N_25105,N_19429,N_20728);
or U25106 (N_25106,N_22787,N_18251);
or U25107 (N_25107,N_18573,N_22402);
and U25108 (N_25108,N_20074,N_23280);
nor U25109 (N_25109,N_22193,N_21747);
xnor U25110 (N_25110,N_21017,N_21807);
nor U25111 (N_25111,N_21523,N_23767);
xor U25112 (N_25112,N_18984,N_19645);
nand U25113 (N_25113,N_18563,N_22314);
nor U25114 (N_25114,N_18055,N_23163);
xnor U25115 (N_25115,N_23263,N_22342);
and U25116 (N_25116,N_22725,N_22564);
nor U25117 (N_25117,N_23888,N_20026);
or U25118 (N_25118,N_18188,N_23674);
or U25119 (N_25119,N_21226,N_21010);
nor U25120 (N_25120,N_18218,N_21718);
and U25121 (N_25121,N_20664,N_22160);
or U25122 (N_25122,N_22408,N_23841);
or U25123 (N_25123,N_19650,N_20245);
nand U25124 (N_25124,N_22958,N_21538);
nor U25125 (N_25125,N_18308,N_20020);
nand U25126 (N_25126,N_20270,N_20170);
nor U25127 (N_25127,N_23741,N_18825);
nand U25128 (N_25128,N_18021,N_21398);
and U25129 (N_25129,N_21114,N_21212);
nand U25130 (N_25130,N_18352,N_23819);
nor U25131 (N_25131,N_19477,N_18014);
nor U25132 (N_25132,N_22241,N_23712);
nand U25133 (N_25133,N_22760,N_18677);
xnor U25134 (N_25134,N_19235,N_23205);
xor U25135 (N_25135,N_18527,N_23820);
nand U25136 (N_25136,N_18426,N_22316);
or U25137 (N_25137,N_19994,N_23840);
or U25138 (N_25138,N_21725,N_23188);
and U25139 (N_25139,N_18667,N_22710);
nor U25140 (N_25140,N_19562,N_18586);
nand U25141 (N_25141,N_20764,N_23962);
or U25142 (N_25142,N_21478,N_21373);
nand U25143 (N_25143,N_18800,N_21780);
xnor U25144 (N_25144,N_23050,N_19942);
and U25145 (N_25145,N_21582,N_21753);
or U25146 (N_25146,N_22595,N_19399);
nor U25147 (N_25147,N_19632,N_18127);
xnor U25148 (N_25148,N_20051,N_19712);
xnor U25149 (N_25149,N_20691,N_21911);
and U25150 (N_25150,N_21203,N_21973);
nor U25151 (N_25151,N_18503,N_18572);
xnor U25152 (N_25152,N_21330,N_20903);
or U25153 (N_25153,N_22421,N_22019);
nand U25154 (N_25154,N_19590,N_19279);
xor U25155 (N_25155,N_23029,N_19742);
and U25156 (N_25156,N_20359,N_21391);
xor U25157 (N_25157,N_23204,N_22621);
and U25158 (N_25158,N_21687,N_20497);
nor U25159 (N_25159,N_21690,N_18182);
nor U25160 (N_25160,N_23138,N_21846);
xor U25161 (N_25161,N_23091,N_21983);
nor U25162 (N_25162,N_20616,N_18882);
or U25163 (N_25163,N_22569,N_18682);
and U25164 (N_25164,N_19276,N_19595);
nor U25165 (N_25165,N_19155,N_21219);
and U25166 (N_25166,N_18691,N_20355);
nor U25167 (N_25167,N_19168,N_18028);
or U25168 (N_25168,N_23386,N_19532);
xnor U25169 (N_25169,N_21240,N_18399);
and U25170 (N_25170,N_19340,N_20300);
or U25171 (N_25171,N_18391,N_18174);
nor U25172 (N_25172,N_18529,N_19533);
and U25173 (N_25173,N_23327,N_19384);
or U25174 (N_25174,N_23224,N_18192);
or U25175 (N_25175,N_21186,N_21269);
and U25176 (N_25176,N_23783,N_21992);
and U25177 (N_25177,N_20712,N_19799);
and U25178 (N_25178,N_22192,N_20406);
nor U25179 (N_25179,N_20292,N_21179);
nand U25180 (N_25180,N_20630,N_22005);
or U25181 (N_25181,N_19900,N_23856);
and U25182 (N_25182,N_23465,N_21916);
nor U25183 (N_25183,N_19120,N_22924);
nor U25184 (N_25184,N_19602,N_20356);
nand U25185 (N_25185,N_22190,N_20954);
nor U25186 (N_25186,N_23881,N_23234);
and U25187 (N_25187,N_18652,N_18193);
xnor U25188 (N_25188,N_22890,N_20909);
xnor U25189 (N_25189,N_21087,N_19391);
xor U25190 (N_25190,N_21336,N_20528);
nor U25191 (N_25191,N_23788,N_19091);
nor U25192 (N_25192,N_18303,N_23120);
nand U25193 (N_25193,N_23639,N_22617);
or U25194 (N_25194,N_22058,N_21540);
nor U25195 (N_25195,N_19879,N_18520);
nand U25196 (N_25196,N_20384,N_19838);
nor U25197 (N_25197,N_21436,N_20538);
or U25198 (N_25198,N_21000,N_20262);
or U25199 (N_25199,N_19096,N_23640);
nor U25200 (N_25200,N_21337,N_19167);
and U25201 (N_25201,N_23953,N_19471);
and U25202 (N_25202,N_23958,N_21913);
and U25203 (N_25203,N_23824,N_19355);
and U25204 (N_25204,N_23907,N_20849);
or U25205 (N_25205,N_18947,N_18969);
xnor U25206 (N_25206,N_19707,N_20401);
nor U25207 (N_25207,N_23176,N_23521);
xor U25208 (N_25208,N_22861,N_18558);
xnor U25209 (N_25209,N_22642,N_19197);
nor U25210 (N_25210,N_22227,N_21292);
and U25211 (N_25211,N_22669,N_19441);
nor U25212 (N_25212,N_23553,N_18982);
or U25213 (N_25213,N_20605,N_21090);
or U25214 (N_25214,N_21769,N_21294);
xnor U25215 (N_25215,N_23676,N_22115);
and U25216 (N_25216,N_20875,N_20705);
nand U25217 (N_25217,N_22334,N_18212);
or U25218 (N_25218,N_18880,N_21546);
nand U25219 (N_25219,N_22088,N_23330);
xnor U25220 (N_25220,N_19817,N_20715);
or U25221 (N_25221,N_18246,N_21439);
nand U25222 (N_25222,N_18605,N_21545);
nand U25223 (N_25223,N_22637,N_20976);
xnor U25224 (N_25224,N_23693,N_19786);
and U25225 (N_25225,N_19766,N_19945);
xnor U25226 (N_25226,N_20870,N_23406);
nor U25227 (N_25227,N_18575,N_21750);
nand U25228 (N_25228,N_18389,N_20007);
nor U25229 (N_25229,N_18460,N_23615);
nand U25230 (N_25230,N_19375,N_18371);
xnor U25231 (N_25231,N_19311,N_20295);
xor U25232 (N_25232,N_22042,N_23341);
or U25233 (N_25233,N_19496,N_18350);
xnor U25234 (N_25234,N_21057,N_18830);
and U25235 (N_25235,N_21567,N_18397);
nand U25236 (N_25236,N_18809,N_19976);
nand U25237 (N_25237,N_22155,N_18796);
nand U25238 (N_25238,N_23628,N_22475);
and U25239 (N_25239,N_19034,N_22167);
nand U25240 (N_25240,N_21850,N_23476);
xor U25241 (N_25241,N_23125,N_18284);
or U25242 (N_25242,N_18073,N_22810);
nand U25243 (N_25243,N_22091,N_20335);
and U25244 (N_25244,N_22368,N_22168);
and U25245 (N_25245,N_20205,N_19641);
nand U25246 (N_25246,N_22015,N_21279);
nand U25247 (N_25247,N_21796,N_20347);
and U25248 (N_25248,N_18657,N_21500);
and U25249 (N_25249,N_20928,N_21729);
and U25250 (N_25250,N_22481,N_23591);
nor U25251 (N_25251,N_21599,N_20817);
xor U25252 (N_25252,N_19927,N_21508);
and U25253 (N_25253,N_19915,N_22039);
xor U25254 (N_25254,N_21910,N_19726);
or U25255 (N_25255,N_23939,N_19002);
or U25256 (N_25256,N_18870,N_22581);
and U25257 (N_25257,N_21374,N_23697);
nor U25258 (N_25258,N_21387,N_22245);
and U25259 (N_25259,N_21465,N_21744);
and U25260 (N_25260,N_18639,N_20502);
nor U25261 (N_25261,N_20942,N_22313);
xnor U25262 (N_25262,N_18679,N_22875);
or U25263 (N_25263,N_22656,N_22534);
and U25264 (N_25264,N_23678,N_18619);
nor U25265 (N_25265,N_20136,N_23729);
nand U25266 (N_25266,N_20052,N_18042);
xor U25267 (N_25267,N_18213,N_23556);
and U25268 (N_25268,N_19618,N_22828);
nor U25269 (N_25269,N_22973,N_19258);
xnor U25270 (N_25270,N_20651,N_23141);
xnor U25271 (N_25271,N_22782,N_21233);
and U25272 (N_25272,N_21860,N_21419);
xor U25273 (N_25273,N_21353,N_18666);
xor U25274 (N_25274,N_19987,N_20627);
xnor U25275 (N_25275,N_21459,N_21471);
or U25276 (N_25276,N_21805,N_19475);
and U25277 (N_25277,N_18263,N_19221);
xor U25278 (N_25278,N_21617,N_21407);
nor U25279 (N_25279,N_18658,N_23981);
nor U25280 (N_25280,N_23001,N_21351);
or U25281 (N_25281,N_20176,N_19361);
xnor U25282 (N_25282,N_22178,N_22698);
and U25283 (N_25283,N_22963,N_20070);
nor U25284 (N_25284,N_22683,N_20927);
xnor U25285 (N_25285,N_23862,N_18487);
and U25286 (N_25286,N_23966,N_18993);
nand U25287 (N_25287,N_18446,N_21800);
or U25288 (N_25288,N_21573,N_18877);
or U25289 (N_25289,N_23936,N_18243);
xnor U25290 (N_25290,N_18114,N_19930);
or U25291 (N_25291,N_18578,N_23283);
or U25292 (N_25292,N_22301,N_19011);
xor U25293 (N_25293,N_19137,N_18478);
and U25294 (N_25294,N_21004,N_20518);
nand U25295 (N_25295,N_19069,N_20048);
or U25296 (N_25296,N_19440,N_19911);
xnor U25297 (N_25297,N_18928,N_19271);
xor U25298 (N_25298,N_20047,N_21899);
and U25299 (N_25299,N_22081,N_20140);
nand U25300 (N_25300,N_22671,N_23486);
nor U25301 (N_25301,N_22960,N_23664);
or U25302 (N_25302,N_22552,N_23268);
xor U25303 (N_25303,N_19589,N_23087);
nand U25304 (N_25304,N_20327,N_20944);
nand U25305 (N_25305,N_20376,N_19469);
nand U25306 (N_25306,N_19960,N_18444);
and U25307 (N_25307,N_18134,N_22153);
or U25308 (N_25308,N_18785,N_22779);
nand U25309 (N_25309,N_18961,N_22265);
nor U25310 (N_25310,N_21959,N_21050);
or U25311 (N_25311,N_22364,N_18893);
xor U25312 (N_25312,N_23836,N_22068);
nand U25313 (N_25313,N_23332,N_18689);
xor U25314 (N_25314,N_21491,N_20913);
and U25315 (N_25315,N_23753,N_20552);
or U25316 (N_25316,N_23348,N_20797);
or U25317 (N_25317,N_23201,N_20938);
nor U25318 (N_25318,N_18951,N_18789);
and U25319 (N_25319,N_22793,N_23127);
or U25320 (N_25320,N_22347,N_20023);
nor U25321 (N_25321,N_19557,N_18858);
nor U25322 (N_25322,N_20830,N_18103);
or U25323 (N_25323,N_19709,N_18039);
or U25324 (N_25324,N_23909,N_21592);
or U25325 (N_25325,N_19673,N_21517);
nor U25326 (N_25326,N_22366,N_19048);
or U25327 (N_25327,N_18169,N_23334);
or U25328 (N_25328,N_21965,N_18236);
or U25329 (N_25329,N_23536,N_18024);
or U25330 (N_25330,N_21068,N_21963);
nor U25331 (N_25331,N_23151,N_21903);
and U25332 (N_25332,N_23740,N_18853);
and U25333 (N_25333,N_20354,N_22307);
and U25334 (N_25334,N_23035,N_21049);
and U25335 (N_25335,N_18508,N_20178);
nor U25336 (N_25336,N_22928,N_18332);
nor U25337 (N_25337,N_23276,N_21839);
xnor U25338 (N_25338,N_21659,N_23278);
and U25339 (N_25339,N_23105,N_19829);
nand U25340 (N_25340,N_23686,N_22852);
nand U25341 (N_25341,N_18383,N_18562);
nand U25342 (N_25342,N_23495,N_18978);
nor U25343 (N_25343,N_20613,N_18512);
or U25344 (N_25344,N_21683,N_18828);
nor U25345 (N_25345,N_19128,N_22048);
xor U25346 (N_25346,N_21596,N_20776);
xor U25347 (N_25347,N_20191,N_23344);
and U25348 (N_25348,N_20173,N_23279);
nand U25349 (N_25349,N_20125,N_22517);
nand U25350 (N_25350,N_19567,N_23973);
or U25351 (N_25351,N_22405,N_20602);
nand U25352 (N_25352,N_19644,N_23422);
or U25353 (N_25353,N_20947,N_21467);
xnor U25354 (N_25354,N_18831,N_21199);
and U25355 (N_25355,N_21411,N_22032);
nand U25356 (N_25356,N_23427,N_21283);
and U25357 (N_25357,N_21412,N_23271);
xnor U25358 (N_25358,N_21124,N_18582);
nand U25359 (N_25359,N_23076,N_20264);
nor U25360 (N_25360,N_23409,N_22741);
nand U25361 (N_25361,N_23937,N_23895);
or U25362 (N_25362,N_19670,N_22897);
and U25363 (N_25363,N_21835,N_23292);
and U25364 (N_25364,N_22422,N_21344);
xnor U25365 (N_25365,N_22242,N_20441);
and U25366 (N_25366,N_18091,N_19816);
and U25367 (N_25367,N_19330,N_20013);
nand U25368 (N_25368,N_18881,N_20992);
nand U25369 (N_25369,N_19213,N_22770);
xor U25370 (N_25370,N_21678,N_20859);
xnor U25371 (N_25371,N_22677,N_18556);
nand U25372 (N_25372,N_21721,N_22209);
or U25373 (N_25373,N_22831,N_22855);
xor U25374 (N_25374,N_20390,N_18170);
xnor U25375 (N_25375,N_22358,N_18515);
nand U25376 (N_25376,N_19257,N_21384);
or U25377 (N_25377,N_18076,N_22226);
or U25378 (N_25378,N_23809,N_22374);
nor U25379 (N_25379,N_23977,N_18943);
nand U25380 (N_25380,N_22772,N_20899);
or U25381 (N_25381,N_19586,N_20868);
or U25382 (N_25382,N_21249,N_22713);
xnor U25383 (N_25383,N_22965,N_22300);
nand U25384 (N_25384,N_18228,N_21483);
nor U25385 (N_25385,N_23033,N_21779);
or U25386 (N_25386,N_21995,N_23062);
xnor U25387 (N_25387,N_23030,N_21464);
nand U25388 (N_25388,N_22055,N_19135);
nor U25389 (N_25389,N_20805,N_21191);
nor U25390 (N_25390,N_23930,N_23656);
and U25391 (N_25391,N_18777,N_21932);
xor U25392 (N_25392,N_20965,N_23111);
xor U25393 (N_25393,N_18797,N_19635);
or U25394 (N_25394,N_21905,N_20977);
xor U25395 (N_25395,N_21414,N_19906);
xor U25396 (N_25396,N_21189,N_22947);
and U25397 (N_25397,N_22372,N_18394);
nor U25398 (N_25398,N_19438,N_19317);
and U25399 (N_25399,N_19768,N_23998);
and U25400 (N_25400,N_19389,N_20073);
nor U25401 (N_25401,N_21694,N_20940);
and U25402 (N_25402,N_23219,N_20873);
xnor U25403 (N_25403,N_22746,N_20930);
nand U25404 (N_25404,N_20318,N_20388);
and U25405 (N_25405,N_19625,N_22716);
nor U25406 (N_25406,N_21257,N_20467);
and U25407 (N_25407,N_20228,N_18476);
or U25408 (N_25408,N_19990,N_21266);
or U25409 (N_25409,N_22246,N_21201);
or U25410 (N_25410,N_21894,N_19928);
nand U25411 (N_25411,N_20109,N_19781);
nand U25412 (N_25412,N_18734,N_19405);
and U25413 (N_25413,N_21949,N_20813);
or U25414 (N_25414,N_23772,N_21590);
or U25415 (N_25415,N_19682,N_21912);
nand U25416 (N_25416,N_19217,N_22322);
and U25417 (N_25417,N_18043,N_22365);
or U25418 (N_25418,N_21605,N_20445);
and U25419 (N_25419,N_21428,N_19484);
nand U25420 (N_25420,N_19125,N_20534);
and U25421 (N_25421,N_21250,N_18111);
and U25422 (N_25422,N_18721,N_23237);
nand U25423 (N_25423,N_18987,N_19924);
nand U25424 (N_25424,N_18815,N_21440);
or U25425 (N_25425,N_20031,N_22428);
or U25426 (N_25426,N_21512,N_23721);
xor U25427 (N_25427,N_22291,N_19319);
nor U25428 (N_25428,N_21162,N_21073);
nand U25429 (N_25429,N_23306,N_19643);
xnor U25430 (N_25430,N_20533,N_20215);
or U25431 (N_25431,N_18205,N_18953);
nor U25432 (N_25432,N_20989,N_22045);
and U25433 (N_25433,N_23720,N_23545);
xor U25434 (N_25434,N_22525,N_22566);
or U25435 (N_25435,N_18798,N_18669);
xnor U25436 (N_25436,N_23808,N_20810);
or U25437 (N_25437,N_21032,N_21409);
and U25438 (N_25438,N_19366,N_20666);
and U25439 (N_25439,N_18427,N_20863);
nor U25440 (N_25440,N_22094,N_21320);
nor U25441 (N_25441,N_18759,N_23594);
or U25442 (N_25442,N_19302,N_18659);
xnor U25443 (N_25443,N_18637,N_22515);
nand U25444 (N_25444,N_18726,N_22479);
or U25445 (N_25445,N_21697,N_23040);
nor U25446 (N_25446,N_19604,N_22845);
and U25447 (N_25447,N_20653,N_20427);
nor U25448 (N_25448,N_20381,N_20482);
xor U25449 (N_25449,N_21811,N_22102);
and U25450 (N_25450,N_20432,N_19734);
nor U25451 (N_25451,N_20956,N_20692);
xnor U25452 (N_25452,N_19515,N_19236);
xor U25453 (N_25453,N_20476,N_18649);
or U25454 (N_25454,N_21035,N_22618);
xor U25455 (N_25455,N_19129,N_18275);
and U25456 (N_25456,N_22580,N_18414);
nand U25457 (N_25457,N_22575,N_22528);
nor U25458 (N_25458,N_20260,N_22100);
or U25459 (N_25459,N_21227,N_23781);
xnor U25460 (N_25460,N_22862,N_20725);
nor U25461 (N_25461,N_21229,N_21176);
and U25462 (N_25462,N_21089,N_22201);
nand U25463 (N_25463,N_18775,N_23150);
and U25464 (N_25464,N_20966,N_18118);
and U25465 (N_25465,N_18402,N_21628);
nor U25466 (N_25466,N_22985,N_23657);
and U25467 (N_25467,N_22223,N_20836);
and U25468 (N_25468,N_19531,N_20038);
nand U25469 (N_25469,N_19962,N_21055);
nand U25470 (N_25470,N_22304,N_22375);
or U25471 (N_25471,N_19055,N_18545);
and U25472 (N_25472,N_18156,N_21541);
xnor U25473 (N_25473,N_19419,N_23185);
nand U25474 (N_25474,N_22057,N_20396);
and U25475 (N_25475,N_18754,N_20974);
xor U25476 (N_25476,N_22903,N_23661);
xor U25477 (N_25477,N_18198,N_20835);
or U25478 (N_25478,N_23777,N_20858);
or U25479 (N_25479,N_21550,N_19139);
or U25480 (N_25480,N_18544,N_19828);
and U25481 (N_25481,N_21549,N_19315);
xor U25482 (N_25482,N_22884,N_22630);
xor U25483 (N_25483,N_22259,N_22695);
xor U25484 (N_25484,N_19882,N_23103);
xor U25485 (N_25485,N_21534,N_21643);
and U25486 (N_25486,N_21759,N_23704);
or U25487 (N_25487,N_22349,N_23063);
nand U25488 (N_25488,N_20419,N_23257);
or U25489 (N_25489,N_22684,N_22249);
and U25490 (N_25490,N_22919,N_18690);
xor U25491 (N_25491,N_19566,N_22554);
nand U25492 (N_25492,N_23653,N_18202);
nor U25493 (N_25493,N_19473,N_21914);
xor U25494 (N_25494,N_21994,N_21268);
and U25495 (N_25495,N_20779,N_18923);
nor U25496 (N_25496,N_18752,N_22053);
nand U25497 (N_25497,N_22009,N_23261);
and U25498 (N_25498,N_18501,N_22207);
nor U25499 (N_25499,N_22908,N_19372);
or U25500 (N_25500,N_21614,N_23875);
or U25501 (N_25501,N_22820,N_23733);
nand U25502 (N_25502,N_20945,N_18711);
and U25503 (N_25503,N_21989,N_22413);
xor U25504 (N_25504,N_19482,N_23885);
nand U25505 (N_25505,N_20357,N_19631);
nor U25506 (N_25506,N_18027,N_21235);
xnor U25507 (N_25507,N_21063,N_18088);
and U25508 (N_25508,N_22234,N_19804);
nand U25509 (N_25509,N_19580,N_18926);
xnor U25510 (N_25510,N_18868,N_22458);
and U25511 (N_25511,N_18696,N_18477);
xor U25512 (N_25512,N_23756,N_21429);
nand U25513 (N_25513,N_21430,N_18920);
nand U25514 (N_25514,N_20607,N_20059);
xnor U25515 (N_25515,N_23101,N_23823);
nand U25516 (N_25516,N_19057,N_21972);
nor U25517 (N_25517,N_18958,N_23776);
or U25518 (N_25518,N_19503,N_20620);
or U25519 (N_25519,N_22013,N_19743);
nand U25520 (N_25520,N_22182,N_20549);
and U25521 (N_25521,N_23032,N_22293);
and U25522 (N_25522,N_18490,N_23950);
or U25523 (N_25523,N_23223,N_21077);
or U25524 (N_25524,N_21248,N_18555);
xor U25525 (N_25525,N_22702,N_22980);
nor U25526 (N_25526,N_20622,N_21103);
or U25527 (N_25527,N_20604,N_18016);
and U25528 (N_25528,N_19611,N_22662);
nor U25529 (N_25529,N_21159,N_18321);
nor U25530 (N_25530,N_23448,N_18439);
nand U25531 (N_25531,N_22557,N_21633);
xor U25532 (N_25532,N_20407,N_20498);
or U25533 (N_25533,N_21462,N_22359);
nand U25534 (N_25534,N_19536,N_22140);
and U25535 (N_25535,N_19685,N_18179);
or U25536 (N_25536,N_19961,N_19028);
nand U25537 (N_25537,N_18884,N_20067);
xnor U25538 (N_25538,N_22798,N_22012);
nor U25539 (N_25539,N_22591,N_19951);
nand U25540 (N_25540,N_23000,N_22385);
and U25541 (N_25541,N_18168,N_23372);
xor U25542 (N_25542,N_22921,N_23117);
nor U25543 (N_25543,N_18875,N_19821);
nor U25544 (N_25544,N_19117,N_22146);
nand U25545 (N_25545,N_19827,N_22511);
and U25546 (N_25546,N_22395,N_18857);
or U25547 (N_25547,N_19460,N_18701);
xor U25548 (N_25548,N_21648,N_20579);
and U25549 (N_25549,N_20637,N_23146);
nand U25550 (N_25550,N_19374,N_18909);
or U25551 (N_25551,N_18151,N_18097);
and U25552 (N_25552,N_22948,N_23621);
nand U25553 (N_25553,N_21808,N_19095);
nor U25554 (N_25554,N_19023,N_20152);
nor U25555 (N_25555,N_22936,N_18995);
or U25556 (N_25556,N_23945,N_20694);
and U25557 (N_25557,N_18165,N_21034);
nor U25558 (N_25558,N_20599,N_19263);
xnor U25559 (N_25559,N_21695,N_21253);
xor U25560 (N_25560,N_23393,N_18025);
nor U25561 (N_25561,N_20838,N_18099);
and U25562 (N_25562,N_22253,N_23663);
nand U25563 (N_25563,N_21698,N_20255);
xnor U25564 (N_25564,N_23295,N_20097);
xor U25565 (N_25565,N_22112,N_19426);
or U25566 (N_25566,N_20603,N_18225);
nand U25567 (N_25567,N_21967,N_22523);
nor U25568 (N_25568,N_20296,N_23090);
nand U25569 (N_25569,N_19774,N_19480);
xnor U25570 (N_25570,N_23675,N_23533);
and U25571 (N_25571,N_18655,N_20242);
nor U25572 (N_25572,N_18991,N_18530);
or U25573 (N_25573,N_23226,N_20466);
xnor U25574 (N_25574,N_21139,N_22022);
xnor U25575 (N_25575,N_22641,N_19858);
nand U25576 (N_25576,N_22614,N_23307);
nor U25577 (N_25577,N_18086,N_21898);
and U25578 (N_25578,N_20134,N_20050);
nor U25579 (N_25579,N_18438,N_20907);
or U25580 (N_25580,N_23898,N_20304);
nor U25581 (N_25581,N_21503,N_23519);
nor U25582 (N_25582,N_20470,N_19718);
xnor U25583 (N_25583,N_20792,N_19424);
or U25584 (N_25584,N_21295,N_18368);
nor U25585 (N_25585,N_21236,N_23199);
nand U25586 (N_25586,N_19101,N_18260);
xor U25587 (N_25587,N_21327,N_19622);
nor U25588 (N_25588,N_22518,N_21601);
xor U25589 (N_25589,N_22709,N_21492);
and U25590 (N_25590,N_19324,N_19215);
xor U25591 (N_25591,N_21613,N_18313);
xor U25592 (N_25592,N_19825,N_19264);
nor U25593 (N_25593,N_23642,N_19422);
or U25594 (N_25594,N_18615,N_22049);
nor U25595 (N_25595,N_20481,N_20884);
or U25596 (N_25596,N_21979,N_20433);
xor U25597 (N_25597,N_23801,N_22509);
and U25598 (N_25598,N_19759,N_21709);
nor U25599 (N_25599,N_21872,N_22186);
xor U25600 (N_25600,N_18548,N_20923);
xor U25601 (N_25601,N_19921,N_23559);
or U25602 (N_25602,N_22062,N_21572);
and U25603 (N_25603,N_23383,N_18713);
nor U25604 (N_25604,N_18354,N_20371);
xor U25605 (N_25605,N_23695,N_19919);
and U25606 (N_25606,N_21766,N_19014);
nor U25607 (N_25607,N_23255,N_22237);
and U25608 (N_25608,N_23554,N_20107);
xor U25609 (N_25609,N_18375,N_22036);
and U25610 (N_25610,N_19185,N_22067);
xor U25611 (N_25611,N_19411,N_19748);
or U25612 (N_25612,N_20449,N_18456);
nand U25613 (N_25613,N_21406,N_21654);
or U25614 (N_25614,N_22521,N_20452);
nand U25615 (N_25615,N_23471,N_22326);
nor U25616 (N_25616,N_23585,N_23584);
nand U25617 (N_25617,N_20351,N_21506);
nand U25618 (N_25618,N_22771,N_23919);
and U25619 (N_25619,N_18454,N_19984);
xor U25620 (N_25620,N_23900,N_18739);
or U25621 (N_25621,N_18137,N_18373);
nor U25622 (N_25622,N_19639,N_22232);
nor U25623 (N_25623,N_20856,N_20998);
xnor U25624 (N_25624,N_23326,N_23423);
nor U25625 (N_25625,N_23245,N_21510);
nand U25626 (N_25626,N_20686,N_21999);
xor U25627 (N_25627,N_22212,N_18057);
xnor U25628 (N_25628,N_23810,N_20036);
and U25629 (N_25629,N_23509,N_19878);
and U25630 (N_25630,N_18906,N_23026);
nand U25631 (N_25631,N_18207,N_19719);
xor U25632 (N_25632,N_18407,N_23768);
or U25633 (N_25633,N_19207,N_22812);
xnor U25634 (N_25634,N_19811,N_22466);
or U25635 (N_25635,N_20234,N_23217);
nor U25636 (N_25636,N_20898,N_21488);
xor U25637 (N_25637,N_21576,N_22281);
nand U25638 (N_25638,N_19123,N_23155);
nor U25639 (N_25639,N_21828,N_21889);
or U25640 (N_25640,N_18418,N_22397);
nor U25641 (N_25641,N_23660,N_22189);
nand U25642 (N_25642,N_18237,N_20282);
and U25643 (N_25643,N_21842,N_23002);
nor U25644 (N_25644,N_21134,N_20410);
nand U25645 (N_25645,N_23317,N_20003);
xnor U25646 (N_25646,N_20122,N_20591);
or U25647 (N_25647,N_21094,N_23735);
nor U25648 (N_25648,N_19118,N_22931);
and U25649 (N_25649,N_22613,N_23066);
and U25650 (N_25650,N_21366,N_23243);
and U25651 (N_25651,N_21542,N_19009);
and U25652 (N_25652,N_23691,N_21481);
xor U25653 (N_25653,N_23270,N_22697);
xnor U25654 (N_25654,N_23136,N_19691);
or U25655 (N_25655,N_19815,N_19394);
or U25656 (N_25656,N_22804,N_21190);
or U25657 (N_25657,N_21799,N_23622);
and U25658 (N_25658,N_21376,N_23963);
or U25659 (N_25659,N_22111,N_20756);
and U25660 (N_25660,N_20617,N_22079);
and U25661 (N_25661,N_20087,N_21847);
nor U25662 (N_25662,N_19554,N_21526);
xor U25663 (N_25663,N_19757,N_18938);
or U25664 (N_25664,N_19871,N_22836);
nand U25665 (N_25665,N_22376,N_18506);
and U25666 (N_25666,N_21308,N_21022);
xnor U25667 (N_25667,N_21285,N_18787);
and U25668 (N_25668,N_19314,N_19671);
xor U25669 (N_25669,N_19971,N_23434);
nor U25670 (N_25670,N_20897,N_20080);
xor U25671 (N_25671,N_23082,N_21700);
nand U25672 (N_25672,N_19076,N_21417);
and U25673 (N_25673,N_18964,N_20172);
nand U25674 (N_25674,N_21907,N_19977);
and U25675 (N_25675,N_19342,N_23876);
and U25676 (N_25676,N_18143,N_21018);
and U25677 (N_25677,N_19767,N_23563);
xor U25678 (N_25678,N_21730,N_23184);
or U25679 (N_25679,N_19401,N_23980);
and U25680 (N_25680,N_21075,N_21974);
or U25681 (N_25681,N_21194,N_22786);
and U25682 (N_25682,N_20910,N_18329);
nor U25683 (N_25683,N_23290,N_19922);
and U25684 (N_25684,N_18933,N_18838);
or U25685 (N_25685,N_20258,N_22286);
and U25686 (N_25686,N_23927,N_23424);
nand U25687 (N_25687,N_23929,N_22915);
nor U25688 (N_25688,N_21346,N_19245);
nand U25689 (N_25689,N_21312,N_18595);
nor U25690 (N_25690,N_20241,N_22625);
nor U25691 (N_25691,N_20145,N_21757);
nand U25692 (N_25692,N_22390,N_18588);
nor U25693 (N_25693,N_23104,N_21619);
or U25694 (N_25694,N_22346,N_18315);
xnor U25695 (N_25695,N_19680,N_18030);
or U25696 (N_25696,N_22686,N_19303);
xnor U25697 (N_25697,N_21149,N_21132);
nand U25698 (N_25698,N_19917,N_22455);
nor U25699 (N_25699,N_22629,N_21982);
or U25700 (N_25700,N_23550,N_20808);
nor U25701 (N_25701,N_22781,N_18160);
or U25702 (N_25702,N_22325,N_20968);
and U25703 (N_25703,N_19126,N_20744);
xor U25704 (N_25704,N_23248,N_20102);
nand U25705 (N_25705,N_19826,N_21881);
nand U25706 (N_25706,N_18436,N_23947);
nand U25707 (N_25707,N_22801,N_21274);
or U25708 (N_25708,N_23075,N_21254);
nor U25709 (N_25709,N_20723,N_22089);
nand U25710 (N_25710,N_22688,N_23378);
nor U25711 (N_25711,N_19835,N_18059);
nor U25712 (N_25712,N_23934,N_22262);
nand U25713 (N_25713,N_21918,N_20320);
and U25714 (N_25714,N_20569,N_23282);
nand U25715 (N_25715,N_21672,N_23380);
nand U25716 (N_25716,N_23558,N_21469);
and U25717 (N_25717,N_18799,N_18528);
nor U25718 (N_25718,N_22767,N_18398);
or U25719 (N_25719,N_19229,N_21045);
and U25720 (N_25720,N_19110,N_20932);
and U25721 (N_25721,N_23859,N_22840);
nand U25722 (N_25722,N_20213,N_19052);
nor U25723 (N_25723,N_23466,N_21902);
nor U25724 (N_25724,N_21857,N_20428);
or U25725 (N_25725,N_18762,N_23569);
or U25726 (N_25726,N_18763,N_23022);
or U25727 (N_25727,N_18340,N_22379);
nor U25728 (N_25728,N_20293,N_23905);
nand U25729 (N_25729,N_23179,N_21002);
xnor U25730 (N_25730,N_20815,N_19998);
xnor U25731 (N_25731,N_18570,N_22093);
nor U25732 (N_25732,N_22217,N_22537);
nand U25733 (N_25733,N_20115,N_20834);
nor U25734 (N_25734,N_23251,N_21123);
nor U25735 (N_25735,N_20854,N_22176);
nor U25736 (N_25736,N_18200,N_20439);
nor U25737 (N_25737,N_23760,N_21038);
and U25738 (N_25738,N_22611,N_21873);
nand U25739 (N_25739,N_23446,N_21765);
nand U25740 (N_25740,N_20261,N_22231);
nor U25741 (N_25741,N_21071,N_18223);
or U25742 (N_25742,N_23053,N_23683);
nand U25743 (N_25743,N_18764,N_23335);
or U25744 (N_25744,N_22639,N_22343);
nor U25745 (N_25745,N_23181,N_23328);
nor U25746 (N_25746,N_18820,N_21609);
and U25747 (N_25747,N_21362,N_18668);
or U25748 (N_25748,N_21988,N_18623);
nor U25749 (N_25749,N_22438,N_20088);
nand U25750 (N_25750,N_22872,N_22953);
nor U25751 (N_25751,N_19131,N_21290);
nor U25752 (N_25752,N_23419,N_21877);
nand U25753 (N_25753,N_20740,N_20594);
or U25754 (N_25754,N_19173,N_18965);
or U25755 (N_25755,N_19376,N_19608);
xor U25756 (N_25756,N_18392,N_20548);
or U25757 (N_25757,N_22942,N_18335);
xnor U25758 (N_25758,N_21615,N_20132);
xor U25759 (N_25759,N_20916,N_19331);
xor U25760 (N_25760,N_19163,N_21205);
nand U25761 (N_25761,N_21147,N_20248);
nand U25762 (N_25762,N_18351,N_23716);
xnor U25763 (N_25763,N_21909,N_19284);
xor U25764 (N_25764,N_19654,N_18079);
or U25765 (N_25765,N_18277,N_21583);
or U25766 (N_25766,N_22895,N_18369);
nor U25767 (N_25767,N_20997,N_20483);
nand U25768 (N_25768,N_23514,N_19985);
and U25769 (N_25769,N_23436,N_19400);
and U25770 (N_25770,N_21390,N_20822);
and U25771 (N_25771,N_19839,N_18492);
nor U25772 (N_25772,N_21655,N_21639);
nand U25773 (N_25773,N_23080,N_18052);
nand U25774 (N_25774,N_20317,N_19876);
nand U25775 (N_25775,N_18496,N_18247);
nand U25776 (N_25776,N_19294,N_19150);
or U25777 (N_25777,N_22833,N_20519);
nor U25778 (N_25778,N_22171,N_21612);
nor U25779 (N_25779,N_20499,N_21357);
nor U25780 (N_25780,N_21302,N_22174);
or U25781 (N_25781,N_19883,N_18505);
xor U25782 (N_25782,N_21888,N_21231);
or U25783 (N_25783,N_20012,N_20005);
or U25784 (N_25784,N_18539,N_22932);
xor U25785 (N_25785,N_20717,N_18625);
or U25786 (N_25786,N_23830,N_18012);
nor U25787 (N_25787,N_18092,N_19820);
nand U25788 (N_25788,N_22156,N_20539);
xor U25789 (N_25789,N_22877,N_22655);
and U25790 (N_25790,N_22107,N_18180);
and U25791 (N_25791,N_18096,N_23285);
nand U25792 (N_25792,N_23770,N_23083);
nand U25793 (N_25793,N_23399,N_18807);
and U25794 (N_25794,N_19669,N_18396);
nor U25795 (N_25795,N_23815,N_18597);
nor U25796 (N_25796,N_21665,N_19403);
and U25797 (N_25797,N_23067,N_20961);
nor U25798 (N_25798,N_20746,N_18718);
and U25799 (N_25799,N_19677,N_22310);
and U25800 (N_25800,N_21131,N_18026);
xor U25801 (N_25801,N_20186,N_23879);
or U25802 (N_25802,N_19796,N_19099);
and U25803 (N_25803,N_20864,N_22540);
xnor U25804 (N_25804,N_23428,N_18058);
and U25805 (N_25805,N_19478,N_20029);
nand U25806 (N_25806,N_22279,N_18643);
and U25807 (N_25807,N_21193,N_22930);
or U25808 (N_25808,N_21728,N_22085);
nand U25809 (N_25809,N_19087,N_20148);
xnor U25810 (N_25810,N_23112,N_21475);
xor U25811 (N_25811,N_23333,N_22162);
xor U25812 (N_25812,N_22001,N_20227);
xnor U25813 (N_25813,N_19075,N_23311);
nand U25814 (N_25814,N_21129,N_19731);
xor U25815 (N_25815,N_19676,N_22729);
and U25816 (N_25816,N_20557,N_19459);
nand U25817 (N_25817,N_19824,N_21931);
and U25818 (N_25818,N_18925,N_18683);
xnor U25819 (N_25819,N_18911,N_18589);
or U25820 (N_25820,N_20642,N_18907);
and U25821 (N_25821,N_18940,N_19582);
nand U25822 (N_25822,N_20823,N_21689);
xnor U25823 (N_25823,N_21088,N_19094);
xnor U25824 (N_25824,N_18068,N_21410);
xor U25825 (N_25825,N_20021,N_22027);
nand U25826 (N_25826,N_19909,N_23619);
nor U25827 (N_25827,N_21836,N_19205);
xnor U25828 (N_25828,N_19599,N_21893);
xor U25829 (N_25829,N_23955,N_23310);
nand U25830 (N_25830,N_20766,N_21891);
xor U25831 (N_25831,N_20625,N_19703);
nand U25832 (N_25832,N_21395,N_20268);
nor U25833 (N_25833,N_19427,N_21433);
xor U25834 (N_25834,N_22484,N_23889);
and U25835 (N_25835,N_18206,N_21023);
nand U25836 (N_25836,N_23059,N_19642);
and U25837 (N_25837,N_22028,N_19568);
and U25838 (N_25838,N_22051,N_18804);
and U25839 (N_25839,N_21603,N_23043);
nand U25840 (N_25840,N_19395,N_19396);
or U25841 (N_25841,N_22650,N_23620);
nand U25842 (N_25842,N_19913,N_20298);
xor U25843 (N_25843,N_22199,N_22761);
nand U25844 (N_25844,N_23700,N_22658);
and U25845 (N_25845,N_20741,N_21472);
or U25846 (N_25846,N_18550,N_21246);
xnor U25847 (N_25847,N_21165,N_19404);
nor U25848 (N_25848,N_19797,N_19371);
xnor U25849 (N_25849,N_18761,N_20659);
or U25850 (N_25850,N_19024,N_19291);
or U25851 (N_25851,N_19530,N_22901);
and U25852 (N_25852,N_19901,N_22807);
or U25853 (N_25853,N_22324,N_22690);
or U25854 (N_25854,N_19454,N_18239);
xnor U25855 (N_25855,N_20737,N_23193);
and U25856 (N_25856,N_21198,N_18537);
nand U25857 (N_25857,N_22740,N_20581);
and U25858 (N_25858,N_21815,N_18421);
and U25859 (N_25859,N_19428,N_18936);
xor U25860 (N_25860,N_21316,N_19583);
and U25861 (N_25861,N_22473,N_23203);
or U25862 (N_25862,N_22818,N_23651);
nor U25863 (N_25863,N_18841,N_18393);
and U25864 (N_25864,N_19407,N_21896);
and U25865 (N_25865,N_18581,N_19329);
nand U25866 (N_25866,N_20237,N_18176);
nand U25867 (N_25867,N_22319,N_21781);
or U25868 (N_25868,N_22914,N_23366);
or U25869 (N_25869,N_19410,N_20096);
and U25870 (N_25870,N_21375,N_20839);
xnor U25871 (N_25871,N_23122,N_19109);
nor U25872 (N_25872,N_21457,N_21772);
nand U25873 (N_25873,N_18325,N_23645);
xnor U25874 (N_25874,N_20490,N_23865);
xor U25875 (N_25875,N_20345,N_23828);
nand U25876 (N_25876,N_18896,N_23336);
and U25877 (N_25877,N_18495,N_21555);
nand U25878 (N_25878,N_18301,N_18047);
nor U25879 (N_25879,N_20857,N_21392);
and U25880 (N_25880,N_18956,N_23342);
or U25881 (N_25881,N_23451,N_19609);
nand U25882 (N_25882,N_19398,N_19299);
or U25883 (N_25883,N_22927,N_22181);
xor U25884 (N_25884,N_20055,N_19439);
or U25885 (N_25885,N_23156,N_22288);
xnor U25886 (N_25886,N_21970,N_23438);
nor U25887 (N_25887,N_20951,N_19100);
or U25888 (N_25888,N_21394,N_20435);
and U25889 (N_25889,N_23586,N_22707);
nor U25890 (N_25890,N_18681,N_21287);
xor U25891 (N_25891,N_21040,N_21760);
and U25892 (N_25892,N_20442,N_19313);
nor U25893 (N_25893,N_21444,N_19899);
and U25894 (N_25894,N_23361,N_22060);
and U25895 (N_25895,N_20143,N_19353);
xnor U25896 (N_25896,N_22749,N_22687);
or U25897 (N_25897,N_19941,N_23321);
nor U25898 (N_25898,N_20301,N_21053);
xnor U25899 (N_25899,N_22803,N_20473);
and U25900 (N_25900,N_21403,N_21108);
xor U25901 (N_25901,N_23641,N_19464);
nor U25902 (N_25902,N_19432,N_21447);
and U25903 (N_25903,N_20216,N_18968);
nor U25904 (N_25904,N_21477,N_23308);
nand U25905 (N_25905,N_21110,N_20378);
xor U25906 (N_25906,N_20914,N_20353);
nand U25907 (N_25907,N_18227,N_18208);
xnor U25908 (N_25908,N_23527,N_19539);
and U25909 (N_25909,N_23038,N_20844);
xor U25910 (N_25910,N_22783,N_19617);
and U25911 (N_25911,N_21143,N_18840);
or U25912 (N_25912,N_22933,N_23345);
nand U25913 (N_25913,N_22830,N_19846);
or U25914 (N_25914,N_21632,N_22229);
xnor U25915 (N_25915,N_21210,N_19937);
xnor U25916 (N_25916,N_18189,N_20414);
nand U25917 (N_25917,N_23707,N_21563);
xor U25918 (N_25918,N_20949,N_19378);
or U25919 (N_25919,N_23731,N_21361);
nor U25920 (N_25920,N_23167,N_20131);
nor U25921 (N_25921,N_21589,N_20157);
or U25922 (N_25922,N_23440,N_20361);
nand U25923 (N_25923,N_22827,N_20784);
nor U25924 (N_25924,N_18390,N_21452);
nor U25925 (N_25925,N_19765,N_18697);
or U25926 (N_25926,N_20374,N_18732);
nand U25927 (N_25927,N_23983,N_21127);
nor U25928 (N_25928,N_23816,N_22896);
and U25929 (N_25929,N_21037,N_22544);
xnor U25930 (N_25930,N_23701,N_23296);
xnor U25931 (N_25931,N_18644,N_18001);
and U25932 (N_25932,N_19068,N_20331);
xnor U25933 (N_25933,N_22469,N_21736);
xnor U25934 (N_25934,N_20397,N_20510);
or U25935 (N_25935,N_23233,N_21978);
nor U25936 (N_25936,N_22247,N_20825);
or U25937 (N_25937,N_19005,N_22260);
and U25938 (N_25938,N_20085,N_23081);
nor U25939 (N_25939,N_19895,N_23009);
xor U25940 (N_25940,N_18035,N_22240);
or U25941 (N_25941,N_18453,N_20734);
nor U25942 (N_25942,N_23088,N_18767);
xnor U25943 (N_25943,N_18832,N_18116);
and U25944 (N_25944,N_19104,N_20098);
nand U25945 (N_25945,N_22072,N_21637);
nand U25946 (N_25946,N_19970,N_18386);
and U25947 (N_25947,N_18546,N_20895);
nor U25948 (N_25948,N_22255,N_20568);
nor U25949 (N_25949,N_19544,N_23916);
or U25950 (N_25950,N_23314,N_23159);
and U25951 (N_25951,N_18482,N_23718);
and U25952 (N_25952,N_21195,N_19160);
xor U25953 (N_25953,N_19065,N_19421);
or U25954 (N_25954,N_19003,N_19232);
nand U25955 (N_25955,N_18613,N_20888);
or U25956 (N_25956,N_18155,N_18401);
nor U25957 (N_25957,N_20016,N_19059);
and U25958 (N_25958,N_20240,N_23844);
nor U25959 (N_25959,N_21322,N_20960);
nand U25960 (N_25960,N_23390,N_21707);
nand U25961 (N_25961,N_19016,N_23124);
and U25962 (N_25962,N_23115,N_20015);
and U25963 (N_25963,N_20124,N_23573);
xor U25964 (N_25964,N_20297,N_19242);
nand U25965 (N_25965,N_19281,N_21137);
xor U25966 (N_25966,N_22294,N_20075);
xnor U25967 (N_25967,N_19847,N_19413);
nor U25968 (N_25968,N_19321,N_18053);
nand U25969 (N_25969,N_22542,N_18717);
xor U25970 (N_25970,N_21957,N_22133);
xnor U25971 (N_25971,N_21518,N_21297);
or U25972 (N_25972,N_20454,N_19887);
and U25973 (N_25973,N_20391,N_21106);
and U25974 (N_25974,N_22691,N_23848);
nand U25975 (N_25975,N_18442,N_20072);
nor U25976 (N_25976,N_21437,N_20647);
nor U25977 (N_25977,N_23266,N_23595);
nand U25978 (N_25978,N_23078,N_23194);
nand U25979 (N_25979,N_19431,N_22414);
or U25980 (N_25980,N_19497,N_19187);
nand U25981 (N_25981,N_23496,N_21880);
nor U25982 (N_25982,N_18291,N_19558);
nor U25983 (N_25983,N_18988,N_20824);
nor U25984 (N_25984,N_22082,N_21930);
or U25985 (N_25985,N_21173,N_20277);
and U25986 (N_25986,N_19581,N_22696);
and U25987 (N_25987,N_19770,N_22737);
xnor U25988 (N_25988,N_20027,N_18885);
or U25989 (N_25989,N_19259,N_18594);
nand U25990 (N_25990,N_19573,N_20198);
xnor U25991 (N_25991,N_19283,N_23375);
or U25992 (N_25992,N_20500,N_19492);
and U25993 (N_25993,N_23951,N_19175);
and U25994 (N_25994,N_22457,N_20537);
and U25995 (N_25995,N_22456,N_22582);
nor U25996 (N_25996,N_21434,N_20946);
nor U25997 (N_25997,N_18484,N_22035);
or U25998 (N_25998,N_23042,N_18483);
xor U25999 (N_25999,N_20468,N_19189);
nand U26000 (N_26000,N_23987,N_20308);
or U26001 (N_26001,N_19211,N_21692);
and U26002 (N_26002,N_20423,N_20064);
nor U26003 (N_26003,N_22934,N_21420);
and U26004 (N_26004,N_18048,N_19549);
xor U26005 (N_26005,N_18747,N_22805);
xor U26006 (N_26006,N_22822,N_19277);
xnor U26007 (N_26007,N_18081,N_20319);
or U26008 (N_26008,N_19751,N_22185);
xor U26009 (N_26009,N_19046,N_20920);
xor U26010 (N_26010,N_21962,N_21070);
and U26011 (N_26011,N_18624,N_20980);
and U26012 (N_26012,N_20763,N_21746);
nor U26013 (N_26013,N_18101,N_19383);
xnor U26014 (N_26014,N_23549,N_23762);
nand U26015 (N_26015,N_20675,N_21125);
xnor U26016 (N_26016,N_18466,N_19190);
nor U26017 (N_26017,N_18836,N_22900);
nand U26018 (N_26018,N_22720,N_21180);
nor U26019 (N_26019,N_19144,N_22865);
nand U26020 (N_26020,N_21499,N_21923);
nor U26021 (N_26021,N_20367,N_23920);
xnor U26022 (N_26022,N_22703,N_20201);
and U26023 (N_26023,N_22978,N_20771);
or U26024 (N_26024,N_22541,N_18626);
nor U26025 (N_26025,N_23305,N_22730);
and U26026 (N_26026,N_21791,N_20802);
nand U26027 (N_26027,N_18331,N_22267);
and U26028 (N_26028,N_23957,N_21764);
xnor U26029 (N_26029,N_20338,N_18793);
and U26030 (N_26030,N_18065,N_20742);
or U26031 (N_26031,N_18576,N_22533);
and U26032 (N_26032,N_20146,N_20448);
xnor U26033 (N_26033,N_18776,N_21310);
and U26034 (N_26034,N_20560,N_19880);
or U26035 (N_26035,N_22398,N_22416);
or U26036 (N_26036,N_19717,N_20409);
and U26037 (N_26037,N_20443,N_23178);
nand U26038 (N_26038,N_18935,N_21646);
xor U26039 (N_26039,N_20577,N_21586);
nor U26040 (N_26040,N_22576,N_22560);
nand U26041 (N_26041,N_21200,N_23589);
and U26042 (N_26042,N_21151,N_20615);
or U26043 (N_26043,N_21300,N_19886);
nand U26044 (N_26044,N_20288,N_20829);
nor U26045 (N_26045,N_23302,N_19660);
nor U26046 (N_26046,N_23826,N_22508);
and U26047 (N_26047,N_19730,N_22136);
xnor U26048 (N_26048,N_21187,N_22502);
nor U26049 (N_26049,N_19822,N_19365);
nor U26050 (N_26050,N_18186,N_20563);
and U26051 (N_26051,N_21084,N_18288);
xnor U26052 (N_26052,N_22498,N_21291);
or U26053 (N_26053,N_22159,N_18252);
nand U26054 (N_26054,N_23638,N_18574);
or U26055 (N_26055,N_22556,N_22382);
nand U26056 (N_26056,N_19801,N_20758);
xnor U26057 (N_26057,N_22966,N_18071);
nand U26058 (N_26058,N_22188,N_21122);
or U26059 (N_26059,N_22796,N_20377);
nand U26060 (N_26060,N_18540,N_20730);
or U26061 (N_26061,N_20285,N_18955);
nand U26062 (N_26062,N_21862,N_19904);
xnor U26063 (N_26063,N_20463,N_18140);
nor U26064 (N_26064,N_20244,N_18154);
xor U26065 (N_26065,N_23800,N_19402);
and U26066 (N_26066,N_23825,N_18745);
and U26067 (N_26067,N_20632,N_21553);
nand U26068 (N_26068,N_19121,N_23537);
xnor U26069 (N_26069,N_19621,N_23158);
nor U26070 (N_26070,N_22272,N_22287);
or U26071 (N_26071,N_22999,N_20196);
nor U26072 (N_26072,N_18327,N_21786);
nand U26073 (N_26073,N_23024,N_18821);
nand U26074 (N_26074,N_23265,N_21755);
and U26075 (N_26075,N_22378,N_20696);
and U26076 (N_26076,N_22037,N_21527);
and U26077 (N_26077,N_20876,N_20082);
and U26078 (N_26078,N_23320,N_23717);
and U26079 (N_26079,N_21146,N_18510);
or U26080 (N_26080,N_23036,N_20719);
nor U26081 (N_26081,N_21625,N_23834);
or U26082 (N_26082,N_22762,N_23995);
nor U26083 (N_26083,N_21875,N_23482);
and U26084 (N_26084,N_20456,N_18282);
or U26085 (N_26085,N_23908,N_20202);
nor U26086 (N_26086,N_23408,N_22665);
or U26087 (N_26087,N_23351,N_21951);
or U26088 (N_26088,N_18699,N_22263);
xnor U26089 (N_26089,N_21154,N_21858);
xor U26090 (N_26090,N_20646,N_22800);
and U26091 (N_26091,N_21790,N_18023);
xor U26092 (N_26092,N_22177,N_21871);
xor U26093 (N_26093,N_20010,N_22173);
or U26094 (N_26094,N_20095,N_21580);
nor U26095 (N_26095,N_18670,N_23012);
nand U26096 (N_26096,N_23503,N_18146);
nor U26097 (N_26097,N_21496,N_18422);
xor U26098 (N_26098,N_22718,N_20963);
nor U26099 (N_26099,N_22816,N_19955);
nand U26100 (N_26100,N_23100,N_21326);
or U26101 (N_26101,N_23682,N_21921);
nand U26102 (N_26102,N_18663,N_20990);
xnor U26103 (N_26103,N_19874,N_23784);
or U26104 (N_26104,N_22996,N_19244);
nand U26105 (N_26105,N_23529,N_23212);
nor U26106 (N_26106,N_18784,N_19978);
xnor U26107 (N_26107,N_20714,N_18120);
nor U26108 (N_26108,N_22252,N_22447);
nor U26109 (N_26109,N_18553,N_21460);
xor U26110 (N_26110,N_18740,N_23575);
xor U26111 (N_26111,N_19015,N_18675);
nor U26112 (N_26112,N_18379,N_19006);
nor U26113 (N_26113,N_22476,N_22340);
nand U26114 (N_26114,N_22879,N_22424);
nor U26115 (N_26115,N_23322,N_22110);
and U26116 (N_26116,N_20504,N_20702);
xor U26117 (N_26117,N_23359,N_22869);
nor U26118 (N_26118,N_22006,N_18883);
nand U26119 (N_26119,N_23394,N_20342);
and U26120 (N_26120,N_23152,N_23049);
xnor U26121 (N_26121,N_23044,N_20816);
nor U26122 (N_26122,N_18126,N_19304);
or U26123 (N_26123,N_18265,N_21564);
nor U26124 (N_26124,N_23189,N_18062);
nor U26125 (N_26125,N_23835,N_21990);
and U26126 (N_26126,N_22844,N_20121);
nor U26127 (N_26127,N_21245,N_22129);
and U26128 (N_26128,N_22943,N_21650);
nor U26129 (N_26129,N_22215,N_22442);
and U26130 (N_26130,N_23349,N_21082);
nand U26131 (N_26131,N_21816,N_20525);
or U26132 (N_26132,N_18743,N_18518);
or U26133 (N_26133,N_22607,N_21155);
nor U26134 (N_26134,N_20091,N_18428);
or U26135 (N_26135,N_23719,N_21792);
or U26136 (N_26136,N_19947,N_20188);
nand U26137 (N_26137,N_21705,N_21535);
nand U26138 (N_26138,N_19357,N_21784);
or U26139 (N_26139,N_21756,N_19040);
or U26140 (N_26140,N_23552,N_19752);
nand U26141 (N_26141,N_19033,N_22411);
nor U26142 (N_26142,N_22419,N_23921);
nand U26143 (N_26143,N_18240,N_22753);
or U26144 (N_26144,N_22539,N_23587);
and U26145 (N_26145,N_20495,N_21741);
or U26146 (N_26146,N_22097,N_19447);
nand U26147 (N_26147,N_22163,N_20128);
and U26148 (N_26148,N_18616,N_23917);
xor U26149 (N_26149,N_23166,N_21966);
xor U26150 (N_26150,N_22271,N_21832);
nand U26151 (N_26151,N_23684,N_19507);
nand U26152 (N_26152,N_23441,N_18806);
nand U26153 (N_26153,N_18536,N_21841);
nor U26154 (N_26154,N_22997,N_21493);
xor U26155 (N_26155,N_23315,N_18095);
nor U26156 (N_26156,N_19898,N_22075);
and U26157 (N_26157,N_22734,N_20210);
or U26158 (N_26158,N_21158,N_19940);
and U26159 (N_26159,N_22530,N_20129);
nor U26160 (N_26160,N_20706,N_23391);
nor U26161 (N_26161,N_22228,N_19463);
xnor U26162 (N_26162,N_20851,N_19261);
xor U26163 (N_26163,N_23388,N_18019);
xnor U26164 (N_26164,N_22031,N_23985);
nor U26165 (N_26165,N_19090,N_21666);
nor U26166 (N_26166,N_20041,N_20236);
nand U26167 (N_26167,N_21515,N_18782);
or U26168 (N_26168,N_19926,N_21251);
nor U26169 (N_26169,N_21922,N_23139);
nand U26170 (N_26170,N_20544,N_18130);
or U26171 (N_26171,N_23531,N_21498);
xor U26172 (N_26172,N_23108,N_20259);
or U26173 (N_26173,N_20084,N_19624);
nor U26174 (N_26174,N_22064,N_18032);
xor U26175 (N_26175,N_22907,N_22002);
xor U26176 (N_26176,N_20530,N_19272);
and U26177 (N_26177,N_18471,N_18022);
nor U26178 (N_26178,N_22354,N_23363);
nand U26179 (N_26179,N_18997,N_23119);
and U26180 (N_26180,N_20385,N_21048);
nor U26181 (N_26181,N_23324,N_20783);
nor U26182 (N_26182,N_19896,N_19668);
and U26183 (N_26183,N_23751,N_23890);
xnor U26184 (N_26184,N_23490,N_19134);
nor U26185 (N_26185,N_20649,N_18410);
xor U26186 (N_26186,N_18664,N_23593);
xnor U26187 (N_26187,N_21822,N_22224);
nor U26188 (N_26188,N_23376,N_23135);
xor U26189 (N_26189,N_20254,N_18293);
or U26190 (N_26190,N_22468,N_22078);
xor U26191 (N_26191,N_23668,N_19220);
or U26192 (N_26192,N_23853,N_21142);
nand U26193 (N_26193,N_20698,N_20042);
nand U26194 (N_26194,N_20197,N_23190);
xor U26195 (N_26195,N_22040,N_20943);
nor U26196 (N_26196,N_19056,N_19514);
nor U26197 (N_26197,N_22084,N_22763);
and U26198 (N_26198,N_22794,N_19466);
or U26199 (N_26199,N_23402,N_18719);
or U26200 (N_26200,N_20474,N_22429);
nand U26201 (N_26201,N_18526,N_22061);
nor U26202 (N_26202,N_21239,N_22874);
nor U26203 (N_26203,N_19354,N_23116);
nand U26204 (N_26204,N_19704,N_23630);
or U26205 (N_26205,N_18144,N_19563);
nand U26206 (N_26206,N_20905,N_18952);
xor U26207 (N_26207,N_23010,N_21789);
xor U26208 (N_26208,N_18790,N_18561);
and U26209 (N_26209,N_23073,N_22742);
nor U26210 (N_26210,N_22273,N_20438);
nand U26211 (N_26211,N_20881,N_23369);
nor U26212 (N_26212,N_20755,N_18498);
nand U26213 (N_26213,N_20512,N_21726);
xor U26214 (N_26214,N_20716,N_20768);
nor U26215 (N_26215,N_21667,N_18714);
or U26216 (N_26216,N_22532,N_19975);
or U26217 (N_26217,N_21321,N_20787);
xor U26218 (N_26218,N_19966,N_21561);
and U26219 (N_26219,N_18967,N_21885);
and U26220 (N_26220,N_19194,N_18136);
nor U26221 (N_26221,N_19111,N_19969);
and U26222 (N_26222,N_22391,N_18449);
nor U26223 (N_26223,N_18630,N_22758);
nor U26224 (N_26224,N_19338,N_19347);
nand U26225 (N_26225,N_20781,N_19805);
nand U26226 (N_26226,N_23453,N_23214);
nand U26227 (N_26227,N_20800,N_19483);
xnor U26228 (N_26228,N_18813,N_19289);
nand U26229 (N_26229,N_22297,N_19050);
and U26230 (N_26230,N_18230,N_23913);
xor U26231 (N_26231,N_21225,N_21156);
or U26232 (N_26232,N_20153,N_20556);
or U26233 (N_26233,N_20393,N_18509);
or U26234 (N_26234,N_20611,N_20794);
nor U26235 (N_26235,N_22170,N_20144);
nand U26236 (N_26236,N_19020,N_19255);
nor U26237 (N_26237,N_19499,N_22054);
or U26238 (N_26238,N_19932,N_21934);
nor U26239 (N_26239,N_20929,N_22967);
nor U26240 (N_26240,N_21072,N_18916);
xnor U26241 (N_26241,N_21060,N_20326);
and U26242 (N_26242,N_20697,N_19201);
xnor U26243 (N_26243,N_20981,N_18461);
xor U26244 (N_26244,N_20492,N_20472);
xnor U26245 (N_26245,N_19409,N_19227);
nand U26246 (N_26246,N_23343,N_19802);
and U26247 (N_26247,N_19246,N_21111);
or U26248 (N_26248,N_21359,N_23051);
nor U26249 (N_26249,N_22792,N_22296);
nor U26250 (N_26250,N_19842,N_18197);
or U26251 (N_26251,N_23287,N_20526);
or U26252 (N_26252,N_20387,N_18783);
nand U26253 (N_26253,N_22583,N_19079);
and U26254 (N_26254,N_23480,N_22574);
and U26255 (N_26255,N_20158,N_18361);
nand U26256 (N_26256,N_21865,N_20681);
and U26257 (N_26257,N_23398,N_22609);
or U26258 (N_26258,N_22891,N_23272);
nand U26259 (N_26259,N_20760,N_18542);
xor U26260 (N_26260,N_21716,N_21803);
or U26261 (N_26261,N_22585,N_22577);
xnor U26262 (N_26262,N_18610,N_19325);
xor U26263 (N_26263,N_18002,N_23679);
or U26264 (N_26264,N_22204,N_22622);
xnor U26265 (N_26265,N_20229,N_18892);
or U26266 (N_26266,N_21100,N_22472);
and U26267 (N_26267,N_18611,N_18161);
nor U26268 (N_26268,N_18602,N_23967);
xor U26269 (N_26269,N_19574,N_18871);
nand U26270 (N_26270,N_23992,N_19349);
and U26271 (N_26271,N_21296,N_20503);
or U26272 (N_26272,N_18698,N_23046);
xor U26273 (N_26273,N_20804,N_21001);
or U26274 (N_26274,N_23629,N_19305);
nor U26275 (N_26275,N_21479,N_18187);
xnor U26276 (N_26276,N_18312,N_21425);
nand U26277 (N_26277,N_22909,N_23705);
xor U26278 (N_26278,N_22108,N_23463);
nand U26279 (N_26279,N_20281,N_22205);
or U26280 (N_26280,N_19373,N_22603);
nand U26281 (N_26281,N_18238,N_21588);
nor U26282 (N_26282,N_20325,N_22847);
xor U26283 (N_26283,N_20379,N_20083);
nor U26284 (N_26284,N_23312,N_18962);
and U26285 (N_26285,N_18450,N_20263);
nand U26286 (N_26286,N_22954,N_23512);
xnor U26287 (N_26287,N_18898,N_19763);
and U26288 (N_26288,N_19380,N_21658);
xor U26289 (N_26289,N_22144,N_20535);
or U26290 (N_26290,N_20921,N_19952);
nand U26291 (N_26291,N_19663,N_21577);
nand U26292 (N_26292,N_21347,N_22549);
nor U26293 (N_26293,N_23467,N_23487);
and U26294 (N_26294,N_22825,N_23404);
nor U26295 (N_26295,N_18937,N_23241);
nand U26296 (N_26296,N_23699,N_21548);
nor U26297 (N_26297,N_21303,N_22981);
or U26298 (N_26298,N_19140,N_23192);
nor U26299 (N_26299,N_23806,N_21317);
nand U26300 (N_26300,N_19502,N_23145);
nand U26301 (N_26301,N_21271,N_18725);
and U26302 (N_26302,N_22572,N_20906);
or U26303 (N_26303,N_18423,N_20806);
or U26304 (N_26304,N_21958,N_20767);
nand U26305 (N_26305,N_20985,N_22460);
nand U26306 (N_26306,N_22680,N_19495);
nor U26307 (N_26307,N_22312,N_20685);
xnor U26308 (N_26308,N_19851,N_23938);
nor U26309 (N_26309,N_21164,N_18181);
and U26310 (N_26310,N_20891,N_18034);
or U26311 (N_26311,N_22161,N_23497);
and U26312 (N_26312,N_19988,N_20226);
nand U26313 (N_26313,N_19269,N_21968);
nand U26314 (N_26314,N_23507,N_20453);
or U26315 (N_26315,N_18455,N_20554);
or U26316 (N_26316,N_19054,N_20306);
nor U26317 (N_26317,N_18748,N_20798);
or U26318 (N_26318,N_23548,N_20402);
nor U26319 (N_26319,N_21908,N_21521);
xnor U26320 (N_26320,N_21948,N_21211);
or U26321 (N_26321,N_23504,N_21516);
and U26322 (N_26322,N_19388,N_21208);
nand U26323 (N_26323,N_23057,N_18852);
or U26324 (N_26324,N_23649,N_21797);
nand U26325 (N_26325,N_22490,N_18566);
nand U26326 (N_26326,N_19031,N_19772);
or U26327 (N_26327,N_18067,N_21991);
xor U26328 (N_26328,N_22198,N_19737);
xor U26329 (N_26329,N_18457,N_20305);
nand U26330 (N_26330,N_22432,N_20887);
xnor U26331 (N_26331,N_18468,N_23571);
nand U26332 (N_26332,N_21929,N_20333);
nor U26333 (N_26333,N_20922,N_22571);
nand U26334 (N_26334,N_20641,N_23277);
nand U26335 (N_26335,N_23089,N_22880);
nor U26336 (N_26336,N_23873,N_22724);
nand U26337 (N_26337,N_20177,N_19965);
xnor U26338 (N_26338,N_20853,N_19721);
nor U26339 (N_26339,N_20606,N_21115);
and U26340 (N_26340,N_18289,N_20689);
or U26341 (N_26341,N_21745,N_20600);
nor U26342 (N_26342,N_21126,N_19636);
xnor U26343 (N_26343,N_19226,N_23225);
nand U26344 (N_26344,N_18172,N_22412);
and U26345 (N_26345,N_20745,N_21265);
nor U26346 (N_26346,N_18049,N_21324);
xor U26347 (N_26347,N_18158,N_23933);
nor U26348 (N_26348,N_21511,N_21379);
and U26349 (N_26349,N_20933,N_22132);
xnor U26350 (N_26350,N_23524,N_19587);
and U26351 (N_26351,N_23744,N_20425);
xnor U26352 (N_26352,N_23952,N_18948);
or U26353 (N_26353,N_22623,N_19181);
nand U26354 (N_26354,N_21622,N_21192);
nor U26355 (N_26355,N_23133,N_18326);
nand U26356 (N_26356,N_21919,N_21710);
and U26357 (N_26357,N_22220,N_23690);
xnor U26358 (N_26358,N_23444,N_20350);
or U26359 (N_26359,N_21943,N_20078);
and U26360 (N_26360,N_18489,N_20878);
nor U26361 (N_26361,N_23339,N_20114);
nor U26362 (N_26362,N_18257,N_21006);
nand U26363 (N_26363,N_23662,N_20251);
xor U26364 (N_26364,N_19296,N_19840);
or U26365 (N_26365,N_20138,N_21107);
nand U26366 (N_26366,N_19764,N_18387);
and U26367 (N_26367,N_23442,N_19981);
nand U26368 (N_26368,N_20770,N_20973);
nor U26369 (N_26369,N_22645,N_23070);
nor U26370 (N_26370,N_20230,N_23072);
xnor U26371 (N_26371,N_21600,N_18305);
or U26372 (N_26372,N_19866,N_20959);
nand U26373 (N_26373,N_22923,N_22038);
or U26374 (N_26374,N_21424,N_22835);
nor U26375 (N_26375,N_23387,N_22044);
nand U26376 (N_26376,N_22008,N_19667);
or U26377 (N_26377,N_20103,N_20192);
or U26378 (N_26378,N_22633,N_18712);
nand U26379 (N_26379,N_18532,N_20754);
or U26380 (N_26380,N_19812,N_18642);
nor U26381 (N_26381,N_19697,N_20634);
nor U26382 (N_26382,N_21402,N_20640);
or U26383 (N_26383,N_22367,N_20811);
xor U26384 (N_26384,N_18203,N_23778);
nor U26385 (N_26385,N_23099,N_22589);
and U26386 (N_26386,N_20275,N_22023);
nor U26387 (N_26387,N_23780,N_23470);
xnor U26388 (N_26388,N_22906,N_19749);
xor U26389 (N_26389,N_21852,N_23303);
nor U26390 (N_26390,N_19143,N_19027);
and U26391 (N_26391,N_21977,N_19706);
xor U26392 (N_26392,N_22303,N_18872);
or U26393 (N_26393,N_19199,N_22441);
xnor U26394 (N_26394,N_21884,N_20165);
nand U26395 (N_26395,N_20695,N_23692);
or U26396 (N_26396,N_21611,N_23687);
and U26397 (N_26397,N_23435,N_22951);
and U26398 (N_26398,N_22277,N_21169);
or U26399 (N_26399,N_18330,N_18736);
or U26400 (N_26400,N_18768,N_18890);
xor U26401 (N_26401,N_18050,N_22640);
nor U26402 (N_26402,N_18148,N_22095);
nand U26403 (N_26403,N_21466,N_20828);
or U26404 (N_26404,N_23566,N_18378);
and U26405 (N_26405,N_19598,N_18253);
and U26406 (N_26406,N_22152,N_19085);
nand U26407 (N_26407,N_18080,N_22663);
xnor U26408 (N_26408,N_20011,N_20713);
nor U26409 (N_26409,N_23015,N_19506);
and U26410 (N_26410,N_18292,N_23413);
or U26411 (N_26411,N_23337,N_20375);
and U26412 (N_26412,N_18879,N_23567);
and U26413 (N_26413,N_18837,N_22504);
or U26414 (N_26414,N_20009,N_21282);
xor U26415 (N_26415,N_20166,N_23286);
or U26416 (N_26416,N_23457,N_22389);
xor U26417 (N_26417,N_23468,N_22619);
and U26418 (N_26418,N_18112,N_20889);
nor U26419 (N_26419,N_23454,N_19430);
xor U26420 (N_26420,N_23056,N_22461);
or U26421 (N_26421,N_21876,N_21734);
or U26422 (N_26422,N_20759,N_22077);
xnor U26423 (N_26423,N_21559,N_23758);
xnor U26424 (N_26424,N_22597,N_23812);
nand U26425 (N_26425,N_21400,N_22282);
nand U26426 (N_26426,N_18064,N_22998);
nand U26427 (N_26427,N_23506,N_22843);
or U26428 (N_26428,N_19525,N_22952);
xor U26429 (N_26429,N_21883,N_18773);
or U26430 (N_26430,N_22104,N_21170);
or U26431 (N_26431,N_22268,N_20370);
and U26432 (N_26432,N_22141,N_20077);
and U26433 (N_26433,N_21083,N_21036);
xnor U26434 (N_26434,N_20141,N_21706);
or U26435 (N_26435,N_21623,N_22692);
nand U26436 (N_26436,N_21758,N_23940);
nand U26437 (N_26437,N_19700,N_19393);
and U26438 (N_26438,N_20983,N_22257);
nor U26439 (N_26439,N_20867,N_18269);
xor U26440 (N_26440,N_19696,N_22784);
or U26441 (N_26441,N_23539,N_23564);
and U26442 (N_26442,N_21737,N_18750);
or U26443 (N_26443,N_20886,N_23769);
or U26444 (N_26444,N_20343,N_22888);
nand U26445 (N_26445,N_22117,N_23449);
nand U26446 (N_26446,N_21097,N_22986);
nor U26447 (N_26447,N_18145,N_20596);
xor U26448 (N_26448,N_19537,N_19788);
or U26449 (N_26449,N_19149,N_20999);
xnor U26450 (N_26450,N_22945,N_21814);
nand U26451 (N_26451,N_18264,N_18139);
and U26452 (N_26452,N_18221,N_19392);
and U26453 (N_26453,N_21584,N_23415);
nor U26454 (N_26454,N_19769,N_22752);
nand U26455 (N_26455,N_20645,N_21788);
nor U26456 (N_26456,N_18629,N_22858);
xnor U26457 (N_26457,N_20365,N_23239);
nor U26458 (N_26458,N_20431,N_23646);
or U26459 (N_26459,N_22514,N_22274);
nand U26460 (N_26460,N_23523,N_22745);
nand U26461 (N_26461,N_21964,N_21213);
xnor U26462 (N_26462,N_23560,N_21838);
and U26463 (N_26463,N_23894,N_19443);
xor U26464 (N_26464,N_18974,N_23058);
nor U26465 (N_26465,N_23685,N_22941);
or U26466 (N_26466,N_21562,N_21720);
and U26467 (N_26467,N_21843,N_19860);
xor U26468 (N_26468,N_21378,N_23520);
xnor U26469 (N_26469,N_21012,N_20420);
or U26470 (N_26470,N_18949,N_19058);
nor U26471 (N_26471,N_22018,N_21054);
nor U26472 (N_26472,N_22388,N_22588);
nand U26473 (N_26473,N_18939,N_20218);
nand U26474 (N_26474,N_20489,N_21237);
and U26475 (N_26475,N_21047,N_18020);
or U26476 (N_26476,N_18849,N_23377);
nand U26477 (N_26477,N_22606,N_23213);
xor U26478 (N_26478,N_18106,N_18005);
nand U26479 (N_26479,N_22026,N_21763);
and U26480 (N_26480,N_23580,N_22711);
xnor U26481 (N_26481,N_21845,N_21976);
xor U26482 (N_26482,N_23765,N_19929);
xor U26483 (N_26483,N_20529,N_19750);
nand U26484 (N_26484,N_23982,N_21742);
and U26485 (N_26485,N_19656,N_23128);
or U26486 (N_26486,N_22230,N_18406);
nand U26487 (N_26487,N_22506,N_23384);
and U26488 (N_26488,N_18380,N_22435);
nor U26489 (N_26489,N_20484,N_22251);
xnor U26490 (N_26490,N_19386,N_19346);
or U26491 (N_26491,N_22126,N_21221);
nor U26492 (N_26492,N_21519,N_20358);
nor U26493 (N_26493,N_19387,N_18006);
nand U26494 (N_26494,N_20364,N_22066);
nand U26495 (N_26495,N_18497,N_22866);
nor U26496 (N_26496,N_22423,N_22837);
xnor U26497 (N_26497,N_22666,N_23414);
xnor U26498 (N_26498,N_21242,N_22605);
nand U26499 (N_26499,N_19306,N_18420);
and U26500 (N_26500,N_21793,N_20400);
and U26501 (N_26501,N_22311,N_20902);
or U26502 (N_26502,N_23924,N_18316);
and U26503 (N_26503,N_18941,N_20181);
and U26504 (N_26504,N_20316,N_21052);
or U26505 (N_26505,N_18290,N_23609);
or U26506 (N_26506,N_21985,N_19638);
nor U26507 (N_26507,N_20572,N_20791);
or U26508 (N_26508,N_19723,N_22099);
xor U26509 (N_26509,N_22258,N_21450);
and U26510 (N_26510,N_21754,N_18636);
nor U26511 (N_26511,N_19450,N_22003);
nor U26512 (N_26512,N_19260,N_22893);
and U26513 (N_26513,N_22109,N_23412);
nand U26514 (N_26514,N_19164,N_22329);
and U26515 (N_26515,N_23168,N_21102);
nand U26516 (N_26516,N_23474,N_21181);
nor U26517 (N_26517,N_20272,N_19416);
nand U26518 (N_26518,N_23433,N_18448);
nor U26519 (N_26519,N_23473,N_19474);
nor U26520 (N_26520,N_19151,N_18488);
xor U26521 (N_26521,N_20123,N_19967);
nor U26522 (N_26522,N_19884,N_21031);
and U26523 (N_26523,N_23365,N_22393);
or U26524 (N_26524,N_22396,N_20670);
or U26525 (N_26525,N_20917,N_19080);
nor U26526 (N_26526,N_21261,N_18817);
or U26527 (N_26527,N_18362,N_18452);
or U26528 (N_26528,N_20668,N_18687);
nand U26529 (N_26529,N_19437,N_23833);
nand U26530 (N_26530,N_23612,N_23522);
xnor U26531 (N_26531,N_20380,N_22426);
xnor U26532 (N_26532,N_22125,N_19265);
or U26533 (N_26533,N_18286,N_21827);
xnor U26534 (N_26534,N_23708,N_21007);
and U26535 (N_26535,N_21080,N_20093);
nor U26536 (N_26536,N_22179,N_18596);
or U26537 (N_26537,N_23143,N_23922);
or U26538 (N_26538,N_21095,N_22485);
xnor U26539 (N_26539,N_19864,N_22203);
nand U26540 (N_26540,N_23899,N_21241);
or U26541 (N_26541,N_21782,N_20720);
nand U26542 (N_26542,N_19253,N_18494);
nand U26543 (N_26543,N_23055,N_18910);
and U26544 (N_26544,N_21547,N_20046);
nor U26545 (N_26545,N_21696,N_23319);
or U26546 (N_26546,N_21396,N_18864);
and U26547 (N_26547,N_23147,N_22592);
or U26548 (N_26548,N_18036,N_23483);
or U26549 (N_26549,N_19078,N_21897);
xnor U26550 (N_26550,N_22969,N_21386);
xnor U26551 (N_26551,N_19830,N_18131);
nor U26552 (N_26552,N_20574,N_18835);
or U26553 (N_26553,N_23211,N_23447);
or U26554 (N_26554,N_20120,N_21487);
nor U26555 (N_26555,N_21260,N_21058);
xor U26556 (N_26556,N_19728,N_22169);
or U26557 (N_26557,N_22598,N_19993);
nor U26558 (N_26558,N_18184,N_23371);
xnor U26559 (N_26559,N_18590,N_23485);
nand U26560 (N_26560,N_22802,N_22477);
and U26561 (N_26561,N_22950,N_22643);
or U26562 (N_26562,N_22213,N_19470);
nor U26563 (N_26563,N_19818,N_18737);
xnor U26564 (N_26564,N_22370,N_21713);
nand U26565 (N_26565,N_20386,N_23714);
xnor U26566 (N_26566,N_18998,N_20223);
nand U26567 (N_26567,N_20609,N_19195);
nor U26568 (N_26568,N_21947,N_20575);
nand U26569 (N_26569,N_23637,N_19021);
xor U26570 (N_26570,N_18818,N_20635);
xor U26571 (N_26571,N_20399,N_20748);
and U26572 (N_26572,N_22278,N_21214);
nand U26573 (N_26573,N_18531,N_22780);
nor U26574 (N_26574,N_22401,N_20462);
nand U26575 (N_26575,N_23014,N_18829);
nor U26576 (N_26576,N_23231,N_21130);
nor U26577 (N_26577,N_22119,N_21014);
nor U26578 (N_26578,N_21661,N_18592);
xnor U26579 (N_26579,N_20662,N_22149);
nor U26580 (N_26580,N_21272,N_21715);
xnor U26581 (N_26581,N_21350,N_18119);
nand U26582 (N_26582,N_19510,N_19526);
nand U26583 (N_26583,N_19519,N_23941);
and U26584 (N_26584,N_21360,N_21660);
or U26585 (N_26585,N_18194,N_18108);
or U26586 (N_26586,N_20200,N_23658);
nand U26587 (N_26587,N_23732,N_18694);
and U26588 (N_26588,N_18093,N_21339);
or U26589 (N_26589,N_21749,N_19012);
or U26590 (N_26590,N_21539,N_22722);
and U26591 (N_26591,N_23200,N_23389);
nand U26592 (N_26592,N_22309,N_23562);
nand U26593 (N_26593,N_19018,N_20106);
nand U26594 (N_26594,N_19848,N_23688);
nand U26595 (N_26595,N_20801,N_19171);
or U26596 (N_26596,N_20547,N_22685);
xnor U26597 (N_26597,N_19585,N_23672);
and U26598 (N_26598,N_22206,N_18803);
xor U26599 (N_26599,N_20688,N_20493);
xor U26600 (N_26600,N_18824,N_20584);
and U26601 (N_26601,N_19780,N_21618);
and U26602 (N_26602,N_21594,N_23003);
nor U26603 (N_26603,N_20303,N_20458);
or U26604 (N_26604,N_19564,N_23607);
xnor U26605 (N_26605,N_23754,N_19524);
nand U26606 (N_26606,N_20852,N_22594);
or U26607 (N_26607,N_18638,N_19963);
and U26608 (N_26608,N_18741,N_20311);
xnor U26609 (N_26609,N_18045,N_22652);
and U26610 (N_26610,N_18954,N_20565);
or U26611 (N_26611,N_23766,N_18989);
and U26612 (N_26612,N_20970,N_21076);
and U26613 (N_26613,N_19341,N_20757);
nand U26614 (N_26614,N_19992,N_19648);
nand U26615 (N_26615,N_19902,N_18250);
xnor U26616 (N_26616,N_18579,N_23805);
or U26617 (N_26617,N_19852,N_23355);
nand U26618 (N_26618,N_23728,N_19368);
xor U26619 (N_26619,N_18500,N_22704);
and U26620 (N_26620,N_22225,N_21668);
nand U26621 (N_26621,N_23604,N_23606);
or U26622 (N_26622,N_23618,N_18913);
or U26623 (N_26623,N_23689,N_22675);
or U26624 (N_26624,N_22105,N_22860);
nand U26625 (N_26625,N_20598,N_23715);
nor U26626 (N_26626,N_23972,N_21166);
nand U26627 (N_26627,N_21638,N_21935);
or U26628 (N_26628,N_18056,N_21399);
nand U26629 (N_26629,N_18523,N_22765);
or U26630 (N_26630,N_23455,N_19651);
or U26631 (N_26631,N_18985,N_18142);
nand U26632 (N_26632,N_18464,N_23577);
and U26633 (N_26633,N_22492,N_23978);
nand U26634 (N_26634,N_19724,N_20159);
or U26635 (N_26635,N_19060,N_23123);
and U26636 (N_26636,N_19931,N_22531);
xor U26637 (N_26637,N_22838,N_22824);
nand U26638 (N_26638,N_19013,N_23854);
and U26639 (N_26639,N_22431,N_23246);
nor U26640 (N_26640,N_20671,N_18357);
or U26641 (N_26641,N_22976,N_22459);
nor U26642 (N_26642,N_22280,N_18769);
nor U26643 (N_26643,N_22991,N_19834);
and U26644 (N_26644,N_21882,N_20957);
and U26645 (N_26645,N_18756,N_18472);
and U26646 (N_26646,N_19877,N_22715);
nor U26647 (N_26647,N_18356,N_20790);
or U26648 (N_26648,N_20780,N_23903);
or U26649 (N_26649,N_19295,N_18261);
nand U26650 (N_26650,N_22409,N_20394);
or U26651 (N_26651,N_22317,N_19219);
xnor U26652 (N_26652,N_23773,N_19077);
or U26653 (N_26653,N_23748,N_18905);
nand U26654 (N_26654,N_19541,N_18175);
xnor U26655 (N_26655,N_19204,N_22318);
xor U26656 (N_26656,N_18254,N_21677);
xnor U26657 (N_26657,N_18233,N_18648);
and U26658 (N_26658,N_19316,N_18600);
nand U26659 (N_26659,N_23016,N_19379);
nand U26660 (N_26660,N_19230,N_19298);
xor U26661 (N_26661,N_19288,N_18435);
nor U26662 (N_26662,N_20590,N_18443);
xnor U26663 (N_26663,N_21157,N_20373);
and U26664 (N_26664,N_23114,N_22092);
or U26665 (N_26665,N_22881,N_18960);
or U26666 (N_26666,N_18932,N_18551);
nor U26667 (N_26667,N_18304,N_22014);
and U26668 (N_26668,N_23350,N_20587);
xor U26669 (N_26669,N_20509,N_21981);
and U26670 (N_26670,N_22501,N_22726);
nand U26671 (N_26671,N_23294,N_22353);
nand U26672 (N_26672,N_18132,N_19996);
nand U26673 (N_26673,N_20883,N_23574);
and U26674 (N_26674,N_20408,N_22470);
and U26675 (N_26675,N_20412,N_23988);
nand U26676 (N_26676,N_23557,N_19147);
nand U26677 (N_26677,N_21141,N_20060);
and U26678 (N_26678,N_23866,N_18242);
nor U26679 (N_26679,N_21364,N_18585);
nand U26680 (N_26680,N_23703,N_21701);
nand U26681 (N_26681,N_20926,N_22196);
nor U26682 (N_26682,N_23725,N_22145);
xnor U26683 (N_26683,N_21168,N_22250);
and U26684 (N_26684,N_18901,N_18710);
xnor U26685 (N_26685,N_22128,N_23624);
nand U26686 (N_26686,N_19130,N_21640);
xnor U26687 (N_26687,N_18692,N_18232);
nor U26688 (N_26688,N_22776,N_22073);
nand U26689 (N_26689,N_22545,N_18310);
nand U26690 (N_26690,N_21591,N_19870);
nand U26691 (N_26691,N_22010,N_20151);
and U26692 (N_26692,N_20278,N_23069);
and U26693 (N_26693,N_20861,N_20550);
nor U26694 (N_26694,N_18268,N_19606);
or U26695 (N_26695,N_19249,N_18294);
nor U26696 (N_26696,N_19713,N_20733);
xnor U26697 (N_26697,N_22184,N_19795);
and U26698 (N_26698,N_21381,N_20267);
nor U26699 (N_26699,N_23134,N_19991);
xnor U26700 (N_26700,N_19865,N_19819);
nor U26701 (N_26701,N_21969,N_22214);
nor U26702 (N_26702,N_23250,N_20652);
xnor U26703 (N_26703,N_23882,N_21104);
nor U26704 (N_26704,N_23582,N_23358);
nand U26705 (N_26705,N_18425,N_22610);
xnor U26706 (N_26706,N_23706,N_19736);
nor U26707 (N_26707,N_23515,N_18281);
nand U26708 (N_26708,N_22427,N_19072);
and U26709 (N_26709,N_22788,N_22512);
xor U26710 (N_26710,N_20567,N_21207);
nor U26711 (N_26711,N_22000,N_23827);
and U26712 (N_26712,N_20655,N_23079);
xor U26713 (N_26713,N_23786,N_19806);
and U26714 (N_26714,N_21443,N_21284);
nand U26715 (N_26715,N_19733,N_18856);
or U26716 (N_26716,N_18859,N_22854);
xnor U26717 (N_26717,N_18680,N_19192);
nand U26718 (N_26718,N_19293,N_22559);
nor U26719 (N_26719,N_22628,N_23868);
nand U26720 (N_26720,N_22493,N_21128);
nor U26721 (N_26721,N_20673,N_22024);
xor U26722 (N_26722,N_23818,N_19425);
nand U26723 (N_26723,N_21820,N_19857);
nor U26724 (N_26724,N_22568,N_22882);
or U26725 (N_26725,N_21042,N_19153);
xnor U26726 (N_26726,N_18345,N_21938);
and U26727 (N_26727,N_19672,N_23631);
nand U26728 (N_26728,N_21135,N_21906);
nand U26729 (N_26729,N_21682,N_22505);
and U26730 (N_26730,N_18147,N_20068);
nand U26731 (N_26731,N_19914,N_18684);
and U26732 (N_26732,N_22106,N_23617);
xnor U26733 (N_26733,N_23946,N_18618);
or U26734 (N_26734,N_22601,N_23572);
nor U26735 (N_26735,N_19777,N_18041);
xor U26736 (N_26736,N_18167,N_23232);
xnor U26737 (N_26737,N_23464,N_20874);
nand U26738 (N_26738,N_18708,N_21798);
and U26739 (N_26739,N_19170,N_22360);
xor U26740 (N_26740,N_20283,N_21711);
nor U26741 (N_26741,N_22331,N_23863);
nor U26742 (N_26742,N_22113,N_19753);
or U26743 (N_26743,N_20703,N_19063);
and U26744 (N_26744,N_21041,N_18889);
and U26745 (N_26745,N_21953,N_20517);
and U26746 (N_26746,N_21019,N_22638);
xnor U26747 (N_26747,N_21258,N_20253);
or U26748 (N_26748,N_20890,N_21028);
and U26749 (N_26749,N_23173,N_20570);
or U26750 (N_26750,N_20464,N_18729);
nor U26751 (N_26751,N_23643,N_20934);
xor U26752 (N_26752,N_18751,N_23007);
nor U26753 (N_26753,N_18475,N_19105);
xor U26754 (N_26754,N_23611,N_23479);
xnor U26755 (N_26755,N_18833,N_23530);
nand U26756 (N_26756,N_21092,N_21684);
or U26757 (N_26757,N_21522,N_21993);
nor U26758 (N_26758,N_21371,N_18105);
and U26759 (N_26759,N_23061,N_23670);
nand U26760 (N_26760,N_20772,N_18365);
and U26761 (N_26761,N_23493,N_22627);
or U26762 (N_26762,N_20323,N_22939);
nor U26763 (N_26763,N_23247,N_19891);
nand U26764 (N_26764,N_23392,N_20515);
xnor U26765 (N_26765,N_23164,N_19136);
and U26766 (N_26766,N_18015,N_18614);
or U26767 (N_26767,N_18270,N_18685);
and U26768 (N_26768,N_19161,N_22832);
or U26769 (N_26769,N_19613,N_19290);
nand U26770 (N_26770,N_22450,N_23546);
nor U26771 (N_26771,N_20369,N_18381);
nor U26772 (N_26772,N_18411,N_23298);
and U26773 (N_26773,N_23025,N_22721);
xnor U26774 (N_26774,N_21340,N_18069);
nand U26775 (N_26775,N_23437,N_19875);
and U26776 (N_26776,N_20732,N_22856);
nor U26777 (N_26777,N_20185,N_20315);
and U26778 (N_26778,N_18337,N_19689);
nor U26779 (N_26779,N_22719,N_19698);
nand U26780 (N_26780,N_19381,N_20840);
nor U26781 (N_26781,N_23625,N_20612);
or U26782 (N_26782,N_18981,N_18622);
nor U26783 (N_26783,N_22351,N_19782);
and U26784 (N_26784,N_23206,N_20786);
and U26785 (N_26785,N_18306,N_22551);
or U26786 (N_26786,N_20032,N_23031);
nor U26787 (N_26787,N_18317,N_22982);
or U26788 (N_26788,N_18135,N_19508);
nor U26789 (N_26789,N_23450,N_18846);
nor U26790 (N_26790,N_23870,N_19989);
and U26791 (N_26791,N_19044,N_18665);
nand U26792 (N_26792,N_21936,N_22983);
or U26793 (N_26793,N_19623,N_21404);
nand U26794 (N_26794,N_18564,N_19074);
nand U26795 (N_26795,N_23017,N_20411);
or U26796 (N_26796,N_20879,N_22670);
nand U26797 (N_26797,N_23724,N_22323);
and U26798 (N_26798,N_19262,N_20341);
nand U26799 (N_26799,N_23269,N_18121);
xor U26800 (N_26800,N_20187,N_22764);
nor U26801 (N_26801,N_18693,N_18300);
nand U26802 (N_26802,N_20514,N_19203);
xor U26803 (N_26803,N_21630,N_23749);
and U26804 (N_26804,N_18919,N_21062);
xor U26805 (N_26805,N_21456,N_20168);
and U26806 (N_26806,N_23694,N_20918);
nand U26807 (N_26807,N_18129,N_22910);
and U26808 (N_26808,N_18702,N_19647);
nor U26809 (N_26809,N_23175,N_18778);
xor U26810 (N_26810,N_23086,N_19760);
nand U26811 (N_26811,N_23659,N_19218);
xor U26812 (N_26812,N_18070,N_19810);
nand U26813 (N_26813,N_18185,N_22867);
and U26814 (N_26814,N_23207,N_20636);
nand U26815 (N_26815,N_22308,N_18220);
or U26816 (N_26816,N_20971,N_18661);
or U26817 (N_26817,N_18844,N_19831);
and U26818 (N_26818,N_23723,N_19657);
xor U26819 (N_26819,N_21497,N_23852);
and U26820 (N_26820,N_21653,N_21216);
xnor U26821 (N_26821,N_22298,N_21079);
xnor U26822 (N_26822,N_22392,N_23849);
nand U26823 (N_26823,N_20775,N_21422);
xnor U26824 (N_26824,N_20793,N_21649);
nand U26825 (N_26825,N_22992,N_18245);
and U26826 (N_26826,N_18534,N_20195);
and U26827 (N_26827,N_19223,N_21145);
and U26828 (N_26828,N_23884,N_21044);
nand U26829 (N_26829,N_21349,N_23601);
or U26830 (N_26830,N_19529,N_18810);
and U26831 (N_26831,N_21867,N_19444);
nand U26832 (N_26832,N_23739,N_18400);
or U26833 (N_26833,N_23918,N_18716);
and U26834 (N_26834,N_23074,N_22946);
or U26835 (N_26835,N_23568,N_23382);
and U26836 (N_26836,N_23004,N_20225);
nor U26837 (N_26837,N_22527,N_22593);
and U26838 (N_26838,N_20161,N_19370);
nand U26839 (N_26839,N_19182,N_22491);
nor U26840 (N_26840,N_19184,N_21064);
xnor U26841 (N_26841,N_22363,N_23596);
nor U26842 (N_26842,N_20190,N_22956);
or U26843 (N_26843,N_19152,N_21804);
nor U26844 (N_26844,N_23095,N_22046);
nor U26845 (N_26845,N_19362,N_19177);
and U26846 (N_26846,N_21473,N_20299);
or U26847 (N_26847,N_22743,N_23210);
xor U26848 (N_26848,N_19903,N_21204);
or U26849 (N_26849,N_23842,N_23944);
nor U26850 (N_26850,N_19007,N_23275);
or U26851 (N_26851,N_20588,N_22529);
and U26852 (N_26852,N_19448,N_22116);
and U26853 (N_26853,N_20079,N_19889);
xnor U26854 (N_26854,N_18983,N_20222);
and U26855 (N_26855,N_23505,N_18113);
nor U26856 (N_26856,N_18226,N_23838);
nor U26857 (N_26857,N_19045,N_19920);
nand U26858 (N_26858,N_21393,N_19908);
nor U26859 (N_26859,N_21864,N_19859);
xor U26860 (N_26860,N_23300,N_21837);
or U26861 (N_26861,N_23745,N_19493);
or U26862 (N_26862,N_19092,N_18054);
or U26863 (N_26863,N_20982,N_20028);
nand U26864 (N_26864,N_23005,N_23547);
and U26865 (N_26865,N_19208,N_18082);
and U26866 (N_26866,N_18921,N_22706);
nand U26867 (N_26867,N_19106,N_18010);
xor U26868 (N_26868,N_20246,N_23666);
and U26869 (N_26869,N_19814,N_18791);
nor U26870 (N_26870,N_22817,N_22087);
nand U26871 (N_26871,N_22352,N_21174);
nand U26872 (N_26872,N_19534,N_19442);
or U26873 (N_26873,N_18720,N_18333);
and U26874 (N_26874,N_18792,N_19888);
xnor U26875 (N_26875,N_18822,N_23481);
or U26876 (N_26876,N_19946,N_19714);
and U26877 (N_26877,N_20991,N_21878);
or U26878 (N_26878,N_20911,N_23931);
nand U26879 (N_26879,N_18934,N_21446);
nand U26880 (N_26880,N_20522,N_23959);
or U26881 (N_26881,N_22139,N_22987);
xnor U26882 (N_26882,N_21441,N_21276);
nand U26883 (N_26883,N_19943,N_23240);
nor U26884 (N_26884,N_23439,N_20661);
and U26885 (N_26885,N_22596,N_23822);
xnor U26886 (N_26886,N_21560,N_18355);
xnor U26887 (N_26887,N_20964,N_22221);
nor U26888 (N_26888,N_23532,N_19540);
or U26889 (N_26889,N_19968,N_23632);
nand U26890 (N_26890,N_22339,N_21813);
xnor U26891 (N_26891,N_19809,N_23738);
xor U26892 (N_26892,N_21342,N_22474);
and U26893 (N_26893,N_21809,N_18415);
nand U26894 (N_26894,N_18324,N_22819);
nand U26895 (N_26895,N_19948,N_23489);
nand U26896 (N_26896,N_19066,N_20291);
nand U26897 (N_26897,N_23425,N_20269);
and U26898 (N_26898,N_18772,N_19047);
xor U26899 (N_26899,N_19545,N_22321);
nor U26900 (N_26900,N_22041,N_20209);
or U26901 (N_26901,N_22821,N_19364);
xnor U26902 (N_26902,N_20404,N_21278);
and U26903 (N_26903,N_23709,N_20127);
xnor U26904 (N_26904,N_20017,N_20279);
or U26905 (N_26905,N_21030,N_19980);
xnor U26906 (N_26906,N_21098,N_20289);
nand U26907 (N_26907,N_21085,N_23511);
nor U26908 (N_26908,N_20896,N_19251);
and U26909 (N_26909,N_21945,N_19433);
nor U26910 (N_26910,N_19446,N_18705);
nand U26911 (N_26911,N_18744,N_20543);
nor U26912 (N_26912,N_23829,N_23860);
nand U26913 (N_26913,N_18405,N_20110);
nor U26914 (N_26914,N_19174,N_22437);
or U26915 (N_26915,N_21280,N_23872);
nor U26916 (N_26916,N_23667,N_20175);
nor U26917 (N_26917,N_22751,N_22499);
and U26918 (N_26918,N_19873,N_19614);
nand U26919 (N_26919,N_22208,N_19787);
and U26920 (N_26920,N_19339,N_23304);
or U26921 (N_26921,N_20426,N_21975);
nor U26922 (N_26922,N_21762,N_22774);
or U26923 (N_26923,N_23710,N_18507);
xnor U26924 (N_26924,N_22635,N_19986);
and U26925 (N_26925,N_20819,N_18432);
xor U26926 (N_26926,N_22519,N_18621);
or U26927 (N_26927,N_19097,N_22809);
or U26928 (N_26928,N_19307,N_18018);
nand U26929 (N_26929,N_19578,N_19061);
nor U26930 (N_26930,N_21299,N_23544);
nor U26931 (N_26931,N_19868,N_21306);
nand U26932 (N_26932,N_23968,N_22507);
nor U26933 (N_26933,N_22578,N_18376);
nand U26934 (N_26934,N_20219,N_20116);
and U26935 (N_26935,N_23293,N_23140);
and U26936 (N_26936,N_23915,N_21029);
and U26937 (N_26937,N_23979,N_23997);
or U26938 (N_26938,N_20486,N_20749);
or U26939 (N_26939,N_18318,N_19133);
and U26940 (N_26940,N_18224,N_19973);
or U26941 (N_26941,N_23374,N_19280);
or U26942 (N_26942,N_18502,N_21313);
nor U26943 (N_26943,N_20231,N_20221);
or U26944 (N_26944,N_18874,N_21163);
xor U26945 (N_26945,N_19559,N_23019);
xor U26946 (N_26946,N_23020,N_23202);
xnor U26947 (N_26947,N_22739,N_23845);
and U26948 (N_26948,N_22248,N_20383);
and U26949 (N_26949,N_23928,N_20372);
xor U26950 (N_26950,N_21960,N_20039);
xor U26951 (N_26951,N_20809,N_20302);
and U26952 (N_26952,N_20465,N_22283);
or U26953 (N_26953,N_23911,N_18973);
xor U26954 (N_26954,N_20546,N_19699);
xnor U26955 (N_26955,N_20206,N_22216);
and U26956 (N_26956,N_23986,N_23965);
nor U26957 (N_26957,N_20217,N_20788);
xor U26958 (N_26958,N_23154,N_20208);
xnor U26959 (N_26959,N_19083,N_18554);
xnor U26960 (N_26960,N_21086,N_21305);
and U26961 (N_26961,N_18924,N_20650);
nand U26962 (N_26962,N_20919,N_18886);
nand U26963 (N_26963,N_19451,N_19435);
nand U26964 (N_26964,N_23215,N_18654);
nand U26965 (N_26965,N_18038,N_21348);
xnor U26966 (N_26966,N_21679,N_18342);
nor U26967 (N_26967,N_21552,N_23354);
and U26968 (N_26968,N_21833,N_20111);
xor U26969 (N_26969,N_20618,N_23407);
or U26970 (N_26970,N_22151,N_19308);
or U26971 (N_26971,N_23209,N_22175);
and U26972 (N_26972,N_18848,N_19553);
or U26973 (N_26973,N_18343,N_19666);
or U26974 (N_26974,N_18704,N_18980);
or U26975 (N_26975,N_22154,N_21739);
and U26976 (N_26976,N_21262,N_23804);
nor U26977 (N_26977,N_20337,N_21081);
xor U26978 (N_26978,N_19756,N_21574);
nand U26979 (N_26979,N_19620,N_18709);
nand U26980 (N_26980,N_22337,N_22295);
xnor U26981 (N_26981,N_23698,N_21513);
nand U26982 (N_26982,N_21490,N_21463);
xor U26983 (N_26983,N_23197,N_19634);
or U26984 (N_26984,N_23994,N_23299);
or U26985 (N_26985,N_20593,N_19465);
and U26986 (N_26986,N_20885,N_20164);
and U26987 (N_26987,N_21485,N_21372);
xor U26988 (N_26988,N_22813,N_18867);
or U26989 (N_26989,N_18009,N_19855);
nand U26990 (N_26990,N_18779,N_22011);
and U26991 (N_26991,N_18017,N_21900);
nand U26992 (N_26992,N_19972,N_19523);
nand U26993 (N_26993,N_20833,N_22700);
xor U26994 (N_26994,N_18794,N_23491);
nor U26995 (N_26995,N_22183,N_22857);
xnor U26996 (N_26996,N_19022,N_21581);
xor U26997 (N_26997,N_20735,N_21046);
or U26998 (N_26998,N_21621,N_23129);
and U26999 (N_26999,N_18735,N_20392);
and U27000 (N_27000,N_21962,N_19627);
xnor U27001 (N_27001,N_21145,N_18623);
xor U27002 (N_27002,N_23773,N_18624);
and U27003 (N_27003,N_20379,N_21277);
or U27004 (N_27004,N_23625,N_18941);
or U27005 (N_27005,N_18843,N_20062);
xnor U27006 (N_27006,N_22015,N_20330);
nor U27007 (N_27007,N_18569,N_21252);
or U27008 (N_27008,N_19819,N_23869);
nand U27009 (N_27009,N_21863,N_23511);
or U27010 (N_27010,N_21430,N_21758);
and U27011 (N_27011,N_22639,N_20190);
nor U27012 (N_27012,N_22858,N_19695);
and U27013 (N_27013,N_20732,N_18704);
nand U27014 (N_27014,N_22603,N_18095);
or U27015 (N_27015,N_18734,N_19528);
or U27016 (N_27016,N_18075,N_21064);
and U27017 (N_27017,N_23148,N_20402);
nand U27018 (N_27018,N_23701,N_23613);
or U27019 (N_27019,N_20118,N_23807);
nand U27020 (N_27020,N_21854,N_22622);
nor U27021 (N_27021,N_23579,N_19008);
and U27022 (N_27022,N_19046,N_21131);
nor U27023 (N_27023,N_23901,N_22252);
or U27024 (N_27024,N_20108,N_18786);
nand U27025 (N_27025,N_23068,N_21548);
nand U27026 (N_27026,N_20106,N_20022);
nor U27027 (N_27027,N_21605,N_19231);
nand U27028 (N_27028,N_22502,N_21797);
nor U27029 (N_27029,N_19324,N_22121);
or U27030 (N_27030,N_19257,N_23157);
nor U27031 (N_27031,N_19696,N_22870);
xor U27032 (N_27032,N_23011,N_21446);
nand U27033 (N_27033,N_19224,N_19088);
nand U27034 (N_27034,N_21630,N_22448);
nor U27035 (N_27035,N_19613,N_23585);
or U27036 (N_27036,N_19796,N_20707);
or U27037 (N_27037,N_22090,N_18073);
or U27038 (N_27038,N_22315,N_20751);
nand U27039 (N_27039,N_23830,N_18159);
xnor U27040 (N_27040,N_21147,N_18219);
or U27041 (N_27041,N_21323,N_22850);
nand U27042 (N_27042,N_18457,N_21030);
or U27043 (N_27043,N_18790,N_22013);
nand U27044 (N_27044,N_22368,N_20365);
or U27045 (N_27045,N_19576,N_22480);
and U27046 (N_27046,N_22079,N_20533);
nor U27047 (N_27047,N_22313,N_18007);
xnor U27048 (N_27048,N_20049,N_21940);
nor U27049 (N_27049,N_19870,N_18461);
or U27050 (N_27050,N_21209,N_19024);
and U27051 (N_27051,N_23909,N_18583);
nand U27052 (N_27052,N_21928,N_21812);
xor U27053 (N_27053,N_22063,N_22406);
nor U27054 (N_27054,N_20738,N_22497);
or U27055 (N_27055,N_23296,N_19141);
xnor U27056 (N_27056,N_19346,N_21617);
and U27057 (N_27057,N_21251,N_18379);
xor U27058 (N_27058,N_19566,N_21583);
nor U27059 (N_27059,N_21200,N_18619);
nor U27060 (N_27060,N_23521,N_23485);
or U27061 (N_27061,N_19527,N_18677);
nor U27062 (N_27062,N_21500,N_19823);
and U27063 (N_27063,N_22558,N_22466);
nor U27064 (N_27064,N_20251,N_18587);
xor U27065 (N_27065,N_18294,N_23423);
or U27066 (N_27066,N_23371,N_21161);
xnor U27067 (N_27067,N_21338,N_19263);
and U27068 (N_27068,N_21112,N_19635);
or U27069 (N_27069,N_22980,N_19094);
and U27070 (N_27070,N_21019,N_18946);
or U27071 (N_27071,N_20682,N_21512);
or U27072 (N_27072,N_19745,N_19507);
nand U27073 (N_27073,N_22746,N_23405);
or U27074 (N_27074,N_23935,N_18886);
nand U27075 (N_27075,N_19448,N_23766);
nand U27076 (N_27076,N_22270,N_23657);
and U27077 (N_27077,N_22236,N_18539);
nor U27078 (N_27078,N_21381,N_23772);
xor U27079 (N_27079,N_22597,N_18605);
or U27080 (N_27080,N_22204,N_20511);
nand U27081 (N_27081,N_23203,N_20651);
nor U27082 (N_27082,N_20181,N_23213);
nor U27083 (N_27083,N_20118,N_22951);
nand U27084 (N_27084,N_18653,N_22990);
xnor U27085 (N_27085,N_18770,N_22261);
or U27086 (N_27086,N_21250,N_21564);
nor U27087 (N_27087,N_20900,N_20678);
and U27088 (N_27088,N_22513,N_23992);
nor U27089 (N_27089,N_22231,N_20925);
and U27090 (N_27090,N_18591,N_23890);
nor U27091 (N_27091,N_19662,N_22846);
xor U27092 (N_27092,N_18009,N_18632);
nand U27093 (N_27093,N_19221,N_18922);
nand U27094 (N_27094,N_20498,N_23008);
nor U27095 (N_27095,N_23901,N_22589);
nand U27096 (N_27096,N_20411,N_20540);
and U27097 (N_27097,N_20454,N_21568);
xnor U27098 (N_27098,N_21821,N_22229);
nor U27099 (N_27099,N_19656,N_19691);
xor U27100 (N_27100,N_18270,N_23993);
and U27101 (N_27101,N_23043,N_23903);
or U27102 (N_27102,N_19926,N_22165);
nor U27103 (N_27103,N_18483,N_21067);
nand U27104 (N_27104,N_18572,N_23761);
and U27105 (N_27105,N_21049,N_20911);
nor U27106 (N_27106,N_23657,N_20526);
xor U27107 (N_27107,N_19216,N_18649);
nor U27108 (N_27108,N_22277,N_19326);
nor U27109 (N_27109,N_21349,N_19446);
xor U27110 (N_27110,N_20086,N_22902);
or U27111 (N_27111,N_20760,N_18853);
nor U27112 (N_27112,N_23436,N_20589);
xor U27113 (N_27113,N_19557,N_20633);
or U27114 (N_27114,N_20477,N_21326);
nand U27115 (N_27115,N_22618,N_22802);
and U27116 (N_27116,N_22782,N_23122);
xnor U27117 (N_27117,N_20156,N_22894);
nor U27118 (N_27118,N_18703,N_23995);
or U27119 (N_27119,N_21052,N_23656);
and U27120 (N_27120,N_19001,N_18776);
xor U27121 (N_27121,N_22279,N_21660);
or U27122 (N_27122,N_18976,N_21983);
nand U27123 (N_27123,N_21767,N_18045);
nor U27124 (N_27124,N_21761,N_19473);
nand U27125 (N_27125,N_19504,N_22303);
xnor U27126 (N_27126,N_18213,N_23763);
and U27127 (N_27127,N_21997,N_20073);
nand U27128 (N_27128,N_23659,N_20071);
nand U27129 (N_27129,N_20155,N_23344);
xnor U27130 (N_27130,N_23287,N_18805);
and U27131 (N_27131,N_21202,N_19398);
or U27132 (N_27132,N_22108,N_21822);
and U27133 (N_27133,N_21153,N_18496);
or U27134 (N_27134,N_18137,N_21420);
or U27135 (N_27135,N_22881,N_22621);
xnor U27136 (N_27136,N_22191,N_22682);
xor U27137 (N_27137,N_22682,N_21251);
and U27138 (N_27138,N_19709,N_21013);
nor U27139 (N_27139,N_23030,N_18844);
or U27140 (N_27140,N_18692,N_18038);
nor U27141 (N_27141,N_23018,N_20770);
or U27142 (N_27142,N_22528,N_18743);
or U27143 (N_27143,N_21005,N_23057);
nor U27144 (N_27144,N_21610,N_18915);
xor U27145 (N_27145,N_21850,N_21837);
or U27146 (N_27146,N_23829,N_21759);
nor U27147 (N_27147,N_19409,N_23611);
nand U27148 (N_27148,N_21265,N_21882);
and U27149 (N_27149,N_20260,N_22250);
and U27150 (N_27150,N_19014,N_19372);
xnor U27151 (N_27151,N_18477,N_19219);
and U27152 (N_27152,N_20244,N_18216);
nor U27153 (N_27153,N_22752,N_22460);
and U27154 (N_27154,N_18387,N_21308);
and U27155 (N_27155,N_21817,N_19578);
or U27156 (N_27156,N_23964,N_22873);
and U27157 (N_27157,N_18912,N_22215);
nor U27158 (N_27158,N_19643,N_23043);
nor U27159 (N_27159,N_19263,N_23700);
or U27160 (N_27160,N_21473,N_19086);
or U27161 (N_27161,N_18155,N_22896);
xor U27162 (N_27162,N_22748,N_21479);
and U27163 (N_27163,N_20196,N_18061);
or U27164 (N_27164,N_23711,N_21073);
or U27165 (N_27165,N_21125,N_20726);
nand U27166 (N_27166,N_19382,N_20657);
and U27167 (N_27167,N_21240,N_23977);
and U27168 (N_27168,N_21353,N_18281);
nand U27169 (N_27169,N_20255,N_20527);
or U27170 (N_27170,N_23366,N_22677);
nand U27171 (N_27171,N_20732,N_18930);
and U27172 (N_27172,N_21445,N_21314);
xor U27173 (N_27173,N_18001,N_21929);
nor U27174 (N_27174,N_23885,N_18213);
nand U27175 (N_27175,N_19917,N_19652);
nand U27176 (N_27176,N_20012,N_18732);
and U27177 (N_27177,N_19716,N_19867);
and U27178 (N_27178,N_19113,N_23845);
nand U27179 (N_27179,N_18054,N_18560);
nand U27180 (N_27180,N_23109,N_22424);
and U27181 (N_27181,N_18833,N_18654);
or U27182 (N_27182,N_19448,N_23003);
or U27183 (N_27183,N_18327,N_19080);
nor U27184 (N_27184,N_19314,N_20119);
or U27185 (N_27185,N_19758,N_23588);
xor U27186 (N_27186,N_23806,N_22792);
nand U27187 (N_27187,N_19835,N_23279);
nand U27188 (N_27188,N_22310,N_23175);
and U27189 (N_27189,N_18554,N_20111);
nor U27190 (N_27190,N_18833,N_19398);
and U27191 (N_27191,N_20043,N_22874);
nor U27192 (N_27192,N_21896,N_21575);
nand U27193 (N_27193,N_18408,N_19313);
nand U27194 (N_27194,N_19001,N_21404);
nand U27195 (N_27195,N_23607,N_21599);
nor U27196 (N_27196,N_23410,N_20201);
nor U27197 (N_27197,N_19856,N_18654);
nor U27198 (N_27198,N_22344,N_21725);
xor U27199 (N_27199,N_21564,N_18220);
nor U27200 (N_27200,N_21850,N_23454);
or U27201 (N_27201,N_22150,N_20831);
nand U27202 (N_27202,N_21212,N_19234);
nand U27203 (N_27203,N_19066,N_20599);
xnor U27204 (N_27204,N_22422,N_21992);
nor U27205 (N_27205,N_18182,N_19929);
xor U27206 (N_27206,N_21585,N_21046);
nand U27207 (N_27207,N_21381,N_21955);
and U27208 (N_27208,N_19135,N_19320);
nor U27209 (N_27209,N_19220,N_23619);
xor U27210 (N_27210,N_21329,N_18611);
xnor U27211 (N_27211,N_23502,N_19577);
and U27212 (N_27212,N_21308,N_21379);
and U27213 (N_27213,N_22854,N_18457);
nor U27214 (N_27214,N_18366,N_18448);
xor U27215 (N_27215,N_23762,N_21673);
nor U27216 (N_27216,N_22498,N_21660);
or U27217 (N_27217,N_21687,N_22555);
nand U27218 (N_27218,N_19186,N_21334);
and U27219 (N_27219,N_20505,N_23111);
and U27220 (N_27220,N_22655,N_23765);
nor U27221 (N_27221,N_20944,N_21972);
nand U27222 (N_27222,N_20433,N_21503);
and U27223 (N_27223,N_19989,N_22231);
nor U27224 (N_27224,N_19185,N_22811);
or U27225 (N_27225,N_19841,N_21707);
xor U27226 (N_27226,N_19197,N_18915);
xnor U27227 (N_27227,N_22220,N_19083);
and U27228 (N_27228,N_23580,N_18129);
xor U27229 (N_27229,N_18349,N_21472);
and U27230 (N_27230,N_18988,N_19859);
xnor U27231 (N_27231,N_21127,N_21324);
xnor U27232 (N_27232,N_20976,N_21328);
xnor U27233 (N_27233,N_21952,N_21886);
nor U27234 (N_27234,N_19733,N_19439);
nand U27235 (N_27235,N_18231,N_22390);
nand U27236 (N_27236,N_21227,N_20024);
nor U27237 (N_27237,N_21495,N_23584);
and U27238 (N_27238,N_19577,N_23109);
nand U27239 (N_27239,N_22819,N_18260);
or U27240 (N_27240,N_20357,N_21313);
or U27241 (N_27241,N_22419,N_20566);
nor U27242 (N_27242,N_21009,N_23424);
and U27243 (N_27243,N_20037,N_22494);
and U27244 (N_27244,N_18330,N_20795);
nand U27245 (N_27245,N_23901,N_19097);
nor U27246 (N_27246,N_19720,N_23859);
nor U27247 (N_27247,N_21116,N_19266);
nand U27248 (N_27248,N_19587,N_18448);
xnor U27249 (N_27249,N_18648,N_22157);
nand U27250 (N_27250,N_18135,N_22077);
xor U27251 (N_27251,N_23410,N_21533);
or U27252 (N_27252,N_21943,N_21750);
or U27253 (N_27253,N_18747,N_20944);
nor U27254 (N_27254,N_23662,N_21598);
and U27255 (N_27255,N_19753,N_21035);
xor U27256 (N_27256,N_18822,N_19609);
xor U27257 (N_27257,N_21828,N_21710);
xor U27258 (N_27258,N_19250,N_20409);
and U27259 (N_27259,N_20813,N_19892);
nor U27260 (N_27260,N_23811,N_19391);
nand U27261 (N_27261,N_18426,N_22786);
nor U27262 (N_27262,N_22738,N_19353);
xnor U27263 (N_27263,N_18252,N_20807);
and U27264 (N_27264,N_18221,N_21816);
nor U27265 (N_27265,N_23054,N_21240);
nor U27266 (N_27266,N_18138,N_19699);
xnor U27267 (N_27267,N_20093,N_19359);
xnor U27268 (N_27268,N_22218,N_18059);
and U27269 (N_27269,N_19621,N_20544);
nor U27270 (N_27270,N_23065,N_22149);
or U27271 (N_27271,N_23084,N_23440);
or U27272 (N_27272,N_18951,N_22678);
nor U27273 (N_27273,N_19562,N_22634);
or U27274 (N_27274,N_23695,N_21462);
or U27275 (N_27275,N_22661,N_20973);
and U27276 (N_27276,N_21508,N_18383);
xnor U27277 (N_27277,N_21717,N_18866);
nor U27278 (N_27278,N_18409,N_22907);
and U27279 (N_27279,N_19209,N_19334);
or U27280 (N_27280,N_23295,N_22493);
and U27281 (N_27281,N_22458,N_23291);
nand U27282 (N_27282,N_18764,N_19706);
nor U27283 (N_27283,N_23462,N_19821);
nor U27284 (N_27284,N_18897,N_18438);
nor U27285 (N_27285,N_20757,N_20703);
or U27286 (N_27286,N_20940,N_22243);
nor U27287 (N_27287,N_22461,N_21514);
nand U27288 (N_27288,N_18553,N_20191);
xor U27289 (N_27289,N_18518,N_23497);
or U27290 (N_27290,N_20946,N_23138);
or U27291 (N_27291,N_20026,N_22009);
and U27292 (N_27292,N_18117,N_19460);
nor U27293 (N_27293,N_23895,N_22002);
nor U27294 (N_27294,N_23700,N_22386);
nor U27295 (N_27295,N_22759,N_19594);
nor U27296 (N_27296,N_22017,N_23314);
nor U27297 (N_27297,N_22427,N_19403);
or U27298 (N_27298,N_22913,N_18000);
nand U27299 (N_27299,N_23963,N_21609);
or U27300 (N_27300,N_21650,N_18375);
and U27301 (N_27301,N_22274,N_20843);
and U27302 (N_27302,N_21362,N_22643);
xor U27303 (N_27303,N_21212,N_22178);
or U27304 (N_27304,N_18313,N_18059);
xnor U27305 (N_27305,N_21982,N_23321);
or U27306 (N_27306,N_21000,N_23034);
or U27307 (N_27307,N_21578,N_23528);
xnor U27308 (N_27308,N_19691,N_18780);
or U27309 (N_27309,N_19392,N_20046);
and U27310 (N_27310,N_21066,N_23446);
or U27311 (N_27311,N_23377,N_20428);
nand U27312 (N_27312,N_22033,N_22340);
xor U27313 (N_27313,N_23553,N_22836);
and U27314 (N_27314,N_19163,N_23417);
and U27315 (N_27315,N_22322,N_23699);
or U27316 (N_27316,N_20198,N_22091);
nand U27317 (N_27317,N_19336,N_19862);
nand U27318 (N_27318,N_21988,N_21546);
or U27319 (N_27319,N_20581,N_22132);
xnor U27320 (N_27320,N_23452,N_21057);
nand U27321 (N_27321,N_23492,N_18961);
nor U27322 (N_27322,N_23415,N_23315);
xor U27323 (N_27323,N_21562,N_23852);
or U27324 (N_27324,N_18230,N_23722);
nor U27325 (N_27325,N_22698,N_22439);
nor U27326 (N_27326,N_21475,N_23279);
and U27327 (N_27327,N_21754,N_22346);
xnor U27328 (N_27328,N_20135,N_19357);
xor U27329 (N_27329,N_19312,N_23528);
nand U27330 (N_27330,N_20991,N_23902);
nand U27331 (N_27331,N_18670,N_23531);
or U27332 (N_27332,N_22096,N_23459);
nor U27333 (N_27333,N_19879,N_21391);
or U27334 (N_27334,N_18636,N_18668);
or U27335 (N_27335,N_20866,N_19905);
nand U27336 (N_27336,N_22700,N_21323);
nor U27337 (N_27337,N_18229,N_23770);
or U27338 (N_27338,N_20000,N_22202);
nor U27339 (N_27339,N_21021,N_20502);
nor U27340 (N_27340,N_18659,N_23259);
nor U27341 (N_27341,N_23372,N_22758);
nand U27342 (N_27342,N_20624,N_20183);
nor U27343 (N_27343,N_22317,N_22374);
and U27344 (N_27344,N_18948,N_21537);
and U27345 (N_27345,N_20800,N_20971);
nor U27346 (N_27346,N_19450,N_22479);
nand U27347 (N_27347,N_22172,N_21198);
nor U27348 (N_27348,N_23431,N_23016);
or U27349 (N_27349,N_20654,N_23384);
nand U27350 (N_27350,N_19736,N_23747);
xnor U27351 (N_27351,N_19661,N_18222);
xnor U27352 (N_27352,N_18599,N_19158);
nand U27353 (N_27353,N_23004,N_18503);
nand U27354 (N_27354,N_19813,N_22078);
xor U27355 (N_27355,N_18426,N_19831);
nor U27356 (N_27356,N_18262,N_18029);
nor U27357 (N_27357,N_21646,N_20561);
or U27358 (N_27358,N_23608,N_19930);
nand U27359 (N_27359,N_23552,N_18630);
nor U27360 (N_27360,N_22748,N_22846);
and U27361 (N_27361,N_20711,N_23087);
nand U27362 (N_27362,N_22769,N_23943);
or U27363 (N_27363,N_19082,N_19620);
nand U27364 (N_27364,N_22306,N_23187);
nand U27365 (N_27365,N_19991,N_21052);
and U27366 (N_27366,N_23310,N_21966);
and U27367 (N_27367,N_19714,N_21062);
nand U27368 (N_27368,N_20781,N_19259);
xor U27369 (N_27369,N_22073,N_23988);
and U27370 (N_27370,N_20629,N_23578);
nor U27371 (N_27371,N_23692,N_18736);
or U27372 (N_27372,N_19940,N_22669);
nor U27373 (N_27373,N_23808,N_22907);
nor U27374 (N_27374,N_19343,N_21913);
xor U27375 (N_27375,N_20272,N_19326);
and U27376 (N_27376,N_19458,N_23549);
and U27377 (N_27377,N_20602,N_21517);
and U27378 (N_27378,N_20863,N_20065);
nand U27379 (N_27379,N_22479,N_23521);
and U27380 (N_27380,N_23964,N_20440);
or U27381 (N_27381,N_18969,N_22118);
and U27382 (N_27382,N_21221,N_21837);
or U27383 (N_27383,N_22451,N_19995);
xor U27384 (N_27384,N_20134,N_19280);
xor U27385 (N_27385,N_19165,N_18505);
or U27386 (N_27386,N_19826,N_18491);
nor U27387 (N_27387,N_21459,N_18418);
nand U27388 (N_27388,N_20047,N_22598);
xnor U27389 (N_27389,N_19121,N_20590);
or U27390 (N_27390,N_19704,N_18989);
nand U27391 (N_27391,N_20177,N_18100);
nor U27392 (N_27392,N_18175,N_18228);
and U27393 (N_27393,N_18729,N_21215);
nand U27394 (N_27394,N_20481,N_20809);
and U27395 (N_27395,N_20878,N_20140);
and U27396 (N_27396,N_18345,N_18869);
or U27397 (N_27397,N_22324,N_22716);
nor U27398 (N_27398,N_21899,N_21361);
xor U27399 (N_27399,N_23045,N_19577);
xnor U27400 (N_27400,N_19007,N_23461);
nor U27401 (N_27401,N_20149,N_21653);
nor U27402 (N_27402,N_22838,N_23288);
nor U27403 (N_27403,N_20837,N_23132);
xnor U27404 (N_27404,N_21321,N_20288);
xnor U27405 (N_27405,N_21476,N_18686);
nor U27406 (N_27406,N_21770,N_21495);
or U27407 (N_27407,N_21051,N_20067);
and U27408 (N_27408,N_22803,N_21253);
nor U27409 (N_27409,N_19937,N_20141);
xor U27410 (N_27410,N_18736,N_23183);
nand U27411 (N_27411,N_18785,N_19077);
nor U27412 (N_27412,N_20718,N_21282);
and U27413 (N_27413,N_19863,N_23104);
and U27414 (N_27414,N_21005,N_22734);
or U27415 (N_27415,N_21121,N_19804);
nor U27416 (N_27416,N_21650,N_19668);
xor U27417 (N_27417,N_20602,N_19761);
or U27418 (N_27418,N_22903,N_20009);
and U27419 (N_27419,N_19856,N_21707);
or U27420 (N_27420,N_23491,N_19058);
nor U27421 (N_27421,N_19065,N_22944);
nor U27422 (N_27422,N_19317,N_20763);
or U27423 (N_27423,N_19066,N_20881);
nor U27424 (N_27424,N_22933,N_19656);
nor U27425 (N_27425,N_20349,N_22714);
or U27426 (N_27426,N_22591,N_19171);
xnor U27427 (N_27427,N_18420,N_23952);
nand U27428 (N_27428,N_23361,N_18606);
and U27429 (N_27429,N_22149,N_19714);
or U27430 (N_27430,N_20605,N_21568);
xnor U27431 (N_27431,N_22075,N_23248);
or U27432 (N_27432,N_22176,N_21221);
and U27433 (N_27433,N_20168,N_20765);
nand U27434 (N_27434,N_20141,N_20726);
and U27435 (N_27435,N_22672,N_21285);
and U27436 (N_27436,N_20897,N_22708);
xnor U27437 (N_27437,N_18255,N_18585);
nor U27438 (N_27438,N_21476,N_22690);
nor U27439 (N_27439,N_22460,N_22598);
nor U27440 (N_27440,N_19376,N_19301);
nor U27441 (N_27441,N_21131,N_18831);
or U27442 (N_27442,N_18629,N_19959);
nand U27443 (N_27443,N_22587,N_20636);
nand U27444 (N_27444,N_22899,N_23818);
and U27445 (N_27445,N_21388,N_18335);
nand U27446 (N_27446,N_22760,N_22816);
and U27447 (N_27447,N_22595,N_23940);
nand U27448 (N_27448,N_23488,N_22834);
or U27449 (N_27449,N_22415,N_18097);
xnor U27450 (N_27450,N_23003,N_19513);
xnor U27451 (N_27451,N_22733,N_19799);
nor U27452 (N_27452,N_19065,N_21284);
xnor U27453 (N_27453,N_22296,N_22991);
nor U27454 (N_27454,N_18944,N_22510);
xnor U27455 (N_27455,N_20552,N_20370);
and U27456 (N_27456,N_20994,N_21930);
and U27457 (N_27457,N_23826,N_18624);
or U27458 (N_27458,N_18125,N_22738);
or U27459 (N_27459,N_19558,N_20907);
nand U27460 (N_27460,N_21759,N_18635);
xor U27461 (N_27461,N_21855,N_18795);
xnor U27462 (N_27462,N_20543,N_18399);
or U27463 (N_27463,N_20966,N_19059);
nand U27464 (N_27464,N_21836,N_20038);
and U27465 (N_27465,N_20564,N_20873);
nor U27466 (N_27466,N_19669,N_22055);
xnor U27467 (N_27467,N_18450,N_19355);
or U27468 (N_27468,N_22401,N_23126);
and U27469 (N_27469,N_19213,N_22695);
xnor U27470 (N_27470,N_20710,N_23755);
or U27471 (N_27471,N_23169,N_20044);
or U27472 (N_27472,N_20576,N_22846);
nand U27473 (N_27473,N_22241,N_20197);
or U27474 (N_27474,N_21788,N_19830);
and U27475 (N_27475,N_18084,N_19654);
nor U27476 (N_27476,N_23202,N_23971);
nor U27477 (N_27477,N_22978,N_23999);
and U27478 (N_27478,N_19046,N_19654);
nor U27479 (N_27479,N_21131,N_21625);
xor U27480 (N_27480,N_18615,N_20777);
nor U27481 (N_27481,N_19711,N_23792);
or U27482 (N_27482,N_18500,N_23160);
or U27483 (N_27483,N_22001,N_22544);
nor U27484 (N_27484,N_23323,N_19455);
or U27485 (N_27485,N_21739,N_22142);
nand U27486 (N_27486,N_20564,N_19383);
or U27487 (N_27487,N_23647,N_20724);
xor U27488 (N_27488,N_20440,N_18246);
and U27489 (N_27489,N_21185,N_21952);
xor U27490 (N_27490,N_18316,N_18403);
xor U27491 (N_27491,N_19450,N_20476);
nand U27492 (N_27492,N_19832,N_20201);
or U27493 (N_27493,N_21568,N_18509);
and U27494 (N_27494,N_18332,N_18942);
nor U27495 (N_27495,N_19037,N_18878);
nor U27496 (N_27496,N_19439,N_18870);
nand U27497 (N_27497,N_22110,N_23788);
nand U27498 (N_27498,N_18487,N_21019);
nand U27499 (N_27499,N_18923,N_20839);
xor U27500 (N_27500,N_21296,N_22994);
nand U27501 (N_27501,N_20301,N_20291);
or U27502 (N_27502,N_20899,N_19905);
and U27503 (N_27503,N_20478,N_23245);
nor U27504 (N_27504,N_18957,N_20484);
nand U27505 (N_27505,N_19102,N_21398);
nor U27506 (N_27506,N_21349,N_18411);
or U27507 (N_27507,N_21909,N_19217);
and U27508 (N_27508,N_22754,N_21605);
nand U27509 (N_27509,N_20996,N_22512);
nand U27510 (N_27510,N_21430,N_23395);
or U27511 (N_27511,N_20442,N_23658);
and U27512 (N_27512,N_21275,N_19084);
or U27513 (N_27513,N_20558,N_22993);
nor U27514 (N_27514,N_23306,N_19430);
nand U27515 (N_27515,N_18237,N_21908);
nor U27516 (N_27516,N_22997,N_20288);
and U27517 (N_27517,N_19538,N_21824);
and U27518 (N_27518,N_18519,N_23441);
and U27519 (N_27519,N_21242,N_20909);
and U27520 (N_27520,N_21291,N_23864);
nand U27521 (N_27521,N_23461,N_22269);
xnor U27522 (N_27522,N_20282,N_23398);
and U27523 (N_27523,N_21289,N_18473);
xor U27524 (N_27524,N_21095,N_19389);
xor U27525 (N_27525,N_23291,N_23431);
nand U27526 (N_27526,N_22520,N_23404);
nor U27527 (N_27527,N_19445,N_23993);
nand U27528 (N_27528,N_22480,N_18256);
xnor U27529 (N_27529,N_23234,N_21749);
xnor U27530 (N_27530,N_20373,N_22481);
or U27531 (N_27531,N_18613,N_22431);
xnor U27532 (N_27532,N_20523,N_22179);
xor U27533 (N_27533,N_19588,N_18552);
nor U27534 (N_27534,N_21823,N_19562);
nor U27535 (N_27535,N_19082,N_23148);
xor U27536 (N_27536,N_19240,N_21885);
or U27537 (N_27537,N_19574,N_20190);
xor U27538 (N_27538,N_18875,N_18799);
xor U27539 (N_27539,N_18195,N_21752);
or U27540 (N_27540,N_22058,N_19176);
or U27541 (N_27541,N_19673,N_20651);
and U27542 (N_27542,N_18357,N_23130);
nor U27543 (N_27543,N_22316,N_19413);
nor U27544 (N_27544,N_22989,N_18992);
nand U27545 (N_27545,N_23986,N_19743);
xor U27546 (N_27546,N_21218,N_18947);
and U27547 (N_27547,N_20170,N_20657);
nor U27548 (N_27548,N_19540,N_18925);
xnor U27549 (N_27549,N_20038,N_22064);
and U27550 (N_27550,N_18630,N_19206);
nor U27551 (N_27551,N_19106,N_21283);
or U27552 (N_27552,N_23770,N_20728);
xnor U27553 (N_27553,N_22736,N_22224);
or U27554 (N_27554,N_18054,N_23535);
nand U27555 (N_27555,N_23934,N_18694);
or U27556 (N_27556,N_18146,N_19190);
nor U27557 (N_27557,N_18818,N_19038);
and U27558 (N_27558,N_20506,N_21645);
or U27559 (N_27559,N_19379,N_22332);
xnor U27560 (N_27560,N_18409,N_19581);
and U27561 (N_27561,N_23188,N_19737);
and U27562 (N_27562,N_21109,N_21483);
or U27563 (N_27563,N_18004,N_22518);
or U27564 (N_27564,N_22518,N_19980);
or U27565 (N_27565,N_21856,N_19312);
and U27566 (N_27566,N_20934,N_19907);
or U27567 (N_27567,N_23747,N_19709);
nor U27568 (N_27568,N_23738,N_18268);
and U27569 (N_27569,N_19658,N_20546);
and U27570 (N_27570,N_22329,N_18131);
nor U27571 (N_27571,N_21369,N_20105);
or U27572 (N_27572,N_20909,N_21227);
nor U27573 (N_27573,N_23698,N_23817);
nor U27574 (N_27574,N_20518,N_21456);
nor U27575 (N_27575,N_21347,N_20156);
nand U27576 (N_27576,N_20348,N_23603);
nor U27577 (N_27577,N_22737,N_18083);
and U27578 (N_27578,N_18959,N_19055);
nand U27579 (N_27579,N_18187,N_23804);
and U27580 (N_27580,N_21376,N_21407);
nor U27581 (N_27581,N_19770,N_20596);
xnor U27582 (N_27582,N_22421,N_18581);
and U27583 (N_27583,N_21660,N_20774);
xor U27584 (N_27584,N_22912,N_18867);
and U27585 (N_27585,N_18742,N_22881);
nor U27586 (N_27586,N_20159,N_22340);
nand U27587 (N_27587,N_21057,N_22471);
or U27588 (N_27588,N_18590,N_18034);
xnor U27589 (N_27589,N_18685,N_21743);
and U27590 (N_27590,N_23499,N_22435);
nand U27591 (N_27591,N_21644,N_22274);
or U27592 (N_27592,N_23100,N_18517);
xnor U27593 (N_27593,N_21056,N_19471);
nand U27594 (N_27594,N_23609,N_18661);
or U27595 (N_27595,N_20457,N_21294);
and U27596 (N_27596,N_23687,N_22195);
nor U27597 (N_27597,N_23655,N_21560);
and U27598 (N_27598,N_21798,N_23149);
or U27599 (N_27599,N_18572,N_18438);
xor U27600 (N_27600,N_18583,N_21157);
nand U27601 (N_27601,N_22245,N_21997);
or U27602 (N_27602,N_21098,N_21917);
and U27603 (N_27603,N_19451,N_23604);
and U27604 (N_27604,N_18021,N_21277);
xor U27605 (N_27605,N_18884,N_22107);
and U27606 (N_27606,N_18176,N_21102);
nor U27607 (N_27607,N_20378,N_19779);
nand U27608 (N_27608,N_19110,N_21414);
xnor U27609 (N_27609,N_23100,N_22877);
xnor U27610 (N_27610,N_21507,N_20875);
or U27611 (N_27611,N_23171,N_21960);
and U27612 (N_27612,N_21886,N_20680);
nand U27613 (N_27613,N_20057,N_23765);
or U27614 (N_27614,N_21302,N_18950);
nand U27615 (N_27615,N_21190,N_21481);
xnor U27616 (N_27616,N_18510,N_19260);
nand U27617 (N_27617,N_19506,N_23784);
and U27618 (N_27618,N_23508,N_19796);
nand U27619 (N_27619,N_19501,N_18773);
nor U27620 (N_27620,N_18945,N_23245);
nor U27621 (N_27621,N_21633,N_21457);
xnor U27622 (N_27622,N_21511,N_18391);
xor U27623 (N_27623,N_18589,N_21431);
and U27624 (N_27624,N_23660,N_21654);
or U27625 (N_27625,N_19609,N_19744);
and U27626 (N_27626,N_23132,N_19642);
nor U27627 (N_27627,N_22229,N_20251);
xnor U27628 (N_27628,N_19222,N_19494);
or U27629 (N_27629,N_23456,N_20657);
nand U27630 (N_27630,N_20689,N_18529);
xnor U27631 (N_27631,N_21999,N_23596);
nand U27632 (N_27632,N_21776,N_23994);
xor U27633 (N_27633,N_20099,N_18041);
nor U27634 (N_27634,N_19554,N_20217);
nand U27635 (N_27635,N_19191,N_19024);
and U27636 (N_27636,N_21126,N_23132);
nor U27637 (N_27637,N_22548,N_19575);
nand U27638 (N_27638,N_22871,N_18556);
and U27639 (N_27639,N_21330,N_22801);
and U27640 (N_27640,N_19098,N_23117);
or U27641 (N_27641,N_18590,N_20821);
xor U27642 (N_27642,N_20992,N_21135);
nor U27643 (N_27643,N_18630,N_23880);
nor U27644 (N_27644,N_18304,N_19510);
nand U27645 (N_27645,N_20782,N_18613);
or U27646 (N_27646,N_18172,N_22147);
nand U27647 (N_27647,N_23813,N_18491);
and U27648 (N_27648,N_23444,N_21209);
nor U27649 (N_27649,N_23544,N_21472);
nor U27650 (N_27650,N_22278,N_18315);
or U27651 (N_27651,N_19546,N_22873);
or U27652 (N_27652,N_23190,N_20822);
nor U27653 (N_27653,N_20567,N_18876);
and U27654 (N_27654,N_20752,N_22049);
or U27655 (N_27655,N_23640,N_19251);
nor U27656 (N_27656,N_23674,N_23216);
nor U27657 (N_27657,N_22406,N_19032);
and U27658 (N_27658,N_18043,N_20202);
or U27659 (N_27659,N_18656,N_21029);
xnor U27660 (N_27660,N_18622,N_23827);
nor U27661 (N_27661,N_22714,N_21240);
and U27662 (N_27662,N_20240,N_23699);
nand U27663 (N_27663,N_20081,N_23743);
nor U27664 (N_27664,N_19999,N_23961);
nand U27665 (N_27665,N_20820,N_19277);
nor U27666 (N_27666,N_19872,N_19500);
nand U27667 (N_27667,N_21221,N_18250);
xor U27668 (N_27668,N_18628,N_22252);
or U27669 (N_27669,N_21180,N_18488);
nand U27670 (N_27670,N_23860,N_22197);
nand U27671 (N_27671,N_19164,N_20205);
and U27672 (N_27672,N_22300,N_20029);
nand U27673 (N_27673,N_19190,N_18415);
nand U27674 (N_27674,N_21046,N_19829);
and U27675 (N_27675,N_23061,N_20718);
or U27676 (N_27676,N_19553,N_20054);
xnor U27677 (N_27677,N_19966,N_19232);
nor U27678 (N_27678,N_19891,N_20214);
nor U27679 (N_27679,N_21678,N_22318);
or U27680 (N_27680,N_18403,N_18855);
xor U27681 (N_27681,N_21001,N_23768);
or U27682 (N_27682,N_21793,N_23613);
and U27683 (N_27683,N_21382,N_19004);
nor U27684 (N_27684,N_21477,N_23474);
and U27685 (N_27685,N_21425,N_20388);
or U27686 (N_27686,N_22012,N_18737);
nor U27687 (N_27687,N_18465,N_19648);
or U27688 (N_27688,N_19437,N_18427);
and U27689 (N_27689,N_21659,N_19704);
or U27690 (N_27690,N_20734,N_22912);
nor U27691 (N_27691,N_19550,N_20704);
nand U27692 (N_27692,N_22520,N_18184);
nor U27693 (N_27693,N_23971,N_18240);
and U27694 (N_27694,N_22178,N_18266);
xor U27695 (N_27695,N_19776,N_19043);
nand U27696 (N_27696,N_20090,N_20780);
and U27697 (N_27697,N_21752,N_18543);
nand U27698 (N_27698,N_19155,N_23485);
nor U27699 (N_27699,N_22234,N_18544);
and U27700 (N_27700,N_20573,N_18448);
xor U27701 (N_27701,N_19576,N_19591);
or U27702 (N_27702,N_21536,N_21968);
xnor U27703 (N_27703,N_23832,N_22453);
nand U27704 (N_27704,N_19681,N_18089);
and U27705 (N_27705,N_21213,N_22614);
xor U27706 (N_27706,N_21557,N_18984);
or U27707 (N_27707,N_22510,N_18207);
xnor U27708 (N_27708,N_20269,N_23482);
xor U27709 (N_27709,N_19137,N_19138);
nand U27710 (N_27710,N_23491,N_23584);
and U27711 (N_27711,N_18578,N_18783);
nand U27712 (N_27712,N_19444,N_18607);
nand U27713 (N_27713,N_22273,N_20077);
nand U27714 (N_27714,N_23621,N_18884);
and U27715 (N_27715,N_22242,N_20947);
or U27716 (N_27716,N_22445,N_23654);
and U27717 (N_27717,N_20205,N_21669);
nor U27718 (N_27718,N_19910,N_23117);
and U27719 (N_27719,N_23108,N_23778);
and U27720 (N_27720,N_19394,N_20632);
or U27721 (N_27721,N_18482,N_20758);
xnor U27722 (N_27722,N_21014,N_20817);
xnor U27723 (N_27723,N_18172,N_18352);
xor U27724 (N_27724,N_21192,N_19041);
xor U27725 (N_27725,N_19673,N_21267);
nand U27726 (N_27726,N_18305,N_20391);
or U27727 (N_27727,N_18967,N_22144);
and U27728 (N_27728,N_20168,N_21026);
or U27729 (N_27729,N_22151,N_18382);
or U27730 (N_27730,N_18803,N_20792);
or U27731 (N_27731,N_21821,N_22869);
or U27732 (N_27732,N_18934,N_22298);
nor U27733 (N_27733,N_23700,N_18400);
and U27734 (N_27734,N_22450,N_22083);
nand U27735 (N_27735,N_21811,N_21406);
or U27736 (N_27736,N_23444,N_21588);
or U27737 (N_27737,N_18843,N_22694);
and U27738 (N_27738,N_21945,N_20480);
nand U27739 (N_27739,N_20347,N_20288);
or U27740 (N_27740,N_19822,N_20501);
and U27741 (N_27741,N_20066,N_20531);
or U27742 (N_27742,N_21108,N_22841);
nand U27743 (N_27743,N_21711,N_21688);
nand U27744 (N_27744,N_23304,N_19988);
nand U27745 (N_27745,N_21527,N_19543);
and U27746 (N_27746,N_20013,N_19676);
and U27747 (N_27747,N_23126,N_22475);
xnor U27748 (N_27748,N_20947,N_23343);
or U27749 (N_27749,N_19347,N_23858);
xnor U27750 (N_27750,N_23855,N_21462);
nor U27751 (N_27751,N_20667,N_21433);
and U27752 (N_27752,N_19499,N_19095);
xnor U27753 (N_27753,N_23934,N_20338);
nand U27754 (N_27754,N_20935,N_21217);
nor U27755 (N_27755,N_20037,N_23189);
and U27756 (N_27756,N_22546,N_21385);
xnor U27757 (N_27757,N_18653,N_21363);
nand U27758 (N_27758,N_22696,N_22757);
xnor U27759 (N_27759,N_23390,N_19623);
nor U27760 (N_27760,N_23372,N_19813);
and U27761 (N_27761,N_23393,N_19195);
or U27762 (N_27762,N_19479,N_20510);
nand U27763 (N_27763,N_22396,N_18808);
or U27764 (N_27764,N_20318,N_22260);
or U27765 (N_27765,N_22935,N_22835);
xor U27766 (N_27766,N_20877,N_22258);
nand U27767 (N_27767,N_19055,N_23282);
xor U27768 (N_27768,N_19650,N_19246);
nand U27769 (N_27769,N_22323,N_20316);
nand U27770 (N_27770,N_20814,N_21556);
nor U27771 (N_27771,N_19580,N_20448);
nor U27772 (N_27772,N_20573,N_22304);
nand U27773 (N_27773,N_19831,N_21351);
xor U27774 (N_27774,N_18429,N_22605);
and U27775 (N_27775,N_23285,N_19096);
nand U27776 (N_27776,N_22357,N_20734);
or U27777 (N_27777,N_19018,N_20855);
xor U27778 (N_27778,N_23972,N_22744);
or U27779 (N_27779,N_18877,N_21192);
and U27780 (N_27780,N_22132,N_20670);
xnor U27781 (N_27781,N_22666,N_21595);
xor U27782 (N_27782,N_19282,N_19070);
nor U27783 (N_27783,N_22221,N_19606);
and U27784 (N_27784,N_21877,N_23777);
nor U27785 (N_27785,N_21155,N_21053);
nor U27786 (N_27786,N_18851,N_19487);
or U27787 (N_27787,N_21938,N_18323);
or U27788 (N_27788,N_19651,N_18285);
and U27789 (N_27789,N_23861,N_23372);
and U27790 (N_27790,N_20829,N_18021);
xor U27791 (N_27791,N_20458,N_18337);
nand U27792 (N_27792,N_23614,N_21316);
xor U27793 (N_27793,N_22847,N_20930);
and U27794 (N_27794,N_21607,N_20535);
or U27795 (N_27795,N_21265,N_18419);
xnor U27796 (N_27796,N_23388,N_18166);
nor U27797 (N_27797,N_19681,N_23054);
and U27798 (N_27798,N_18299,N_19488);
nand U27799 (N_27799,N_21654,N_22136);
xor U27800 (N_27800,N_21048,N_18253);
xor U27801 (N_27801,N_21989,N_22570);
xnor U27802 (N_27802,N_19681,N_18708);
nor U27803 (N_27803,N_22973,N_22558);
nor U27804 (N_27804,N_19122,N_18375);
xnor U27805 (N_27805,N_23155,N_21150);
xnor U27806 (N_27806,N_21506,N_22627);
nor U27807 (N_27807,N_19042,N_22107);
xor U27808 (N_27808,N_19309,N_20707);
nor U27809 (N_27809,N_18998,N_20849);
xnor U27810 (N_27810,N_20350,N_19978);
and U27811 (N_27811,N_21359,N_18003);
or U27812 (N_27812,N_18160,N_18016);
and U27813 (N_27813,N_23675,N_19432);
nand U27814 (N_27814,N_19088,N_18798);
and U27815 (N_27815,N_19216,N_22049);
xor U27816 (N_27816,N_22639,N_21616);
or U27817 (N_27817,N_19779,N_19735);
nand U27818 (N_27818,N_19064,N_18089);
and U27819 (N_27819,N_21091,N_20643);
and U27820 (N_27820,N_22625,N_19813);
xnor U27821 (N_27821,N_18108,N_20136);
nand U27822 (N_27822,N_19901,N_23930);
nand U27823 (N_27823,N_18524,N_22545);
and U27824 (N_27824,N_22149,N_22584);
xnor U27825 (N_27825,N_18431,N_21774);
nand U27826 (N_27826,N_18361,N_20200);
or U27827 (N_27827,N_19086,N_20057);
or U27828 (N_27828,N_18221,N_19936);
and U27829 (N_27829,N_22482,N_22485);
and U27830 (N_27830,N_20478,N_19190);
nor U27831 (N_27831,N_23064,N_19583);
and U27832 (N_27832,N_21258,N_19534);
xor U27833 (N_27833,N_19505,N_19657);
nor U27834 (N_27834,N_20862,N_23235);
and U27835 (N_27835,N_23933,N_23946);
or U27836 (N_27836,N_20910,N_18627);
or U27837 (N_27837,N_19753,N_20976);
and U27838 (N_27838,N_21820,N_23903);
nand U27839 (N_27839,N_18062,N_23990);
and U27840 (N_27840,N_22233,N_19104);
xor U27841 (N_27841,N_18524,N_21615);
nor U27842 (N_27842,N_23252,N_20383);
nor U27843 (N_27843,N_20217,N_22642);
nand U27844 (N_27844,N_20871,N_20778);
nor U27845 (N_27845,N_23013,N_20662);
and U27846 (N_27846,N_23394,N_18978);
xnor U27847 (N_27847,N_23712,N_20397);
nor U27848 (N_27848,N_20022,N_21816);
and U27849 (N_27849,N_20554,N_21291);
and U27850 (N_27850,N_18758,N_20565);
xnor U27851 (N_27851,N_19090,N_21285);
xnor U27852 (N_27852,N_23759,N_20987);
and U27853 (N_27853,N_19836,N_22778);
or U27854 (N_27854,N_20769,N_19394);
or U27855 (N_27855,N_22635,N_19389);
or U27856 (N_27856,N_19169,N_21444);
nand U27857 (N_27857,N_20307,N_23153);
nor U27858 (N_27858,N_18987,N_22024);
xnor U27859 (N_27859,N_18184,N_21765);
xnor U27860 (N_27860,N_18799,N_21613);
and U27861 (N_27861,N_19587,N_20635);
nand U27862 (N_27862,N_18111,N_21206);
nand U27863 (N_27863,N_19274,N_20761);
or U27864 (N_27864,N_22098,N_20567);
nor U27865 (N_27865,N_23362,N_23070);
and U27866 (N_27866,N_21486,N_19872);
and U27867 (N_27867,N_23478,N_21957);
and U27868 (N_27868,N_19013,N_20666);
nor U27869 (N_27869,N_23348,N_23951);
and U27870 (N_27870,N_20622,N_23251);
xnor U27871 (N_27871,N_18714,N_22573);
nor U27872 (N_27872,N_18825,N_19202);
nor U27873 (N_27873,N_19579,N_22982);
or U27874 (N_27874,N_23426,N_22338);
nor U27875 (N_27875,N_20329,N_19263);
xnor U27876 (N_27876,N_18056,N_23360);
nor U27877 (N_27877,N_23160,N_21944);
nor U27878 (N_27878,N_19167,N_20164);
or U27879 (N_27879,N_22345,N_21347);
or U27880 (N_27880,N_20388,N_22465);
and U27881 (N_27881,N_20319,N_19755);
nor U27882 (N_27882,N_23075,N_22457);
or U27883 (N_27883,N_21568,N_20668);
nand U27884 (N_27884,N_21360,N_22202);
nor U27885 (N_27885,N_23407,N_22073);
nor U27886 (N_27886,N_18171,N_18464);
nor U27887 (N_27887,N_22954,N_20908);
or U27888 (N_27888,N_18645,N_19503);
nor U27889 (N_27889,N_23277,N_18324);
nor U27890 (N_27890,N_18415,N_18021);
nand U27891 (N_27891,N_18462,N_23438);
nor U27892 (N_27892,N_18699,N_18567);
and U27893 (N_27893,N_23590,N_23427);
nor U27894 (N_27894,N_23157,N_22755);
nand U27895 (N_27895,N_23897,N_20901);
xor U27896 (N_27896,N_22603,N_23006);
xnor U27897 (N_27897,N_21256,N_19495);
nand U27898 (N_27898,N_21048,N_21230);
nand U27899 (N_27899,N_19776,N_22463);
xor U27900 (N_27900,N_22780,N_23616);
nand U27901 (N_27901,N_20261,N_20899);
or U27902 (N_27902,N_22307,N_23114);
and U27903 (N_27903,N_19599,N_18257);
or U27904 (N_27904,N_22862,N_18180);
xnor U27905 (N_27905,N_22596,N_19783);
nand U27906 (N_27906,N_20794,N_18256);
or U27907 (N_27907,N_19238,N_18665);
or U27908 (N_27908,N_21938,N_18092);
nand U27909 (N_27909,N_20852,N_22900);
or U27910 (N_27910,N_18282,N_22610);
nor U27911 (N_27911,N_23217,N_23493);
and U27912 (N_27912,N_22450,N_21192);
xnor U27913 (N_27913,N_18949,N_18490);
nand U27914 (N_27914,N_21928,N_22847);
nand U27915 (N_27915,N_19276,N_19441);
or U27916 (N_27916,N_20618,N_23966);
and U27917 (N_27917,N_18569,N_22262);
and U27918 (N_27918,N_19644,N_22720);
xor U27919 (N_27919,N_21405,N_21795);
nor U27920 (N_27920,N_18472,N_21457);
xnor U27921 (N_27921,N_22738,N_21216);
xor U27922 (N_27922,N_23074,N_18951);
nor U27923 (N_27923,N_19499,N_22989);
and U27924 (N_27924,N_18483,N_18381);
xnor U27925 (N_27925,N_21031,N_21400);
nor U27926 (N_27926,N_23028,N_21227);
xor U27927 (N_27927,N_23568,N_23114);
and U27928 (N_27928,N_23282,N_18652);
or U27929 (N_27929,N_23568,N_21927);
xnor U27930 (N_27930,N_22694,N_18282);
and U27931 (N_27931,N_18522,N_19589);
and U27932 (N_27932,N_21884,N_18533);
nand U27933 (N_27933,N_23606,N_23632);
and U27934 (N_27934,N_22416,N_22317);
or U27935 (N_27935,N_19642,N_20676);
xnor U27936 (N_27936,N_21586,N_23353);
nand U27937 (N_27937,N_23337,N_23004);
nand U27938 (N_27938,N_23398,N_21101);
nor U27939 (N_27939,N_19837,N_18987);
xor U27940 (N_27940,N_20190,N_21514);
nand U27941 (N_27941,N_19557,N_19026);
or U27942 (N_27942,N_18897,N_20499);
nand U27943 (N_27943,N_21221,N_19349);
xnor U27944 (N_27944,N_20614,N_23560);
or U27945 (N_27945,N_22358,N_20531);
xnor U27946 (N_27946,N_19297,N_19236);
xor U27947 (N_27947,N_20908,N_19083);
nor U27948 (N_27948,N_20950,N_20133);
or U27949 (N_27949,N_19106,N_19584);
or U27950 (N_27950,N_19851,N_20618);
nor U27951 (N_27951,N_21430,N_18019);
and U27952 (N_27952,N_21346,N_18251);
xor U27953 (N_27953,N_22999,N_21163);
xor U27954 (N_27954,N_23927,N_21260);
xnor U27955 (N_27955,N_21052,N_19773);
xor U27956 (N_27956,N_23961,N_21373);
or U27957 (N_27957,N_23956,N_20173);
nor U27958 (N_27958,N_21285,N_19583);
xor U27959 (N_27959,N_22430,N_21875);
nor U27960 (N_27960,N_19671,N_22910);
or U27961 (N_27961,N_19231,N_19698);
or U27962 (N_27962,N_21716,N_20313);
and U27963 (N_27963,N_23902,N_20484);
nand U27964 (N_27964,N_23366,N_22835);
xnor U27965 (N_27965,N_18383,N_23036);
or U27966 (N_27966,N_22290,N_21131);
nand U27967 (N_27967,N_20132,N_20062);
nor U27968 (N_27968,N_23827,N_19324);
and U27969 (N_27969,N_22042,N_19469);
nor U27970 (N_27970,N_18828,N_23434);
or U27971 (N_27971,N_19156,N_23494);
or U27972 (N_27972,N_18978,N_20324);
or U27973 (N_27973,N_21207,N_22132);
and U27974 (N_27974,N_18137,N_18641);
and U27975 (N_27975,N_18108,N_19580);
xor U27976 (N_27976,N_18903,N_22162);
xnor U27977 (N_27977,N_23466,N_21011);
nor U27978 (N_27978,N_18364,N_21155);
nor U27979 (N_27979,N_20571,N_22233);
xnor U27980 (N_27980,N_18371,N_20309);
or U27981 (N_27981,N_23556,N_20358);
nor U27982 (N_27982,N_21255,N_18906);
nand U27983 (N_27983,N_23394,N_21981);
or U27984 (N_27984,N_22530,N_18757);
nor U27985 (N_27985,N_20427,N_19788);
nand U27986 (N_27986,N_23391,N_21386);
or U27987 (N_27987,N_19585,N_19458);
nor U27988 (N_27988,N_18625,N_19375);
nor U27989 (N_27989,N_23534,N_22565);
or U27990 (N_27990,N_19976,N_19406);
nor U27991 (N_27991,N_23728,N_22813);
and U27992 (N_27992,N_18255,N_20458);
and U27993 (N_27993,N_23605,N_18119);
nor U27994 (N_27994,N_21228,N_18479);
nand U27995 (N_27995,N_21806,N_22897);
xnor U27996 (N_27996,N_21032,N_23075);
or U27997 (N_27997,N_19379,N_21617);
and U27998 (N_27998,N_18510,N_22244);
xnor U27999 (N_27999,N_19312,N_20930);
nor U28000 (N_28000,N_22413,N_18373);
nand U28001 (N_28001,N_22646,N_19000);
xor U28002 (N_28002,N_20777,N_19264);
nand U28003 (N_28003,N_20233,N_22135);
nor U28004 (N_28004,N_21560,N_22999);
xor U28005 (N_28005,N_20422,N_19564);
xor U28006 (N_28006,N_19913,N_23141);
or U28007 (N_28007,N_21914,N_20339);
nor U28008 (N_28008,N_22487,N_21701);
or U28009 (N_28009,N_19165,N_19729);
or U28010 (N_28010,N_20246,N_19003);
xnor U28011 (N_28011,N_21418,N_23070);
nor U28012 (N_28012,N_20420,N_18686);
or U28013 (N_28013,N_19154,N_19219);
nor U28014 (N_28014,N_22089,N_22144);
nor U28015 (N_28015,N_20351,N_20675);
xor U28016 (N_28016,N_22128,N_19326);
and U28017 (N_28017,N_21528,N_22671);
nand U28018 (N_28018,N_23323,N_23217);
xnor U28019 (N_28019,N_22986,N_20562);
xnor U28020 (N_28020,N_20903,N_18655);
nand U28021 (N_28021,N_18847,N_23175);
nor U28022 (N_28022,N_20651,N_18239);
nor U28023 (N_28023,N_20140,N_22410);
or U28024 (N_28024,N_19114,N_23183);
and U28025 (N_28025,N_22658,N_18650);
nand U28026 (N_28026,N_18113,N_22098);
nor U28027 (N_28027,N_21718,N_20933);
or U28028 (N_28028,N_23355,N_22075);
and U28029 (N_28029,N_22032,N_18133);
and U28030 (N_28030,N_20126,N_23441);
nand U28031 (N_28031,N_18416,N_21444);
nand U28032 (N_28032,N_20235,N_20200);
or U28033 (N_28033,N_20436,N_21321);
xnor U28034 (N_28034,N_20596,N_22313);
and U28035 (N_28035,N_23961,N_23050);
or U28036 (N_28036,N_21326,N_21637);
nor U28037 (N_28037,N_23859,N_22023);
or U28038 (N_28038,N_22139,N_22670);
xnor U28039 (N_28039,N_20434,N_22376);
nor U28040 (N_28040,N_18759,N_20101);
nor U28041 (N_28041,N_18883,N_18411);
and U28042 (N_28042,N_20425,N_18191);
nand U28043 (N_28043,N_18023,N_23256);
and U28044 (N_28044,N_20006,N_19102);
nor U28045 (N_28045,N_19059,N_23678);
and U28046 (N_28046,N_19170,N_20842);
and U28047 (N_28047,N_18747,N_22793);
nor U28048 (N_28048,N_19826,N_19650);
nand U28049 (N_28049,N_23106,N_20784);
nand U28050 (N_28050,N_18427,N_18171);
nand U28051 (N_28051,N_21184,N_19628);
and U28052 (N_28052,N_19095,N_20165);
and U28053 (N_28053,N_21814,N_21245);
nand U28054 (N_28054,N_23343,N_21941);
nor U28055 (N_28055,N_23458,N_19308);
xnor U28056 (N_28056,N_18096,N_23597);
and U28057 (N_28057,N_19795,N_19369);
xnor U28058 (N_28058,N_22373,N_23963);
nor U28059 (N_28059,N_20928,N_18765);
and U28060 (N_28060,N_21364,N_23369);
nor U28061 (N_28061,N_22374,N_19239);
or U28062 (N_28062,N_20224,N_18790);
or U28063 (N_28063,N_23679,N_23801);
xnor U28064 (N_28064,N_22031,N_21529);
and U28065 (N_28065,N_21251,N_19370);
nor U28066 (N_28066,N_20175,N_19016);
nand U28067 (N_28067,N_21197,N_20863);
or U28068 (N_28068,N_22633,N_23065);
nor U28069 (N_28069,N_22987,N_22160);
and U28070 (N_28070,N_21478,N_18365);
and U28071 (N_28071,N_21755,N_22721);
xor U28072 (N_28072,N_20762,N_18853);
or U28073 (N_28073,N_21469,N_19625);
or U28074 (N_28074,N_18967,N_19421);
xor U28075 (N_28075,N_18990,N_22992);
nor U28076 (N_28076,N_19443,N_21056);
and U28077 (N_28077,N_20015,N_19009);
and U28078 (N_28078,N_20047,N_20069);
nor U28079 (N_28079,N_20230,N_22555);
nor U28080 (N_28080,N_23669,N_19346);
nand U28081 (N_28081,N_23472,N_23919);
xnor U28082 (N_28082,N_23348,N_23934);
and U28083 (N_28083,N_20324,N_18062);
nor U28084 (N_28084,N_21141,N_20011);
nor U28085 (N_28085,N_22736,N_23127);
and U28086 (N_28086,N_21015,N_23063);
or U28087 (N_28087,N_19104,N_18018);
nand U28088 (N_28088,N_18407,N_19214);
nand U28089 (N_28089,N_20069,N_21317);
nand U28090 (N_28090,N_18633,N_23670);
and U28091 (N_28091,N_22871,N_22832);
or U28092 (N_28092,N_23871,N_20843);
and U28093 (N_28093,N_18194,N_22598);
and U28094 (N_28094,N_19533,N_21811);
xnor U28095 (N_28095,N_19802,N_20353);
and U28096 (N_28096,N_22000,N_20007);
or U28097 (N_28097,N_23536,N_18326);
nor U28098 (N_28098,N_18379,N_19776);
or U28099 (N_28099,N_23245,N_21374);
and U28100 (N_28100,N_19410,N_21979);
and U28101 (N_28101,N_23092,N_23504);
and U28102 (N_28102,N_20624,N_18004);
and U28103 (N_28103,N_20740,N_20716);
and U28104 (N_28104,N_23647,N_22072);
nor U28105 (N_28105,N_21060,N_22203);
nand U28106 (N_28106,N_21575,N_23747);
nor U28107 (N_28107,N_22197,N_21479);
and U28108 (N_28108,N_23412,N_21717);
nand U28109 (N_28109,N_22763,N_21674);
or U28110 (N_28110,N_20454,N_18103);
xnor U28111 (N_28111,N_18358,N_19552);
or U28112 (N_28112,N_20977,N_19978);
xnor U28113 (N_28113,N_23393,N_18984);
or U28114 (N_28114,N_21782,N_21469);
nor U28115 (N_28115,N_22469,N_23348);
nand U28116 (N_28116,N_18778,N_22090);
or U28117 (N_28117,N_21961,N_22671);
or U28118 (N_28118,N_19521,N_22727);
xnor U28119 (N_28119,N_21947,N_21943);
nand U28120 (N_28120,N_23870,N_21906);
or U28121 (N_28121,N_22562,N_22008);
or U28122 (N_28122,N_21313,N_23269);
or U28123 (N_28123,N_18787,N_21050);
and U28124 (N_28124,N_23452,N_22830);
xnor U28125 (N_28125,N_20197,N_19514);
nor U28126 (N_28126,N_19155,N_21926);
nor U28127 (N_28127,N_19750,N_23867);
and U28128 (N_28128,N_22531,N_21778);
xor U28129 (N_28129,N_18020,N_23330);
or U28130 (N_28130,N_21271,N_23306);
and U28131 (N_28131,N_18496,N_20234);
and U28132 (N_28132,N_21544,N_20600);
nor U28133 (N_28133,N_19358,N_20948);
or U28134 (N_28134,N_22390,N_21283);
and U28135 (N_28135,N_19708,N_23764);
nand U28136 (N_28136,N_23232,N_18304);
nor U28137 (N_28137,N_22040,N_22593);
xnor U28138 (N_28138,N_18096,N_22195);
xor U28139 (N_28139,N_23102,N_18178);
xnor U28140 (N_28140,N_19695,N_20780);
or U28141 (N_28141,N_22786,N_20773);
and U28142 (N_28142,N_18905,N_23875);
nor U28143 (N_28143,N_21033,N_21408);
and U28144 (N_28144,N_20962,N_20327);
or U28145 (N_28145,N_21075,N_18815);
xnor U28146 (N_28146,N_21655,N_19199);
or U28147 (N_28147,N_23197,N_22397);
nand U28148 (N_28148,N_19843,N_21808);
or U28149 (N_28149,N_20451,N_18367);
nor U28150 (N_28150,N_20494,N_23166);
nand U28151 (N_28151,N_21327,N_22305);
xnor U28152 (N_28152,N_21747,N_18150);
xor U28153 (N_28153,N_18963,N_19067);
or U28154 (N_28154,N_18303,N_21948);
nand U28155 (N_28155,N_20194,N_22768);
nand U28156 (N_28156,N_23704,N_23120);
nor U28157 (N_28157,N_21449,N_22064);
and U28158 (N_28158,N_21914,N_23278);
or U28159 (N_28159,N_23157,N_20136);
xor U28160 (N_28160,N_20008,N_18196);
nor U28161 (N_28161,N_22378,N_23629);
or U28162 (N_28162,N_20210,N_19741);
nand U28163 (N_28163,N_23361,N_22629);
xnor U28164 (N_28164,N_18676,N_22006);
nor U28165 (N_28165,N_21778,N_19944);
xnor U28166 (N_28166,N_23864,N_19202);
nand U28167 (N_28167,N_23056,N_22904);
nor U28168 (N_28168,N_19276,N_20841);
or U28169 (N_28169,N_18563,N_20801);
and U28170 (N_28170,N_19773,N_21746);
nand U28171 (N_28171,N_20533,N_21424);
or U28172 (N_28172,N_19088,N_19681);
or U28173 (N_28173,N_20720,N_18281);
and U28174 (N_28174,N_18503,N_18378);
nor U28175 (N_28175,N_22805,N_23799);
and U28176 (N_28176,N_18948,N_21510);
nor U28177 (N_28177,N_21906,N_22696);
or U28178 (N_28178,N_22435,N_21558);
and U28179 (N_28179,N_20906,N_19999);
or U28180 (N_28180,N_21106,N_21344);
nand U28181 (N_28181,N_19710,N_22832);
xnor U28182 (N_28182,N_22893,N_21520);
nor U28183 (N_28183,N_20509,N_23679);
nor U28184 (N_28184,N_23782,N_20776);
or U28185 (N_28185,N_22710,N_20624);
or U28186 (N_28186,N_20575,N_18536);
xnor U28187 (N_28187,N_18731,N_20081);
nor U28188 (N_28188,N_21522,N_19066);
or U28189 (N_28189,N_19938,N_20252);
nand U28190 (N_28190,N_22742,N_20826);
nand U28191 (N_28191,N_20740,N_21897);
and U28192 (N_28192,N_19399,N_21262);
nor U28193 (N_28193,N_23922,N_19627);
or U28194 (N_28194,N_18761,N_20100);
and U28195 (N_28195,N_20796,N_18031);
and U28196 (N_28196,N_23988,N_19063);
nand U28197 (N_28197,N_18008,N_21150);
and U28198 (N_28198,N_19858,N_19254);
nor U28199 (N_28199,N_23657,N_21841);
nand U28200 (N_28200,N_18698,N_21086);
and U28201 (N_28201,N_18539,N_18611);
nor U28202 (N_28202,N_18476,N_20304);
or U28203 (N_28203,N_21359,N_18698);
and U28204 (N_28204,N_19697,N_23605);
nor U28205 (N_28205,N_20704,N_23072);
nand U28206 (N_28206,N_23385,N_23625);
and U28207 (N_28207,N_19874,N_22113);
xnor U28208 (N_28208,N_19145,N_20232);
nand U28209 (N_28209,N_23750,N_19795);
and U28210 (N_28210,N_23048,N_18855);
and U28211 (N_28211,N_20048,N_18756);
xnor U28212 (N_28212,N_18424,N_21375);
or U28213 (N_28213,N_23077,N_19802);
xnor U28214 (N_28214,N_22058,N_21955);
nor U28215 (N_28215,N_22063,N_18660);
or U28216 (N_28216,N_22880,N_18458);
or U28217 (N_28217,N_20757,N_18673);
or U28218 (N_28218,N_22222,N_20606);
nor U28219 (N_28219,N_21163,N_19171);
nand U28220 (N_28220,N_22964,N_21739);
nor U28221 (N_28221,N_23258,N_23052);
nor U28222 (N_28222,N_20683,N_21555);
xor U28223 (N_28223,N_19225,N_22996);
or U28224 (N_28224,N_23722,N_21934);
xor U28225 (N_28225,N_21932,N_22062);
and U28226 (N_28226,N_23852,N_21289);
and U28227 (N_28227,N_23167,N_23942);
xor U28228 (N_28228,N_19876,N_23409);
xor U28229 (N_28229,N_21670,N_19176);
nand U28230 (N_28230,N_21922,N_23032);
xnor U28231 (N_28231,N_21909,N_19269);
nor U28232 (N_28232,N_19728,N_23276);
and U28233 (N_28233,N_23846,N_23719);
and U28234 (N_28234,N_19887,N_19093);
and U28235 (N_28235,N_21549,N_23848);
nand U28236 (N_28236,N_20505,N_21400);
and U28237 (N_28237,N_21378,N_21795);
nand U28238 (N_28238,N_22987,N_20663);
nor U28239 (N_28239,N_19681,N_23266);
nand U28240 (N_28240,N_22100,N_23012);
and U28241 (N_28241,N_18846,N_18031);
and U28242 (N_28242,N_19560,N_23257);
nor U28243 (N_28243,N_19616,N_22055);
or U28244 (N_28244,N_20545,N_22414);
or U28245 (N_28245,N_18550,N_22471);
xor U28246 (N_28246,N_18240,N_23528);
nor U28247 (N_28247,N_18477,N_23933);
xnor U28248 (N_28248,N_20895,N_20043);
nor U28249 (N_28249,N_21933,N_18985);
and U28250 (N_28250,N_20048,N_19300);
or U28251 (N_28251,N_23175,N_20701);
xor U28252 (N_28252,N_18141,N_22396);
and U28253 (N_28253,N_22022,N_23029);
xor U28254 (N_28254,N_22828,N_23010);
nor U28255 (N_28255,N_20397,N_20629);
nand U28256 (N_28256,N_23786,N_20328);
nor U28257 (N_28257,N_23416,N_20506);
xnor U28258 (N_28258,N_18638,N_18658);
nand U28259 (N_28259,N_21379,N_22218);
nor U28260 (N_28260,N_23308,N_21256);
and U28261 (N_28261,N_20507,N_23336);
or U28262 (N_28262,N_23998,N_18661);
nand U28263 (N_28263,N_21212,N_21657);
and U28264 (N_28264,N_19596,N_18631);
nand U28265 (N_28265,N_22148,N_23722);
nor U28266 (N_28266,N_20670,N_22626);
or U28267 (N_28267,N_20848,N_23765);
and U28268 (N_28268,N_22048,N_21266);
nor U28269 (N_28269,N_19126,N_21868);
xnor U28270 (N_28270,N_18821,N_22827);
nor U28271 (N_28271,N_21832,N_23539);
or U28272 (N_28272,N_22413,N_22056);
nand U28273 (N_28273,N_21592,N_21759);
nor U28274 (N_28274,N_18102,N_23861);
or U28275 (N_28275,N_19325,N_23256);
nand U28276 (N_28276,N_22214,N_21404);
nand U28277 (N_28277,N_19443,N_23128);
nand U28278 (N_28278,N_18999,N_22882);
xor U28279 (N_28279,N_20308,N_23503);
nand U28280 (N_28280,N_23848,N_23748);
and U28281 (N_28281,N_21125,N_19091);
nor U28282 (N_28282,N_20828,N_21570);
or U28283 (N_28283,N_23002,N_22284);
and U28284 (N_28284,N_22016,N_21408);
and U28285 (N_28285,N_21658,N_18224);
nand U28286 (N_28286,N_22225,N_19926);
or U28287 (N_28287,N_23986,N_18962);
xnor U28288 (N_28288,N_22427,N_20963);
xnor U28289 (N_28289,N_22934,N_22166);
nand U28290 (N_28290,N_22774,N_19327);
and U28291 (N_28291,N_22154,N_21352);
xor U28292 (N_28292,N_21245,N_21318);
and U28293 (N_28293,N_21564,N_18202);
xor U28294 (N_28294,N_20328,N_19164);
and U28295 (N_28295,N_21733,N_19085);
nand U28296 (N_28296,N_19119,N_21255);
nand U28297 (N_28297,N_18819,N_20391);
and U28298 (N_28298,N_19711,N_22467);
and U28299 (N_28299,N_23732,N_18008);
xnor U28300 (N_28300,N_20153,N_19378);
xor U28301 (N_28301,N_19755,N_18530);
or U28302 (N_28302,N_23595,N_18728);
and U28303 (N_28303,N_20062,N_18568);
and U28304 (N_28304,N_21898,N_19885);
xor U28305 (N_28305,N_21868,N_23592);
or U28306 (N_28306,N_18395,N_23675);
xor U28307 (N_28307,N_22499,N_21604);
xor U28308 (N_28308,N_20817,N_19154);
nor U28309 (N_28309,N_22395,N_21453);
xor U28310 (N_28310,N_19076,N_18771);
xnor U28311 (N_28311,N_18996,N_22615);
nor U28312 (N_28312,N_21576,N_21969);
or U28313 (N_28313,N_22042,N_22697);
xor U28314 (N_28314,N_19358,N_19614);
or U28315 (N_28315,N_18630,N_23304);
xor U28316 (N_28316,N_23694,N_21744);
nand U28317 (N_28317,N_19737,N_19188);
and U28318 (N_28318,N_22592,N_19198);
nand U28319 (N_28319,N_23847,N_21098);
nor U28320 (N_28320,N_20421,N_19894);
nand U28321 (N_28321,N_23900,N_20747);
xnor U28322 (N_28322,N_23623,N_21517);
or U28323 (N_28323,N_22213,N_23041);
nor U28324 (N_28324,N_20988,N_20375);
xor U28325 (N_28325,N_18048,N_22939);
or U28326 (N_28326,N_22657,N_23175);
or U28327 (N_28327,N_21094,N_22774);
nor U28328 (N_28328,N_21699,N_23070);
xnor U28329 (N_28329,N_18395,N_21302);
nor U28330 (N_28330,N_23891,N_19671);
xor U28331 (N_28331,N_22182,N_21790);
or U28332 (N_28332,N_22373,N_19916);
nor U28333 (N_28333,N_22486,N_21945);
and U28334 (N_28334,N_22115,N_20963);
or U28335 (N_28335,N_21027,N_21949);
and U28336 (N_28336,N_21976,N_20250);
nor U28337 (N_28337,N_20602,N_23792);
or U28338 (N_28338,N_19231,N_20068);
or U28339 (N_28339,N_19801,N_22180);
xnor U28340 (N_28340,N_23283,N_18418);
nor U28341 (N_28341,N_23008,N_19684);
nor U28342 (N_28342,N_21636,N_22895);
nand U28343 (N_28343,N_22070,N_18698);
xor U28344 (N_28344,N_21512,N_21135);
xnor U28345 (N_28345,N_23108,N_19221);
and U28346 (N_28346,N_23357,N_22842);
or U28347 (N_28347,N_20519,N_22981);
nand U28348 (N_28348,N_22927,N_20539);
nor U28349 (N_28349,N_18623,N_18977);
and U28350 (N_28350,N_23077,N_21075);
and U28351 (N_28351,N_21019,N_21178);
or U28352 (N_28352,N_21559,N_23056);
nand U28353 (N_28353,N_19297,N_19826);
and U28354 (N_28354,N_21681,N_22979);
and U28355 (N_28355,N_21608,N_22599);
or U28356 (N_28356,N_19793,N_23005);
xnor U28357 (N_28357,N_23841,N_23886);
or U28358 (N_28358,N_18990,N_23818);
xor U28359 (N_28359,N_21174,N_18589);
nor U28360 (N_28360,N_20154,N_22651);
nand U28361 (N_28361,N_19121,N_21665);
and U28362 (N_28362,N_22967,N_21616);
and U28363 (N_28363,N_21706,N_23142);
or U28364 (N_28364,N_22067,N_20676);
nand U28365 (N_28365,N_22790,N_21502);
nand U28366 (N_28366,N_23824,N_22971);
nand U28367 (N_28367,N_20265,N_22288);
nand U28368 (N_28368,N_22486,N_22812);
or U28369 (N_28369,N_20666,N_22907);
nor U28370 (N_28370,N_19488,N_20846);
nor U28371 (N_28371,N_23172,N_21546);
and U28372 (N_28372,N_19604,N_21205);
nor U28373 (N_28373,N_19742,N_23958);
xnor U28374 (N_28374,N_23787,N_23811);
nor U28375 (N_28375,N_21887,N_23346);
and U28376 (N_28376,N_23979,N_22449);
xor U28377 (N_28377,N_21410,N_18488);
nand U28378 (N_28378,N_22557,N_21260);
xor U28379 (N_28379,N_21834,N_18198);
nand U28380 (N_28380,N_20769,N_19646);
nor U28381 (N_28381,N_21021,N_18974);
and U28382 (N_28382,N_19419,N_20261);
and U28383 (N_28383,N_23837,N_23316);
and U28384 (N_28384,N_23685,N_18926);
nand U28385 (N_28385,N_19361,N_21198);
nand U28386 (N_28386,N_18933,N_19006);
and U28387 (N_28387,N_22248,N_20056);
xor U28388 (N_28388,N_18360,N_21419);
nand U28389 (N_28389,N_21215,N_21326);
nor U28390 (N_28390,N_23196,N_21047);
and U28391 (N_28391,N_23149,N_21455);
nor U28392 (N_28392,N_22986,N_21203);
nand U28393 (N_28393,N_22109,N_18948);
nand U28394 (N_28394,N_23813,N_23474);
nor U28395 (N_28395,N_21788,N_20680);
nand U28396 (N_28396,N_22319,N_19315);
nor U28397 (N_28397,N_18472,N_22543);
or U28398 (N_28398,N_23844,N_21043);
and U28399 (N_28399,N_21829,N_20831);
or U28400 (N_28400,N_23768,N_18535);
and U28401 (N_28401,N_22233,N_23160);
and U28402 (N_28402,N_22604,N_20931);
and U28403 (N_28403,N_22053,N_18520);
or U28404 (N_28404,N_23495,N_23996);
or U28405 (N_28405,N_22574,N_22756);
or U28406 (N_28406,N_22058,N_21363);
nand U28407 (N_28407,N_21217,N_23471);
nor U28408 (N_28408,N_19974,N_19169);
nor U28409 (N_28409,N_22591,N_22447);
nand U28410 (N_28410,N_18317,N_21544);
nand U28411 (N_28411,N_18071,N_19709);
nor U28412 (N_28412,N_19723,N_20444);
nand U28413 (N_28413,N_21602,N_20983);
nor U28414 (N_28414,N_18352,N_19054);
nand U28415 (N_28415,N_20026,N_23266);
and U28416 (N_28416,N_18784,N_21556);
or U28417 (N_28417,N_23275,N_19136);
and U28418 (N_28418,N_18848,N_21397);
and U28419 (N_28419,N_22325,N_19683);
or U28420 (N_28420,N_18448,N_22850);
xnor U28421 (N_28421,N_22566,N_23142);
or U28422 (N_28422,N_22786,N_19661);
xnor U28423 (N_28423,N_18869,N_22298);
nor U28424 (N_28424,N_23144,N_22302);
or U28425 (N_28425,N_22444,N_20659);
and U28426 (N_28426,N_23601,N_20764);
and U28427 (N_28427,N_20676,N_18441);
or U28428 (N_28428,N_22819,N_19832);
and U28429 (N_28429,N_23853,N_18357);
nor U28430 (N_28430,N_23226,N_19202);
nand U28431 (N_28431,N_18304,N_23010);
nand U28432 (N_28432,N_23178,N_21189);
or U28433 (N_28433,N_20631,N_19484);
or U28434 (N_28434,N_19484,N_18138);
or U28435 (N_28435,N_18225,N_19805);
and U28436 (N_28436,N_19645,N_22266);
or U28437 (N_28437,N_21534,N_20771);
and U28438 (N_28438,N_21362,N_22345);
or U28439 (N_28439,N_22948,N_18895);
nor U28440 (N_28440,N_18981,N_20958);
nor U28441 (N_28441,N_23239,N_23621);
nand U28442 (N_28442,N_18580,N_20748);
or U28443 (N_28443,N_19108,N_20993);
and U28444 (N_28444,N_19732,N_18369);
xor U28445 (N_28445,N_19795,N_23813);
nand U28446 (N_28446,N_20784,N_20189);
xnor U28447 (N_28447,N_18928,N_22201);
xnor U28448 (N_28448,N_22401,N_20354);
xnor U28449 (N_28449,N_22778,N_22791);
and U28450 (N_28450,N_21919,N_20785);
nand U28451 (N_28451,N_19092,N_22069);
or U28452 (N_28452,N_20384,N_22249);
xnor U28453 (N_28453,N_19614,N_18800);
and U28454 (N_28454,N_19667,N_21884);
xnor U28455 (N_28455,N_20011,N_21575);
and U28456 (N_28456,N_22256,N_19041);
and U28457 (N_28457,N_18298,N_23316);
nand U28458 (N_28458,N_22291,N_20884);
nand U28459 (N_28459,N_18705,N_19723);
nand U28460 (N_28460,N_18943,N_23979);
xnor U28461 (N_28461,N_22352,N_23297);
nand U28462 (N_28462,N_19949,N_18797);
and U28463 (N_28463,N_23614,N_19046);
nor U28464 (N_28464,N_18875,N_22823);
or U28465 (N_28465,N_22925,N_18371);
nor U28466 (N_28466,N_20398,N_22397);
and U28467 (N_28467,N_18590,N_20121);
and U28468 (N_28468,N_20880,N_19718);
or U28469 (N_28469,N_19559,N_23734);
or U28470 (N_28470,N_22162,N_18928);
nor U28471 (N_28471,N_22338,N_20038);
xor U28472 (N_28472,N_23215,N_23556);
or U28473 (N_28473,N_20603,N_19911);
nor U28474 (N_28474,N_22929,N_23877);
or U28475 (N_28475,N_23200,N_21949);
or U28476 (N_28476,N_19576,N_19798);
and U28477 (N_28477,N_21739,N_22484);
and U28478 (N_28478,N_23388,N_22120);
or U28479 (N_28479,N_19880,N_19574);
and U28480 (N_28480,N_21478,N_19487);
and U28481 (N_28481,N_20478,N_21730);
xor U28482 (N_28482,N_23926,N_18677);
and U28483 (N_28483,N_22497,N_19299);
xnor U28484 (N_28484,N_23873,N_23408);
nor U28485 (N_28485,N_21872,N_21764);
nor U28486 (N_28486,N_20721,N_19263);
or U28487 (N_28487,N_20116,N_19978);
nor U28488 (N_28488,N_23313,N_21225);
and U28489 (N_28489,N_22485,N_22808);
or U28490 (N_28490,N_23568,N_21583);
or U28491 (N_28491,N_20688,N_22511);
or U28492 (N_28492,N_20045,N_23334);
nand U28493 (N_28493,N_19724,N_18323);
xnor U28494 (N_28494,N_23913,N_19781);
and U28495 (N_28495,N_19752,N_21383);
xnor U28496 (N_28496,N_19341,N_19472);
xnor U28497 (N_28497,N_20468,N_22518);
xnor U28498 (N_28498,N_20019,N_20749);
and U28499 (N_28499,N_23615,N_21988);
and U28500 (N_28500,N_19628,N_23046);
or U28501 (N_28501,N_20438,N_20469);
xnor U28502 (N_28502,N_20674,N_18468);
or U28503 (N_28503,N_20077,N_21723);
xor U28504 (N_28504,N_21384,N_18678);
xor U28505 (N_28505,N_21190,N_20413);
and U28506 (N_28506,N_23769,N_20830);
nand U28507 (N_28507,N_19704,N_18965);
nor U28508 (N_28508,N_18904,N_18661);
xor U28509 (N_28509,N_18933,N_18182);
xor U28510 (N_28510,N_19198,N_23655);
xnor U28511 (N_28511,N_18617,N_19142);
nor U28512 (N_28512,N_22569,N_23774);
and U28513 (N_28513,N_23291,N_21880);
nand U28514 (N_28514,N_20471,N_22603);
xnor U28515 (N_28515,N_23851,N_21565);
and U28516 (N_28516,N_22191,N_18438);
nor U28517 (N_28517,N_22840,N_19726);
xor U28518 (N_28518,N_18593,N_21284);
nand U28519 (N_28519,N_20668,N_19853);
nand U28520 (N_28520,N_21020,N_20530);
or U28521 (N_28521,N_18507,N_20995);
nor U28522 (N_28522,N_22563,N_18859);
xnor U28523 (N_28523,N_18145,N_19102);
xor U28524 (N_28524,N_22055,N_20589);
nor U28525 (N_28525,N_18091,N_21647);
nor U28526 (N_28526,N_20335,N_19244);
xor U28527 (N_28527,N_22433,N_19593);
nand U28528 (N_28528,N_23648,N_23199);
or U28529 (N_28529,N_22583,N_19728);
or U28530 (N_28530,N_20405,N_22576);
and U28531 (N_28531,N_20873,N_19511);
nand U28532 (N_28532,N_20301,N_19584);
nor U28533 (N_28533,N_23177,N_22595);
nor U28534 (N_28534,N_20879,N_23970);
xor U28535 (N_28535,N_22261,N_21494);
nor U28536 (N_28536,N_20242,N_18764);
nor U28537 (N_28537,N_21120,N_23106);
nand U28538 (N_28538,N_19801,N_21203);
or U28539 (N_28539,N_20146,N_23374);
xnor U28540 (N_28540,N_21200,N_21352);
nor U28541 (N_28541,N_18522,N_23990);
nor U28542 (N_28542,N_21460,N_19355);
xor U28543 (N_28543,N_22715,N_23919);
nand U28544 (N_28544,N_22029,N_22764);
xnor U28545 (N_28545,N_23165,N_20065);
nor U28546 (N_28546,N_21770,N_18588);
or U28547 (N_28547,N_23479,N_23302);
and U28548 (N_28548,N_20191,N_19711);
and U28549 (N_28549,N_23885,N_21022);
xnor U28550 (N_28550,N_21455,N_21861);
xor U28551 (N_28551,N_21890,N_22657);
or U28552 (N_28552,N_18748,N_20896);
or U28553 (N_28553,N_22879,N_19398);
or U28554 (N_28554,N_23741,N_22096);
or U28555 (N_28555,N_20177,N_22931);
or U28556 (N_28556,N_18037,N_23895);
and U28557 (N_28557,N_18830,N_18754);
nor U28558 (N_28558,N_21982,N_21635);
and U28559 (N_28559,N_18945,N_18751);
xnor U28560 (N_28560,N_21922,N_21396);
nand U28561 (N_28561,N_23227,N_21349);
xnor U28562 (N_28562,N_19629,N_23581);
nand U28563 (N_28563,N_19376,N_20786);
xor U28564 (N_28564,N_22721,N_23799);
nor U28565 (N_28565,N_21892,N_21154);
or U28566 (N_28566,N_20124,N_23514);
and U28567 (N_28567,N_22711,N_22819);
nand U28568 (N_28568,N_18861,N_19515);
nor U28569 (N_28569,N_19105,N_20416);
xor U28570 (N_28570,N_18197,N_23875);
xor U28571 (N_28571,N_21277,N_23625);
or U28572 (N_28572,N_22809,N_20077);
nand U28573 (N_28573,N_22774,N_21404);
nor U28574 (N_28574,N_23056,N_19019);
or U28575 (N_28575,N_18182,N_21283);
and U28576 (N_28576,N_22410,N_23111);
xnor U28577 (N_28577,N_21006,N_20222);
nor U28578 (N_28578,N_20843,N_23977);
or U28579 (N_28579,N_18901,N_19838);
nand U28580 (N_28580,N_18078,N_23033);
or U28581 (N_28581,N_21797,N_21929);
xor U28582 (N_28582,N_18048,N_19947);
nor U28583 (N_28583,N_21341,N_20429);
xnor U28584 (N_28584,N_23620,N_21429);
nor U28585 (N_28585,N_20355,N_19244);
and U28586 (N_28586,N_19557,N_20229);
nand U28587 (N_28587,N_18412,N_18035);
xnor U28588 (N_28588,N_22016,N_22134);
or U28589 (N_28589,N_19027,N_20819);
nand U28590 (N_28590,N_21681,N_20255);
xor U28591 (N_28591,N_21180,N_23619);
and U28592 (N_28592,N_20601,N_19680);
or U28593 (N_28593,N_23186,N_18701);
nor U28594 (N_28594,N_20240,N_22169);
xnor U28595 (N_28595,N_22400,N_19466);
and U28596 (N_28596,N_21139,N_22982);
nor U28597 (N_28597,N_18435,N_22980);
nand U28598 (N_28598,N_19824,N_23853);
and U28599 (N_28599,N_20855,N_23826);
and U28600 (N_28600,N_22032,N_22613);
nand U28601 (N_28601,N_21331,N_20186);
xor U28602 (N_28602,N_19568,N_22036);
xnor U28603 (N_28603,N_18377,N_23760);
xnor U28604 (N_28604,N_20933,N_18246);
xnor U28605 (N_28605,N_20475,N_20523);
nand U28606 (N_28606,N_23530,N_23733);
xor U28607 (N_28607,N_19447,N_18321);
xnor U28608 (N_28608,N_18779,N_21567);
nand U28609 (N_28609,N_19673,N_19847);
and U28610 (N_28610,N_23874,N_23438);
nand U28611 (N_28611,N_19464,N_18800);
nand U28612 (N_28612,N_18624,N_18656);
nand U28613 (N_28613,N_19523,N_21646);
and U28614 (N_28614,N_20663,N_21631);
or U28615 (N_28615,N_21551,N_19054);
nand U28616 (N_28616,N_23219,N_21809);
nand U28617 (N_28617,N_21972,N_19301);
and U28618 (N_28618,N_22236,N_18892);
nor U28619 (N_28619,N_19979,N_18395);
or U28620 (N_28620,N_20728,N_19991);
nor U28621 (N_28621,N_19362,N_18516);
nor U28622 (N_28622,N_23745,N_18536);
and U28623 (N_28623,N_20405,N_20521);
or U28624 (N_28624,N_21570,N_21300);
or U28625 (N_28625,N_20855,N_18288);
nand U28626 (N_28626,N_20306,N_20591);
nand U28627 (N_28627,N_18140,N_19933);
and U28628 (N_28628,N_20804,N_22563);
and U28629 (N_28629,N_18410,N_20209);
nand U28630 (N_28630,N_19777,N_19535);
and U28631 (N_28631,N_21871,N_22131);
nor U28632 (N_28632,N_23328,N_20849);
nor U28633 (N_28633,N_22290,N_22288);
xnor U28634 (N_28634,N_21756,N_22773);
or U28635 (N_28635,N_20642,N_21702);
or U28636 (N_28636,N_23569,N_23119);
nand U28637 (N_28637,N_19469,N_20567);
xnor U28638 (N_28638,N_22895,N_23053);
nor U28639 (N_28639,N_20609,N_20987);
and U28640 (N_28640,N_22029,N_23386);
nor U28641 (N_28641,N_23098,N_20866);
and U28642 (N_28642,N_22070,N_20987);
nor U28643 (N_28643,N_21892,N_19866);
xor U28644 (N_28644,N_21225,N_23086);
and U28645 (N_28645,N_22215,N_18947);
nand U28646 (N_28646,N_21749,N_19261);
or U28647 (N_28647,N_22106,N_22132);
and U28648 (N_28648,N_22589,N_18009);
and U28649 (N_28649,N_23563,N_21415);
and U28650 (N_28650,N_23067,N_20242);
xor U28651 (N_28651,N_19565,N_21635);
xnor U28652 (N_28652,N_19584,N_19440);
and U28653 (N_28653,N_21218,N_18054);
nand U28654 (N_28654,N_23561,N_18358);
and U28655 (N_28655,N_22355,N_19748);
xnor U28656 (N_28656,N_23016,N_19178);
or U28657 (N_28657,N_23076,N_19800);
or U28658 (N_28658,N_23939,N_23471);
xor U28659 (N_28659,N_20023,N_19728);
or U28660 (N_28660,N_21612,N_18101);
or U28661 (N_28661,N_22859,N_23859);
or U28662 (N_28662,N_21308,N_19356);
nor U28663 (N_28663,N_21568,N_22308);
xnor U28664 (N_28664,N_21909,N_21654);
nor U28665 (N_28665,N_22982,N_21875);
nand U28666 (N_28666,N_19907,N_20633);
or U28667 (N_28667,N_20647,N_21266);
and U28668 (N_28668,N_20395,N_23451);
xor U28669 (N_28669,N_23782,N_22649);
nor U28670 (N_28670,N_22923,N_19176);
or U28671 (N_28671,N_22215,N_22657);
nand U28672 (N_28672,N_23492,N_18341);
nor U28673 (N_28673,N_21928,N_21535);
or U28674 (N_28674,N_18737,N_18453);
xnor U28675 (N_28675,N_20395,N_20688);
and U28676 (N_28676,N_20367,N_18256);
or U28677 (N_28677,N_20848,N_18547);
nor U28678 (N_28678,N_23248,N_21475);
or U28679 (N_28679,N_20823,N_18621);
xor U28680 (N_28680,N_18747,N_20199);
nand U28681 (N_28681,N_19415,N_20629);
nor U28682 (N_28682,N_21388,N_20665);
or U28683 (N_28683,N_18925,N_19296);
nor U28684 (N_28684,N_21827,N_22908);
or U28685 (N_28685,N_21238,N_21630);
xnor U28686 (N_28686,N_18945,N_20735);
xor U28687 (N_28687,N_22114,N_19653);
nor U28688 (N_28688,N_22798,N_18469);
nand U28689 (N_28689,N_20126,N_19298);
xor U28690 (N_28690,N_18742,N_20127);
and U28691 (N_28691,N_23409,N_23046);
xor U28692 (N_28692,N_19156,N_23223);
xnor U28693 (N_28693,N_18341,N_20445);
or U28694 (N_28694,N_22726,N_19639);
or U28695 (N_28695,N_23755,N_23857);
nor U28696 (N_28696,N_18224,N_21617);
xor U28697 (N_28697,N_21164,N_20161);
nand U28698 (N_28698,N_21653,N_21730);
nor U28699 (N_28699,N_22583,N_20276);
nand U28700 (N_28700,N_21732,N_18136);
nor U28701 (N_28701,N_20443,N_19444);
and U28702 (N_28702,N_22600,N_20327);
nor U28703 (N_28703,N_22566,N_21567);
or U28704 (N_28704,N_20071,N_21939);
nor U28705 (N_28705,N_19600,N_18234);
and U28706 (N_28706,N_23268,N_22673);
and U28707 (N_28707,N_19712,N_20582);
nand U28708 (N_28708,N_22261,N_18605);
xor U28709 (N_28709,N_22873,N_18359);
or U28710 (N_28710,N_23585,N_18697);
nand U28711 (N_28711,N_20752,N_23109);
nand U28712 (N_28712,N_22154,N_19072);
nand U28713 (N_28713,N_19245,N_19654);
or U28714 (N_28714,N_21392,N_20146);
or U28715 (N_28715,N_18101,N_19513);
or U28716 (N_28716,N_19882,N_21634);
or U28717 (N_28717,N_19990,N_22774);
nor U28718 (N_28718,N_18477,N_21892);
xor U28719 (N_28719,N_22836,N_20562);
and U28720 (N_28720,N_19927,N_23512);
and U28721 (N_28721,N_23619,N_22640);
xnor U28722 (N_28722,N_21760,N_23774);
nor U28723 (N_28723,N_23384,N_18671);
and U28724 (N_28724,N_21836,N_19771);
or U28725 (N_28725,N_20708,N_20611);
xnor U28726 (N_28726,N_22723,N_18895);
xnor U28727 (N_28727,N_19681,N_22551);
xor U28728 (N_28728,N_18868,N_19217);
or U28729 (N_28729,N_21186,N_21488);
nand U28730 (N_28730,N_20270,N_23392);
nand U28731 (N_28731,N_18829,N_20554);
nor U28732 (N_28732,N_20011,N_23407);
xnor U28733 (N_28733,N_21154,N_21809);
xnor U28734 (N_28734,N_21697,N_20209);
and U28735 (N_28735,N_18183,N_19728);
nand U28736 (N_28736,N_18337,N_20918);
or U28737 (N_28737,N_20744,N_22043);
nand U28738 (N_28738,N_18390,N_18057);
nor U28739 (N_28739,N_20030,N_23551);
xor U28740 (N_28740,N_22428,N_22679);
nand U28741 (N_28741,N_21912,N_22214);
nand U28742 (N_28742,N_18138,N_18600);
xor U28743 (N_28743,N_20284,N_19301);
nand U28744 (N_28744,N_22951,N_18451);
xnor U28745 (N_28745,N_20735,N_21838);
nand U28746 (N_28746,N_19000,N_22459);
xor U28747 (N_28747,N_22834,N_22667);
nand U28748 (N_28748,N_23157,N_23326);
nand U28749 (N_28749,N_18866,N_23980);
nand U28750 (N_28750,N_18375,N_22631);
nand U28751 (N_28751,N_18590,N_18538);
xor U28752 (N_28752,N_20729,N_21516);
and U28753 (N_28753,N_21379,N_18039);
or U28754 (N_28754,N_19730,N_18219);
or U28755 (N_28755,N_22242,N_18068);
nand U28756 (N_28756,N_21847,N_19607);
xnor U28757 (N_28757,N_19178,N_23111);
nor U28758 (N_28758,N_21285,N_18147);
nor U28759 (N_28759,N_21316,N_21561);
or U28760 (N_28760,N_21687,N_21307);
xnor U28761 (N_28761,N_19349,N_21579);
nor U28762 (N_28762,N_18961,N_19249);
nand U28763 (N_28763,N_22109,N_21659);
or U28764 (N_28764,N_18147,N_22484);
nor U28765 (N_28765,N_18667,N_19005);
and U28766 (N_28766,N_18114,N_18024);
and U28767 (N_28767,N_23434,N_20934);
or U28768 (N_28768,N_20341,N_21587);
nor U28769 (N_28769,N_20677,N_22338);
nor U28770 (N_28770,N_20511,N_18496);
and U28771 (N_28771,N_18504,N_22515);
nand U28772 (N_28772,N_18382,N_23609);
xnor U28773 (N_28773,N_23528,N_19313);
xnor U28774 (N_28774,N_21230,N_21151);
nand U28775 (N_28775,N_20278,N_20025);
and U28776 (N_28776,N_20810,N_23602);
or U28777 (N_28777,N_20026,N_21939);
and U28778 (N_28778,N_18408,N_22735);
nand U28779 (N_28779,N_18863,N_19796);
nand U28780 (N_28780,N_21072,N_18811);
and U28781 (N_28781,N_23616,N_19919);
nor U28782 (N_28782,N_19825,N_20824);
or U28783 (N_28783,N_22780,N_21389);
and U28784 (N_28784,N_21132,N_23666);
and U28785 (N_28785,N_22779,N_20131);
xor U28786 (N_28786,N_23583,N_19848);
or U28787 (N_28787,N_22104,N_20016);
nand U28788 (N_28788,N_20180,N_21648);
xor U28789 (N_28789,N_23931,N_22433);
nand U28790 (N_28790,N_22794,N_23150);
nand U28791 (N_28791,N_22872,N_22980);
nor U28792 (N_28792,N_19430,N_20313);
or U28793 (N_28793,N_20681,N_22960);
xnor U28794 (N_28794,N_18446,N_19125);
or U28795 (N_28795,N_21705,N_21855);
or U28796 (N_28796,N_22379,N_20698);
xnor U28797 (N_28797,N_21359,N_19997);
nand U28798 (N_28798,N_22288,N_20773);
and U28799 (N_28799,N_19348,N_18337);
and U28800 (N_28800,N_22708,N_21551);
xnor U28801 (N_28801,N_23006,N_20730);
or U28802 (N_28802,N_23835,N_21030);
nor U28803 (N_28803,N_21131,N_21908);
xnor U28804 (N_28804,N_21221,N_20745);
nand U28805 (N_28805,N_19391,N_21551);
or U28806 (N_28806,N_19096,N_22040);
xnor U28807 (N_28807,N_18103,N_20143);
and U28808 (N_28808,N_20872,N_19559);
xnor U28809 (N_28809,N_21738,N_19356);
nor U28810 (N_28810,N_20626,N_21441);
or U28811 (N_28811,N_23358,N_18184);
xor U28812 (N_28812,N_22052,N_21980);
nand U28813 (N_28813,N_23045,N_22901);
and U28814 (N_28814,N_22595,N_23521);
nor U28815 (N_28815,N_22776,N_20539);
or U28816 (N_28816,N_20100,N_23689);
nand U28817 (N_28817,N_19793,N_18125);
nor U28818 (N_28818,N_22681,N_22882);
nand U28819 (N_28819,N_21832,N_23752);
nor U28820 (N_28820,N_23448,N_22761);
or U28821 (N_28821,N_23461,N_23469);
nor U28822 (N_28822,N_21014,N_23800);
xor U28823 (N_28823,N_21909,N_20467);
nand U28824 (N_28824,N_21105,N_22067);
nor U28825 (N_28825,N_18190,N_20485);
nor U28826 (N_28826,N_23080,N_18083);
or U28827 (N_28827,N_21796,N_21424);
nand U28828 (N_28828,N_21132,N_20504);
or U28829 (N_28829,N_22820,N_19991);
nor U28830 (N_28830,N_22688,N_20602);
nor U28831 (N_28831,N_18564,N_22743);
or U28832 (N_28832,N_21080,N_21475);
and U28833 (N_28833,N_18343,N_22618);
nand U28834 (N_28834,N_20937,N_18063);
or U28835 (N_28835,N_23711,N_20226);
nand U28836 (N_28836,N_22782,N_22506);
nand U28837 (N_28837,N_19398,N_21157);
nand U28838 (N_28838,N_21174,N_18975);
nand U28839 (N_28839,N_20776,N_21623);
xnor U28840 (N_28840,N_19731,N_22902);
nor U28841 (N_28841,N_23588,N_21859);
and U28842 (N_28842,N_18631,N_18179);
or U28843 (N_28843,N_22108,N_22625);
nand U28844 (N_28844,N_19805,N_18870);
and U28845 (N_28845,N_19788,N_19172);
or U28846 (N_28846,N_21896,N_18968);
or U28847 (N_28847,N_22317,N_20898);
and U28848 (N_28848,N_20620,N_18931);
nor U28849 (N_28849,N_19762,N_21946);
nand U28850 (N_28850,N_23227,N_22120);
nor U28851 (N_28851,N_23982,N_22134);
nor U28852 (N_28852,N_23641,N_22066);
xnor U28853 (N_28853,N_21122,N_20624);
or U28854 (N_28854,N_21889,N_19599);
xnor U28855 (N_28855,N_19909,N_23750);
nand U28856 (N_28856,N_19756,N_21296);
nor U28857 (N_28857,N_18088,N_19930);
nand U28858 (N_28858,N_18286,N_18676);
and U28859 (N_28859,N_23206,N_19268);
and U28860 (N_28860,N_22354,N_21832);
nand U28861 (N_28861,N_21596,N_21908);
and U28862 (N_28862,N_23494,N_21757);
xnor U28863 (N_28863,N_23072,N_18888);
or U28864 (N_28864,N_19980,N_20463);
and U28865 (N_28865,N_22429,N_22670);
nand U28866 (N_28866,N_20773,N_23307);
and U28867 (N_28867,N_22241,N_23051);
nand U28868 (N_28868,N_21266,N_19421);
nor U28869 (N_28869,N_18914,N_19758);
xor U28870 (N_28870,N_19882,N_22495);
and U28871 (N_28871,N_19659,N_18159);
and U28872 (N_28872,N_23323,N_20174);
and U28873 (N_28873,N_18755,N_22231);
nor U28874 (N_28874,N_21538,N_21929);
or U28875 (N_28875,N_18861,N_19616);
nand U28876 (N_28876,N_18100,N_18078);
or U28877 (N_28877,N_22681,N_23155);
nor U28878 (N_28878,N_21011,N_22274);
or U28879 (N_28879,N_21518,N_19527);
xor U28880 (N_28880,N_21564,N_22990);
or U28881 (N_28881,N_20744,N_19766);
xor U28882 (N_28882,N_19531,N_23947);
xnor U28883 (N_28883,N_21684,N_21678);
nand U28884 (N_28884,N_19847,N_23631);
nand U28885 (N_28885,N_22289,N_20813);
xor U28886 (N_28886,N_19773,N_22361);
and U28887 (N_28887,N_18352,N_19631);
xor U28888 (N_28888,N_18026,N_19706);
or U28889 (N_28889,N_23615,N_20310);
nor U28890 (N_28890,N_21006,N_18873);
and U28891 (N_28891,N_18007,N_18076);
xor U28892 (N_28892,N_20194,N_20377);
nor U28893 (N_28893,N_20073,N_21793);
and U28894 (N_28894,N_23281,N_23091);
and U28895 (N_28895,N_21263,N_22039);
or U28896 (N_28896,N_21483,N_22869);
nand U28897 (N_28897,N_23694,N_18309);
xor U28898 (N_28898,N_21082,N_22057);
nor U28899 (N_28899,N_23013,N_19530);
and U28900 (N_28900,N_18564,N_18769);
nand U28901 (N_28901,N_18037,N_23034);
or U28902 (N_28902,N_23085,N_18318);
xnor U28903 (N_28903,N_19653,N_21195);
nor U28904 (N_28904,N_19025,N_21718);
and U28905 (N_28905,N_22023,N_23598);
xor U28906 (N_28906,N_20652,N_19444);
nor U28907 (N_28907,N_22666,N_18588);
nor U28908 (N_28908,N_22454,N_22243);
nand U28909 (N_28909,N_18212,N_19829);
nand U28910 (N_28910,N_18855,N_20956);
and U28911 (N_28911,N_18449,N_21023);
and U28912 (N_28912,N_22828,N_21561);
xor U28913 (N_28913,N_18369,N_20447);
xor U28914 (N_28914,N_19805,N_18200);
and U28915 (N_28915,N_19531,N_19061);
xnor U28916 (N_28916,N_20017,N_18688);
nand U28917 (N_28917,N_21246,N_23815);
and U28918 (N_28918,N_18169,N_19674);
or U28919 (N_28919,N_20140,N_22079);
nor U28920 (N_28920,N_22923,N_20188);
or U28921 (N_28921,N_20329,N_20735);
or U28922 (N_28922,N_18563,N_19414);
nor U28923 (N_28923,N_18857,N_20113);
xor U28924 (N_28924,N_22002,N_21140);
nor U28925 (N_28925,N_23556,N_19202);
nor U28926 (N_28926,N_20840,N_22963);
xor U28927 (N_28927,N_22732,N_19905);
xor U28928 (N_28928,N_22403,N_20093);
nor U28929 (N_28929,N_19720,N_20349);
or U28930 (N_28930,N_22998,N_21244);
xor U28931 (N_28931,N_18184,N_20678);
xor U28932 (N_28932,N_22334,N_23488);
xor U28933 (N_28933,N_22772,N_23050);
xor U28934 (N_28934,N_18639,N_23907);
or U28935 (N_28935,N_18921,N_21134);
and U28936 (N_28936,N_23339,N_21274);
nand U28937 (N_28937,N_22149,N_23382);
or U28938 (N_28938,N_21664,N_23039);
and U28939 (N_28939,N_23903,N_21519);
or U28940 (N_28940,N_22139,N_18990);
or U28941 (N_28941,N_18249,N_22916);
xor U28942 (N_28942,N_21496,N_23882);
xnor U28943 (N_28943,N_20201,N_21547);
and U28944 (N_28944,N_20123,N_20481);
nand U28945 (N_28945,N_21102,N_21127);
nand U28946 (N_28946,N_22969,N_20347);
or U28947 (N_28947,N_20166,N_22430);
or U28948 (N_28948,N_19293,N_22330);
nand U28949 (N_28949,N_19463,N_20118);
xnor U28950 (N_28950,N_23576,N_23350);
and U28951 (N_28951,N_21170,N_18085);
or U28952 (N_28952,N_21084,N_20505);
and U28953 (N_28953,N_23080,N_23899);
nand U28954 (N_28954,N_20504,N_18469);
nand U28955 (N_28955,N_20361,N_22917);
nor U28956 (N_28956,N_19667,N_18897);
nand U28957 (N_28957,N_22050,N_18698);
nand U28958 (N_28958,N_20374,N_18936);
nor U28959 (N_28959,N_20368,N_19907);
nand U28960 (N_28960,N_19071,N_21563);
nor U28961 (N_28961,N_20988,N_22170);
or U28962 (N_28962,N_20965,N_21858);
nand U28963 (N_28963,N_19572,N_21183);
and U28964 (N_28964,N_23982,N_20397);
or U28965 (N_28965,N_21091,N_23069);
or U28966 (N_28966,N_18725,N_21319);
and U28967 (N_28967,N_20055,N_20517);
xor U28968 (N_28968,N_23166,N_18340);
xnor U28969 (N_28969,N_20741,N_18857);
nor U28970 (N_28970,N_20727,N_23714);
xor U28971 (N_28971,N_20752,N_19688);
and U28972 (N_28972,N_23483,N_23787);
xor U28973 (N_28973,N_22720,N_18415);
or U28974 (N_28974,N_21709,N_23772);
nand U28975 (N_28975,N_18140,N_18255);
nand U28976 (N_28976,N_21501,N_23136);
xnor U28977 (N_28977,N_23588,N_22736);
and U28978 (N_28978,N_23555,N_21302);
xnor U28979 (N_28979,N_21466,N_23577);
and U28980 (N_28980,N_20631,N_22041);
and U28981 (N_28981,N_23228,N_21574);
or U28982 (N_28982,N_21262,N_19972);
and U28983 (N_28983,N_18621,N_23557);
and U28984 (N_28984,N_19020,N_21353);
nor U28985 (N_28985,N_18234,N_21906);
xnor U28986 (N_28986,N_18982,N_23338);
nand U28987 (N_28987,N_23729,N_19954);
or U28988 (N_28988,N_18774,N_21625);
or U28989 (N_28989,N_21955,N_23111);
nand U28990 (N_28990,N_20032,N_20271);
xor U28991 (N_28991,N_18699,N_21865);
or U28992 (N_28992,N_21513,N_18676);
and U28993 (N_28993,N_23507,N_18085);
nand U28994 (N_28994,N_22141,N_20858);
nand U28995 (N_28995,N_23912,N_20030);
and U28996 (N_28996,N_23098,N_21590);
and U28997 (N_28997,N_23413,N_19321);
nor U28998 (N_28998,N_21429,N_22962);
xnor U28999 (N_28999,N_22839,N_22808);
nor U29000 (N_29000,N_21132,N_20871);
and U29001 (N_29001,N_21879,N_18005);
and U29002 (N_29002,N_23578,N_20623);
and U29003 (N_29003,N_21130,N_22802);
xor U29004 (N_29004,N_23979,N_21791);
or U29005 (N_29005,N_20968,N_18037);
nor U29006 (N_29006,N_19137,N_22953);
nand U29007 (N_29007,N_20070,N_20677);
nor U29008 (N_29008,N_20185,N_20258);
or U29009 (N_29009,N_19301,N_19600);
nand U29010 (N_29010,N_19122,N_21418);
nand U29011 (N_29011,N_21896,N_22420);
xor U29012 (N_29012,N_18852,N_19116);
nor U29013 (N_29013,N_21414,N_19887);
or U29014 (N_29014,N_22504,N_18704);
or U29015 (N_29015,N_19863,N_23144);
or U29016 (N_29016,N_20281,N_23911);
nor U29017 (N_29017,N_23323,N_22568);
nand U29018 (N_29018,N_20015,N_23933);
or U29019 (N_29019,N_23302,N_22941);
nand U29020 (N_29020,N_18958,N_20118);
and U29021 (N_29021,N_22881,N_22194);
or U29022 (N_29022,N_22526,N_23927);
and U29023 (N_29023,N_20477,N_18364);
xor U29024 (N_29024,N_21759,N_19586);
xnor U29025 (N_29025,N_21693,N_20749);
nor U29026 (N_29026,N_18713,N_20092);
nor U29027 (N_29027,N_19110,N_22218);
and U29028 (N_29028,N_19329,N_20924);
xnor U29029 (N_29029,N_20407,N_18045);
xnor U29030 (N_29030,N_20754,N_23467);
or U29031 (N_29031,N_18199,N_23511);
xor U29032 (N_29032,N_19267,N_22333);
nor U29033 (N_29033,N_23330,N_22231);
xor U29034 (N_29034,N_23901,N_19746);
nor U29035 (N_29035,N_20741,N_20082);
xnor U29036 (N_29036,N_23138,N_19310);
xnor U29037 (N_29037,N_18628,N_21825);
nor U29038 (N_29038,N_20468,N_18153);
nor U29039 (N_29039,N_19902,N_20407);
or U29040 (N_29040,N_18543,N_19139);
and U29041 (N_29041,N_20097,N_23826);
or U29042 (N_29042,N_22883,N_19845);
or U29043 (N_29043,N_19641,N_21722);
xnor U29044 (N_29044,N_22146,N_23386);
xnor U29045 (N_29045,N_20767,N_19457);
or U29046 (N_29046,N_21739,N_22250);
xor U29047 (N_29047,N_19787,N_19002);
nand U29048 (N_29048,N_23437,N_19597);
nand U29049 (N_29049,N_19381,N_18532);
nor U29050 (N_29050,N_23823,N_21034);
and U29051 (N_29051,N_23633,N_18180);
or U29052 (N_29052,N_22170,N_23250);
or U29053 (N_29053,N_18282,N_19671);
nor U29054 (N_29054,N_21299,N_20777);
and U29055 (N_29055,N_23514,N_18403);
or U29056 (N_29056,N_19558,N_20630);
xnor U29057 (N_29057,N_20918,N_23939);
nand U29058 (N_29058,N_20710,N_18239);
xor U29059 (N_29059,N_23555,N_18468);
xor U29060 (N_29060,N_22159,N_19373);
xnor U29061 (N_29061,N_20226,N_20822);
and U29062 (N_29062,N_22435,N_19931);
and U29063 (N_29063,N_18721,N_20561);
nand U29064 (N_29064,N_22407,N_21606);
or U29065 (N_29065,N_18227,N_19519);
nand U29066 (N_29066,N_20491,N_19072);
and U29067 (N_29067,N_18197,N_19817);
nand U29068 (N_29068,N_20524,N_20825);
and U29069 (N_29069,N_19837,N_20156);
nor U29070 (N_29070,N_20031,N_19783);
and U29071 (N_29071,N_20520,N_22543);
or U29072 (N_29072,N_20488,N_23094);
nor U29073 (N_29073,N_18336,N_23218);
nand U29074 (N_29074,N_21061,N_19552);
nor U29075 (N_29075,N_18851,N_21502);
xor U29076 (N_29076,N_23173,N_20730);
and U29077 (N_29077,N_20167,N_20079);
nand U29078 (N_29078,N_20415,N_21872);
and U29079 (N_29079,N_23011,N_20200);
xnor U29080 (N_29080,N_23786,N_23130);
nand U29081 (N_29081,N_20312,N_23641);
nor U29082 (N_29082,N_20540,N_22415);
nand U29083 (N_29083,N_23674,N_18306);
xnor U29084 (N_29084,N_22525,N_18804);
xor U29085 (N_29085,N_21707,N_23110);
xor U29086 (N_29086,N_23546,N_18387);
and U29087 (N_29087,N_22946,N_21274);
nor U29088 (N_29088,N_23764,N_20859);
nor U29089 (N_29089,N_22349,N_18228);
or U29090 (N_29090,N_23325,N_20740);
nand U29091 (N_29091,N_18339,N_22330);
xor U29092 (N_29092,N_22331,N_22037);
nor U29093 (N_29093,N_21694,N_21082);
or U29094 (N_29094,N_18804,N_21927);
nor U29095 (N_29095,N_22869,N_22999);
nor U29096 (N_29096,N_21485,N_18653);
nand U29097 (N_29097,N_22847,N_22612);
and U29098 (N_29098,N_23844,N_21547);
or U29099 (N_29099,N_19773,N_19930);
xnor U29100 (N_29100,N_22252,N_21009);
nand U29101 (N_29101,N_20316,N_23352);
xor U29102 (N_29102,N_22073,N_20714);
xor U29103 (N_29103,N_23220,N_22161);
nor U29104 (N_29104,N_19611,N_18134);
xnor U29105 (N_29105,N_19687,N_22344);
nand U29106 (N_29106,N_22764,N_20935);
nand U29107 (N_29107,N_23784,N_21480);
xnor U29108 (N_29108,N_20370,N_21509);
nand U29109 (N_29109,N_20028,N_18051);
xor U29110 (N_29110,N_23875,N_23405);
nor U29111 (N_29111,N_19336,N_19061);
or U29112 (N_29112,N_23942,N_22873);
or U29113 (N_29113,N_21090,N_22976);
nand U29114 (N_29114,N_20225,N_21672);
xor U29115 (N_29115,N_19905,N_21258);
or U29116 (N_29116,N_23678,N_19615);
or U29117 (N_29117,N_22991,N_19529);
and U29118 (N_29118,N_22195,N_19221);
and U29119 (N_29119,N_22138,N_19087);
nor U29120 (N_29120,N_18155,N_20566);
nand U29121 (N_29121,N_18679,N_20913);
nor U29122 (N_29122,N_21261,N_18084);
or U29123 (N_29123,N_22033,N_20146);
or U29124 (N_29124,N_19320,N_21550);
nor U29125 (N_29125,N_23248,N_23110);
nand U29126 (N_29126,N_22603,N_20917);
or U29127 (N_29127,N_23257,N_22635);
nand U29128 (N_29128,N_20957,N_20913);
and U29129 (N_29129,N_20899,N_21601);
nand U29130 (N_29130,N_23722,N_20808);
and U29131 (N_29131,N_19011,N_22595);
nand U29132 (N_29132,N_18778,N_19447);
nor U29133 (N_29133,N_19877,N_22894);
xnor U29134 (N_29134,N_23070,N_21869);
and U29135 (N_29135,N_21234,N_19332);
and U29136 (N_29136,N_22606,N_19828);
nor U29137 (N_29137,N_21369,N_22797);
nand U29138 (N_29138,N_20540,N_18480);
and U29139 (N_29139,N_22564,N_18592);
nand U29140 (N_29140,N_22926,N_20605);
or U29141 (N_29141,N_22037,N_20749);
and U29142 (N_29142,N_21466,N_20112);
or U29143 (N_29143,N_22834,N_21664);
and U29144 (N_29144,N_22617,N_22549);
or U29145 (N_29145,N_18223,N_19163);
nand U29146 (N_29146,N_19250,N_21302);
nand U29147 (N_29147,N_19927,N_20605);
or U29148 (N_29148,N_20708,N_20128);
and U29149 (N_29149,N_22866,N_21695);
nor U29150 (N_29150,N_19477,N_23427);
and U29151 (N_29151,N_18580,N_23852);
nand U29152 (N_29152,N_19753,N_18604);
xnor U29153 (N_29153,N_18667,N_22144);
nand U29154 (N_29154,N_23127,N_22975);
and U29155 (N_29155,N_23353,N_23032);
and U29156 (N_29156,N_20026,N_22646);
and U29157 (N_29157,N_22365,N_18874);
and U29158 (N_29158,N_23031,N_20469);
or U29159 (N_29159,N_19454,N_18731);
and U29160 (N_29160,N_18432,N_20198);
nand U29161 (N_29161,N_23259,N_18852);
or U29162 (N_29162,N_19126,N_19586);
or U29163 (N_29163,N_23503,N_22758);
nand U29164 (N_29164,N_20814,N_18226);
nand U29165 (N_29165,N_21150,N_23227);
or U29166 (N_29166,N_22103,N_23346);
or U29167 (N_29167,N_21978,N_18544);
or U29168 (N_29168,N_20037,N_21191);
or U29169 (N_29169,N_20750,N_22402);
or U29170 (N_29170,N_20744,N_22711);
xnor U29171 (N_29171,N_19550,N_22180);
or U29172 (N_29172,N_22061,N_20561);
nand U29173 (N_29173,N_20535,N_18918);
and U29174 (N_29174,N_19807,N_20894);
nor U29175 (N_29175,N_22792,N_20464);
or U29176 (N_29176,N_23773,N_20190);
nor U29177 (N_29177,N_22404,N_23183);
nand U29178 (N_29178,N_23245,N_19319);
xnor U29179 (N_29179,N_18187,N_21757);
xnor U29180 (N_29180,N_19422,N_22537);
nand U29181 (N_29181,N_18011,N_22579);
and U29182 (N_29182,N_19366,N_20313);
nand U29183 (N_29183,N_22692,N_22914);
or U29184 (N_29184,N_20132,N_20544);
or U29185 (N_29185,N_23469,N_22433);
or U29186 (N_29186,N_22852,N_18766);
nor U29187 (N_29187,N_19596,N_23236);
and U29188 (N_29188,N_21170,N_21225);
xor U29189 (N_29189,N_19864,N_21528);
nor U29190 (N_29190,N_22676,N_20093);
xor U29191 (N_29191,N_23875,N_21714);
and U29192 (N_29192,N_19858,N_18085);
or U29193 (N_29193,N_20314,N_19501);
and U29194 (N_29194,N_18641,N_21420);
and U29195 (N_29195,N_22192,N_19262);
or U29196 (N_29196,N_23220,N_21757);
nor U29197 (N_29197,N_19091,N_20185);
nand U29198 (N_29198,N_21063,N_23785);
xnor U29199 (N_29199,N_21381,N_21776);
nor U29200 (N_29200,N_21637,N_23415);
or U29201 (N_29201,N_22005,N_19995);
nand U29202 (N_29202,N_23595,N_21417);
and U29203 (N_29203,N_19777,N_22990);
and U29204 (N_29204,N_23727,N_19274);
xnor U29205 (N_29205,N_22435,N_23648);
nor U29206 (N_29206,N_18290,N_20583);
and U29207 (N_29207,N_23921,N_20046);
and U29208 (N_29208,N_18776,N_21036);
xor U29209 (N_29209,N_22227,N_18234);
xor U29210 (N_29210,N_22304,N_22138);
or U29211 (N_29211,N_20075,N_20324);
nand U29212 (N_29212,N_22878,N_22397);
and U29213 (N_29213,N_18938,N_21082);
nor U29214 (N_29214,N_19047,N_18005);
or U29215 (N_29215,N_23641,N_18955);
or U29216 (N_29216,N_21110,N_21218);
nor U29217 (N_29217,N_21069,N_19283);
nand U29218 (N_29218,N_20618,N_20398);
and U29219 (N_29219,N_22164,N_23253);
nor U29220 (N_29220,N_22919,N_19999);
nand U29221 (N_29221,N_22112,N_21492);
nand U29222 (N_29222,N_23611,N_20580);
or U29223 (N_29223,N_21070,N_23927);
nand U29224 (N_29224,N_20752,N_18674);
nor U29225 (N_29225,N_18297,N_23176);
nor U29226 (N_29226,N_19982,N_19352);
and U29227 (N_29227,N_20780,N_18532);
nor U29228 (N_29228,N_19091,N_22871);
xor U29229 (N_29229,N_21531,N_22696);
nand U29230 (N_29230,N_18448,N_20026);
xor U29231 (N_29231,N_20512,N_22368);
or U29232 (N_29232,N_19114,N_19139);
nand U29233 (N_29233,N_19655,N_19654);
nand U29234 (N_29234,N_18193,N_19116);
nand U29235 (N_29235,N_19468,N_22341);
nand U29236 (N_29236,N_22058,N_19831);
xor U29237 (N_29237,N_19410,N_21878);
xnor U29238 (N_29238,N_18293,N_21853);
nor U29239 (N_29239,N_21840,N_21580);
nand U29240 (N_29240,N_18375,N_19139);
nand U29241 (N_29241,N_18258,N_23213);
xnor U29242 (N_29242,N_23932,N_23725);
or U29243 (N_29243,N_22447,N_18512);
or U29244 (N_29244,N_22239,N_20644);
nor U29245 (N_29245,N_22870,N_21039);
nor U29246 (N_29246,N_21469,N_19221);
and U29247 (N_29247,N_22447,N_23068);
nor U29248 (N_29248,N_22442,N_19979);
nand U29249 (N_29249,N_19778,N_18108);
and U29250 (N_29250,N_21551,N_23501);
nand U29251 (N_29251,N_22800,N_20888);
or U29252 (N_29252,N_19128,N_22003);
nand U29253 (N_29253,N_23912,N_20589);
xor U29254 (N_29254,N_18587,N_18528);
nand U29255 (N_29255,N_18216,N_23728);
xnor U29256 (N_29256,N_20350,N_20496);
nand U29257 (N_29257,N_23202,N_20636);
xor U29258 (N_29258,N_22973,N_20036);
or U29259 (N_29259,N_22529,N_18213);
xnor U29260 (N_29260,N_21716,N_22299);
or U29261 (N_29261,N_18863,N_21631);
and U29262 (N_29262,N_19932,N_22399);
or U29263 (N_29263,N_22261,N_22386);
xor U29264 (N_29264,N_20820,N_18180);
and U29265 (N_29265,N_21881,N_23909);
nor U29266 (N_29266,N_23212,N_23305);
nor U29267 (N_29267,N_21790,N_22564);
xor U29268 (N_29268,N_22195,N_23139);
and U29269 (N_29269,N_23694,N_23161);
xnor U29270 (N_29270,N_20160,N_19364);
nor U29271 (N_29271,N_22539,N_19953);
nor U29272 (N_29272,N_18417,N_18805);
and U29273 (N_29273,N_18523,N_23340);
or U29274 (N_29274,N_19798,N_20246);
nand U29275 (N_29275,N_19530,N_23304);
and U29276 (N_29276,N_18393,N_18893);
nand U29277 (N_29277,N_19894,N_22517);
xnor U29278 (N_29278,N_21715,N_22567);
and U29279 (N_29279,N_21301,N_21547);
or U29280 (N_29280,N_19927,N_20787);
xnor U29281 (N_29281,N_18195,N_19052);
xor U29282 (N_29282,N_19065,N_21065);
nand U29283 (N_29283,N_19772,N_19309);
or U29284 (N_29284,N_22772,N_20222);
and U29285 (N_29285,N_18595,N_22985);
xor U29286 (N_29286,N_19334,N_22577);
nand U29287 (N_29287,N_19919,N_23992);
nor U29288 (N_29288,N_19751,N_18660);
or U29289 (N_29289,N_23327,N_21390);
or U29290 (N_29290,N_23010,N_18953);
nor U29291 (N_29291,N_19695,N_23417);
nand U29292 (N_29292,N_20288,N_19953);
nor U29293 (N_29293,N_18163,N_21183);
and U29294 (N_29294,N_23818,N_23626);
xor U29295 (N_29295,N_22802,N_19705);
and U29296 (N_29296,N_21376,N_20068);
nor U29297 (N_29297,N_22007,N_23130);
nor U29298 (N_29298,N_18572,N_21994);
and U29299 (N_29299,N_19924,N_22092);
nor U29300 (N_29300,N_20759,N_23527);
and U29301 (N_29301,N_22166,N_21336);
nor U29302 (N_29302,N_20473,N_21493);
xor U29303 (N_29303,N_20374,N_23613);
nor U29304 (N_29304,N_22344,N_22889);
xor U29305 (N_29305,N_19785,N_21295);
nand U29306 (N_29306,N_21147,N_19577);
nor U29307 (N_29307,N_19742,N_18902);
xor U29308 (N_29308,N_23841,N_18707);
xor U29309 (N_29309,N_18548,N_19821);
xnor U29310 (N_29310,N_19384,N_19167);
xor U29311 (N_29311,N_20444,N_20221);
or U29312 (N_29312,N_22636,N_19067);
xnor U29313 (N_29313,N_19883,N_20567);
nand U29314 (N_29314,N_19958,N_23441);
xnor U29315 (N_29315,N_21336,N_19668);
and U29316 (N_29316,N_22869,N_22619);
or U29317 (N_29317,N_22220,N_18768);
nand U29318 (N_29318,N_18795,N_18685);
nand U29319 (N_29319,N_19298,N_20997);
or U29320 (N_29320,N_20756,N_18795);
and U29321 (N_29321,N_20398,N_22537);
xor U29322 (N_29322,N_20208,N_18639);
xor U29323 (N_29323,N_21714,N_21625);
or U29324 (N_29324,N_22531,N_19304);
xor U29325 (N_29325,N_18968,N_18951);
and U29326 (N_29326,N_21059,N_19447);
nor U29327 (N_29327,N_19768,N_21137);
nor U29328 (N_29328,N_22464,N_21154);
xor U29329 (N_29329,N_21025,N_22031);
nand U29330 (N_29330,N_21210,N_19661);
or U29331 (N_29331,N_20184,N_23869);
nor U29332 (N_29332,N_20407,N_22830);
nand U29333 (N_29333,N_18493,N_23670);
and U29334 (N_29334,N_19751,N_19069);
and U29335 (N_29335,N_18159,N_19296);
or U29336 (N_29336,N_20242,N_23780);
nand U29337 (N_29337,N_23193,N_21827);
and U29338 (N_29338,N_19339,N_22467);
xnor U29339 (N_29339,N_19227,N_23648);
or U29340 (N_29340,N_22528,N_21786);
xnor U29341 (N_29341,N_21314,N_22858);
xor U29342 (N_29342,N_19119,N_23778);
nand U29343 (N_29343,N_20918,N_20616);
and U29344 (N_29344,N_21492,N_23295);
or U29345 (N_29345,N_22558,N_18196);
nor U29346 (N_29346,N_22772,N_22734);
nand U29347 (N_29347,N_21128,N_21798);
or U29348 (N_29348,N_18225,N_23665);
nor U29349 (N_29349,N_19930,N_18547);
or U29350 (N_29350,N_19095,N_18781);
nor U29351 (N_29351,N_23079,N_20776);
or U29352 (N_29352,N_20023,N_18404);
xnor U29353 (N_29353,N_20832,N_18356);
nand U29354 (N_29354,N_21337,N_19046);
nand U29355 (N_29355,N_23271,N_18321);
xor U29356 (N_29356,N_18163,N_23700);
nand U29357 (N_29357,N_18926,N_21664);
or U29358 (N_29358,N_19694,N_22487);
nor U29359 (N_29359,N_22009,N_20360);
xor U29360 (N_29360,N_21391,N_18268);
nor U29361 (N_29361,N_18092,N_19356);
nand U29362 (N_29362,N_20723,N_20681);
and U29363 (N_29363,N_22794,N_21143);
xnor U29364 (N_29364,N_21002,N_18723);
nor U29365 (N_29365,N_21675,N_19769);
and U29366 (N_29366,N_22751,N_22012);
and U29367 (N_29367,N_23228,N_20175);
or U29368 (N_29368,N_21371,N_23764);
nand U29369 (N_29369,N_20206,N_23281);
xor U29370 (N_29370,N_21769,N_23977);
xor U29371 (N_29371,N_23582,N_22881);
nand U29372 (N_29372,N_18090,N_23883);
xnor U29373 (N_29373,N_19336,N_19784);
xor U29374 (N_29374,N_18196,N_18411);
and U29375 (N_29375,N_20889,N_19736);
nand U29376 (N_29376,N_18283,N_20772);
nor U29377 (N_29377,N_21671,N_19914);
and U29378 (N_29378,N_22910,N_18343);
nor U29379 (N_29379,N_18131,N_23625);
or U29380 (N_29380,N_19624,N_22130);
nand U29381 (N_29381,N_23528,N_19456);
nand U29382 (N_29382,N_23948,N_19521);
or U29383 (N_29383,N_21786,N_23843);
and U29384 (N_29384,N_21312,N_21347);
and U29385 (N_29385,N_20538,N_20713);
or U29386 (N_29386,N_19071,N_22406);
or U29387 (N_29387,N_20662,N_18402);
nor U29388 (N_29388,N_20050,N_18547);
and U29389 (N_29389,N_20085,N_19773);
nor U29390 (N_29390,N_20747,N_23223);
or U29391 (N_29391,N_22476,N_18962);
or U29392 (N_29392,N_19137,N_22811);
or U29393 (N_29393,N_21397,N_22745);
or U29394 (N_29394,N_19089,N_22502);
and U29395 (N_29395,N_19598,N_18306);
nor U29396 (N_29396,N_19037,N_19152);
or U29397 (N_29397,N_22401,N_21420);
xor U29398 (N_29398,N_20972,N_23560);
nand U29399 (N_29399,N_20830,N_19510);
nor U29400 (N_29400,N_20629,N_19453);
and U29401 (N_29401,N_20636,N_20828);
or U29402 (N_29402,N_22304,N_23715);
nand U29403 (N_29403,N_19994,N_19459);
and U29404 (N_29404,N_18498,N_18338);
and U29405 (N_29405,N_23984,N_18967);
nand U29406 (N_29406,N_21765,N_21397);
nor U29407 (N_29407,N_20785,N_20410);
nor U29408 (N_29408,N_21455,N_19107);
xor U29409 (N_29409,N_18993,N_23466);
and U29410 (N_29410,N_20335,N_23306);
nor U29411 (N_29411,N_21558,N_19452);
xor U29412 (N_29412,N_20384,N_23707);
and U29413 (N_29413,N_19019,N_21622);
nor U29414 (N_29414,N_20473,N_18748);
nand U29415 (N_29415,N_20136,N_21121);
nor U29416 (N_29416,N_22371,N_18795);
or U29417 (N_29417,N_22339,N_20297);
or U29418 (N_29418,N_23850,N_22087);
and U29419 (N_29419,N_20045,N_21606);
nand U29420 (N_29420,N_19927,N_23099);
or U29421 (N_29421,N_19160,N_23269);
nand U29422 (N_29422,N_20570,N_20788);
xnor U29423 (N_29423,N_19271,N_19898);
nor U29424 (N_29424,N_21113,N_23139);
xor U29425 (N_29425,N_23467,N_19009);
xnor U29426 (N_29426,N_21662,N_19711);
or U29427 (N_29427,N_23358,N_23925);
xor U29428 (N_29428,N_23058,N_22846);
nand U29429 (N_29429,N_18188,N_22896);
nand U29430 (N_29430,N_22423,N_20676);
nor U29431 (N_29431,N_18404,N_21998);
xor U29432 (N_29432,N_21417,N_21263);
xnor U29433 (N_29433,N_23586,N_18420);
xnor U29434 (N_29434,N_22874,N_23205);
and U29435 (N_29435,N_19863,N_23768);
nand U29436 (N_29436,N_23956,N_21210);
nand U29437 (N_29437,N_22900,N_20750);
nand U29438 (N_29438,N_18250,N_22025);
nor U29439 (N_29439,N_23610,N_23601);
nand U29440 (N_29440,N_19539,N_18305);
xnor U29441 (N_29441,N_23564,N_21352);
nor U29442 (N_29442,N_19184,N_19437);
or U29443 (N_29443,N_22917,N_18893);
nand U29444 (N_29444,N_22831,N_23714);
nand U29445 (N_29445,N_22888,N_20842);
nor U29446 (N_29446,N_21745,N_18867);
and U29447 (N_29447,N_22401,N_23096);
or U29448 (N_29448,N_20264,N_23525);
or U29449 (N_29449,N_22686,N_19711);
and U29450 (N_29450,N_23079,N_21091);
or U29451 (N_29451,N_18082,N_23818);
and U29452 (N_29452,N_23649,N_19599);
nand U29453 (N_29453,N_18898,N_21351);
nor U29454 (N_29454,N_22094,N_22592);
and U29455 (N_29455,N_19793,N_19999);
nand U29456 (N_29456,N_19298,N_18128);
or U29457 (N_29457,N_21911,N_19331);
xor U29458 (N_29458,N_22076,N_23064);
and U29459 (N_29459,N_23656,N_22802);
nand U29460 (N_29460,N_20066,N_23381);
nor U29461 (N_29461,N_18899,N_22883);
or U29462 (N_29462,N_23138,N_23739);
nand U29463 (N_29463,N_23066,N_22563);
nand U29464 (N_29464,N_19563,N_21573);
xor U29465 (N_29465,N_22945,N_18098);
or U29466 (N_29466,N_21697,N_20050);
nand U29467 (N_29467,N_23108,N_20290);
nand U29468 (N_29468,N_18881,N_20080);
or U29469 (N_29469,N_23956,N_23845);
nand U29470 (N_29470,N_18455,N_23430);
and U29471 (N_29471,N_23126,N_20309);
and U29472 (N_29472,N_23884,N_21650);
xnor U29473 (N_29473,N_19161,N_23817);
nor U29474 (N_29474,N_20588,N_21734);
or U29475 (N_29475,N_21021,N_21472);
xnor U29476 (N_29476,N_23806,N_22283);
and U29477 (N_29477,N_20559,N_19800);
or U29478 (N_29478,N_23491,N_20579);
xor U29479 (N_29479,N_18259,N_20327);
xor U29480 (N_29480,N_23536,N_18385);
xnor U29481 (N_29481,N_19070,N_19435);
and U29482 (N_29482,N_20177,N_22176);
nor U29483 (N_29483,N_22659,N_18315);
nor U29484 (N_29484,N_21486,N_18921);
nand U29485 (N_29485,N_19622,N_21975);
nand U29486 (N_29486,N_19420,N_23815);
nand U29487 (N_29487,N_19022,N_19260);
nand U29488 (N_29488,N_22696,N_22713);
nand U29489 (N_29489,N_22095,N_19223);
or U29490 (N_29490,N_19244,N_23119);
or U29491 (N_29491,N_20954,N_21180);
nand U29492 (N_29492,N_20750,N_18104);
and U29493 (N_29493,N_20248,N_23431);
xor U29494 (N_29494,N_22435,N_22053);
nand U29495 (N_29495,N_20171,N_19241);
and U29496 (N_29496,N_18817,N_18727);
nor U29497 (N_29497,N_18007,N_23801);
or U29498 (N_29498,N_19818,N_23143);
and U29499 (N_29499,N_22884,N_21132);
or U29500 (N_29500,N_23435,N_22900);
nor U29501 (N_29501,N_21130,N_21165);
and U29502 (N_29502,N_21369,N_18975);
or U29503 (N_29503,N_23930,N_20558);
nor U29504 (N_29504,N_22150,N_18955);
and U29505 (N_29505,N_23976,N_19902);
nor U29506 (N_29506,N_23192,N_18269);
xnor U29507 (N_29507,N_21984,N_21708);
or U29508 (N_29508,N_23937,N_21029);
nand U29509 (N_29509,N_19876,N_20239);
or U29510 (N_29510,N_22174,N_18239);
or U29511 (N_29511,N_20451,N_21632);
or U29512 (N_29512,N_19379,N_22689);
or U29513 (N_29513,N_18409,N_21953);
and U29514 (N_29514,N_21682,N_20083);
xnor U29515 (N_29515,N_22920,N_21461);
and U29516 (N_29516,N_21159,N_22208);
and U29517 (N_29517,N_20925,N_20864);
xor U29518 (N_29518,N_19233,N_20282);
xor U29519 (N_29519,N_23301,N_18354);
or U29520 (N_29520,N_20468,N_23312);
xor U29521 (N_29521,N_22714,N_19298);
nor U29522 (N_29522,N_20167,N_21622);
nand U29523 (N_29523,N_21403,N_19896);
or U29524 (N_29524,N_19252,N_20303);
nand U29525 (N_29525,N_22234,N_23793);
and U29526 (N_29526,N_20766,N_21446);
nor U29527 (N_29527,N_20737,N_19165);
and U29528 (N_29528,N_18935,N_18453);
nand U29529 (N_29529,N_22006,N_19143);
and U29530 (N_29530,N_20911,N_22239);
xor U29531 (N_29531,N_20488,N_21800);
xnor U29532 (N_29532,N_19593,N_18406);
nor U29533 (N_29533,N_20094,N_19735);
nor U29534 (N_29534,N_20636,N_23172);
or U29535 (N_29535,N_18242,N_20542);
or U29536 (N_29536,N_23235,N_22339);
nand U29537 (N_29537,N_18317,N_22523);
or U29538 (N_29538,N_23140,N_20710);
xor U29539 (N_29539,N_19301,N_18614);
xnor U29540 (N_29540,N_20497,N_19279);
or U29541 (N_29541,N_21722,N_23493);
nand U29542 (N_29542,N_22808,N_23967);
nand U29543 (N_29543,N_19274,N_19241);
nor U29544 (N_29544,N_21615,N_19587);
and U29545 (N_29545,N_18838,N_20494);
and U29546 (N_29546,N_22267,N_21556);
or U29547 (N_29547,N_20832,N_21193);
and U29548 (N_29548,N_23984,N_18088);
nor U29549 (N_29549,N_23375,N_20021);
and U29550 (N_29550,N_23075,N_22318);
and U29551 (N_29551,N_23068,N_23776);
and U29552 (N_29552,N_22696,N_18471);
and U29553 (N_29553,N_23686,N_22688);
nor U29554 (N_29554,N_18690,N_22338);
or U29555 (N_29555,N_19947,N_22300);
nor U29556 (N_29556,N_19473,N_19495);
nor U29557 (N_29557,N_19711,N_20375);
and U29558 (N_29558,N_18922,N_22370);
or U29559 (N_29559,N_23818,N_22550);
or U29560 (N_29560,N_20063,N_20881);
nor U29561 (N_29561,N_20713,N_20493);
or U29562 (N_29562,N_20026,N_19467);
nor U29563 (N_29563,N_22621,N_23714);
nand U29564 (N_29564,N_21110,N_20295);
xor U29565 (N_29565,N_19277,N_19126);
nor U29566 (N_29566,N_21163,N_19915);
or U29567 (N_29567,N_19266,N_22362);
nor U29568 (N_29568,N_21974,N_22258);
and U29569 (N_29569,N_23411,N_18059);
nand U29570 (N_29570,N_22729,N_20685);
and U29571 (N_29571,N_21755,N_20613);
xnor U29572 (N_29572,N_18943,N_19952);
nor U29573 (N_29573,N_20581,N_22057);
nor U29574 (N_29574,N_19800,N_19508);
xor U29575 (N_29575,N_18536,N_21892);
nor U29576 (N_29576,N_21834,N_20737);
or U29577 (N_29577,N_21619,N_23650);
xor U29578 (N_29578,N_21555,N_20410);
nor U29579 (N_29579,N_18671,N_18765);
or U29580 (N_29580,N_22357,N_20959);
nand U29581 (N_29581,N_18828,N_20836);
or U29582 (N_29582,N_20045,N_22108);
xnor U29583 (N_29583,N_19453,N_20034);
xor U29584 (N_29584,N_18351,N_21306);
nor U29585 (N_29585,N_21566,N_21806);
nor U29586 (N_29586,N_21007,N_19161);
and U29587 (N_29587,N_22894,N_18900);
nor U29588 (N_29588,N_20732,N_20303);
and U29589 (N_29589,N_21611,N_20548);
xor U29590 (N_29590,N_21658,N_18715);
xor U29591 (N_29591,N_21949,N_22852);
and U29592 (N_29592,N_23952,N_18324);
or U29593 (N_29593,N_23812,N_22555);
xnor U29594 (N_29594,N_19116,N_21187);
or U29595 (N_29595,N_23926,N_21538);
xnor U29596 (N_29596,N_18394,N_21641);
nand U29597 (N_29597,N_18629,N_20837);
nand U29598 (N_29598,N_20938,N_18240);
nor U29599 (N_29599,N_21398,N_19876);
nor U29600 (N_29600,N_20372,N_18174);
or U29601 (N_29601,N_19484,N_20977);
nor U29602 (N_29602,N_22915,N_23940);
nor U29603 (N_29603,N_23932,N_19847);
nand U29604 (N_29604,N_19235,N_22324);
nor U29605 (N_29605,N_19445,N_22951);
and U29606 (N_29606,N_23843,N_18268);
and U29607 (N_29607,N_20238,N_18620);
xor U29608 (N_29608,N_21499,N_21215);
nor U29609 (N_29609,N_20043,N_22973);
nand U29610 (N_29610,N_18189,N_18397);
xor U29611 (N_29611,N_22259,N_21503);
nand U29612 (N_29612,N_21129,N_21032);
or U29613 (N_29613,N_20051,N_22031);
and U29614 (N_29614,N_18193,N_20037);
or U29615 (N_29615,N_22692,N_20844);
and U29616 (N_29616,N_20906,N_20970);
or U29617 (N_29617,N_21656,N_21346);
nor U29618 (N_29618,N_22401,N_23342);
nor U29619 (N_29619,N_19110,N_20491);
or U29620 (N_29620,N_20645,N_19883);
and U29621 (N_29621,N_18908,N_22844);
nand U29622 (N_29622,N_19528,N_19860);
and U29623 (N_29623,N_19838,N_23971);
or U29624 (N_29624,N_22287,N_23332);
nor U29625 (N_29625,N_23617,N_21013);
nor U29626 (N_29626,N_21232,N_23526);
nor U29627 (N_29627,N_21674,N_18766);
nor U29628 (N_29628,N_20696,N_21250);
nand U29629 (N_29629,N_18238,N_19752);
nand U29630 (N_29630,N_18841,N_18326);
xor U29631 (N_29631,N_22648,N_21542);
or U29632 (N_29632,N_18481,N_22975);
and U29633 (N_29633,N_22356,N_19141);
or U29634 (N_29634,N_20774,N_23075);
and U29635 (N_29635,N_22695,N_22582);
and U29636 (N_29636,N_22051,N_22025);
nor U29637 (N_29637,N_20603,N_18575);
and U29638 (N_29638,N_22622,N_21549);
nor U29639 (N_29639,N_19016,N_22240);
and U29640 (N_29640,N_18147,N_19468);
xnor U29641 (N_29641,N_23981,N_22263);
and U29642 (N_29642,N_19602,N_22434);
and U29643 (N_29643,N_21358,N_23630);
nand U29644 (N_29644,N_23210,N_23239);
xnor U29645 (N_29645,N_21739,N_20564);
nor U29646 (N_29646,N_21814,N_23114);
xor U29647 (N_29647,N_18218,N_21703);
nor U29648 (N_29648,N_21481,N_22975);
nor U29649 (N_29649,N_21488,N_23527);
nor U29650 (N_29650,N_22998,N_22458);
and U29651 (N_29651,N_22856,N_20690);
or U29652 (N_29652,N_19860,N_20046);
nor U29653 (N_29653,N_21708,N_19277);
nor U29654 (N_29654,N_19082,N_23061);
nand U29655 (N_29655,N_18338,N_22479);
or U29656 (N_29656,N_22540,N_21958);
and U29657 (N_29657,N_20263,N_20700);
xor U29658 (N_29658,N_23141,N_23563);
xnor U29659 (N_29659,N_21861,N_22468);
or U29660 (N_29660,N_21705,N_22919);
and U29661 (N_29661,N_23741,N_23895);
nor U29662 (N_29662,N_21747,N_19930);
nor U29663 (N_29663,N_21353,N_19427);
nor U29664 (N_29664,N_20120,N_21954);
and U29665 (N_29665,N_21593,N_22204);
or U29666 (N_29666,N_21411,N_20485);
and U29667 (N_29667,N_20834,N_21407);
or U29668 (N_29668,N_19610,N_21832);
xor U29669 (N_29669,N_22101,N_22988);
nor U29670 (N_29670,N_22865,N_18150);
nor U29671 (N_29671,N_23188,N_23095);
or U29672 (N_29672,N_22789,N_21583);
nand U29673 (N_29673,N_23575,N_21879);
nand U29674 (N_29674,N_22496,N_19367);
xor U29675 (N_29675,N_21104,N_19394);
or U29676 (N_29676,N_19330,N_22266);
xnor U29677 (N_29677,N_18456,N_23921);
nand U29678 (N_29678,N_19051,N_21838);
nand U29679 (N_29679,N_22372,N_21880);
and U29680 (N_29680,N_21882,N_19399);
nor U29681 (N_29681,N_22087,N_21706);
nand U29682 (N_29682,N_20225,N_22894);
and U29683 (N_29683,N_18158,N_21430);
nor U29684 (N_29684,N_22501,N_21238);
xnor U29685 (N_29685,N_18963,N_22950);
nand U29686 (N_29686,N_20178,N_21617);
nand U29687 (N_29687,N_18281,N_19644);
nand U29688 (N_29688,N_19497,N_22969);
nand U29689 (N_29689,N_22810,N_20819);
nand U29690 (N_29690,N_22709,N_21870);
nor U29691 (N_29691,N_18534,N_20526);
xnor U29692 (N_29692,N_23823,N_20487);
xnor U29693 (N_29693,N_20077,N_21554);
or U29694 (N_29694,N_19117,N_22713);
nand U29695 (N_29695,N_21079,N_23943);
or U29696 (N_29696,N_22283,N_21241);
nand U29697 (N_29697,N_23302,N_20289);
and U29698 (N_29698,N_23741,N_23646);
nand U29699 (N_29699,N_22435,N_19299);
xnor U29700 (N_29700,N_19086,N_18089);
xor U29701 (N_29701,N_22042,N_23652);
or U29702 (N_29702,N_21957,N_19813);
nor U29703 (N_29703,N_22352,N_21124);
or U29704 (N_29704,N_18976,N_23710);
nand U29705 (N_29705,N_22537,N_21642);
and U29706 (N_29706,N_19948,N_21719);
xnor U29707 (N_29707,N_23502,N_21986);
or U29708 (N_29708,N_21475,N_21535);
nand U29709 (N_29709,N_20206,N_19586);
or U29710 (N_29710,N_19101,N_18348);
and U29711 (N_29711,N_20752,N_20112);
nand U29712 (N_29712,N_21443,N_21679);
and U29713 (N_29713,N_19861,N_21381);
xnor U29714 (N_29714,N_22027,N_21957);
nor U29715 (N_29715,N_20445,N_22451);
or U29716 (N_29716,N_22523,N_21911);
nor U29717 (N_29717,N_18813,N_21474);
xnor U29718 (N_29718,N_22378,N_19553);
or U29719 (N_29719,N_19209,N_22375);
xnor U29720 (N_29720,N_19093,N_20243);
and U29721 (N_29721,N_21546,N_22142);
and U29722 (N_29722,N_23485,N_22114);
nor U29723 (N_29723,N_23544,N_23104);
or U29724 (N_29724,N_23491,N_20566);
xor U29725 (N_29725,N_22191,N_20095);
xnor U29726 (N_29726,N_18936,N_21478);
and U29727 (N_29727,N_22465,N_21425);
or U29728 (N_29728,N_19778,N_19687);
nor U29729 (N_29729,N_21409,N_20440);
xnor U29730 (N_29730,N_18545,N_22864);
nor U29731 (N_29731,N_20156,N_18967);
and U29732 (N_29732,N_20351,N_19402);
and U29733 (N_29733,N_23333,N_20461);
nor U29734 (N_29734,N_20246,N_19990);
and U29735 (N_29735,N_21757,N_23404);
or U29736 (N_29736,N_20263,N_19155);
and U29737 (N_29737,N_20197,N_19796);
nor U29738 (N_29738,N_21371,N_18345);
and U29739 (N_29739,N_20619,N_23837);
xor U29740 (N_29740,N_18913,N_23037);
or U29741 (N_29741,N_18468,N_22842);
or U29742 (N_29742,N_20446,N_21272);
nor U29743 (N_29743,N_18150,N_18369);
and U29744 (N_29744,N_20226,N_21082);
xor U29745 (N_29745,N_21540,N_23453);
nand U29746 (N_29746,N_23169,N_21575);
xor U29747 (N_29747,N_19783,N_18730);
nand U29748 (N_29748,N_21060,N_20731);
xor U29749 (N_29749,N_23680,N_21045);
nand U29750 (N_29750,N_18211,N_22181);
nor U29751 (N_29751,N_20106,N_20954);
nor U29752 (N_29752,N_19821,N_20144);
or U29753 (N_29753,N_23171,N_20705);
xor U29754 (N_29754,N_22859,N_20823);
xnor U29755 (N_29755,N_23354,N_18934);
nand U29756 (N_29756,N_19453,N_20241);
or U29757 (N_29757,N_19033,N_21682);
xnor U29758 (N_29758,N_18945,N_21192);
or U29759 (N_29759,N_19996,N_19616);
or U29760 (N_29760,N_19735,N_21776);
and U29761 (N_29761,N_18943,N_18697);
nand U29762 (N_29762,N_20625,N_18961);
and U29763 (N_29763,N_21730,N_22571);
nand U29764 (N_29764,N_22344,N_21651);
xor U29765 (N_29765,N_18401,N_19193);
and U29766 (N_29766,N_22905,N_20960);
xor U29767 (N_29767,N_22567,N_19371);
nand U29768 (N_29768,N_19471,N_21991);
and U29769 (N_29769,N_23010,N_23628);
nor U29770 (N_29770,N_22688,N_23575);
nor U29771 (N_29771,N_22921,N_21715);
or U29772 (N_29772,N_20516,N_19339);
and U29773 (N_29773,N_20384,N_22399);
xor U29774 (N_29774,N_19531,N_23191);
and U29775 (N_29775,N_20588,N_21479);
nor U29776 (N_29776,N_23775,N_22272);
nand U29777 (N_29777,N_19464,N_22370);
and U29778 (N_29778,N_23725,N_23974);
or U29779 (N_29779,N_18357,N_23361);
xor U29780 (N_29780,N_20193,N_23350);
nand U29781 (N_29781,N_23735,N_20741);
or U29782 (N_29782,N_21497,N_20529);
xnor U29783 (N_29783,N_23443,N_18569);
or U29784 (N_29784,N_23686,N_20043);
or U29785 (N_29785,N_22588,N_18054);
and U29786 (N_29786,N_18046,N_22747);
and U29787 (N_29787,N_21236,N_21650);
and U29788 (N_29788,N_18314,N_23449);
nor U29789 (N_29789,N_20779,N_20451);
nand U29790 (N_29790,N_18269,N_20613);
nand U29791 (N_29791,N_23432,N_20891);
xor U29792 (N_29792,N_23638,N_21122);
nor U29793 (N_29793,N_23344,N_21009);
nor U29794 (N_29794,N_18125,N_21075);
or U29795 (N_29795,N_21165,N_20787);
nor U29796 (N_29796,N_18765,N_18114);
nand U29797 (N_29797,N_20414,N_22481);
or U29798 (N_29798,N_20746,N_18140);
nand U29799 (N_29799,N_19707,N_22417);
nor U29800 (N_29800,N_22262,N_22703);
xor U29801 (N_29801,N_23130,N_22388);
or U29802 (N_29802,N_19750,N_21200);
nor U29803 (N_29803,N_20976,N_22205);
and U29804 (N_29804,N_19638,N_21006);
and U29805 (N_29805,N_22007,N_22770);
nor U29806 (N_29806,N_20145,N_19951);
nand U29807 (N_29807,N_19516,N_19382);
nor U29808 (N_29808,N_22054,N_19629);
nor U29809 (N_29809,N_18342,N_20877);
nand U29810 (N_29810,N_19284,N_19563);
xor U29811 (N_29811,N_22241,N_21003);
nand U29812 (N_29812,N_21658,N_23905);
nor U29813 (N_29813,N_20915,N_19548);
and U29814 (N_29814,N_19815,N_21707);
or U29815 (N_29815,N_23714,N_18958);
or U29816 (N_29816,N_19432,N_19788);
and U29817 (N_29817,N_22206,N_23494);
nand U29818 (N_29818,N_20010,N_18236);
xnor U29819 (N_29819,N_23315,N_18380);
nor U29820 (N_29820,N_21906,N_18468);
and U29821 (N_29821,N_23872,N_19277);
xnor U29822 (N_29822,N_22524,N_18347);
nand U29823 (N_29823,N_20368,N_21356);
and U29824 (N_29824,N_23854,N_21426);
or U29825 (N_29825,N_21083,N_21585);
and U29826 (N_29826,N_23432,N_22381);
xnor U29827 (N_29827,N_21950,N_23657);
nand U29828 (N_29828,N_21008,N_19246);
or U29829 (N_29829,N_18977,N_22624);
nor U29830 (N_29830,N_19693,N_21466);
xnor U29831 (N_29831,N_21984,N_18491);
or U29832 (N_29832,N_18996,N_22979);
nor U29833 (N_29833,N_22534,N_18848);
and U29834 (N_29834,N_19187,N_18979);
nand U29835 (N_29835,N_19249,N_19324);
or U29836 (N_29836,N_19948,N_21581);
nand U29837 (N_29837,N_21859,N_21246);
and U29838 (N_29838,N_22155,N_18699);
nand U29839 (N_29839,N_22839,N_23745);
and U29840 (N_29840,N_18375,N_21088);
or U29841 (N_29841,N_18137,N_20989);
nand U29842 (N_29842,N_21670,N_22748);
and U29843 (N_29843,N_18873,N_19606);
nor U29844 (N_29844,N_20939,N_22502);
xnor U29845 (N_29845,N_20641,N_23138);
nor U29846 (N_29846,N_22880,N_21311);
nor U29847 (N_29847,N_18105,N_18012);
and U29848 (N_29848,N_21431,N_19720);
nand U29849 (N_29849,N_18326,N_23188);
or U29850 (N_29850,N_21464,N_23903);
nand U29851 (N_29851,N_21692,N_21394);
or U29852 (N_29852,N_23689,N_23416);
or U29853 (N_29853,N_21014,N_20006);
nand U29854 (N_29854,N_19576,N_21929);
or U29855 (N_29855,N_18654,N_23189);
nor U29856 (N_29856,N_20998,N_20124);
and U29857 (N_29857,N_21187,N_19034);
or U29858 (N_29858,N_22911,N_19581);
and U29859 (N_29859,N_18876,N_21238);
nor U29860 (N_29860,N_21666,N_19872);
nor U29861 (N_29861,N_20212,N_20726);
xnor U29862 (N_29862,N_20178,N_21677);
or U29863 (N_29863,N_18016,N_22897);
xnor U29864 (N_29864,N_18847,N_22761);
nor U29865 (N_29865,N_20842,N_20908);
or U29866 (N_29866,N_23612,N_19286);
nor U29867 (N_29867,N_22655,N_18180);
xnor U29868 (N_29868,N_23547,N_19808);
and U29869 (N_29869,N_23074,N_18135);
nand U29870 (N_29870,N_22178,N_22206);
or U29871 (N_29871,N_21948,N_20424);
xor U29872 (N_29872,N_18016,N_19479);
and U29873 (N_29873,N_22701,N_21937);
nand U29874 (N_29874,N_22483,N_22415);
xor U29875 (N_29875,N_21560,N_20696);
and U29876 (N_29876,N_23655,N_21811);
xnor U29877 (N_29877,N_22221,N_23807);
or U29878 (N_29878,N_19232,N_22114);
or U29879 (N_29879,N_21352,N_18595);
nor U29880 (N_29880,N_21352,N_18043);
or U29881 (N_29881,N_21005,N_20910);
xor U29882 (N_29882,N_19216,N_19179);
and U29883 (N_29883,N_23587,N_19484);
and U29884 (N_29884,N_19922,N_21020);
nand U29885 (N_29885,N_18268,N_19008);
or U29886 (N_29886,N_20566,N_20055);
nand U29887 (N_29887,N_19066,N_20248);
nand U29888 (N_29888,N_21698,N_19120);
or U29889 (N_29889,N_19131,N_23343);
nand U29890 (N_29890,N_23727,N_21116);
and U29891 (N_29891,N_18965,N_18155);
xor U29892 (N_29892,N_19041,N_19251);
nor U29893 (N_29893,N_19315,N_20187);
or U29894 (N_29894,N_22154,N_23993);
and U29895 (N_29895,N_21395,N_21936);
nor U29896 (N_29896,N_21123,N_19385);
and U29897 (N_29897,N_23984,N_19641);
nor U29898 (N_29898,N_19437,N_19889);
nand U29899 (N_29899,N_22183,N_22963);
or U29900 (N_29900,N_19737,N_19875);
xor U29901 (N_29901,N_22756,N_18594);
or U29902 (N_29902,N_22469,N_22021);
nor U29903 (N_29903,N_20852,N_22289);
nor U29904 (N_29904,N_21369,N_20462);
nand U29905 (N_29905,N_22822,N_23058);
nand U29906 (N_29906,N_18444,N_23218);
and U29907 (N_29907,N_23607,N_22964);
xnor U29908 (N_29908,N_23395,N_21927);
nand U29909 (N_29909,N_18758,N_20971);
or U29910 (N_29910,N_21248,N_21417);
nor U29911 (N_29911,N_19358,N_23025);
or U29912 (N_29912,N_20944,N_22955);
or U29913 (N_29913,N_22339,N_21885);
and U29914 (N_29914,N_21093,N_18502);
nor U29915 (N_29915,N_20966,N_23357);
xnor U29916 (N_29916,N_21757,N_23542);
xnor U29917 (N_29917,N_18069,N_18163);
xor U29918 (N_29918,N_21448,N_23208);
or U29919 (N_29919,N_23667,N_23883);
and U29920 (N_29920,N_21273,N_21010);
nor U29921 (N_29921,N_22833,N_18153);
or U29922 (N_29922,N_19901,N_20911);
nand U29923 (N_29923,N_21284,N_22225);
or U29924 (N_29924,N_22869,N_18264);
and U29925 (N_29925,N_18449,N_23308);
nand U29926 (N_29926,N_23533,N_18527);
nand U29927 (N_29927,N_18011,N_19179);
and U29928 (N_29928,N_21537,N_19672);
nor U29929 (N_29929,N_18444,N_19823);
nor U29930 (N_29930,N_22468,N_22003);
nor U29931 (N_29931,N_19085,N_19563);
nor U29932 (N_29932,N_21085,N_18489);
nand U29933 (N_29933,N_21683,N_18043);
xnor U29934 (N_29934,N_20279,N_21461);
or U29935 (N_29935,N_19547,N_22646);
nor U29936 (N_29936,N_20409,N_21713);
or U29937 (N_29937,N_21565,N_18817);
or U29938 (N_29938,N_20494,N_19646);
nand U29939 (N_29939,N_22596,N_19427);
and U29940 (N_29940,N_23245,N_21830);
and U29941 (N_29941,N_23934,N_23772);
and U29942 (N_29942,N_22232,N_22791);
and U29943 (N_29943,N_22703,N_18761);
and U29944 (N_29944,N_21061,N_19752);
or U29945 (N_29945,N_21929,N_21093);
nand U29946 (N_29946,N_19343,N_22047);
or U29947 (N_29947,N_22508,N_19657);
and U29948 (N_29948,N_19172,N_18679);
nor U29949 (N_29949,N_19679,N_22251);
or U29950 (N_29950,N_23912,N_20284);
nor U29951 (N_29951,N_19556,N_20591);
and U29952 (N_29952,N_23578,N_20063);
nand U29953 (N_29953,N_20971,N_19113);
or U29954 (N_29954,N_23290,N_20688);
nand U29955 (N_29955,N_22999,N_23539);
nor U29956 (N_29956,N_21508,N_18219);
and U29957 (N_29957,N_20012,N_21848);
nor U29958 (N_29958,N_20537,N_22735);
nor U29959 (N_29959,N_23756,N_21830);
nor U29960 (N_29960,N_20450,N_19710);
or U29961 (N_29961,N_19832,N_19160);
or U29962 (N_29962,N_23320,N_19741);
and U29963 (N_29963,N_23864,N_22256);
or U29964 (N_29964,N_20343,N_22392);
nand U29965 (N_29965,N_20692,N_21347);
nand U29966 (N_29966,N_19014,N_19669);
or U29967 (N_29967,N_22193,N_20254);
or U29968 (N_29968,N_19494,N_21408);
xor U29969 (N_29969,N_22328,N_23471);
xnor U29970 (N_29970,N_21966,N_20440);
and U29971 (N_29971,N_22270,N_18989);
and U29972 (N_29972,N_21500,N_21869);
nand U29973 (N_29973,N_19874,N_22142);
xor U29974 (N_29974,N_21807,N_21092);
nor U29975 (N_29975,N_18198,N_19273);
or U29976 (N_29976,N_18021,N_21727);
nor U29977 (N_29977,N_23178,N_22931);
or U29978 (N_29978,N_18826,N_21942);
nor U29979 (N_29979,N_20094,N_22496);
nand U29980 (N_29980,N_23789,N_19395);
xor U29981 (N_29981,N_20331,N_22049);
and U29982 (N_29982,N_20015,N_21531);
or U29983 (N_29983,N_20132,N_22847);
nor U29984 (N_29984,N_22657,N_23413);
xor U29985 (N_29985,N_22273,N_22439);
nand U29986 (N_29986,N_21793,N_20119);
or U29987 (N_29987,N_21250,N_19724);
xor U29988 (N_29988,N_19050,N_19092);
xor U29989 (N_29989,N_20331,N_19663);
or U29990 (N_29990,N_23372,N_23599);
nor U29991 (N_29991,N_19677,N_23863);
or U29992 (N_29992,N_19667,N_20116);
or U29993 (N_29993,N_23919,N_19297);
and U29994 (N_29994,N_18453,N_23746);
nand U29995 (N_29995,N_21630,N_20226);
xnor U29996 (N_29996,N_19389,N_23642);
xor U29997 (N_29997,N_19765,N_18723);
and U29998 (N_29998,N_23829,N_19452);
xor U29999 (N_29999,N_19201,N_20108);
or UO_0 (O_0,N_25167,N_26947);
xnor UO_1 (O_1,N_26641,N_27483);
nand UO_2 (O_2,N_25672,N_25484);
or UO_3 (O_3,N_26527,N_29554);
nor UO_4 (O_4,N_27955,N_25849);
nand UO_5 (O_5,N_28041,N_29871);
xor UO_6 (O_6,N_28834,N_24573);
or UO_7 (O_7,N_28868,N_28142);
xor UO_8 (O_8,N_28362,N_25041);
nor UO_9 (O_9,N_25286,N_29791);
or UO_10 (O_10,N_27951,N_29570);
nor UO_11 (O_11,N_24539,N_26737);
nand UO_12 (O_12,N_24789,N_26176);
xnor UO_13 (O_13,N_25401,N_25520);
and UO_14 (O_14,N_24688,N_27715);
or UO_15 (O_15,N_24517,N_29120);
xnor UO_16 (O_16,N_25026,N_25179);
xnor UO_17 (O_17,N_28522,N_24015);
and UO_18 (O_18,N_29395,N_26608);
xnor UO_19 (O_19,N_29321,N_26366);
and UO_20 (O_20,N_28226,N_24715);
or UO_21 (O_21,N_27708,N_28819);
or UO_22 (O_22,N_26490,N_28640);
or UO_23 (O_23,N_25854,N_28582);
and UO_24 (O_24,N_24048,N_25066);
nand UO_25 (O_25,N_25755,N_29641);
nor UO_26 (O_26,N_28778,N_25614);
nand UO_27 (O_27,N_28480,N_26107);
nand UO_28 (O_28,N_27645,N_26790);
xor UO_29 (O_29,N_28239,N_24492);
nor UO_30 (O_30,N_26014,N_27423);
and UO_31 (O_31,N_29543,N_25525);
or UO_32 (O_32,N_27647,N_27936);
or UO_33 (O_33,N_26864,N_28175);
nand UO_34 (O_34,N_27772,N_29031);
nor UO_35 (O_35,N_28323,N_29854);
xor UO_36 (O_36,N_28675,N_24974);
or UO_37 (O_37,N_24075,N_26673);
or UO_38 (O_38,N_26343,N_24775);
or UO_39 (O_39,N_27519,N_29184);
xnor UO_40 (O_40,N_26997,N_27249);
nor UO_41 (O_41,N_26536,N_26516);
nor UO_42 (O_42,N_25339,N_26636);
nand UO_43 (O_43,N_29469,N_28987);
and UO_44 (O_44,N_27864,N_26349);
nand UO_45 (O_45,N_28287,N_26091);
nor UO_46 (O_46,N_27334,N_29172);
and UO_47 (O_47,N_27059,N_25120);
xnor UO_48 (O_48,N_28598,N_27041);
and UO_49 (O_49,N_28276,N_26786);
nor UO_50 (O_50,N_28790,N_24147);
nand UO_51 (O_51,N_26991,N_27841);
and UO_52 (O_52,N_29107,N_26310);
and UO_53 (O_53,N_26239,N_29348);
xnor UO_54 (O_54,N_28900,N_29899);
nor UO_55 (O_55,N_24818,N_26478);
or UO_56 (O_56,N_24244,N_28935);
and UO_57 (O_57,N_24289,N_28406);
xor UO_58 (O_58,N_26395,N_25280);
or UO_59 (O_59,N_25661,N_26746);
nand UO_60 (O_60,N_27252,N_26347);
xor UO_61 (O_61,N_26162,N_26062);
and UO_62 (O_62,N_27893,N_29676);
or UO_63 (O_63,N_25669,N_25512);
xnor UO_64 (O_64,N_29287,N_26160);
nor UO_65 (O_65,N_24078,N_24521);
nor UO_66 (O_66,N_26015,N_29093);
xor UO_67 (O_67,N_25343,N_27798);
nor UO_68 (O_68,N_24997,N_24723);
nor UO_69 (O_69,N_24845,N_25338);
or UO_70 (O_70,N_24023,N_29531);
xnor UO_71 (O_71,N_27711,N_24493);
and UO_72 (O_72,N_27834,N_25933);
xnor UO_73 (O_73,N_25981,N_27712);
nor UO_74 (O_74,N_27793,N_27648);
and UO_75 (O_75,N_28456,N_26992);
xnor UO_76 (O_76,N_28973,N_25535);
or UO_77 (O_77,N_27944,N_29041);
nand UO_78 (O_78,N_27346,N_24941);
and UO_79 (O_79,N_26892,N_27828);
nand UO_80 (O_80,N_29516,N_29908);
and UO_81 (O_81,N_25402,N_28433);
nor UO_82 (O_82,N_29923,N_24219);
or UO_83 (O_83,N_29955,N_26494);
nand UO_84 (O_84,N_25270,N_29198);
and UO_85 (O_85,N_24594,N_28812);
and UO_86 (O_86,N_29176,N_27923);
nand UO_87 (O_87,N_27010,N_27759);
xnor UO_88 (O_88,N_27921,N_28628);
or UO_89 (O_89,N_27734,N_29070);
or UO_90 (O_90,N_24519,N_25962);
and UO_91 (O_91,N_26030,N_28391);
nor UO_92 (O_92,N_24740,N_25992);
or UO_93 (O_93,N_26482,N_25435);
nor UO_94 (O_94,N_25150,N_26426);
or UO_95 (O_95,N_26534,N_24704);
or UO_96 (O_96,N_24861,N_26671);
or UO_97 (O_97,N_24165,N_27452);
nor UO_98 (O_98,N_28886,N_27998);
xnor UO_99 (O_99,N_27342,N_28477);
and UO_100 (O_100,N_25096,N_25998);
nand UO_101 (O_101,N_25900,N_28903);
xor UO_102 (O_102,N_25376,N_29616);
xor UO_103 (O_103,N_29998,N_24033);
xnor UO_104 (O_104,N_27007,N_24378);
xnor UO_105 (O_105,N_28629,N_24647);
or UO_106 (O_106,N_24524,N_26092);
nor UO_107 (O_107,N_27593,N_25634);
nor UO_108 (O_108,N_26268,N_25508);
nand UO_109 (O_109,N_27453,N_25194);
or UO_110 (O_110,N_24070,N_28368);
xor UO_111 (O_111,N_26204,N_24153);
nand UO_112 (O_112,N_27698,N_26948);
and UO_113 (O_113,N_25304,N_25380);
xor UO_114 (O_114,N_24605,N_28849);
xor UO_115 (O_115,N_24295,N_29745);
or UO_116 (O_116,N_26812,N_24267);
or UO_117 (O_117,N_26101,N_29402);
nand UO_118 (O_118,N_26587,N_27705);
nand UO_119 (O_119,N_27961,N_26566);
nand UO_120 (O_120,N_28594,N_29628);
nand UO_121 (O_121,N_28850,N_28082);
nor UO_122 (O_122,N_29410,N_29349);
xnor UO_123 (O_123,N_27178,N_26927);
or UO_124 (O_124,N_25146,N_27092);
xor UO_125 (O_125,N_29234,N_29891);
nor UO_126 (O_126,N_25616,N_24472);
or UO_127 (O_127,N_25209,N_24619);
nand UO_128 (O_128,N_29413,N_25511);
and UO_129 (O_129,N_25526,N_26080);
nor UO_130 (O_130,N_25187,N_24104);
and UO_131 (O_131,N_26362,N_27722);
and UO_132 (O_132,N_26049,N_29480);
nor UO_133 (O_133,N_25815,N_26582);
xor UO_134 (O_134,N_24156,N_29209);
or UO_135 (O_135,N_29930,N_27157);
xnor UO_136 (O_136,N_27596,N_28359);
or UO_137 (O_137,N_25673,N_28417);
or UO_138 (O_138,N_29390,N_29577);
nand UO_139 (O_139,N_25638,N_26010);
and UO_140 (O_140,N_25922,N_28939);
nand UO_141 (O_141,N_29169,N_29449);
xor UO_142 (O_142,N_29486,N_25784);
nand UO_143 (O_143,N_27384,N_27467);
and UO_144 (O_144,N_28783,N_25206);
nand UO_145 (O_145,N_26396,N_25622);
nand UO_146 (O_146,N_25252,N_24520);
nand UO_147 (O_147,N_24136,N_24178);
or UO_148 (O_148,N_24606,N_26957);
nand UO_149 (O_149,N_26398,N_27605);
nor UO_150 (O_150,N_26038,N_29769);
and UO_151 (O_151,N_27977,N_28038);
and UO_152 (O_152,N_28355,N_24393);
and UO_153 (O_153,N_27589,N_25300);
nor UO_154 (O_154,N_25572,N_25603);
nand UO_155 (O_155,N_24037,N_25950);
and UO_156 (O_156,N_24877,N_28552);
nand UO_157 (O_157,N_27883,N_26949);
or UO_158 (O_158,N_24461,N_27969);
or UO_159 (O_159,N_25073,N_27775);
or UO_160 (O_160,N_28086,N_27665);
nor UO_161 (O_161,N_28986,N_25919);
or UO_162 (O_162,N_28632,N_27463);
nand UO_163 (O_163,N_28774,N_29478);
and UO_164 (O_164,N_25116,N_24194);
or UO_165 (O_165,N_24551,N_27690);
nand UO_166 (O_166,N_28025,N_26959);
or UO_167 (O_167,N_28578,N_28780);
nand UO_168 (O_168,N_24210,N_26755);
nor UO_169 (O_169,N_27782,N_26810);
and UO_170 (O_170,N_25968,N_26690);
and UO_171 (O_171,N_24898,N_24570);
nor UO_172 (O_172,N_29537,N_24678);
and UO_173 (O_173,N_25879,N_26900);
and UO_174 (O_174,N_29695,N_24248);
nand UO_175 (O_175,N_26238,N_27513);
and UO_176 (O_176,N_29091,N_24249);
nand UO_177 (O_177,N_26215,N_25394);
and UO_178 (O_178,N_25009,N_24060);
nand UO_179 (O_179,N_25643,N_27225);
nand UO_180 (O_180,N_25524,N_29709);
or UO_181 (O_181,N_28198,N_24724);
nand UO_182 (O_182,N_25698,N_29645);
nand UO_183 (O_183,N_24263,N_26389);
or UO_184 (O_184,N_27383,N_24375);
and UO_185 (O_185,N_24039,N_27022);
nand UO_186 (O_186,N_24176,N_29126);
and UO_187 (O_187,N_25322,N_26245);
nand UO_188 (O_188,N_24428,N_25607);
or UO_189 (O_189,N_24245,N_27580);
xor UO_190 (O_190,N_28408,N_29821);
and UO_191 (O_191,N_24301,N_28777);
nor UO_192 (O_192,N_24691,N_25001);
nand UO_193 (O_193,N_27680,N_24951);
nor UO_194 (O_194,N_28394,N_26454);
nor UO_195 (O_195,N_27840,N_27332);
xor UO_196 (O_196,N_27014,N_28474);
and UO_197 (O_197,N_29197,N_27694);
nor UO_198 (O_198,N_25248,N_26439);
or UO_199 (O_199,N_28074,N_24872);
nand UO_200 (O_200,N_27094,N_24402);
nand UO_201 (O_201,N_24126,N_29991);
and UO_202 (O_202,N_24484,N_28670);
and UO_203 (O_203,N_24068,N_29263);
nand UO_204 (O_204,N_26056,N_28566);
and UO_205 (O_205,N_27867,N_25264);
nor UO_206 (O_206,N_27473,N_28214);
nor UO_207 (O_207,N_28450,N_25540);
or UO_208 (O_208,N_28716,N_28428);
nor UO_209 (O_209,N_26921,N_24534);
nor UO_210 (O_210,N_28584,N_29672);
xor UO_211 (O_211,N_27741,N_25753);
xor UO_212 (O_212,N_28424,N_26477);
nor UO_213 (O_213,N_29522,N_27839);
nor UO_214 (O_214,N_26971,N_28662);
nand UO_215 (O_215,N_24038,N_28472);
or UO_216 (O_216,N_29850,N_25365);
and UO_217 (O_217,N_26441,N_25792);
nor UO_218 (O_218,N_29778,N_27151);
nor UO_219 (O_219,N_25573,N_26094);
nand UO_220 (O_220,N_25040,N_27899);
xnor UO_221 (O_221,N_25650,N_25044);
and UO_222 (O_222,N_27458,N_26951);
nor UO_223 (O_223,N_24591,N_28139);
nor UO_224 (O_224,N_24299,N_29274);
nand UO_225 (O_225,N_28397,N_26473);
and UO_226 (O_226,N_25710,N_25692);
and UO_227 (O_227,N_24003,N_28998);
and UO_228 (O_228,N_28343,N_27750);
nor UO_229 (O_229,N_29648,N_26313);
xor UO_230 (O_230,N_28878,N_25825);
or UO_231 (O_231,N_25993,N_26603);
or UO_232 (O_232,N_25881,N_28170);
or UO_233 (O_233,N_27307,N_26065);
nand UO_234 (O_234,N_25314,N_25481);
xnor UO_235 (O_235,N_27379,N_25766);
xor UO_236 (O_236,N_29838,N_24433);
xor UO_237 (O_237,N_29824,N_27790);
nand UO_238 (O_238,N_27214,N_29611);
nand UO_239 (O_239,N_27636,N_27613);
and UO_240 (O_240,N_27510,N_27975);
xnor UO_241 (O_241,N_25004,N_24749);
nand UO_242 (O_242,N_29314,N_24696);
or UO_243 (O_243,N_24705,N_25822);
or UO_244 (O_244,N_26303,N_29690);
or UO_245 (O_245,N_28311,N_26639);
nand UO_246 (O_246,N_27373,N_27603);
and UO_247 (O_247,N_28246,N_28217);
nand UO_248 (O_248,N_25081,N_29897);
xor UO_249 (O_249,N_27988,N_29830);
xnor UO_250 (O_250,N_27305,N_25449);
nand UO_251 (O_251,N_29889,N_27770);
or UO_252 (O_252,N_24702,N_25362);
xnor UO_253 (O_253,N_29067,N_27742);
or UO_254 (O_254,N_29843,N_27766);
nand UO_255 (O_255,N_24954,N_27093);
nand UO_256 (O_256,N_25901,N_28898);
or UO_257 (O_257,N_27582,N_27492);
and UO_258 (O_258,N_28667,N_25970);
xor UO_259 (O_259,N_24306,N_27304);
or UO_260 (O_260,N_26644,N_28680);
nor UO_261 (O_261,N_27845,N_29608);
nor UO_262 (O_262,N_29175,N_28729);
nor UO_263 (O_263,N_25729,N_27223);
nor UO_264 (O_264,N_27555,N_25364);
or UO_265 (O_265,N_25451,N_24292);
nor UO_266 (O_266,N_28719,N_24827);
nor UO_267 (O_267,N_25445,N_25611);
or UO_268 (O_268,N_29189,N_27043);
or UO_269 (O_269,N_24857,N_26481);
nor UO_270 (O_270,N_24773,N_27161);
xnor UO_271 (O_271,N_27488,N_24737);
xnor UO_272 (O_272,N_29751,N_26497);
nand UO_273 (O_273,N_27166,N_24367);
or UO_274 (O_274,N_27894,N_24149);
nand UO_275 (O_275,N_29905,N_24985);
nand UO_276 (O_276,N_29494,N_29153);
xor UO_277 (O_277,N_29151,N_29202);
or UO_278 (O_278,N_24457,N_25291);
xor UO_279 (O_279,N_24173,N_27737);
nor UO_280 (O_280,N_26938,N_27856);
nand UO_281 (O_281,N_25728,N_29810);
xnor UO_282 (O_282,N_25757,N_26631);
or UO_283 (O_283,N_26844,N_28854);
and UO_284 (O_284,N_27032,N_24382);
and UO_285 (O_285,N_24386,N_26550);
and UO_286 (O_286,N_26336,N_24533);
and UO_287 (O_287,N_27788,N_29619);
and UO_288 (O_288,N_28661,N_28194);
nand UO_289 (O_289,N_27604,N_26901);
xnor UO_290 (O_290,N_29772,N_25235);
xor UO_291 (O_291,N_27374,N_27701);
and UO_292 (O_292,N_24734,N_27105);
nor UO_293 (O_293,N_27993,N_26674);
nand UO_294 (O_294,N_26664,N_27460);
or UO_295 (O_295,N_28208,N_26384);
nor UO_296 (O_296,N_29039,N_26431);
or UO_297 (O_297,N_25140,N_24069);
and UO_298 (O_298,N_26139,N_28965);
nor UO_299 (O_299,N_26841,N_28943);
nand UO_300 (O_300,N_28934,N_25907);
nand UO_301 (O_301,N_24733,N_25318);
nand UO_302 (O_302,N_28296,N_27208);
and UO_303 (O_303,N_25884,N_28023);
or UO_304 (O_304,N_29677,N_27297);
nand UO_305 (O_305,N_26262,N_25668);
nor UO_306 (O_306,N_27338,N_25243);
and UO_307 (O_307,N_24975,N_26643);
and UO_308 (O_308,N_27704,N_28007);
or UO_309 (O_309,N_27552,N_24383);
xor UO_310 (O_310,N_25736,N_24644);
nor UO_311 (O_311,N_26577,N_29927);
xnor UO_312 (O_312,N_27842,N_27106);
xnor UO_313 (O_313,N_24050,N_25958);
and UO_314 (O_314,N_28814,N_27326);
nand UO_315 (O_315,N_24955,N_24736);
nor UO_316 (O_316,N_27940,N_29180);
xnor UO_317 (O_317,N_25608,N_24275);
nor UO_318 (O_318,N_26999,N_25459);
nor UO_319 (O_319,N_24589,N_24663);
and UO_320 (O_320,N_29773,N_26593);
xor UO_321 (O_321,N_29737,N_27080);
nand UO_322 (O_322,N_26213,N_24247);
xor UO_323 (O_323,N_24344,N_27641);
xnor UO_324 (O_324,N_28330,N_24446);
or UO_325 (O_325,N_25383,N_29393);
xnor UO_326 (O_326,N_29845,N_28409);
nor UO_327 (O_327,N_26289,N_24811);
nand UO_328 (O_328,N_25115,N_26409);
nor UO_329 (O_329,N_26205,N_28195);
nand UO_330 (O_330,N_24675,N_25470);
xnor UO_331 (O_331,N_24727,N_26722);
nor UO_332 (O_332,N_27746,N_26504);
or UO_333 (O_333,N_26203,N_24303);
nor UO_334 (O_334,N_25400,N_29163);
nor UO_335 (O_335,N_24047,N_24636);
and UO_336 (O_336,N_26500,N_25082);
and UO_337 (O_337,N_29140,N_27008);
and UO_338 (O_338,N_28867,N_25105);
xor UO_339 (O_339,N_24915,N_29675);
nand UO_340 (O_340,N_27402,N_24735);
xnor UO_341 (O_341,N_25932,N_26965);
and UO_342 (O_342,N_26299,N_28315);
xor UO_343 (O_343,N_29062,N_26899);
xor UO_344 (O_344,N_24346,N_28067);
xor UO_345 (O_345,N_25791,N_26653);
nor UO_346 (O_346,N_24262,N_29514);
or UO_347 (O_347,N_29158,N_25424);
xnor UO_348 (O_348,N_25012,N_29765);
or UO_349 (O_349,N_29228,N_24909);
and UO_350 (O_350,N_27239,N_29674);
xnor UO_351 (O_351,N_28024,N_24876);
nand UO_352 (O_352,N_24187,N_24622);
xor UO_353 (O_353,N_24381,N_25055);
or UO_354 (O_354,N_27231,N_25709);
nand UO_355 (O_355,N_25779,N_25561);
nand UO_356 (O_356,N_24259,N_25442);
nand UO_357 (O_357,N_29444,N_28379);
xor UO_358 (O_358,N_29361,N_27897);
and UO_359 (O_359,N_25934,N_29162);
nand UO_360 (O_360,N_29559,N_25054);
and UO_361 (O_361,N_25378,N_28029);
or UO_362 (O_362,N_29079,N_29763);
nand UO_363 (O_363,N_27137,N_29989);
or UO_364 (O_364,N_27058,N_26161);
or UO_365 (O_365,N_27443,N_27753);
and UO_366 (O_366,N_25103,N_29711);
nor UO_367 (O_367,N_28981,N_24616);
and UO_368 (O_368,N_24512,N_29309);
xor UO_369 (O_369,N_29591,N_27274);
xor UO_370 (O_370,N_27428,N_24193);
or UO_371 (O_371,N_27122,N_26698);
nand UO_372 (O_372,N_28752,N_27550);
nand UO_373 (O_373,N_25615,N_26843);
and UO_374 (O_374,N_29461,N_28283);
and UO_375 (O_375,N_27996,N_29131);
xor UO_376 (O_376,N_25326,N_24508);
nor UO_377 (O_377,N_29397,N_25689);
nor UO_378 (O_378,N_24894,N_29336);
or UO_379 (O_379,N_28003,N_27065);
or UO_380 (O_380,N_25068,N_26106);
or UO_381 (O_381,N_28060,N_24442);
or UO_382 (O_382,N_24336,N_26917);
nor UO_383 (O_383,N_25530,N_25931);
xnor UO_384 (O_384,N_28238,N_29731);
nand UO_385 (O_385,N_24559,N_28180);
nand UO_386 (O_386,N_28122,N_28700);
or UO_387 (O_387,N_28295,N_24170);
or UO_388 (O_388,N_26694,N_25016);
and UO_389 (O_389,N_27123,N_24198);
nor UO_390 (O_390,N_26302,N_28995);
nor UO_391 (O_391,N_27812,N_26090);
and UO_392 (O_392,N_28960,N_27529);
xnor UO_393 (O_393,N_27077,N_24342);
xor UO_394 (O_394,N_24300,N_27203);
nand UO_395 (O_395,N_29220,N_26538);
nand UO_396 (O_396,N_25379,N_25397);
and UO_397 (O_397,N_24026,N_25085);
xor UO_398 (O_398,N_27395,N_27578);
nor UO_399 (O_399,N_25551,N_27250);
nand UO_400 (O_400,N_26064,N_27210);
nor UO_401 (O_401,N_25808,N_24942);
xor UO_402 (O_402,N_28843,N_27344);
or UO_403 (O_403,N_26661,N_24405);
xnor UO_404 (O_404,N_28173,N_28524);
and UO_405 (O_405,N_25684,N_26931);
xnor UO_406 (O_406,N_28366,N_27321);
or UO_407 (O_407,N_25346,N_29226);
and UO_408 (O_408,N_26480,N_26613);
or UO_409 (O_409,N_29057,N_25034);
nand UO_410 (O_410,N_29982,N_27827);
nand UO_411 (O_411,N_24482,N_28095);
nor UO_412 (O_412,N_26624,N_27258);
and UO_413 (O_413,N_24217,N_24797);
nand UO_414 (O_414,N_29756,N_29868);
and UO_415 (O_415,N_24453,N_25565);
nor UO_416 (O_416,N_27586,N_27324);
and UO_417 (O_417,N_26476,N_29383);
or UO_418 (O_418,N_28571,N_29650);
nand UO_419 (O_419,N_28461,N_27090);
xnor UO_420 (O_420,N_26640,N_24255);
and UO_421 (O_421,N_29476,N_27789);
xor UO_422 (O_422,N_29999,N_28388);
nor UO_423 (O_423,N_26535,N_24196);
and UO_424 (O_424,N_26712,N_24285);
nand UO_425 (O_425,N_24222,N_27530);
and UO_426 (O_426,N_25559,N_28831);
or UO_427 (O_427,N_29415,N_26430);
xnor UO_428 (O_428,N_29742,N_26129);
nor UO_429 (O_429,N_27282,N_27234);
nand UO_430 (O_430,N_24803,N_29225);
nand UO_431 (O_431,N_24786,N_29853);
nand UO_432 (O_432,N_25290,N_24816);
or UO_433 (O_433,N_26216,N_28400);
nor UO_434 (O_434,N_28922,N_27034);
and UO_435 (O_435,N_29268,N_27179);
xnor UO_436 (O_436,N_25456,N_28909);
xor UO_437 (O_437,N_28896,N_26327);
and UO_438 (O_438,N_29892,N_26960);
nand UO_439 (O_439,N_29735,N_24969);
nor UO_440 (O_440,N_28457,N_28150);
nand UO_441 (O_441,N_24349,N_25949);
nor UO_442 (O_442,N_29481,N_25464);
nor UO_443 (O_443,N_29520,N_29432);
and UO_444 (O_444,N_26276,N_28604);
and UO_445 (O_445,N_29656,N_27614);
and UO_446 (O_446,N_29059,N_25628);
nand UO_447 (O_447,N_26976,N_29177);
xnor UO_448 (O_448,N_26709,N_25171);
or UO_449 (O_449,N_26217,N_27335);
xnor UO_450 (O_450,N_28743,N_29776);
nor UO_451 (O_451,N_26058,N_29870);
nor UO_452 (O_452,N_27643,N_26159);
nand UO_453 (O_453,N_29692,N_26849);
nand UO_454 (O_454,N_25963,N_26375);
and UO_455 (O_455,N_28492,N_28297);
xnor UO_456 (O_456,N_24338,N_28663);
or UO_457 (O_457,N_26073,N_27664);
nand UO_458 (O_458,N_24698,N_29622);
or UO_459 (O_459,N_25189,N_29109);
nand UO_460 (O_460,N_24662,N_29026);
and UO_461 (O_461,N_24110,N_28145);
and UO_462 (O_462,N_25353,N_24327);
and UO_463 (O_463,N_25035,N_29893);
nor UO_464 (O_464,N_28855,N_26108);
nand UO_465 (O_465,N_24326,N_27806);
xor UO_466 (O_466,N_24030,N_28065);
and UO_467 (O_467,N_25880,N_29990);
or UO_468 (O_468,N_28022,N_26393);
and UO_469 (O_469,N_28742,N_28241);
nand UO_470 (O_470,N_24755,N_28345);
or UO_471 (O_471,N_26022,N_25771);
or UO_472 (O_472,N_29241,N_25308);
xnor UO_473 (O_473,N_27539,N_28070);
nand UO_474 (O_474,N_28623,N_25796);
nand UO_475 (O_475,N_29369,N_24523);
nand UO_476 (O_476,N_28906,N_24837);
and UO_477 (O_477,N_28316,N_28757);
and UO_478 (O_478,N_29956,N_29113);
and UO_479 (O_479,N_27477,N_29582);
nor UO_480 (O_480,N_24793,N_26702);
nor UO_481 (O_481,N_27378,N_28452);
nand UO_482 (O_482,N_25373,N_27066);
nor UO_483 (O_483,N_28063,N_28470);
nor UO_484 (O_484,N_27255,N_26183);
and UO_485 (O_485,N_24408,N_26253);
xnor UO_486 (O_486,N_26318,N_24652);
xnor UO_487 (O_487,N_28779,N_28149);
xnor UO_488 (O_488,N_27033,N_28390);
nand UO_489 (O_489,N_26874,N_28487);
nor UO_490 (O_490,N_27037,N_24764);
and UO_491 (O_491,N_29096,N_25956);
nand UO_492 (O_492,N_25460,N_25872);
and UO_493 (O_493,N_24307,N_28620);
or UO_494 (O_494,N_29327,N_29803);
xor UO_495 (O_495,N_24946,N_26676);
nor UO_496 (O_496,N_29513,N_26320);
and UO_497 (O_497,N_28832,N_24653);
and UO_498 (O_498,N_25544,N_29707);
xor UO_499 (O_499,N_24464,N_26131);
or UO_500 (O_500,N_28042,N_25089);
or UO_501 (O_501,N_24831,N_26221);
and UO_502 (O_502,N_24416,N_27676);
or UO_503 (O_503,N_25560,N_24592);
or UO_504 (O_504,N_24322,N_25910);
nand UO_505 (O_505,N_25153,N_27259);
or UO_506 (O_506,N_27963,N_26592);
xor UO_507 (O_507,N_28507,N_27269);
or UO_508 (O_508,N_28310,N_27703);
nand UO_509 (O_509,N_28785,N_25321);
xnor UO_510 (O_510,N_24302,N_27667);
nand UO_511 (O_511,N_24041,N_24777);
or UO_512 (O_512,N_26803,N_29022);
nand UO_513 (O_513,N_25246,N_26607);
or UO_514 (O_514,N_27646,N_28563);
or UO_515 (O_515,N_26436,N_29418);
and UO_516 (O_516,N_29382,N_27079);
or UO_517 (O_517,N_24753,N_25802);
and UO_518 (O_518,N_24265,N_29414);
xor UO_519 (O_519,N_27632,N_24542);
or UO_520 (O_520,N_28091,N_26188);
or UO_521 (O_521,N_25492,N_27273);
and UO_522 (O_522,N_29748,N_27217);
and UO_523 (O_523,N_28044,N_24602);
nand UO_524 (O_524,N_24171,N_24708);
or UO_525 (O_525,N_25823,N_27086);
xor UO_526 (O_526,N_24612,N_28749);
nor UO_527 (O_527,N_24889,N_25770);
or UO_528 (O_528,N_24369,N_25967);
xnor UO_529 (O_529,N_24438,N_28876);
or UO_530 (O_530,N_25760,N_25899);
nand UO_531 (O_531,N_24918,N_27296);
or UO_532 (O_532,N_27764,N_27301);
xnor UO_533 (O_533,N_29210,N_24325);
or UO_534 (O_534,N_28941,N_29952);
xnor UO_535 (O_535,N_25635,N_25162);
nand UO_536 (O_536,N_25557,N_26605);
xnor UO_537 (O_537,N_29121,N_28518);
or UO_538 (O_538,N_25629,N_28872);
nor UO_539 (O_539,N_25230,N_25349);
xor UO_540 (O_540,N_29195,N_26048);
nor UO_541 (O_541,N_27526,N_29993);
and UO_542 (O_542,N_24479,N_26881);
nor UO_543 (O_543,N_25393,N_26595);
nand UO_544 (O_544,N_25840,N_25022);
or UO_545 (O_545,N_28146,N_28706);
or UO_546 (O_546,N_24162,N_25363);
or UO_547 (O_547,N_24967,N_27655);
nand UO_548 (O_548,N_29583,N_28155);
nand UO_549 (O_549,N_28054,N_24473);
nor UO_550 (O_550,N_29833,N_27745);
or UO_551 (O_551,N_29515,N_26778);
or UO_552 (O_552,N_29396,N_24328);
nand UO_553 (O_553,N_24529,N_29028);
nor UO_554 (O_554,N_29814,N_27849);
and UO_555 (O_555,N_29823,N_27442);
xor UO_556 (O_556,N_27823,N_25439);
nor UO_557 (O_557,N_28553,N_24990);
nand UO_558 (O_558,N_27837,N_28575);
and UO_559 (O_559,N_25656,N_24175);
nor UO_560 (O_560,N_29655,N_25957);
or UO_561 (O_561,N_28422,N_26867);
xnor UO_562 (O_562,N_26135,N_27459);
nand UO_563 (O_563,N_29947,N_25275);
or UO_564 (O_564,N_27628,N_24091);
nor UO_565 (O_565,N_24899,N_29416);
nand UO_566 (O_566,N_28616,N_28593);
xor UO_567 (O_567,N_27414,N_24574);
nor UO_568 (O_568,N_27315,N_25360);
nand UO_569 (O_569,N_26513,N_28143);
xor UO_570 (O_570,N_27240,N_24413);
and UO_571 (O_571,N_24053,N_27887);
and UO_572 (O_572,N_28410,N_25306);
or UO_573 (O_573,N_28674,N_29135);
nor UO_574 (O_574,N_29722,N_28611);
nor UO_575 (O_575,N_28665,N_29596);
xnor UO_576 (O_576,N_29483,N_27811);
nor UO_577 (O_577,N_24759,N_28817);
nor UO_578 (O_578,N_24567,N_25909);
and UO_579 (O_579,N_24415,N_27497);
or UO_580 (O_580,N_28336,N_29100);
nor UO_581 (O_581,N_29876,N_26471);
and UO_582 (O_582,N_27286,N_27594);
and UO_583 (O_583,N_26710,N_28685);
nor UO_584 (O_584,N_24134,N_25604);
or UO_585 (O_585,N_26686,N_26440);
and UO_586 (O_586,N_29171,N_29652);
and UO_587 (O_587,N_24809,N_29101);
nor UO_588 (O_588,N_29917,N_26332);
xor UO_589 (O_589,N_25592,N_25332);
nand UO_590 (O_590,N_28874,N_24599);
nor UO_591 (O_591,N_25785,N_27242);
or UO_592 (O_592,N_24019,N_26779);
nor UO_593 (O_593,N_25818,N_28482);
nand UO_594 (O_594,N_25472,N_25260);
nand UO_595 (O_595,N_24182,N_26359);
or UO_596 (O_596,N_25504,N_29261);
nor UO_597 (O_597,N_26856,N_25858);
xor UO_598 (O_598,N_27169,N_26903);
and UO_599 (O_599,N_29474,N_25505);
xor UO_600 (O_600,N_26335,N_24407);
xnor UO_601 (O_601,N_26123,N_26011);
and UO_602 (O_602,N_26155,N_29574);
and UO_603 (O_603,N_24425,N_29159);
or UO_604 (O_604,N_25575,N_27386);
nand UO_605 (O_605,N_26793,N_24447);
xnor UO_606 (O_606,N_25838,N_26241);
and UO_607 (O_607,N_25168,N_25323);
xnor UO_608 (O_608,N_25977,N_29482);
nor UO_609 (O_609,N_24791,N_27243);
nor UO_610 (O_610,N_25392,N_26732);
nor UO_611 (O_611,N_29613,N_26224);
and UO_612 (O_612,N_27795,N_26708);
and UO_613 (O_613,N_28755,N_27470);
nor UO_614 (O_614,N_25904,N_28801);
and UO_615 (O_615,N_27009,N_27499);
nand UO_616 (O_616,N_24631,N_25023);
and UO_617 (O_617,N_24229,N_28727);
or UO_618 (O_618,N_29292,N_24431);
and UO_619 (O_619,N_25118,N_27303);
or UO_620 (O_620,N_28434,N_29428);
and UO_621 (O_621,N_28810,N_25108);
and UO_622 (O_622,N_25176,N_27455);
nor UO_623 (O_623,N_27207,N_24858);
nor UO_624 (O_624,N_26469,N_24751);
and UO_625 (O_625,N_29680,N_28971);
and UO_626 (O_626,N_24970,N_26039);
or UO_627 (O_627,N_26312,N_25251);
nor UO_628 (O_628,N_27343,N_28595);
and UO_629 (O_629,N_27310,N_29528);
and UO_630 (O_630,N_29598,N_27192);
nor UO_631 (O_631,N_27075,N_29165);
and UO_632 (O_632,N_27997,N_25427);
or UO_633 (O_633,N_27480,N_27778);
xnor UO_634 (O_634,N_26758,N_29953);
xor UO_635 (O_635,N_28268,N_28374);
or UO_636 (O_636,N_29715,N_25386);
nand UO_637 (O_637,N_24991,N_28105);
or UO_638 (O_638,N_29164,N_28321);
xor UO_639 (O_639,N_24203,N_28833);
xor UO_640 (O_640,N_25469,N_28159);
xnor UO_641 (O_641,N_28228,N_28017);
and UO_642 (O_642,N_29533,N_26908);
or UO_643 (O_643,N_29014,N_25283);
nand UO_644 (O_644,N_24769,N_28207);
or UO_645 (O_645,N_24496,N_25694);
xnor UO_646 (O_646,N_24471,N_25891);
nor UO_647 (O_647,N_25101,N_25478);
or UO_648 (O_648,N_25088,N_29848);
or UO_649 (O_649,N_28333,N_26255);
nor UO_650 (O_650,N_26143,N_24423);
xor UO_651 (O_651,N_27222,N_26567);
or UO_652 (O_652,N_25074,N_27405);
or UO_653 (O_653,N_29951,N_27903);
xnor UO_654 (O_654,N_29130,N_29018);
nor UO_655 (O_655,N_29585,N_24499);
and UO_656 (O_656,N_29005,N_25974);
nand UO_657 (O_657,N_28291,N_28196);
nand UO_658 (O_658,N_25036,N_28197);
and UO_659 (O_659,N_28356,N_24131);
nand UO_660 (O_660,N_24707,N_26173);
nor UO_661 (O_661,N_27661,N_24532);
nor UO_662 (O_662,N_27965,N_27724);
and UO_663 (O_663,N_29271,N_28750);
nand UO_664 (O_664,N_26875,N_26752);
nand UO_665 (O_665,N_26602,N_24297);
nor UO_666 (O_666,N_27723,N_25987);
xnor UO_667 (O_667,N_29123,N_25446);
and UO_668 (O_668,N_28157,N_24308);
nor UO_669 (O_669,N_29787,N_25384);
or UO_670 (O_670,N_29755,N_28510);
and UO_671 (O_671,N_26337,N_29029);
or UO_672 (O_672,N_25679,N_29352);
nor UO_673 (O_673,N_25991,N_28799);
xnor UO_674 (O_674,N_24829,N_28491);
or UO_675 (O_675,N_26958,N_25370);
nor UO_676 (O_676,N_24331,N_29152);
nor UO_677 (O_677,N_24172,N_26095);
nor UO_678 (O_678,N_25011,N_29251);
nor UO_679 (O_679,N_25501,N_29985);
and UO_680 (O_680,N_26879,N_29030);
nand UO_681 (O_681,N_26590,N_27781);
and UO_682 (O_682,N_26324,N_24699);
nand UO_683 (O_683,N_25644,N_26912);
and UO_684 (O_684,N_26723,N_28164);
xnor UO_685 (O_685,N_27061,N_29712);
nor UO_686 (O_686,N_29146,N_25325);
nand UO_687 (O_687,N_26824,N_29566);
nor UO_688 (O_688,N_27263,N_25843);
nor UO_689 (O_689,N_24002,N_24546);
nor UO_690 (O_690,N_27517,N_28349);
xnor UO_691 (O_691,N_24659,N_29119);
and UO_692 (O_692,N_24904,N_28579);
and UO_693 (O_693,N_27859,N_25262);
or UO_694 (O_694,N_24324,N_25609);
and UO_695 (O_695,N_26925,N_28289);
nor UO_696 (O_696,N_26380,N_24368);
nand UO_697 (O_697,N_28458,N_29412);
nor UO_698 (O_698,N_26168,N_25651);
nor UO_699 (O_699,N_28169,N_25666);
nor UO_700 (O_700,N_27364,N_26558);
and UO_701 (O_701,N_25758,N_28097);
xnor UO_702 (O_702,N_27548,N_25057);
and UO_703 (O_703,N_26377,N_27126);
or UO_704 (O_704,N_26933,N_26611);
and UO_705 (O_705,N_27410,N_27896);
or UO_706 (O_706,N_25936,N_27462);
nor UO_707 (O_707,N_27919,N_26493);
and UO_708 (O_708,N_24127,N_26986);
or UO_709 (O_709,N_29359,N_29311);
nor UO_710 (O_710,N_29726,N_29017);
or UO_711 (O_711,N_24335,N_29553);
xnor UO_712 (O_712,N_28708,N_27544);
and UO_713 (O_713,N_24364,N_25959);
or UO_714 (O_714,N_28002,N_25437);
and UO_715 (O_715,N_25324,N_26071);
nand UO_716 (O_716,N_29325,N_25149);
xnor UO_717 (O_717,N_26279,N_26663);
xnor UO_718 (O_718,N_25898,N_29536);
and UO_719 (O_719,N_27472,N_26435);
and UO_720 (O_720,N_25491,N_29685);
or UO_721 (O_721,N_27830,N_29550);
or UO_722 (O_722,N_24634,N_27779);
and UO_723 (O_723,N_26460,N_27657);
and UO_724 (O_724,N_27729,N_28193);
nand UO_725 (O_725,N_29367,N_27440);
nand UO_726 (O_726,N_29042,N_26678);
nor UO_727 (O_727,N_26919,N_27736);
and UO_728 (O_728,N_28201,N_27658);
nor UO_729 (O_729,N_25582,N_27777);
xor UO_730 (O_730,N_27960,N_28529);
nor UO_731 (O_731,N_29943,N_27767);
xor UO_732 (O_732,N_26531,N_27162);
nor UO_733 (O_733,N_29555,N_25761);
nand UO_734 (O_734,N_25221,N_29063);
nor UO_735 (O_735,N_24034,N_26304);
xnor UO_736 (O_736,N_26647,N_29388);
or UO_737 (O_737,N_28609,N_24848);
xnor UO_738 (O_738,N_26928,N_29970);
or UO_739 (O_739,N_27999,N_27654);
and UO_740 (O_740,N_27116,N_27748);
and UO_741 (O_741,N_26799,N_26163);
nor UO_742 (O_742,N_28737,N_24008);
nor UO_743 (O_743,N_27370,N_25214);
xor UO_744 (O_744,N_24073,N_29913);
nand UO_745 (O_745,N_27540,N_26290);
or UO_746 (O_746,N_26984,N_25045);
or UO_747 (O_747,N_24912,N_27436);
nand UO_748 (O_748,N_25161,N_24875);
or UO_749 (O_749,N_28701,N_28996);
and UO_750 (O_750,N_26832,N_26057);
nor UO_751 (O_751,N_24554,N_28933);
nor UO_752 (O_752,N_25871,N_27278);
and UO_753 (O_753,N_24434,N_28104);
or UO_754 (O_754,N_28747,N_28370);
nand UO_755 (O_755,N_28532,N_28715);
and UO_756 (O_756,N_25507,N_24483);
or UO_757 (O_757,N_29303,N_25047);
xor UO_758 (O_758,N_28741,N_27922);
or UO_759 (O_759,N_24743,N_28978);
nor UO_760 (O_760,N_28884,N_26939);
or UO_761 (O_761,N_25072,N_26724);
or UO_762 (O_762,N_28690,N_28364);
xor UO_763 (O_763,N_26305,N_28040);
and UO_764 (O_764,N_29285,N_27159);
nor UO_765 (O_765,N_26581,N_28676);
xnor UO_766 (O_766,N_27356,N_24076);
xnor UO_767 (O_767,N_28800,N_27291);
xor UO_768 (O_768,N_26059,N_26625);
and UO_769 (O_769,N_25762,N_24293);
nand UO_770 (O_770,N_27142,N_26272);
nor UO_771 (O_771,N_28754,N_27229);
or UO_772 (O_772,N_28853,N_29132);
or UO_773 (O_773,N_26868,N_29662);
nand UO_774 (O_774,N_26616,N_28630);
xor UO_775 (O_775,N_29201,N_24609);
nor UO_776 (O_776,N_27127,N_24205);
xor UO_777 (O_777,N_24832,N_26223);
nor UO_778 (O_778,N_24052,N_26465);
or UO_779 (O_779,N_27285,N_29006);
nor UO_780 (O_780,N_25233,N_25225);
or UO_781 (O_781,N_28905,N_24879);
or UO_782 (O_782,N_28365,N_26475);
xnor UO_783 (O_783,N_24279,N_26271);
nor UO_784 (O_784,N_25313,N_28930);
nor UO_785 (O_785,N_24107,N_25164);
xnor UO_786 (O_786,N_28484,N_26964);
and UO_787 (O_787,N_26498,N_24916);
nand UO_788 (O_788,N_26032,N_25687);
xnor UO_789 (O_789,N_29021,N_26153);
or UO_790 (O_790,N_27649,N_29922);
nand UO_791 (O_791,N_26578,N_26070);
nand UO_792 (O_792,N_27546,N_28446);
nand UO_793 (O_793,N_28636,N_25050);
or UO_794 (O_794,N_28983,N_24621);
nand UO_795 (O_795,N_25806,N_24891);
xor UO_796 (O_796,N_26894,N_27618);
and UO_797 (O_797,N_29051,N_24866);
or UO_798 (O_798,N_25357,N_25003);
nor UO_799 (O_799,N_27005,N_27391);
or UO_800 (O_800,N_24932,N_28231);
nand UO_801 (O_801,N_27564,N_27444);
xor UO_802 (O_802,N_25404,N_24814);
and UO_803 (O_803,N_28907,N_29340);
nand UO_804 (O_804,N_24487,N_24613);
nor UO_805 (O_805,N_26142,N_27966);
or UO_806 (O_806,N_28761,N_24319);
or UO_807 (O_807,N_28686,N_25447);
nor UO_808 (O_808,N_28966,N_27396);
xnor UO_809 (O_809,N_25000,N_24371);
nand UO_810 (O_810,N_29704,N_26834);
nand UO_811 (O_811,N_26177,N_26387);
xor UO_812 (O_812,N_26099,N_29266);
and UO_813 (O_813,N_25265,N_24045);
nor UO_814 (O_814,N_25348,N_26701);
xnor UO_815 (O_815,N_29589,N_29784);
and UO_816 (O_816,N_27487,N_29061);
nand UO_817 (O_817,N_27184,N_29799);
xor UO_818 (O_818,N_28352,N_24506);
nand UO_819 (O_819,N_29007,N_25617);
nor UO_820 (O_820,N_25069,N_27568);
or UO_821 (O_821,N_25930,N_25916);
nor UO_822 (O_822,N_25902,N_24728);
and UO_823 (O_823,N_26425,N_29442);
nor UO_824 (O_824,N_24226,N_25856);
nand UO_825 (O_825,N_25063,N_28829);
and UO_826 (O_826,N_26987,N_26418);
nand UO_827 (O_827,N_29435,N_26932);
xnor UO_828 (O_828,N_29089,N_29971);
and UO_829 (O_829,N_27727,N_29542);
and UO_830 (O_830,N_25124,N_24151);
nand UO_831 (O_831,N_29549,N_27865);
nor UO_832 (O_832,N_27785,N_25395);
nand UO_833 (O_833,N_25517,N_29950);
nor UO_834 (O_834,N_24418,N_28371);
or UO_835 (O_835,N_29752,N_29812);
and UO_836 (O_836,N_25499,N_25033);
or UO_837 (O_837,N_27974,N_24937);
and UO_838 (O_838,N_28649,N_27675);
nor UO_839 (O_839,N_29693,N_27064);
nand UO_840 (O_840,N_29199,N_26774);
or UO_841 (O_841,N_29139,N_29665);
or UO_842 (O_842,N_28625,N_26817);
and UO_843 (O_843,N_26474,N_24711);
xnor UO_844 (O_844,N_28631,N_27484);
nand UO_845 (O_845,N_28072,N_27024);
xor UO_846 (O_846,N_26240,N_29078);
or UO_847 (O_847,N_27716,N_29670);
xnor UO_848 (O_848,N_26006,N_25037);
or UO_849 (O_849,N_25623,N_24142);
and UO_850 (O_850,N_29925,N_27740);
or UO_851 (O_851,N_27085,N_25801);
or UO_852 (O_852,N_29055,N_24206);
nor UO_853 (O_853,N_26734,N_24139);
and UO_854 (O_854,N_27399,N_26730);
nand UO_855 (O_855,N_26942,N_24593);
nor UO_856 (O_856,N_26254,N_28006);
nand UO_857 (O_857,N_28895,N_28324);
xnor UO_858 (O_858,N_25166,N_27995);
nor UO_859 (O_859,N_26348,N_24054);
and UO_860 (O_860,N_29054,N_27031);
or UO_861 (O_861,N_27451,N_28528);
nor UO_862 (O_862,N_29420,N_24213);
nand UO_863 (O_863,N_29387,N_27104);
nand UO_864 (O_864,N_27121,N_29038);
and UO_865 (O_865,N_25078,N_25172);
or UO_866 (O_866,N_24584,N_27773);
xnor UO_867 (O_867,N_25155,N_29479);
or UO_868 (O_868,N_24065,N_26739);
nand UO_869 (O_869,N_27481,N_29157);
or UO_870 (O_870,N_27979,N_24223);
or UO_871 (O_871,N_26628,N_24195);
or UO_872 (O_872,N_25704,N_24933);
xnor UO_873 (O_873,N_29614,N_26025);
or UO_874 (O_874,N_24116,N_28650);
xor UO_875 (O_875,N_29283,N_24525);
nand UO_876 (O_876,N_25268,N_27515);
xnor UO_877 (O_877,N_27412,N_24046);
nor UO_878 (O_878,N_27206,N_28688);
or UO_879 (O_879,N_25208,N_25245);
or UO_880 (O_880,N_29534,N_28009);
nand UO_881 (O_881,N_28918,N_24489);
and UO_882 (O_882,N_26145,N_25913);
nor UO_883 (O_883,N_24531,N_26645);
nand UO_884 (O_884,N_28722,N_25630);
and UO_885 (O_885,N_26761,N_25654);
xor UO_886 (O_886,N_26680,N_26189);
or UO_887 (O_887,N_26004,N_26784);
xnor UO_888 (O_888,N_25866,N_25752);
and UO_889 (O_889,N_29638,N_29954);
and UO_890 (O_890,N_28189,N_28064);
xnor UO_891 (O_891,N_24782,N_25855);
xnor UO_892 (O_892,N_28633,N_29607);
or UO_893 (O_893,N_27447,N_27637);
nor UO_894 (O_894,N_24449,N_28709);
nand UO_895 (O_895,N_27520,N_25800);
xnor UO_896 (O_896,N_24236,N_26260);
nor UO_897 (O_897,N_25080,N_28443);
and UO_898 (O_898,N_25328,N_28842);
nor UO_899 (O_899,N_29400,N_26413);
or UO_900 (O_900,N_25523,N_27393);
and UO_901 (O_901,N_27873,N_26808);
nor UO_902 (O_902,N_27553,N_24216);
or UO_903 (O_903,N_26278,N_26926);
xor UO_904 (O_904,N_25599,N_28877);
nand UO_905 (O_905,N_26697,N_29230);
xor UO_906 (O_906,N_27877,N_27191);
or UO_907 (O_907,N_26234,N_29231);
xnor UO_908 (O_908,N_27264,N_27928);
or UO_909 (O_909,N_28448,N_24598);
xnor UO_910 (O_910,N_28257,N_26858);
and UO_911 (O_911,N_27339,N_27407);
nor UO_912 (O_912,N_27890,N_27171);
nor UO_913 (O_913,N_25886,N_25125);
xor UO_914 (O_914,N_29828,N_24128);
nand UO_915 (O_915,N_24746,N_25202);
nor UO_916 (O_916,N_29565,N_24849);
or UO_917 (O_917,N_27971,N_26795);
or UO_918 (O_918,N_28427,N_26453);
nor UO_919 (O_919,N_24796,N_27309);
nand UO_920 (O_920,N_26061,N_29262);
nand UO_921 (O_921,N_26017,N_24987);
xor UO_922 (O_922,N_25862,N_26167);
or UO_923 (O_923,N_24077,N_27015);
nor UO_924 (O_924,N_29380,N_24140);
xnor UO_925 (O_925,N_27702,N_29024);
nor UO_926 (O_926,N_28658,N_26533);
and UO_927 (O_927,N_25031,N_25019);
or UO_928 (O_928,N_29240,N_26983);
nor UO_929 (O_929,N_25345,N_26495);
nor UO_930 (O_930,N_25329,N_28634);
or UO_931 (O_931,N_24420,N_28758);
and UO_932 (O_932,N_24097,N_26132);
or UO_933 (O_933,N_25632,N_24863);
nand UO_934 (O_934,N_28694,N_28547);
and UO_935 (O_935,N_25610,N_29438);
nor UO_936 (O_936,N_25028,N_25964);
xnor UO_937 (O_937,N_26777,N_24360);
nor UO_938 (O_938,N_28956,N_24007);
nor UO_939 (O_939,N_29076,N_24029);
xnor UO_940 (O_940,N_28493,N_28375);
and UO_941 (O_941,N_29250,N_26688);
or UO_942 (O_942,N_29819,N_24463);
nor UO_943 (O_943,N_24370,N_29003);
xor UO_944 (O_944,N_25060,N_26519);
and UO_945 (O_945,N_26633,N_28353);
xnor UO_946 (O_946,N_24873,N_24838);
and UO_947 (O_947,N_27933,N_24424);
or UO_948 (O_948,N_26368,N_27011);
xnor UO_949 (O_949,N_29546,N_24982);
nand UO_950 (O_950,N_29944,N_26081);
and UO_951 (O_951,N_25600,N_24778);
xor UO_952 (O_952,N_24092,N_28840);
or UO_953 (O_953,N_26668,N_28498);
and UO_954 (O_954,N_28564,N_26316);
xnor UO_955 (O_955,N_24815,N_29842);
nand UO_956 (O_956,N_24667,N_25653);
and UO_957 (O_957,N_28659,N_25875);
or UO_958 (O_958,N_28429,N_26136);
nor UO_959 (O_959,N_28771,N_28859);
nor UO_960 (O_960,N_26112,N_25493);
nor UO_961 (O_961,N_26767,N_25121);
and UO_962 (O_962,N_26658,N_29817);
or UO_963 (O_963,N_26677,N_27056);
nor UO_964 (O_964,N_28865,N_26023);
and UO_965 (O_965,N_29487,N_26950);
nor UO_966 (O_966,N_28047,N_28726);
xnor UO_967 (O_967,N_29783,N_25699);
and UO_968 (O_968,N_27341,N_29182);
and UO_969 (O_969,N_27147,N_25591);
xor UO_970 (O_970,N_29181,N_29724);
nor UO_971 (O_971,N_28913,N_26574);
xor UO_972 (O_972,N_29966,N_26416);
and UO_973 (O_973,N_29278,N_27493);
xnor UO_974 (O_974,N_24422,N_26544);
nor UO_975 (O_975,N_26282,N_26609);
or UO_976 (O_976,N_28653,N_29847);
nor UO_977 (O_977,N_27498,N_26077);
and UO_978 (O_978,N_29260,N_27060);
and UO_979 (O_979,N_27140,N_28802);
xor UO_980 (O_980,N_29593,N_29295);
nand UO_981 (O_981,N_28118,N_25414);
and UO_982 (O_982,N_27287,N_26610);
and UO_983 (O_983,N_27895,N_26164);
nor UO_984 (O_984,N_25895,N_24466);
xor UO_985 (O_985,N_24081,N_29903);
nor UO_986 (O_986,N_24670,N_28991);
and UO_987 (O_987,N_27084,N_24742);
and UO_988 (O_988,N_27874,N_26514);
xor UO_989 (O_989,N_25798,N_28932);
nor UO_990 (O_990,N_24188,N_29716);
xnor UO_991 (O_991,N_24893,N_28121);
nor UO_992 (O_992,N_24716,N_26764);
xnor UO_993 (O_993,N_27554,N_27316);
nor UO_994 (O_994,N_26447,N_27183);
xnor UO_995 (O_995,N_26954,N_25953);
and UO_996 (O_996,N_27733,N_26499);
or UO_997 (O_997,N_26172,N_29430);
xor UO_998 (O_998,N_29935,N_26972);
or UO_999 (O_999,N_29304,N_28079);
or UO_1000 (O_1000,N_24395,N_26295);
xnor UO_1001 (O_1001,N_28166,N_26386);
xnor UO_1002 (O_1002,N_29102,N_27331);
nor UO_1003 (O_1003,N_28124,N_25835);
and UO_1004 (O_1004,N_27138,N_24132);
and UO_1005 (O_1005,N_28698,N_27292);
and UO_1006 (O_1006,N_25126,N_28953);
nand UO_1007 (O_1007,N_29404,N_26549);
xor UO_1008 (O_1008,N_24490,N_29429);
xnor UO_1009 (O_1009,N_28839,N_26369);
or UO_1010 (O_1010,N_25972,N_25718);
xnor UO_1011 (O_1011,N_29111,N_28432);
xnor UO_1012 (O_1012,N_26003,N_29807);
or UO_1013 (O_1013,N_26281,N_29658);
or UO_1014 (O_1014,N_28894,N_24785);
and UO_1015 (O_1015,N_24960,N_28467);
xor UO_1016 (O_1016,N_29247,N_28475);
and UO_1017 (O_1017,N_24648,N_29493);
xnor UO_1018 (O_1018,N_25278,N_26148);
nand UO_1019 (O_1019,N_27926,N_25220);
or UO_1020 (O_1020,N_25897,N_26110);
nand UO_1021 (O_1021,N_29590,N_28857);
and UO_1022 (O_1022,N_29385,N_29185);
and UO_1023 (O_1023,N_24561,N_25090);
nand UO_1024 (O_1024,N_28245,N_28451);
and UO_1025 (O_1025,N_27070,N_27419);
nand UO_1026 (O_1026,N_26363,N_29506);
xnor UO_1027 (O_1027,N_28893,N_25861);
and UO_1028 (O_1028,N_28026,N_26715);
nand UO_1029 (O_1029,N_24577,N_25940);
xor UO_1030 (O_1030,N_26736,N_26109);
xor UO_1031 (O_1031,N_25311,N_29901);
and UO_1032 (O_1032,N_27475,N_26819);
and UO_1033 (O_1033,N_28085,N_28537);
nand UO_1034 (O_1034,N_28441,N_28637);
nand UO_1035 (O_1035,N_26687,N_27495);
and UO_1036 (O_1036,N_25642,N_29979);
or UO_1037 (O_1037,N_29997,N_24406);
or UO_1038 (O_1038,N_24826,N_26751);
nor UO_1039 (O_1039,N_28190,N_28760);
nor UO_1040 (O_1040,N_24477,N_26792);
and UO_1041 (O_1041,N_26511,N_25803);
nand UO_1042 (O_1042,N_24251,N_28403);
nand UO_1043 (O_1043,N_29912,N_29867);
or UO_1044 (O_1044,N_29049,N_29798);
xnor UO_1045 (O_1045,N_27879,N_27622);
nand UO_1046 (O_1046,N_28186,N_27083);
nand UO_1047 (O_1047,N_25529,N_27609);
xor UO_1048 (O_1048,N_27862,N_25462);
and UO_1049 (O_1049,N_28416,N_26187);
or UO_1050 (O_1050,N_27124,N_24840);
and UO_1051 (O_1051,N_26019,N_27599);
xnor UO_1052 (O_1052,N_29746,N_24957);
nand UO_1053 (O_1053,N_24385,N_29379);
xnor UO_1054 (O_1054,N_24852,N_27109);
xor UO_1055 (O_1055,N_27565,N_28738);
and UO_1056 (O_1056,N_29727,N_25477);
nor UO_1057 (O_1057,N_29747,N_24779);
nor UO_1058 (O_1058,N_29488,N_29368);
xnor UO_1059 (O_1059,N_29307,N_28535);
and UO_1060 (O_1060,N_27021,N_25226);
or UO_1061 (O_1061,N_24160,N_27067);
xnor UO_1062 (O_1062,N_28606,N_28168);
nor UO_1063 (O_1063,N_26275,N_28975);
or UO_1064 (O_1064,N_25982,N_28519);
xor UO_1065 (O_1065,N_28092,N_27446);
nor UO_1066 (O_1066,N_25312,N_27131);
or UO_1067 (O_1067,N_29910,N_25431);
nor UO_1068 (O_1068,N_24819,N_25197);
and UO_1069 (O_1069,N_26659,N_25839);
xnor UO_1070 (O_1070,N_28980,N_28723);
and UO_1071 (O_1071,N_26382,N_27115);
and UO_1072 (O_1072,N_27575,N_27445);
or UO_1073 (O_1073,N_28469,N_25946);
nor UO_1074 (O_1074,N_26552,N_29338);
or UO_1075 (O_1075,N_25765,N_29104);
and UO_1076 (O_1076,N_26696,N_28967);
and UO_1077 (O_1077,N_26745,N_27361);
and UO_1078 (O_1078,N_29491,N_29405);
nor UO_1079 (O_1079,N_28271,N_28221);
nor UO_1080 (O_1080,N_29217,N_24956);
and UO_1081 (O_1081,N_28077,N_25662);
nand UO_1082 (O_1082,N_25344,N_24958);
nor UO_1083 (O_1083,N_24031,N_29223);
and UO_1084 (O_1084,N_28030,N_25244);
nand UO_1085 (O_1085,N_28073,N_24939);
nand UO_1086 (O_1086,N_24578,N_27177);
or UO_1087 (O_1087,N_27769,N_25776);
and UO_1088 (O_1088,N_28337,N_28259);
nand UO_1089 (O_1089,N_27110,N_29594);
nor UO_1090 (O_1090,N_28147,N_25377);
and UO_1091 (O_1091,N_24309,N_27078);
nand UO_1092 (O_1092,N_25334,N_25749);
nand UO_1093 (O_1093,N_29191,N_26853);
xnor UO_1094 (O_1094,N_28010,N_28638);
nor UO_1095 (O_1095,N_27561,N_27108);
xor UO_1096 (O_1096,N_24035,N_25834);
and UO_1097 (O_1097,N_29646,N_28938);
nor UO_1098 (O_1098,N_25302,N_24200);
or UO_1099 (O_1099,N_29218,N_26351);
or UO_1100 (O_1100,N_25231,N_26809);
nor UO_1101 (O_1101,N_28851,N_26264);
and UO_1102 (O_1102,N_25814,N_27422);
xnor UO_1103 (O_1103,N_24329,N_25708);
and UO_1104 (O_1104,N_29992,N_28341);
nand UO_1105 (O_1105,N_29212,N_26796);
xnor UO_1106 (O_1106,N_29073,N_29541);
or UO_1107 (O_1107,N_24071,N_27017);
nor UO_1108 (O_1108,N_26307,N_26557);
or UO_1109 (O_1109,N_29332,N_26907);
nand UO_1110 (O_1110,N_24082,N_24362);
xor UO_1111 (O_1111,N_28976,N_28234);
and UO_1112 (O_1112,N_27329,N_28151);
xnor UO_1113 (O_1113,N_29279,N_28982);
xnor UO_1114 (O_1114,N_24770,N_25240);
xnor UO_1115 (O_1115,N_28807,N_27826);
nand UO_1116 (O_1116,N_27398,N_28013);
and UO_1117 (O_1117,N_26484,N_24579);
nor UO_1118 (O_1118,N_29238,N_24450);
nor UO_1119 (O_1119,N_25025,N_29839);
and UO_1120 (O_1120,N_29431,N_26996);
or UO_1121 (O_1121,N_28687,N_24747);
xor UO_1122 (O_1122,N_28782,N_29371);
xnor UO_1123 (O_1123,N_29629,N_25249);
and UO_1124 (O_1124,N_27491,N_29540);
or UO_1125 (O_1125,N_29378,N_26442);
nand UO_1126 (O_1126,N_29227,N_24509);
nand UO_1127 (O_1127,N_28032,N_24212);
nand UO_1128 (O_1128,N_27340,N_26354);
nand UO_1129 (O_1129,N_29453,N_29239);
nor UO_1130 (O_1130,N_25882,N_29422);
nand UO_1131 (O_1131,N_28001,N_29771);
and UO_1132 (O_1132,N_28615,N_28950);
nand UO_1133 (O_1133,N_27245,N_24515);
xnor UO_1134 (O_1134,N_27595,N_29535);
nand UO_1135 (O_1135,N_26882,N_28137);
xor UO_1136 (O_1136,N_26360,N_27382);
and UO_1137 (O_1137,N_24270,N_28731);
and UO_1138 (O_1138,N_28642,N_29085);
and UO_1139 (O_1139,N_27429,N_24057);
or UO_1140 (O_1140,N_28130,N_28551);
nor UO_1141 (O_1141,N_29691,N_27592);
nand UO_1142 (O_1142,N_24113,N_24706);
and UO_1143 (O_1143,N_26766,N_25942);
and UO_1144 (O_1144,N_25659,N_28796);
xor UO_1145 (O_1145,N_26813,N_29170);
nand UO_1146 (O_1146,N_25132,N_24672);
and UO_1147 (O_1147,N_25374,N_24027);
xnor UO_1148 (O_1148,N_29035,N_28338);
nor UO_1149 (O_1149,N_25691,N_29841);
nand UO_1150 (O_1150,N_24268,N_29661);
and UO_1151 (O_1151,N_25369,N_25988);
nor UO_1152 (O_1152,N_29502,N_28215);
xor UO_1153 (O_1153,N_26831,N_27461);
nand UO_1154 (O_1154,N_25048,N_25454);
or UO_1155 (O_1155,N_28587,N_26209);
nand UO_1156 (O_1156,N_27682,N_28931);
nor UO_1157 (O_1157,N_28384,N_28573);
and UO_1158 (O_1158,N_27579,N_25495);
or UO_1159 (O_1159,N_29467,N_25284);
and UO_1160 (O_1160,N_24448,N_29112);
nor UO_1161 (O_1161,N_28942,N_28572);
xor UO_1162 (O_1162,N_25141,N_29060);
nand UO_1163 (O_1163,N_25317,N_25488);
nor UO_1164 (O_1164,N_24022,N_24588);
xnor UO_1165 (O_1165,N_25455,N_29710);
nor UO_1166 (O_1166,N_26780,N_28795);
nand UO_1167 (O_1167,N_28300,N_26515);
and UO_1168 (O_1168,N_27898,N_24089);
and UO_1169 (O_1169,N_29595,N_28612);
nor UO_1170 (O_1170,N_27300,N_28772);
nand UO_1171 (O_1171,N_26995,N_26691);
xnor UO_1172 (O_1172,N_27294,N_27813);
xnor UO_1173 (O_1173,N_29782,N_29363);
nand UO_1174 (O_1174,N_25099,N_29673);
xor UO_1175 (O_1175,N_29995,N_28962);
and UO_1176 (O_1176,N_29863,N_26138);
and UO_1177 (O_1177,N_28200,N_27288);
nand UO_1178 (O_1178,N_28911,N_27311);
or UO_1179 (O_1179,N_28501,N_28944);
nand UO_1180 (O_1180,N_24305,N_28014);
nand UO_1181 (O_1181,N_24973,N_24851);
xnor UO_1182 (O_1182,N_25678,N_29606);
and UO_1183 (O_1183,N_29668,N_29934);
nand UO_1184 (O_1184,N_29719,N_29904);
or UO_1185 (O_1185,N_28334,N_28635);
and UO_1186 (O_1186,N_25675,N_24730);
nand UO_1187 (O_1187,N_24885,N_27330);
and UO_1188 (O_1188,N_25224,N_27707);
nor UO_1189 (O_1189,N_29978,N_24282);
and UO_1190 (O_1190,N_24714,N_29044);
xor UO_1191 (O_1191,N_29468,N_27992);
nor UO_1192 (O_1192,N_24090,N_24871);
nand UO_1193 (O_1193,N_28920,N_25918);
nand UO_1194 (O_1194,N_27886,N_27521);
xor UO_1195 (O_1195,N_24610,N_25713);
nor UO_1196 (O_1196,N_26657,N_27144);
nor UO_1197 (O_1197,N_29118,N_25519);
nor UO_1198 (O_1198,N_25183,N_24507);
nor UO_1199 (O_1199,N_27002,N_25285);
and UO_1200 (O_1200,N_26270,N_26706);
or UO_1201 (O_1201,N_28664,N_29046);
and UO_1202 (O_1202,N_29013,N_28702);
or UO_1203 (O_1203,N_24553,N_25812);
or UO_1204 (O_1204,N_26198,N_27585);
nor UO_1205 (O_1205,N_29933,N_27362);
nand UO_1206 (O_1206,N_26747,N_28230);
or UO_1207 (O_1207,N_29206,N_26420);
or UO_1208 (O_1208,N_26267,N_29381);
xnor UO_1209 (O_1209,N_29584,N_29684);
and UO_1210 (O_1210,N_29911,N_25079);
or UO_1211 (O_1211,N_24938,N_24972);
and UO_1212 (O_1212,N_25342,N_28497);
xor UO_1213 (O_1213,N_28405,N_27929);
or UO_1214 (O_1214,N_29781,N_25543);
or UO_1215 (O_1215,N_27129,N_28273);
xnor UO_1216 (O_1216,N_25203,N_25158);
and UO_1217 (O_1217,N_28813,N_29600);
nand UO_1218 (O_1218,N_25714,N_24562);
and UO_1219 (O_1219,N_28514,N_27541);
or UO_1220 (O_1220,N_25865,N_26974);
nor UO_1221 (O_1221,N_27111,N_28657);
nand UO_1222 (O_1222,N_28119,N_28822);
nor UO_1223 (O_1223,N_26561,N_28672);
nor UO_1224 (O_1224,N_29654,N_27016);
or UO_1225 (O_1225,N_25747,N_27760);
or UO_1226 (O_1226,N_24676,N_24788);
and UO_1227 (O_1227,N_28088,N_28693);
xnor UO_1228 (O_1228,N_24260,N_27739);
nand UO_1229 (O_1229,N_29647,N_25819);
and UO_1230 (O_1230,N_27934,N_25948);
nor UO_1231 (O_1231,N_25624,N_24928);
nand UO_1232 (O_1232,N_28928,N_29053);
nor UO_1233 (O_1233,N_29229,N_25748);
nor UO_1234 (O_1234,N_24595,N_26871);
and UO_1235 (O_1235,N_29568,N_27917);
nor UO_1236 (O_1236,N_28294,N_29532);
nand UO_1237 (O_1237,N_25301,N_26280);
and UO_1238 (O_1238,N_29446,N_29306);
nand UO_1239 (O_1239,N_29374,N_27700);
nand UO_1240 (O_1240,N_27503,N_26119);
nor UO_1241 (O_1241,N_24497,N_27145);
nand UO_1242 (O_1242,N_24148,N_27559);
and UO_1243 (O_1243,N_25434,N_25541);
or UO_1244 (O_1244,N_26072,N_26456);
xnor UO_1245 (O_1245,N_27511,N_25331);
nand UO_1246 (O_1246,N_28590,N_26355);
nor UO_1247 (O_1247,N_28314,N_28993);
nand UO_1248 (O_1248,N_24929,N_29888);
xnor UO_1249 (O_1249,N_24158,N_29688);
or UO_1250 (O_1250,N_29445,N_29750);
nor UO_1251 (O_1251,N_24094,N_29644);
and UO_1252 (O_1252,N_26589,N_29980);
or UO_1253 (O_1253,N_24168,N_29844);
and UO_1254 (O_1254,N_29122,N_28125);
xnor UO_1255 (O_1255,N_26257,N_26556);
nand UO_1256 (O_1256,N_26895,N_28574);
and UO_1257 (O_1257,N_27039,N_27876);
and UO_1258 (O_1258,N_26617,N_25589);
nor UO_1259 (O_1259,N_26692,N_26953);
xor UO_1260 (O_1260,N_26945,N_26920);
nand UO_1261 (O_1261,N_26314,N_27755);
and UO_1262 (O_1262,N_27684,N_25503);
and UO_1263 (O_1263,N_25117,N_28994);
and UO_1264 (O_1264,N_29377,N_28011);
and UO_1265 (O_1265,N_25002,N_27730);
and UO_1266 (O_1266,N_27128,N_26103);
or UO_1267 (O_1267,N_27418,N_26412);
and UO_1268 (O_1268,N_27102,N_29441);
xor UO_1269 (O_1269,N_26127,N_28112);
xor UO_1270 (O_1270,N_24906,N_28732);
or UO_1271 (O_1271,N_28483,N_27763);
nand UO_1272 (O_1272,N_28279,N_27253);
or UO_1273 (O_1273,N_24294,N_26297);
or UO_1274 (O_1274,N_26598,N_27174);
nor UO_1275 (O_1275,N_28205,N_28847);
nor UO_1276 (O_1276,N_29071,N_24961);
nand UO_1277 (O_1277,N_26762,N_26905);
nor UO_1278 (O_1278,N_24888,N_28227);
xor UO_1279 (O_1279,N_28585,N_27761);
or UO_1280 (O_1280,N_24977,N_25809);
or UO_1281 (O_1281,N_26704,N_26580);
xor UO_1282 (O_1282,N_27947,N_27821);
nand UO_1283 (O_1283,N_27967,N_28647);
xor UO_1284 (O_1284,N_27215,N_29573);
nand UO_1285 (O_1285,N_29215,N_26507);
or UO_1286 (O_1286,N_24124,N_27780);
xnor UO_1287 (O_1287,N_25744,N_26893);
xor UO_1288 (O_1288,N_27132,N_24080);
xor UO_1289 (O_1289,N_27866,N_29759);
xor UO_1290 (O_1290,N_24807,N_27660);
nand UO_1291 (O_1291,N_29255,N_26269);
nor UO_1292 (O_1292,N_24629,N_28548);
nor UO_1293 (O_1293,N_25677,N_28825);
and UO_1294 (O_1294,N_24180,N_29766);
nor UO_1295 (O_1295,N_24566,N_26001);
xor UO_1296 (O_1296,N_25738,N_27380);
xor UO_1297 (O_1297,N_27196,N_27468);
or UO_1298 (O_1298,N_27099,N_25190);
nor UO_1299 (O_1299,N_26961,N_26488);
xnor UO_1300 (O_1300,N_27687,N_26904);
or UO_1301 (O_1301,N_26235,N_28765);
or UO_1302 (O_1302,N_27531,N_28710);
or UO_1303 (O_1303,N_26423,N_25482);
and UO_1304 (O_1304,N_24454,N_24374);
or UO_1305 (O_1305,N_26693,N_24596);
nor UO_1306 (O_1306,N_28614,N_24287);
nand UO_1307 (O_1307,N_25980,N_24834);
nand UO_1308 (O_1308,N_24980,N_27638);
xnor UO_1309 (O_1309,N_26261,N_28945);
nor UO_1310 (O_1310,N_24014,N_26098);
and UO_1311 (O_1311,N_26707,N_25920);
nor UO_1312 (O_1312,N_25279,N_28533);
or UO_1313 (O_1313,N_25657,N_25911);
or UO_1314 (O_1314,N_26943,N_26193);
nor UO_1315 (O_1315,N_28109,N_29873);
xnor UO_1316 (O_1316,N_25546,N_29643);
xor UO_1317 (O_1317,N_24626,N_29886);
xnor UO_1318 (O_1318,N_29504,N_25021);
nor UO_1319 (O_1319,N_25152,N_29762);
xor UO_1320 (O_1320,N_27148,N_27363);
or UO_1321 (O_1321,N_26096,N_27625);
and UO_1322 (O_1322,N_27328,N_29423);
or UO_1323 (O_1323,N_27327,N_28282);
nor UO_1324 (O_1324,N_25584,N_27822);
xor UO_1325 (O_1325,N_29270,N_25914);
and UO_1326 (O_1326,N_27199,N_28045);
nor UO_1327 (O_1327,N_25042,N_27101);
nand UO_1328 (O_1328,N_24443,N_26356);
or UO_1329 (O_1329,N_29517,N_29115);
nor UO_1330 (O_1330,N_29160,N_28835);
or UO_1331 (O_1331,N_27377,N_28915);
or UO_1332 (O_1332,N_27945,N_25463);
and UO_1333 (O_1333,N_25686,N_24351);
nor UO_1334 (O_1334,N_25550,N_28912);
nand UO_1335 (O_1335,N_28099,N_25211);
nor UO_1336 (O_1336,N_27634,N_28969);
nand UO_1337 (O_1337,N_25453,N_28711);
and UO_1338 (O_1338,N_24009,N_25100);
and UO_1339 (O_1339,N_24350,N_24332);
xnor UO_1340 (O_1340,N_25461,N_28331);
nor UO_1341 (O_1341,N_28272,N_27525);
xnor UO_1342 (O_1342,N_26835,N_25406);
or UO_1343 (O_1343,N_29019,N_28502);
xor UO_1344 (O_1344,N_27946,N_24850);
xor UO_1345 (O_1345,N_26104,N_28240);
or UO_1346 (O_1346,N_27421,N_26563);
and UO_1347 (O_1347,N_28730,N_29440);
xnor UO_1348 (O_1348,N_26911,N_25038);
nor UO_1349 (O_1349,N_24995,N_25128);
nor UO_1350 (O_1350,N_29615,N_27185);
or UO_1351 (O_1351,N_28404,N_29452);
nand UO_1352 (O_1352,N_27352,N_28517);
nor UO_1353 (O_1353,N_26811,N_29392);
or UO_1354 (O_1354,N_27049,N_27611);
and UO_1355 (O_1355,N_28419,N_28618);
or UO_1356 (O_1356,N_29968,N_27857);
xor UO_1357 (O_1357,N_28059,N_24164);
nor UO_1358 (O_1358,N_29907,N_28043);
or UO_1359 (O_1359,N_27091,N_28773);
nand UO_1360 (O_1360,N_25631,N_26765);
and UO_1361 (O_1361,N_28828,N_24024);
xor UO_1362 (O_1362,N_24119,N_25569);
or UO_1363 (O_1363,N_25663,N_24590);
xor UO_1364 (O_1364,N_27794,N_24810);
or UO_1365 (O_1365,N_27299,N_27502);
and UO_1366 (O_1366,N_29741,N_24086);
xor UO_1367 (O_1367,N_25768,N_29624);
or UO_1368 (O_1368,N_25945,N_29631);
and UO_1369 (O_1369,N_27656,N_27829);
nand UO_1370 (O_1370,N_25649,N_25282);
nand UO_1371 (O_1371,N_27796,N_28624);
nand UO_1372 (O_1372,N_26031,N_26719);
nand UO_1373 (O_1373,N_29946,N_25597);
or UO_1374 (O_1374,N_24643,N_27256);
nor UO_1375 (O_1375,N_29249,N_25497);
xor UO_1376 (O_1376,N_27855,N_27392);
or UO_1377 (O_1377,N_25912,N_25852);
xor UO_1378 (O_1378,N_29194,N_26035);
xor UO_1379 (O_1379,N_25636,N_29166);
and UO_1380 (O_1380,N_27617,N_29025);
nor UO_1381 (O_1381,N_24836,N_25741);
nor UO_1382 (O_1382,N_28815,N_28459);
nand UO_1383 (O_1383,N_28046,N_29544);
xnor UO_1384 (O_1384,N_25721,N_29065);
xnor UO_1385 (O_1385,N_27053,N_24535);
xnor UO_1386 (O_1386,N_25842,N_26763);
and UO_1387 (O_1387,N_27430,N_24722);
and UO_1388 (O_1388,N_25432,N_24697);
xor UO_1389 (O_1389,N_29880,N_28751);
nand UO_1390 (O_1390,N_26055,N_24230);
or UO_1391 (O_1391,N_26448,N_28021);
nor UO_1392 (O_1392,N_29257,N_28179);
nor UO_1393 (O_1393,N_27807,N_24994);
nor UO_1394 (O_1394,N_28387,N_24854);
or UO_1395 (O_1395,N_28447,N_24185);
or UO_1396 (O_1396,N_27743,N_26222);
nand UO_1397 (O_1397,N_26685,N_24358);
xor UO_1398 (O_1398,N_28823,N_26827);
and UO_1399 (O_1399,N_26776,N_27406);
nand UO_1400 (O_1400,N_26788,N_29941);
nor UO_1401 (O_1401,N_24741,N_28861);
or UO_1402 (O_1402,N_25836,N_27901);
nand UO_1403 (O_1403,N_25198,N_29334);
nand UO_1404 (O_1404,N_27348,N_26757);
xor UO_1405 (O_1405,N_28096,N_29312);
nor UO_1406 (O_1406,N_27885,N_27871);
nor UO_1407 (O_1407,N_28301,N_28204);
xor UO_1408 (O_1408,N_27146,N_26036);
xnor UO_1409 (O_1409,N_29964,N_29083);
nor UO_1410 (O_1410,N_25829,N_24280);
and UO_1411 (O_1411,N_27717,N_26956);
nand UO_1412 (O_1412,N_24537,N_27238);
or UO_1413 (O_1413,N_27983,N_26909);
xor UO_1414 (O_1414,N_29087,N_27532);
nor UO_1415 (O_1415,N_28018,N_29822);
and UO_1416 (O_1416,N_26768,N_27799);
xor UO_1417 (O_1417,N_29333,N_29353);
or UO_1418 (O_1418,N_24138,N_27276);
xnor UO_1419 (O_1419,N_26872,N_28561);
and UO_1420 (O_1420,N_28252,N_25163);
and UO_1421 (O_1421,N_26277,N_29190);
xnor UO_1422 (O_1422,N_28304,N_26542);
nand UO_1423 (O_1423,N_29496,N_29826);
and UO_1424 (O_1424,N_25618,N_27284);
xor UO_1425 (O_1425,N_26750,N_24056);
and UO_1426 (O_1426,N_27679,N_28107);
nand UO_1427 (O_1427,N_26740,N_28972);
or UO_1428 (O_1428,N_26422,N_29507);
nand UO_1429 (O_1429,N_28206,N_27591);
nor UO_1430 (O_1430,N_28348,N_28312);
or UO_1431 (O_1431,N_29605,N_29068);
nand UO_1432 (O_1432,N_25954,N_24808);
nor UO_1433 (O_1433,N_28415,N_29451);
and UO_1434 (O_1434,N_29734,N_26760);
or UO_1435 (O_1435,N_29267,N_28875);
and UO_1436 (O_1436,N_26434,N_27881);
nand UO_1437 (O_1437,N_24587,N_26401);
nor UO_1438 (O_1438,N_29849,N_26731);
nand UO_1439 (O_1439,N_28346,N_29914);
and UO_1440 (O_1440,N_26526,N_28856);
nand UO_1441 (O_1441,N_25821,N_27369);
or UO_1442 (O_1442,N_29702,N_24353);
or UO_1443 (O_1443,N_28237,N_29155);
or UO_1444 (O_1444,N_27689,N_28769);
and UO_1445 (O_1445,N_28897,N_26399);
or UO_1446 (O_1446,N_28577,N_29552);
xnor UO_1447 (O_1447,N_29809,N_24549);
nand UO_1448 (O_1448,N_24919,N_26800);
nor UO_1449 (O_1449,N_25127,N_27644);
or UO_1450 (O_1450,N_28984,N_25247);
nor UO_1451 (O_1451,N_27726,N_25924);
nor UO_1452 (O_1452,N_28516,N_24234);
nor UO_1453 (O_1453,N_29586,N_24214);
and UO_1454 (O_1454,N_24085,N_27991);
and UO_1455 (O_1455,N_26847,N_26821);
nand UO_1456 (O_1456,N_28717,N_24016);
nand UO_1457 (O_1457,N_29269,N_26237);
nor UO_1458 (O_1458,N_29699,N_26772);
nand UO_1459 (O_1459,N_24435,N_29940);
and UO_1460 (O_1460,N_28793,N_26450);
xor UO_1461 (O_1461,N_28775,N_24115);
xor UO_1462 (O_1462,N_27449,N_28411);
nand UO_1463 (O_1463,N_27200,N_24209);
xor UO_1464 (O_1464,N_26433,N_25727);
or UO_1465 (O_1465,N_24376,N_24390);
nand UO_1466 (O_1466,N_29874,N_25107);
nor UO_1467 (O_1467,N_28592,N_25773);
xnor UO_1468 (O_1468,N_25259,N_29000);
nor UO_1469 (O_1469,N_29894,N_28264);
xnor UO_1470 (O_1470,N_26147,N_25111);
xor UO_1471 (O_1471,N_25450,N_29345);
and UO_1472 (O_1472,N_26829,N_27671);
nor UO_1473 (O_1473,N_28622,N_24718);
nand UO_1474 (O_1474,N_27068,N_27850);
xnor UO_1475 (O_1475,N_28285,N_29983);
and UO_1476 (O_1476,N_27013,N_27251);
and UO_1477 (O_1477,N_27524,N_28203);
xor UO_1478 (O_1478,N_29969,N_27815);
nand UO_1479 (O_1479,N_24557,N_26988);
xor UO_1480 (O_1480,N_29074,N_29300);
xor UO_1481 (O_1481,N_25368,N_24298);
nand UO_1482 (O_1482,N_24660,N_28558);
xnor UO_1483 (O_1483,N_27359,N_26026);
or UO_1484 (O_1484,N_29790,N_28530);
and UO_1485 (O_1485,N_24224,N_25428);
xnor UO_1486 (O_1486,N_25794,N_29508);
or UO_1487 (O_1487,N_27277,N_27265);
xnor UO_1488 (O_1488,N_24694,N_25444);
nand UO_1489 (O_1489,N_29183,N_24028);
nor UO_1490 (O_1490,N_25975,N_27125);
nor UO_1491 (O_1491,N_24480,N_27809);
and UO_1492 (O_1492,N_27653,N_25999);
or UO_1493 (O_1493,N_29805,N_26977);
or UO_1494 (O_1494,N_25564,N_27953);
xnor UO_1495 (O_1495,N_25170,N_25015);
nand UO_1496 (O_1496,N_28671,N_28899);
nor UO_1497 (O_1497,N_24976,N_25706);
and UO_1498 (O_1498,N_27351,N_28678);
or UO_1499 (O_1499,N_28050,N_29597);
nand UO_1500 (O_1500,N_29617,N_24805);
and UO_1501 (O_1501,N_24548,N_27219);
and UO_1502 (O_1502,N_29436,N_26781);
or UO_1503 (O_1503,N_25723,N_25210);
nand UO_1504 (O_1504,N_24456,N_27267);
nand UO_1505 (O_1505,N_24558,N_24513);
or UO_1506 (O_1506,N_28339,N_26807);
or UO_1507 (O_1507,N_25763,N_24813);
nand UO_1508 (O_1508,N_24189,N_28970);
nor UO_1509 (O_1509,N_24585,N_24765);
nor UO_1510 (O_1510,N_26888,N_25429);
xor UO_1511 (O_1511,N_25097,N_26367);
or UO_1512 (O_1512,N_27816,N_24186);
and UO_1513 (O_1513,N_24635,N_29409);
xor UO_1514 (O_1514,N_25876,N_24669);
nor UO_1515 (O_1515,N_25585,N_25489);
xor UO_1516 (O_1516,N_29462,N_24944);
xor UO_1517 (O_1517,N_26524,N_25966);
xor UO_1518 (O_1518,N_28152,N_24790);
and UO_1519 (O_1519,N_25641,N_29835);
nor UO_1520 (O_1520,N_27875,N_27485);
or UO_1521 (O_1521,N_26929,N_28570);
and UO_1522 (O_1522,N_26468,N_29732);
or UO_1523 (O_1523,N_29846,N_24042);
and UO_1524 (O_1524,N_24824,N_27560);
nor UO_1525 (O_1525,N_25532,N_25288);
and UO_1526 (O_1526,N_29244,N_28216);
nand UO_1527 (O_1527,N_27154,N_28549);
or UO_1528 (O_1528,N_26539,N_27052);
nor UO_1529 (O_1529,N_29523,N_26202);
xor UO_1530 (O_1530,N_26140,N_25952);
xor UO_1531 (O_1531,N_29864,N_25017);
or UO_1532 (O_1532,N_24005,N_27908);
or UO_1533 (O_1533,N_28545,N_25205);
and UO_1534 (O_1534,N_29343,N_24163);
xor UO_1535 (O_1535,N_25498,N_27044);
or UO_1536 (O_1536,N_24847,N_26591);
or UO_1537 (O_1537,N_28012,N_29077);
nand UO_1538 (O_1538,N_24352,N_25976);
and UO_1539 (O_1539,N_27673,N_28440);
nand UO_1540 (O_1540,N_28378,N_27358);
xor UO_1541 (O_1541,N_26084,N_29401);
or UO_1542 (O_1542,N_25528,N_24971);
nand UO_1543 (O_1543,N_25536,N_26323);
or UO_1544 (O_1544,N_28542,N_26485);
nor UO_1545 (O_1545,N_25077,N_28580);
and UO_1546 (O_1546,N_24231,N_24881);
and UO_1547 (O_1547,N_26884,N_28033);
nor UO_1548 (O_1548,N_28398,N_27266);
nor UO_1549 (O_1549,N_28412,N_28811);
nand UO_1550 (O_1550,N_28048,N_24379);
nor UO_1551 (O_1551,N_24756,N_25813);
or UO_1552 (O_1552,N_28515,N_29640);
nor UO_1553 (O_1553,N_25915,N_27375);
and UO_1554 (O_1554,N_28952,N_28380);
nand UO_1555 (O_1555,N_26669,N_27308);
or UO_1556 (O_1556,N_26975,N_27295);
xnor UO_1557 (O_1557,N_24685,N_27870);
and UO_1558 (O_1558,N_26637,N_24580);
xnor UO_1559 (O_1559,N_24988,N_28114);
or UO_1560 (O_1560,N_28809,N_28220);
and UO_1561 (O_1561,N_29986,N_26554);
nand UO_1562 (O_1562,N_29796,N_28951);
nand UO_1563 (O_1563,N_26878,N_29777);
xnor UO_1564 (O_1564,N_25754,N_25408);
nand UO_1565 (O_1565,N_25086,N_24661);
and UO_1566 (O_1566,N_29319,N_25648);
and UO_1567 (O_1567,N_29341,N_27904);
nand UO_1568 (O_1568,N_28720,N_29317);
and UO_1569 (O_1569,N_24830,N_25388);
nor UO_1570 (O_1570,N_28565,N_27141);
nor UO_1571 (O_1571,N_28053,N_25216);
xor UO_1572 (O_1572,N_26973,N_25261);
and UO_1573 (O_1573,N_25186,N_26682);
and UO_1574 (O_1574,N_24414,N_28977);
or UO_1575 (O_1575,N_28550,N_28087);
nor UO_1576 (O_1576,N_28126,N_25358);
nor UO_1577 (O_1577,N_26461,N_29273);
nor UO_1578 (O_1578,N_26315,N_25319);
nand UO_1579 (O_1579,N_29322,N_28805);
and UO_1580 (O_1580,N_25745,N_26863);
and UO_1581 (O_1581,N_28120,N_26308);
or UO_1582 (O_1582,N_26082,N_25413);
xnor UO_1583 (O_1583,N_28613,N_27153);
and UO_1584 (O_1584,N_29498,N_25867);
nor UO_1585 (O_1585,N_27394,N_27542);
xnor UO_1586 (O_1586,N_26374,N_25352);
xnor UO_1587 (O_1587,N_28392,N_25574);
and UO_1588 (O_1588,N_26458,N_27317);
nand UO_1589 (O_1589,N_24556,N_29033);
and UO_1590 (O_1590,N_28766,N_28873);
and UO_1591 (O_1591,N_28202,N_25441);
xnor UO_1592 (O_1592,N_29562,N_24846);
and UO_1593 (O_1593,N_29313,N_25579);
or UO_1594 (O_1594,N_28133,N_24310);
nor UO_1595 (O_1595,N_27836,N_29232);
nand UO_1596 (O_1596,N_27204,N_29527);
xor UO_1597 (O_1597,N_28357,N_26725);
and UO_1598 (O_1598,N_24357,N_25295);
nand UO_1599 (O_1599,N_27134,N_26726);
nor UO_1600 (O_1600,N_24040,N_25142);
and UO_1601 (O_1601,N_26560,N_24505);
nand UO_1602 (O_1602,N_25212,N_26880);
and UO_1603 (O_1603,N_25740,N_26891);
nand UO_1604 (O_1604,N_25094,N_24825);
nor UO_1605 (O_1605,N_25483,N_26530);
nand UO_1606 (O_1606,N_28185,N_28286);
xor UO_1607 (O_1607,N_25647,N_28354);
nor UO_1608 (O_1608,N_28162,N_25356);
xnor UO_1609 (O_1609,N_25058,N_25869);
or UO_1610 (O_1610,N_24677,N_28619);
nand UO_1611 (O_1611,N_25405,N_26185);
nor UO_1612 (O_1612,N_24717,N_27372);
nor UO_1613 (O_1613,N_28892,N_24445);
nor UO_1614 (O_1614,N_27448,N_27218);
and UO_1615 (O_1615,N_29682,N_29072);
xnor UO_1616 (O_1616,N_29618,N_29588);
nand UO_1617 (O_1617,N_26331,N_29124);
or UO_1618 (O_1618,N_26405,N_29500);
xor UO_1619 (O_1619,N_29802,N_29282);
nor UO_1620 (O_1620,N_27195,N_25294);
and UO_1621 (O_1621,N_25350,N_26814);
and UO_1622 (O_1622,N_26394,N_28923);
xor UO_1623 (O_1623,N_28236,N_28395);
nand UO_1624 (O_1624,N_25870,N_27494);
nor UO_1625 (O_1625,N_26285,N_28066);
or UO_1626 (O_1626,N_27272,N_27543);
nor UO_1627 (O_1627,N_25181,N_28888);
nand UO_1628 (O_1628,N_26652,N_26600);
and UO_1629 (O_1629,N_24654,N_29156);
xnor UO_1630 (O_1630,N_28902,N_29355);
or UO_1631 (O_1631,N_27713,N_25119);
nor UO_1632 (O_1632,N_28055,N_29497);
xnor UO_1633 (O_1633,N_29612,N_26924);
nand UO_1634 (O_1634,N_25739,N_27597);
nand UO_1635 (O_1635,N_25682,N_28455);
and UO_1636 (O_1636,N_29207,N_27892);
or UO_1637 (O_1637,N_26154,N_28864);
or UO_1638 (O_1638,N_28222,N_26564);
or UO_1639 (O_1639,N_29757,N_24380);
or UO_1640 (O_1640,N_25515,N_27744);
and UO_1641 (O_1641,N_29651,N_24455);
nand UO_1642 (O_1642,N_24563,N_29906);
xor UO_1643 (O_1643,N_27350,N_28648);
xor UO_1644 (O_1644,N_24064,N_27757);
or UO_1645 (O_1645,N_29698,N_25165);
nor UO_1646 (O_1646,N_27918,N_26074);
nand UO_1647 (O_1647,N_25730,N_27925);
and UO_1648 (O_1648,N_29344,N_28531);
and UO_1649 (O_1649,N_29635,N_27868);
nor UO_1650 (O_1650,N_28049,N_27160);
xor UO_1651 (O_1651,N_24417,N_29539);
or UO_1652 (O_1652,N_27835,N_24945);
xor UO_1653 (O_1653,N_24388,N_28160);
and UO_1654 (O_1654,N_24930,N_27413);
nor UO_1655 (O_1655,N_25480,N_24343);
or UO_1656 (O_1656,N_24924,N_26985);
nand UO_1657 (O_1657,N_25372,N_26012);
xor UO_1658 (O_1658,N_24738,N_25680);
nand UO_1659 (O_1659,N_27948,N_29318);
or UO_1660 (O_1660,N_26211,N_28396);
or UO_1661 (O_1661,N_27456,N_28165);
nand UO_1662 (O_1662,N_28360,N_29898);
nor UO_1663 (O_1663,N_24377,N_26679);
or UO_1664 (O_1664,N_26491,N_26575);
xnor UO_1665 (O_1665,N_29425,N_27964);
nor UO_1666 (O_1666,N_25436,N_25148);
xnor UO_1667 (O_1667,N_26594,N_28881);
or UO_1668 (O_1668,N_28376,N_26738);
nand UO_1669 (O_1669,N_28250,N_26968);
or UO_1670 (O_1670,N_28901,N_26459);
nand UO_1671 (O_1671,N_25725,N_29296);
xnor UO_1672 (O_1672,N_25746,N_24257);
nand UO_1673 (O_1673,N_26445,N_24296);
nand UO_1674 (O_1674,N_29825,N_26296);
or UO_1675 (O_1675,N_27268,N_28712);
nor UO_1676 (O_1676,N_27784,N_28768);
nor UO_1677 (O_1677,N_26918,N_24844);
or UO_1678 (O_1678,N_24884,N_29560);
xor UO_1679 (O_1679,N_28108,N_25908);
nor UO_1680 (O_1680,N_28386,N_27551);
nor UO_1681 (O_1681,N_27051,N_26462);
xor UO_1682 (O_1682,N_24207,N_27538);
xnor UO_1683 (O_1683,N_29689,N_28588);
nand UO_1684 (O_1684,N_24155,N_28028);
and UO_1685 (O_1685,N_27457,N_26408);
xor UO_1686 (O_1686,N_24144,N_28261);
or UO_1687 (O_1687,N_26068,N_29350);
and UO_1688 (O_1688,N_28914,N_29581);
nor UO_1689 (O_1689,N_25850,N_25941);
or UO_1690 (O_1690,N_29138,N_28936);
or UO_1691 (O_1691,N_28539,N_24671);
and UO_1692 (O_1692,N_25788,N_25136);
nor UO_1693 (O_1693,N_24527,N_27385);
or UO_1694 (O_1694,N_26705,N_25354);
xor UO_1695 (O_1695,N_26028,N_27749);
xnor UO_1696 (O_1696,N_27621,N_24998);
and UO_1697 (O_1697,N_24321,N_27063);
or UO_1698 (O_1698,N_25700,N_28679);
xor UO_1699 (O_1699,N_24981,N_29761);
or UO_1700 (O_1700,N_29356,N_24317);
nand UO_1701 (O_1701,N_26749,N_26522);
nor UO_1702 (O_1702,N_27198,N_28167);
xor UO_1703 (O_1703,N_26877,N_27012);
or UO_1704 (O_1704,N_25399,N_26156);
or UO_1705 (O_1705,N_27139,N_26833);
or UO_1706 (O_1706,N_28153,N_28223);
nand UO_1707 (O_1707,N_25874,N_27025);
or UO_1708 (O_1708,N_26443,N_28544);
and UO_1709 (O_1709,N_26963,N_29623);
and UO_1710 (O_1710,N_29080,N_26883);
and UO_1711 (O_1711,N_27230,N_27851);
nor UO_1712 (O_1712,N_28538,N_25683);
nand UO_1713 (O_1713,N_24429,N_25774);
nand UO_1714 (O_1714,N_26400,N_27168);
nand UO_1715 (O_1715,N_29505,N_25795);
xor UO_1716 (O_1716,N_28256,N_25786);
or UO_1717 (O_1717,N_29154,N_26079);
nand UO_1718 (O_1718,N_29976,N_26190);
and UO_1719 (O_1719,N_24021,N_26325);
xnor UO_1720 (O_1720,N_26196,N_24617);
or UO_1721 (O_1721,N_25665,N_29896);
or UO_1722 (O_1722,N_28435,N_29302);
or UO_1723 (O_1723,N_29284,N_24901);
or UO_1724 (O_1724,N_29975,N_25553);
xnor UO_1725 (O_1725,N_24668,N_28292);
and UO_1726 (O_1726,N_28344,N_26649);
xor UO_1727 (O_1727,N_25122,N_24895);
and UO_1728 (O_1728,N_25549,N_29681);
and UO_1729 (O_1729,N_29454,N_25637);
or UO_1730 (O_1730,N_27801,N_26845);
nand UO_1731 (O_1731,N_27281,N_27986);
or UO_1732 (O_1732,N_24646,N_25797);
nor UO_1733 (O_1733,N_25695,N_29720);
xor UO_1734 (O_1734,N_25857,N_26681);
or UO_1735 (O_1735,N_26247,N_29339);
xnor UO_1736 (O_1736,N_29472,N_25013);
and UO_1737 (O_1737,N_25778,N_28465);
nand UO_1738 (O_1738,N_26816,N_26930);
xor UO_1739 (O_1739,N_27972,N_24639);
nand UO_1740 (O_1740,N_25391,N_26967);
nand UO_1741 (O_1741,N_28326,N_26802);
or UO_1742 (O_1742,N_26955,N_26182);
nor UO_1743 (O_1743,N_26288,N_28255);
xor UO_1744 (O_1744,N_24101,N_25423);
nor UO_1745 (O_1745,N_27615,N_25846);
nor UO_1746 (O_1746,N_24476,N_29775);
and UO_1747 (O_1747,N_28557,N_28937);
or UO_1748 (O_1748,N_28218,N_29211);
nand UO_1749 (O_1749,N_26860,N_25626);
xnor UO_1750 (O_1750,N_24084,N_27566);
and UO_1751 (O_1751,N_28313,N_27158);
xnor UO_1752 (O_1752,N_28845,N_26902);
xor UO_1753 (O_1753,N_26801,N_25095);
or UO_1754 (O_1754,N_26935,N_26759);
nor UO_1755 (O_1755,N_26854,N_26830);
xnor UO_1756 (O_1756,N_29545,N_26886);
or UO_1757 (O_1757,N_27787,N_29463);
nor UO_1758 (O_1758,N_28113,N_28791);
or UO_1759 (O_1759,N_26966,N_26292);
nand UO_1760 (O_1760,N_28525,N_26117);
xor UO_1761 (O_1761,N_25702,N_27409);
nand UO_1762 (O_1762,N_26381,N_26370);
nor UO_1763 (O_1763,N_25341,N_25735);
nor UO_1764 (O_1764,N_27213,N_24726);
nor UO_1765 (O_1765,N_24485,N_26449);
or UO_1766 (O_1766,N_26166,N_29128);
and UO_1767 (O_1767,N_27432,N_24748);
or UO_1768 (O_1768,N_27884,N_24133);
and UO_1769 (O_1769,N_25135,N_24823);
nand UO_1770 (O_1770,N_29253,N_27117);
nor UO_1771 (O_1771,N_24059,N_25790);
or UO_1772 (O_1772,N_27469,N_25670);
or UO_1773 (O_1773,N_28957,N_28989);
and UO_1774 (O_1774,N_27583,N_29963);
nor UO_1775 (O_1775,N_29626,N_29866);
xnor UO_1776 (O_1776,N_28879,N_25418);
nand UO_1777 (O_1777,N_28926,N_28681);
nor UO_1778 (O_1778,N_26169,N_24258);
and UO_1779 (O_1779,N_27441,N_27119);
and UO_1780 (O_1780,N_26105,N_29919);
and UO_1781 (O_1781,N_26446,N_26785);
or UO_1782 (O_1782,N_27706,N_27293);
xnor UO_1783 (O_1783,N_29967,N_27938);
and UO_1784 (O_1784,N_28644,N_24665);
nand UO_1785 (O_1785,N_27825,N_26840);
xnor UO_1786 (O_1786,N_25983,N_26876);
nor UO_1787 (O_1787,N_24341,N_26555);
nor UO_1788 (O_1788,N_27710,N_28586);
nor UO_1789 (O_1789,N_25024,N_26149);
nor UO_1790 (O_1790,N_28560,N_27927);
xnor UO_1791 (O_1791,N_24812,N_26113);
or UO_1792 (O_1792,N_26870,N_24137);
nor UO_1793 (O_1793,N_24235,N_29920);
or UO_1794 (O_1794,N_25720,N_28707);
nand UO_1795 (O_1795,N_26791,N_29767);
and UO_1796 (O_1796,N_27549,N_27434);
xnor UO_1797 (O_1797,N_29208,N_24143);
nor UO_1798 (O_1798,N_24404,N_24821);
nor UO_1799 (O_1799,N_25894,N_28235);
or UO_1800 (O_1800,N_25289,N_25847);
and UO_1801 (O_1801,N_26852,N_26941);
or UO_1802 (O_1802,N_25440,N_24266);
nor UO_1803 (O_1803,N_27982,N_27133);
nand UO_1804 (O_1804,N_25257,N_24902);
xor UO_1805 (O_1805,N_27211,N_27588);
or UO_1806 (O_1806,N_24122,N_27989);
nand UO_1807 (O_1807,N_24440,N_29040);
nor UO_1808 (O_1808,N_27693,N_26195);
and UO_1809 (O_1809,N_24291,N_29834);
nor UO_1810 (O_1810,N_27831,N_24964);
nand UO_1811 (O_1811,N_28136,N_27516);
xnor UO_1812 (O_1812,N_27535,N_27071);
or UO_1813 (O_1813,N_25200,N_28669);
nand UO_1814 (O_1814,N_28541,N_27924);
nor UO_1815 (O_1815,N_25256,N_28974);
nor UO_1816 (O_1816,N_25296,N_29299);
nand UO_1817 (O_1817,N_24693,N_28129);
nor UO_1818 (O_1818,N_24682,N_28039);
nor UO_1819 (O_1819,N_27425,N_27765);
nand UO_1820 (O_1820,N_25777,N_25452);
or UO_1821 (O_1821,N_24650,N_29188);
xnor UO_1822 (O_1822,N_27572,N_25971);
nand UO_1823 (O_1823,N_29373,N_29915);
nand UO_1824 (O_1824,N_24774,N_25775);
and UO_1825 (O_1825,N_29027,N_24560);
and UO_1826 (O_1826,N_27681,N_29926);
nand UO_1827 (O_1827,N_24935,N_24108);
or UO_1828 (O_1828,N_25204,N_25169);
nor UO_1829 (O_1829,N_27620,N_27216);
xor UO_1830 (O_1830,N_29793,N_27797);
or UO_1831 (O_1831,N_25674,N_26754);
or UO_1832 (O_1832,N_28568,N_25996);
nand UO_1833 (O_1833,N_27289,N_25506);
and UO_1834 (O_1834,N_25056,N_27937);
nor UO_1835 (O_1835,N_26419,N_27920);
xor UO_1836 (O_1836,N_29178,N_27607);
or UO_1837 (O_1837,N_27783,N_29433);
nand UO_1838 (O_1838,N_29780,N_24552);
nor UO_1839 (O_1839,N_29900,N_24323);
or UO_1840 (O_1840,N_25742,N_29161);
nand UO_1841 (O_1841,N_28449,N_29110);
and UO_1842 (O_1842,N_26869,N_28243);
or UO_1843 (O_1843,N_29331,N_26358);
nor UO_1844 (O_1844,N_28733,N_29948);
nand UO_1845 (O_1845,N_27235,N_25232);
nand UO_1846 (O_1846,N_29960,N_28479);
and UO_1847 (O_1847,N_28476,N_24754);
nand UO_1848 (O_1848,N_27163,N_25494);
and UO_1849 (O_1849,N_28281,N_24470);
xor UO_1850 (O_1850,N_29499,N_28075);
nand UO_1851 (O_1851,N_24798,N_26626);
and UO_1852 (O_1852,N_26116,N_26998);
or UO_1853 (O_1853,N_26634,N_24098);
xor UO_1854 (O_1854,N_26219,N_26120);
and UO_1855 (O_1855,N_27426,N_25864);
and UO_1856 (O_1856,N_29708,N_24043);
and UO_1857 (O_1857,N_29399,N_29256);
and UO_1858 (O_1858,N_24571,N_27968);
nand UO_1859 (O_1859,N_24154,N_25430);
xnor UO_1860 (O_1860,N_24806,N_24271);
and UO_1861 (O_1861,N_29004,N_25487);
xnor UO_1862 (O_1862,N_29439,N_26543);
or UO_1863 (O_1863,N_26192,N_25236);
or UO_1864 (O_1864,N_29320,N_28383);
nand UO_1865 (O_1865,N_28925,N_29235);
nand UO_1866 (O_1866,N_28061,N_28887);
or UO_1867 (O_1867,N_28481,N_26300);
nand UO_1868 (O_1868,N_24686,N_25751);
and UO_1869 (O_1869,N_26122,N_28090);
xor UO_1870 (O_1870,N_28526,N_26597);
nor UO_1871 (O_1871,N_28418,N_26376);
nand UO_1872 (O_1872,N_26804,N_24683);
xnor UO_1873 (O_1873,N_25887,N_28820);
xor UO_1874 (O_1874,N_25688,N_25014);
or UO_1875 (O_1875,N_27718,N_29086);
and UO_1876 (O_1876,N_27692,N_27902);
nor UO_1877 (O_1877,N_26085,N_27833);
nand UO_1878 (O_1878,N_28232,N_26334);
xor UO_1879 (O_1879,N_25715,N_24607);
nor UO_1880 (O_1880,N_26457,N_24221);
nor UO_1881 (O_1881,N_26121,N_25537);
xor UO_1882 (O_1882,N_28363,N_27678);
or UO_1883 (O_1883,N_29460,N_25005);
xor UO_1884 (O_1884,N_25696,N_24666);
and UO_1885 (O_1885,N_26509,N_29297);
or UO_1886 (O_1886,N_25269,N_25878);
or UO_1887 (O_1887,N_29391,N_27336);
xor UO_1888 (O_1888,N_25191,N_26206);
xor UO_1889 (O_1889,N_29519,N_28019);
nand UO_1890 (O_1890,N_29298,N_25367);
nand UO_1891 (O_1891,N_24799,N_28274);
xor UO_1892 (O_1892,N_24664,N_25984);
xnor UO_1893 (O_1893,N_28891,N_29921);
or UO_1894 (O_1894,N_24550,N_27167);
or UO_1895 (O_1895,N_27464,N_24095);
or UO_1896 (O_1896,N_25921,N_25253);
and UO_1897 (O_1897,N_25335,N_29878);
nor UO_1898 (O_1898,N_27508,N_26672);
nand UO_1899 (O_1899,N_29290,N_26717);
nor UO_1900 (O_1900,N_28626,N_27504);
nor UO_1901 (O_1901,N_27728,N_26787);
xor UO_1902 (O_1902,N_26053,N_24780);
and UO_1903 (O_1903,N_27598,N_28794);
nand UO_1904 (O_1904,N_25237,N_29082);
xor UO_1905 (O_1905,N_26246,N_29526);
and UO_1906 (O_1906,N_26250,N_26783);
nor UO_1907 (O_1907,N_28852,N_26371);
or UO_1908 (O_1908,N_27354,N_25241);
or UO_1909 (O_1909,N_24146,N_29511);
nand UO_1910 (O_1910,N_28513,N_24835);
xor UO_1911 (O_1911,N_25923,N_24731);
nand UO_1912 (O_1912,N_27685,N_26207);
and UO_1913 (O_1913,N_27095,N_26517);
nor UO_1914 (O_1914,N_24502,N_25138);
nand UO_1915 (O_1915,N_26568,N_27869);
or UO_1916 (O_1916,N_29036,N_29272);
and UO_1917 (O_1917,N_27792,N_24878);
xnor UO_1918 (O_1918,N_29938,N_27118);
or UO_1919 (O_1919,N_29503,N_24526);
nor UO_1920 (O_1920,N_29509,N_25411);
and UO_1921 (O_1921,N_24181,N_29961);
nand UO_1922 (O_1922,N_28369,N_27978);
nand UO_1923 (O_1923,N_28078,N_28192);
nand UO_1924 (O_1924,N_29090,N_27619);
or UO_1925 (O_1925,N_26152,N_28885);
or UO_1926 (O_1926,N_26714,N_26989);
xor UO_1927 (O_1927,N_27973,N_24862);
nor UO_1928 (O_1928,N_26018,N_29417);
xor UO_1929 (O_1929,N_27170,N_27047);
or UO_1930 (O_1930,N_24281,N_26027);
nand UO_1931 (O_1931,N_24760,N_26005);
nand UO_1932 (O_1932,N_25973,N_24684);
xnor UO_1933 (O_1933,N_29167,N_24855);
or UO_1934 (O_1934,N_28027,N_29818);
xnor UO_1935 (O_1935,N_26866,N_28691);
or UO_1936 (O_1936,N_26619,N_26532);
or UO_1937 (O_1937,N_27435,N_28051);
xnor UO_1938 (O_1938,N_27323,N_29219);
nor UO_1939 (O_1939,N_26181,N_29108);
nor UO_1940 (O_1940,N_27843,N_25065);
or UO_1941 (O_1941,N_25892,N_26937);
nand UO_1942 (O_1942,N_28838,N_24936);
and UO_1943 (O_1943,N_26729,N_28260);
xnor UO_1944 (O_1944,N_24111,N_28008);
nor UO_1945 (O_1945,N_24999,N_25465);
nor UO_1946 (O_1946,N_28381,N_25518);
and UO_1947 (O_1947,N_29204,N_28559);
and UO_1948 (O_1948,N_27567,N_25496);
xor UO_1949 (O_1949,N_28660,N_24011);
nor UO_1950 (O_1950,N_27349,N_28382);
nand UO_1951 (O_1951,N_28621,N_27633);
nand UO_1952 (O_1952,N_29936,N_28753);
nand UO_1953 (O_1953,N_24333,N_25711);
nand UO_1954 (O_1954,N_27006,N_27156);
nand UO_1955 (O_1955,N_26088,N_29937);
nand UO_1956 (O_1956,N_28106,N_25832);
or UO_1957 (O_1957,N_26472,N_29525);
xor UO_1958 (O_1958,N_26306,N_29276);
or UO_1959 (O_1959,N_28445,N_29630);
and UO_1960 (O_1960,N_24649,N_26397);
and UO_1961 (O_1961,N_28248,N_25731);
nor UO_1962 (O_1962,N_29259,N_25310);
xnor UO_1963 (O_1963,N_24276,N_28399);
and UO_1964 (O_1964,N_28682,N_25733);
or UO_1965 (O_1965,N_27074,N_24000);
nand UO_1966 (O_1966,N_28373,N_29547);
nand UO_1967 (O_1967,N_27916,N_24491);
nor UO_1968 (O_1968,N_28466,N_28020);
nor UO_1969 (O_1969,N_25570,N_26236);
nand UO_1970 (O_1970,N_24689,N_24432);
and UO_1971 (O_1971,N_24540,N_25703);
xor UO_1972 (O_1972,N_28597,N_28233);
nand UO_1973 (O_1973,N_29744,N_28724);
nor UO_1974 (O_1974,N_25157,N_28495);
xnor UO_1975 (O_1975,N_27474,N_25960);
xor UO_1976 (O_1976,N_24348,N_24833);
nor UO_1977 (O_1977,N_24865,N_25889);
xor UO_1978 (O_1978,N_26388,N_24242);
xnor UO_1979 (O_1979,N_29529,N_24963);
xor UO_1980 (O_1980,N_24870,N_25137);
or UO_1981 (O_1981,N_27368,N_29127);
or UO_1982 (O_1982,N_28478,N_27450);
nand UO_1983 (O_1983,N_26225,N_29996);
and UO_1984 (O_1984,N_26890,N_24658);
or UO_1985 (O_1985,N_29895,N_25577);
xnor UO_1986 (O_1986,N_24167,N_24345);
or UO_1987 (O_1987,N_27221,N_26842);
xnor UO_1988 (O_1988,N_24253,N_26741);
and UO_1989 (O_1989,N_24330,N_29411);
xor UO_1990 (O_1990,N_25787,N_26716);
nand UO_1991 (O_1991,N_25359,N_28827);
xnor UO_1992 (O_1992,N_24992,N_24274);
nand UO_1993 (O_1993,N_27089,N_24313);
nor UO_1994 (O_1994,N_29563,N_24114);
nor UO_1995 (O_1995,N_27563,N_26773);
nor UO_1996 (O_1996,N_24006,N_26372);
nor UO_1997 (O_1997,N_24135,N_26606);
nor UO_1998 (O_1998,N_27257,N_24125);
xor UO_1999 (O_1999,N_24462,N_29855);
nor UO_2000 (O_2000,N_25258,N_25613);
xor UO_2001 (O_2001,N_29437,N_24959);
xnor UO_2002 (O_2002,N_25555,N_27189);
xnor UO_2003 (O_2003,N_29084,N_24083);
nor UO_2004 (O_2004,N_25724,N_28247);
xor UO_2005 (O_2005,N_24709,N_26212);
xnor UO_2006 (O_2006,N_29364,N_25417);
and UO_2007 (O_2007,N_27980,N_25500);
and UO_2008 (O_2008,N_28641,N_28309);
nand UO_2009 (O_2009,N_28298,N_25409);
xnor UO_2010 (O_2010,N_29883,N_25947);
nand UO_2011 (O_2011,N_26897,N_26067);
or UO_2012 (O_2012,N_24701,N_24943);
xnor UO_2013 (O_2013,N_26815,N_28277);
xnor UO_2014 (O_2014,N_26665,N_26828);
nand UO_2015 (O_2015,N_28762,N_28188);
or UO_2016 (O_2016,N_26851,N_25716);
nand UO_2017 (O_2017,N_28496,N_24966);
xor UO_2018 (O_2018,N_25671,N_26565);
nand UO_2019 (O_2019,N_25007,N_26233);
nor UO_2020 (O_2020,N_24500,N_27949);
nor UO_2021 (O_2021,N_26861,N_24792);
or UO_2022 (O_2022,N_28258,N_29265);
or UO_2023 (O_2023,N_26848,N_25008);
and UO_2024 (O_2024,N_25185,N_29501);
nor UO_2025 (O_2025,N_24721,N_25660);
or UO_2026 (O_2026,N_27228,N_26496);
xnor UO_2027 (O_2027,N_27040,N_26487);
nand UO_2028 (O_2028,N_29557,N_25726);
or UO_2029 (O_2029,N_26350,N_28494);
nor UO_2030 (O_2030,N_26621,N_26547);
and UO_2031 (O_2031,N_29125,N_24238);
nor UO_2032 (O_2032,N_24444,N_26191);
nor UO_2033 (O_2033,N_26391,N_29877);
and UO_2034 (O_2034,N_24729,N_27984);
and UO_2035 (O_2035,N_24347,N_29587);
nor UO_2036 (O_2036,N_25906,N_29275);
nor UO_2037 (O_2037,N_29291,N_28138);
nor UO_2038 (O_2038,N_28358,N_25562);
nand UO_2039 (O_2039,N_28031,N_26243);
or UO_2040 (O_2040,N_27029,N_24087);
nor UO_2041 (O_2041,N_29222,N_25046);
nor UO_2042 (O_2042,N_26044,N_25375);
or UO_2043 (O_2043,N_26666,N_24401);
xnor UO_2044 (O_2044,N_27558,N_29447);
and UO_2045 (O_2045,N_27500,N_26421);
xnor UO_2046 (O_2046,N_24908,N_25531);
nor UO_2047 (O_2047,N_28735,N_28423);
and UO_2048 (O_2048,N_27188,N_26700);
nor UO_2049 (O_2049,N_28161,N_27732);
nor UO_2050 (O_2050,N_24947,N_25750);
and UO_2051 (O_2051,N_26046,N_28062);
or UO_2052 (O_2052,N_24396,N_24739);
or UO_2053 (O_2053,N_27246,N_25180);
or UO_2054 (O_2054,N_27306,N_25986);
nor UO_2055 (O_2055,N_29962,N_27227);
nand UO_2056 (O_2056,N_27337,N_28299);
xor UO_2057 (O_2057,N_26284,N_28599);
nand UO_2058 (O_2058,N_26174,N_27439);
nand UO_2059 (O_2059,N_29621,N_26855);
xnor UO_2060 (O_2060,N_24922,N_26782);
nand UO_2061 (O_2061,N_25273,N_27652);
nor UO_2062 (O_2062,N_28591,N_28442);
nand UO_2063 (O_2063,N_24801,N_24419);
and UO_2064 (O_2064,N_25188,N_25389);
nor UO_2065 (O_2065,N_28746,N_26319);
nand UO_2066 (O_2066,N_29801,N_28540);
nor UO_2067 (O_2067,N_24679,N_27808);
xor UO_2068 (O_2068,N_26021,N_29459);
xor UO_2069 (O_2069,N_26689,N_27417);
xnor UO_2070 (O_2070,N_25336,N_27714);
nand UO_2071 (O_2071,N_26404,N_29723);
xnor UO_2072 (O_2072,N_27518,N_26483);
nor UO_2073 (O_2073,N_26969,N_28656);
and UO_2074 (O_2074,N_25139,N_29236);
nor UO_2075 (O_2075,N_24392,N_27818);
and UO_2076 (O_2076,N_28955,N_26873);
and UO_2077 (O_2077,N_26050,N_25830);
nor UO_2078 (O_2078,N_29758,N_27747);
or UO_2079 (O_2079,N_28115,N_28890);
nand UO_2080 (O_2080,N_24511,N_28425);
nor UO_2081 (O_2081,N_25473,N_28504);
and UO_2082 (O_2082,N_24910,N_24458);
xor UO_2083 (O_2083,N_26571,N_27357);
nor UO_2084 (O_2084,N_27627,N_27325);
and UO_2085 (O_2085,N_24105,N_29458);
nor UO_2086 (O_2086,N_28610,N_24109);
nor UO_2087 (O_2087,N_28187,N_28439);
xor UO_2088 (O_2088,N_26922,N_26158);
and UO_2089 (O_2089,N_24522,N_26184);
and UO_2090 (O_2090,N_28347,N_27768);
nor UO_2091 (O_2091,N_26438,N_27482);
nor UO_2092 (O_2092,N_24256,N_26615);
nor UO_2093 (O_2093,N_29610,N_24655);
or UO_2094 (O_2094,N_26365,N_24681);
or UO_2095 (O_2095,N_26797,N_26466);
or UO_2096 (O_2096,N_25664,N_26402);
xnor UO_2097 (O_2097,N_28181,N_26266);
nand UO_2098 (O_2098,N_24968,N_25083);
and UO_2099 (O_2099,N_28351,N_26822);
and UO_2100 (O_2100,N_26352,N_24771);
xnor UO_2101 (O_2101,N_24129,N_26274);
xnor UO_2102 (O_2102,N_25213,N_28265);
and UO_2103 (O_2103,N_25837,N_26518);
xnor UO_2104 (O_2104,N_26338,N_26063);
or UO_2105 (O_2105,N_24001,N_27097);
or UO_2106 (O_2106,N_26906,N_26651);
nor UO_2107 (O_2107,N_25051,N_26525);
nor UO_2108 (O_2108,N_29902,N_27853);
xnor UO_2109 (O_2109,N_29066,N_27212);
and UO_2110 (O_2110,N_24608,N_28083);
or UO_2111 (O_2111,N_26007,N_25697);
and UO_2112 (O_2112,N_29032,N_25421);
nor UO_2113 (O_2113,N_24984,N_28303);
nand UO_2114 (O_2114,N_24757,N_28728);
nand UO_2115 (O_2115,N_25606,N_27522);
nand UO_2116 (O_2116,N_24102,N_26562);
nand UO_2117 (O_2117,N_28627,N_26157);
or UO_2118 (O_2118,N_24892,N_28117);
xor UO_2119 (O_2119,N_25433,N_29095);
nor UO_2120 (O_2120,N_24304,N_29394);
or UO_2121 (O_2121,N_27318,N_25410);
and UO_2122 (O_2122,N_24201,N_29362);
nand UO_2123 (O_2123,N_26579,N_28767);
nor UO_2124 (O_2124,N_28505,N_25330);
nand UO_2125 (O_2125,N_29840,N_29424);
or UO_2126 (O_2126,N_27906,N_25315);
nor UO_2127 (O_2127,N_26379,N_26632);
and UO_2128 (O_2128,N_24934,N_24498);
nand UO_2129 (O_2129,N_29330,N_29324);
and UO_2130 (O_2130,N_28110,N_26570);
and UO_2131 (O_2131,N_28444,N_29224);
or UO_2132 (O_2132,N_26489,N_25681);
or UO_2133 (O_2133,N_24692,N_26756);
or UO_2134 (O_2134,N_24763,N_25390);
nor UO_2135 (O_2135,N_29714,N_25938);
nor UO_2136 (O_2136,N_26505,N_24478);
and UO_2137 (O_2137,N_26642,N_27465);
xor UO_2138 (O_2138,N_28350,N_28904);
and UO_2139 (O_2139,N_28080,N_26718);
and UO_2140 (O_2140,N_29434,N_25175);
xnor UO_2141 (O_2141,N_26695,N_29034);
nor UO_2142 (O_2142,N_24869,N_24013);
xnor UO_2143 (O_2143,N_26301,N_25371);
xor UO_2144 (O_2144,N_28596,N_27735);
nand UO_2145 (O_2145,N_24117,N_26100);
xnor UO_2146 (O_2146,N_28569,N_27910);
and UO_2147 (O_2147,N_27533,N_29326);
or UO_2148 (O_2148,N_29729,N_26052);
or UO_2149 (O_2149,N_26727,N_24501);
and UO_2150 (O_2150,N_28968,N_26373);
nor UO_2151 (O_2151,N_27226,N_24628);
xnor UO_2152 (O_2152,N_26294,N_27642);
nor UO_2153 (O_2153,N_28826,N_28929);
nand UO_2154 (O_2154,N_25883,N_26218);
and UO_2155 (O_2155,N_27624,N_24208);
xor UO_2156 (O_2156,N_26463,N_25059);
xnor UO_2157 (O_2157,N_27100,N_28468);
nand UO_2158 (O_2158,N_24072,N_28673);
or UO_2159 (O_2159,N_25266,N_24044);
and UO_2160 (O_2160,N_27042,N_24228);
nand UO_2161 (O_2161,N_26229,N_28489);
nand UO_2162 (O_2162,N_27244,N_25514);
nor UO_2163 (O_2163,N_27345,N_26915);
nand UO_2164 (O_2164,N_25145,N_25810);
and UO_2165 (O_2165,N_28131,N_27489);
and UO_2166 (O_2166,N_26329,N_24290);
nor UO_2167 (O_2167,N_26008,N_27241);
and UO_2168 (O_2168,N_29510,N_25347);
or UO_2169 (O_2169,N_29001,N_29168);
xor UO_2170 (O_2170,N_28148,N_24575);
xor UO_2171 (O_2171,N_26194,N_28302);
nand UO_2172 (O_2172,N_25193,N_27630);
or UO_2173 (O_2173,N_26770,N_27570);
nand UO_2174 (O_2174,N_24494,N_29671);
or UO_2175 (O_2175,N_28985,N_24403);
or UO_2176 (O_2176,N_27832,N_25509);
nand UO_2177 (O_2177,N_29149,N_27683);
nor UO_2178 (O_2178,N_29075,N_25195);
and UO_2179 (O_2179,N_28666,N_28792);
or UO_2180 (O_2180,N_28172,N_25873);
nand UO_2181 (O_2181,N_24903,N_28319);
xnor UO_2182 (O_2182,N_28385,N_24623);
nor UO_2183 (O_2183,N_24516,N_24586);
or UO_2184 (O_2184,N_29098,N_29421);
and UO_2185 (O_2185,N_25965,N_27912);
and UO_2186 (O_2186,N_26980,N_25566);
nor UO_2187 (O_2187,N_29376,N_29088);
nand UO_2188 (O_2188,N_27020,N_28713);
nand UO_2189 (O_2189,N_26407,N_27496);
nor UO_2190 (O_2190,N_26151,N_25845);
or UO_2191 (O_2191,N_28908,N_29800);
nand UO_2192 (O_2192,N_27819,N_29669);
or UO_2193 (O_2193,N_29856,N_27194);
nand UO_2194 (O_2194,N_29567,N_29293);
and UO_2195 (O_2195,N_24569,N_28437);
and UO_2196 (O_2196,N_29572,N_24640);
nor UO_2197 (O_2197,N_27677,N_27754);
xor UO_2198 (O_2198,N_28035,N_25485);
xor UO_2199 (O_2199,N_26042,N_28144);
nor UO_2200 (O_2200,N_26585,N_28278);
nor UO_2201 (O_2201,N_26576,N_24632);
nor UO_2202 (O_2202,N_24239,N_24340);
nand UO_2203 (O_2203,N_29470,N_29408);
nor UO_2204 (O_2204,N_24066,N_26208);
xnor UO_2205 (O_2205,N_25928,N_24441);
nor UO_2206 (O_2206,N_28556,N_27233);
xor UO_2207 (O_2207,N_26230,N_24320);
nand UO_2208 (O_2208,N_29308,N_28860);
xnor UO_2209 (O_2209,N_27416,N_28414);
xor UO_2210 (O_2210,N_29484,N_26291);
nand UO_2211 (O_2211,N_27688,N_29145);
nor UO_2212 (O_2212,N_29806,N_28601);
and UO_2213 (O_2213,N_29419,N_29832);
xor UO_2214 (O_2214,N_25303,N_24695);
or UO_2215 (O_2215,N_24572,N_26599);
or UO_2216 (O_2216,N_25534,N_24436);
or UO_2217 (O_2217,N_27408,N_25783);
xor UO_2218 (O_2218,N_26850,N_28837);
xnor UO_2219 (O_2219,N_28081,N_28177);
or UO_2220 (O_2220,N_26076,N_29703);
xnor UO_2221 (O_2221,N_26728,N_29277);
and UO_2222 (O_2222,N_25563,N_24278);
and UO_2223 (O_2223,N_28128,N_24481);
xnor UO_2224 (O_2224,N_24191,N_28361);
nor UO_2225 (O_2225,N_24820,N_27036);
nand UO_2226 (O_2226,N_25147,N_24657);
or UO_2227 (O_2227,N_29094,N_28393);
nor UO_2228 (O_2228,N_25403,N_24264);
or UO_2229 (O_2229,N_26622,N_26321);
xnor UO_2230 (O_2230,N_29683,N_26896);
nor UO_2231 (O_2231,N_29974,N_25580);
nand UO_2232 (O_2232,N_26769,N_25587);
or UO_2233 (O_2233,N_29328,N_24179);
xor UO_2234 (O_2234,N_26551,N_24204);
nand UO_2235 (O_2235,N_24421,N_26197);
nor UO_2236 (O_2236,N_28210,N_25594);
xor UO_2237 (O_2237,N_26263,N_29949);
nor UO_2238 (O_2238,N_26344,N_26265);
xor UO_2239 (O_2239,N_25554,N_26411);
xnor UO_2240 (O_2240,N_27663,N_27130);
nand UO_2241 (O_2241,N_29663,N_25831);
nor UO_2242 (O_2242,N_28463,N_26646);
nand UO_2243 (O_2243,N_28057,N_24882);
nor UO_2244 (O_2244,N_26141,N_24240);
xnor UO_2245 (O_2245,N_26721,N_24633);
and UO_2246 (O_2246,N_27237,N_25978);
nand UO_2247 (O_2247,N_28199,N_26660);
xnor UO_2248 (O_2248,N_25184,N_26170);
xor UO_2249 (O_2249,N_24890,N_27057);
xor UO_2250 (O_2250,N_25276,N_29627);
and UO_2251 (O_2251,N_26910,N_27490);
and UO_2252 (O_2252,N_29254,N_24641);
and UO_2253 (O_2253,N_27466,N_28464);
and UO_2254 (O_2254,N_24058,N_28818);
nor UO_2255 (O_2255,N_25633,N_25123);
and UO_2256 (O_2256,N_27696,N_25793);
xnor UO_2257 (O_2257,N_24314,N_26820);
xnor UO_2258 (O_2258,N_24993,N_25612);
or UO_2259 (O_2259,N_26914,N_24169);
nand UO_2260 (O_2260,N_28005,N_24564);
and UO_2261 (O_2261,N_29885,N_25979);
nand UO_2262 (O_2262,N_24339,N_27143);
xor UO_2263 (O_2263,N_26051,N_28797);
nand UO_2264 (O_2264,N_24927,N_25571);
xnor UO_2265 (O_2265,N_29728,N_29455);
nand UO_2266 (O_2266,N_25640,N_26540);
xnor UO_2267 (O_2267,N_28534,N_29475);
nand UO_2268 (O_2268,N_24920,N_24568);
and UO_2269 (O_2269,N_26124,N_28862);
or UO_2270 (O_2270,N_26000,N_28948);
or UO_2271 (O_2271,N_25943,N_25130);
and UO_2272 (O_2272,N_26630,N_28695);
nor UO_2273 (O_2273,N_28178,N_28069);
nand UO_2274 (O_2274,N_27271,N_29174);
xnor UO_2275 (O_2275,N_24953,N_25307);
or UO_2276 (O_2276,N_25351,N_25420);
or UO_2277 (O_2277,N_24106,N_24603);
and UO_2278 (O_2278,N_25927,N_26428);
nor UO_2279 (O_2279,N_26638,N_24055);
xor UO_2280 (O_2280,N_27650,N_24067);
nand UO_2281 (O_2281,N_26451,N_28284);
nor UO_2282 (O_2282,N_26806,N_24690);
or UO_2283 (O_2283,N_27415,N_26244);
nor UO_2284 (O_2284,N_28372,N_24914);
and UO_2285 (O_2285,N_29398,N_24900);
nand UO_2286 (O_2286,N_28844,N_27302);
and UO_2287 (O_2287,N_25926,N_28089);
nor UO_2288 (O_2288,N_25281,N_25989);
nor UO_2289 (O_2289,N_24192,N_25701);
nor UO_2290 (O_2290,N_27931,N_28689);
and UO_2291 (O_2291,N_24620,N_27054);
nand UO_2292 (O_2292,N_27844,N_25833);
nand UO_2293 (O_2293,N_28320,N_24917);
or UO_2294 (O_2294,N_27387,N_24359);
xnor UO_2295 (O_2295,N_26083,N_29792);
or UO_2296 (O_2296,N_26548,N_25896);
or UO_2297 (O_2297,N_28959,N_28520);
xor UO_2298 (O_2298,N_24316,N_28808);
or UO_2299 (O_2299,N_29512,N_24983);
and UO_2300 (O_2300,N_28332,N_25029);
and UO_2301 (O_2301,N_26865,N_29686);
nor UO_2302 (O_2302,N_26326,N_24822);
or UO_2303 (O_2303,N_27322,N_26180);
nor UO_2304 (O_2304,N_25098,N_29521);
nand UO_2305 (O_2305,N_29406,N_26137);
nand UO_2306 (O_2306,N_25780,N_26993);
and UO_2307 (O_2307,N_29216,N_24459);
nand UO_2308 (O_2308,N_27035,N_26520);
or UO_2309 (O_2309,N_29143,N_25756);
nand UO_2310 (O_2310,N_29575,N_25705);
or UO_2311 (O_2311,N_28132,N_26889);
nand UO_2312 (O_2312,N_27858,N_26503);
nor UO_2313 (O_2313,N_28744,N_27666);
nand UO_2314 (O_2314,N_27424,N_26165);
xor UO_2315 (O_2315,N_27175,N_24355);
nor UO_2316 (O_2316,N_24781,N_27527);
xnor UO_2317 (O_2317,N_28275,N_27283);
nor UO_2318 (O_2318,N_24582,N_26283);
nand UO_2319 (O_2319,N_24615,N_29117);
nor UO_2320 (O_2320,N_25605,N_24197);
xnor UO_2321 (O_2321,N_27631,N_29192);
nand UO_2322 (O_2322,N_24651,N_25426);
xnor UO_2323 (O_2323,N_24541,N_24925);
nor UO_2324 (O_2324,N_25737,N_25583);
nor UO_2325 (O_2325,N_28816,N_28262);
nor UO_2326 (O_2326,N_27479,N_25581);
nand UO_2327 (O_2327,N_28251,N_25598);
xor UO_2328 (O_2328,N_24318,N_27397);
or UO_2329 (O_2329,N_27360,N_29764);
and UO_2330 (O_2330,N_29489,N_27939);
nand UO_2331 (O_2331,N_24700,N_25676);
xnor UO_2332 (O_2332,N_25903,N_29016);
or UO_2333 (O_2333,N_25052,N_27062);
or UO_2334 (O_2334,N_24233,N_27569);
nor UO_2335 (O_2335,N_26111,N_29718);
nand UO_2336 (O_2336,N_26069,N_25228);
nand UO_2337 (O_2337,N_25381,N_27390);
nor UO_2338 (O_2338,N_24841,N_25129);
nor UO_2339 (O_2339,N_27320,N_25824);
or UO_2340 (O_2340,N_28225,N_28512);
and UO_2341 (O_2341,N_28102,N_26043);
and UO_2342 (O_2342,N_24150,N_27981);
xor UO_2343 (O_2343,N_27076,N_26492);
nor UO_2344 (O_2344,N_27026,N_28100);
nand UO_2345 (O_2345,N_26298,N_26078);
nor UO_2346 (O_2346,N_24062,N_29965);
and UO_2347 (O_2347,N_28191,N_26249);
xor UO_2348 (O_2348,N_29456,N_25154);
and UO_2349 (O_2349,N_27958,N_29815);
nor UO_2350 (O_2350,N_29571,N_29518);
and UO_2351 (O_2351,N_29133,N_29214);
nor UO_2352 (O_2352,N_29713,N_24288);
nand UO_2353 (O_2353,N_29697,N_25767);
xnor UO_2354 (O_2354,N_28111,N_29609);
or UO_2355 (O_2355,N_24625,N_28947);
or UO_2356 (O_2356,N_26675,N_26521);
and UO_2357 (O_2357,N_26410,N_26898);
nand UO_2358 (O_2358,N_25053,N_29246);
and UO_2359 (O_2359,N_25178,N_26559);
nor UO_2360 (O_2360,N_27838,N_27371);
nor UO_2361 (O_2361,N_29660,N_26114);
and UO_2362 (O_2362,N_28328,N_27411);
or UO_2363 (O_2363,N_24637,N_24099);
or UO_2364 (O_2364,N_24225,N_25070);
nand UO_2365 (O_2365,N_26231,N_29636);
xor UO_2366 (O_2366,N_25219,N_24286);
or UO_2367 (O_2367,N_26390,N_29857);
and UO_2368 (O_2368,N_26024,N_27149);
nor UO_2369 (O_2369,N_28438,N_26944);
and UO_2370 (O_2370,N_28880,N_26125);
or UO_2371 (O_2371,N_27804,N_26179);
xor UO_2372 (O_2372,N_29556,N_24032);
nor UO_2373 (O_2373,N_26836,N_27771);
xnor UO_2374 (O_2374,N_28770,N_29492);
nor UO_2375 (O_2375,N_24772,N_24828);
xor UO_2376 (O_2376,N_24246,N_28317);
nand UO_2377 (O_2377,N_24063,N_26311);
nand UO_2378 (O_2378,N_29389,N_24510);
xnor UO_2379 (O_2379,N_27709,N_26444);
nand UO_2380 (O_2380,N_26979,N_29811);
nor UO_2381 (O_2381,N_27854,N_27400);
nand UO_2382 (O_2382,N_29099,N_28866);
xor UO_2383 (O_2383,N_28787,N_29069);
or UO_2384 (O_2384,N_29945,N_26383);
nor UO_2385 (O_2385,N_24120,N_29258);
nor UO_2386 (O_2386,N_28699,N_26047);
or UO_2387 (O_2387,N_25995,N_24100);
nor UO_2388 (O_2388,N_28318,N_24079);
and UO_2389 (O_2389,N_26486,N_28266);
nor UO_2390 (O_2390,N_28267,N_24989);
or UO_2391 (O_2391,N_27672,N_28602);
xor UO_2392 (O_2392,N_26134,N_29881);
xnor UO_2393 (O_2393,N_24926,N_27606);
nor UO_2394 (O_2394,N_26199,N_27557);
nand UO_2395 (O_2395,N_24486,N_26838);
nand UO_2396 (O_2396,N_24387,N_29603);
xnor UO_2397 (O_2397,N_24093,N_24183);
and UO_2398 (O_2398,N_28500,N_26743);
nor UO_2399 (O_2399,N_24719,N_29048);
and UO_2400 (O_2400,N_28037,N_24547);
and UO_2401 (O_2401,N_27319,N_27669);
nand UO_2402 (O_2402,N_24732,N_26251);
nand UO_2403 (O_2403,N_25340,N_29733);
nor UO_2404 (O_2404,N_29150,N_26273);
or UO_2405 (O_2405,N_27262,N_25764);
nor UO_2406 (O_2406,N_24962,N_29186);
nor UO_2407 (O_2407,N_27662,N_26037);
nand UO_2408 (O_2408,N_29705,N_26794);
xnor UO_2409 (O_2409,N_29770,N_25961);
nand UO_2410 (O_2410,N_25396,N_27878);
or UO_2411 (O_2411,N_24157,N_26214);
nand UO_2412 (O_2412,N_28883,N_29837);
xor UO_2413 (O_2413,N_25734,N_26054);
nand UO_2414 (O_2414,N_26699,N_27861);
nand UO_2415 (O_2415,N_25071,N_27731);
nor UO_2416 (O_2416,N_24315,N_28718);
nor UO_2417 (O_2417,N_24853,N_24710);
nand UO_2418 (O_2418,N_28697,N_24400);
xor UO_2419 (O_2419,N_27182,N_26146);
xnor UO_2420 (O_2420,N_28889,N_27135);
nand UO_2421 (O_2421,N_24389,N_28421);
nand UO_2422 (O_2422,N_29450,N_28645);
nand UO_2423 (O_2423,N_27956,N_28543);
xnor UO_2424 (O_2424,N_28871,N_26635);
and UO_2425 (O_2425,N_26150,N_28736);
and UO_2426 (O_2426,N_28958,N_26994);
and UO_2427 (O_2427,N_25109,N_28158);
xnor UO_2428 (O_2428,N_28798,N_29137);
or UO_2429 (O_2429,N_28058,N_28270);
and UO_2430 (O_2430,N_28600,N_25316);
and UO_2431 (O_2431,N_29653,N_24356);
nor UO_2432 (O_2432,N_25627,N_28327);
and UO_2433 (O_2433,N_25277,N_25227);
nand UO_2434 (O_2434,N_28325,N_25234);
xnor UO_2435 (O_2435,N_29779,N_28589);
and UO_2436 (O_2436,N_25552,N_25412);
nand UO_2437 (O_2437,N_25468,N_29464);
nor UO_2438 (O_2438,N_24074,N_25422);
and UO_2439 (O_2439,N_24673,N_28116);
nand UO_2440 (O_2440,N_28927,N_25717);
nand UO_2441 (O_2441,N_27616,N_26529);
and UO_2442 (O_2442,N_29875,N_27186);
nand UO_2443 (O_2443,N_29869,N_28652);
nor UO_2444 (O_2444,N_29002,N_29753);
nand UO_2445 (O_2445,N_29357,N_28503);
or UO_2446 (O_2446,N_28471,N_29957);
and UO_2447 (O_2447,N_28135,N_26934);
and UO_2448 (O_2448,N_29736,N_25333);
or UO_2449 (O_2449,N_29994,N_26333);
and UO_2450 (O_2450,N_24543,N_26573);
nor UO_2451 (O_2451,N_25621,N_27389);
and UO_2452 (O_2452,N_24949,N_29740);
nand UO_2453 (O_2453,N_29056,N_26415);
xnor UO_2454 (O_2454,N_25092,N_28910);
and UO_2455 (O_2455,N_25955,N_29129);
nor UO_2456 (O_2456,N_24061,N_28213);
nand UO_2457 (O_2457,N_29221,N_26186);
or UO_2458 (O_2458,N_27659,N_29457);
nor UO_2459 (O_2459,N_26178,N_27907);
nand UO_2460 (O_2460,N_25398,N_25620);
and UO_2461 (O_2461,N_25156,N_27082);
and UO_2462 (O_2462,N_29797,N_24638);
xor UO_2463 (O_2463,N_29639,N_25593);
nor UO_2464 (O_2464,N_24474,N_24614);
and UO_2465 (O_2465,N_27431,N_25242);
nor UO_2466 (O_2466,N_25645,N_24411);
xnor UO_2467 (O_2467,N_24583,N_26357);
and UO_2468 (O_2468,N_28997,N_28306);
or UO_2469 (O_2469,N_27152,N_29785);
xnor UO_2470 (O_2470,N_26201,N_24254);
nand UO_2471 (O_2471,N_27098,N_28249);
and UO_2472 (O_2472,N_29485,N_26060);
and UO_2473 (O_2473,N_24518,N_25255);
xor UO_2474 (O_2474,N_27950,N_29335);
nor UO_2475 (O_2475,N_27719,N_26962);
nor UO_2476 (O_2476,N_24802,N_26470);
nor UO_2477 (O_2477,N_29637,N_25027);
nand UO_2478 (O_2478,N_28140,N_24096);
or UO_2479 (O_2479,N_24190,N_25588);
nand UO_2480 (O_2480,N_26034,N_27050);
nand UO_2481 (O_2481,N_28141,N_28639);
xor UO_2482 (O_2482,N_26952,N_28420);
or UO_2483 (O_2483,N_27173,N_26330);
or UO_2484 (O_2484,N_28824,N_27055);
nor UO_2485 (O_2485,N_29987,N_28603);
and UO_2486 (O_2486,N_24025,N_25062);
nor UO_2487 (O_2487,N_27686,N_26601);
nor UO_2488 (O_2488,N_27994,N_28608);
nand UO_2489 (O_2489,N_29659,N_25807);
and UO_2490 (O_2490,N_27562,N_26287);
xnor UO_2491 (O_2491,N_27501,N_28488);
or UO_2492 (O_2492,N_27275,N_28004);
nor UO_2493 (O_2493,N_26604,N_26467);
xnor UO_2494 (O_2494,N_29301,N_24656);
nand UO_2495 (O_2495,N_26045,N_25271);
nand UO_2496 (O_2496,N_29700,N_29477);
xnor UO_2497 (O_2497,N_26452,N_24886);
and UO_2498 (O_2498,N_29795,N_27817);
or UO_2499 (O_2499,N_27814,N_28654);
xnor UO_2500 (O_2500,N_26713,N_28921);
nand UO_2501 (O_2501,N_29337,N_25658);
nand UO_2502 (O_2502,N_28290,N_26102);
xor UO_2503 (O_2503,N_26742,N_24391);
xor UO_2504 (O_2504,N_26437,N_25309);
or UO_2505 (O_2505,N_26629,N_29564);
nor UO_2506 (O_2506,N_27353,N_28127);
nor UO_2507 (O_2507,N_26837,N_28242);
nor UO_2508 (O_2508,N_26846,N_27019);
nand UO_2509 (O_2509,N_25114,N_28263);
and UO_2510 (O_2510,N_24794,N_24018);
xnor UO_2511 (O_2511,N_29649,N_27623);
nor UO_2512 (O_2512,N_29193,N_29351);
xnor UO_2513 (O_2513,N_27576,N_27190);
or UO_2514 (O_2514,N_27547,N_29678);
nor UO_2515 (O_2515,N_25619,N_28954);
nor UO_2516 (O_2516,N_24864,N_29248);
nand UO_2517 (O_2517,N_27800,N_25578);
xnor UO_2518 (O_2518,N_24860,N_27987);
nand UO_2519 (O_2519,N_27914,N_27721);
xnor UO_2520 (O_2520,N_25595,N_28846);
nor UO_2521 (O_2521,N_26226,N_25272);
nand UO_2522 (O_2522,N_27478,N_26033);
nor UO_2523 (O_2523,N_24576,N_27201);
nand UO_2524 (O_2524,N_27941,N_27695);
nand UO_2525 (O_2525,N_26093,N_29173);
or UO_2526 (O_2526,N_26584,N_29884);
and UO_2527 (O_2527,N_28174,N_27376);
or UO_2528 (O_2528,N_26703,N_27610);
or UO_2529 (O_2529,N_24565,N_27114);
and UO_2530 (O_2530,N_25652,N_28000);
xor UO_2531 (O_2531,N_26523,N_24911);
xnor UO_2532 (O_2532,N_26839,N_27420);
nor UO_2533 (O_2533,N_29865,N_25471);
and UO_2534 (O_2534,N_27205,N_29366);
nand UO_2535 (O_2535,N_29530,N_28101);
and UO_2536 (O_2536,N_29179,N_28725);
nor UO_2537 (O_2537,N_28288,N_25885);
xor UO_2538 (O_2538,N_29142,N_25781);
and UO_2539 (O_2539,N_25844,N_27486);
nand UO_2540 (O_2540,N_24088,N_29384);
nand UO_2541 (O_2541,N_24758,N_24965);
nor UO_2542 (O_2542,N_29243,N_25820);
nand UO_2543 (O_2543,N_25937,N_28869);
or UO_2544 (O_2544,N_25102,N_28335);
and UO_2545 (O_2545,N_26684,N_24784);
and UO_2546 (O_2546,N_26130,N_28696);
or UO_2547 (O_2547,N_27756,N_27534);
nand UO_2548 (O_2548,N_26887,N_25851);
nor UO_2549 (O_2549,N_28536,N_27150);
or UO_2550 (O_2550,N_24036,N_26118);
or UO_2551 (O_2551,N_29471,N_29579);
nor UO_2552 (O_2552,N_29280,N_26455);
or UO_2553 (O_2553,N_25067,N_27962);
and UO_2554 (O_2554,N_28163,N_28340);
nor UO_2555 (O_2555,N_28183,N_26923);
xnor UO_2556 (O_2556,N_25888,N_27248);
nor UO_2557 (O_2557,N_25805,N_29551);
or UO_2558 (O_2558,N_27312,N_29852);
xor UO_2559 (O_2559,N_24642,N_28646);
or UO_2560 (O_2560,N_25994,N_25743);
xnor UO_2561 (O_2561,N_24725,N_28764);
or UO_2562 (O_2562,N_28508,N_24243);
nand UO_2563 (O_2563,N_26248,N_29738);
nand UO_2564 (O_2564,N_29942,N_24530);
nor UO_2565 (O_2565,N_29289,N_25539);
and UO_2566 (O_2566,N_26627,N_24284);
nand UO_2567 (O_2567,N_25320,N_24017);
nand UO_2568 (O_2568,N_25853,N_26946);
nand UO_2569 (O_2569,N_26097,N_27930);
and UO_2570 (O_2570,N_24272,N_29370);
and UO_2571 (O_2571,N_28776,N_29023);
and UO_2572 (O_2572,N_26322,N_29346);
and UO_2573 (O_2573,N_25732,N_25039);
or UO_2574 (O_2574,N_29116,N_24581);
nor UO_2575 (O_2575,N_27030,N_28683);
nor UO_2576 (O_2576,N_28462,N_26970);
nand UO_2577 (O_2577,N_29008,N_28788);
nor UO_2578 (O_2578,N_24218,N_26429);
and UO_2579 (O_2579,N_25997,N_24460);
or UO_2580 (O_2580,N_26353,N_25104);
and UO_2581 (O_2581,N_24409,N_26029);
nand UO_2582 (O_2582,N_24887,N_27120);
nor UO_2583 (O_2583,N_25355,N_27427);
or UO_2584 (O_2584,N_29859,N_27193);
nand UO_2585 (O_2585,N_27581,N_29687);
nand UO_2586 (O_2586,N_25238,N_26654);
or UO_2587 (O_2587,N_26667,N_27810);
nand UO_2588 (O_2588,N_24624,N_24130);
or UO_2589 (O_2589,N_27942,N_27905);
xor UO_2590 (O_2590,N_25929,N_28490);
nor UO_2591 (O_2591,N_25061,N_24495);
nor UO_2592 (O_2592,N_25438,N_29064);
nor UO_2593 (O_2593,N_29147,N_25712);
nor UO_2594 (O_2594,N_26175,N_25860);
nand UO_2595 (O_2595,N_28034,N_29213);
nand UO_2596 (O_2596,N_26256,N_29816);
or UO_2597 (O_2597,N_26586,N_24184);
or UO_2598 (O_2598,N_25828,N_27197);
nor UO_2599 (O_2599,N_24112,N_28068);
nor UO_2600 (O_2600,N_27863,N_27601);
xor UO_2601 (O_2601,N_24211,N_25877);
or UO_2602 (O_2602,N_26340,N_28076);
and UO_2603 (O_2603,N_27280,N_25466);
or UO_2604 (O_2604,N_25133,N_26798);
nor UO_2605 (O_2605,N_29020,N_28804);
nand UO_2606 (O_2606,N_27900,N_29495);
and UO_2607 (O_2607,N_25305,N_24334);
xor UO_2608 (O_2608,N_25772,N_27577);
nand UO_2609 (O_2609,N_28562,N_28401);
and UO_2610 (O_2610,N_24010,N_28567);
or UO_2611 (O_2611,N_24049,N_29569);
or UO_2612 (O_2612,N_29760,N_29725);
or UO_2613 (O_2613,N_28015,N_29561);
xnor UO_2614 (O_2614,N_25951,N_28734);
xnor UO_2615 (O_2615,N_29592,N_28527);
or UO_2616 (O_2616,N_25917,N_29604);
or UO_2617 (O_2617,N_24277,N_26328);
nand UO_2618 (O_2618,N_25841,N_24159);
nand UO_2619 (O_2619,N_28617,N_24536);
nand UO_2620 (O_2620,N_27651,N_24161);
xor UO_2621 (O_2621,N_25292,N_28436);
nand UO_2622 (O_2622,N_28949,N_24923);
and UO_2623 (O_2623,N_27181,N_25218);
and UO_2624 (O_2624,N_26510,N_28229);
or UO_2625 (O_2625,N_28576,N_24761);
xor UO_2626 (O_2626,N_24868,N_27027);
and UO_2627 (O_2627,N_24399,N_28431);
xor UO_2628 (O_2628,N_27584,N_24469);
or UO_2629 (O_2629,N_28244,N_25299);
nand UO_2630 (O_2630,N_26775,N_26546);
nor UO_2631 (O_2631,N_29448,N_29403);
and UO_2632 (O_2632,N_27725,N_29294);
nor UO_2633 (O_2633,N_29386,N_27670);
or UO_2634 (O_2634,N_27889,N_29148);
nand UO_2635 (O_2635,N_26916,N_28607);
nor UO_2636 (O_2636,N_24986,N_27626);
nor UO_2637 (O_2637,N_24412,N_28821);
or UO_2638 (O_2638,N_24766,N_25032);
nand UO_2639 (O_2639,N_26771,N_28848);
or UO_2640 (O_2640,N_24504,N_24630);
nand UO_2641 (O_2641,N_28916,N_29443);
nor UO_2642 (O_2642,N_27187,N_25064);
and UO_2643 (O_2643,N_24121,N_24555);
nor UO_2644 (O_2644,N_24950,N_28605);
nor UO_2645 (O_2645,N_28721,N_29664);
and UO_2646 (O_2646,N_27298,N_25223);
nand UO_2647 (O_2647,N_29959,N_27913);
xnor UO_2648 (O_2648,N_27209,N_26040);
and UO_2649 (O_2649,N_28305,N_28219);
nor UO_2650 (O_2650,N_29958,N_27000);
nand UO_2651 (O_2651,N_29315,N_27247);
or UO_2652 (O_2652,N_28293,N_26655);
or UO_2653 (O_2653,N_28056,N_29264);
nor UO_2654 (O_2654,N_28917,N_25113);
nand UO_2655 (O_2655,N_27454,N_27909);
nor UO_2656 (O_2656,N_24398,N_28963);
nand UO_2657 (O_2657,N_28924,N_28329);
nor UO_2658 (O_2658,N_24528,N_28961);
nand UO_2659 (O_2659,N_29860,N_25131);
and UO_2660 (O_2660,N_25567,N_25586);
xor UO_2661 (O_2661,N_28739,N_28863);
nor UO_2662 (O_2662,N_24004,N_25719);
nand UO_2663 (O_2663,N_24940,N_27640);
nor UO_2664 (O_2664,N_27537,N_28212);
xnor UO_2665 (O_2665,N_27635,N_28413);
nor UO_2666 (O_2666,N_25263,N_29754);
xnor UO_2667 (O_2667,N_29360,N_27403);
nand UO_2668 (O_2668,N_27046,N_28098);
or UO_2669 (O_2669,N_27172,N_27433);
xnor UO_2670 (O_2670,N_26002,N_27674);
and UO_2671 (O_2671,N_26936,N_25690);
nand UO_2672 (O_2672,N_25144,N_26479);
nand UO_2673 (O_2673,N_26990,N_28655);
xnor UO_2674 (O_2674,N_29667,N_26733);
nor UO_2675 (O_2675,N_29092,N_29721);
nand UO_2676 (O_2676,N_24843,N_27888);
or UO_2677 (O_2677,N_27103,N_27943);
and UO_2678 (O_2678,N_27752,N_24856);
nor UO_2679 (O_2679,N_25939,N_24905);
nand UO_2680 (O_2680,N_24762,N_26528);
nand UO_2681 (O_2681,N_27957,N_25811);
xor UO_2682 (O_2682,N_29233,N_28182);
nand UO_2683 (O_2683,N_24768,N_24227);
nand UO_2684 (O_2684,N_26978,N_26823);
or UO_2685 (O_2685,N_29701,N_28546);
xor UO_2686 (O_2686,N_26862,N_25905);
or UO_2687 (O_2687,N_27028,N_25486);
nor UO_2688 (O_2688,N_29354,N_28377);
and UO_2689 (O_2689,N_27073,N_28882);
or UO_2690 (O_2690,N_29794,N_28071);
and UO_2691 (O_2691,N_25173,N_25759);
xor UO_2692 (O_2692,N_26115,N_24597);
nor UO_2693 (O_2693,N_27507,N_24776);
nor UO_2694 (O_2694,N_26341,N_27891);
nor UO_2695 (O_2695,N_29242,N_24874);
and UO_2696 (O_2696,N_24103,N_27001);
and UO_2697 (O_2697,N_29836,N_29749);
nand UO_2698 (O_2698,N_26293,N_24787);
nor UO_2699 (O_2699,N_24465,N_29310);
nor UO_2700 (O_2700,N_25049,N_28704);
nor UO_2701 (O_2701,N_27112,N_29196);
xnor UO_2702 (O_2702,N_26361,N_24427);
nand UO_2703 (O_2703,N_24627,N_29730);
or UO_2704 (O_2704,N_28036,N_27107);
or UO_2705 (O_2705,N_27514,N_26805);
nor UO_2706 (O_2706,N_25601,N_27333);
nand UO_2707 (O_2707,N_25192,N_27404);
xor UO_2708 (O_2708,N_24883,N_24921);
and UO_2709 (O_2709,N_28740,N_29827);
nor UO_2710 (O_2710,N_24475,N_27820);
and UO_2711 (O_2711,N_27751,N_26020);
nand UO_2712 (O_2712,N_29252,N_27528);
or UO_2713 (O_2713,N_27932,N_25207);
and UO_2714 (O_2714,N_25475,N_26009);
nand UO_2715 (O_2715,N_24978,N_24604);
or UO_2716 (O_2716,N_29358,N_29858);
or UO_2717 (O_2717,N_28123,N_24373);
and UO_2718 (O_2718,N_26066,N_27388);
or UO_2719 (O_2719,N_26128,N_26583);
and UO_2720 (O_2720,N_27505,N_25516);
and UO_2721 (O_2721,N_27852,N_26683);
and UO_2722 (O_2722,N_27438,N_24703);
nor UO_2723 (O_2723,N_24611,N_25337);
and UO_2724 (O_2724,N_24430,N_24199);
xor UO_2725 (O_2725,N_28084,N_24795);
xor UO_2726 (O_2726,N_25415,N_25254);
nand UO_2727 (O_2727,N_24842,N_27220);
and UO_2728 (O_2728,N_28322,N_24750);
nor UO_2729 (O_2729,N_27590,N_26913);
nand UO_2730 (O_2730,N_29916,N_29011);
and UO_2731 (O_2731,N_28453,N_28103);
and UO_2732 (O_2732,N_25222,N_27600);
nor UO_2733 (O_2733,N_29323,N_25387);
nor UO_2734 (O_2734,N_24372,N_27401);
nor UO_2735 (O_2735,N_24337,N_29407);
nand UO_2736 (O_2736,N_29694,N_28407);
or UO_2737 (O_2737,N_27691,N_28830);
nand UO_2738 (O_2738,N_25817,N_26618);
xor UO_2739 (O_2739,N_28473,N_25287);
nand UO_2740 (O_2740,N_27985,N_24767);
nor UO_2741 (O_2741,N_28509,N_24745);
nor UO_2742 (O_2742,N_25110,N_24361);
nor UO_2743 (O_2743,N_24397,N_24544);
nand UO_2744 (O_2744,N_27314,N_24618);
and UO_2745 (O_2745,N_27018,N_29305);
nor UO_2746 (O_2746,N_29200,N_24645);
and UO_2747 (O_2747,N_25667,N_25925);
or UO_2748 (O_2748,N_25030,N_25215);
and UO_2749 (O_2749,N_24366,N_25625);
or UO_2750 (O_2750,N_25327,N_26545);
nand UO_2751 (O_2751,N_29768,N_27366);
nor UO_2752 (O_2752,N_24467,N_26392);
and UO_2753 (O_2753,N_26317,N_28784);
xnor UO_2754 (O_2754,N_25093,N_24680);
or UO_2755 (O_2755,N_25890,N_27911);
nand UO_2756 (O_2756,N_29890,N_25868);
or UO_2757 (O_2757,N_25297,N_27880);
xor UO_2758 (O_2758,N_25020,N_27236);
nor UO_2759 (O_2759,N_26982,N_28763);
nand UO_2760 (O_2760,N_24426,N_28940);
and UO_2761 (O_2761,N_25490,N_26432);
and UO_2762 (O_2762,N_24283,N_25827);
xnor UO_2763 (O_2763,N_27164,N_26171);
and UO_2764 (O_2764,N_29580,N_28705);
and UO_2765 (O_2765,N_26818,N_29696);
nor UO_2766 (O_2766,N_29105,N_28342);
nand UO_2767 (O_2767,N_28389,N_25804);
nand UO_2768 (O_2768,N_27668,N_29136);
and UO_2769 (O_2769,N_29058,N_27224);
xnor UO_2770 (O_2770,N_26013,N_26501);
or UO_2771 (O_2771,N_24394,N_26342);
and UO_2772 (O_2772,N_26859,N_28759);
or UO_2773 (O_2773,N_27180,N_29203);
xor UO_2774 (O_2774,N_25199,N_29601);
nor UO_2775 (O_2775,N_29045,N_27776);
nor UO_2776 (O_2776,N_28134,N_28184);
xnor UO_2777 (O_2777,N_27365,N_26258);
or UO_2778 (O_2778,N_29739,N_27512);
or UO_2779 (O_2779,N_29010,N_25545);
xnor UO_2780 (O_2780,N_29932,N_24177);
or UO_2781 (O_2781,N_28789,N_26744);
and UO_2782 (O_2782,N_29862,N_25448);
or UO_2783 (O_2783,N_29037,N_26086);
and UO_2784 (O_2784,N_28521,N_25576);
or UO_2785 (O_2785,N_29887,N_29578);
and UO_2786 (O_2786,N_27959,N_28426);
nor UO_2787 (O_2787,N_25239,N_29820);
and UO_2788 (O_2788,N_28454,N_24311);
nor UO_2789 (O_2789,N_29187,N_24250);
or UO_2790 (O_2790,N_29879,N_27860);
nor UO_2791 (O_2791,N_28581,N_27699);
or UO_2792 (O_2792,N_28052,N_26596);
xor UO_2793 (O_2793,N_26378,N_27990);
or UO_2794 (O_2794,N_28964,N_29081);
nor UO_2795 (O_2795,N_26126,N_25196);
xor UO_2796 (O_2796,N_28988,N_26825);
nor UO_2797 (O_2797,N_28858,N_24252);
and UO_2798 (O_2798,N_26210,N_26748);
nand UO_2799 (O_2799,N_28992,N_26885);
nand UO_2800 (O_2800,N_28485,N_25010);
xor UO_2801 (O_2801,N_25533,N_29347);
and UO_2802 (O_2802,N_24363,N_26662);
xnor UO_2803 (O_2803,N_29789,N_24897);
nor UO_2804 (O_2804,N_28919,N_29538);
nand UO_2805 (O_2805,N_27113,N_26656);
or UO_2806 (O_2806,N_28803,N_28781);
xor UO_2807 (O_2807,N_29043,N_25789);
nand UO_2808 (O_2808,N_28156,N_27791);
xnor UO_2809 (O_2809,N_26087,N_29427);
or UO_2810 (O_2810,N_29602,N_28643);
or UO_2811 (O_2811,N_29286,N_25655);
nand UO_2812 (O_2812,N_28786,N_24261);
nand UO_2813 (O_2813,N_26220,N_25160);
xor UO_2814 (O_2814,N_27803,N_26502);
xnor UO_2815 (O_2815,N_29633,N_26144);
nor UO_2816 (O_2816,N_29813,N_26089);
and UO_2817 (O_2817,N_26826,N_25087);
xnor UO_2818 (O_2818,N_27355,N_29918);
or UO_2819 (O_2819,N_29548,N_25361);
or UO_2820 (O_2820,N_28555,N_29634);
nor UO_2821 (O_2821,N_28171,N_26259);
nand UO_2822 (O_2822,N_24720,N_27786);
nor UO_2823 (O_2823,N_24880,N_27954);
and UO_2824 (O_2824,N_29929,N_25935);
xor UO_2825 (O_2825,N_26200,N_29576);
and UO_2826 (O_2826,N_25707,N_26620);
nand UO_2827 (O_2827,N_26623,N_27824);
xor UO_2828 (O_2828,N_25990,N_26735);
and UO_2829 (O_2829,N_27882,N_29973);
xnor UO_2830 (O_2830,N_27848,N_26506);
nand UO_2831 (O_2831,N_29666,N_25548);
or UO_2832 (O_2832,N_24545,N_29774);
and UO_2833 (O_2833,N_27872,N_25693);
nand UO_2834 (O_2834,N_24713,N_29052);
nor UO_2835 (O_2835,N_24384,N_28209);
nor UO_2836 (O_2836,N_27846,N_29804);
xor UO_2837 (O_2837,N_26286,N_24687);
nor UO_2838 (O_2838,N_25143,N_24804);
nor UO_2839 (O_2839,N_28253,N_27571);
nand UO_2840 (O_2840,N_25542,N_28499);
xnor UO_2841 (O_2841,N_27437,N_25084);
or UO_2842 (O_2842,N_25969,N_25985);
nand UO_2843 (O_2843,N_26572,N_26857);
nand UO_2844 (O_2844,N_28430,N_24141);
or UO_2845 (O_2845,N_27629,N_25769);
nand UO_2846 (O_2846,N_26753,N_27762);
nand UO_2847 (O_2847,N_29972,N_27155);
or UO_2848 (O_2848,N_28367,N_25457);
or UO_2849 (O_2849,N_25182,N_25174);
nand UO_2850 (O_2850,N_25407,N_24365);
xor UO_2851 (O_2851,N_27290,N_28668);
xor UO_2852 (O_2852,N_29988,N_26075);
and UO_2853 (O_2853,N_25527,N_24220);
and UO_2854 (O_2854,N_28308,N_28677);
nand UO_2855 (O_2855,N_27545,N_26588);
and UO_2856 (O_2856,N_24118,N_24237);
nand UO_2857 (O_2857,N_27254,N_24503);
nor UO_2858 (O_2858,N_27381,N_25502);
nor UO_2859 (O_2859,N_26981,N_27004);
xnor UO_2860 (O_2860,N_29931,N_26614);
and UO_2861 (O_2861,N_29114,N_29134);
or UO_2862 (O_2862,N_27802,N_29831);
xor UO_2863 (O_2863,N_27476,N_27952);
and UO_2864 (O_2864,N_26414,N_26508);
xnor UO_2865 (O_2865,N_29365,N_24896);
xnor UO_2866 (O_2866,N_27072,N_28506);
or UO_2867 (O_2867,N_24166,N_27003);
xor UO_2868 (O_2868,N_26670,N_26537);
and UO_2869 (O_2869,N_29141,N_25859);
and UO_2870 (O_2870,N_26252,N_28307);
or UO_2871 (O_2871,N_24354,N_28946);
and UO_2872 (O_2872,N_25151,N_29050);
nand UO_2873 (O_2873,N_28651,N_26346);
or UO_2874 (O_2874,N_27081,N_26612);
nor UO_2875 (O_2875,N_27602,N_25293);
xnor UO_2876 (O_2876,N_29632,N_26016);
nor UO_2877 (O_2877,N_24996,N_25479);
xnor UO_2878 (O_2878,N_29939,N_25476);
and UO_2879 (O_2879,N_28692,N_25018);
nor UO_2880 (O_2880,N_25513,N_24674);
nor UO_2881 (O_2881,N_26424,N_29205);
nor UO_2882 (O_2882,N_27202,N_24979);
nor UO_2883 (O_2883,N_24601,N_29851);
and UO_2884 (O_2884,N_28093,N_28211);
or UO_2885 (O_2885,N_25267,N_26385);
or UO_2886 (O_2886,N_25443,N_26309);
and UO_2887 (O_2887,N_26417,N_29788);
and UO_2888 (O_2888,N_29599,N_25568);
nand UO_2889 (O_2889,N_25091,N_25076);
and UO_2890 (O_2890,N_24174,N_25510);
xnor UO_2891 (O_2891,N_27260,N_29786);
nor UO_2892 (O_2892,N_25826,N_29984);
xnor UO_2893 (O_2893,N_26403,N_26242);
and UO_2894 (O_2894,N_27471,N_25556);
nand UO_2895 (O_2895,N_26720,N_26339);
nor UO_2896 (O_2896,N_24145,N_27069);
xor UO_2897 (O_2897,N_28745,N_25217);
xor UO_2898 (O_2898,N_26569,N_24800);
xor UO_2899 (O_2899,N_26512,N_27720);
nand UO_2900 (O_2900,N_26364,N_29524);
or UO_2901 (O_2901,N_28684,N_25558);
and UO_2902 (O_2902,N_28714,N_28402);
nor UO_2903 (O_2903,N_25419,N_26041);
or UO_2904 (O_2904,N_24241,N_25467);
nor UO_2905 (O_2905,N_29473,N_24488);
nand UO_2906 (O_2906,N_24712,N_27023);
or UO_2907 (O_2907,N_27536,N_24931);
xnor UO_2908 (O_2908,N_24600,N_29829);
and UO_2909 (O_2909,N_27976,N_29009);
or UO_2910 (O_2910,N_28703,N_29372);
xnor UO_2911 (O_2911,N_29924,N_29861);
or UO_2912 (O_2912,N_25229,N_28756);
and UO_2913 (O_2913,N_26345,N_28224);
xnor UO_2914 (O_2914,N_24020,N_29281);
or UO_2915 (O_2915,N_27367,N_29097);
nor UO_2916 (O_2916,N_28016,N_27587);
nand UO_2917 (O_2917,N_26464,N_29743);
or UO_2918 (O_2918,N_27165,N_25646);
nor UO_2919 (O_2919,N_25522,N_24514);
nor UO_2920 (O_2920,N_24152,N_28806);
nor UO_2921 (O_2921,N_24202,N_25177);
nand UO_2922 (O_2922,N_26227,N_24439);
and UO_2923 (O_2923,N_25816,N_25159);
or UO_2924 (O_2924,N_25547,N_29706);
and UO_2925 (O_2925,N_29882,N_28836);
xor UO_2926 (O_2926,N_25863,N_24273);
or UO_2927 (O_2927,N_25944,N_25848);
or UO_2928 (O_2928,N_29329,N_24452);
or UO_2929 (O_2929,N_25425,N_29808);
or UO_2930 (O_2930,N_29625,N_29872);
xor UO_2931 (O_2931,N_24451,N_25521);
nand UO_2932 (O_2932,N_28154,N_25385);
nor UO_2933 (O_2933,N_24312,N_24817);
nand UO_2934 (O_2934,N_26711,N_25602);
nand UO_2935 (O_2935,N_27096,N_24215);
xor UO_2936 (O_2936,N_29466,N_27523);
and UO_2937 (O_2937,N_29245,N_25274);
nor UO_2938 (O_2938,N_29237,N_29047);
and UO_2939 (O_2939,N_27612,N_28870);
or UO_2940 (O_2940,N_27048,N_29679);
and UO_2941 (O_2941,N_29426,N_27774);
xor UO_2942 (O_2942,N_29103,N_28460);
xor UO_2943 (O_2943,N_27045,N_25416);
and UO_2944 (O_2944,N_25043,N_28523);
xnor UO_2945 (O_2945,N_27270,N_29012);
or UO_2946 (O_2946,N_28841,N_29717);
and UO_2947 (O_2947,N_25201,N_25782);
nor UO_2948 (O_2948,N_28254,N_24952);
and UO_2949 (O_2949,N_29642,N_26427);
xor UO_2950 (O_2950,N_28176,N_25474);
and UO_2951 (O_2951,N_28999,N_27279);
xor UO_2952 (O_2952,N_27347,N_29342);
nor UO_2953 (O_2953,N_29977,N_27509);
nor UO_2954 (O_2954,N_27176,N_29490);
xor UO_2955 (O_2955,N_29015,N_24859);
nand UO_2956 (O_2956,N_27738,N_27573);
xnor UO_2957 (O_2957,N_29657,N_26133);
xnor UO_2958 (O_2958,N_24839,N_25685);
and UO_2959 (O_2959,N_27556,N_26553);
or UO_2960 (O_2960,N_26648,N_29909);
xor UO_2961 (O_2961,N_27847,N_25075);
xnor UO_2962 (O_2962,N_26940,N_25458);
xor UO_2963 (O_2963,N_25722,N_29558);
and UO_2964 (O_2964,N_27087,N_24783);
and UO_2965 (O_2965,N_28990,N_26541);
xnor UO_2966 (O_2966,N_25893,N_25596);
nor UO_2967 (O_2967,N_28748,N_25590);
xnor UO_2968 (O_2968,N_28269,N_24437);
nand UO_2969 (O_2969,N_29981,N_29144);
and UO_2970 (O_2970,N_27506,N_28554);
nor UO_2971 (O_2971,N_24913,N_25382);
or UO_2972 (O_2972,N_27232,N_25799);
xnor UO_2973 (O_2973,N_28979,N_27038);
nand UO_2974 (O_2974,N_25006,N_27935);
and UO_2975 (O_2975,N_25134,N_27697);
xnor UO_2976 (O_2976,N_26232,N_27805);
and UO_2977 (O_2977,N_24752,N_28511);
nand UO_2978 (O_2978,N_25538,N_24538);
xor UO_2979 (O_2979,N_28583,N_28094);
or UO_2980 (O_2980,N_28486,N_29620);
or UO_2981 (O_2981,N_27915,N_25366);
nand UO_2982 (O_2982,N_24269,N_27088);
or UO_2983 (O_2983,N_25106,N_24948);
and UO_2984 (O_2984,N_29106,N_26228);
xnor UO_2985 (O_2985,N_27970,N_24744);
nand UO_2986 (O_2986,N_28280,N_26789);
and UO_2987 (O_2987,N_29288,N_25112);
xnor UO_2988 (O_2988,N_25298,N_24232);
and UO_2989 (O_2989,N_29375,N_24012);
xnor UO_2990 (O_2990,N_29928,N_26406);
or UO_2991 (O_2991,N_27639,N_29465);
nor UO_2992 (O_2992,N_25250,N_24867);
xnor UO_2993 (O_2993,N_24468,N_29316);
or UO_2994 (O_2994,N_27758,N_25639);
or UO_2995 (O_2995,N_26650,N_24907);
xnor UO_2996 (O_2996,N_27136,N_24051);
nand UO_2997 (O_2997,N_24410,N_27261);
and UO_2998 (O_2998,N_27574,N_27608);
xor UO_2999 (O_2999,N_24123,N_27313);
and UO_3000 (O_3000,N_24193,N_25862);
nand UO_3001 (O_3001,N_27757,N_27394);
and UO_3002 (O_3002,N_29793,N_27990);
and UO_3003 (O_3003,N_25433,N_27238);
or UO_3004 (O_3004,N_26991,N_25085);
xor UO_3005 (O_3005,N_26913,N_24857);
nor UO_3006 (O_3006,N_25450,N_27219);
nor UO_3007 (O_3007,N_29371,N_28484);
and UO_3008 (O_3008,N_29728,N_25382);
nor UO_3009 (O_3009,N_27435,N_28198);
or UO_3010 (O_3010,N_28684,N_28009);
or UO_3011 (O_3011,N_27391,N_27610);
nor UO_3012 (O_3012,N_26933,N_29235);
nand UO_3013 (O_3013,N_26527,N_24579);
nor UO_3014 (O_3014,N_28359,N_26562);
xor UO_3015 (O_3015,N_25580,N_24899);
and UO_3016 (O_3016,N_25846,N_27085);
nor UO_3017 (O_3017,N_24303,N_24818);
nand UO_3018 (O_3018,N_29593,N_28018);
nor UO_3019 (O_3019,N_27949,N_25414);
nand UO_3020 (O_3020,N_26356,N_28783);
xor UO_3021 (O_3021,N_24521,N_28253);
and UO_3022 (O_3022,N_26666,N_27422);
xnor UO_3023 (O_3023,N_24212,N_24745);
and UO_3024 (O_3024,N_28546,N_27974);
nor UO_3025 (O_3025,N_26537,N_27869);
and UO_3026 (O_3026,N_28899,N_24447);
and UO_3027 (O_3027,N_26154,N_29156);
or UO_3028 (O_3028,N_29127,N_29212);
or UO_3029 (O_3029,N_26524,N_26309);
nor UO_3030 (O_3030,N_26816,N_25259);
and UO_3031 (O_3031,N_27942,N_29267);
xnor UO_3032 (O_3032,N_27778,N_28374);
xnor UO_3033 (O_3033,N_25655,N_28824);
xnor UO_3034 (O_3034,N_29652,N_29920);
nor UO_3035 (O_3035,N_24822,N_29539);
and UO_3036 (O_3036,N_24816,N_28328);
nor UO_3037 (O_3037,N_26995,N_27595);
and UO_3038 (O_3038,N_28047,N_29622);
xor UO_3039 (O_3039,N_25935,N_29844);
nor UO_3040 (O_3040,N_25372,N_29244);
xor UO_3041 (O_3041,N_24660,N_27307);
or UO_3042 (O_3042,N_25592,N_29787);
nand UO_3043 (O_3043,N_28597,N_26668);
nor UO_3044 (O_3044,N_24394,N_26952);
xnor UO_3045 (O_3045,N_28966,N_28502);
nor UO_3046 (O_3046,N_29121,N_24074);
nand UO_3047 (O_3047,N_29583,N_29332);
xnor UO_3048 (O_3048,N_24068,N_28874);
xnor UO_3049 (O_3049,N_28536,N_25232);
nor UO_3050 (O_3050,N_29507,N_24407);
or UO_3051 (O_3051,N_25283,N_24222);
and UO_3052 (O_3052,N_28941,N_24310);
nor UO_3053 (O_3053,N_26864,N_29959);
nand UO_3054 (O_3054,N_26015,N_28467);
or UO_3055 (O_3055,N_25278,N_25956);
or UO_3056 (O_3056,N_27888,N_29790);
nor UO_3057 (O_3057,N_29924,N_24070);
or UO_3058 (O_3058,N_27823,N_24811);
and UO_3059 (O_3059,N_27669,N_28128);
xnor UO_3060 (O_3060,N_29210,N_28889);
nor UO_3061 (O_3061,N_29264,N_25037);
xor UO_3062 (O_3062,N_24490,N_27010);
nor UO_3063 (O_3063,N_28639,N_29483);
or UO_3064 (O_3064,N_27513,N_27734);
or UO_3065 (O_3065,N_28370,N_25534);
and UO_3066 (O_3066,N_27824,N_24489);
and UO_3067 (O_3067,N_26371,N_27724);
xnor UO_3068 (O_3068,N_25959,N_29846);
nor UO_3069 (O_3069,N_29163,N_29104);
xor UO_3070 (O_3070,N_26356,N_28373);
xnor UO_3071 (O_3071,N_29213,N_26790);
xor UO_3072 (O_3072,N_26384,N_25591);
xor UO_3073 (O_3073,N_26986,N_29224);
xnor UO_3074 (O_3074,N_25464,N_25371);
xnor UO_3075 (O_3075,N_28673,N_25915);
and UO_3076 (O_3076,N_25944,N_26078);
or UO_3077 (O_3077,N_25933,N_27873);
and UO_3078 (O_3078,N_26875,N_27847);
xor UO_3079 (O_3079,N_28312,N_24149);
and UO_3080 (O_3080,N_24881,N_29078);
xnor UO_3081 (O_3081,N_26351,N_29924);
and UO_3082 (O_3082,N_24626,N_26228);
xnor UO_3083 (O_3083,N_25972,N_25452);
nand UO_3084 (O_3084,N_26950,N_28814);
xnor UO_3085 (O_3085,N_27690,N_27707);
and UO_3086 (O_3086,N_28706,N_26483);
xor UO_3087 (O_3087,N_26891,N_26326);
or UO_3088 (O_3088,N_29814,N_29315);
or UO_3089 (O_3089,N_26706,N_25935);
or UO_3090 (O_3090,N_27343,N_26559);
xor UO_3091 (O_3091,N_27854,N_25977);
nand UO_3092 (O_3092,N_26304,N_28876);
nand UO_3093 (O_3093,N_26746,N_25185);
nor UO_3094 (O_3094,N_29995,N_26182);
nor UO_3095 (O_3095,N_28251,N_27498);
nand UO_3096 (O_3096,N_29280,N_28288);
nor UO_3097 (O_3097,N_29095,N_26577);
nand UO_3098 (O_3098,N_27276,N_25486);
nand UO_3099 (O_3099,N_26730,N_29940);
nor UO_3100 (O_3100,N_28010,N_24171);
or UO_3101 (O_3101,N_26812,N_28916);
nor UO_3102 (O_3102,N_25247,N_26821);
and UO_3103 (O_3103,N_27044,N_28986);
xor UO_3104 (O_3104,N_29261,N_27039);
nand UO_3105 (O_3105,N_27291,N_28397);
and UO_3106 (O_3106,N_29587,N_26501);
xor UO_3107 (O_3107,N_25129,N_24091);
nor UO_3108 (O_3108,N_24134,N_25680);
or UO_3109 (O_3109,N_24307,N_28480);
nand UO_3110 (O_3110,N_26190,N_29000);
and UO_3111 (O_3111,N_29607,N_25283);
or UO_3112 (O_3112,N_24835,N_26693);
or UO_3113 (O_3113,N_24145,N_28397);
nor UO_3114 (O_3114,N_26466,N_28892);
or UO_3115 (O_3115,N_25725,N_24447);
and UO_3116 (O_3116,N_25443,N_29776);
and UO_3117 (O_3117,N_24802,N_24269);
nand UO_3118 (O_3118,N_26095,N_25961);
and UO_3119 (O_3119,N_26652,N_29708);
or UO_3120 (O_3120,N_25206,N_27837);
and UO_3121 (O_3121,N_28582,N_27045);
or UO_3122 (O_3122,N_27415,N_29034);
nor UO_3123 (O_3123,N_28415,N_28381);
or UO_3124 (O_3124,N_28537,N_25369);
nor UO_3125 (O_3125,N_27782,N_28683);
nor UO_3126 (O_3126,N_29263,N_25637);
or UO_3127 (O_3127,N_29287,N_24401);
and UO_3128 (O_3128,N_26658,N_28205);
xor UO_3129 (O_3129,N_26700,N_27083);
xnor UO_3130 (O_3130,N_28738,N_26866);
xnor UO_3131 (O_3131,N_24926,N_28331);
and UO_3132 (O_3132,N_28091,N_28582);
nor UO_3133 (O_3133,N_27481,N_24928);
nand UO_3134 (O_3134,N_29104,N_28725);
or UO_3135 (O_3135,N_24030,N_25295);
nand UO_3136 (O_3136,N_28764,N_24836);
or UO_3137 (O_3137,N_27809,N_29851);
nor UO_3138 (O_3138,N_29807,N_24923);
and UO_3139 (O_3139,N_24733,N_28869);
nor UO_3140 (O_3140,N_27522,N_25780);
and UO_3141 (O_3141,N_29080,N_27446);
and UO_3142 (O_3142,N_29579,N_29000);
and UO_3143 (O_3143,N_28139,N_28929);
and UO_3144 (O_3144,N_29370,N_25230);
and UO_3145 (O_3145,N_28225,N_29337);
nand UO_3146 (O_3146,N_26976,N_27117);
nor UO_3147 (O_3147,N_28038,N_29276);
and UO_3148 (O_3148,N_25973,N_25758);
or UO_3149 (O_3149,N_25106,N_26306);
nor UO_3150 (O_3150,N_26063,N_29025);
nand UO_3151 (O_3151,N_28930,N_25578);
or UO_3152 (O_3152,N_24902,N_29375);
or UO_3153 (O_3153,N_24836,N_25904);
xnor UO_3154 (O_3154,N_26929,N_27243);
and UO_3155 (O_3155,N_25151,N_24201);
or UO_3156 (O_3156,N_26778,N_25775);
or UO_3157 (O_3157,N_29249,N_29627);
nand UO_3158 (O_3158,N_28382,N_27841);
nor UO_3159 (O_3159,N_26194,N_26190);
or UO_3160 (O_3160,N_28236,N_24243);
nand UO_3161 (O_3161,N_27119,N_29168);
and UO_3162 (O_3162,N_29821,N_29038);
and UO_3163 (O_3163,N_27828,N_24885);
xnor UO_3164 (O_3164,N_24320,N_24568);
or UO_3165 (O_3165,N_25173,N_25426);
xor UO_3166 (O_3166,N_29455,N_28641);
xnor UO_3167 (O_3167,N_29263,N_28168);
xnor UO_3168 (O_3168,N_28016,N_27413);
nor UO_3169 (O_3169,N_29752,N_26290);
nand UO_3170 (O_3170,N_24243,N_29929);
or UO_3171 (O_3171,N_29014,N_24925);
nand UO_3172 (O_3172,N_27216,N_25654);
nand UO_3173 (O_3173,N_29552,N_25617);
xnor UO_3174 (O_3174,N_29306,N_26487);
or UO_3175 (O_3175,N_25699,N_27240);
and UO_3176 (O_3176,N_25542,N_24153);
and UO_3177 (O_3177,N_29781,N_26448);
nor UO_3178 (O_3178,N_27998,N_27240);
xnor UO_3179 (O_3179,N_27230,N_29954);
or UO_3180 (O_3180,N_27562,N_26477);
or UO_3181 (O_3181,N_28624,N_27701);
nand UO_3182 (O_3182,N_26842,N_29763);
and UO_3183 (O_3183,N_27829,N_24574);
and UO_3184 (O_3184,N_28141,N_27339);
nor UO_3185 (O_3185,N_26254,N_29158);
xor UO_3186 (O_3186,N_26926,N_24925);
xor UO_3187 (O_3187,N_26494,N_29588);
xnor UO_3188 (O_3188,N_28118,N_28598);
and UO_3189 (O_3189,N_28981,N_28466);
or UO_3190 (O_3190,N_27017,N_27755);
or UO_3191 (O_3191,N_26938,N_25767);
or UO_3192 (O_3192,N_27631,N_28883);
or UO_3193 (O_3193,N_25659,N_24130);
xnor UO_3194 (O_3194,N_27925,N_25185);
and UO_3195 (O_3195,N_27268,N_24669);
or UO_3196 (O_3196,N_27459,N_25989);
nor UO_3197 (O_3197,N_28184,N_27782);
nand UO_3198 (O_3198,N_29984,N_29809);
xnor UO_3199 (O_3199,N_25918,N_29590);
nor UO_3200 (O_3200,N_28510,N_24186);
or UO_3201 (O_3201,N_24557,N_27806);
or UO_3202 (O_3202,N_26226,N_28073);
xnor UO_3203 (O_3203,N_25491,N_29018);
or UO_3204 (O_3204,N_26154,N_26193);
nor UO_3205 (O_3205,N_25761,N_26804);
nand UO_3206 (O_3206,N_25867,N_29751);
or UO_3207 (O_3207,N_29474,N_26898);
and UO_3208 (O_3208,N_26302,N_24060);
nor UO_3209 (O_3209,N_25861,N_24564);
and UO_3210 (O_3210,N_24819,N_29257);
or UO_3211 (O_3211,N_24820,N_25380);
nor UO_3212 (O_3212,N_25369,N_26429);
nor UO_3213 (O_3213,N_29545,N_29218);
xor UO_3214 (O_3214,N_27386,N_25096);
nor UO_3215 (O_3215,N_25468,N_28677);
nand UO_3216 (O_3216,N_27530,N_27756);
or UO_3217 (O_3217,N_26940,N_27813);
and UO_3218 (O_3218,N_29899,N_24663);
nor UO_3219 (O_3219,N_26555,N_29892);
and UO_3220 (O_3220,N_26968,N_29181);
or UO_3221 (O_3221,N_27462,N_26659);
xor UO_3222 (O_3222,N_25695,N_29885);
or UO_3223 (O_3223,N_24427,N_28369);
nand UO_3224 (O_3224,N_29577,N_26019);
or UO_3225 (O_3225,N_27849,N_28626);
nand UO_3226 (O_3226,N_29921,N_26504);
nor UO_3227 (O_3227,N_28681,N_24003);
and UO_3228 (O_3228,N_27953,N_26059);
or UO_3229 (O_3229,N_27423,N_28825);
nand UO_3230 (O_3230,N_26924,N_24662);
nor UO_3231 (O_3231,N_29015,N_28339);
or UO_3232 (O_3232,N_28461,N_29262);
or UO_3233 (O_3233,N_24963,N_27504);
xor UO_3234 (O_3234,N_28079,N_24014);
or UO_3235 (O_3235,N_24753,N_28621);
or UO_3236 (O_3236,N_28279,N_29856);
nor UO_3237 (O_3237,N_24377,N_27587);
or UO_3238 (O_3238,N_24399,N_27997);
or UO_3239 (O_3239,N_27247,N_29424);
nor UO_3240 (O_3240,N_26851,N_28885);
nand UO_3241 (O_3241,N_27470,N_24414);
and UO_3242 (O_3242,N_29876,N_28567);
nor UO_3243 (O_3243,N_26082,N_25233);
nor UO_3244 (O_3244,N_26393,N_28841);
xnor UO_3245 (O_3245,N_27044,N_29827);
xor UO_3246 (O_3246,N_29316,N_27254);
or UO_3247 (O_3247,N_28524,N_29257);
nand UO_3248 (O_3248,N_26498,N_28029);
nand UO_3249 (O_3249,N_29086,N_25100);
and UO_3250 (O_3250,N_25554,N_28465);
and UO_3251 (O_3251,N_27096,N_24204);
nand UO_3252 (O_3252,N_29846,N_28788);
nand UO_3253 (O_3253,N_25727,N_27213);
and UO_3254 (O_3254,N_28235,N_28568);
nand UO_3255 (O_3255,N_28964,N_29586);
xor UO_3256 (O_3256,N_24910,N_29355);
nor UO_3257 (O_3257,N_26871,N_29614);
and UO_3258 (O_3258,N_28073,N_25118);
nor UO_3259 (O_3259,N_28819,N_25462);
nand UO_3260 (O_3260,N_28291,N_29380);
xor UO_3261 (O_3261,N_25388,N_24149);
or UO_3262 (O_3262,N_26171,N_28324);
and UO_3263 (O_3263,N_25349,N_25924);
and UO_3264 (O_3264,N_24167,N_25719);
and UO_3265 (O_3265,N_29753,N_24482);
and UO_3266 (O_3266,N_29103,N_28203);
nor UO_3267 (O_3267,N_24279,N_27600);
nor UO_3268 (O_3268,N_25714,N_25311);
and UO_3269 (O_3269,N_28983,N_26975);
nand UO_3270 (O_3270,N_28916,N_27095);
or UO_3271 (O_3271,N_27656,N_29514);
or UO_3272 (O_3272,N_28864,N_28013);
nand UO_3273 (O_3273,N_27937,N_25987);
and UO_3274 (O_3274,N_25135,N_25127);
nor UO_3275 (O_3275,N_29053,N_27495);
or UO_3276 (O_3276,N_24873,N_26568);
xor UO_3277 (O_3277,N_26069,N_24288);
xor UO_3278 (O_3278,N_29244,N_29104);
nor UO_3279 (O_3279,N_28193,N_26442);
nand UO_3280 (O_3280,N_28713,N_27937);
nor UO_3281 (O_3281,N_26703,N_27409);
nand UO_3282 (O_3282,N_26974,N_28433);
or UO_3283 (O_3283,N_24757,N_27269);
or UO_3284 (O_3284,N_25764,N_27289);
nor UO_3285 (O_3285,N_29672,N_28519);
and UO_3286 (O_3286,N_29686,N_24646);
and UO_3287 (O_3287,N_29509,N_25017);
or UO_3288 (O_3288,N_26069,N_28942);
xnor UO_3289 (O_3289,N_28891,N_29553);
xor UO_3290 (O_3290,N_26775,N_29421);
nand UO_3291 (O_3291,N_25132,N_24513);
nand UO_3292 (O_3292,N_27000,N_26803);
and UO_3293 (O_3293,N_26477,N_26985);
and UO_3294 (O_3294,N_24622,N_27582);
or UO_3295 (O_3295,N_28968,N_29280);
or UO_3296 (O_3296,N_28909,N_25931);
nand UO_3297 (O_3297,N_29692,N_25528);
and UO_3298 (O_3298,N_27431,N_24100);
and UO_3299 (O_3299,N_27040,N_25900);
xor UO_3300 (O_3300,N_28573,N_29043);
nor UO_3301 (O_3301,N_26727,N_26885);
nand UO_3302 (O_3302,N_24235,N_24379);
and UO_3303 (O_3303,N_27645,N_26437);
and UO_3304 (O_3304,N_25352,N_27205);
nor UO_3305 (O_3305,N_29217,N_25077);
or UO_3306 (O_3306,N_29761,N_25335);
nor UO_3307 (O_3307,N_26057,N_29674);
or UO_3308 (O_3308,N_28898,N_29205);
nor UO_3309 (O_3309,N_24125,N_28904);
xor UO_3310 (O_3310,N_28983,N_25735);
or UO_3311 (O_3311,N_26482,N_27923);
xor UO_3312 (O_3312,N_26349,N_29714);
or UO_3313 (O_3313,N_27349,N_25097);
nand UO_3314 (O_3314,N_27362,N_25666);
or UO_3315 (O_3315,N_28739,N_27404);
and UO_3316 (O_3316,N_29600,N_25204);
nand UO_3317 (O_3317,N_28163,N_27054);
nor UO_3318 (O_3318,N_27242,N_29421);
nand UO_3319 (O_3319,N_26490,N_26542);
nor UO_3320 (O_3320,N_29898,N_26748);
nor UO_3321 (O_3321,N_28146,N_24494);
nor UO_3322 (O_3322,N_28045,N_27267);
or UO_3323 (O_3323,N_26923,N_26753);
nor UO_3324 (O_3324,N_26145,N_25634);
xnor UO_3325 (O_3325,N_26188,N_29214);
nor UO_3326 (O_3326,N_27232,N_29547);
nor UO_3327 (O_3327,N_24143,N_29018);
or UO_3328 (O_3328,N_25955,N_27514);
and UO_3329 (O_3329,N_29587,N_27060);
nor UO_3330 (O_3330,N_26860,N_25322);
or UO_3331 (O_3331,N_26639,N_29767);
nand UO_3332 (O_3332,N_25282,N_24131);
nor UO_3333 (O_3333,N_25125,N_29465);
nand UO_3334 (O_3334,N_28317,N_29718);
or UO_3335 (O_3335,N_29006,N_29699);
nand UO_3336 (O_3336,N_24455,N_29955);
and UO_3337 (O_3337,N_25432,N_28472);
nor UO_3338 (O_3338,N_29597,N_24936);
nand UO_3339 (O_3339,N_27862,N_27408);
nand UO_3340 (O_3340,N_28967,N_26122);
nor UO_3341 (O_3341,N_28604,N_26933);
nand UO_3342 (O_3342,N_28198,N_26118);
xnor UO_3343 (O_3343,N_27437,N_25373);
and UO_3344 (O_3344,N_24159,N_29741);
and UO_3345 (O_3345,N_29604,N_29531);
and UO_3346 (O_3346,N_29346,N_28758);
nand UO_3347 (O_3347,N_24577,N_27032);
and UO_3348 (O_3348,N_26642,N_27099);
and UO_3349 (O_3349,N_25152,N_26031);
and UO_3350 (O_3350,N_29662,N_24140);
and UO_3351 (O_3351,N_26354,N_27470);
xor UO_3352 (O_3352,N_29107,N_25200);
xnor UO_3353 (O_3353,N_29172,N_27779);
nand UO_3354 (O_3354,N_29501,N_27413);
or UO_3355 (O_3355,N_25211,N_29935);
nor UO_3356 (O_3356,N_25371,N_26192);
or UO_3357 (O_3357,N_24147,N_27400);
and UO_3358 (O_3358,N_24434,N_29502);
nand UO_3359 (O_3359,N_26618,N_24087);
and UO_3360 (O_3360,N_24248,N_29451);
or UO_3361 (O_3361,N_25028,N_27436);
and UO_3362 (O_3362,N_28087,N_26155);
xnor UO_3363 (O_3363,N_26961,N_25505);
or UO_3364 (O_3364,N_25822,N_25874);
xnor UO_3365 (O_3365,N_29951,N_25030);
and UO_3366 (O_3366,N_24737,N_24253);
xnor UO_3367 (O_3367,N_25417,N_24780);
and UO_3368 (O_3368,N_27406,N_25092);
and UO_3369 (O_3369,N_24420,N_25689);
or UO_3370 (O_3370,N_27504,N_29821);
xnor UO_3371 (O_3371,N_28018,N_27648);
or UO_3372 (O_3372,N_24262,N_24710);
nor UO_3373 (O_3373,N_25791,N_26809);
nand UO_3374 (O_3374,N_24860,N_27879);
nor UO_3375 (O_3375,N_29019,N_26317);
xnor UO_3376 (O_3376,N_24503,N_25752);
or UO_3377 (O_3377,N_29255,N_24193);
nand UO_3378 (O_3378,N_26649,N_26512);
or UO_3379 (O_3379,N_26878,N_29963);
xnor UO_3380 (O_3380,N_25844,N_26599);
nand UO_3381 (O_3381,N_27439,N_24972);
and UO_3382 (O_3382,N_27405,N_25796);
nand UO_3383 (O_3383,N_27979,N_28085);
or UO_3384 (O_3384,N_26611,N_26804);
or UO_3385 (O_3385,N_26479,N_24207);
xnor UO_3386 (O_3386,N_24860,N_26581);
and UO_3387 (O_3387,N_27181,N_28775);
and UO_3388 (O_3388,N_28017,N_24946);
nor UO_3389 (O_3389,N_26012,N_27364);
xnor UO_3390 (O_3390,N_27698,N_24841);
nand UO_3391 (O_3391,N_28112,N_26715);
and UO_3392 (O_3392,N_24014,N_26090);
xor UO_3393 (O_3393,N_24584,N_26181);
and UO_3394 (O_3394,N_29930,N_26516);
and UO_3395 (O_3395,N_29285,N_27359);
xnor UO_3396 (O_3396,N_26632,N_24415);
nor UO_3397 (O_3397,N_28872,N_24811);
nand UO_3398 (O_3398,N_29055,N_25604);
xnor UO_3399 (O_3399,N_24371,N_24871);
nand UO_3400 (O_3400,N_28699,N_29115);
nor UO_3401 (O_3401,N_24583,N_25293);
nor UO_3402 (O_3402,N_27942,N_29533);
and UO_3403 (O_3403,N_28344,N_29206);
or UO_3404 (O_3404,N_26104,N_27052);
and UO_3405 (O_3405,N_29112,N_28485);
nand UO_3406 (O_3406,N_26793,N_24131);
xnor UO_3407 (O_3407,N_25893,N_24382);
xnor UO_3408 (O_3408,N_25511,N_25903);
and UO_3409 (O_3409,N_29261,N_26563);
xor UO_3410 (O_3410,N_26989,N_29239);
nand UO_3411 (O_3411,N_27962,N_24662);
or UO_3412 (O_3412,N_28172,N_26355);
and UO_3413 (O_3413,N_25362,N_29822);
and UO_3414 (O_3414,N_24100,N_24072);
or UO_3415 (O_3415,N_29945,N_29275);
nor UO_3416 (O_3416,N_24055,N_24541);
nor UO_3417 (O_3417,N_25789,N_25687);
or UO_3418 (O_3418,N_28594,N_28569);
nand UO_3419 (O_3419,N_25653,N_26978);
or UO_3420 (O_3420,N_26978,N_25745);
and UO_3421 (O_3421,N_29449,N_24537);
xor UO_3422 (O_3422,N_25718,N_27768);
or UO_3423 (O_3423,N_26133,N_29441);
nor UO_3424 (O_3424,N_27296,N_29063);
and UO_3425 (O_3425,N_29244,N_25879);
or UO_3426 (O_3426,N_24681,N_28085);
xnor UO_3427 (O_3427,N_28876,N_24723);
or UO_3428 (O_3428,N_25286,N_27837);
nand UO_3429 (O_3429,N_25508,N_28204);
and UO_3430 (O_3430,N_25100,N_27052);
and UO_3431 (O_3431,N_28807,N_28453);
nor UO_3432 (O_3432,N_24096,N_29099);
xnor UO_3433 (O_3433,N_26217,N_26770);
nor UO_3434 (O_3434,N_28895,N_26776);
nand UO_3435 (O_3435,N_27181,N_26881);
and UO_3436 (O_3436,N_28992,N_25403);
xor UO_3437 (O_3437,N_24861,N_25945);
or UO_3438 (O_3438,N_29268,N_29018);
nor UO_3439 (O_3439,N_26400,N_25772);
and UO_3440 (O_3440,N_28743,N_25505);
or UO_3441 (O_3441,N_28318,N_28886);
nor UO_3442 (O_3442,N_27587,N_28472);
or UO_3443 (O_3443,N_25850,N_29234);
nand UO_3444 (O_3444,N_28040,N_25461);
nand UO_3445 (O_3445,N_27859,N_28485);
or UO_3446 (O_3446,N_24278,N_25940);
nand UO_3447 (O_3447,N_24459,N_26364);
and UO_3448 (O_3448,N_29922,N_29678);
nor UO_3449 (O_3449,N_26071,N_27005);
and UO_3450 (O_3450,N_26980,N_25997);
xor UO_3451 (O_3451,N_24516,N_26346);
xnor UO_3452 (O_3452,N_29112,N_26707);
nand UO_3453 (O_3453,N_26944,N_29704);
nand UO_3454 (O_3454,N_24787,N_27815);
and UO_3455 (O_3455,N_24984,N_24559);
nand UO_3456 (O_3456,N_26964,N_24243);
or UO_3457 (O_3457,N_27604,N_29485);
or UO_3458 (O_3458,N_24502,N_26451);
nand UO_3459 (O_3459,N_24332,N_25901);
and UO_3460 (O_3460,N_28195,N_29070);
nor UO_3461 (O_3461,N_29605,N_24889);
nor UO_3462 (O_3462,N_27919,N_25461);
xnor UO_3463 (O_3463,N_29684,N_27437);
or UO_3464 (O_3464,N_27117,N_25077);
or UO_3465 (O_3465,N_26770,N_27770);
and UO_3466 (O_3466,N_25342,N_25826);
or UO_3467 (O_3467,N_24045,N_29110);
and UO_3468 (O_3468,N_26282,N_29976);
and UO_3469 (O_3469,N_25549,N_28196);
nand UO_3470 (O_3470,N_25592,N_25470);
nor UO_3471 (O_3471,N_29183,N_28630);
xor UO_3472 (O_3472,N_25686,N_24210);
nor UO_3473 (O_3473,N_27343,N_24752);
or UO_3474 (O_3474,N_28350,N_24795);
xnor UO_3475 (O_3475,N_26820,N_27925);
xor UO_3476 (O_3476,N_26019,N_28678);
nor UO_3477 (O_3477,N_24094,N_28792);
or UO_3478 (O_3478,N_28641,N_27327);
nor UO_3479 (O_3479,N_29119,N_27427);
nor UO_3480 (O_3480,N_28714,N_26851);
xor UO_3481 (O_3481,N_28787,N_25572);
xor UO_3482 (O_3482,N_29177,N_25971);
and UO_3483 (O_3483,N_24624,N_28641);
nand UO_3484 (O_3484,N_29366,N_26563);
nor UO_3485 (O_3485,N_28726,N_24436);
nand UO_3486 (O_3486,N_26756,N_24152);
nand UO_3487 (O_3487,N_25471,N_26587);
xnor UO_3488 (O_3488,N_29660,N_26916);
nor UO_3489 (O_3489,N_25928,N_29519);
nor UO_3490 (O_3490,N_27733,N_29549);
and UO_3491 (O_3491,N_27198,N_25983);
nand UO_3492 (O_3492,N_27462,N_28674);
and UO_3493 (O_3493,N_27999,N_25599);
nor UO_3494 (O_3494,N_29710,N_26870);
nand UO_3495 (O_3495,N_28538,N_26415);
or UO_3496 (O_3496,N_28870,N_28969);
and UO_3497 (O_3497,N_25011,N_25759);
and UO_3498 (O_3498,N_24944,N_29943);
xor UO_3499 (O_3499,N_28589,N_26832);
endmodule