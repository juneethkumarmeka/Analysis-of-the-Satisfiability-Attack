module basic_2000_20000_2500_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1957,In_1544);
xor U1 (N_1,In_1240,In_332);
xnor U2 (N_2,In_1537,In_1701);
nand U3 (N_3,In_265,In_1505);
xnor U4 (N_4,In_1115,In_1777);
xor U5 (N_5,In_1885,In_1074);
nor U6 (N_6,In_1134,In_731);
nor U7 (N_7,In_1809,In_339);
xnor U8 (N_8,In_1439,In_1198);
xnor U9 (N_9,In_302,In_1990);
and U10 (N_10,In_1410,In_206);
or U11 (N_11,In_631,In_978);
nand U12 (N_12,In_659,In_506);
xor U13 (N_13,In_1652,In_1868);
nor U14 (N_14,In_859,In_1284);
nand U15 (N_15,In_1586,In_176);
xor U16 (N_16,In_1668,In_1994);
nor U17 (N_17,In_584,In_563);
nand U18 (N_18,In_359,In_855);
nor U19 (N_19,In_1760,In_1727);
and U20 (N_20,In_1566,In_1318);
xor U21 (N_21,In_1210,In_353);
and U22 (N_22,In_1008,In_536);
and U23 (N_23,In_883,In_1889);
xor U24 (N_24,In_1390,In_1817);
and U25 (N_25,In_1780,In_212);
xnor U26 (N_26,In_860,In_907);
and U27 (N_27,In_1445,In_1097);
nand U28 (N_28,In_1186,In_1419);
nand U29 (N_29,In_1144,In_692);
or U30 (N_30,In_1906,In_361);
nand U31 (N_31,In_834,In_1430);
nor U32 (N_32,In_1549,In_511);
nor U33 (N_33,In_1814,In_299);
nor U34 (N_34,In_981,In_1917);
xnor U35 (N_35,In_1570,In_86);
nand U36 (N_36,In_1355,In_1496);
and U37 (N_37,In_310,In_1995);
nand U38 (N_38,In_555,In_1781);
or U39 (N_39,In_533,In_1278);
nand U40 (N_40,In_451,In_1229);
nor U41 (N_41,In_923,In_235);
or U42 (N_42,In_1215,In_1317);
nand U43 (N_43,In_1993,In_226);
xnor U44 (N_44,In_598,In_131);
xnor U45 (N_45,In_843,In_1138);
nor U46 (N_46,In_1294,In_788);
xnor U47 (N_47,In_297,In_1477);
or U48 (N_48,In_79,In_266);
nor U49 (N_49,In_831,In_1293);
xor U50 (N_50,In_223,In_1821);
and U51 (N_51,In_626,In_3);
nor U52 (N_52,In_1107,In_190);
or U53 (N_53,In_1599,In_273);
nand U54 (N_54,In_1216,In_1203);
xor U55 (N_55,In_576,In_1458);
xnor U56 (N_56,In_1504,In_973);
nor U57 (N_57,In_1037,In_1704);
nor U58 (N_58,In_1258,In_930);
or U59 (N_59,In_957,In_1329);
nand U60 (N_60,In_1481,In_61);
nand U61 (N_61,In_524,In_360);
or U62 (N_62,In_16,In_368);
or U63 (N_63,In_459,In_1334);
nor U64 (N_64,In_586,In_1793);
or U65 (N_65,In_1673,In_1248);
and U66 (N_66,In_1232,In_1618);
xnor U67 (N_67,In_1971,In_1491);
xnor U68 (N_68,In_1040,In_285);
and U69 (N_69,In_162,In_307);
and U70 (N_70,In_1782,In_1071);
or U71 (N_71,In_349,In_160);
and U72 (N_72,In_750,In_1531);
or U73 (N_73,In_661,In_1576);
xnor U74 (N_74,In_1879,In_399);
or U75 (N_75,In_962,In_1579);
and U76 (N_76,In_658,In_1363);
nand U77 (N_77,In_1444,In_879);
and U78 (N_78,In_747,In_1436);
xnor U79 (N_79,In_1722,In_1041);
or U80 (N_80,In_1979,In_337);
nor U81 (N_81,In_1280,In_1195);
or U82 (N_82,In_249,In_1651);
and U83 (N_83,In_1453,In_400);
or U84 (N_84,In_1752,In_727);
nand U85 (N_85,In_327,In_836);
and U86 (N_86,In_677,In_84);
nand U87 (N_87,In_874,In_927);
and U88 (N_88,In_1913,In_352);
xnor U89 (N_89,In_968,In_113);
nand U90 (N_90,In_1922,In_1620);
nor U91 (N_91,In_581,In_1452);
xor U92 (N_92,In_293,In_1978);
and U93 (N_93,In_443,In_1540);
nor U94 (N_94,In_1724,In_1158);
xor U95 (N_95,In_1242,In_1762);
nand U96 (N_96,In_34,In_1102);
or U97 (N_97,In_292,In_1985);
nor U98 (N_98,In_1660,In_759);
and U99 (N_99,In_1154,In_758);
or U100 (N_100,In_838,In_1245);
and U101 (N_101,In_1842,In_276);
nand U102 (N_102,In_562,In_322);
or U103 (N_103,In_1779,In_1147);
nand U104 (N_104,In_440,In_699);
nor U105 (N_105,In_940,In_1698);
or U106 (N_106,In_100,In_1327);
and U107 (N_107,In_493,In_1970);
nor U108 (N_108,In_1328,In_189);
xnor U109 (N_109,In_766,In_1233);
and U110 (N_110,In_802,In_1636);
xor U111 (N_111,In_549,In_1870);
and U112 (N_112,In_1702,In_680);
nor U113 (N_113,In_1123,In_1918);
xnor U114 (N_114,In_1022,In_1079);
nand U115 (N_115,In_1563,In_575);
xor U116 (N_116,In_1498,In_1472);
xor U117 (N_117,In_577,In_167);
nor U118 (N_118,In_719,In_1713);
or U119 (N_119,In_247,In_1823);
nor U120 (N_120,In_535,In_1356);
xor U121 (N_121,In_350,In_77);
and U122 (N_122,In_743,In_1562);
or U123 (N_123,In_1470,In_1473);
and U124 (N_124,In_670,In_1737);
and U125 (N_125,In_1556,In_130);
nor U126 (N_126,In_599,In_45);
nor U127 (N_127,In_1499,In_1747);
nor U128 (N_128,In_73,In_509);
or U129 (N_129,In_881,In_1333);
nand U130 (N_130,In_1853,In_787);
xor U131 (N_131,In_1070,In_126);
xnor U132 (N_132,In_1068,In_1638);
nor U133 (N_133,In_229,In_119);
or U134 (N_134,In_354,In_1613);
xor U135 (N_135,In_1690,In_716);
nand U136 (N_136,In_539,In_984);
nand U137 (N_137,In_1083,In_1406);
nor U138 (N_138,In_282,In_983);
nor U139 (N_139,In_1016,In_1625);
and U140 (N_140,In_1207,In_711);
xor U141 (N_141,In_122,In_364);
nor U142 (N_142,In_965,In_1503);
or U143 (N_143,In_1302,In_343);
and U144 (N_144,In_288,In_889);
nor U145 (N_145,In_1886,In_305);
xnor U146 (N_146,In_455,In_156);
nand U147 (N_147,In_1986,In_414);
or U148 (N_148,In_1408,In_1188);
nor U149 (N_149,In_262,In_418);
and U150 (N_150,In_604,In_324);
nand U151 (N_151,In_830,In_1373);
nor U152 (N_152,In_268,In_919);
nor U153 (N_153,In_92,In_1916);
nand U154 (N_154,In_1682,In_1276);
nor U155 (N_155,In_1880,In_425);
or U156 (N_156,In_1301,In_1120);
xor U157 (N_157,In_633,In_817);
and U158 (N_158,In_939,In_308);
or U159 (N_159,In_908,In_1735);
nor U160 (N_160,In_1688,In_1623);
nand U161 (N_161,In_42,In_325);
xor U162 (N_162,In_1801,In_1536);
xor U163 (N_163,In_1253,In_173);
nand U164 (N_164,In_1377,In_500);
and U165 (N_165,In_39,In_538);
nand U166 (N_166,In_592,In_1768);
or U167 (N_167,In_1657,In_820);
or U168 (N_168,In_688,In_784);
or U169 (N_169,In_1644,In_1155);
or U170 (N_170,In_1681,In_1667);
or U171 (N_171,In_1105,In_1009);
nand U172 (N_172,In_1368,In_707);
and U173 (N_173,In_81,In_1897);
or U174 (N_174,In_24,In_1568);
xor U175 (N_175,In_1595,In_989);
nand U176 (N_176,In_526,In_776);
or U177 (N_177,In_291,In_95);
or U178 (N_178,In_281,In_1121);
nand U179 (N_179,In_452,In_579);
nand U180 (N_180,In_1739,In_1740);
nand U181 (N_181,In_503,In_1420);
nand U182 (N_182,In_1231,In_470);
nor U183 (N_183,In_1340,In_56);
nor U184 (N_184,In_1963,In_1849);
xor U185 (N_185,In_1583,In_1672);
nand U186 (N_186,In_1542,In_952);
or U187 (N_187,In_234,In_1422);
or U188 (N_188,In_306,In_208);
xor U189 (N_189,In_1012,In_1708);
xnor U190 (N_190,In_1087,In_1244);
or U191 (N_191,In_793,In_85);
and U192 (N_192,In_1141,In_1018);
or U193 (N_193,In_377,In_717);
nor U194 (N_194,In_1630,In_1414);
and U195 (N_195,In_313,In_1789);
nand U196 (N_196,In_821,In_611);
xnor U197 (N_197,In_1136,In_1127);
xor U198 (N_198,In_124,In_1733);
and U199 (N_199,In_147,In_431);
nand U200 (N_200,In_497,In_429);
and U201 (N_201,In_1157,In_567);
xnor U202 (N_202,In_1820,In_730);
and U203 (N_203,In_623,In_1602);
and U204 (N_204,In_605,In_72);
or U205 (N_205,In_1863,In_594);
and U206 (N_206,In_636,In_912);
xnor U207 (N_207,In_225,In_70);
xnor U208 (N_208,In_553,In_1310);
nand U209 (N_209,In_1146,In_315);
or U210 (N_210,In_734,In_329);
xor U211 (N_211,In_155,In_1940);
and U212 (N_212,In_1588,In_871);
nand U213 (N_213,In_1175,In_217);
nand U214 (N_214,In_620,In_774);
nand U215 (N_215,In_1714,In_1920);
nand U216 (N_216,In_182,In_681);
xor U217 (N_217,In_1129,In_667);
or U218 (N_218,In_1168,In_810);
nor U219 (N_219,In_1605,In_896);
nand U220 (N_220,In_1169,In_1749);
and U221 (N_221,In_1265,In_1560);
nor U222 (N_222,In_294,In_675);
xor U223 (N_223,In_1398,In_1217);
or U224 (N_224,In_238,In_78);
nor U225 (N_225,In_33,In_1559);
or U226 (N_226,In_71,In_852);
or U227 (N_227,In_150,In_1862);
nor U228 (N_228,In_1221,In_1174);
nor U229 (N_229,In_1696,In_906);
and U230 (N_230,In_15,In_1104);
or U231 (N_231,In_442,In_1639);
nor U232 (N_232,In_404,In_1488);
nand U233 (N_233,In_972,In_1263);
xnor U234 (N_234,In_1944,In_20);
xor U235 (N_235,In_1828,In_649);
or U236 (N_236,In_1236,In_1808);
or U237 (N_237,In_1791,In_1553);
or U238 (N_238,In_237,In_369);
xnor U239 (N_239,In_1839,In_746);
and U240 (N_240,In_1590,In_856);
nor U241 (N_241,In_1815,In_961);
or U242 (N_242,In_461,In_139);
nor U243 (N_243,In_284,In_1474);
xor U244 (N_244,In_1019,In_1227);
and U245 (N_245,In_997,In_1982);
nand U246 (N_246,In_1856,In_964);
or U247 (N_247,In_203,In_1836);
nand U248 (N_248,In_597,In_1500);
or U249 (N_249,In_1860,In_462);
xnor U250 (N_250,In_1561,In_1824);
xor U251 (N_251,In_1324,In_1440);
nor U252 (N_252,In_1335,In_1264);
nand U253 (N_253,In_260,In_1797);
or U254 (N_254,In_502,In_1988);
or U255 (N_255,In_1787,In_1023);
and U256 (N_256,In_1750,In_1521);
nand U257 (N_257,In_1254,In_481);
nor U258 (N_258,In_1058,In_1711);
xor U259 (N_259,In_1585,In_663);
or U260 (N_260,In_557,In_263);
and U261 (N_261,In_1366,In_19);
nand U262 (N_262,In_1725,In_1872);
xor U263 (N_263,In_1770,In_1530);
and U264 (N_264,In_1803,In_1984);
and U265 (N_265,In_1395,In_1790);
and U266 (N_266,In_1743,In_1734);
nor U267 (N_267,In_1364,In_1197);
nor U268 (N_268,In_127,In_791);
nor U269 (N_269,In_861,In_104);
xor U270 (N_270,In_648,In_777);
and U271 (N_271,In_1901,In_521);
nand U272 (N_272,In_862,In_753);
and U273 (N_273,In_1126,In_1788);
nand U274 (N_274,In_931,In_708);
or U275 (N_275,In_1180,In_1151);
xnor U276 (N_276,In_1048,In_606);
or U277 (N_277,In_1965,In_660);
xnor U278 (N_278,In_715,In_1748);
nor U279 (N_279,In_93,In_827);
xnor U280 (N_280,In_1628,In_546);
xnor U281 (N_281,In_995,In_705);
nor U282 (N_282,In_1816,In_600);
and U283 (N_283,In_1592,In_1035);
or U284 (N_284,In_1867,In_832);
and U285 (N_285,In_825,In_1225);
or U286 (N_286,In_635,In_1156);
xor U287 (N_287,In_388,In_517);
nand U288 (N_288,In_1109,In_1234);
and U289 (N_289,In_391,In_1581);
and U290 (N_290,In_565,In_1894);
and U291 (N_291,In_693,In_653);
nor U292 (N_292,In_1977,In_1832);
or U293 (N_293,In_488,In_1966);
and U294 (N_294,In_419,In_185);
nor U295 (N_295,In_1761,In_1947);
and U296 (N_296,In_573,In_18);
and U297 (N_297,In_69,In_1371);
xnor U298 (N_298,In_762,In_813);
xor U299 (N_299,In_1851,In_1831);
nor U300 (N_300,In_1285,In_897);
nor U301 (N_301,In_1376,In_650);
or U302 (N_302,In_240,In_1846);
xnor U303 (N_303,In_1066,In_1767);
nor U304 (N_304,In_1273,In_1053);
or U305 (N_305,In_1381,In_1999);
or U306 (N_306,In_654,In_566);
or U307 (N_307,In_27,In_890);
nand U308 (N_308,In_314,In_428);
and U309 (N_309,In_152,In_1418);
nand U310 (N_310,In_363,In_724);
or U311 (N_311,In_823,In_1962);
or U312 (N_312,In_1142,In_1635);
nand U313 (N_313,In_1929,In_105);
and U314 (N_314,In_950,In_1457);
nor U315 (N_315,In_1666,In_1312);
or U316 (N_316,In_1116,In_1818);
xor U317 (N_317,In_942,In_1766);
nor U318 (N_318,In_1380,In_424);
and U319 (N_319,In_1323,In_197);
or U320 (N_320,In_745,In_1359);
nand U321 (N_321,In_1061,In_1170);
nand U322 (N_322,In_910,In_14);
xnor U323 (N_323,In_1214,In_1833);
xor U324 (N_324,In_628,In_1172);
nand U325 (N_325,In_389,In_1044);
and U326 (N_326,In_239,In_1336);
or U327 (N_327,In_1425,In_1526);
or U328 (N_328,In_1547,In_1492);
or U329 (N_329,In_1098,In_687);
or U330 (N_330,In_1130,In_133);
nand U331 (N_331,In_172,In_1523);
xnor U332 (N_332,In_1572,In_1143);
xor U333 (N_333,In_1352,In_1091);
xnor U334 (N_334,In_1389,In_900);
nor U335 (N_335,In_800,In_1358);
or U336 (N_336,In_996,In_204);
xnor U337 (N_337,In_178,In_245);
and U338 (N_338,In_1677,In_454);
or U339 (N_339,In_1346,In_334);
or U340 (N_340,In_617,In_1813);
and U341 (N_341,In_191,In_1297);
and U342 (N_342,In_928,In_495);
or U343 (N_343,In_1490,In_578);
xor U344 (N_344,In_68,In_1065);
xnor U345 (N_345,In_679,In_1616);
xor U346 (N_346,In_619,In_607);
nand U347 (N_347,In_603,In_601);
nor U348 (N_348,In_1881,In_1517);
and U349 (N_349,In_1938,In_902);
and U350 (N_350,In_1026,In_1369);
nand U351 (N_351,In_484,In_312);
and U352 (N_352,In_1153,In_755);
xnor U353 (N_353,In_241,In_1348);
xnor U354 (N_354,In_188,In_463);
and U355 (N_355,In_1096,In_1004);
nand U356 (N_356,In_209,In_955);
nor U357 (N_357,In_174,In_102);
nor U358 (N_358,In_621,In_602);
or U359 (N_359,In_228,In_271);
nand U360 (N_360,In_1594,In_1837);
xor U361 (N_361,In_406,In_1307);
nand U362 (N_362,In_1942,In_1875);
and U363 (N_363,In_1838,In_394);
or U364 (N_364,In_729,In_783);
xor U365 (N_365,In_1309,In_1006);
nor U366 (N_366,In_770,In_28);
or U367 (N_367,In_1235,In_59);
xor U368 (N_368,In_351,In_445);
xor U369 (N_369,In_1896,In_819);
nand U370 (N_370,In_111,In_316);
and U371 (N_371,In_494,In_1511);
or U372 (N_372,In_709,In_1683);
and U373 (N_373,In_1279,In_151);
and U374 (N_374,In_686,In_88);
nor U375 (N_375,In_21,In_103);
or U376 (N_376,In_630,In_1039);
nor U377 (N_377,In_1912,In_595);
nand U378 (N_378,In_159,In_118);
and U379 (N_379,In_1438,In_924);
nand U380 (N_380,In_1241,In_519);
xnor U381 (N_381,In_574,In_1956);
xnor U382 (N_382,In_227,In_64);
nor U383 (N_383,In_1150,In_1139);
nor U384 (N_384,In_275,In_1397);
nand U385 (N_385,In_1367,In_466);
xor U386 (N_386,In_264,In_1567);
nand U387 (N_387,In_330,In_67);
xor U388 (N_388,In_1795,In_1306);
and U389 (N_389,In_1758,In_1357);
or U390 (N_390,In_1101,In_1303);
nor U391 (N_391,In_618,In_572);
nand U392 (N_392,In_1784,In_387);
and U393 (N_393,In_725,In_1753);
nand U394 (N_394,In_846,In_358);
and U395 (N_395,In_547,In_1953);
nand U396 (N_396,In_1205,In_640);
xnor U397 (N_397,In_742,In_1194);
nor U398 (N_398,In_1421,In_1786);
or U399 (N_399,In_971,In_1718);
or U400 (N_400,In_804,In_1140);
nand U401 (N_401,In_1338,In_1300);
xor U402 (N_402,In_1384,In_1314);
nor U403 (N_403,In_1372,In_5);
and U404 (N_404,In_1036,In_435);
and U405 (N_405,In_1100,In_175);
nand U406 (N_406,In_1428,In_1259);
nand U407 (N_407,In_1122,In_769);
nor U408 (N_408,In_714,In_427);
and U409 (N_409,In_829,In_1654);
nand U410 (N_410,In_1196,In_485);
xor U411 (N_411,In_878,In_588);
nand U412 (N_412,In_1876,In_1250);
xnor U413 (N_413,In_1723,In_1665);
or U414 (N_414,In_137,In_967);
or U415 (N_415,In_1295,In_1270);
xnor U416 (N_416,In_1024,In_1810);
nand U417 (N_417,In_1484,In_1843);
nor U418 (N_418,In_416,In_785);
and U419 (N_419,In_1238,In_401);
and U420 (N_420,In_438,In_624);
and U421 (N_421,In_977,In_544);
and U422 (N_422,In_1399,In_1528);
and U423 (N_423,In_183,In_884);
or U424 (N_424,In_918,In_483);
xnor U425 (N_425,In_664,In_1013);
nor U426 (N_426,In_976,In_13);
nor U427 (N_427,In_559,In_885);
and U428 (N_428,In_158,In_380);
nor U429 (N_429,In_1007,In_458);
nand U430 (N_430,In_356,In_1936);
nand U431 (N_431,In_953,In_789);
nand U432 (N_432,In_430,In_921);
nand U433 (N_433,In_157,In_1742);
and U434 (N_434,In_1633,In_279);
nand U435 (N_435,In_1441,In_37);
and U436 (N_436,In_477,In_1337);
or U437 (N_437,In_556,In_1057);
and U438 (N_438,In_1516,In_710);
nor U439 (N_439,In_876,In_1471);
nand U440 (N_440,In_1951,In_641);
nand U441 (N_441,In_946,In_523);
nand U442 (N_442,In_627,In_943);
nand U443 (N_443,In_32,In_1981);
xor U444 (N_444,In_722,In_1111);
xor U445 (N_445,In_1805,In_213);
and U446 (N_446,In_165,In_1765);
and U447 (N_447,In_145,In_933);
xor U448 (N_448,In_537,In_917);
xor U449 (N_449,In_672,In_1908);
nand U450 (N_450,In_1755,In_1883);
and U451 (N_451,In_589,In_1432);
and U452 (N_452,In_1538,In_1514);
nor U453 (N_453,In_1510,In_1525);
nand U454 (N_454,In_858,In_1968);
and U455 (N_455,In_1298,In_765);
nand U456 (N_456,In_925,In_1974);
and U457 (N_457,In_2,In_1365);
nand U458 (N_458,In_696,In_1859);
nor U459 (N_459,In_242,In_1165);
and U460 (N_460,In_844,In_25);
xor U461 (N_461,In_1051,In_1463);
nor U462 (N_462,In_583,In_491);
nand U463 (N_463,In_1550,In_453);
nor U464 (N_464,In_920,In_1220);
or U465 (N_465,In_1653,In_1532);
and U466 (N_466,In_1078,In_1596);
nor U467 (N_467,In_405,In_1417);
and U468 (N_468,In_1774,In_1326);
nand U469 (N_469,In_259,In_935);
or U470 (N_470,In_1729,In_1494);
xor U471 (N_471,In_1485,In_1189);
nor U472 (N_472,In_340,In_398);
and U473 (N_473,In_1032,In_1331);
xnor U474 (N_474,In_616,In_773);
and U475 (N_475,In_1513,In_433);
nand U476 (N_476,In_1060,In_1449);
nor U477 (N_477,In_593,In_170);
xor U478 (N_478,In_916,In_6);
xor U479 (N_479,In_1015,In_210);
and U480 (N_480,In_36,In_1475);
xnor U481 (N_481,In_1476,In_1631);
or U482 (N_482,In_694,In_1267);
xnor U483 (N_483,In_1448,In_975);
nor U484 (N_484,In_1315,In_1923);
nand U485 (N_485,In_525,In_872);
and U486 (N_486,In_468,In_1607);
or U487 (N_487,In_437,In_1900);
and U488 (N_488,In_796,In_1822);
and U489 (N_489,In_1268,In_196);
or U490 (N_490,In_1429,In_1899);
and U491 (N_491,In_300,In_501);
xnor U492 (N_492,In_1756,In_840);
xor U493 (N_493,In_1558,In_963);
nand U494 (N_494,In_1159,In_1002);
xor U495 (N_495,In_610,In_736);
nor U496 (N_496,In_657,In_90);
nand U497 (N_497,In_1728,In_409);
nor U498 (N_498,In_1396,In_1663);
nand U499 (N_499,In_1686,In_274);
xnor U500 (N_500,In_744,In_9);
nand U501 (N_501,In_1861,In_637);
nor U502 (N_502,In_1311,In_1112);
nor U503 (N_503,In_1459,In_1073);
xor U504 (N_504,In_1261,In_1997);
nand U505 (N_505,In_1726,In_1387);
nor U506 (N_506,In_551,In_141);
xnor U507 (N_507,In_768,In_1705);
nor U508 (N_508,In_1769,In_512);
and U509 (N_509,In_8,In_591);
nand U510 (N_510,In_934,In_63);
nand U511 (N_511,In_4,In_396);
xnor U512 (N_512,In_1462,In_1000);
nand U513 (N_513,In_450,In_666);
nand U514 (N_514,In_1684,In_1132);
nand U515 (N_515,In_1160,In_941);
and U516 (N_516,In_83,In_1489);
or U517 (N_517,In_761,In_1577);
or U518 (N_518,In_201,In_1687);
nand U519 (N_519,In_898,In_473);
and U520 (N_520,In_230,In_1152);
nor U521 (N_521,In_480,In_1252);
or U522 (N_522,In_1075,In_1502);
nand U523 (N_523,In_1845,In_342);
nor U524 (N_524,In_423,In_1678);
nand U525 (N_525,In_187,In_1800);
and U526 (N_526,In_1928,In_991);
xor U527 (N_527,In_1092,In_988);
nor U528 (N_528,In_718,In_1296);
or U529 (N_529,In_1179,In_1247);
or U530 (N_530,In_1052,In_1598);
or U531 (N_531,In_1394,In_257);
nor U532 (N_532,In_1290,In_1939);
nand U533 (N_533,In_780,In_1110);
or U534 (N_534,In_842,In_854);
or U535 (N_535,In_1676,In_571);
nand U536 (N_536,In_1289,In_1719);
xnor U537 (N_537,In_936,In_1834);
nand U538 (N_538,In_1266,In_94);
and U539 (N_539,In_1877,In_1757);
and U540 (N_540,In_1930,In_1308);
xor U541 (N_541,In_662,In_298);
nand U542 (N_542,In_146,In_1520);
or U543 (N_543,In_1148,In_469);
xor U544 (N_544,In_1771,In_1063);
nand U545 (N_545,In_134,In_508);
xor U546 (N_546,In_311,In_875);
nand U547 (N_547,In_1802,In_1089);
or U548 (N_548,In_1325,In_1622);
or U549 (N_549,In_1647,In_214);
or U550 (N_550,In_1534,In_254);
nand U551 (N_551,In_1171,In_937);
nor U552 (N_552,In_471,In_1487);
nor U553 (N_553,In_1855,In_514);
xnor U554 (N_554,In_895,In_1183);
and U555 (N_555,In_622,In_1555);
nor U556 (N_556,In_1891,In_10);
nand U557 (N_557,In_1996,In_614);
nor U558 (N_558,In_1949,In_179);
or U559 (N_559,In_1679,In_763);
xor U560 (N_560,In_956,In_1641);
nand U561 (N_561,In_893,In_395);
nand U562 (N_562,In_96,In_1621);
or U563 (N_563,In_1385,In_1330);
xnor U564 (N_564,In_48,In_570);
or U565 (N_565,In_911,In_1648);
nor U566 (N_566,In_982,In_140);
and U567 (N_567,In_1321,In_1269);
and U568 (N_568,In_1017,In_1460);
or U569 (N_569,In_74,In_582);
xor U570 (N_570,In_1543,In_1082);
nand U571 (N_571,In_712,In_397);
nand U572 (N_572,In_193,In_1580);
nor U573 (N_573,In_1292,In_1745);
xnor U574 (N_574,In_1131,In_1578);
nand U575 (N_575,In_865,In_1149);
nand U576 (N_576,In_1694,In_1626);
xnor U577 (N_577,In_1712,In_1405);
nand U578 (N_578,In_732,In_23);
nand U579 (N_579,In_1468,In_1050);
or U580 (N_580,In_913,In_1840);
and U581 (N_581,In_1461,In_548);
nand U582 (N_582,In_1339,In_1415);
xor U583 (N_583,In_510,In_120);
xor U584 (N_584,In_1099,In_674);
and U585 (N_585,In_993,In_1119);
nor U586 (N_586,In_690,In_1721);
nor U587 (N_587,In_1030,In_901);
and U588 (N_588,In_252,In_945);
or U589 (N_589,In_1424,In_702);
nand U590 (N_590,In_1167,In_221);
nor U591 (N_591,In_1858,In_642);
and U592 (N_592,In_1427,In_467);
nor U593 (N_593,In_1176,In_1);
nor U594 (N_594,In_905,In_1969);
or U595 (N_595,In_985,In_698);
nand U596 (N_596,In_1084,In_1360);
xor U597 (N_597,In_587,In_1045);
and U598 (N_598,In_949,In_771);
nand U599 (N_599,In_1222,In_1569);
xor U600 (N_600,In_366,In_951);
nand U601 (N_601,In_1118,In_371);
nand U602 (N_602,In_128,In_1844);
or U603 (N_603,In_720,In_1031);
or U604 (N_604,In_1529,In_180);
or U605 (N_605,In_1034,In_775);
xnor U606 (N_606,In_1691,In_478);
nor U607 (N_607,In_248,In_489);
nor U608 (N_608,In_1905,In_1201);
xnor U609 (N_609,In_457,In_1926);
or U610 (N_610,In_1509,In_43);
nand U611 (N_611,In_1043,In_1643);
nand U612 (N_612,In_415,In_319);
nor U613 (N_613,In_1975,In_1709);
xnor U614 (N_614,In_1890,In_323);
nor U615 (N_615,In_1237,In_749);
or U616 (N_616,In_1014,In_1888);
xor U617 (N_617,In_1190,In_805);
or U618 (N_618,In_689,In_1316);
nor U619 (N_619,In_1640,In_560);
and U620 (N_620,In_116,In_1403);
or U621 (N_621,In_1114,In_513);
nand U622 (N_622,In_1533,In_669);
nor U623 (N_623,In_222,In_1804);
nor U624 (N_624,In_1230,In_184);
xor U625 (N_625,In_256,In_1442);
xor U626 (N_626,In_1893,In_652);
nand U627 (N_627,In_1806,In_381);
or U628 (N_628,In_1857,In_82);
nor U629 (N_629,In_384,In_1869);
xor U630 (N_630,In_434,In_1072);
and U631 (N_631,In_1703,In_1882);
xor U632 (N_632,In_1286,In_11);
and U633 (N_633,In_1206,In_772);
nor U634 (N_634,In_969,In_612);
or U635 (N_635,In_283,In_1961);
xnor U636 (N_636,In_1163,In_1483);
xor U637 (N_637,In_472,In_199);
and U638 (N_638,In_695,In_1907);
or U639 (N_639,In_1632,In_46);
and U640 (N_640,In_1671,In_1224);
nor U641 (N_641,In_795,In_166);
xor U642 (N_642,In_161,In_833);
nor U643 (N_643,In_1211,In_1412);
and U644 (N_644,In_764,In_99);
nand U645 (N_645,In_841,In_751);
nand U646 (N_646,In_290,In_346);
nand U647 (N_647,In_338,In_1674);
xnor U648 (N_648,In_1850,In_168);
xnor U649 (N_649,In_1256,In_101);
xor U650 (N_650,In_1645,In_1927);
xnor U651 (N_651,In_849,In_164);
nor U652 (N_652,In_1934,In_863);
nor U653 (N_653,In_1305,In_1914);
nand U654 (N_654,In_613,In_320);
or U655 (N_655,In_194,In_947);
nor U656 (N_656,In_1069,In_704);
and U657 (N_657,In_1778,In_1539);
and U658 (N_658,In_80,In_421);
nand U659 (N_659,In_125,In_987);
nand U660 (N_660,In_1873,In_706);
or U661 (N_661,In_1212,In_1950);
nor U662 (N_662,In_1164,In_723);
xnor U663 (N_663,In_375,In_891);
nand U664 (N_664,In_420,In_596);
or U665 (N_665,In_236,In_171);
xnor U666 (N_666,In_870,In_1407);
nand U667 (N_667,In_107,In_1973);
nor U668 (N_668,In_108,In_839);
and U669 (N_669,In_1178,In_1741);
nand U670 (N_670,In_824,In_873);
nand U671 (N_671,In_656,In_1124);
nand U672 (N_672,In_1895,In_867);
nor U673 (N_673,In_685,In_1085);
nand U674 (N_674,In_808,In_1716);
and U675 (N_675,In_899,In_30);
nand U676 (N_676,In_866,In_1108);
and U677 (N_677,In_149,In_60);
or U678 (N_678,In_446,In_1299);
xor U679 (N_679,In_1067,In_1670);
nand U680 (N_680,In_1600,In_1960);
nor U681 (N_681,In_1662,In_1464);
and U682 (N_682,In_1388,In_417);
nand U683 (N_683,In_1161,In_738);
xor U684 (N_684,In_721,In_1541);
nand U685 (N_685,In_561,In_1557);
and U686 (N_686,In_143,In_278);
nor U687 (N_687,In_816,In_1606);
nor U688 (N_688,In_309,In_385);
and U689 (N_689,In_317,In_1386);
nand U690 (N_690,In_98,In_938);
nand U691 (N_691,In_782,In_1379);
or U692 (N_692,In_1847,In_1257);
and U693 (N_693,In_1958,In_1255);
and U694 (N_694,In_379,In_38);
and U695 (N_695,In_1411,In_1251);
nand U696 (N_696,In_1362,In_944);
xor U697 (N_697,In_136,In_1038);
nor U698 (N_698,In_531,In_643);
nand U699 (N_699,In_1699,In_1706);
nor U700 (N_700,In_1759,In_392);
and U701 (N_701,In_1482,In_1608);
nand U702 (N_702,In_1864,In_154);
nor U703 (N_703,In_568,In_1564);
nand U704 (N_704,In_413,In_106);
xor U705 (N_705,In_914,In_1402);
nor U706 (N_706,In_794,In_528);
or U707 (N_707,In_1937,In_1954);
or U708 (N_708,In_673,In_12);
or U709 (N_709,In_1401,In_1943);
or U710 (N_710,In_726,In_1903);
and U711 (N_711,In_1413,In_684);
or U712 (N_712,In_1952,In_1835);
nor U713 (N_713,In_786,In_703);
or U714 (N_714,In_91,In_518);
nor U715 (N_715,In_651,In_1056);
or U716 (N_716,In_1451,In_550);
and U717 (N_717,In_22,In_1046);
and U718 (N_718,In_757,In_748);
nand U719 (N_719,In_713,In_1054);
and U720 (N_720,In_1825,In_894);
nand U721 (N_721,In_1811,In_1349);
and U722 (N_722,In_545,In_847);
nor U723 (N_723,In_1746,In_296);
nor U724 (N_724,In_1799,In_809);
xor U725 (N_725,In_1456,In_1426);
or U726 (N_726,In_534,In_287);
xor U727 (N_727,In_1546,In_1772);
and U728 (N_728,In_1001,In_1497);
nand U729 (N_729,In_378,In_1343);
xor U730 (N_730,In_1522,In_1898);
xnor U731 (N_731,In_1219,In_382);
nor U732 (N_732,In_1033,In_1697);
xnor U733 (N_733,In_57,In_1524);
nor U734 (N_734,In_778,In_752);
nand U735 (N_735,In_691,In_701);
and U736 (N_736,In_932,In_682);
nor U737 (N_737,In_1059,In_1493);
and U738 (N_738,In_625,In_65);
or U739 (N_739,In_244,In_1935);
nand U740 (N_740,In_135,In_1117);
or U741 (N_741,In_348,In_1027);
nand U742 (N_742,In_376,In_1223);
and U743 (N_743,In_552,In_1573);
nor U744 (N_744,In_474,In_218);
and U745 (N_745,In_233,In_286);
nor U746 (N_746,In_1103,In_114);
or U747 (N_747,In_1827,In_1361);
nand U748 (N_748,In_163,In_1187);
and U749 (N_749,In_1466,In_632);
xor U750 (N_750,In_515,In_1593);
nand U751 (N_751,In_1707,In_115);
nand U752 (N_752,In_529,In_410);
nand U753 (N_753,In_869,In_1955);
nor U754 (N_754,In_1715,In_639);
nor U755 (N_755,In_644,In_1518);
nand U756 (N_756,In_1551,In_960);
nor U757 (N_757,In_357,In_877);
xnor U758 (N_758,In_1736,In_1508);
nand U759 (N_759,In_1400,In_798);
and U760 (N_760,In_41,In_1288);
nor U761 (N_761,In_1661,In_1437);
nand U762 (N_762,In_50,In_365);
nand U763 (N_763,In_1382,In_1617);
nor U764 (N_764,In_1611,In_1246);
and U765 (N_765,In_1610,In_1304);
or U766 (N_766,In_1945,In_1931);
nand U767 (N_767,In_564,In_1785);
nand U768 (N_768,In_522,In_970);
nand U769 (N_769,In_1775,In_558);
nor U770 (N_770,In_1319,In_1347);
xor U771 (N_771,In_1932,In_1341);
and U772 (N_772,In_1933,In_456);
nor U773 (N_773,In_487,In_1731);
xor U774 (N_774,In_1005,In_1848);
nor U775 (N_775,In_1910,In_29);
nor U776 (N_776,In_1627,In_1047);
nor U777 (N_777,In_0,In_781);
and U778 (N_778,In_1077,In_1807);
xnor U779 (N_779,In_507,In_1011);
or U780 (N_780,In_1064,In_1552);
nand U781 (N_781,In_1967,In_1450);
or U782 (N_782,In_251,In_1271);
nor U783 (N_783,In_295,In_1987);
nor U784 (N_784,In_1480,In_1375);
or U785 (N_785,In_1313,In_1744);
xnor U786 (N_786,In_492,In_1689);
or U787 (N_787,In_1878,In_1991);
nand U788 (N_788,In_1865,In_1275);
or U789 (N_789,In_1650,In_1055);
and U790 (N_790,In_540,In_460);
or U791 (N_791,In_1792,In_1609);
nor U792 (N_792,In_215,In_580);
nand U793 (N_793,In_1423,In_926);
and U794 (N_794,In_345,In_737);
nor U795 (N_795,In_207,In_1416);
and U796 (N_796,In_1911,In_475);
nand U797 (N_797,In_1656,In_1614);
nand U798 (N_798,In_615,In_1003);
xor U799 (N_799,In_634,In_129);
nor U800 (N_800,In_326,In_1919);
xor U801 (N_801,In_1946,In_1925);
nand U802 (N_802,In_1446,In_882);
and U803 (N_803,In_1983,In_390);
xnor U804 (N_804,In_1776,In_205);
and U805 (N_805,In_246,In_1637);
xnor U806 (N_806,In_328,In_756);
xor U807 (N_807,In_144,In_1332);
and U808 (N_808,In_1433,In_1584);
and U809 (N_809,In_697,In_498);
xnor U810 (N_810,In_35,In_992);
nand U811 (N_811,In_1717,In_1972);
nor U812 (N_812,In_422,In_958);
nand U813 (N_813,In_887,In_1921);
or U814 (N_814,In_811,In_1200);
nor U815 (N_815,In_1272,In_123);
and U816 (N_816,In_1571,In_1479);
nor U817 (N_817,In_1852,In_1353);
nor U818 (N_818,In_303,In_1020);
and U819 (N_819,In_504,In_321);
or U820 (N_820,In_1213,In_845);
nand U821 (N_821,In_826,In_52);
nor U822 (N_822,In_1128,In_1658);
and U823 (N_823,In_1454,In_1764);
nor U824 (N_824,In_1655,In_1826);
nand U825 (N_825,In_1841,In_1094);
nor U826 (N_826,In_231,In_948);
nand U827 (N_827,In_383,In_1763);
nor U828 (N_828,In_426,In_1080);
and U829 (N_829,In_1320,In_1209);
nand U830 (N_830,In_17,In_289);
nand U831 (N_831,In_886,In_1992);
nand U832 (N_832,In_1989,In_1021);
and U833 (N_833,In_1535,In_1204);
or U834 (N_834,In_97,In_1182);
nand U835 (N_835,In_700,In_676);
nand U836 (N_836,In_1391,In_1486);
xnor U837 (N_837,In_272,In_1730);
nand U838 (N_838,In_432,In_110);
xor U839 (N_839,In_754,In_465);
and U840 (N_840,In_444,In_1612);
xnor U841 (N_841,In_220,In_915);
xnor U842 (N_842,In_341,In_412);
xnor U843 (N_843,In_888,In_646);
nor U844 (N_844,In_1345,In_797);
or U845 (N_845,In_1948,In_966);
or U846 (N_846,In_590,In_31);
and U847 (N_847,In_1695,In_505);
or U848 (N_848,In_733,In_232);
nor U849 (N_849,In_1495,In_998);
or U850 (N_850,In_903,In_1909);
nand U851 (N_851,In_1393,In_1469);
or U852 (N_852,In_922,In_301);
nand U853 (N_853,In_402,In_1192);
and U854 (N_854,In_1344,In_954);
nand U855 (N_855,In_647,In_261);
or U856 (N_856,In_1202,In_1512);
nor U857 (N_857,In_270,In_54);
nand U858 (N_858,In_569,In_1354);
nor U859 (N_859,In_55,In_1964);
xnor U860 (N_860,In_543,In_479);
nand U861 (N_861,In_1693,In_1941);
nand U862 (N_862,In_441,In_608);
and U863 (N_863,In_1601,In_267);
or U864 (N_864,In_1049,In_386);
nand U865 (N_865,In_1819,In_40);
and U866 (N_866,In_1591,In_1738);
nand U867 (N_867,In_250,In_408);
or U868 (N_868,In_1404,In_851);
nor U869 (N_869,In_224,In_779);
or U870 (N_870,In_344,In_1025);
or U871 (N_871,In_58,In_1871);
xor U872 (N_872,In_464,In_1587);
or U873 (N_873,In_258,In_986);
nor U874 (N_874,In_857,In_1283);
and U875 (N_875,In_304,In_1904);
nand U876 (N_876,In_269,In_1081);
nor U877 (N_877,In_148,In_1434);
xor U878 (N_878,In_585,In_1249);
nand U879 (N_879,In_665,In_1199);
nor U880 (N_880,In_1754,In_1392);
xnor U881 (N_881,In_1646,In_436);
nand U882 (N_882,In_1642,In_1076);
nor U883 (N_883,In_198,In_541);
xnor U884 (N_884,In_448,In_999);
or U885 (N_885,In_1976,In_219);
nand U886 (N_886,In_1603,In_959);
xor U887 (N_887,In_1383,In_1409);
nand U888 (N_888,In_1575,In_818);
nor U889 (N_889,In_142,In_1443);
nand U890 (N_890,In_372,In_1515);
nor U891 (N_891,In_1435,In_1243);
and U892 (N_892,In_1548,In_336);
nand U893 (N_893,In_1629,In_1342);
and U894 (N_894,In_407,In_799);
or U895 (N_895,In_1277,In_49);
nand U896 (N_896,In_807,In_1680);
or U897 (N_897,In_1664,In_76);
xor U898 (N_898,In_1260,In_1892);
and U899 (N_899,In_476,In_1924);
nand U900 (N_900,In_1604,In_1884);
xor U901 (N_901,In_1378,In_814);
and U902 (N_902,In_1874,In_850);
nor U903 (N_903,In_1113,In_1507);
nand U904 (N_904,In_904,In_1565);
nand U905 (N_905,In_1135,In_121);
nand U906 (N_906,In_1854,In_1322);
or U907 (N_907,In_1137,In_994);
xor U908 (N_908,In_169,In_1262);
nor U909 (N_909,In_192,In_51);
or U910 (N_910,In_554,In_1088);
nand U911 (N_911,In_801,In_89);
nand U912 (N_912,In_211,In_1184);
nor U913 (N_913,In_47,In_741);
nand U914 (N_914,In_880,In_132);
xnor U915 (N_915,In_1794,In_837);
nand U916 (N_916,In_496,In_1720);
nand U917 (N_917,In_1239,In_370);
and U918 (N_918,In_44,In_1287);
and U919 (N_919,In_1431,In_835);
and U920 (N_920,In_66,In_112);
nor U921 (N_921,In_815,In_1998);
nand U922 (N_922,In_1959,In_806);
xor U923 (N_923,In_1042,In_75);
and U924 (N_924,In_767,In_1634);
and U925 (N_925,In_1185,In_1181);
nor U926 (N_926,In_929,In_1812);
xnor U927 (N_927,In_1291,In_740);
nand U928 (N_928,In_542,In_1783);
or U929 (N_929,In_1597,In_87);
and U930 (N_930,In_490,In_1028);
or U931 (N_931,In_1465,In_792);
nand U932 (N_932,In_530,In_1582);
and U933 (N_933,In_449,In_1351);
xor U934 (N_934,In_373,In_181);
nand U935 (N_935,In_1095,In_974);
xor U936 (N_936,In_678,In_195);
or U937 (N_937,In_1615,In_683);
or U938 (N_938,In_26,In_1455);
xor U939 (N_939,In_1350,In_109);
nor U940 (N_940,In_318,In_1830);
or U941 (N_941,In_1700,In_516);
or U942 (N_942,In_760,In_186);
nand U943 (N_943,In_1191,In_1685);
xor U944 (N_944,In_1796,In_1829);
nor U945 (N_945,In_1010,In_980);
xor U946 (N_946,In_1649,In_868);
nand U947 (N_947,In_482,In_892);
nand U948 (N_948,In_1086,In_1062);
nor U949 (N_949,In_1208,In_979);
xnor U950 (N_950,In_645,In_1282);
nor U951 (N_951,In_1659,In_671);
nand U952 (N_952,In_1980,In_803);
xnor U953 (N_953,In_739,In_1370);
nor U954 (N_954,In_62,In_447);
and U955 (N_955,In_335,In_1374);
nand U956 (N_956,In_7,In_1274);
and U957 (N_957,In_848,In_1177);
and U958 (N_958,In_1619,In_138);
nor U959 (N_959,In_277,In_117);
nand U960 (N_960,In_864,In_1866);
nor U961 (N_961,In_790,In_1106);
or U962 (N_962,In_1090,In_202);
nor U963 (N_963,In_486,In_243);
xnor U964 (N_964,In_1527,In_216);
nor U965 (N_965,In_53,In_668);
nand U966 (N_966,In_1193,In_1589);
and U967 (N_967,In_331,In_1166);
and U968 (N_968,In_1029,In_367);
nand U969 (N_969,In_499,In_1773);
xnor U970 (N_970,In_200,In_1478);
nor U971 (N_971,In_439,In_1162);
or U972 (N_972,In_1226,In_280);
xnor U973 (N_973,In_1751,In_1732);
or U974 (N_974,In_909,In_1218);
and U975 (N_975,In_638,In_1467);
nand U976 (N_976,In_177,In_520);
nor U977 (N_977,In_1506,In_1501);
xor U978 (N_978,In_853,In_355);
and U979 (N_979,In_153,In_374);
nand U980 (N_980,In_828,In_655);
or U981 (N_981,In_347,In_1093);
and U982 (N_982,In_393,In_1710);
nand U983 (N_983,In_362,In_1675);
xnor U984 (N_984,In_1519,In_1545);
or U985 (N_985,In_728,In_1133);
or U986 (N_986,In_532,In_1173);
xnor U987 (N_987,In_629,In_1145);
or U988 (N_988,In_1574,In_1692);
xnor U989 (N_989,In_990,In_822);
nand U990 (N_990,In_735,In_1554);
or U991 (N_991,In_253,In_1447);
or U992 (N_992,In_255,In_1125);
nand U993 (N_993,In_1228,In_1669);
xor U994 (N_994,In_411,In_1281);
and U995 (N_995,In_1624,In_1887);
nand U996 (N_996,In_1902,In_1915);
xnor U997 (N_997,In_333,In_403);
nor U998 (N_998,In_1798,In_812);
or U999 (N_999,In_527,In_609);
nand U1000 (N_1000,In_1537,In_1885);
nor U1001 (N_1001,In_1855,In_1978);
nor U1002 (N_1002,In_1975,In_286);
nor U1003 (N_1003,In_1312,In_1695);
and U1004 (N_1004,In_455,In_1053);
or U1005 (N_1005,In_1500,In_1374);
nor U1006 (N_1006,In_256,In_542);
or U1007 (N_1007,In_1658,In_806);
xor U1008 (N_1008,In_827,In_239);
nor U1009 (N_1009,In_298,In_1314);
nand U1010 (N_1010,In_1192,In_1017);
nor U1011 (N_1011,In_1331,In_345);
or U1012 (N_1012,In_1007,In_1332);
and U1013 (N_1013,In_459,In_1085);
xor U1014 (N_1014,In_734,In_1459);
xor U1015 (N_1015,In_1012,In_1923);
xor U1016 (N_1016,In_368,In_1925);
nand U1017 (N_1017,In_1846,In_1558);
nor U1018 (N_1018,In_1944,In_1031);
xnor U1019 (N_1019,In_745,In_570);
or U1020 (N_1020,In_772,In_245);
nand U1021 (N_1021,In_1706,In_213);
and U1022 (N_1022,In_1555,In_148);
or U1023 (N_1023,In_1964,In_1818);
or U1024 (N_1024,In_4,In_1052);
nand U1025 (N_1025,In_1042,In_1555);
nor U1026 (N_1026,In_1843,In_754);
nor U1027 (N_1027,In_1733,In_468);
or U1028 (N_1028,In_359,In_1408);
nand U1029 (N_1029,In_94,In_568);
xnor U1030 (N_1030,In_487,In_64);
nand U1031 (N_1031,In_1715,In_304);
nor U1032 (N_1032,In_154,In_116);
xnor U1033 (N_1033,In_1602,In_605);
or U1034 (N_1034,In_484,In_1205);
xor U1035 (N_1035,In_1600,In_1337);
nand U1036 (N_1036,In_82,In_968);
nor U1037 (N_1037,In_945,In_973);
and U1038 (N_1038,In_1108,In_1592);
xnor U1039 (N_1039,In_1323,In_1722);
and U1040 (N_1040,In_50,In_1272);
nor U1041 (N_1041,In_1039,In_1280);
nand U1042 (N_1042,In_772,In_67);
xor U1043 (N_1043,In_411,In_517);
xor U1044 (N_1044,In_1451,In_1492);
xnor U1045 (N_1045,In_1919,In_938);
nand U1046 (N_1046,In_1328,In_1591);
or U1047 (N_1047,In_1973,In_1468);
nor U1048 (N_1048,In_632,In_104);
or U1049 (N_1049,In_1434,In_606);
xnor U1050 (N_1050,In_1103,In_295);
xnor U1051 (N_1051,In_1288,In_161);
and U1052 (N_1052,In_761,In_638);
nor U1053 (N_1053,In_667,In_86);
xnor U1054 (N_1054,In_1817,In_1732);
and U1055 (N_1055,In_158,In_1312);
xnor U1056 (N_1056,In_1219,In_1683);
nor U1057 (N_1057,In_682,In_1156);
or U1058 (N_1058,In_1558,In_1832);
xnor U1059 (N_1059,In_1240,In_1574);
nor U1060 (N_1060,In_759,In_1079);
xnor U1061 (N_1061,In_557,In_1951);
and U1062 (N_1062,In_419,In_1816);
nor U1063 (N_1063,In_400,In_523);
nor U1064 (N_1064,In_1802,In_533);
nor U1065 (N_1065,In_1571,In_1471);
nand U1066 (N_1066,In_1437,In_71);
nor U1067 (N_1067,In_1742,In_1985);
nand U1068 (N_1068,In_981,In_1433);
nand U1069 (N_1069,In_893,In_1592);
and U1070 (N_1070,In_1181,In_1159);
or U1071 (N_1071,In_724,In_63);
xnor U1072 (N_1072,In_421,In_1323);
and U1073 (N_1073,In_362,In_1226);
or U1074 (N_1074,In_675,In_1507);
nor U1075 (N_1075,In_414,In_1872);
nor U1076 (N_1076,In_277,In_389);
xor U1077 (N_1077,In_44,In_404);
xor U1078 (N_1078,In_1699,In_1);
xor U1079 (N_1079,In_381,In_1503);
xnor U1080 (N_1080,In_1005,In_299);
nor U1081 (N_1081,In_51,In_830);
or U1082 (N_1082,In_1510,In_342);
nor U1083 (N_1083,In_1801,In_969);
and U1084 (N_1084,In_1423,In_542);
and U1085 (N_1085,In_561,In_1134);
and U1086 (N_1086,In_1228,In_1306);
nor U1087 (N_1087,In_1136,In_1093);
nand U1088 (N_1088,In_906,In_1161);
nand U1089 (N_1089,In_276,In_1434);
xor U1090 (N_1090,In_1769,In_629);
or U1091 (N_1091,In_1724,In_1057);
xnor U1092 (N_1092,In_1559,In_230);
or U1093 (N_1093,In_1335,In_890);
nand U1094 (N_1094,In_1181,In_527);
or U1095 (N_1095,In_399,In_1565);
nor U1096 (N_1096,In_1890,In_376);
and U1097 (N_1097,In_950,In_46);
nand U1098 (N_1098,In_1888,In_626);
and U1099 (N_1099,In_1322,In_1998);
nor U1100 (N_1100,In_362,In_1450);
nor U1101 (N_1101,In_835,In_711);
or U1102 (N_1102,In_1784,In_344);
and U1103 (N_1103,In_256,In_90);
nor U1104 (N_1104,In_1548,In_806);
xnor U1105 (N_1105,In_1263,In_1921);
or U1106 (N_1106,In_1489,In_860);
and U1107 (N_1107,In_990,In_442);
and U1108 (N_1108,In_1776,In_1070);
xor U1109 (N_1109,In_282,In_732);
or U1110 (N_1110,In_405,In_763);
nor U1111 (N_1111,In_1077,In_1107);
or U1112 (N_1112,In_310,In_663);
nor U1113 (N_1113,In_766,In_1004);
xnor U1114 (N_1114,In_3,In_572);
and U1115 (N_1115,In_1107,In_140);
nor U1116 (N_1116,In_292,In_1742);
or U1117 (N_1117,In_959,In_1700);
nand U1118 (N_1118,In_1960,In_753);
nor U1119 (N_1119,In_226,In_867);
or U1120 (N_1120,In_626,In_313);
xor U1121 (N_1121,In_634,In_172);
xnor U1122 (N_1122,In_955,In_444);
and U1123 (N_1123,In_937,In_401);
nor U1124 (N_1124,In_1118,In_31);
or U1125 (N_1125,In_1006,In_1960);
or U1126 (N_1126,In_1517,In_1021);
and U1127 (N_1127,In_500,In_636);
and U1128 (N_1128,In_1955,In_1298);
xor U1129 (N_1129,In_1598,In_1225);
nand U1130 (N_1130,In_1656,In_570);
or U1131 (N_1131,In_1184,In_1596);
nand U1132 (N_1132,In_649,In_703);
and U1133 (N_1133,In_1150,In_1746);
and U1134 (N_1134,In_1448,In_1283);
or U1135 (N_1135,In_849,In_55);
xor U1136 (N_1136,In_845,In_20);
nor U1137 (N_1137,In_843,In_572);
and U1138 (N_1138,In_1816,In_676);
and U1139 (N_1139,In_1144,In_502);
nor U1140 (N_1140,In_1553,In_1264);
xnor U1141 (N_1141,In_1623,In_415);
or U1142 (N_1142,In_360,In_423);
or U1143 (N_1143,In_165,In_908);
xor U1144 (N_1144,In_920,In_4);
or U1145 (N_1145,In_1094,In_1892);
and U1146 (N_1146,In_7,In_1448);
xor U1147 (N_1147,In_1466,In_1950);
xor U1148 (N_1148,In_792,In_1687);
nand U1149 (N_1149,In_1621,In_1549);
xnor U1150 (N_1150,In_1066,In_1463);
nand U1151 (N_1151,In_434,In_645);
nor U1152 (N_1152,In_1999,In_1899);
nor U1153 (N_1153,In_1170,In_937);
xnor U1154 (N_1154,In_652,In_489);
nand U1155 (N_1155,In_1858,In_863);
and U1156 (N_1156,In_766,In_1051);
and U1157 (N_1157,In_726,In_1426);
and U1158 (N_1158,In_1740,In_238);
and U1159 (N_1159,In_351,In_1389);
and U1160 (N_1160,In_155,In_727);
nand U1161 (N_1161,In_1420,In_1077);
xnor U1162 (N_1162,In_270,In_6);
nand U1163 (N_1163,In_804,In_1319);
or U1164 (N_1164,In_1676,In_1372);
and U1165 (N_1165,In_1126,In_687);
or U1166 (N_1166,In_1309,In_1596);
and U1167 (N_1167,In_921,In_1627);
or U1168 (N_1168,In_1263,In_459);
and U1169 (N_1169,In_1605,In_1004);
or U1170 (N_1170,In_31,In_913);
and U1171 (N_1171,In_28,In_1759);
and U1172 (N_1172,In_1708,In_1177);
nand U1173 (N_1173,In_281,In_374);
or U1174 (N_1174,In_372,In_1890);
nor U1175 (N_1175,In_275,In_588);
and U1176 (N_1176,In_870,In_295);
or U1177 (N_1177,In_123,In_1126);
nor U1178 (N_1178,In_905,In_191);
or U1179 (N_1179,In_1952,In_869);
nor U1180 (N_1180,In_639,In_1076);
xnor U1181 (N_1181,In_1348,In_768);
nor U1182 (N_1182,In_1353,In_280);
nor U1183 (N_1183,In_1211,In_1636);
nor U1184 (N_1184,In_486,In_1484);
or U1185 (N_1185,In_1174,In_847);
nand U1186 (N_1186,In_407,In_1551);
nand U1187 (N_1187,In_443,In_756);
xnor U1188 (N_1188,In_1921,In_1458);
nand U1189 (N_1189,In_1874,In_248);
or U1190 (N_1190,In_735,In_10);
nor U1191 (N_1191,In_80,In_1556);
nor U1192 (N_1192,In_1782,In_465);
nor U1193 (N_1193,In_1022,In_1347);
or U1194 (N_1194,In_19,In_189);
nor U1195 (N_1195,In_132,In_992);
nand U1196 (N_1196,In_297,In_1074);
nand U1197 (N_1197,In_1262,In_394);
or U1198 (N_1198,In_720,In_1153);
nor U1199 (N_1199,In_951,In_185);
xnor U1200 (N_1200,In_657,In_969);
nor U1201 (N_1201,In_119,In_1955);
or U1202 (N_1202,In_1522,In_610);
and U1203 (N_1203,In_1037,In_1635);
nor U1204 (N_1204,In_1105,In_1284);
xor U1205 (N_1205,In_444,In_1538);
xnor U1206 (N_1206,In_1293,In_315);
nand U1207 (N_1207,In_254,In_718);
and U1208 (N_1208,In_1879,In_482);
or U1209 (N_1209,In_1774,In_761);
nor U1210 (N_1210,In_1574,In_457);
and U1211 (N_1211,In_704,In_1998);
and U1212 (N_1212,In_215,In_485);
nand U1213 (N_1213,In_274,In_1799);
or U1214 (N_1214,In_1474,In_1478);
nor U1215 (N_1215,In_1945,In_1537);
xnor U1216 (N_1216,In_355,In_33);
xnor U1217 (N_1217,In_197,In_1833);
nand U1218 (N_1218,In_550,In_192);
or U1219 (N_1219,In_429,In_14);
nand U1220 (N_1220,In_132,In_394);
or U1221 (N_1221,In_1892,In_1956);
nor U1222 (N_1222,In_575,In_66);
or U1223 (N_1223,In_659,In_164);
or U1224 (N_1224,In_701,In_782);
or U1225 (N_1225,In_465,In_638);
nor U1226 (N_1226,In_1343,In_1199);
xor U1227 (N_1227,In_1158,In_1750);
and U1228 (N_1228,In_100,In_1298);
nor U1229 (N_1229,In_1806,In_1653);
and U1230 (N_1230,In_1620,In_1955);
and U1231 (N_1231,In_683,In_1877);
or U1232 (N_1232,In_1315,In_1706);
nand U1233 (N_1233,In_1078,In_377);
or U1234 (N_1234,In_117,In_1541);
and U1235 (N_1235,In_556,In_764);
xnor U1236 (N_1236,In_420,In_837);
and U1237 (N_1237,In_617,In_807);
or U1238 (N_1238,In_578,In_1481);
or U1239 (N_1239,In_1636,In_412);
xnor U1240 (N_1240,In_1985,In_737);
nand U1241 (N_1241,In_470,In_1809);
nand U1242 (N_1242,In_277,In_1818);
xnor U1243 (N_1243,In_663,In_799);
nor U1244 (N_1244,In_202,In_1532);
or U1245 (N_1245,In_1687,In_1888);
or U1246 (N_1246,In_834,In_1055);
nand U1247 (N_1247,In_1715,In_665);
nor U1248 (N_1248,In_1325,In_1018);
or U1249 (N_1249,In_1673,In_532);
nand U1250 (N_1250,In_780,In_426);
nor U1251 (N_1251,In_1625,In_1672);
or U1252 (N_1252,In_445,In_457);
nand U1253 (N_1253,In_1780,In_276);
xor U1254 (N_1254,In_861,In_1984);
nand U1255 (N_1255,In_1434,In_981);
and U1256 (N_1256,In_475,In_1055);
or U1257 (N_1257,In_1045,In_171);
nand U1258 (N_1258,In_1233,In_1319);
and U1259 (N_1259,In_1094,In_1531);
or U1260 (N_1260,In_652,In_363);
nor U1261 (N_1261,In_547,In_1741);
xor U1262 (N_1262,In_1398,In_1274);
or U1263 (N_1263,In_1875,In_1192);
nor U1264 (N_1264,In_1221,In_847);
nand U1265 (N_1265,In_708,In_1307);
nand U1266 (N_1266,In_486,In_307);
nor U1267 (N_1267,In_39,In_1656);
xnor U1268 (N_1268,In_588,In_180);
nor U1269 (N_1269,In_1383,In_1494);
xnor U1270 (N_1270,In_360,In_1920);
nand U1271 (N_1271,In_112,In_1875);
nor U1272 (N_1272,In_988,In_461);
or U1273 (N_1273,In_1979,In_699);
xnor U1274 (N_1274,In_1060,In_1965);
and U1275 (N_1275,In_1048,In_395);
or U1276 (N_1276,In_352,In_1419);
and U1277 (N_1277,In_934,In_333);
nand U1278 (N_1278,In_1859,In_1008);
nor U1279 (N_1279,In_805,In_1925);
or U1280 (N_1280,In_512,In_1096);
and U1281 (N_1281,In_1676,In_1863);
nor U1282 (N_1282,In_1029,In_12);
xor U1283 (N_1283,In_1805,In_1524);
nand U1284 (N_1284,In_916,In_1916);
nor U1285 (N_1285,In_1426,In_966);
and U1286 (N_1286,In_32,In_1594);
xnor U1287 (N_1287,In_750,In_296);
nor U1288 (N_1288,In_1277,In_467);
xnor U1289 (N_1289,In_334,In_1116);
xnor U1290 (N_1290,In_1844,In_1038);
nand U1291 (N_1291,In_1418,In_519);
nor U1292 (N_1292,In_923,In_45);
nor U1293 (N_1293,In_306,In_1749);
and U1294 (N_1294,In_352,In_1263);
xor U1295 (N_1295,In_238,In_673);
xor U1296 (N_1296,In_186,In_1650);
nand U1297 (N_1297,In_1386,In_351);
or U1298 (N_1298,In_1671,In_1864);
nor U1299 (N_1299,In_1151,In_1648);
nor U1300 (N_1300,In_1661,In_849);
nand U1301 (N_1301,In_1031,In_1517);
or U1302 (N_1302,In_133,In_1956);
nor U1303 (N_1303,In_367,In_1954);
or U1304 (N_1304,In_293,In_1385);
nor U1305 (N_1305,In_413,In_324);
xnor U1306 (N_1306,In_825,In_439);
nor U1307 (N_1307,In_1373,In_150);
xor U1308 (N_1308,In_382,In_1907);
xor U1309 (N_1309,In_625,In_419);
and U1310 (N_1310,In_609,In_1327);
or U1311 (N_1311,In_1288,In_1786);
or U1312 (N_1312,In_1522,In_1174);
xnor U1313 (N_1313,In_610,In_1438);
and U1314 (N_1314,In_1589,In_35);
xor U1315 (N_1315,In_1704,In_532);
and U1316 (N_1316,In_1520,In_1603);
nor U1317 (N_1317,In_568,In_542);
nor U1318 (N_1318,In_852,In_195);
nor U1319 (N_1319,In_1742,In_930);
and U1320 (N_1320,In_255,In_435);
nand U1321 (N_1321,In_216,In_6);
and U1322 (N_1322,In_1783,In_1657);
and U1323 (N_1323,In_790,In_245);
xnor U1324 (N_1324,In_898,In_1510);
xnor U1325 (N_1325,In_656,In_575);
xor U1326 (N_1326,In_1481,In_239);
nand U1327 (N_1327,In_1119,In_1620);
nor U1328 (N_1328,In_159,In_1447);
or U1329 (N_1329,In_654,In_1710);
xor U1330 (N_1330,In_154,In_1426);
and U1331 (N_1331,In_476,In_1234);
nand U1332 (N_1332,In_1108,In_663);
nand U1333 (N_1333,In_844,In_346);
or U1334 (N_1334,In_1594,In_262);
nand U1335 (N_1335,In_1141,In_1317);
nand U1336 (N_1336,In_1964,In_316);
nand U1337 (N_1337,In_659,In_1680);
and U1338 (N_1338,In_992,In_1789);
and U1339 (N_1339,In_474,In_121);
nor U1340 (N_1340,In_811,In_1775);
and U1341 (N_1341,In_1836,In_975);
nand U1342 (N_1342,In_156,In_190);
and U1343 (N_1343,In_734,In_1289);
xor U1344 (N_1344,In_1642,In_1936);
xnor U1345 (N_1345,In_1115,In_518);
and U1346 (N_1346,In_1626,In_911);
nand U1347 (N_1347,In_862,In_368);
and U1348 (N_1348,In_1575,In_1477);
or U1349 (N_1349,In_806,In_765);
nor U1350 (N_1350,In_859,In_562);
nor U1351 (N_1351,In_531,In_1854);
or U1352 (N_1352,In_506,In_1967);
and U1353 (N_1353,In_1772,In_462);
or U1354 (N_1354,In_97,In_594);
and U1355 (N_1355,In_1518,In_516);
or U1356 (N_1356,In_1614,In_82);
xnor U1357 (N_1357,In_188,In_16);
nor U1358 (N_1358,In_601,In_586);
or U1359 (N_1359,In_728,In_1899);
nor U1360 (N_1360,In_109,In_1629);
and U1361 (N_1361,In_1296,In_1150);
nand U1362 (N_1362,In_1797,In_1416);
or U1363 (N_1363,In_346,In_1143);
nor U1364 (N_1364,In_735,In_297);
and U1365 (N_1365,In_189,In_1669);
and U1366 (N_1366,In_1912,In_105);
nor U1367 (N_1367,In_308,In_385);
nor U1368 (N_1368,In_154,In_1395);
and U1369 (N_1369,In_1549,In_1490);
or U1370 (N_1370,In_1132,In_1213);
or U1371 (N_1371,In_1550,In_390);
or U1372 (N_1372,In_1790,In_1467);
nor U1373 (N_1373,In_550,In_1936);
xor U1374 (N_1374,In_807,In_972);
and U1375 (N_1375,In_603,In_1800);
nor U1376 (N_1376,In_655,In_1367);
and U1377 (N_1377,In_1112,In_714);
and U1378 (N_1378,In_1841,In_830);
and U1379 (N_1379,In_1187,In_1278);
xor U1380 (N_1380,In_178,In_1193);
nand U1381 (N_1381,In_1319,In_732);
xor U1382 (N_1382,In_1335,In_877);
and U1383 (N_1383,In_1871,In_873);
nor U1384 (N_1384,In_676,In_1742);
or U1385 (N_1385,In_599,In_89);
nor U1386 (N_1386,In_366,In_1453);
xnor U1387 (N_1387,In_1641,In_881);
or U1388 (N_1388,In_1592,In_1535);
nand U1389 (N_1389,In_406,In_1376);
or U1390 (N_1390,In_1797,In_1331);
or U1391 (N_1391,In_619,In_1321);
nand U1392 (N_1392,In_601,In_292);
xnor U1393 (N_1393,In_225,In_355);
and U1394 (N_1394,In_245,In_1102);
nor U1395 (N_1395,In_1512,In_1714);
nand U1396 (N_1396,In_826,In_583);
nor U1397 (N_1397,In_1205,In_1034);
nor U1398 (N_1398,In_814,In_1920);
nand U1399 (N_1399,In_1734,In_8);
nand U1400 (N_1400,In_1115,In_279);
nor U1401 (N_1401,In_982,In_570);
or U1402 (N_1402,In_1035,In_1378);
xor U1403 (N_1403,In_1619,In_457);
or U1404 (N_1404,In_165,In_1689);
or U1405 (N_1405,In_366,In_768);
xnor U1406 (N_1406,In_149,In_58);
nor U1407 (N_1407,In_553,In_1950);
nor U1408 (N_1408,In_1196,In_836);
nor U1409 (N_1409,In_1490,In_1844);
nor U1410 (N_1410,In_478,In_1892);
and U1411 (N_1411,In_1892,In_1975);
or U1412 (N_1412,In_1723,In_170);
nor U1413 (N_1413,In_686,In_292);
nor U1414 (N_1414,In_1762,In_1964);
xnor U1415 (N_1415,In_801,In_27);
nand U1416 (N_1416,In_1853,In_1507);
xor U1417 (N_1417,In_1544,In_714);
xor U1418 (N_1418,In_319,In_1241);
and U1419 (N_1419,In_1889,In_1750);
nand U1420 (N_1420,In_1663,In_208);
or U1421 (N_1421,In_1566,In_371);
and U1422 (N_1422,In_370,In_1097);
xor U1423 (N_1423,In_490,In_862);
nor U1424 (N_1424,In_1809,In_1291);
xnor U1425 (N_1425,In_1675,In_465);
or U1426 (N_1426,In_1328,In_1644);
or U1427 (N_1427,In_1570,In_1185);
xor U1428 (N_1428,In_1449,In_825);
xnor U1429 (N_1429,In_1195,In_993);
nand U1430 (N_1430,In_231,In_1051);
nor U1431 (N_1431,In_1159,In_1467);
nand U1432 (N_1432,In_278,In_86);
nand U1433 (N_1433,In_1633,In_1416);
and U1434 (N_1434,In_1258,In_169);
xor U1435 (N_1435,In_135,In_414);
nand U1436 (N_1436,In_1878,In_1927);
nand U1437 (N_1437,In_1145,In_521);
xnor U1438 (N_1438,In_1606,In_1987);
xnor U1439 (N_1439,In_649,In_1871);
and U1440 (N_1440,In_140,In_1001);
nor U1441 (N_1441,In_559,In_933);
nand U1442 (N_1442,In_54,In_1540);
and U1443 (N_1443,In_721,In_1806);
nor U1444 (N_1444,In_1905,In_1036);
nor U1445 (N_1445,In_483,In_1511);
or U1446 (N_1446,In_73,In_362);
nand U1447 (N_1447,In_788,In_214);
and U1448 (N_1448,In_1962,In_1553);
nor U1449 (N_1449,In_335,In_1364);
xnor U1450 (N_1450,In_1871,In_933);
or U1451 (N_1451,In_1913,In_1216);
xor U1452 (N_1452,In_1550,In_659);
xnor U1453 (N_1453,In_1460,In_1770);
nor U1454 (N_1454,In_706,In_149);
and U1455 (N_1455,In_786,In_155);
nand U1456 (N_1456,In_1120,In_248);
nor U1457 (N_1457,In_1541,In_1871);
nor U1458 (N_1458,In_1321,In_589);
or U1459 (N_1459,In_1138,In_613);
and U1460 (N_1460,In_1994,In_1173);
nand U1461 (N_1461,In_998,In_1237);
nor U1462 (N_1462,In_1111,In_87);
nor U1463 (N_1463,In_135,In_1153);
and U1464 (N_1464,In_499,In_1103);
nor U1465 (N_1465,In_608,In_1334);
xnor U1466 (N_1466,In_641,In_642);
xor U1467 (N_1467,In_251,In_1157);
xnor U1468 (N_1468,In_1119,In_1730);
xor U1469 (N_1469,In_941,In_888);
and U1470 (N_1470,In_1966,In_187);
nand U1471 (N_1471,In_134,In_1639);
and U1472 (N_1472,In_1713,In_1420);
and U1473 (N_1473,In_44,In_1542);
nand U1474 (N_1474,In_1816,In_225);
and U1475 (N_1475,In_1626,In_1723);
nand U1476 (N_1476,In_1677,In_272);
and U1477 (N_1477,In_1518,In_1996);
xor U1478 (N_1478,In_1845,In_1364);
or U1479 (N_1479,In_1168,In_865);
nand U1480 (N_1480,In_321,In_1906);
nor U1481 (N_1481,In_1038,In_407);
and U1482 (N_1482,In_1222,In_559);
and U1483 (N_1483,In_102,In_1332);
and U1484 (N_1484,In_1221,In_1661);
xor U1485 (N_1485,In_1674,In_1780);
or U1486 (N_1486,In_62,In_1526);
xnor U1487 (N_1487,In_901,In_837);
and U1488 (N_1488,In_1016,In_1910);
or U1489 (N_1489,In_1046,In_1940);
nor U1490 (N_1490,In_1164,In_540);
or U1491 (N_1491,In_1493,In_796);
and U1492 (N_1492,In_1870,In_1171);
and U1493 (N_1493,In_1200,In_104);
xor U1494 (N_1494,In_849,In_703);
xor U1495 (N_1495,In_1412,In_537);
or U1496 (N_1496,In_492,In_1047);
nor U1497 (N_1497,In_146,In_1369);
or U1498 (N_1498,In_110,In_756);
xnor U1499 (N_1499,In_1255,In_1691);
xnor U1500 (N_1500,In_1036,In_1399);
or U1501 (N_1501,In_1038,In_1661);
nor U1502 (N_1502,In_995,In_1271);
xnor U1503 (N_1503,In_214,In_170);
xor U1504 (N_1504,In_1413,In_183);
xnor U1505 (N_1505,In_1863,In_1260);
nand U1506 (N_1506,In_1241,In_1125);
xor U1507 (N_1507,In_540,In_141);
nor U1508 (N_1508,In_1795,In_1682);
nand U1509 (N_1509,In_1622,In_1392);
or U1510 (N_1510,In_1090,In_1034);
or U1511 (N_1511,In_475,In_1414);
xor U1512 (N_1512,In_1566,In_1393);
and U1513 (N_1513,In_148,In_1841);
nor U1514 (N_1514,In_1806,In_1885);
xor U1515 (N_1515,In_48,In_367);
and U1516 (N_1516,In_1494,In_1873);
xor U1517 (N_1517,In_21,In_1041);
or U1518 (N_1518,In_1239,In_1586);
nor U1519 (N_1519,In_222,In_1349);
xnor U1520 (N_1520,In_989,In_1739);
xor U1521 (N_1521,In_1255,In_400);
nand U1522 (N_1522,In_205,In_1186);
or U1523 (N_1523,In_1955,In_256);
or U1524 (N_1524,In_359,In_934);
xnor U1525 (N_1525,In_523,In_1855);
xor U1526 (N_1526,In_604,In_269);
and U1527 (N_1527,In_117,In_1762);
nor U1528 (N_1528,In_1728,In_523);
and U1529 (N_1529,In_1452,In_1308);
nand U1530 (N_1530,In_930,In_310);
nand U1531 (N_1531,In_518,In_1410);
nand U1532 (N_1532,In_88,In_1701);
xor U1533 (N_1533,In_1087,In_154);
nor U1534 (N_1534,In_192,In_105);
nand U1535 (N_1535,In_1021,In_1094);
nand U1536 (N_1536,In_436,In_1833);
xnor U1537 (N_1537,In_419,In_150);
and U1538 (N_1538,In_1079,In_299);
or U1539 (N_1539,In_804,In_1074);
or U1540 (N_1540,In_958,In_415);
xor U1541 (N_1541,In_1361,In_372);
or U1542 (N_1542,In_971,In_242);
and U1543 (N_1543,In_1038,In_779);
nand U1544 (N_1544,In_854,In_1357);
and U1545 (N_1545,In_215,In_493);
nor U1546 (N_1546,In_617,In_1096);
nand U1547 (N_1547,In_1796,In_1113);
or U1548 (N_1548,In_246,In_262);
or U1549 (N_1549,In_737,In_150);
or U1550 (N_1550,In_1115,In_170);
and U1551 (N_1551,In_1950,In_106);
and U1552 (N_1552,In_1741,In_1837);
nor U1553 (N_1553,In_250,In_1959);
and U1554 (N_1554,In_99,In_1412);
xor U1555 (N_1555,In_1083,In_163);
nor U1556 (N_1556,In_706,In_1215);
or U1557 (N_1557,In_828,In_1179);
nand U1558 (N_1558,In_566,In_213);
or U1559 (N_1559,In_1561,In_1062);
xor U1560 (N_1560,In_493,In_1181);
nor U1561 (N_1561,In_894,In_1403);
and U1562 (N_1562,In_1130,In_1957);
nand U1563 (N_1563,In_966,In_559);
nor U1564 (N_1564,In_1447,In_510);
and U1565 (N_1565,In_1966,In_1104);
xor U1566 (N_1566,In_1743,In_1198);
xor U1567 (N_1567,In_1624,In_910);
nor U1568 (N_1568,In_29,In_1144);
or U1569 (N_1569,In_381,In_616);
xnor U1570 (N_1570,In_1147,In_364);
nand U1571 (N_1571,In_557,In_1406);
xnor U1572 (N_1572,In_1063,In_1654);
and U1573 (N_1573,In_1404,In_55);
nand U1574 (N_1574,In_195,In_888);
or U1575 (N_1575,In_343,In_1280);
and U1576 (N_1576,In_1487,In_1852);
xor U1577 (N_1577,In_406,In_837);
nor U1578 (N_1578,In_1860,In_1384);
nand U1579 (N_1579,In_1341,In_1359);
xnor U1580 (N_1580,In_296,In_1763);
nor U1581 (N_1581,In_1544,In_1874);
xor U1582 (N_1582,In_1090,In_758);
nand U1583 (N_1583,In_1320,In_1237);
nor U1584 (N_1584,In_1237,In_368);
nor U1585 (N_1585,In_290,In_1073);
nand U1586 (N_1586,In_1786,In_1546);
xnor U1587 (N_1587,In_974,In_365);
and U1588 (N_1588,In_1948,In_676);
or U1589 (N_1589,In_624,In_1350);
or U1590 (N_1590,In_1342,In_1595);
xor U1591 (N_1591,In_1634,In_250);
nand U1592 (N_1592,In_1253,In_413);
or U1593 (N_1593,In_1965,In_609);
or U1594 (N_1594,In_1465,In_1700);
or U1595 (N_1595,In_1311,In_329);
xnor U1596 (N_1596,In_859,In_253);
and U1597 (N_1597,In_1594,In_904);
nor U1598 (N_1598,In_105,In_1527);
xor U1599 (N_1599,In_1457,In_1847);
nand U1600 (N_1600,In_1382,In_129);
or U1601 (N_1601,In_881,In_1035);
xor U1602 (N_1602,In_1760,In_1925);
or U1603 (N_1603,In_455,In_1313);
xnor U1604 (N_1604,In_1935,In_514);
or U1605 (N_1605,In_747,In_979);
and U1606 (N_1606,In_1982,In_681);
xnor U1607 (N_1607,In_1275,In_519);
nor U1608 (N_1608,In_1843,In_1207);
nor U1609 (N_1609,In_1214,In_1440);
or U1610 (N_1610,In_1578,In_990);
nor U1611 (N_1611,In_1918,In_588);
or U1612 (N_1612,In_1772,In_1323);
xor U1613 (N_1613,In_1024,In_1710);
and U1614 (N_1614,In_290,In_1876);
xnor U1615 (N_1615,In_821,In_1642);
nor U1616 (N_1616,In_706,In_1626);
and U1617 (N_1617,In_862,In_138);
or U1618 (N_1618,In_715,In_864);
xor U1619 (N_1619,In_251,In_341);
or U1620 (N_1620,In_764,In_746);
or U1621 (N_1621,In_1392,In_1142);
and U1622 (N_1622,In_743,In_1584);
or U1623 (N_1623,In_828,In_126);
and U1624 (N_1624,In_1417,In_1292);
or U1625 (N_1625,In_68,In_156);
nor U1626 (N_1626,In_1289,In_1856);
nor U1627 (N_1627,In_525,In_671);
or U1628 (N_1628,In_1896,In_1856);
and U1629 (N_1629,In_920,In_1671);
xor U1630 (N_1630,In_1406,In_304);
nand U1631 (N_1631,In_1334,In_824);
xor U1632 (N_1632,In_764,In_1216);
nor U1633 (N_1633,In_1433,In_983);
or U1634 (N_1634,In_1826,In_1124);
and U1635 (N_1635,In_309,In_1378);
xnor U1636 (N_1636,In_1317,In_1273);
xnor U1637 (N_1637,In_139,In_549);
nor U1638 (N_1638,In_702,In_214);
nor U1639 (N_1639,In_1738,In_1707);
nand U1640 (N_1640,In_1144,In_543);
and U1641 (N_1641,In_1407,In_1778);
or U1642 (N_1642,In_324,In_1046);
xnor U1643 (N_1643,In_872,In_318);
and U1644 (N_1644,In_944,In_1160);
nand U1645 (N_1645,In_266,In_83);
nand U1646 (N_1646,In_1913,In_1476);
nand U1647 (N_1647,In_874,In_1522);
and U1648 (N_1648,In_1224,In_263);
and U1649 (N_1649,In_497,In_955);
and U1650 (N_1650,In_262,In_1926);
and U1651 (N_1651,In_918,In_961);
nand U1652 (N_1652,In_396,In_667);
nor U1653 (N_1653,In_532,In_985);
or U1654 (N_1654,In_359,In_819);
nor U1655 (N_1655,In_939,In_886);
or U1656 (N_1656,In_1600,In_1235);
nand U1657 (N_1657,In_414,In_1747);
nor U1658 (N_1658,In_1927,In_1618);
nor U1659 (N_1659,In_1486,In_1937);
or U1660 (N_1660,In_1784,In_47);
xnor U1661 (N_1661,In_1593,In_161);
xor U1662 (N_1662,In_1453,In_1790);
nand U1663 (N_1663,In_832,In_742);
and U1664 (N_1664,In_839,In_40);
nor U1665 (N_1665,In_1796,In_276);
xor U1666 (N_1666,In_679,In_1948);
nor U1667 (N_1667,In_1249,In_1960);
nor U1668 (N_1668,In_1351,In_1443);
or U1669 (N_1669,In_1744,In_1492);
and U1670 (N_1670,In_378,In_1088);
or U1671 (N_1671,In_972,In_381);
and U1672 (N_1672,In_758,In_5);
nand U1673 (N_1673,In_1782,In_1946);
nor U1674 (N_1674,In_610,In_1778);
and U1675 (N_1675,In_1657,In_237);
nor U1676 (N_1676,In_1414,In_1642);
nand U1677 (N_1677,In_271,In_631);
xor U1678 (N_1678,In_1600,In_1453);
xnor U1679 (N_1679,In_1979,In_789);
nor U1680 (N_1680,In_407,In_1841);
or U1681 (N_1681,In_194,In_1124);
or U1682 (N_1682,In_914,In_189);
and U1683 (N_1683,In_985,In_186);
nor U1684 (N_1684,In_1103,In_1617);
or U1685 (N_1685,In_563,In_1416);
xnor U1686 (N_1686,In_1995,In_610);
xor U1687 (N_1687,In_1112,In_1786);
nor U1688 (N_1688,In_1835,In_567);
and U1689 (N_1689,In_52,In_474);
and U1690 (N_1690,In_1090,In_11);
or U1691 (N_1691,In_1844,In_1499);
xnor U1692 (N_1692,In_1961,In_982);
nand U1693 (N_1693,In_549,In_1703);
nand U1694 (N_1694,In_1287,In_214);
nand U1695 (N_1695,In_1969,In_1287);
nand U1696 (N_1696,In_129,In_1859);
nand U1697 (N_1697,In_227,In_288);
or U1698 (N_1698,In_178,In_401);
or U1699 (N_1699,In_684,In_1138);
nand U1700 (N_1700,In_1821,In_638);
or U1701 (N_1701,In_1200,In_358);
nand U1702 (N_1702,In_1633,In_1356);
and U1703 (N_1703,In_921,In_145);
xnor U1704 (N_1704,In_656,In_1855);
xnor U1705 (N_1705,In_1405,In_563);
and U1706 (N_1706,In_81,In_1035);
or U1707 (N_1707,In_1532,In_319);
nor U1708 (N_1708,In_684,In_569);
xnor U1709 (N_1709,In_16,In_1445);
nor U1710 (N_1710,In_135,In_180);
nor U1711 (N_1711,In_265,In_752);
nor U1712 (N_1712,In_1188,In_414);
and U1713 (N_1713,In_57,In_691);
nor U1714 (N_1714,In_1683,In_546);
nor U1715 (N_1715,In_654,In_1503);
nand U1716 (N_1716,In_1814,In_1673);
xor U1717 (N_1717,In_50,In_1115);
and U1718 (N_1718,In_9,In_350);
nand U1719 (N_1719,In_1470,In_1982);
or U1720 (N_1720,In_528,In_1511);
xnor U1721 (N_1721,In_1663,In_1853);
nand U1722 (N_1722,In_316,In_0);
xnor U1723 (N_1723,In_746,In_568);
xor U1724 (N_1724,In_1749,In_1167);
and U1725 (N_1725,In_435,In_918);
and U1726 (N_1726,In_488,In_863);
nand U1727 (N_1727,In_548,In_1656);
nand U1728 (N_1728,In_464,In_479);
nand U1729 (N_1729,In_225,In_1888);
nand U1730 (N_1730,In_1533,In_158);
or U1731 (N_1731,In_1229,In_358);
nand U1732 (N_1732,In_1367,In_98);
nor U1733 (N_1733,In_559,In_379);
and U1734 (N_1734,In_1038,In_1553);
xor U1735 (N_1735,In_413,In_959);
or U1736 (N_1736,In_1173,In_991);
and U1737 (N_1737,In_749,In_1313);
and U1738 (N_1738,In_1241,In_977);
xor U1739 (N_1739,In_1727,In_922);
and U1740 (N_1740,In_1462,In_1089);
or U1741 (N_1741,In_850,In_662);
and U1742 (N_1742,In_174,In_1678);
or U1743 (N_1743,In_568,In_1867);
and U1744 (N_1744,In_1977,In_856);
nor U1745 (N_1745,In_1794,In_240);
or U1746 (N_1746,In_915,In_37);
nand U1747 (N_1747,In_282,In_910);
and U1748 (N_1748,In_872,In_972);
or U1749 (N_1749,In_332,In_846);
xnor U1750 (N_1750,In_263,In_1820);
nand U1751 (N_1751,In_1094,In_1264);
nand U1752 (N_1752,In_1398,In_1919);
or U1753 (N_1753,In_89,In_374);
nand U1754 (N_1754,In_999,In_1639);
xor U1755 (N_1755,In_1185,In_673);
and U1756 (N_1756,In_650,In_494);
and U1757 (N_1757,In_1921,In_934);
nor U1758 (N_1758,In_642,In_1358);
nand U1759 (N_1759,In_722,In_455);
nand U1760 (N_1760,In_1375,In_562);
or U1761 (N_1761,In_493,In_992);
nand U1762 (N_1762,In_215,In_325);
xnor U1763 (N_1763,In_1710,In_1144);
nor U1764 (N_1764,In_676,In_1241);
xor U1765 (N_1765,In_582,In_641);
nand U1766 (N_1766,In_1576,In_378);
nand U1767 (N_1767,In_739,In_613);
and U1768 (N_1768,In_1863,In_1017);
xor U1769 (N_1769,In_5,In_714);
or U1770 (N_1770,In_818,In_1006);
or U1771 (N_1771,In_733,In_659);
and U1772 (N_1772,In_696,In_1930);
nand U1773 (N_1773,In_1282,In_1895);
or U1774 (N_1774,In_1889,In_367);
nand U1775 (N_1775,In_176,In_489);
nor U1776 (N_1776,In_1252,In_1679);
xnor U1777 (N_1777,In_175,In_407);
nor U1778 (N_1778,In_89,In_1356);
nor U1779 (N_1779,In_1093,In_1303);
nor U1780 (N_1780,In_380,In_1326);
nor U1781 (N_1781,In_1384,In_577);
nand U1782 (N_1782,In_1204,In_1873);
xnor U1783 (N_1783,In_744,In_226);
nand U1784 (N_1784,In_1218,In_263);
nor U1785 (N_1785,In_1500,In_1947);
xnor U1786 (N_1786,In_1984,In_1154);
xor U1787 (N_1787,In_1608,In_459);
nor U1788 (N_1788,In_323,In_741);
and U1789 (N_1789,In_641,In_828);
and U1790 (N_1790,In_26,In_1377);
xor U1791 (N_1791,In_1707,In_1669);
or U1792 (N_1792,In_548,In_324);
or U1793 (N_1793,In_880,In_1879);
or U1794 (N_1794,In_755,In_1131);
nand U1795 (N_1795,In_1766,In_691);
nor U1796 (N_1796,In_1588,In_1133);
nand U1797 (N_1797,In_1962,In_1083);
and U1798 (N_1798,In_805,In_178);
nor U1799 (N_1799,In_1370,In_223);
nor U1800 (N_1800,In_1424,In_896);
nor U1801 (N_1801,In_1359,In_284);
or U1802 (N_1802,In_1774,In_1662);
and U1803 (N_1803,In_954,In_196);
xor U1804 (N_1804,In_74,In_1906);
or U1805 (N_1805,In_1521,In_434);
nand U1806 (N_1806,In_63,In_1521);
or U1807 (N_1807,In_1591,In_44);
or U1808 (N_1808,In_1158,In_1471);
nand U1809 (N_1809,In_1886,In_1475);
and U1810 (N_1810,In_140,In_931);
and U1811 (N_1811,In_1651,In_1593);
and U1812 (N_1812,In_45,In_1712);
and U1813 (N_1813,In_419,In_1727);
nand U1814 (N_1814,In_1375,In_593);
or U1815 (N_1815,In_86,In_1353);
nor U1816 (N_1816,In_464,In_1698);
xor U1817 (N_1817,In_867,In_1887);
nor U1818 (N_1818,In_687,In_1140);
and U1819 (N_1819,In_556,In_961);
or U1820 (N_1820,In_1058,In_1364);
nor U1821 (N_1821,In_1271,In_1010);
or U1822 (N_1822,In_650,In_533);
xnor U1823 (N_1823,In_1395,In_1989);
nor U1824 (N_1824,In_824,In_882);
or U1825 (N_1825,In_1468,In_1032);
nor U1826 (N_1826,In_351,In_108);
and U1827 (N_1827,In_1354,In_1249);
xnor U1828 (N_1828,In_711,In_1276);
xor U1829 (N_1829,In_573,In_140);
and U1830 (N_1830,In_863,In_882);
nor U1831 (N_1831,In_1131,In_730);
nand U1832 (N_1832,In_662,In_149);
nand U1833 (N_1833,In_1105,In_1063);
or U1834 (N_1834,In_634,In_428);
nand U1835 (N_1835,In_812,In_1815);
xnor U1836 (N_1836,In_875,In_1281);
and U1837 (N_1837,In_498,In_1313);
or U1838 (N_1838,In_1714,In_1063);
xor U1839 (N_1839,In_1689,In_1214);
nand U1840 (N_1840,In_174,In_1755);
or U1841 (N_1841,In_980,In_831);
and U1842 (N_1842,In_1997,In_715);
xnor U1843 (N_1843,In_1961,In_578);
nand U1844 (N_1844,In_993,In_1333);
or U1845 (N_1845,In_1258,In_1011);
or U1846 (N_1846,In_989,In_83);
nor U1847 (N_1847,In_237,In_930);
and U1848 (N_1848,In_1570,In_739);
and U1849 (N_1849,In_1161,In_1717);
or U1850 (N_1850,In_1537,In_122);
nor U1851 (N_1851,In_1041,In_266);
or U1852 (N_1852,In_1106,In_594);
and U1853 (N_1853,In_1498,In_851);
nand U1854 (N_1854,In_1351,In_1385);
xnor U1855 (N_1855,In_48,In_1969);
or U1856 (N_1856,In_1663,In_1609);
or U1857 (N_1857,In_1369,In_468);
and U1858 (N_1858,In_727,In_1115);
and U1859 (N_1859,In_327,In_1958);
and U1860 (N_1860,In_1578,In_501);
and U1861 (N_1861,In_1822,In_253);
or U1862 (N_1862,In_68,In_1656);
nand U1863 (N_1863,In_1770,In_1637);
nand U1864 (N_1864,In_1949,In_1027);
xor U1865 (N_1865,In_1844,In_459);
and U1866 (N_1866,In_746,In_901);
xor U1867 (N_1867,In_1431,In_771);
and U1868 (N_1868,In_1843,In_966);
and U1869 (N_1869,In_883,In_191);
xnor U1870 (N_1870,In_1795,In_1314);
or U1871 (N_1871,In_1771,In_222);
nand U1872 (N_1872,In_355,In_1806);
nand U1873 (N_1873,In_1464,In_847);
nor U1874 (N_1874,In_1418,In_1333);
and U1875 (N_1875,In_1323,In_1166);
or U1876 (N_1876,In_410,In_22);
or U1877 (N_1877,In_116,In_882);
nor U1878 (N_1878,In_1609,In_774);
nand U1879 (N_1879,In_131,In_1926);
xnor U1880 (N_1880,In_498,In_1340);
nand U1881 (N_1881,In_1769,In_1013);
and U1882 (N_1882,In_1720,In_1539);
nor U1883 (N_1883,In_953,In_1998);
or U1884 (N_1884,In_1894,In_128);
nor U1885 (N_1885,In_1207,In_1475);
xor U1886 (N_1886,In_986,In_509);
nor U1887 (N_1887,In_1697,In_435);
xnor U1888 (N_1888,In_573,In_1640);
xor U1889 (N_1889,In_1966,In_1661);
xnor U1890 (N_1890,In_812,In_768);
nor U1891 (N_1891,In_579,In_901);
nor U1892 (N_1892,In_187,In_953);
nor U1893 (N_1893,In_934,In_1453);
or U1894 (N_1894,In_530,In_296);
or U1895 (N_1895,In_357,In_246);
xnor U1896 (N_1896,In_1762,In_682);
xnor U1897 (N_1897,In_1680,In_477);
and U1898 (N_1898,In_1616,In_497);
or U1899 (N_1899,In_1048,In_568);
or U1900 (N_1900,In_1248,In_819);
nand U1901 (N_1901,In_965,In_808);
nor U1902 (N_1902,In_1298,In_467);
nand U1903 (N_1903,In_194,In_1527);
and U1904 (N_1904,In_1973,In_232);
xor U1905 (N_1905,In_167,In_59);
and U1906 (N_1906,In_298,In_321);
nor U1907 (N_1907,In_1574,In_485);
nor U1908 (N_1908,In_1821,In_1181);
and U1909 (N_1909,In_1304,In_524);
nor U1910 (N_1910,In_653,In_451);
xor U1911 (N_1911,In_1284,In_760);
and U1912 (N_1912,In_770,In_1369);
nand U1913 (N_1913,In_720,In_641);
nor U1914 (N_1914,In_1291,In_1479);
and U1915 (N_1915,In_1934,In_786);
and U1916 (N_1916,In_1219,In_997);
or U1917 (N_1917,In_1420,In_1434);
xnor U1918 (N_1918,In_907,In_203);
nand U1919 (N_1919,In_124,In_478);
nor U1920 (N_1920,In_177,In_1338);
and U1921 (N_1921,In_134,In_479);
and U1922 (N_1922,In_877,In_1091);
or U1923 (N_1923,In_93,In_1044);
or U1924 (N_1924,In_925,In_794);
nand U1925 (N_1925,In_1574,In_945);
xnor U1926 (N_1926,In_473,In_454);
and U1927 (N_1927,In_413,In_1664);
or U1928 (N_1928,In_560,In_1914);
or U1929 (N_1929,In_346,In_1590);
nor U1930 (N_1930,In_127,In_1697);
or U1931 (N_1931,In_817,In_1251);
and U1932 (N_1932,In_1233,In_693);
nand U1933 (N_1933,In_1819,In_225);
nor U1934 (N_1934,In_1577,In_959);
nand U1935 (N_1935,In_795,In_1491);
or U1936 (N_1936,In_1462,In_1381);
and U1937 (N_1937,In_759,In_813);
or U1938 (N_1938,In_738,In_243);
xnor U1939 (N_1939,In_763,In_1866);
xor U1940 (N_1940,In_798,In_1179);
nor U1941 (N_1941,In_336,In_1279);
and U1942 (N_1942,In_532,In_1556);
or U1943 (N_1943,In_800,In_78);
nand U1944 (N_1944,In_1505,In_1720);
nand U1945 (N_1945,In_622,In_433);
or U1946 (N_1946,In_488,In_1833);
nor U1947 (N_1947,In_1421,In_1638);
and U1948 (N_1948,In_1015,In_1610);
nor U1949 (N_1949,In_1664,In_673);
nand U1950 (N_1950,In_1977,In_1621);
nand U1951 (N_1951,In_969,In_119);
or U1952 (N_1952,In_68,In_1281);
nand U1953 (N_1953,In_514,In_1806);
xnor U1954 (N_1954,In_645,In_1760);
xnor U1955 (N_1955,In_1717,In_474);
or U1956 (N_1956,In_764,In_1961);
or U1957 (N_1957,In_1396,In_799);
or U1958 (N_1958,In_138,In_1402);
nor U1959 (N_1959,In_404,In_1627);
or U1960 (N_1960,In_1624,In_797);
nand U1961 (N_1961,In_624,In_230);
or U1962 (N_1962,In_1621,In_305);
nor U1963 (N_1963,In_858,In_627);
or U1964 (N_1964,In_1450,In_1584);
or U1965 (N_1965,In_1620,In_1987);
nand U1966 (N_1966,In_124,In_1759);
nand U1967 (N_1967,In_1181,In_1089);
xnor U1968 (N_1968,In_1306,In_376);
nor U1969 (N_1969,In_1420,In_208);
nor U1970 (N_1970,In_1800,In_839);
nand U1971 (N_1971,In_1732,In_438);
xor U1972 (N_1972,In_1592,In_1496);
nand U1973 (N_1973,In_1203,In_438);
nor U1974 (N_1974,In_1648,In_182);
and U1975 (N_1975,In_511,In_925);
nand U1976 (N_1976,In_1718,In_1519);
nor U1977 (N_1977,In_1971,In_32);
and U1978 (N_1978,In_1629,In_171);
xnor U1979 (N_1979,In_1039,In_1452);
and U1980 (N_1980,In_124,In_121);
xor U1981 (N_1981,In_314,In_871);
xor U1982 (N_1982,In_564,In_1956);
nand U1983 (N_1983,In_1933,In_726);
nand U1984 (N_1984,In_1925,In_208);
nand U1985 (N_1985,In_122,In_1425);
nand U1986 (N_1986,In_1478,In_1100);
or U1987 (N_1987,In_554,In_1973);
xor U1988 (N_1988,In_1152,In_1669);
or U1989 (N_1989,In_162,In_138);
or U1990 (N_1990,In_706,In_1858);
nor U1991 (N_1991,In_1638,In_290);
and U1992 (N_1992,In_337,In_1392);
or U1993 (N_1993,In_1809,In_1991);
xor U1994 (N_1994,In_169,In_520);
nor U1995 (N_1995,In_273,In_575);
and U1996 (N_1996,In_301,In_1181);
and U1997 (N_1997,In_1689,In_1229);
or U1998 (N_1998,In_1531,In_617);
xnor U1999 (N_1999,In_1318,In_1375);
xnor U2000 (N_2000,N_813,N_1644);
nand U2001 (N_2001,N_242,N_144);
xnor U2002 (N_2002,N_771,N_1159);
nand U2003 (N_2003,N_1950,N_1322);
nor U2004 (N_2004,N_670,N_1015);
and U2005 (N_2005,N_1674,N_1711);
nor U2006 (N_2006,N_1925,N_1839);
or U2007 (N_2007,N_247,N_977);
or U2008 (N_2008,N_1891,N_1774);
or U2009 (N_2009,N_40,N_654);
or U2010 (N_2010,N_947,N_349);
or U2011 (N_2011,N_93,N_1107);
xnor U2012 (N_2012,N_1768,N_94);
nand U2013 (N_2013,N_1027,N_1135);
xor U2014 (N_2014,N_1100,N_24);
nor U2015 (N_2015,N_625,N_338);
and U2016 (N_2016,N_1084,N_1113);
nor U2017 (N_2017,N_1718,N_1779);
nand U2018 (N_2018,N_196,N_1974);
nor U2019 (N_2019,N_1985,N_36);
nand U2020 (N_2020,N_1365,N_846);
or U2021 (N_2021,N_1271,N_1907);
nor U2022 (N_2022,N_1241,N_1227);
and U2023 (N_2023,N_1225,N_1286);
xor U2024 (N_2024,N_32,N_1805);
nor U2025 (N_2025,N_1118,N_839);
xnor U2026 (N_2026,N_908,N_1369);
nand U2027 (N_2027,N_1445,N_1428);
nand U2028 (N_2028,N_1809,N_1359);
xnor U2029 (N_2029,N_1813,N_1494);
xor U2030 (N_2030,N_163,N_667);
and U2031 (N_2031,N_589,N_1512);
nand U2032 (N_2032,N_68,N_1206);
nand U2033 (N_2033,N_1513,N_460);
nand U2034 (N_2034,N_957,N_1811);
nand U2035 (N_2035,N_1753,N_1052);
xnor U2036 (N_2036,N_231,N_781);
or U2037 (N_2037,N_1914,N_1928);
xnor U2038 (N_2038,N_1977,N_1888);
nor U2039 (N_2039,N_619,N_282);
and U2040 (N_2040,N_77,N_1821);
nand U2041 (N_2041,N_427,N_7);
and U2042 (N_2042,N_1540,N_1059);
nor U2043 (N_2043,N_1122,N_1838);
or U2044 (N_2044,N_1128,N_1742);
nor U2045 (N_2045,N_284,N_1617);
nand U2046 (N_2046,N_882,N_565);
xor U2047 (N_2047,N_1012,N_835);
xnor U2048 (N_2048,N_216,N_689);
nor U2049 (N_2049,N_56,N_772);
or U2050 (N_2050,N_486,N_1406);
xor U2051 (N_2051,N_678,N_1333);
and U2052 (N_2052,N_1904,N_1381);
or U2053 (N_2053,N_1973,N_1851);
and U2054 (N_2054,N_9,N_1347);
and U2055 (N_2055,N_506,N_29);
nor U2056 (N_2056,N_1859,N_1345);
nand U2057 (N_2057,N_661,N_1475);
and U2058 (N_2058,N_1583,N_1498);
xnor U2059 (N_2059,N_1425,N_1987);
or U2060 (N_2060,N_645,N_1267);
nor U2061 (N_2061,N_1775,N_1873);
xnor U2062 (N_2062,N_1731,N_652);
nor U2063 (N_2063,N_1455,N_274);
or U2064 (N_2064,N_816,N_83);
nand U2065 (N_2065,N_1854,N_1575);
nand U2066 (N_2066,N_1554,N_27);
or U2067 (N_2067,N_564,N_159);
xor U2068 (N_2068,N_1087,N_491);
and U2069 (N_2069,N_1156,N_1899);
nand U2070 (N_2070,N_1000,N_1901);
nor U2071 (N_2071,N_770,N_1088);
and U2072 (N_2072,N_1185,N_122);
nor U2073 (N_2073,N_422,N_1641);
nand U2074 (N_2074,N_991,N_883);
nand U2075 (N_2075,N_579,N_861);
or U2076 (N_2076,N_191,N_243);
xnor U2077 (N_2077,N_1189,N_515);
or U2078 (N_2078,N_389,N_222);
xnor U2079 (N_2079,N_1092,N_1256);
xor U2080 (N_2080,N_86,N_1177);
xor U2081 (N_2081,N_692,N_1684);
or U2082 (N_2082,N_1618,N_71);
and U2083 (N_2083,N_1588,N_246);
xnor U2084 (N_2084,N_503,N_473);
and U2085 (N_2085,N_694,N_975);
or U2086 (N_2086,N_1566,N_370);
nand U2087 (N_2087,N_874,N_890);
or U2088 (N_2088,N_969,N_1221);
or U2089 (N_2089,N_853,N_1508);
nand U2090 (N_2090,N_948,N_1106);
and U2091 (N_2091,N_1294,N_236);
and U2092 (N_2092,N_1228,N_744);
and U2093 (N_2093,N_1665,N_1074);
nor U2094 (N_2094,N_562,N_604);
nor U2095 (N_2095,N_875,N_887);
nand U2096 (N_2096,N_1739,N_450);
nand U2097 (N_2097,N_1143,N_1034);
xor U2098 (N_2098,N_372,N_1968);
xnor U2099 (N_2099,N_444,N_691);
nand U2100 (N_2100,N_1023,N_1773);
nand U2101 (N_2101,N_1410,N_82);
or U2102 (N_2102,N_702,N_1491);
and U2103 (N_2103,N_843,N_171);
nand U2104 (N_2104,N_1929,N_149);
xor U2105 (N_2105,N_1824,N_714);
or U2106 (N_2106,N_307,N_886);
nor U2107 (N_2107,N_736,N_409);
nor U2108 (N_2108,N_1943,N_337);
xnor U2109 (N_2109,N_119,N_631);
nand U2110 (N_2110,N_1955,N_956);
or U2111 (N_2111,N_1252,N_1944);
or U2112 (N_2112,N_1981,N_452);
and U2113 (N_2113,N_34,N_1701);
xor U2114 (N_2114,N_1650,N_737);
or U2115 (N_2115,N_239,N_1536);
nand U2116 (N_2116,N_404,N_1876);
nor U2117 (N_2117,N_301,N_1963);
or U2118 (N_2118,N_799,N_1148);
and U2119 (N_2119,N_659,N_1523);
or U2120 (N_2120,N_1865,N_433);
and U2121 (N_2121,N_761,N_252);
and U2122 (N_2122,N_845,N_1780);
nor U2123 (N_2123,N_1833,N_273);
and U2124 (N_2124,N_1857,N_617);
nor U2125 (N_2125,N_1367,N_189);
or U2126 (N_2126,N_92,N_791);
xnor U2127 (N_2127,N_1200,N_1042);
nand U2128 (N_2128,N_1157,N_374);
or U2129 (N_2129,N_1817,N_276);
and U2130 (N_2130,N_219,N_1712);
nand U2131 (N_2131,N_148,N_440);
nand U2132 (N_2132,N_367,N_1026);
nor U2133 (N_2133,N_1037,N_576);
xnor U2134 (N_2134,N_1013,N_855);
or U2135 (N_2135,N_1884,N_1667);
nand U2136 (N_2136,N_660,N_129);
or U2137 (N_2137,N_1336,N_623);
xnor U2138 (N_2138,N_675,N_209);
and U2139 (N_2139,N_1158,N_111);
xnor U2140 (N_2140,N_821,N_1502);
nor U2141 (N_2141,N_626,N_303);
xor U2142 (N_2142,N_1442,N_651);
xnor U2143 (N_2143,N_1457,N_1687);
nor U2144 (N_2144,N_850,N_260);
xor U2145 (N_2145,N_286,N_1850);
nor U2146 (N_2146,N_745,N_54);
nor U2147 (N_2147,N_930,N_1078);
nand U2148 (N_2148,N_1936,N_526);
nor U2149 (N_2149,N_451,N_1916);
or U2150 (N_2150,N_193,N_1982);
and U2151 (N_2151,N_1184,N_704);
and U2152 (N_2152,N_6,N_378);
and U2153 (N_2153,N_300,N_766);
and U2154 (N_2154,N_1161,N_1440);
xnor U2155 (N_2155,N_1994,N_929);
and U2156 (N_2156,N_375,N_346);
nand U2157 (N_2157,N_1331,N_616);
or U2158 (N_2158,N_1598,N_1570);
xnor U2159 (N_2159,N_922,N_69);
nand U2160 (N_2160,N_342,N_1182);
or U2161 (N_2161,N_642,N_188);
nand U2162 (N_2162,N_1474,N_641);
or U2163 (N_2163,N_508,N_199);
xnor U2164 (N_2164,N_1880,N_11);
xnor U2165 (N_2165,N_0,N_1255);
and U2166 (N_2166,N_1056,N_1595);
and U2167 (N_2167,N_156,N_757);
and U2168 (N_2168,N_51,N_1902);
xor U2169 (N_2169,N_904,N_1);
or U2170 (N_2170,N_1790,N_743);
and U2171 (N_2171,N_1145,N_728);
nand U2172 (N_2172,N_1745,N_1793);
nand U2173 (N_2173,N_1728,N_637);
nor U2174 (N_2174,N_559,N_1877);
nand U2175 (N_2175,N_650,N_1082);
and U2176 (N_2176,N_89,N_946);
and U2177 (N_2177,N_1139,N_1908);
nor U2178 (N_2178,N_803,N_1911);
and U2179 (N_2179,N_1213,N_461);
and U2180 (N_2180,N_1480,N_1131);
nor U2181 (N_2181,N_352,N_167);
nand U2182 (N_2182,N_1462,N_1108);
and U2183 (N_2183,N_1453,N_1342);
or U2184 (N_2184,N_471,N_225);
or U2185 (N_2185,N_1668,N_1299);
or U2186 (N_2186,N_747,N_1863);
xor U2187 (N_2187,N_973,N_1297);
xor U2188 (N_2188,N_1849,N_1534);
or U2189 (N_2189,N_1556,N_306);
or U2190 (N_2190,N_1298,N_399);
xnor U2191 (N_2191,N_419,N_848);
or U2192 (N_2192,N_458,N_1160);
xor U2193 (N_2193,N_1707,N_1852);
nor U2194 (N_2194,N_47,N_1637);
xor U2195 (N_2195,N_1886,N_481);
nor U2196 (N_2196,N_125,N_1756);
nand U2197 (N_2197,N_976,N_794);
or U2198 (N_2198,N_1964,N_1676);
or U2199 (N_2199,N_112,N_487);
xnor U2200 (N_2200,N_1530,N_1679);
or U2201 (N_2201,N_1577,N_121);
xor U2202 (N_2202,N_416,N_1452);
nor U2203 (N_2203,N_681,N_865);
xnor U2204 (N_2204,N_1953,N_1077);
nand U2205 (N_2205,N_1235,N_994);
and U2206 (N_2206,N_1520,N_1828);
or U2207 (N_2207,N_76,N_1446);
or U2208 (N_2208,N_750,N_1431);
and U2209 (N_2209,N_1592,N_868);
and U2210 (N_2210,N_1152,N_1682);
xnor U2211 (N_2211,N_390,N_1239);
or U2212 (N_2212,N_1028,N_1589);
nand U2213 (N_2213,N_1353,N_412);
and U2214 (N_2214,N_1105,N_1253);
nand U2215 (N_2215,N_1210,N_1121);
and U2216 (N_2216,N_319,N_1262);
or U2217 (N_2217,N_1533,N_366);
and U2218 (N_2218,N_632,N_758);
nor U2219 (N_2219,N_573,N_46);
xor U2220 (N_2220,N_1169,N_1747);
nand U2221 (N_2221,N_634,N_1630);
or U2222 (N_2222,N_1600,N_1320);
xnor U2223 (N_2223,N_1903,N_1721);
xor U2224 (N_2224,N_1883,N_879);
xnor U2225 (N_2225,N_993,N_1318);
and U2226 (N_2226,N_1532,N_423);
xor U2227 (N_2227,N_1896,N_1041);
xor U2228 (N_2228,N_1319,N_588);
nor U2229 (N_2229,N_1675,N_708);
nor U2230 (N_2230,N_1275,N_863);
and U2231 (N_2231,N_888,N_392);
nand U2232 (N_2232,N_1439,N_428);
xnor U2233 (N_2233,N_1632,N_469);
xor U2234 (N_2234,N_1371,N_847);
xnor U2235 (N_2235,N_327,N_834);
or U2236 (N_2236,N_194,N_1710);
and U2237 (N_2237,N_158,N_295);
nand U2238 (N_2238,N_334,N_1386);
nor U2239 (N_2239,N_729,N_1434);
and U2240 (N_2240,N_437,N_902);
or U2241 (N_2241,N_1504,N_1163);
xnor U2242 (N_2242,N_1196,N_725);
nor U2243 (N_2243,N_1801,N_1102);
nor U2244 (N_2244,N_1807,N_1702);
nor U2245 (N_2245,N_990,N_1538);
nor U2246 (N_2246,N_949,N_1958);
or U2247 (N_2247,N_1218,N_1547);
xnor U2248 (N_2248,N_201,N_1065);
nor U2249 (N_2249,N_1083,N_1476);
or U2250 (N_2250,N_213,N_590);
and U2251 (N_2251,N_12,N_74);
or U2252 (N_2252,N_734,N_1537);
nand U2253 (N_2253,N_1199,N_1594);
nor U2254 (N_2254,N_1578,N_272);
nor U2255 (N_2255,N_1389,N_115);
and U2256 (N_2256,N_26,N_321);
xnor U2257 (N_2257,N_719,N_436);
nand U2258 (N_2258,N_1243,N_1040);
nand U2259 (N_2259,N_1961,N_1941);
and U2260 (N_2260,N_95,N_1999);
nand U2261 (N_2261,N_1719,N_493);
and U2262 (N_2262,N_249,N_1097);
and U2263 (N_2263,N_1751,N_707);
or U2264 (N_2264,N_867,N_1268);
or U2265 (N_2265,N_502,N_120);
and U2266 (N_2266,N_14,N_1094);
and U2267 (N_2267,N_629,N_997);
xor U2268 (N_2268,N_1970,N_656);
nand U2269 (N_2269,N_1378,N_897);
or U2270 (N_2270,N_383,N_1060);
and U2271 (N_2271,N_1260,N_355);
nor U2272 (N_2272,N_1610,N_1330);
xnor U2273 (N_2273,N_699,N_557);
and U2274 (N_2274,N_1146,N_1920);
and U2275 (N_2275,N_860,N_1463);
xnor U2276 (N_2276,N_1586,N_1655);
nor U2277 (N_2277,N_1869,N_1251);
xnor U2278 (N_2278,N_1705,N_1979);
and U2279 (N_2279,N_1678,N_647);
and U2280 (N_2280,N_1208,N_368);
and U2281 (N_2281,N_359,N_1284);
nand U2282 (N_2282,N_107,N_800);
and U2283 (N_2283,N_256,N_1390);
or U2284 (N_2284,N_1729,N_1061);
nand U2285 (N_2285,N_400,N_797);
and U2286 (N_2286,N_1400,N_1288);
or U2287 (N_2287,N_75,N_126);
and U2288 (N_2288,N_205,N_1456);
xor U2289 (N_2289,N_1653,N_435);
xor U2290 (N_2290,N_1274,N_1664);
nor U2291 (N_2291,N_305,N_763);
xnor U2292 (N_2292,N_1261,N_41);
or U2293 (N_2293,N_1215,N_104);
nor U2294 (N_2294,N_1680,N_4);
nand U2295 (N_2295,N_1940,N_684);
nor U2296 (N_2296,N_1421,N_1549);
or U2297 (N_2297,N_1794,N_690);
nor U2298 (N_2298,N_1214,N_1623);
nor U2299 (N_2299,N_1130,N_698);
nand U2300 (N_2300,N_103,N_1002);
xnor U2301 (N_2301,N_1693,N_913);
or U2302 (N_2302,N_873,N_200);
or U2303 (N_2303,N_1767,N_1690);
and U2304 (N_2304,N_620,N_685);
nand U2305 (N_2305,N_459,N_141);
nor U2306 (N_2306,N_280,N_281);
or U2307 (N_2307,N_1848,N_106);
and U2308 (N_2308,N_1301,N_1220);
nor U2309 (N_2309,N_1173,N_1415);
xnor U2310 (N_2310,N_1272,N_1868);
or U2311 (N_2311,N_784,N_872);
nor U2312 (N_2312,N_1355,N_903);
nand U2313 (N_2313,N_1007,N_1295);
xor U2314 (N_2314,N_1226,N_1976);
xor U2315 (N_2315,N_1487,N_248);
xnor U2316 (N_2316,N_1124,N_484);
and U2317 (N_2317,N_1277,N_227);
nor U2318 (N_2318,N_939,N_1071);
or U2319 (N_2319,N_228,N_1114);
or U2320 (N_2320,N_517,N_139);
and U2321 (N_2321,N_601,N_1709);
nor U2322 (N_2322,N_1633,N_1168);
nor U2323 (N_2323,N_657,N_391);
or U2324 (N_2324,N_1489,N_988);
nor U2325 (N_2325,N_1795,N_1783);
nand U2326 (N_2326,N_906,N_836);
or U2327 (N_2327,N_1921,N_1064);
or U2328 (N_2328,N_769,N_195);
xor U2329 (N_2329,N_212,N_1815);
or U2330 (N_2330,N_1560,N_1329);
xnor U2331 (N_2331,N_153,N_1458);
nand U2332 (N_2332,N_1864,N_1376);
or U2333 (N_2333,N_15,N_709);
nor U2334 (N_2334,N_1413,N_1244);
xor U2335 (N_2335,N_1397,N_1306);
and U2336 (N_2336,N_217,N_131);
or U2337 (N_2337,N_25,N_497);
xnor U2338 (N_2338,N_438,N_688);
nor U2339 (N_2339,N_1505,N_901);
and U2340 (N_2340,N_748,N_1069);
xnor U2341 (N_2341,N_1713,N_1831);
and U2342 (N_2342,N_945,N_1531);
and U2343 (N_2343,N_756,N_418);
nor U2344 (N_2344,N_1760,N_135);
xnor U2345 (N_2345,N_958,N_525);
xnor U2346 (N_2346,N_268,N_254);
nand U2347 (N_2347,N_639,N_1066);
and U2348 (N_2348,N_474,N_168);
xor U2349 (N_2349,N_1621,N_806);
nand U2350 (N_2350,N_814,N_1989);
or U2351 (N_2351,N_155,N_1695);
and U2352 (N_2352,N_1889,N_1231);
nand U2353 (N_2353,N_1614,N_1969);
nor U2354 (N_2354,N_1482,N_339);
and U2355 (N_2355,N_1735,N_72);
nor U2356 (N_2356,N_1539,N_916);
or U2357 (N_2357,N_802,N_1216);
and U2358 (N_2358,N_1932,N_1259);
xnor U2359 (N_2359,N_445,N_1829);
nor U2360 (N_2360,N_356,N_607);
xnor U2361 (N_2361,N_292,N_1411);
nor U2362 (N_2362,N_1792,N_432);
nand U2363 (N_2363,N_1038,N_1154);
xnor U2364 (N_2364,N_241,N_1939);
and U2365 (N_2365,N_380,N_298);
xnor U2366 (N_2366,N_1616,N_1321);
and U2367 (N_2367,N_1062,N_1493);
nand U2368 (N_2368,N_127,N_1054);
nor U2369 (N_2369,N_1375,N_154);
nor U2370 (N_2370,N_1599,N_1129);
nor U2371 (N_2371,N_116,N_145);
or U2372 (N_2372,N_1096,N_1111);
nand U2373 (N_2373,N_439,N_488);
or U2374 (N_2374,N_1287,N_876);
or U2375 (N_2375,N_1263,N_1138);
or U2376 (N_2376,N_825,N_1978);
and U2377 (N_2377,N_1835,N_1784);
xnor U2378 (N_2378,N_420,N_1652);
xor U2379 (N_2379,N_705,N_933);
nor U2380 (N_2380,N_182,N_539);
nand U2381 (N_2381,N_950,N_100);
nor U2382 (N_2382,N_1689,N_1232);
or U2383 (N_2383,N_467,N_840);
and U2384 (N_2384,N_1862,N_563);
nor U2385 (N_2385,N_1478,N_932);
or U2386 (N_2386,N_1361,N_759);
nor U2387 (N_2387,N_1245,N_123);
and U2388 (N_2388,N_1820,N_871);
xor U2389 (N_2389,N_1382,N_202);
nor U2390 (N_2390,N_1723,N_885);
nor U2391 (N_2391,N_1464,N_1646);
nand U2392 (N_2392,N_952,N_1211);
or U2393 (N_2393,N_1572,N_1209);
nand U2394 (N_2394,N_569,N_1089);
or U2395 (N_2395,N_489,N_597);
nand U2396 (N_2396,N_1604,N_925);
nor U2397 (N_2397,N_336,N_414);
or U2398 (N_2398,N_1307,N_118);
nor U2399 (N_2399,N_584,N_1699);
or U2400 (N_2400,N_1224,N_1327);
or U2401 (N_2401,N_1433,N_1596);
or U2402 (N_2402,N_1469,N_1303);
or U2403 (N_2403,N_870,N_571);
nand U2404 (N_2404,N_1696,N_1727);
xor U2405 (N_2405,N_161,N_1956);
nand U2406 (N_2406,N_1593,N_240);
nor U2407 (N_2407,N_931,N_316);
nor U2408 (N_2408,N_788,N_900);
or U2409 (N_2409,N_1219,N_877);
xnor U2410 (N_2410,N_567,N_1882);
nand U2411 (N_2411,N_1407,N_755);
or U2412 (N_2412,N_1308,N_754);
nand U2413 (N_2413,N_223,N_627);
nand U2414 (N_2414,N_1363,N_826);
or U2415 (N_2415,N_1965,N_388);
nor U2416 (N_2416,N_1079,N_1519);
xor U2417 (N_2417,N_880,N_621);
xnor U2418 (N_2418,N_1647,N_226);
nand U2419 (N_2419,N_1048,N_1913);
xnor U2420 (N_2420,N_110,N_1426);
nor U2421 (N_2421,N_1264,N_108);
and U2422 (N_2422,N_1887,N_1204);
xnor U2423 (N_2423,N_1934,N_210);
or U2424 (N_2424,N_968,N_1856);
nor U2425 (N_2425,N_152,N_500);
and U2426 (N_2426,N_1070,N_1229);
nor U2427 (N_2427,N_133,N_136);
xnor U2428 (N_2428,N_454,N_1893);
xor U2429 (N_2429,N_1972,N_1959);
xnor U2430 (N_2430,N_1110,N_434);
xor U2431 (N_2431,N_790,N_1346);
nor U2432 (N_2432,N_1119,N_1559);
and U2433 (N_2433,N_1890,N_73);
nor U2434 (N_2434,N_1666,N_1372);
nand U2435 (N_2435,N_1726,N_496);
or U2436 (N_2436,N_1834,N_787);
and U2437 (N_2437,N_1924,N_1484);
xor U2438 (N_2438,N_117,N_942);
or U2439 (N_2439,N_878,N_232);
or U2440 (N_2440,N_960,N_648);
xor U2441 (N_2441,N_1651,N_1561);
or U2442 (N_2442,N_1870,N_1836);
xnor U2443 (N_2443,N_1075,N_13);
xnor U2444 (N_2444,N_1658,N_465);
xor U2445 (N_2445,N_1465,N_1481);
nand U2446 (N_2446,N_1496,N_777);
xor U2447 (N_2447,N_266,N_449);
nand U2448 (N_2448,N_1861,N_238);
nand U2449 (N_2449,N_710,N_190);
xnor U2450 (N_2450,N_1155,N_371);
and U2451 (N_2451,N_45,N_838);
or U2452 (N_2452,N_446,N_197);
nor U2453 (N_2453,N_1142,N_329);
xnor U2454 (N_2454,N_475,N_832);
or U2455 (N_2455,N_1846,N_425);
nor U2456 (N_2456,N_177,N_1186);
nor U2457 (N_2457,N_789,N_1187);
or U2458 (N_2458,N_33,N_1104);
or U2459 (N_2459,N_653,N_1640);
nand U2460 (N_2460,N_1053,N_527);
or U2461 (N_2461,N_1276,N_1418);
and U2462 (N_2462,N_203,N_1766);
nor U2463 (N_2463,N_1283,N_1725);
xnor U2464 (N_2464,N_1919,N_230);
nand U2465 (N_2465,N_250,N_1581);
nand U2466 (N_2466,N_1591,N_893);
or U2467 (N_2467,N_841,N_1351);
and U2468 (N_2468,N_1125,N_550);
or U2469 (N_2469,N_1479,N_987);
or U2470 (N_2470,N_669,N_1952);
and U2471 (N_2471,N_53,N_765);
and U2472 (N_2472,N_996,N_752);
nor U2473 (N_2473,N_1238,N_796);
nand U2474 (N_2474,N_58,N_1230);
xnor U2475 (N_2475,N_537,N_1697);
xor U2476 (N_2476,N_1500,N_38);
nand U2477 (N_2477,N_1009,N_348);
or U2478 (N_2478,N_1918,N_1279);
xor U2479 (N_2479,N_151,N_1730);
and U2480 (N_2480,N_570,N_1222);
xor U2481 (N_2481,N_1761,N_558);
nand U2482 (N_2482,N_1005,N_856);
or U2483 (N_2483,N_507,N_1894);
and U2484 (N_2484,N_164,N_1752);
nor U2485 (N_2485,N_864,N_1998);
and U2486 (N_2486,N_288,N_1170);
nand U2487 (N_2487,N_1349,N_379);
nor U2488 (N_2488,N_70,N_1879);
nand U2489 (N_2489,N_472,N_1832);
nor U2490 (N_2490,N_686,N_1354);
and U2491 (N_2491,N_181,N_1278);
nand U2492 (N_2492,N_1018,N_934);
or U2493 (N_2493,N_322,N_1194);
and U2494 (N_2494,N_1432,N_1542);
nand U2495 (N_2495,N_980,N_178);
and U2496 (N_2496,N_1627,N_1845);
xor U2497 (N_2497,N_124,N_1967);
xor U2498 (N_2498,N_1471,N_1923);
nand U2499 (N_2499,N_923,N_1466);
or U2500 (N_2500,N_1419,N_1607);
and U2501 (N_2501,N_723,N_1337);
nand U2502 (N_2502,N_1514,N_1391);
or U2503 (N_2503,N_130,N_1492);
or U2504 (N_2504,N_1585,N_309);
nor U2505 (N_2505,N_964,N_1765);
nand U2506 (N_2506,N_1328,N_780);
and U2507 (N_2507,N_706,N_381);
and U2508 (N_2508,N_514,N_1044);
and U2509 (N_2509,N_353,N_1802);
nand U2510 (N_2510,N_1569,N_1459);
nor U2511 (N_2511,N_594,N_97);
or U2512 (N_2512,N_1039,N_1499);
and U2513 (N_2513,N_62,N_1149);
and U2514 (N_2514,N_296,N_1625);
nor U2515 (N_2515,N_1648,N_290);
and U2516 (N_2516,N_519,N_1700);
nor U2517 (N_2517,N_674,N_955);
and U2518 (N_2518,N_1764,N_521);
xnor U2519 (N_2519,N_251,N_478);
and U2520 (N_2520,N_1343,N_1414);
and U2521 (N_2521,N_140,N_753);
xor U2522 (N_2522,N_1991,N_1543);
xor U2523 (N_2523,N_480,N_505);
nor U2524 (N_2524,N_943,N_716);
nor U2525 (N_2525,N_1387,N_1769);
and U2526 (N_2526,N_43,N_1344);
xnor U2527 (N_2527,N_1313,N_701);
nor U2528 (N_2528,N_1654,N_1624);
nand U2529 (N_2529,N_522,N_820);
nand U2530 (N_2530,N_767,N_608);
nand U2531 (N_2531,N_941,N_1202);
and U2532 (N_2532,N_1134,N_1992);
nor U2533 (N_2533,N_1635,N_1368);
nor U2534 (N_2534,N_1388,N_1778);
nor U2535 (N_2535,N_30,N_1055);
or U2536 (N_2536,N_1150,N_1293);
nand U2537 (N_2537,N_668,N_396);
and U2538 (N_2538,N_1384,N_1922);
xor U2539 (N_2539,N_1657,N_265);
nand U2540 (N_2540,N_2,N_580);
xor U2541 (N_2541,N_1010,N_1030);
nor U2542 (N_2542,N_463,N_1825);
nand U2543 (N_2543,N_914,N_591);
nand U2544 (N_2544,N_1423,N_429);
and U2545 (N_2545,N_16,N_1527);
nor U2546 (N_2546,N_160,N_1123);
or U2547 (N_2547,N_35,N_715);
nor U2548 (N_2548,N_90,N_636);
nand U2549 (N_2549,N_1067,N_1704);
xnor U2550 (N_2550,N_1582,N_393);
and U2551 (N_2551,N_1485,N_237);
nand U2552 (N_2552,N_1960,N_48);
nor U2553 (N_2553,N_560,N_1162);
nor U2554 (N_2554,N_1203,N_852);
and U2555 (N_2555,N_312,N_333);
or U2556 (N_2556,N_311,N_299);
and U2557 (N_2557,N_63,N_1247);
and U2558 (N_2558,N_1806,N_1910);
nor U2559 (N_2559,N_717,N_1257);
and U2560 (N_2560,N_1133,N_1223);
and U2561 (N_2561,N_324,N_1364);
nor U2562 (N_2562,N_376,N_1050);
xor U2563 (N_2563,N_1685,N_917);
nor U2564 (N_2564,N_132,N_1291);
and U2565 (N_2565,N_361,N_1947);
or U2566 (N_2566,N_1477,N_1686);
nand U2567 (N_2567,N_1317,N_1734);
or U2568 (N_2568,N_1109,N_1659);
and U2569 (N_2569,N_614,N_259);
nand U2570 (N_2570,N_1091,N_1178);
nand U2571 (N_2571,N_1193,N_677);
or U2572 (N_2572,N_566,N_1003);
xnor U2573 (N_2573,N_278,N_102);
nor U2574 (N_2574,N_1460,N_1473);
or U2575 (N_2575,N_974,N_732);
nand U2576 (N_2576,N_91,N_1662);
xor U2577 (N_2577,N_735,N_866);
xor U2578 (N_2578,N_1993,N_61);
xor U2579 (N_2579,N_918,N_532);
nand U2580 (N_2580,N_673,N_829);
xnor U2581 (N_2581,N_905,N_1296);
and U2582 (N_2582,N_1757,N_1240);
xor U2583 (N_2583,N_364,N_1417);
or U2584 (N_2584,N_257,N_1788);
nor U2585 (N_2585,N_1524,N_1174);
nor U2586 (N_2586,N_1951,N_270);
or U2587 (N_2587,N_464,N_1776);
xnor U2588 (N_2588,N_1669,N_192);
and U2589 (N_2589,N_830,N_1573);
nand U2590 (N_2590,N_849,N_98);
or U2591 (N_2591,N_545,N_1670);
xnor U2592 (N_2592,N_778,N_1454);
and U2593 (N_2593,N_561,N_1302);
xnor U2594 (N_2594,N_644,N_1181);
nand U2595 (N_2595,N_1076,N_413);
and U2596 (N_2596,N_1782,N_1603);
nand U2597 (N_2597,N_808,N_1495);
and U2598 (N_2598,N_1290,N_1098);
nor U2599 (N_2599,N_165,N_1198);
nand U2600 (N_2600,N_1885,N_1093);
or U2601 (N_2601,N_1691,N_703);
xor U2602 (N_2602,N_1036,N_1837);
nor U2603 (N_2603,N_801,N_592);
nor U2604 (N_2604,N_1798,N_541);
nand U2605 (N_2605,N_1324,N_186);
xor U2606 (N_2606,N_1450,N_262);
nand U2607 (N_2607,N_805,N_1021);
xnor U2608 (N_2608,N_476,N_80);
nand U2609 (N_2609,N_1855,N_1771);
nand U2610 (N_2610,N_1732,N_99);
or U2611 (N_2611,N_1004,N_1126);
nand U2612 (N_2612,N_1643,N_424);
nor U2613 (N_2613,N_585,N_662);
nor U2614 (N_2614,N_1785,N_492);
and U2615 (N_2615,N_857,N_1019);
nand U2616 (N_2616,N_162,N_553);
and U2617 (N_2617,N_1571,N_733);
or U2618 (N_2618,N_297,N_1606);
xor U2619 (N_2619,N_462,N_1912);
nor U2620 (N_2620,N_1141,N_724);
nor U2621 (N_2621,N_516,N_810);
or U2622 (N_2622,N_1190,N_1437);
xor U2623 (N_2623,N_599,N_546);
nand U2624 (N_2624,N_938,N_544);
or U2625 (N_2625,N_1938,N_1946);
nor U2626 (N_2626,N_937,N_554);
xor U2627 (N_2627,N_340,N_1995);
or U2628 (N_2628,N_1584,N_1167);
nand U2629 (N_2629,N_78,N_972);
and U2630 (N_2630,N_1217,N_1808);
xnor U2631 (N_2631,N_1755,N_166);
nand U2632 (N_2632,N_1740,N_1348);
nand U2633 (N_2633,N_989,N_741);
and U2634 (N_2634,N_959,N_1017);
xor U2635 (N_2635,N_137,N_1326);
nand U2636 (N_2636,N_809,N_1866);
nor U2637 (N_2637,N_609,N_530);
and U2638 (N_2638,N_1871,N_638);
nor U2639 (N_2639,N_920,N_317);
nand U2640 (N_2640,N_1246,N_760);
nor U2641 (N_2641,N_402,N_676);
nor U2642 (N_2642,N_1047,N_1366);
or U2643 (N_2643,N_842,N_1945);
xor U2644 (N_2644,N_1136,N_1472);
xor U2645 (N_2645,N_1304,N_411);
and U2646 (N_2646,N_174,N_105);
nor U2647 (N_2647,N_283,N_578);
and U2648 (N_2648,N_1273,N_1394);
and U2649 (N_2649,N_341,N_18);
or U2650 (N_2650,N_764,N_417);
or U2651 (N_2651,N_172,N_325);
xor U2652 (N_2652,N_373,N_96);
and U2653 (N_2653,N_377,N_431);
nand U2654 (N_2654,N_643,N_406);
nand U2655 (N_2655,N_244,N_1408);
and U2656 (N_2656,N_722,N_548);
nor U2657 (N_2657,N_1430,N_1032);
and U2658 (N_2658,N_1380,N_343);
nor U2659 (N_2659,N_447,N_1441);
nand U2660 (N_2660,N_1515,N_1754);
and U2661 (N_2661,N_470,N_1758);
nand U2662 (N_2662,N_369,N_335);
or U2663 (N_2663,N_87,N_1762);
xor U2664 (N_2664,N_1528,N_207);
nor U2665 (N_2665,N_79,N_277);
nand U2666 (N_2666,N_680,N_635);
xor U2667 (N_2667,N_501,N_1576);
nor U2668 (N_2668,N_1772,N_596);
xor U2669 (N_2669,N_1072,N_382);
and U2670 (N_2670,N_1844,N_1164);
or U2671 (N_2671,N_1781,N_183);
nor U2672 (N_2672,N_81,N_1681);
nor U2673 (N_2673,N_966,N_911);
nor U2674 (N_2674,N_291,N_1557);
or U2675 (N_2675,N_995,N_556);
nor U2676 (N_2676,N_649,N_42);
nor U2677 (N_2677,N_187,N_1443);
or U2678 (N_2678,N_511,N_1615);
or U2679 (N_2679,N_59,N_1103);
and U2680 (N_2680,N_1860,N_267);
or U2681 (N_2681,N_218,N_1063);
xnor U2682 (N_2682,N_1171,N_1242);
xnor U2683 (N_2683,N_927,N_940);
xor U2684 (N_2684,N_807,N_881);
nor U2685 (N_2685,N_1080,N_39);
nor U2686 (N_2686,N_862,N_1878);
and U2687 (N_2687,N_88,N_1248);
nand U2688 (N_2688,N_1180,N_1033);
and U2689 (N_2689,N_1526,N_786);
nor U2690 (N_2690,N_57,N_1447);
and U2691 (N_2691,N_261,N_398);
xor U2692 (N_2692,N_1949,N_540);
nand U2693 (N_2693,N_683,N_31);
nor U2694 (N_2694,N_884,N_185);
and U2695 (N_2695,N_1137,N_1300);
nand U2696 (N_2696,N_721,N_854);
or U2697 (N_2697,N_1525,N_1314);
or U2698 (N_2698,N_263,N_17);
nand U2699 (N_2699,N_19,N_909);
nor U2700 (N_2700,N_1840,N_1081);
nor U2701 (N_2701,N_844,N_583);
and U2702 (N_2702,N_985,N_1715);
nand U2703 (N_2703,N_1045,N_1810);
and U2704 (N_2704,N_739,N_229);
xor U2705 (N_2705,N_289,N_523);
and U2706 (N_2706,N_1212,N_534);
and U2707 (N_2707,N_1120,N_961);
nor U2708 (N_2708,N_1085,N_269);
xor U2709 (N_2709,N_1823,N_979);
nor U2710 (N_2710,N_1580,N_1416);
xor U2711 (N_2711,N_1738,N_1392);
or U2712 (N_2712,N_851,N_509);
nor U2713 (N_2713,N_751,N_1660);
and U2714 (N_2714,N_603,N_211);
xor U2715 (N_2715,N_318,N_895);
or U2716 (N_2716,N_1983,N_1197);
and U2717 (N_2717,N_405,N_387);
and U2718 (N_2718,N_779,N_1468);
and U2719 (N_2719,N_1435,N_101);
and U2720 (N_2720,N_1427,N_1395);
xnor U2721 (N_2721,N_928,N_1843);
nor U2722 (N_2722,N_1770,N_518);
nand U2723 (N_2723,N_1587,N_233);
nand U2724 (N_2724,N_1340,N_255);
nor U2725 (N_2725,N_1613,N_682);
and U2726 (N_2726,N_1620,N_1309);
and U2727 (N_2727,N_494,N_455);
or U2728 (N_2728,N_490,N_1683);
nand U2729 (N_2729,N_1558,N_421);
nand U2730 (N_2730,N_386,N_1176);
nor U2731 (N_2731,N_1352,N_1488);
or U2732 (N_2732,N_785,N_1564);
nand U2733 (N_2733,N_1649,N_776);
nand U2734 (N_2734,N_351,N_1249);
or U2735 (N_2735,N_795,N_658);
nor U2736 (N_2736,N_354,N_1335);
or U2737 (N_2737,N_1611,N_793);
nand U2738 (N_2738,N_1144,N_169);
xnor U2739 (N_2739,N_1694,N_323);
xnor U2740 (N_2740,N_1803,N_1521);
nand U2741 (N_2741,N_762,N_572);
and U2742 (N_2742,N_1270,N_1786);
or U2743 (N_2743,N_924,N_279);
nor U2744 (N_2744,N_293,N_773);
and U2745 (N_2745,N_1043,N_1568);
nor U2746 (N_2746,N_600,N_1827);
xor U2747 (N_2747,N_44,N_1841);
xnor U2748 (N_2748,N_663,N_953);
xnor U2749 (N_2749,N_52,N_1360);
nor U2750 (N_2750,N_912,N_1269);
and U2751 (N_2751,N_1401,N_1645);
nand U2752 (N_2752,N_628,N_828);
xnor U2753 (N_2753,N_66,N_37);
nor U2754 (N_2754,N_302,N_430);
or U2755 (N_2755,N_812,N_214);
nor U2756 (N_2756,N_727,N_1567);
and U2757 (N_2757,N_1562,N_170);
nor U2758 (N_2758,N_1237,N_271);
nand U2759 (N_2759,N_134,N_712);
nand U2760 (N_2760,N_1737,N_1601);
or U2761 (N_2761,N_184,N_1266);
and U2762 (N_2762,N_543,N_528);
nor U2763 (N_2763,N_1529,N_815);
nand U2764 (N_2764,N_971,N_179);
xor U2765 (N_2765,N_1436,N_1948);
or U2766 (N_2766,N_1099,N_700);
xor U2767 (N_2767,N_1897,N_1830);
nand U2768 (N_2768,N_919,N_1663);
nand U2769 (N_2769,N_1265,N_224);
and U2770 (N_2770,N_1073,N_1398);
xor U2771 (N_2771,N_1312,N_1777);
xor U2772 (N_2772,N_347,N_1501);
and U2773 (N_2773,N_287,N_1535);
xnor U2774 (N_2774,N_586,N_630);
or U2775 (N_2775,N_1990,N_443);
or U2776 (N_2776,N_357,N_1867);
or U2777 (N_2777,N_595,N_1814);
or U2778 (N_2778,N_1254,N_220);
nand U2779 (N_2779,N_176,N_666);
or U2780 (N_2780,N_792,N_1201);
or U2781 (N_2781,N_1605,N_466);
and U2782 (N_2782,N_1997,N_1619);
nor U2783 (N_2783,N_1497,N_1553);
or U2784 (N_2784,N_1872,N_1175);
nor U2785 (N_2785,N_671,N_1405);
nand U2786 (N_2786,N_998,N_1634);
nor U2787 (N_2787,N_1172,N_1544);
nand U2788 (N_2788,N_1796,N_713);
xnor U2789 (N_2789,N_310,N_696);
nand U2790 (N_2790,N_551,N_1954);
nor U2791 (N_2791,N_1522,N_1804);
nand U2792 (N_2792,N_1325,N_1671);
or U2793 (N_2793,N_85,N_970);
nand U2794 (N_2794,N_896,N_1858);
xnor U2795 (N_2795,N_1971,N_1011);
nor U2796 (N_2796,N_798,N_611);
or U2797 (N_2797,N_1706,N_1717);
xnor U2798 (N_2798,N_926,N_1826);
and U2799 (N_2799,N_1151,N_1763);
nand U2800 (N_2800,N_1147,N_581);
nor U2801 (N_2801,N_1931,N_245);
xor U2802 (N_2802,N_1818,N_1362);
or U2803 (N_2803,N_679,N_655);
and U2804 (N_2804,N_426,N_819);
nor U2805 (N_2805,N_1986,N_575);
xor U2806 (N_2806,N_1703,N_1819);
nand U2807 (N_2807,N_326,N_1112);
and U2808 (N_2808,N_598,N_1744);
nor U2809 (N_2809,N_1192,N_1024);
nor U2810 (N_2810,N_1579,N_1449);
or U2811 (N_2811,N_574,N_1090);
nor U2812 (N_2812,N_529,N_1356);
nor U2813 (N_2813,N_1510,N_1574);
nor U2814 (N_2814,N_1552,N_394);
and U2815 (N_2815,N_1049,N_1842);
and U2816 (N_2816,N_1688,N_442);
xnor U2817 (N_2817,N_720,N_448);
nand U2818 (N_2818,N_986,N_499);
or U2819 (N_2819,N_1750,N_1789);
or U2820 (N_2820,N_818,N_1937);
and U2821 (N_2821,N_811,N_535);
nor U2822 (N_2822,N_1555,N_1115);
nor U2823 (N_2823,N_294,N_1980);
xnor U2824 (N_2824,N_1377,N_1984);
and U2825 (N_2825,N_1917,N_1357);
or U2826 (N_2826,N_410,N_1179);
nor U2827 (N_2827,N_672,N_1058);
and U2828 (N_2828,N_1117,N_1207);
and U2829 (N_2829,N_1602,N_150);
xnor U2830 (N_2830,N_1608,N_1746);
nand U2831 (N_2831,N_711,N_1677);
or U2832 (N_2832,N_1749,N_1642);
and U2833 (N_2833,N_899,N_235);
and U2834 (N_2834,N_1008,N_859);
xor U2835 (N_2835,N_1516,N_20);
nor U2836 (N_2836,N_1724,N_1509);
nand U2837 (N_2837,N_1258,N_468);
and U2838 (N_2838,N_1930,N_1451);
and U2839 (N_2839,N_1906,N_568);
nand U2840 (N_2840,N_1339,N_823);
nor U2841 (N_2841,N_1517,N_992);
or U2842 (N_2842,N_49,N_10);
nand U2843 (N_2843,N_1140,N_1636);
nor U2844 (N_2844,N_693,N_891);
nor U2845 (N_2845,N_1638,N_1311);
nand U2846 (N_2846,N_206,N_892);
nand U2847 (N_2847,N_1748,N_344);
nand U2848 (N_2848,N_1191,N_221);
nor U2849 (N_2849,N_1281,N_1393);
and U2850 (N_2850,N_1541,N_1565);
xor U2851 (N_2851,N_633,N_1014);
or U2852 (N_2852,N_965,N_1962);
xnor U2853 (N_2853,N_606,N_1195);
nand U2854 (N_2854,N_1101,N_869);
xor U2855 (N_2855,N_542,N_395);
or U2856 (N_2856,N_1183,N_1424);
and U2857 (N_2857,N_1051,N_146);
and U2858 (N_2858,N_746,N_384);
xor U2859 (N_2859,N_718,N_640);
or U2860 (N_2860,N_804,N_999);
or U2861 (N_2861,N_740,N_646);
nand U2862 (N_2862,N_775,N_397);
nand U2863 (N_2863,N_1403,N_360);
or U2864 (N_2864,N_1722,N_1250);
or U2865 (N_2865,N_1518,N_1892);
nand U2866 (N_2866,N_1743,N_1205);
xnor U2867 (N_2867,N_833,N_510);
nand U2868 (N_2868,N_403,N_665);
xnor U2869 (N_2869,N_524,N_1672);
nand U2870 (N_2870,N_824,N_1404);
nor U2871 (N_2871,N_1626,N_593);
or U2872 (N_2872,N_533,N_1396);
and U2873 (N_2873,N_831,N_138);
and U2874 (N_2874,N_1507,N_1412);
nor U2875 (N_2875,N_1853,N_1438);
nand U2876 (N_2876,N_1506,N_1292);
or U2877 (N_2877,N_1095,N_1927);
nand U2878 (N_2878,N_1503,N_1289);
xor U2879 (N_2879,N_180,N_1379);
nor U2880 (N_2880,N_1799,N_441);
and U2881 (N_2881,N_308,N_1188);
xor U2882 (N_2882,N_1399,N_749);
nor U2883 (N_2883,N_822,N_1132);
nor U2884 (N_2884,N_1385,N_768);
xor U2885 (N_2885,N_457,N_1323);
or U2886 (N_2886,N_1622,N_547);
xnor U2887 (N_2887,N_1338,N_1006);
xnor U2888 (N_2888,N_173,N_1716);
or U2889 (N_2889,N_1057,N_320);
nand U2890 (N_2890,N_1847,N_915);
and U2891 (N_2891,N_313,N_1548);
xnor U2892 (N_2892,N_512,N_782);
or U2893 (N_2893,N_1545,N_142);
nor U2894 (N_2894,N_345,N_1341);
xor U2895 (N_2895,N_1905,N_1016);
nor U2896 (N_2896,N_1935,N_485);
or U2897 (N_2897,N_936,N_50);
and U2898 (N_2898,N_1025,N_726);
nand U2899 (N_2899,N_1402,N_1316);
and U2900 (N_2900,N_1511,N_687);
nor U2901 (N_2901,N_363,N_610);
nand U2902 (N_2902,N_577,N_1166);
or U2903 (N_2903,N_1590,N_858);
nand U2904 (N_2904,N_1628,N_482);
nand U2905 (N_2905,N_1791,N_253);
and U2906 (N_2906,N_401,N_1127);
or U2907 (N_2907,N_1673,N_605);
xor U2908 (N_2908,N_1900,N_1031);
nand U2909 (N_2909,N_1692,N_1597);
or U2910 (N_2910,N_1800,N_21);
nor U2911 (N_2911,N_624,N_365);
or U2912 (N_2912,N_285,N_1020);
nor U2913 (N_2913,N_1001,N_582);
and U2914 (N_2914,N_1373,N_783);
and U2915 (N_2915,N_1429,N_314);
nand U2916 (N_2916,N_1720,N_1470);
xor U2917 (N_2917,N_408,N_1915);
and U2918 (N_2918,N_1305,N_264);
nand U2919 (N_2919,N_1374,N_1546);
xor U2920 (N_2920,N_1875,N_742);
or U2921 (N_2921,N_64,N_1086);
and U2922 (N_2922,N_827,N_907);
xnor U2923 (N_2923,N_538,N_175);
and U2924 (N_2924,N_1639,N_1812);
xor U2925 (N_2925,N_1661,N_921);
nand U2926 (N_2926,N_315,N_978);
nor U2927 (N_2927,N_774,N_520);
nand U2928 (N_2928,N_147,N_664);
and U2929 (N_2929,N_983,N_113);
nand U2930 (N_2930,N_1486,N_456);
or U2931 (N_2931,N_1822,N_362);
or U2932 (N_2932,N_1280,N_889);
nand U2933 (N_2933,N_697,N_1233);
or U2934 (N_2934,N_275,N_1551);
nor U2935 (N_2935,N_3,N_981);
and U2936 (N_2936,N_1350,N_258);
or U2937 (N_2937,N_944,N_951);
xnor U2938 (N_2938,N_1612,N_587);
xnor U2939 (N_2939,N_1895,N_963);
or U2940 (N_2940,N_1988,N_1467);
nor U2941 (N_2941,N_1609,N_1234);
or U2942 (N_2942,N_1550,N_8);
nor U2943 (N_2943,N_208,N_1422);
nand U2944 (N_2944,N_1409,N_198);
nor U2945 (N_2945,N_215,N_1631);
nand U2946 (N_2946,N_1490,N_1563);
xor U2947 (N_2947,N_894,N_531);
and U2948 (N_2948,N_407,N_954);
nor U2949 (N_2949,N_1966,N_982);
nand U2950 (N_2950,N_1733,N_1448);
xnor U2951 (N_2951,N_618,N_612);
and U2952 (N_2952,N_128,N_1629);
xor U2953 (N_2953,N_328,N_453);
or U2954 (N_2954,N_1898,N_143);
xnor U2955 (N_2955,N_84,N_1444);
nor U2956 (N_2956,N_304,N_513);
nand U2957 (N_2957,N_1816,N_157);
or U2958 (N_2958,N_898,N_109);
or U2959 (N_2959,N_837,N_1153);
and U2960 (N_2960,N_1483,N_1736);
nand U2961 (N_2961,N_22,N_1698);
and U2962 (N_2962,N_817,N_1029);
nor U2963 (N_2963,N_1282,N_622);
xor U2964 (N_2964,N_1068,N_55);
nand U2965 (N_2965,N_1909,N_28);
and U2966 (N_2966,N_1957,N_1759);
xor U2967 (N_2967,N_1975,N_1165);
nor U2968 (N_2968,N_504,N_1383);
and U2969 (N_2969,N_1926,N_1285);
xnor U2970 (N_2970,N_23,N_415);
xnor U2971 (N_2971,N_602,N_1358);
nand U2972 (N_2972,N_1334,N_536);
or U2973 (N_2973,N_483,N_350);
xnor U2974 (N_2974,N_962,N_332);
and U2975 (N_2975,N_60,N_549);
nor U2976 (N_2976,N_552,N_114);
nand U2977 (N_2977,N_1116,N_615);
or U2978 (N_2978,N_1741,N_1022);
xor U2979 (N_2979,N_910,N_935);
and U2980 (N_2980,N_65,N_731);
nand U2981 (N_2981,N_1933,N_1874);
or U2982 (N_2982,N_555,N_1236);
xor U2983 (N_2983,N_1787,N_67);
xnor U2984 (N_2984,N_1035,N_1332);
and U2985 (N_2985,N_1461,N_695);
nand U2986 (N_2986,N_1420,N_1714);
or U2987 (N_2987,N_738,N_204);
xnor U2988 (N_2988,N_1370,N_613);
and U2989 (N_2989,N_1996,N_477);
nand U2990 (N_2990,N_498,N_5);
nand U2991 (N_2991,N_967,N_358);
nor U2992 (N_2992,N_331,N_234);
xnor U2993 (N_2993,N_330,N_730);
and U2994 (N_2994,N_1881,N_1046);
nand U2995 (N_2995,N_385,N_1797);
and U2996 (N_2996,N_479,N_1315);
nor U2997 (N_2997,N_1942,N_1708);
and U2998 (N_2998,N_495,N_1310);
xnor U2999 (N_2999,N_1656,N_984);
xor U3000 (N_3000,N_432,N_987);
nand U3001 (N_3001,N_0,N_921);
xnor U3002 (N_3002,N_875,N_1303);
nand U3003 (N_3003,N_1064,N_60);
nand U3004 (N_3004,N_102,N_313);
and U3005 (N_3005,N_1358,N_161);
and U3006 (N_3006,N_1971,N_663);
and U3007 (N_3007,N_1846,N_100);
or U3008 (N_3008,N_1676,N_1714);
or U3009 (N_3009,N_1930,N_1712);
or U3010 (N_3010,N_290,N_1091);
nor U3011 (N_3011,N_504,N_1487);
nand U3012 (N_3012,N_1409,N_1394);
nor U3013 (N_3013,N_284,N_1912);
nor U3014 (N_3014,N_1430,N_255);
nor U3015 (N_3015,N_1801,N_1018);
nand U3016 (N_3016,N_1259,N_1563);
nand U3017 (N_3017,N_447,N_1594);
and U3018 (N_3018,N_1029,N_707);
nor U3019 (N_3019,N_48,N_1249);
or U3020 (N_3020,N_418,N_1049);
xnor U3021 (N_3021,N_1660,N_1886);
and U3022 (N_3022,N_1083,N_810);
nor U3023 (N_3023,N_1964,N_562);
or U3024 (N_3024,N_1283,N_209);
nand U3025 (N_3025,N_1919,N_1562);
nand U3026 (N_3026,N_1194,N_1583);
or U3027 (N_3027,N_812,N_52);
nor U3028 (N_3028,N_1257,N_251);
nor U3029 (N_3029,N_269,N_1478);
xor U3030 (N_3030,N_1143,N_927);
xnor U3031 (N_3031,N_1348,N_803);
and U3032 (N_3032,N_756,N_1161);
xnor U3033 (N_3033,N_1635,N_254);
nand U3034 (N_3034,N_725,N_1765);
nand U3035 (N_3035,N_733,N_1034);
nand U3036 (N_3036,N_1759,N_632);
and U3037 (N_3037,N_817,N_1931);
and U3038 (N_3038,N_1794,N_1620);
nand U3039 (N_3039,N_971,N_610);
and U3040 (N_3040,N_441,N_1741);
xnor U3041 (N_3041,N_1694,N_746);
xor U3042 (N_3042,N_1794,N_1868);
xor U3043 (N_3043,N_1266,N_455);
nor U3044 (N_3044,N_16,N_4);
nor U3045 (N_3045,N_339,N_1496);
nor U3046 (N_3046,N_1002,N_1632);
nand U3047 (N_3047,N_532,N_487);
or U3048 (N_3048,N_473,N_829);
or U3049 (N_3049,N_606,N_1499);
xor U3050 (N_3050,N_454,N_195);
nand U3051 (N_3051,N_1411,N_1139);
or U3052 (N_3052,N_1961,N_819);
xnor U3053 (N_3053,N_1579,N_478);
and U3054 (N_3054,N_300,N_707);
and U3055 (N_3055,N_1442,N_86);
or U3056 (N_3056,N_1802,N_1221);
nand U3057 (N_3057,N_118,N_805);
and U3058 (N_3058,N_1382,N_868);
or U3059 (N_3059,N_1855,N_163);
nand U3060 (N_3060,N_575,N_961);
nor U3061 (N_3061,N_1334,N_52);
and U3062 (N_3062,N_525,N_510);
xor U3063 (N_3063,N_1574,N_461);
or U3064 (N_3064,N_809,N_1330);
xnor U3065 (N_3065,N_1073,N_777);
nor U3066 (N_3066,N_594,N_1395);
or U3067 (N_3067,N_1312,N_1653);
nor U3068 (N_3068,N_495,N_1103);
or U3069 (N_3069,N_175,N_1104);
or U3070 (N_3070,N_1187,N_1065);
xnor U3071 (N_3071,N_1412,N_294);
or U3072 (N_3072,N_1883,N_1876);
nand U3073 (N_3073,N_278,N_1222);
or U3074 (N_3074,N_1457,N_67);
and U3075 (N_3075,N_1017,N_455);
or U3076 (N_3076,N_1161,N_636);
or U3077 (N_3077,N_186,N_1547);
nor U3078 (N_3078,N_273,N_369);
or U3079 (N_3079,N_364,N_1272);
xor U3080 (N_3080,N_1615,N_723);
xnor U3081 (N_3081,N_478,N_52);
xor U3082 (N_3082,N_703,N_1359);
xnor U3083 (N_3083,N_1809,N_333);
nand U3084 (N_3084,N_461,N_912);
nor U3085 (N_3085,N_631,N_1171);
or U3086 (N_3086,N_1209,N_247);
nor U3087 (N_3087,N_92,N_291);
or U3088 (N_3088,N_1981,N_963);
xor U3089 (N_3089,N_1348,N_1176);
xnor U3090 (N_3090,N_404,N_408);
or U3091 (N_3091,N_365,N_682);
nand U3092 (N_3092,N_564,N_149);
nor U3093 (N_3093,N_1993,N_1731);
and U3094 (N_3094,N_1143,N_28);
nand U3095 (N_3095,N_971,N_1822);
nand U3096 (N_3096,N_962,N_1408);
and U3097 (N_3097,N_1358,N_1708);
or U3098 (N_3098,N_361,N_603);
or U3099 (N_3099,N_1276,N_176);
and U3100 (N_3100,N_1989,N_1023);
or U3101 (N_3101,N_782,N_1469);
and U3102 (N_3102,N_399,N_1386);
or U3103 (N_3103,N_111,N_1677);
or U3104 (N_3104,N_1518,N_1848);
or U3105 (N_3105,N_1838,N_464);
or U3106 (N_3106,N_1203,N_739);
xnor U3107 (N_3107,N_1645,N_485);
nand U3108 (N_3108,N_1197,N_425);
or U3109 (N_3109,N_155,N_545);
nor U3110 (N_3110,N_1065,N_415);
or U3111 (N_3111,N_991,N_161);
and U3112 (N_3112,N_1540,N_856);
xnor U3113 (N_3113,N_721,N_136);
or U3114 (N_3114,N_10,N_1286);
nand U3115 (N_3115,N_1743,N_174);
xnor U3116 (N_3116,N_524,N_1959);
nor U3117 (N_3117,N_316,N_1289);
and U3118 (N_3118,N_370,N_421);
nor U3119 (N_3119,N_1267,N_64);
or U3120 (N_3120,N_136,N_322);
nor U3121 (N_3121,N_1407,N_1274);
nand U3122 (N_3122,N_291,N_773);
xnor U3123 (N_3123,N_1383,N_233);
xor U3124 (N_3124,N_1613,N_1494);
and U3125 (N_3125,N_1612,N_692);
nor U3126 (N_3126,N_1390,N_839);
nor U3127 (N_3127,N_1555,N_1621);
nand U3128 (N_3128,N_651,N_1633);
nor U3129 (N_3129,N_195,N_1628);
nor U3130 (N_3130,N_930,N_1404);
nor U3131 (N_3131,N_822,N_20);
nor U3132 (N_3132,N_249,N_1688);
xor U3133 (N_3133,N_490,N_567);
and U3134 (N_3134,N_213,N_1681);
and U3135 (N_3135,N_246,N_1602);
nand U3136 (N_3136,N_92,N_55);
xnor U3137 (N_3137,N_516,N_959);
or U3138 (N_3138,N_1091,N_1969);
xor U3139 (N_3139,N_1939,N_1358);
nand U3140 (N_3140,N_870,N_401);
xor U3141 (N_3141,N_1207,N_1591);
or U3142 (N_3142,N_1132,N_966);
and U3143 (N_3143,N_1807,N_1316);
xnor U3144 (N_3144,N_1793,N_1690);
or U3145 (N_3145,N_1924,N_1628);
or U3146 (N_3146,N_972,N_978);
nand U3147 (N_3147,N_649,N_881);
or U3148 (N_3148,N_1935,N_1842);
nand U3149 (N_3149,N_475,N_75);
xnor U3150 (N_3150,N_759,N_245);
xor U3151 (N_3151,N_824,N_495);
xor U3152 (N_3152,N_446,N_1274);
nor U3153 (N_3153,N_1429,N_1266);
nand U3154 (N_3154,N_729,N_1851);
nand U3155 (N_3155,N_512,N_751);
nand U3156 (N_3156,N_1684,N_538);
xor U3157 (N_3157,N_626,N_1458);
and U3158 (N_3158,N_907,N_607);
nor U3159 (N_3159,N_1030,N_70);
nand U3160 (N_3160,N_1161,N_702);
xnor U3161 (N_3161,N_781,N_1664);
nand U3162 (N_3162,N_1346,N_598);
nand U3163 (N_3163,N_722,N_1061);
xnor U3164 (N_3164,N_398,N_94);
or U3165 (N_3165,N_1209,N_765);
or U3166 (N_3166,N_1122,N_1199);
xnor U3167 (N_3167,N_1762,N_1663);
and U3168 (N_3168,N_1498,N_125);
xnor U3169 (N_3169,N_1084,N_1146);
xnor U3170 (N_3170,N_53,N_513);
nor U3171 (N_3171,N_1604,N_1622);
and U3172 (N_3172,N_1728,N_591);
and U3173 (N_3173,N_893,N_1122);
nand U3174 (N_3174,N_582,N_1503);
or U3175 (N_3175,N_1588,N_1544);
xnor U3176 (N_3176,N_1947,N_1556);
and U3177 (N_3177,N_1143,N_509);
or U3178 (N_3178,N_538,N_271);
and U3179 (N_3179,N_775,N_1034);
and U3180 (N_3180,N_205,N_1707);
or U3181 (N_3181,N_86,N_1337);
nand U3182 (N_3182,N_282,N_819);
or U3183 (N_3183,N_536,N_771);
nand U3184 (N_3184,N_1023,N_1721);
or U3185 (N_3185,N_1799,N_1335);
or U3186 (N_3186,N_980,N_710);
and U3187 (N_3187,N_1661,N_1328);
xor U3188 (N_3188,N_468,N_1042);
nor U3189 (N_3189,N_522,N_1020);
nor U3190 (N_3190,N_1923,N_54);
and U3191 (N_3191,N_557,N_75);
nand U3192 (N_3192,N_415,N_811);
nor U3193 (N_3193,N_833,N_726);
and U3194 (N_3194,N_79,N_863);
nand U3195 (N_3195,N_1742,N_476);
or U3196 (N_3196,N_1031,N_1181);
nor U3197 (N_3197,N_1013,N_869);
xor U3198 (N_3198,N_1387,N_1105);
xor U3199 (N_3199,N_1438,N_1984);
nor U3200 (N_3200,N_1842,N_1144);
and U3201 (N_3201,N_1877,N_78);
or U3202 (N_3202,N_334,N_419);
and U3203 (N_3203,N_840,N_766);
xor U3204 (N_3204,N_1373,N_8);
and U3205 (N_3205,N_1851,N_373);
and U3206 (N_3206,N_297,N_1841);
nor U3207 (N_3207,N_1000,N_1209);
nand U3208 (N_3208,N_730,N_481);
nand U3209 (N_3209,N_541,N_421);
nor U3210 (N_3210,N_1406,N_430);
or U3211 (N_3211,N_1221,N_850);
and U3212 (N_3212,N_487,N_286);
xnor U3213 (N_3213,N_1973,N_779);
nand U3214 (N_3214,N_508,N_1775);
or U3215 (N_3215,N_1016,N_1315);
nor U3216 (N_3216,N_1799,N_692);
xor U3217 (N_3217,N_966,N_1021);
nor U3218 (N_3218,N_1708,N_633);
or U3219 (N_3219,N_1763,N_279);
and U3220 (N_3220,N_1005,N_522);
and U3221 (N_3221,N_846,N_1053);
nor U3222 (N_3222,N_740,N_316);
xor U3223 (N_3223,N_1857,N_1991);
xor U3224 (N_3224,N_1130,N_173);
nand U3225 (N_3225,N_696,N_719);
and U3226 (N_3226,N_1407,N_1718);
xnor U3227 (N_3227,N_928,N_535);
xor U3228 (N_3228,N_1458,N_849);
nand U3229 (N_3229,N_1981,N_1915);
xor U3230 (N_3230,N_1704,N_1236);
nand U3231 (N_3231,N_1830,N_364);
xnor U3232 (N_3232,N_448,N_1050);
nor U3233 (N_3233,N_395,N_1586);
and U3234 (N_3234,N_1156,N_53);
nor U3235 (N_3235,N_571,N_1846);
or U3236 (N_3236,N_1155,N_578);
nor U3237 (N_3237,N_1754,N_1968);
and U3238 (N_3238,N_398,N_1947);
nor U3239 (N_3239,N_1656,N_926);
and U3240 (N_3240,N_1532,N_892);
nand U3241 (N_3241,N_949,N_1378);
nor U3242 (N_3242,N_619,N_479);
or U3243 (N_3243,N_445,N_753);
or U3244 (N_3244,N_1712,N_1916);
xor U3245 (N_3245,N_499,N_210);
nor U3246 (N_3246,N_1459,N_1053);
nor U3247 (N_3247,N_1706,N_1383);
xnor U3248 (N_3248,N_838,N_166);
or U3249 (N_3249,N_823,N_514);
and U3250 (N_3250,N_1542,N_837);
xor U3251 (N_3251,N_691,N_84);
nand U3252 (N_3252,N_1159,N_1405);
nor U3253 (N_3253,N_1563,N_188);
nor U3254 (N_3254,N_244,N_1896);
xor U3255 (N_3255,N_937,N_75);
nand U3256 (N_3256,N_435,N_205);
and U3257 (N_3257,N_980,N_1833);
and U3258 (N_3258,N_1392,N_1823);
nor U3259 (N_3259,N_1687,N_1011);
nor U3260 (N_3260,N_1267,N_1464);
nor U3261 (N_3261,N_818,N_520);
xnor U3262 (N_3262,N_891,N_75);
xor U3263 (N_3263,N_1493,N_945);
xor U3264 (N_3264,N_427,N_456);
xor U3265 (N_3265,N_1208,N_665);
or U3266 (N_3266,N_1931,N_1500);
nor U3267 (N_3267,N_1235,N_1854);
and U3268 (N_3268,N_967,N_1169);
nor U3269 (N_3269,N_1805,N_1988);
nor U3270 (N_3270,N_968,N_275);
nand U3271 (N_3271,N_1417,N_1948);
xnor U3272 (N_3272,N_720,N_767);
nor U3273 (N_3273,N_41,N_1168);
xor U3274 (N_3274,N_1402,N_628);
nor U3275 (N_3275,N_426,N_1137);
nor U3276 (N_3276,N_732,N_1357);
and U3277 (N_3277,N_930,N_1998);
nor U3278 (N_3278,N_814,N_32);
nand U3279 (N_3279,N_704,N_1879);
xnor U3280 (N_3280,N_1188,N_1064);
nand U3281 (N_3281,N_476,N_41);
xnor U3282 (N_3282,N_503,N_505);
and U3283 (N_3283,N_1526,N_262);
nor U3284 (N_3284,N_1438,N_821);
or U3285 (N_3285,N_1172,N_1574);
and U3286 (N_3286,N_104,N_1785);
nand U3287 (N_3287,N_701,N_359);
nand U3288 (N_3288,N_1914,N_848);
and U3289 (N_3289,N_1908,N_192);
and U3290 (N_3290,N_1466,N_402);
nand U3291 (N_3291,N_1185,N_1997);
nand U3292 (N_3292,N_1436,N_1074);
and U3293 (N_3293,N_411,N_1273);
nand U3294 (N_3294,N_962,N_1114);
and U3295 (N_3295,N_1725,N_1569);
xnor U3296 (N_3296,N_1877,N_681);
nand U3297 (N_3297,N_116,N_210);
nand U3298 (N_3298,N_1296,N_1773);
xor U3299 (N_3299,N_928,N_728);
or U3300 (N_3300,N_1654,N_787);
nor U3301 (N_3301,N_1861,N_1884);
xor U3302 (N_3302,N_1345,N_974);
or U3303 (N_3303,N_1492,N_481);
xor U3304 (N_3304,N_162,N_264);
or U3305 (N_3305,N_1926,N_1968);
or U3306 (N_3306,N_1605,N_446);
nand U3307 (N_3307,N_972,N_344);
nand U3308 (N_3308,N_590,N_1873);
or U3309 (N_3309,N_1721,N_1698);
or U3310 (N_3310,N_313,N_1056);
xor U3311 (N_3311,N_42,N_420);
and U3312 (N_3312,N_344,N_1828);
and U3313 (N_3313,N_77,N_315);
xor U3314 (N_3314,N_1053,N_958);
and U3315 (N_3315,N_1653,N_123);
nor U3316 (N_3316,N_1287,N_703);
and U3317 (N_3317,N_594,N_475);
or U3318 (N_3318,N_635,N_883);
and U3319 (N_3319,N_1109,N_1144);
xor U3320 (N_3320,N_1737,N_1509);
xnor U3321 (N_3321,N_623,N_1261);
nor U3322 (N_3322,N_780,N_1881);
and U3323 (N_3323,N_942,N_93);
nor U3324 (N_3324,N_246,N_962);
or U3325 (N_3325,N_1682,N_199);
and U3326 (N_3326,N_639,N_1382);
or U3327 (N_3327,N_1971,N_697);
and U3328 (N_3328,N_1286,N_1991);
xor U3329 (N_3329,N_1933,N_1375);
or U3330 (N_3330,N_1426,N_1580);
xor U3331 (N_3331,N_653,N_1049);
or U3332 (N_3332,N_888,N_1694);
nor U3333 (N_3333,N_1673,N_920);
xor U3334 (N_3334,N_955,N_1291);
or U3335 (N_3335,N_1235,N_1774);
nand U3336 (N_3336,N_1553,N_1757);
and U3337 (N_3337,N_574,N_557);
or U3338 (N_3338,N_1846,N_711);
and U3339 (N_3339,N_1990,N_376);
nor U3340 (N_3340,N_1795,N_406);
nand U3341 (N_3341,N_1481,N_20);
xor U3342 (N_3342,N_1902,N_110);
or U3343 (N_3343,N_1032,N_1672);
or U3344 (N_3344,N_383,N_1876);
xor U3345 (N_3345,N_1428,N_352);
nor U3346 (N_3346,N_69,N_1416);
nor U3347 (N_3347,N_1738,N_1377);
and U3348 (N_3348,N_433,N_1537);
and U3349 (N_3349,N_1446,N_279);
xnor U3350 (N_3350,N_1388,N_1709);
nand U3351 (N_3351,N_564,N_1500);
and U3352 (N_3352,N_515,N_311);
nor U3353 (N_3353,N_1166,N_1248);
and U3354 (N_3354,N_1688,N_129);
nand U3355 (N_3355,N_447,N_1373);
nand U3356 (N_3356,N_1200,N_448);
xor U3357 (N_3357,N_1258,N_1324);
and U3358 (N_3358,N_514,N_1967);
nand U3359 (N_3359,N_556,N_1200);
xor U3360 (N_3360,N_1537,N_676);
or U3361 (N_3361,N_847,N_1666);
nand U3362 (N_3362,N_974,N_1535);
or U3363 (N_3363,N_1173,N_1238);
nor U3364 (N_3364,N_1241,N_363);
or U3365 (N_3365,N_863,N_1888);
nand U3366 (N_3366,N_46,N_624);
or U3367 (N_3367,N_827,N_1966);
or U3368 (N_3368,N_510,N_1808);
xnor U3369 (N_3369,N_1402,N_1285);
nand U3370 (N_3370,N_287,N_1404);
and U3371 (N_3371,N_1603,N_1444);
nor U3372 (N_3372,N_8,N_1048);
xnor U3373 (N_3373,N_1196,N_1518);
nor U3374 (N_3374,N_1407,N_812);
or U3375 (N_3375,N_1650,N_331);
nor U3376 (N_3376,N_778,N_1194);
or U3377 (N_3377,N_1479,N_933);
xnor U3378 (N_3378,N_1166,N_1345);
nand U3379 (N_3379,N_315,N_659);
nand U3380 (N_3380,N_1146,N_321);
nor U3381 (N_3381,N_1979,N_1117);
nand U3382 (N_3382,N_907,N_686);
or U3383 (N_3383,N_767,N_1572);
and U3384 (N_3384,N_1643,N_159);
nand U3385 (N_3385,N_1516,N_930);
and U3386 (N_3386,N_1224,N_1281);
and U3387 (N_3387,N_666,N_1427);
and U3388 (N_3388,N_835,N_1131);
xnor U3389 (N_3389,N_671,N_1573);
nor U3390 (N_3390,N_1745,N_1719);
xor U3391 (N_3391,N_607,N_326);
or U3392 (N_3392,N_840,N_1582);
xor U3393 (N_3393,N_1350,N_522);
or U3394 (N_3394,N_1126,N_1476);
nor U3395 (N_3395,N_1192,N_135);
nand U3396 (N_3396,N_1893,N_502);
xnor U3397 (N_3397,N_1161,N_35);
nand U3398 (N_3398,N_805,N_1239);
nand U3399 (N_3399,N_1953,N_812);
and U3400 (N_3400,N_475,N_365);
xnor U3401 (N_3401,N_537,N_996);
nor U3402 (N_3402,N_92,N_1109);
nor U3403 (N_3403,N_1521,N_1571);
xor U3404 (N_3404,N_272,N_1514);
or U3405 (N_3405,N_1346,N_1882);
nand U3406 (N_3406,N_338,N_1196);
and U3407 (N_3407,N_1635,N_1074);
nor U3408 (N_3408,N_1685,N_923);
and U3409 (N_3409,N_449,N_1332);
nor U3410 (N_3410,N_776,N_270);
and U3411 (N_3411,N_204,N_508);
xnor U3412 (N_3412,N_447,N_1175);
or U3413 (N_3413,N_117,N_141);
nor U3414 (N_3414,N_1548,N_423);
xnor U3415 (N_3415,N_1188,N_873);
nor U3416 (N_3416,N_21,N_1381);
xor U3417 (N_3417,N_751,N_1386);
xor U3418 (N_3418,N_1063,N_475);
and U3419 (N_3419,N_677,N_1182);
nand U3420 (N_3420,N_330,N_661);
xnor U3421 (N_3421,N_397,N_628);
nor U3422 (N_3422,N_1396,N_1461);
nor U3423 (N_3423,N_102,N_134);
xor U3424 (N_3424,N_673,N_1276);
xor U3425 (N_3425,N_643,N_1658);
nand U3426 (N_3426,N_1513,N_1399);
xor U3427 (N_3427,N_758,N_735);
xor U3428 (N_3428,N_1379,N_47);
xnor U3429 (N_3429,N_500,N_741);
nand U3430 (N_3430,N_1563,N_1715);
nor U3431 (N_3431,N_1877,N_1268);
nor U3432 (N_3432,N_607,N_1919);
or U3433 (N_3433,N_604,N_117);
nor U3434 (N_3434,N_1906,N_1614);
xnor U3435 (N_3435,N_636,N_577);
xor U3436 (N_3436,N_1477,N_505);
nor U3437 (N_3437,N_927,N_312);
xor U3438 (N_3438,N_403,N_1355);
and U3439 (N_3439,N_1196,N_1960);
nor U3440 (N_3440,N_480,N_897);
or U3441 (N_3441,N_576,N_1719);
or U3442 (N_3442,N_980,N_1753);
nor U3443 (N_3443,N_1644,N_1174);
xnor U3444 (N_3444,N_680,N_669);
nand U3445 (N_3445,N_327,N_1489);
or U3446 (N_3446,N_1524,N_1788);
nor U3447 (N_3447,N_965,N_1821);
and U3448 (N_3448,N_501,N_1212);
nand U3449 (N_3449,N_1479,N_1229);
or U3450 (N_3450,N_1275,N_1103);
xor U3451 (N_3451,N_999,N_1593);
or U3452 (N_3452,N_241,N_1044);
or U3453 (N_3453,N_80,N_959);
nand U3454 (N_3454,N_1927,N_603);
and U3455 (N_3455,N_1169,N_1728);
and U3456 (N_3456,N_829,N_537);
xor U3457 (N_3457,N_632,N_219);
or U3458 (N_3458,N_576,N_535);
or U3459 (N_3459,N_935,N_785);
xor U3460 (N_3460,N_375,N_1851);
xor U3461 (N_3461,N_1443,N_737);
nor U3462 (N_3462,N_328,N_1657);
or U3463 (N_3463,N_1118,N_1307);
xor U3464 (N_3464,N_747,N_1818);
xnor U3465 (N_3465,N_1202,N_1123);
and U3466 (N_3466,N_1590,N_1213);
and U3467 (N_3467,N_997,N_582);
nor U3468 (N_3468,N_149,N_260);
and U3469 (N_3469,N_1905,N_1162);
nor U3470 (N_3470,N_333,N_1086);
xor U3471 (N_3471,N_603,N_9);
nor U3472 (N_3472,N_344,N_1961);
xnor U3473 (N_3473,N_576,N_1750);
nor U3474 (N_3474,N_585,N_1175);
xnor U3475 (N_3475,N_1835,N_1774);
xor U3476 (N_3476,N_1365,N_128);
and U3477 (N_3477,N_845,N_1642);
and U3478 (N_3478,N_504,N_1307);
or U3479 (N_3479,N_1410,N_1392);
nand U3480 (N_3480,N_494,N_1679);
nand U3481 (N_3481,N_404,N_836);
nand U3482 (N_3482,N_329,N_514);
or U3483 (N_3483,N_305,N_311);
and U3484 (N_3484,N_784,N_760);
xnor U3485 (N_3485,N_1769,N_39);
nand U3486 (N_3486,N_216,N_1483);
nor U3487 (N_3487,N_452,N_698);
nand U3488 (N_3488,N_1556,N_693);
xnor U3489 (N_3489,N_476,N_607);
and U3490 (N_3490,N_773,N_1917);
nand U3491 (N_3491,N_1741,N_8);
or U3492 (N_3492,N_1474,N_1193);
or U3493 (N_3493,N_376,N_963);
nand U3494 (N_3494,N_1895,N_918);
or U3495 (N_3495,N_1674,N_50);
and U3496 (N_3496,N_1775,N_123);
or U3497 (N_3497,N_1492,N_1841);
xnor U3498 (N_3498,N_1022,N_670);
or U3499 (N_3499,N_1732,N_1484);
nor U3500 (N_3500,N_596,N_1006);
xor U3501 (N_3501,N_241,N_516);
and U3502 (N_3502,N_1834,N_556);
xor U3503 (N_3503,N_722,N_561);
xnor U3504 (N_3504,N_1999,N_83);
nor U3505 (N_3505,N_338,N_1460);
xnor U3506 (N_3506,N_702,N_982);
or U3507 (N_3507,N_1685,N_66);
nand U3508 (N_3508,N_1405,N_1282);
nor U3509 (N_3509,N_837,N_614);
nor U3510 (N_3510,N_1042,N_1343);
or U3511 (N_3511,N_1503,N_405);
and U3512 (N_3512,N_1372,N_452);
xnor U3513 (N_3513,N_1015,N_330);
nor U3514 (N_3514,N_21,N_1681);
nand U3515 (N_3515,N_224,N_1550);
and U3516 (N_3516,N_1170,N_1363);
and U3517 (N_3517,N_1414,N_851);
or U3518 (N_3518,N_449,N_1535);
nand U3519 (N_3519,N_591,N_1617);
xnor U3520 (N_3520,N_589,N_1549);
and U3521 (N_3521,N_182,N_1756);
and U3522 (N_3522,N_1694,N_265);
or U3523 (N_3523,N_960,N_148);
nand U3524 (N_3524,N_465,N_1827);
xor U3525 (N_3525,N_553,N_634);
and U3526 (N_3526,N_1536,N_1246);
nor U3527 (N_3527,N_240,N_387);
nand U3528 (N_3528,N_1534,N_1147);
nor U3529 (N_3529,N_1382,N_447);
nor U3530 (N_3530,N_1595,N_1072);
nand U3531 (N_3531,N_582,N_988);
or U3532 (N_3532,N_425,N_1876);
or U3533 (N_3533,N_1323,N_849);
nor U3534 (N_3534,N_919,N_286);
and U3535 (N_3535,N_1906,N_297);
xor U3536 (N_3536,N_1524,N_254);
nand U3537 (N_3537,N_447,N_1114);
nor U3538 (N_3538,N_686,N_372);
and U3539 (N_3539,N_87,N_1364);
nor U3540 (N_3540,N_1929,N_355);
xnor U3541 (N_3541,N_260,N_606);
nor U3542 (N_3542,N_57,N_1099);
nor U3543 (N_3543,N_1426,N_1929);
xnor U3544 (N_3544,N_1396,N_1774);
xor U3545 (N_3545,N_1962,N_1411);
nand U3546 (N_3546,N_1422,N_561);
nor U3547 (N_3547,N_276,N_1072);
nand U3548 (N_3548,N_1809,N_1119);
or U3549 (N_3549,N_1472,N_1881);
and U3550 (N_3550,N_134,N_1681);
nor U3551 (N_3551,N_1700,N_1269);
nand U3552 (N_3552,N_604,N_1066);
or U3553 (N_3553,N_0,N_1776);
and U3554 (N_3554,N_1511,N_8);
or U3555 (N_3555,N_804,N_272);
xnor U3556 (N_3556,N_260,N_668);
and U3557 (N_3557,N_1880,N_1778);
nor U3558 (N_3558,N_1778,N_72);
nor U3559 (N_3559,N_854,N_1172);
nor U3560 (N_3560,N_42,N_1874);
nor U3561 (N_3561,N_581,N_884);
and U3562 (N_3562,N_1580,N_1175);
xnor U3563 (N_3563,N_1918,N_119);
and U3564 (N_3564,N_997,N_189);
and U3565 (N_3565,N_626,N_110);
nand U3566 (N_3566,N_1878,N_88);
and U3567 (N_3567,N_713,N_1859);
or U3568 (N_3568,N_157,N_472);
xnor U3569 (N_3569,N_1917,N_159);
and U3570 (N_3570,N_184,N_639);
nand U3571 (N_3571,N_214,N_721);
xnor U3572 (N_3572,N_640,N_1748);
and U3573 (N_3573,N_564,N_1087);
nand U3574 (N_3574,N_1252,N_1481);
or U3575 (N_3575,N_1181,N_1094);
nor U3576 (N_3576,N_1278,N_123);
xor U3577 (N_3577,N_394,N_1489);
nor U3578 (N_3578,N_469,N_1171);
nor U3579 (N_3579,N_1578,N_1237);
nand U3580 (N_3580,N_587,N_1122);
xor U3581 (N_3581,N_464,N_536);
nor U3582 (N_3582,N_818,N_1969);
and U3583 (N_3583,N_988,N_1185);
and U3584 (N_3584,N_490,N_1803);
or U3585 (N_3585,N_1986,N_1500);
nand U3586 (N_3586,N_845,N_105);
nor U3587 (N_3587,N_1883,N_1218);
xor U3588 (N_3588,N_1378,N_1779);
or U3589 (N_3589,N_502,N_595);
xnor U3590 (N_3590,N_1727,N_1614);
nand U3591 (N_3591,N_966,N_163);
nor U3592 (N_3592,N_1402,N_1980);
and U3593 (N_3593,N_192,N_1456);
nand U3594 (N_3594,N_127,N_459);
nand U3595 (N_3595,N_1575,N_650);
or U3596 (N_3596,N_1899,N_1632);
and U3597 (N_3597,N_1745,N_643);
and U3598 (N_3598,N_120,N_846);
or U3599 (N_3599,N_1546,N_1289);
nor U3600 (N_3600,N_170,N_37);
xnor U3601 (N_3601,N_788,N_828);
nand U3602 (N_3602,N_922,N_402);
nor U3603 (N_3603,N_852,N_1627);
xnor U3604 (N_3604,N_1567,N_1825);
xor U3605 (N_3605,N_157,N_1387);
nand U3606 (N_3606,N_43,N_1879);
nor U3607 (N_3607,N_1471,N_1874);
xor U3608 (N_3608,N_1360,N_1025);
xnor U3609 (N_3609,N_1489,N_586);
nor U3610 (N_3610,N_1529,N_1224);
xnor U3611 (N_3611,N_1744,N_467);
and U3612 (N_3612,N_1995,N_484);
nand U3613 (N_3613,N_361,N_551);
and U3614 (N_3614,N_1042,N_1172);
or U3615 (N_3615,N_1561,N_1199);
and U3616 (N_3616,N_852,N_1581);
or U3617 (N_3617,N_1015,N_1939);
and U3618 (N_3618,N_1773,N_377);
or U3619 (N_3619,N_390,N_442);
and U3620 (N_3620,N_1808,N_119);
and U3621 (N_3621,N_1488,N_527);
xnor U3622 (N_3622,N_1392,N_10);
and U3623 (N_3623,N_1139,N_790);
or U3624 (N_3624,N_1494,N_1526);
or U3625 (N_3625,N_1760,N_1112);
nand U3626 (N_3626,N_587,N_53);
xnor U3627 (N_3627,N_1,N_262);
nor U3628 (N_3628,N_1166,N_275);
or U3629 (N_3629,N_480,N_543);
or U3630 (N_3630,N_1421,N_1355);
nand U3631 (N_3631,N_964,N_1448);
and U3632 (N_3632,N_642,N_1286);
xor U3633 (N_3633,N_331,N_119);
and U3634 (N_3634,N_645,N_135);
xor U3635 (N_3635,N_689,N_1675);
and U3636 (N_3636,N_1554,N_1424);
and U3637 (N_3637,N_936,N_1735);
nor U3638 (N_3638,N_1340,N_715);
and U3639 (N_3639,N_797,N_941);
nand U3640 (N_3640,N_191,N_228);
nand U3641 (N_3641,N_786,N_1293);
and U3642 (N_3642,N_1896,N_1620);
nand U3643 (N_3643,N_1991,N_1994);
nand U3644 (N_3644,N_110,N_1237);
nor U3645 (N_3645,N_1379,N_624);
or U3646 (N_3646,N_847,N_33);
and U3647 (N_3647,N_1940,N_56);
nor U3648 (N_3648,N_1268,N_472);
or U3649 (N_3649,N_1029,N_1741);
nand U3650 (N_3650,N_88,N_609);
nand U3651 (N_3651,N_1291,N_1755);
nand U3652 (N_3652,N_366,N_123);
nor U3653 (N_3653,N_1988,N_901);
nor U3654 (N_3654,N_1627,N_350);
or U3655 (N_3655,N_316,N_1575);
nand U3656 (N_3656,N_189,N_1940);
nor U3657 (N_3657,N_302,N_1341);
or U3658 (N_3658,N_1499,N_684);
xnor U3659 (N_3659,N_1040,N_11);
nor U3660 (N_3660,N_1258,N_520);
or U3661 (N_3661,N_222,N_1402);
or U3662 (N_3662,N_889,N_1782);
xnor U3663 (N_3663,N_413,N_959);
and U3664 (N_3664,N_1635,N_1966);
nand U3665 (N_3665,N_1600,N_713);
xnor U3666 (N_3666,N_1776,N_147);
or U3667 (N_3667,N_1386,N_1512);
or U3668 (N_3668,N_553,N_557);
or U3669 (N_3669,N_623,N_441);
or U3670 (N_3670,N_474,N_241);
xor U3671 (N_3671,N_1394,N_294);
nor U3672 (N_3672,N_978,N_831);
xnor U3673 (N_3673,N_1556,N_1697);
and U3674 (N_3674,N_970,N_54);
and U3675 (N_3675,N_911,N_90);
xnor U3676 (N_3676,N_701,N_1284);
xor U3677 (N_3677,N_112,N_1467);
or U3678 (N_3678,N_1995,N_1329);
nand U3679 (N_3679,N_1057,N_1374);
and U3680 (N_3680,N_1629,N_50);
and U3681 (N_3681,N_1811,N_1844);
or U3682 (N_3682,N_1321,N_1187);
and U3683 (N_3683,N_509,N_123);
nor U3684 (N_3684,N_1770,N_1996);
and U3685 (N_3685,N_957,N_693);
or U3686 (N_3686,N_995,N_1397);
nand U3687 (N_3687,N_504,N_1339);
nor U3688 (N_3688,N_869,N_880);
nor U3689 (N_3689,N_476,N_1781);
nor U3690 (N_3690,N_840,N_983);
nor U3691 (N_3691,N_1023,N_1466);
nor U3692 (N_3692,N_1428,N_1683);
nor U3693 (N_3693,N_414,N_1270);
or U3694 (N_3694,N_357,N_645);
nor U3695 (N_3695,N_1889,N_1028);
xor U3696 (N_3696,N_519,N_473);
nand U3697 (N_3697,N_57,N_1873);
nor U3698 (N_3698,N_854,N_934);
and U3699 (N_3699,N_1246,N_1907);
nand U3700 (N_3700,N_1877,N_817);
nand U3701 (N_3701,N_308,N_1949);
xnor U3702 (N_3702,N_1793,N_1861);
and U3703 (N_3703,N_1024,N_1605);
nand U3704 (N_3704,N_455,N_1794);
nand U3705 (N_3705,N_1014,N_123);
and U3706 (N_3706,N_686,N_967);
nand U3707 (N_3707,N_77,N_639);
nand U3708 (N_3708,N_989,N_1005);
xnor U3709 (N_3709,N_1005,N_1367);
nand U3710 (N_3710,N_1618,N_986);
or U3711 (N_3711,N_676,N_1723);
or U3712 (N_3712,N_1612,N_1768);
or U3713 (N_3713,N_1071,N_1817);
and U3714 (N_3714,N_830,N_1900);
or U3715 (N_3715,N_981,N_270);
or U3716 (N_3716,N_1326,N_1218);
xor U3717 (N_3717,N_161,N_134);
nor U3718 (N_3718,N_381,N_1288);
xor U3719 (N_3719,N_219,N_821);
nand U3720 (N_3720,N_739,N_1708);
and U3721 (N_3721,N_782,N_645);
nand U3722 (N_3722,N_239,N_797);
nand U3723 (N_3723,N_754,N_1567);
and U3724 (N_3724,N_267,N_1155);
nor U3725 (N_3725,N_1349,N_1220);
nand U3726 (N_3726,N_717,N_1043);
and U3727 (N_3727,N_1111,N_392);
or U3728 (N_3728,N_1707,N_414);
xor U3729 (N_3729,N_871,N_1094);
nand U3730 (N_3730,N_1121,N_1552);
nand U3731 (N_3731,N_1289,N_1802);
and U3732 (N_3732,N_831,N_1385);
nor U3733 (N_3733,N_1667,N_881);
nand U3734 (N_3734,N_35,N_1203);
and U3735 (N_3735,N_1900,N_875);
and U3736 (N_3736,N_1666,N_284);
and U3737 (N_3737,N_1701,N_690);
xor U3738 (N_3738,N_1489,N_539);
or U3739 (N_3739,N_439,N_461);
and U3740 (N_3740,N_287,N_712);
nand U3741 (N_3741,N_51,N_528);
or U3742 (N_3742,N_381,N_1793);
nand U3743 (N_3743,N_238,N_200);
and U3744 (N_3744,N_395,N_337);
or U3745 (N_3745,N_1530,N_1888);
nor U3746 (N_3746,N_1740,N_599);
or U3747 (N_3747,N_1000,N_1630);
xor U3748 (N_3748,N_1172,N_870);
nor U3749 (N_3749,N_1135,N_1471);
nand U3750 (N_3750,N_999,N_1105);
xor U3751 (N_3751,N_1601,N_735);
xor U3752 (N_3752,N_512,N_1562);
and U3753 (N_3753,N_1725,N_1036);
nand U3754 (N_3754,N_815,N_654);
or U3755 (N_3755,N_1394,N_1112);
or U3756 (N_3756,N_723,N_95);
nor U3757 (N_3757,N_356,N_1342);
nor U3758 (N_3758,N_490,N_865);
and U3759 (N_3759,N_1216,N_1943);
nand U3760 (N_3760,N_1870,N_1607);
xnor U3761 (N_3761,N_1359,N_531);
and U3762 (N_3762,N_1055,N_168);
xor U3763 (N_3763,N_465,N_734);
nor U3764 (N_3764,N_641,N_1170);
nand U3765 (N_3765,N_655,N_1186);
nand U3766 (N_3766,N_1689,N_1403);
xor U3767 (N_3767,N_158,N_328);
or U3768 (N_3768,N_815,N_794);
and U3769 (N_3769,N_1885,N_1567);
nand U3770 (N_3770,N_568,N_1049);
xnor U3771 (N_3771,N_1048,N_1221);
nor U3772 (N_3772,N_1665,N_1851);
and U3773 (N_3773,N_428,N_1290);
xnor U3774 (N_3774,N_1223,N_1337);
nand U3775 (N_3775,N_1197,N_168);
nand U3776 (N_3776,N_1327,N_687);
xor U3777 (N_3777,N_550,N_756);
nor U3778 (N_3778,N_361,N_1174);
and U3779 (N_3779,N_1367,N_149);
xor U3780 (N_3780,N_1622,N_56);
nand U3781 (N_3781,N_1400,N_472);
nand U3782 (N_3782,N_1180,N_1184);
nand U3783 (N_3783,N_1948,N_1257);
nand U3784 (N_3784,N_351,N_49);
nand U3785 (N_3785,N_36,N_995);
and U3786 (N_3786,N_1454,N_614);
nand U3787 (N_3787,N_1284,N_1856);
xnor U3788 (N_3788,N_1277,N_1321);
and U3789 (N_3789,N_245,N_438);
xor U3790 (N_3790,N_786,N_1336);
xor U3791 (N_3791,N_1842,N_444);
or U3792 (N_3792,N_631,N_1031);
nand U3793 (N_3793,N_1067,N_53);
or U3794 (N_3794,N_1048,N_1060);
nor U3795 (N_3795,N_545,N_245);
xnor U3796 (N_3796,N_800,N_104);
xnor U3797 (N_3797,N_1686,N_624);
and U3798 (N_3798,N_1648,N_1204);
nor U3799 (N_3799,N_663,N_900);
xnor U3800 (N_3800,N_1245,N_1225);
nand U3801 (N_3801,N_421,N_192);
and U3802 (N_3802,N_1063,N_193);
nand U3803 (N_3803,N_1641,N_391);
nand U3804 (N_3804,N_187,N_716);
nand U3805 (N_3805,N_671,N_1044);
or U3806 (N_3806,N_864,N_1004);
nand U3807 (N_3807,N_582,N_223);
nor U3808 (N_3808,N_1441,N_1688);
nor U3809 (N_3809,N_1900,N_523);
nand U3810 (N_3810,N_570,N_936);
xnor U3811 (N_3811,N_1148,N_1855);
nor U3812 (N_3812,N_1181,N_1021);
xor U3813 (N_3813,N_750,N_1578);
and U3814 (N_3814,N_1095,N_1087);
nand U3815 (N_3815,N_1523,N_1726);
nor U3816 (N_3816,N_1337,N_1665);
nor U3817 (N_3817,N_137,N_1834);
xor U3818 (N_3818,N_93,N_317);
nand U3819 (N_3819,N_674,N_1218);
and U3820 (N_3820,N_13,N_1107);
nand U3821 (N_3821,N_1338,N_18);
or U3822 (N_3822,N_65,N_185);
nand U3823 (N_3823,N_1710,N_1101);
xor U3824 (N_3824,N_928,N_432);
nand U3825 (N_3825,N_1583,N_1397);
and U3826 (N_3826,N_884,N_1083);
nand U3827 (N_3827,N_947,N_860);
nor U3828 (N_3828,N_862,N_759);
nand U3829 (N_3829,N_188,N_1440);
or U3830 (N_3830,N_520,N_532);
nor U3831 (N_3831,N_1687,N_1294);
xnor U3832 (N_3832,N_1860,N_154);
and U3833 (N_3833,N_1097,N_1724);
and U3834 (N_3834,N_583,N_626);
nand U3835 (N_3835,N_1727,N_1731);
or U3836 (N_3836,N_1507,N_216);
xor U3837 (N_3837,N_573,N_1553);
nor U3838 (N_3838,N_1150,N_369);
nand U3839 (N_3839,N_504,N_1204);
nand U3840 (N_3840,N_743,N_1422);
nor U3841 (N_3841,N_1951,N_32);
xnor U3842 (N_3842,N_167,N_387);
xnor U3843 (N_3843,N_666,N_1696);
or U3844 (N_3844,N_1166,N_1944);
and U3845 (N_3845,N_706,N_740);
and U3846 (N_3846,N_1723,N_1938);
nor U3847 (N_3847,N_1375,N_213);
nand U3848 (N_3848,N_1739,N_602);
nand U3849 (N_3849,N_1162,N_1384);
nand U3850 (N_3850,N_323,N_1273);
and U3851 (N_3851,N_1296,N_546);
and U3852 (N_3852,N_888,N_358);
nor U3853 (N_3853,N_1665,N_201);
nand U3854 (N_3854,N_88,N_1789);
xnor U3855 (N_3855,N_1350,N_1498);
nand U3856 (N_3856,N_163,N_1807);
or U3857 (N_3857,N_1759,N_373);
nand U3858 (N_3858,N_1521,N_1115);
or U3859 (N_3859,N_1736,N_1269);
xnor U3860 (N_3860,N_1100,N_308);
xnor U3861 (N_3861,N_1806,N_1015);
nor U3862 (N_3862,N_772,N_1519);
nor U3863 (N_3863,N_576,N_1322);
xnor U3864 (N_3864,N_1976,N_1607);
and U3865 (N_3865,N_1492,N_828);
or U3866 (N_3866,N_283,N_1596);
xor U3867 (N_3867,N_809,N_349);
xnor U3868 (N_3868,N_1492,N_354);
or U3869 (N_3869,N_1822,N_441);
or U3870 (N_3870,N_439,N_1379);
or U3871 (N_3871,N_584,N_1741);
nor U3872 (N_3872,N_861,N_372);
and U3873 (N_3873,N_578,N_1462);
and U3874 (N_3874,N_344,N_400);
or U3875 (N_3875,N_311,N_173);
and U3876 (N_3876,N_1592,N_500);
nand U3877 (N_3877,N_1244,N_1667);
xor U3878 (N_3878,N_1421,N_106);
and U3879 (N_3879,N_1452,N_1988);
nand U3880 (N_3880,N_499,N_1169);
xnor U3881 (N_3881,N_1697,N_136);
xnor U3882 (N_3882,N_1955,N_1213);
and U3883 (N_3883,N_627,N_751);
and U3884 (N_3884,N_1240,N_1206);
and U3885 (N_3885,N_319,N_1158);
xor U3886 (N_3886,N_19,N_1985);
xor U3887 (N_3887,N_49,N_470);
nor U3888 (N_3888,N_923,N_1350);
or U3889 (N_3889,N_1005,N_1536);
or U3890 (N_3890,N_1675,N_1664);
nor U3891 (N_3891,N_1297,N_1230);
nor U3892 (N_3892,N_461,N_250);
nand U3893 (N_3893,N_1145,N_1830);
and U3894 (N_3894,N_1686,N_675);
or U3895 (N_3895,N_286,N_272);
or U3896 (N_3896,N_1557,N_877);
and U3897 (N_3897,N_1655,N_440);
and U3898 (N_3898,N_1314,N_1109);
xor U3899 (N_3899,N_341,N_767);
or U3900 (N_3900,N_1919,N_962);
xor U3901 (N_3901,N_1442,N_1328);
nor U3902 (N_3902,N_1465,N_226);
xor U3903 (N_3903,N_1742,N_1353);
or U3904 (N_3904,N_145,N_1410);
nor U3905 (N_3905,N_1982,N_489);
nor U3906 (N_3906,N_1651,N_1370);
xor U3907 (N_3907,N_1409,N_1406);
and U3908 (N_3908,N_1432,N_1031);
and U3909 (N_3909,N_426,N_568);
and U3910 (N_3910,N_643,N_490);
nand U3911 (N_3911,N_1607,N_1126);
nor U3912 (N_3912,N_1861,N_1246);
nand U3913 (N_3913,N_397,N_330);
nor U3914 (N_3914,N_4,N_991);
and U3915 (N_3915,N_288,N_1459);
xnor U3916 (N_3916,N_1167,N_520);
nand U3917 (N_3917,N_1161,N_716);
xnor U3918 (N_3918,N_384,N_1020);
or U3919 (N_3919,N_233,N_1393);
or U3920 (N_3920,N_730,N_1264);
nor U3921 (N_3921,N_746,N_1887);
nor U3922 (N_3922,N_576,N_966);
nand U3923 (N_3923,N_326,N_38);
nand U3924 (N_3924,N_1828,N_975);
xor U3925 (N_3925,N_1318,N_1200);
nor U3926 (N_3926,N_607,N_61);
and U3927 (N_3927,N_366,N_1702);
or U3928 (N_3928,N_1466,N_249);
or U3929 (N_3929,N_1869,N_464);
and U3930 (N_3930,N_621,N_825);
nor U3931 (N_3931,N_772,N_258);
xnor U3932 (N_3932,N_168,N_913);
and U3933 (N_3933,N_1553,N_502);
xor U3934 (N_3934,N_46,N_1758);
or U3935 (N_3935,N_1738,N_690);
or U3936 (N_3936,N_511,N_121);
xnor U3937 (N_3937,N_737,N_1276);
nor U3938 (N_3938,N_436,N_1178);
nor U3939 (N_3939,N_1881,N_455);
and U3940 (N_3940,N_1196,N_1186);
or U3941 (N_3941,N_1588,N_1175);
or U3942 (N_3942,N_51,N_1693);
and U3943 (N_3943,N_476,N_1473);
or U3944 (N_3944,N_349,N_652);
nor U3945 (N_3945,N_1368,N_992);
xnor U3946 (N_3946,N_1340,N_1444);
or U3947 (N_3947,N_398,N_1202);
nor U3948 (N_3948,N_1332,N_287);
or U3949 (N_3949,N_1691,N_1725);
nor U3950 (N_3950,N_1294,N_898);
nor U3951 (N_3951,N_603,N_1089);
nor U3952 (N_3952,N_497,N_985);
and U3953 (N_3953,N_1013,N_1006);
or U3954 (N_3954,N_606,N_97);
and U3955 (N_3955,N_1061,N_1640);
or U3956 (N_3956,N_1930,N_942);
nand U3957 (N_3957,N_1408,N_1940);
nand U3958 (N_3958,N_92,N_400);
or U3959 (N_3959,N_872,N_474);
nand U3960 (N_3960,N_1702,N_1462);
nand U3961 (N_3961,N_1516,N_1446);
xor U3962 (N_3962,N_1462,N_768);
nor U3963 (N_3963,N_1560,N_860);
nand U3964 (N_3964,N_1723,N_1430);
nand U3965 (N_3965,N_55,N_985);
nand U3966 (N_3966,N_1050,N_485);
nand U3967 (N_3967,N_99,N_369);
xor U3968 (N_3968,N_545,N_470);
or U3969 (N_3969,N_588,N_1936);
nand U3970 (N_3970,N_996,N_1435);
xor U3971 (N_3971,N_846,N_712);
nor U3972 (N_3972,N_1325,N_1646);
or U3973 (N_3973,N_1042,N_1324);
nand U3974 (N_3974,N_830,N_65);
nor U3975 (N_3975,N_8,N_567);
and U3976 (N_3976,N_214,N_1763);
and U3977 (N_3977,N_204,N_1694);
and U3978 (N_3978,N_3,N_7);
nand U3979 (N_3979,N_414,N_1212);
and U3980 (N_3980,N_1644,N_1303);
nor U3981 (N_3981,N_822,N_406);
xor U3982 (N_3982,N_535,N_238);
or U3983 (N_3983,N_1832,N_312);
xnor U3984 (N_3984,N_893,N_1190);
nand U3985 (N_3985,N_1741,N_1325);
and U3986 (N_3986,N_1869,N_1305);
xnor U3987 (N_3987,N_1837,N_527);
or U3988 (N_3988,N_986,N_66);
nand U3989 (N_3989,N_21,N_1571);
or U3990 (N_3990,N_1132,N_1317);
nand U3991 (N_3991,N_439,N_504);
and U3992 (N_3992,N_1935,N_723);
and U3993 (N_3993,N_1295,N_321);
and U3994 (N_3994,N_1515,N_1464);
nand U3995 (N_3995,N_254,N_491);
xor U3996 (N_3996,N_1214,N_1049);
nand U3997 (N_3997,N_469,N_1048);
nor U3998 (N_3998,N_1785,N_306);
xor U3999 (N_3999,N_934,N_984);
nor U4000 (N_4000,N_3828,N_3905);
and U4001 (N_4001,N_2589,N_3133);
nand U4002 (N_4002,N_3648,N_3332);
and U4003 (N_4003,N_2311,N_2862);
xnor U4004 (N_4004,N_2312,N_3209);
nand U4005 (N_4005,N_2371,N_3459);
and U4006 (N_4006,N_2845,N_3678);
and U4007 (N_4007,N_2203,N_3812);
or U4008 (N_4008,N_2851,N_2536);
nand U4009 (N_4009,N_3617,N_3006);
or U4010 (N_4010,N_2650,N_3676);
and U4011 (N_4011,N_2766,N_2469);
nand U4012 (N_4012,N_2155,N_2901);
xor U4013 (N_4013,N_3119,N_3562);
or U4014 (N_4014,N_3137,N_2376);
and U4015 (N_4015,N_2979,N_2105);
or U4016 (N_4016,N_2359,N_2575);
nor U4017 (N_4017,N_2713,N_3699);
or U4018 (N_4018,N_3327,N_3789);
nor U4019 (N_4019,N_2738,N_3376);
nor U4020 (N_4020,N_3711,N_2982);
nor U4021 (N_4021,N_2206,N_2753);
nor U4022 (N_4022,N_3542,N_2926);
nor U4023 (N_4023,N_2246,N_2394);
nand U4024 (N_4024,N_2912,N_2864);
xnor U4025 (N_4025,N_3107,N_2240);
xnor U4026 (N_4026,N_3943,N_3819);
xor U4027 (N_4027,N_2603,N_3288);
nand U4028 (N_4028,N_2876,N_3419);
or U4029 (N_4029,N_2113,N_3055);
or U4030 (N_4030,N_3815,N_3216);
nand U4031 (N_4031,N_2762,N_3471);
nand U4032 (N_4032,N_3071,N_2387);
nor U4033 (N_4033,N_3974,N_3153);
nor U4034 (N_4034,N_3570,N_3810);
nand U4035 (N_4035,N_3040,N_2290);
xnor U4036 (N_4036,N_2721,N_3507);
and U4037 (N_4037,N_2159,N_2688);
or U4038 (N_4038,N_3840,N_3991);
xor U4039 (N_4039,N_3272,N_2625);
nand U4040 (N_4040,N_2365,N_3850);
nand U4041 (N_4041,N_3920,N_3410);
and U4042 (N_4042,N_2986,N_2509);
nor U4043 (N_4043,N_3377,N_2607);
xor U4044 (N_4044,N_3412,N_3702);
and U4045 (N_4045,N_3366,N_3929);
or U4046 (N_4046,N_2755,N_3132);
nor U4047 (N_4047,N_2343,N_3639);
or U4048 (N_4048,N_2435,N_3803);
or U4049 (N_4049,N_2128,N_3259);
xnor U4050 (N_4050,N_2570,N_3225);
and U4051 (N_4051,N_3844,N_3340);
nor U4052 (N_4052,N_3975,N_3039);
nand U4053 (N_4053,N_3664,N_3368);
and U4054 (N_4054,N_3933,N_2271);
or U4055 (N_4055,N_3169,N_2079);
and U4056 (N_4056,N_3827,N_2835);
or U4057 (N_4057,N_2855,N_2627);
nor U4058 (N_4058,N_2810,N_2141);
nand U4059 (N_4059,N_3788,N_2745);
nor U4060 (N_4060,N_3508,N_3056);
nor U4061 (N_4061,N_2213,N_3482);
and U4062 (N_4062,N_2187,N_3330);
or U4063 (N_4063,N_2587,N_2462);
xnor U4064 (N_4064,N_2396,N_2806);
and U4065 (N_4065,N_3045,N_3388);
or U4066 (N_4066,N_2668,N_2309);
nand U4067 (N_4067,N_3252,N_3506);
nor U4068 (N_4068,N_2406,N_3581);
and U4069 (N_4069,N_2891,N_2740);
nand U4070 (N_4070,N_3762,N_2545);
xor U4071 (N_4071,N_2730,N_2429);
nand U4072 (N_4072,N_2022,N_3020);
nor U4073 (N_4073,N_2774,N_2055);
nor U4074 (N_4074,N_3502,N_2634);
and U4075 (N_4075,N_3060,N_3644);
xor U4076 (N_4076,N_3158,N_3691);
xnor U4077 (N_4077,N_3761,N_3621);
nor U4078 (N_4078,N_3818,N_3725);
and U4079 (N_4079,N_3236,N_3282);
or U4080 (N_4080,N_2189,N_3737);
and U4081 (N_4081,N_2425,N_3050);
nand U4082 (N_4082,N_2940,N_2170);
nor U4083 (N_4083,N_2508,N_2484);
and U4084 (N_4084,N_3892,N_3426);
and U4085 (N_4085,N_2270,N_2599);
nor U4086 (N_4086,N_3635,N_2858);
and U4087 (N_4087,N_3199,N_2330);
nor U4088 (N_4088,N_2717,N_3888);
or U4089 (N_4089,N_2421,N_2499);
nand U4090 (N_4090,N_3479,N_2786);
or U4091 (N_4091,N_2586,N_2772);
nor U4092 (N_4092,N_3918,N_3363);
nor U4093 (N_4093,N_2355,N_2317);
nand U4094 (N_4094,N_3914,N_3928);
xor U4095 (N_4095,N_3014,N_3740);
xor U4096 (N_4096,N_2532,N_3290);
nor U4097 (N_4097,N_3806,N_2734);
nand U4098 (N_4098,N_2594,N_2856);
xor U4099 (N_4099,N_3972,N_2537);
nor U4100 (N_4100,N_2678,N_3160);
and U4101 (N_4101,N_2707,N_3626);
xnor U4102 (N_4102,N_2284,N_3628);
xor U4103 (N_4103,N_2682,N_3012);
xnor U4104 (N_4104,N_2705,N_2944);
nand U4105 (N_4105,N_3895,N_3643);
or U4106 (N_4106,N_3126,N_2943);
nand U4107 (N_4107,N_3183,N_3713);
and U4108 (N_4108,N_3596,N_2455);
nand U4109 (N_4109,N_3284,N_2087);
and U4110 (N_4110,N_2006,N_3712);
xor U4111 (N_4111,N_2889,N_2744);
xnor U4112 (N_4112,N_3666,N_2482);
and U4113 (N_4113,N_2520,N_2723);
and U4114 (N_4114,N_3609,N_2696);
and U4115 (N_4115,N_3960,N_3026);
nor U4116 (N_4116,N_3184,N_2779);
nor U4117 (N_4117,N_3470,N_2885);
or U4118 (N_4118,N_3605,N_2475);
or U4119 (N_4119,N_3215,N_3684);
nor U4120 (N_4120,N_2430,N_2631);
xnor U4121 (N_4121,N_2132,N_3155);
or U4122 (N_4122,N_2630,N_3683);
and U4123 (N_4123,N_3392,N_3662);
xor U4124 (N_4124,N_3099,N_2196);
nor U4125 (N_4125,N_3896,N_3487);
nor U4126 (N_4126,N_3075,N_2946);
or U4127 (N_4127,N_3015,N_3120);
and U4128 (N_4128,N_2528,N_2667);
or U4129 (N_4129,N_3401,N_2692);
and U4130 (N_4130,N_2572,N_2305);
or U4131 (N_4131,N_2641,N_3384);
xnor U4132 (N_4132,N_3185,N_3941);
nor U4133 (N_4133,N_3583,N_2934);
and U4134 (N_4134,N_3607,N_2236);
nor U4135 (N_4135,N_2465,N_2266);
nor U4136 (N_4136,N_3448,N_3886);
nand U4137 (N_4137,N_3496,N_3234);
xor U4138 (N_4138,N_3852,N_3395);
or U4139 (N_4139,N_2061,N_3457);
xor U4140 (N_4140,N_2057,N_3730);
or U4141 (N_4141,N_2837,N_2555);
or U4142 (N_4142,N_3976,N_2001);
nor U4143 (N_4143,N_3212,N_3394);
nand U4144 (N_4144,N_3266,N_3838);
or U4145 (N_4145,N_3357,N_2013);
nor U4146 (N_4146,N_3599,N_2714);
xor U4147 (N_4147,N_3224,N_3182);
xnor U4148 (N_4148,N_3880,N_3616);
nor U4149 (N_4149,N_3796,N_3531);
or U4150 (N_4150,N_3774,N_2582);
nand U4151 (N_4151,N_3343,N_2850);
and U4152 (N_4152,N_2989,N_3518);
and U4153 (N_4153,N_2231,N_2491);
nand U4154 (N_4154,N_3860,N_2296);
xnor U4155 (N_4155,N_3474,N_2951);
nor U4156 (N_4156,N_3032,N_3620);
and U4157 (N_4157,N_3592,N_2259);
nor U4158 (N_4158,N_3987,N_3522);
xor U4159 (N_4159,N_2281,N_2866);
xor U4160 (N_4160,N_3813,N_3795);
xnor U4161 (N_4161,N_2019,N_2732);
nor U4162 (N_4162,N_2158,N_2095);
xnor U4163 (N_4163,N_2872,N_2849);
xnor U4164 (N_4164,N_3980,N_2577);
nand U4165 (N_4165,N_3312,N_2910);
xor U4166 (N_4166,N_2511,N_2778);
nand U4167 (N_4167,N_3049,N_2291);
or U4168 (N_4168,N_3538,N_2632);
xor U4169 (N_4169,N_3858,N_3430);
nand U4170 (N_4170,N_3799,N_2971);
and U4171 (N_4171,N_2184,N_3865);
or U4172 (N_4172,N_2824,N_3841);
nor U4173 (N_4173,N_2743,N_2172);
xor U4174 (N_4174,N_2833,N_2210);
or U4175 (N_4175,N_3552,N_3792);
and U4176 (N_4176,N_2788,N_2892);
nand U4177 (N_4177,N_2268,N_2324);
and U4178 (N_4178,N_3708,N_3811);
xnor U4179 (N_4179,N_3686,N_2710);
xor U4180 (N_4180,N_2785,N_2412);
xor U4181 (N_4181,N_3206,N_2863);
or U4182 (N_4182,N_2925,N_3367);
xor U4183 (N_4183,N_2852,N_3491);
or U4184 (N_4184,N_2831,N_2453);
xnor U4185 (N_4185,N_3034,N_2193);
or U4186 (N_4186,N_2904,N_3629);
or U4187 (N_4187,N_2208,N_2226);
nand U4188 (N_4188,N_2777,N_3624);
or U4189 (N_4189,N_3951,N_3671);
xor U4190 (N_4190,N_2205,N_3217);
nand U4191 (N_4191,N_3362,N_2529);
or U4192 (N_4192,N_2563,N_3484);
and U4193 (N_4193,N_3189,N_2212);
nand U4194 (N_4194,N_3399,N_3842);
nand U4195 (N_4195,N_3753,N_2811);
and U4196 (N_4196,N_3724,N_2990);
or U4197 (N_4197,N_3391,N_3681);
nand U4198 (N_4198,N_2286,N_2816);
xnor U4199 (N_4199,N_2223,N_3735);
nor U4200 (N_4200,N_2662,N_3637);
nor U4201 (N_4201,N_2812,N_2331);
and U4202 (N_4202,N_2611,N_2922);
nand U4203 (N_4203,N_3196,N_2787);
xor U4204 (N_4204,N_3300,N_2722);
nor U4205 (N_4205,N_3510,N_2699);
or U4206 (N_4206,N_3660,N_3539);
or U4207 (N_4207,N_2823,N_3461);
xnor U4208 (N_4208,N_2685,N_2192);
xnor U4209 (N_4209,N_2257,N_3286);
and U4210 (N_4210,N_3279,N_2821);
nor U4211 (N_4211,N_3110,N_2558);
xor U4212 (N_4212,N_3024,N_2628);
nor U4213 (N_4213,N_3109,N_3339);
or U4214 (N_4214,N_3421,N_2794);
xor U4215 (N_4215,N_2334,N_2514);
xnor U4216 (N_4216,N_2372,N_3771);
and U4217 (N_4217,N_3897,N_3798);
nor U4218 (N_4218,N_3065,N_3521);
nor U4219 (N_4219,N_3054,N_3674);
nor U4220 (N_4220,N_2041,N_3543);
nor U4221 (N_4221,N_3988,N_3466);
or U4222 (N_4222,N_3115,N_3760);
or U4223 (N_4223,N_3105,N_2803);
and U4224 (N_4224,N_3128,N_2805);
nor U4225 (N_4225,N_3719,N_2551);
and U4226 (N_4226,N_3940,N_2742);
nor U4227 (N_4227,N_2115,N_3285);
nor U4228 (N_4228,N_3018,N_3499);
nand U4229 (N_4229,N_2588,N_2640);
xor U4230 (N_4230,N_2861,N_2434);
xnor U4231 (N_4231,N_2092,N_3190);
or U4232 (N_4232,N_2503,N_2790);
and U4233 (N_4233,N_3073,N_3064);
nor U4234 (N_4234,N_2679,N_3356);
or U4235 (N_4235,N_3764,N_3194);
or U4236 (N_4236,N_3067,N_2865);
xnor U4237 (N_4237,N_2693,N_3645);
nand U4238 (N_4238,N_3651,N_3910);
and U4239 (N_4239,N_3093,N_2617);
nand U4240 (N_4240,N_3047,N_2706);
nand U4241 (N_4241,N_2695,N_3335);
nand U4242 (N_4242,N_2671,N_3923);
nor U4243 (N_4243,N_2521,N_2496);
nand U4244 (N_4244,N_2486,N_3587);
xnor U4245 (N_4245,N_2201,N_2513);
xnor U4246 (N_4246,N_3350,N_3492);
nand U4247 (N_4247,N_3180,N_2065);
nor U4248 (N_4248,N_3966,N_3763);
nand U4249 (N_4249,N_3559,N_3453);
or U4250 (N_4250,N_2322,N_3211);
or U4251 (N_4251,N_2207,N_3038);
and U4252 (N_4252,N_2897,N_2183);
xor U4253 (N_4253,N_3334,N_2444);
xor U4254 (N_4254,N_3289,N_2568);
nor U4255 (N_4255,N_2357,N_2040);
xor U4256 (N_4256,N_2666,N_2302);
nor U4257 (N_4257,N_2255,N_3118);
nand U4258 (N_4258,N_2871,N_2523);
nor U4259 (N_4259,N_2052,N_3264);
or U4260 (N_4260,N_2538,N_3245);
xnor U4261 (N_4261,N_3879,N_2655);
or U4262 (N_4262,N_3728,N_2522);
xor U4263 (N_4263,N_3072,N_2659);
nor U4264 (N_4264,N_3834,N_3243);
and U4265 (N_4265,N_3536,N_2261);
nand U4266 (N_4266,N_3317,N_3125);
nor U4267 (N_4267,N_3917,N_3833);
xor U4268 (N_4268,N_3585,N_3823);
xnor U4269 (N_4269,N_3374,N_2746);
nand U4270 (N_4270,N_3454,N_3793);
xnor U4271 (N_4271,N_2029,N_3548);
and U4272 (N_4272,N_3240,N_2370);
and U4273 (N_4273,N_2450,N_2358);
nor U4274 (N_4274,N_3375,N_3573);
and U4275 (N_4275,N_2032,N_3705);
nand U4276 (N_4276,N_2163,N_3675);
or U4277 (N_4277,N_2166,N_3787);
or U4278 (N_4278,N_3992,N_3135);
or U4279 (N_4279,N_3292,N_3729);
nand U4280 (N_4280,N_2909,N_2451);
xnor U4281 (N_4281,N_2364,N_3501);
nor U4282 (N_4282,N_2756,N_2247);
xor U4283 (N_4283,N_3411,N_2088);
or U4284 (N_4284,N_2176,N_2410);
nor U4285 (N_4285,N_2648,N_2516);
nand U4286 (N_4286,N_2488,N_2843);
or U4287 (N_4287,N_3074,N_3561);
nor U4288 (N_4288,N_2340,N_2224);
and U4289 (N_4289,N_2842,N_2825);
and U4290 (N_4290,N_2325,N_3130);
nand U4291 (N_4291,N_2140,N_3385);
xnor U4292 (N_4292,N_3436,N_2225);
xnor U4293 (N_4293,N_3566,N_3700);
or U4294 (N_4294,N_2661,N_3364);
or U4295 (N_4295,N_3320,N_3717);
and U4296 (N_4296,N_3044,N_3048);
xnor U4297 (N_4297,N_2160,N_2524);
nand U4298 (N_4298,N_2235,N_2598);
nand U4299 (N_4299,N_2441,N_3344);
and U4300 (N_4300,N_2505,N_3739);
nor U4301 (N_4301,N_2848,N_3916);
xor U4302 (N_4302,N_2426,N_3031);
nor U4303 (N_4303,N_2258,N_2054);
xor U4304 (N_4304,N_2689,N_3167);
or U4305 (N_4305,N_2417,N_3784);
xnor U4306 (N_4306,N_3294,N_2518);
or U4307 (N_4307,N_3076,N_3418);
or U4308 (N_4308,N_3095,N_3756);
nand U4309 (N_4309,N_3801,N_3820);
nor U4310 (N_4310,N_2629,N_2902);
xnor U4311 (N_4311,N_3990,N_3059);
nand U4312 (N_4312,N_3945,N_2307);
nor U4313 (N_4313,N_2420,N_2337);
nor U4314 (N_4314,N_3703,N_3716);
xnor U4315 (N_4315,N_2352,N_3748);
and U4316 (N_4316,N_2719,N_2739);
nand U4317 (N_4317,N_2067,N_2338);
or U4318 (N_4318,N_3451,N_3150);
xor U4319 (N_4319,N_2156,N_3912);
xnor U4320 (N_4320,N_2591,N_2347);
or U4321 (N_4321,N_2253,N_3817);
nand U4322 (N_4322,N_3903,N_3952);
nand U4323 (N_4323,N_3785,N_3558);
or U4324 (N_4324,N_2775,N_3069);
nand U4325 (N_4325,N_3365,N_2799);
or U4326 (N_4326,N_2945,N_2584);
or U4327 (N_4327,N_2660,N_2424);
nor U4328 (N_4328,N_3589,N_3610);
or U4329 (N_4329,N_2216,N_2635);
nand U4330 (N_4330,N_2597,N_3084);
nor U4331 (N_4331,N_3316,N_3349);
nor U4332 (N_4332,N_2470,N_3603);
nand U4333 (N_4333,N_3041,N_3446);
or U4334 (N_4334,N_3857,N_2405);
xor U4335 (N_4335,N_3253,N_3908);
xnor U4336 (N_4336,N_3138,N_2027);
xor U4337 (N_4337,N_2460,N_3379);
nor U4338 (N_4338,N_2737,N_3449);
nor U4339 (N_4339,N_2297,N_3602);
nor U4340 (N_4340,N_2117,N_2708);
and U4341 (N_4341,N_3758,N_2101);
and U4342 (N_4342,N_2828,N_3314);
and U4343 (N_4343,N_3481,N_2178);
or U4344 (N_4344,N_3497,N_2636);
and U4345 (N_4345,N_3647,N_2138);
or U4346 (N_4346,N_3707,N_2557);
or U4347 (N_4347,N_2958,N_2977);
nand U4348 (N_4348,N_2289,N_3866);
nor U4349 (N_4349,N_3393,N_2649);
nand U4350 (N_4350,N_3023,N_2556);
nand U4351 (N_4351,N_3117,N_2877);
or U4352 (N_4352,N_2639,N_3855);
or U4353 (N_4353,N_2830,N_3265);
and U4354 (N_4354,N_3525,N_2750);
and U4355 (N_4355,N_3058,N_2644);
xor U4356 (N_4356,N_3254,N_3821);
xnor U4357 (N_4357,N_2327,N_3352);
xnor U4358 (N_4358,N_2064,N_3094);
nand U4359 (N_4359,N_3995,N_3104);
xnor U4360 (N_4360,N_3846,N_3456);
nor U4361 (N_4361,N_3242,N_3301);
xnor U4362 (N_4362,N_2621,N_2963);
and U4363 (N_4363,N_2249,N_2342);
nand U4364 (N_4364,N_3165,N_3689);
nand U4365 (N_4365,N_2548,N_3582);
or U4366 (N_4366,N_2068,N_3078);
nor U4367 (N_4367,N_2923,N_3822);
xor U4368 (N_4368,N_3455,N_2507);
xnor U4369 (N_4369,N_2919,N_2199);
nand U4370 (N_4370,N_3213,N_3311);
or U4371 (N_4371,N_2991,N_3782);
or U4372 (N_4372,N_3428,N_3092);
nor U4373 (N_4373,N_3371,N_3939);
nand U4374 (N_4374,N_3900,N_2443);
nand U4375 (N_4375,N_3452,N_3519);
xor U4376 (N_4376,N_2807,N_2318);
nor U4377 (N_4377,N_3630,N_2000);
nand U4378 (N_4378,N_3422,N_3627);
xor U4379 (N_4379,N_3460,N_3247);
or U4380 (N_4380,N_2130,N_2221);
nand U4381 (N_4381,N_3089,N_2103);
nor U4382 (N_4382,N_2335,N_3121);
nor U4383 (N_4383,N_3670,N_3273);
and U4384 (N_4384,N_3409,N_3520);
xnor U4385 (N_4385,N_2954,N_2254);
nor U4386 (N_4386,N_2533,N_3495);
or U4387 (N_4387,N_3386,N_2890);
nor U4388 (N_4388,N_3131,N_2604);
nand U4389 (N_4389,N_3985,N_3042);
or U4390 (N_4390,N_3767,N_3554);
xor U4391 (N_4391,N_3218,N_2893);
xor U4392 (N_4392,N_3642,N_3077);
nand U4393 (N_4393,N_3068,N_2432);
nor U4394 (N_4394,N_2964,N_3983);
nand U4395 (N_4395,N_3046,N_2600);
nor U4396 (N_4396,N_3750,N_2677);
and U4397 (N_4397,N_2204,N_2583);
or U4398 (N_4398,N_3523,N_3534);
xor U4399 (N_4399,N_2619,N_3168);
and U4400 (N_4400,N_3540,N_2921);
or U4401 (N_4401,N_2157,N_2733);
and U4402 (N_4402,N_2161,N_3129);
and U4403 (N_4403,N_3261,N_2251);
or U4404 (N_4404,N_3162,N_3141);
nor U4405 (N_4405,N_3274,N_2288);
or U4406 (N_4406,N_3547,N_3275);
xor U4407 (N_4407,N_2094,N_3223);
and U4408 (N_4408,N_3669,N_3696);
or U4409 (N_4409,N_2980,N_2994);
nand U4410 (N_4410,N_2390,N_2917);
nor U4411 (N_4411,N_2814,N_3656);
nand U4412 (N_4412,N_3148,N_2274);
or U4413 (N_4413,N_3477,N_2411);
xor U4414 (N_4414,N_3081,N_3672);
nand U4415 (N_4415,N_2479,N_3687);
xnor U4416 (N_4416,N_2153,N_2200);
xor U4417 (N_4417,N_3576,N_2602);
and U4418 (N_4418,N_3907,N_2916);
xor U4419 (N_4419,N_3932,N_3537);
xnor U4420 (N_4420,N_2606,N_3475);
or U4421 (N_4421,N_3580,N_2581);
nor U4422 (N_4422,N_3953,N_2028);
xor U4423 (N_4423,N_3524,N_3571);
xnor U4424 (N_4424,N_3969,N_3875);
nand U4425 (N_4425,N_3355,N_2961);
xnor U4426 (N_4426,N_3894,N_3000);
or U4427 (N_4427,N_2780,N_2687);
nand U4428 (N_4428,N_3324,N_2546);
and U4429 (N_4429,N_3489,N_3568);
xnor U4430 (N_4430,N_3544,N_3924);
and U4431 (N_4431,N_2093,N_3590);
xnor U4432 (N_4432,N_2433,N_3239);
or U4433 (N_4433,N_3638,N_2082);
xnor U4434 (N_4434,N_2304,N_3512);
xor U4435 (N_4435,N_3341,N_2099);
and U4436 (N_4436,N_3546,N_3329);
nor U4437 (N_4437,N_2947,N_2332);
or U4438 (N_4438,N_2174,N_3063);
xnor U4439 (N_4439,N_3780,N_3515);
nand U4440 (N_4440,N_3052,N_3202);
nor U4441 (N_4441,N_2882,N_2108);
nor U4442 (N_4442,N_2565,N_2495);
or U4443 (N_4443,N_2976,N_2077);
or U4444 (N_4444,N_2836,N_3877);
or U4445 (N_4445,N_3964,N_2676);
nor U4446 (N_4446,N_3443,N_2329);
and U4447 (N_4447,N_2609,N_3397);
and U4448 (N_4448,N_2025,N_3913);
and U4449 (N_4449,N_3978,N_3517);
nor U4450 (N_4450,N_2097,N_3302);
or U4451 (N_4451,N_3634,N_3779);
or U4452 (N_4452,N_3765,N_2709);
and U4453 (N_4453,N_2965,N_2616);
or U4454 (N_4454,N_2764,N_2368);
nor U4455 (N_4455,N_3557,N_2123);
nor U4456 (N_4456,N_2004,N_3003);
nor U4457 (N_4457,N_2264,N_3193);
and U4458 (N_4458,N_2220,N_3017);
or U4459 (N_4459,N_2162,N_3938);
nor U4460 (N_4460,N_3532,N_2996);
nand U4461 (N_4461,N_2754,N_3535);
xor U4462 (N_4462,N_2651,N_3102);
and U4463 (N_4463,N_3321,N_3257);
or U4464 (N_4464,N_2437,N_3387);
xnor U4465 (N_4465,N_3692,N_2459);
or U4466 (N_4466,N_3934,N_3013);
xor U4467 (N_4467,N_2769,N_2096);
nand U4468 (N_4468,N_2860,N_2984);
or U4469 (N_4469,N_3921,N_3066);
and U4470 (N_4470,N_2502,N_2478);
or U4471 (N_4471,N_3112,N_3946);
and U4472 (N_4472,N_3805,N_2485);
and U4473 (N_4473,N_3402,N_2494);
or U4474 (N_4474,N_3749,N_3262);
or U4475 (N_4475,N_3682,N_3550);
nor U4476 (N_4476,N_3230,N_2202);
nor U4477 (N_4477,N_3467,N_3710);
and U4478 (N_4478,N_2905,N_2438);
nor U4479 (N_4479,N_3731,N_3210);
nand U4480 (N_4480,N_3545,N_2826);
or U4481 (N_4481,N_3904,N_2053);
xnor U4482 (N_4482,N_2973,N_3322);
nand U4483 (N_4483,N_3139,N_2792);
nor U4484 (N_4484,N_2319,N_3800);
or U4485 (N_4485,N_3579,N_3468);
and U4486 (N_4486,N_3612,N_2501);
nor U4487 (N_4487,N_3640,N_2124);
nand U4488 (N_4488,N_3694,N_2186);
xor U4489 (N_4489,N_2510,N_3744);
nor U4490 (N_4490,N_3867,N_3458);
nand U4491 (N_4491,N_2915,N_3009);
nor U4492 (N_4492,N_3233,N_2658);
or U4493 (N_4493,N_3595,N_2005);
and U4494 (N_4494,N_2250,N_3114);
nand U4495 (N_4495,N_3197,N_2062);
nor U4496 (N_4496,N_2349,N_3030);
and U4497 (N_4497,N_3087,N_2392);
nor U4498 (N_4498,N_2021,N_3298);
nand U4499 (N_4499,N_3177,N_3679);
or U4500 (N_4500,N_3714,N_2167);
or U4501 (N_4501,N_3600,N_2759);
nor U4502 (N_4502,N_2177,N_2857);
xor U4503 (N_4503,N_3849,N_2768);
and U4504 (N_4504,N_2173,N_3258);
xor U4505 (N_4505,N_2026,N_2798);
xnor U4506 (N_4506,N_2457,N_3514);
xor U4507 (N_4507,N_3698,N_2942);
and U4508 (N_4508,N_2042,N_2552);
and U4509 (N_4509,N_2490,N_3407);
nor U4510 (N_4510,N_2458,N_3837);
xnor U4511 (N_4511,N_3173,N_2561);
nand U4512 (N_4512,N_2820,N_3415);
nor U4513 (N_4513,N_2573,N_3485);
nor U4514 (N_4514,N_2461,N_3623);
nor U4515 (N_4515,N_3593,N_2454);
or U4516 (N_4516,N_2653,N_3227);
nand U4517 (N_4517,N_2953,N_3241);
nand U4518 (N_4518,N_3429,N_2415);
or U4519 (N_4519,N_3308,N_3890);
nor U4520 (N_4520,N_2747,N_3563);
nand U4521 (N_4521,N_3854,N_3530);
nand U4522 (N_4522,N_2933,N_2985);
nor U4523 (N_4523,N_3657,N_3909);
xor U4524 (N_4524,N_3591,N_2643);
xor U4525 (N_4525,N_2397,N_2998);
nand U4526 (N_4526,N_3565,N_3843);
and U4527 (N_4527,N_2883,N_2894);
nor U4528 (N_4528,N_2686,N_3164);
nand U4529 (N_4529,N_2292,N_3337);
or U4530 (N_4530,N_3652,N_2228);
or U4531 (N_4531,N_3493,N_2935);
nand U4532 (N_4532,N_3369,N_3450);
xor U4533 (N_4533,N_2050,N_3174);
nor U4534 (N_4534,N_3769,N_2241);
nor U4535 (N_4535,N_2512,N_3248);
xnor U4536 (N_4536,N_2875,N_3772);
xor U4537 (N_4537,N_3113,N_3999);
or U4538 (N_4538,N_3291,N_2608);
or U4539 (N_4539,N_3297,N_2058);
nand U4540 (N_4540,N_3208,N_3835);
xnor U4541 (N_4541,N_3214,N_3615);
nand U4542 (N_4542,N_2126,N_2749);
nand U4543 (N_4543,N_3685,N_2316);
and U4544 (N_4544,N_2380,N_3606);
and U4545 (N_4545,N_3373,N_3122);
xor U4546 (N_4546,N_2574,N_3342);
and U4547 (N_4547,N_3156,N_2112);
or U4548 (N_4548,N_3228,N_2854);
nor U4549 (N_4549,N_2874,N_2949);
or U4550 (N_4550,N_2481,N_2044);
and U4551 (N_4551,N_2398,N_3295);
and U4552 (N_4552,N_2356,N_2110);
and U4553 (N_4553,N_3235,N_3878);
or U4554 (N_4554,N_2576,N_3016);
and U4555 (N_4555,N_2306,N_3594);
nor U4556 (N_4556,N_3354,N_3108);
xnor U4557 (N_4557,N_2703,N_2023);
nand U4558 (N_4558,N_2147,N_2146);
or U4559 (N_4559,N_3423,N_3336);
or U4560 (N_4560,N_2323,N_2230);
and U4561 (N_4561,N_3555,N_2838);
or U4562 (N_4562,N_2395,N_2165);
and U4563 (N_4563,N_2748,N_3636);
or U4564 (N_4564,N_3057,N_3868);
nor U4565 (N_4565,N_3778,N_2045);
nand U4566 (N_4566,N_3432,N_2321);
nand U4567 (N_4567,N_2477,N_2265);
and U4568 (N_4568,N_2981,N_3830);
xor U4569 (N_4569,N_2729,N_2314);
or U4570 (N_4570,N_3404,N_3622);
nand U4571 (N_4571,N_3333,N_3380);
nand U4572 (N_4572,N_3029,N_2466);
nand U4573 (N_4573,N_2351,N_3965);
nor U4574 (N_4574,N_3134,N_3893);
xnor U4575 (N_4575,N_2066,N_3348);
nor U4576 (N_4576,N_2074,N_2303);
and U4577 (N_4577,N_2983,N_3864);
and U4578 (N_4578,N_2757,N_2974);
or U4579 (N_4579,N_2791,N_2300);
and U4580 (N_4580,N_2776,N_2353);
xnor U4581 (N_4581,N_3653,N_3807);
xnor U4582 (N_4582,N_3277,N_2880);
nor U4583 (N_4583,N_2718,N_2884);
nor U4584 (N_4584,N_3439,N_2393);
and U4585 (N_4585,N_3116,N_2214);
nand U4586 (N_4586,N_2999,N_3433);
nand U4587 (N_4587,N_3201,N_2474);
or U4588 (N_4588,N_3706,N_3996);
nand U4589 (N_4589,N_3560,N_2593);
or U4590 (N_4590,N_2702,N_2154);
nor U4591 (N_4591,N_2758,N_2834);
and U4592 (N_4592,N_3979,N_3962);
and U4593 (N_4593,N_3219,N_3172);
or U4594 (N_4594,N_3673,N_2801);
nand U4595 (N_4595,N_3650,N_3447);
and U4596 (N_4596,N_3614,N_2070);
nand U4597 (N_4597,N_3408,N_3083);
nor U4598 (N_4598,N_2262,N_3915);
xor U4599 (N_4599,N_2149,N_3790);
nand U4600 (N_4600,N_2539,N_2847);
xnor U4601 (N_4601,N_2956,N_2497);
nand U4602 (N_4602,N_2637,N_2034);
and U4603 (N_4603,N_2735,N_2114);
nand U4604 (N_4604,N_2188,N_3768);
nand U4605 (N_4605,N_2272,N_2190);
xnor U4606 (N_4606,N_3305,N_2728);
xnor U4607 (N_4607,N_3181,N_2663);
and U4608 (N_4608,N_2813,N_2211);
xor U4609 (N_4609,N_3151,N_3984);
nand U4610 (N_4610,N_3431,N_3949);
and U4611 (N_4611,N_3578,N_3463);
nand U4612 (N_4612,N_2948,N_3973);
and U4613 (N_4613,N_2260,N_2560);
nor U4614 (N_4614,N_2069,N_2691);
and U4615 (N_4615,N_3526,N_3249);
nand U4616 (N_4616,N_2881,N_2374);
nand U4617 (N_4617,N_2504,N_3977);
nand U4618 (N_4618,N_3935,N_2853);
or U4619 (N_4619,N_2701,N_3863);
nand U4620 (N_4620,N_2090,N_3967);
and U4621 (N_4621,N_2704,N_2654);
xor U4622 (N_4622,N_2400,N_3741);
xor U4623 (N_4623,N_2903,N_2360);
nor U4624 (N_4624,N_2030,N_3661);
and U4625 (N_4625,N_3315,N_2878);
nand U4626 (N_4626,N_2059,N_2638);
or U4627 (N_4627,N_3766,N_2571);
or U4628 (N_4628,N_3147,N_3313);
nand U4629 (N_4629,N_3405,N_2142);
and U4630 (N_4630,N_2385,N_2282);
or U4631 (N_4631,N_3889,N_2169);
nand U4632 (N_4632,N_3632,N_3425);
nand U4633 (N_4633,N_2827,N_3221);
nor U4634 (N_4634,N_3549,N_3963);
nor U4635 (N_4635,N_2506,N_2731);
nand U4636 (N_4636,N_3876,N_2675);
and U4637 (N_4637,N_3851,N_3665);
nor U4638 (N_4638,N_2859,N_2139);
nand U4639 (N_4639,N_2952,N_3871);
xnor U4640 (N_4640,N_2646,N_3086);
nand U4641 (N_4641,N_3659,N_3263);
nand U4642 (N_4642,N_3690,N_3005);
xor U4643 (N_4643,N_3187,N_3154);
xnor U4644 (N_4644,N_3207,N_2404);
or U4645 (N_4645,N_3832,N_2445);
nand U4646 (N_4646,N_3170,N_3186);
or U4647 (N_4647,N_2127,N_3641);
xor U4648 (N_4648,N_2008,N_2081);
or U4649 (N_4649,N_2879,N_3733);
or U4650 (N_4650,N_2822,N_2195);
and U4651 (N_4651,N_2535,N_2369);
nand U4652 (N_4652,N_3572,N_2143);
or U4653 (N_4653,N_2080,N_2817);
and U4654 (N_4654,N_3861,N_2793);
nor U4655 (N_4655,N_3036,N_3891);
xor U4656 (N_4656,N_2447,N_3325);
and U4657 (N_4657,N_2038,N_2642);
nand U4658 (N_4658,N_3942,N_3874);
nand U4659 (N_4659,N_3968,N_2929);
nor U4660 (N_4660,N_2078,N_3677);
xor U4661 (N_4661,N_3658,N_3797);
xor U4662 (N_4662,N_2544,N_3663);
nand U4663 (N_4663,N_2795,N_2540);
or U4664 (N_4664,N_3307,N_2280);
or U4665 (N_4665,N_3802,N_2674);
and U4666 (N_4666,N_2449,N_2237);
xnor U4667 (N_4667,N_3808,N_3633);
or U4668 (N_4668,N_3869,N_3754);
xnor U4669 (N_4669,N_3586,N_2840);
or U4670 (N_4670,N_2547,N_3198);
nand U4671 (N_4671,N_3720,N_2802);
or U4672 (N_4672,N_2972,N_2232);
xor U4673 (N_4673,N_3794,N_2966);
nand U4674 (N_4674,N_2997,N_3505);
and U4675 (N_4675,N_2562,N_2960);
xor U4676 (N_4676,N_3222,N_2233);
nor U4677 (N_4677,N_3601,N_2407);
nor U4678 (N_4678,N_2091,N_3944);
nand U4679 (N_4679,N_2326,N_2084);
or U4680 (N_4680,N_2711,N_3276);
or U4681 (N_4681,N_2525,N_3947);
and U4682 (N_4682,N_2464,N_3303);
xor U4683 (N_4683,N_2294,N_2615);
and U4684 (N_4684,N_2519,N_3529);
or U4685 (N_4685,N_3734,N_3127);
nor U4686 (N_4686,N_3541,N_3511);
nand U4687 (N_4687,N_2950,N_3742);
and U4688 (N_4688,N_3500,N_3556);
and U4689 (N_4689,N_2248,N_3318);
nand U4690 (N_4690,N_2362,N_3751);
or U4691 (N_4691,N_2819,N_2498);
xor U4692 (N_4692,N_3070,N_2134);
and U4693 (N_4693,N_2375,N_2083);
and U4694 (N_4694,N_2987,N_2752);
xnor U4695 (N_4695,N_2913,N_2959);
and U4696 (N_4696,N_2252,N_3613);
and U4697 (N_4697,N_3424,N_3246);
nor U4698 (N_4698,N_2683,N_3435);
nand U4699 (N_4699,N_2071,N_3200);
xnor U4700 (N_4700,N_3142,N_2348);
nand U4701 (N_4701,N_2346,N_3611);
nand U4702 (N_4702,N_3704,N_3035);
xnor U4703 (N_4703,N_3956,N_2527);
and U4704 (N_4704,N_3188,N_3809);
and U4705 (N_4705,N_2423,N_2968);
nand U4706 (N_4706,N_2610,N_2471);
nor U4707 (N_4707,N_3738,N_2336);
nand U4708 (N_4708,N_2017,N_2104);
and U4709 (N_4709,N_3553,N_3237);
xnor U4710 (N_4710,N_2868,N_2182);
and U4711 (N_4711,N_3527,N_3899);
and U4712 (N_4712,N_2647,N_2164);
and U4713 (N_4713,N_2185,N_3926);
nor U4714 (N_4714,N_3143,N_2624);
nand U4715 (N_4715,N_3693,N_3608);
nor U4716 (N_4716,N_3814,N_3445);
and U4717 (N_4717,N_2550,N_2992);
or U4718 (N_4718,N_3251,N_2313);
nand U4719 (N_4719,N_2969,N_3278);
or U4720 (N_4720,N_2569,N_3326);
or U4721 (N_4721,N_3002,N_3588);
xor U4722 (N_4722,N_2622,N_2720);
nand U4723 (N_4723,N_2267,N_2456);
or U4724 (N_4724,N_2378,N_2967);
xnor U4725 (N_4725,N_3856,N_3250);
nand U4726 (N_4726,N_3413,N_3293);
nor U4727 (N_4727,N_2035,N_2970);
nor U4728 (N_4728,N_2037,N_3775);
xnor U4729 (N_4729,N_2446,N_3178);
and U4730 (N_4730,N_3597,N_2151);
xor U4731 (N_4731,N_2796,N_2118);
and U4732 (N_4732,N_2715,N_3280);
and U4733 (N_4733,N_2076,N_2476);
xnor U4734 (N_4734,N_2694,N_2148);
nand U4735 (N_4735,N_2085,N_3372);
xor U4736 (N_4736,N_2133,N_3358);
xor U4737 (N_4737,N_3646,N_2620);
and U4738 (N_4738,N_3486,N_2209);
xnor U4739 (N_4739,N_3478,N_2736);
nor U4740 (N_4740,N_3732,N_3361);
and U4741 (N_4741,N_3791,N_2060);
and U4742 (N_4742,N_2367,N_3001);
and U4743 (N_4743,N_2867,N_2381);
and U4744 (N_4744,N_2416,N_2015);
nor U4745 (N_4745,N_3847,N_3140);
nor U4746 (N_4746,N_2725,N_2783);
nor U4747 (N_4747,N_3862,N_2191);
or U4748 (N_4748,N_3922,N_3577);
or U4749 (N_4749,N_3238,N_2275);
or U4750 (N_4750,N_2238,N_2724);
xor U4751 (N_4751,N_3287,N_2773);
or U4752 (N_4752,N_3345,N_3159);
and U4753 (N_4753,N_3304,N_3145);
nor U4754 (N_4754,N_3604,N_2227);
nand U4755 (N_4755,N_2463,N_2361);
xor U4756 (N_4756,N_3149,N_3872);
xnor U4757 (N_4757,N_2839,N_2333);
or U4758 (N_4758,N_3378,N_3993);
or U4759 (N_4759,N_2782,N_3331);
xnor U4760 (N_4760,N_2383,N_3229);
nand U4761 (N_4761,N_2016,N_2681);
xnor U4762 (N_4762,N_3146,N_2107);
xor U4763 (N_4763,N_2978,N_3400);
xor U4764 (N_4764,N_3299,N_2086);
and U4765 (N_4765,N_3204,N_2256);
and U4766 (N_4766,N_2900,N_3533);
nand U4767 (N_4767,N_3353,N_2580);
and U4768 (N_4768,N_3359,N_3625);
or U4769 (N_4769,N_2386,N_2339);
or U4770 (N_4770,N_3231,N_3025);
nor U4771 (N_4771,N_3360,N_3323);
nor U4772 (N_4772,N_2179,N_2613);
nand U4773 (N_4773,N_2697,N_3564);
nand U4774 (N_4774,N_2039,N_3389);
nor U4775 (N_4775,N_3718,N_3490);
or U4776 (N_4776,N_2809,N_3989);
or U4777 (N_4777,N_2222,N_3715);
xnor U4778 (N_4778,N_3997,N_3296);
nand U4779 (N_4779,N_3270,N_2373);
xnor U4780 (N_4780,N_3007,N_3655);
nor U4781 (N_4781,N_2626,N_3954);
or U4782 (N_4782,N_2242,N_3770);
and U4783 (N_4783,N_3008,N_3406);
nand U4784 (N_4784,N_2239,N_2870);
nand U4785 (N_4785,N_2937,N_2197);
and U4786 (N_4786,N_3881,N_2279);
nor U4787 (N_4787,N_3948,N_2277);
or U4788 (N_4788,N_2886,N_2111);
and U4789 (N_4789,N_3902,N_2601);
xor U4790 (N_4790,N_2043,N_2295);
xnor U4791 (N_4791,N_2287,N_2761);
nand U4792 (N_4792,N_2489,N_3911);
and U4793 (N_4793,N_2168,N_2468);
xnor U4794 (N_4794,N_2567,N_3961);
and U4795 (N_4795,N_3053,N_3898);
nor U4796 (N_4796,N_2727,N_2422);
xor U4797 (N_4797,N_2180,N_3930);
or U4798 (N_4798,N_3021,N_2931);
or U4799 (N_4799,N_2932,N_2656);
or U4800 (N_4800,N_3232,N_2229);
nand U4801 (N_4801,N_3082,N_2487);
and U4802 (N_4802,N_2549,N_3469);
nand U4803 (N_4803,N_3022,N_3444);
xnor U4804 (N_4804,N_2418,N_2150);
nand U4805 (N_4805,N_2818,N_2377);
and U4806 (N_4806,N_3268,N_2751);
or U4807 (N_4807,N_2278,N_3437);
nor U4808 (N_4808,N_3043,N_3370);
and U4809 (N_4809,N_2051,N_2472);
xnor U4810 (N_4810,N_3786,N_3100);
nand U4811 (N_4811,N_2911,N_3981);
and U4812 (N_4812,N_3551,N_3959);
and U4813 (N_4813,N_2308,N_2800);
nand U4814 (N_4814,N_2652,N_3096);
nand U4815 (N_4815,N_3088,N_3970);
nand U4816 (N_4816,N_3776,N_3306);
or U4817 (N_4817,N_3950,N_3171);
and U4818 (N_4818,N_3631,N_3414);
nor U4819 (N_4819,N_3747,N_3870);
and U4820 (N_4820,N_3574,N_2427);
or U4821 (N_4821,N_2941,N_3438);
nor U4822 (N_4822,N_2401,N_3166);
nand U4823 (N_4823,N_3085,N_2328);
nand U4824 (N_4824,N_2924,N_3271);
and U4825 (N_4825,N_3226,N_3680);
nand U4826 (N_4826,N_2181,N_2428);
xnor U4827 (N_4827,N_2056,N_2344);
nor U4828 (N_4828,N_3504,N_3567);
nor U4829 (N_4829,N_2020,N_2440);
and U4830 (N_4830,N_3195,N_3773);
and U4831 (N_4831,N_3010,N_2409);
or U4832 (N_4832,N_2869,N_3887);
nand U4833 (N_4833,N_2927,N_2664);
and U4834 (N_4834,N_2543,N_3416);
nand U4835 (N_4835,N_3090,N_3688);
nand U4836 (N_4836,N_3220,N_2767);
nor U4837 (N_4837,N_3736,N_2125);
or U4838 (N_4838,N_2517,N_2379);
nor U4839 (N_4839,N_2618,N_3513);
nor U4840 (N_4840,N_2135,N_3382);
nor U4841 (N_4841,N_2698,N_2957);
and U4842 (N_4842,N_3998,N_3781);
or U4843 (N_4843,N_3144,N_3124);
xnor U4844 (N_4844,N_2217,N_3831);
or U4845 (N_4845,N_3080,N_2899);
xor U4846 (N_4846,N_2808,N_3829);
and U4847 (N_4847,N_3269,N_3503);
xnor U4848 (N_4848,N_2712,N_3971);
or U4849 (N_4849,N_3256,N_2741);
xor U4850 (N_4850,N_3260,N_3328);
nand U4851 (N_4851,N_2310,N_2585);
nor U4852 (N_4852,N_3465,N_2414);
nor U4853 (N_4853,N_2526,N_2760);
nand U4854 (N_4854,N_2419,N_3873);
nor U4855 (N_4855,N_3569,N_2993);
nor U4856 (N_4856,N_2595,N_2700);
or U4857 (N_4857,N_2672,N_2003);
nand U4858 (N_4858,N_3136,N_3441);
nor U4859 (N_4859,N_3804,N_2106);
nand U4860 (N_4860,N_2770,N_2382);
and U4861 (N_4861,N_3957,N_2136);
or U4862 (N_4862,N_2500,N_3936);
nand U4863 (N_4863,N_3019,N_2633);
nand U4864 (N_4864,N_3347,N_3721);
xor U4865 (N_4865,N_2102,N_3709);
and U4866 (N_4866,N_2137,N_2341);
or U4867 (N_4867,N_2129,N_3927);
or U4868 (N_4868,N_3836,N_2171);
nand U4869 (N_4869,N_2763,N_2283);
and U4870 (N_4870,N_2089,N_2320);
nor U4871 (N_4871,N_3509,N_2841);
xor U4872 (N_4872,N_3826,N_3396);
nand U4873 (N_4873,N_2797,N_2002);
or U4874 (N_4874,N_2408,N_3011);
and U4875 (N_4875,N_2269,N_3309);
nor U4876 (N_4876,N_2467,N_3398);
nand U4877 (N_4877,N_3994,N_3440);
xnor U4878 (N_4878,N_2144,N_2145);
nor U4879 (N_4879,N_2673,N_3777);
or U4880 (N_4880,N_3191,N_2623);
or U4881 (N_4881,N_3098,N_2832);
nand U4882 (N_4882,N_2046,N_2804);
nand U4883 (N_4883,N_3722,N_3062);
nand U4884 (N_4884,N_2530,N_2350);
nand U4885 (N_4885,N_2024,N_2784);
and U4886 (N_4886,N_2244,N_2564);
nand U4887 (N_4887,N_2215,N_3618);
nand U4888 (N_4888,N_3161,N_2559);
nand U4889 (N_4889,N_3883,N_3757);
and U4890 (N_4890,N_2245,N_2120);
nor U4891 (N_4891,N_3033,N_3848);
nor U4892 (N_4892,N_3931,N_2152);
or U4893 (N_4893,N_2887,N_2898);
nor U4894 (N_4894,N_3884,N_3004);
nor U4895 (N_4895,N_3381,N_2198);
xnor U4896 (N_4896,N_3906,N_3783);
and U4897 (N_4897,N_2665,N_3051);
nand U4898 (N_4898,N_2553,N_3937);
and U4899 (N_4899,N_3417,N_3882);
xnor U4900 (N_4900,N_3244,N_2366);
and U4901 (N_4901,N_2888,N_3319);
xnor U4902 (N_4902,N_2011,N_2194);
nor U4903 (N_4903,N_2047,N_3103);
nand U4904 (N_4904,N_2962,N_3434);
nor U4905 (N_4905,N_3179,N_2955);
or U4906 (N_4906,N_2690,N_2846);
xor U4907 (N_4907,N_2975,N_2014);
nor U4908 (N_4908,N_3283,N_2431);
nand U4909 (N_4909,N_2995,N_3152);
or U4910 (N_4910,N_3584,N_3464);
or U4911 (N_4911,N_3494,N_2399);
nor U4912 (N_4912,N_2480,N_2012);
and U4913 (N_4913,N_2938,N_2018);
and U4914 (N_4914,N_2896,N_2121);
and U4915 (N_4915,N_3390,N_3755);
and U4916 (N_4916,N_3743,N_3091);
nand U4917 (N_4917,N_3697,N_2920);
nand U4918 (N_4918,N_2590,N_3476);
and U4919 (N_4919,N_2578,N_2829);
and U4920 (N_4920,N_2098,N_2918);
nand U4921 (N_4921,N_2293,N_2263);
and U4922 (N_4922,N_2273,N_3176);
nor U4923 (N_4923,N_2219,N_2218);
or U4924 (N_4924,N_2781,N_2716);
or U4925 (N_4925,N_2315,N_2914);
xnor U4926 (N_4926,N_2542,N_2680);
and U4927 (N_4927,N_2009,N_2048);
and U4928 (N_4928,N_3816,N_3061);
or U4929 (N_4929,N_2452,N_3824);
xor U4930 (N_4930,N_2669,N_3958);
or U4931 (N_4931,N_3101,N_2403);
nor U4932 (N_4932,N_2285,N_2605);
and U4933 (N_4933,N_3701,N_3383);
or U4934 (N_4934,N_2907,N_2726);
or U4935 (N_4935,N_3442,N_2109);
nor U4936 (N_4936,N_2534,N_2063);
nor U4937 (N_4937,N_3267,N_3462);
nand U4938 (N_4938,N_3472,N_3746);
nor U4939 (N_4939,N_3825,N_3488);
or U4940 (N_4940,N_2939,N_2483);
nor U4941 (N_4941,N_3028,N_3925);
nand U4942 (N_4942,N_3845,N_2930);
nor U4943 (N_4943,N_2073,N_2301);
and U4944 (N_4944,N_3175,N_3106);
nand U4945 (N_4945,N_2049,N_2119);
nand U4946 (N_4946,N_3859,N_2657);
nor U4947 (N_4947,N_2815,N_3919);
or U4948 (N_4948,N_3598,N_2566);
or U4949 (N_4949,N_2391,N_3346);
and U4950 (N_4950,N_2243,N_3480);
xor U4951 (N_4951,N_3203,N_3759);
or U4952 (N_4952,N_2908,N_2075);
nor U4953 (N_4953,N_2906,N_3027);
nand U4954 (N_4954,N_2684,N_3427);
xor U4955 (N_4955,N_2493,N_2771);
nor U4956 (N_4956,N_3668,N_2363);
xnor U4957 (N_4957,N_2116,N_2612);
nor U4958 (N_4958,N_3885,N_3982);
or U4959 (N_4959,N_3619,N_2388);
xor U4960 (N_4960,N_3420,N_2354);
nand U4961 (N_4961,N_3723,N_2789);
or U4962 (N_4962,N_2579,N_2895);
or U4963 (N_4963,N_2596,N_2515);
and U4964 (N_4964,N_2988,N_2928);
nand U4965 (N_4965,N_2276,N_3654);
xor U4966 (N_4966,N_2299,N_3123);
xnor U4967 (N_4967,N_2473,N_2873);
nor U4968 (N_4968,N_2413,N_3205);
nor U4969 (N_4969,N_3839,N_2345);
and U4970 (N_4970,N_3037,N_2389);
and U4971 (N_4971,N_3255,N_2531);
nor U4972 (N_4972,N_2492,N_2436);
and U4973 (N_4973,N_3853,N_3157);
xnor U4974 (N_4974,N_2036,N_3483);
nor U4975 (N_4975,N_3695,N_3281);
or U4976 (N_4976,N_2298,N_2384);
xor U4977 (N_4977,N_3498,N_2033);
xor U4978 (N_4978,N_2100,N_3163);
xor U4979 (N_4979,N_2131,N_2010);
nand U4980 (N_4980,N_2007,N_3649);
xnor U4981 (N_4981,N_3752,N_3901);
nor U4982 (N_4982,N_2402,N_3955);
or U4983 (N_4983,N_3310,N_2175);
xor U4984 (N_4984,N_3726,N_2448);
nor U4985 (N_4985,N_2645,N_2439);
and U4986 (N_4986,N_3079,N_2442);
nand U4987 (N_4987,N_2031,N_2541);
nand U4988 (N_4988,N_2234,N_3575);
nor U4989 (N_4989,N_3473,N_2122);
or U4990 (N_4990,N_2592,N_3986);
nand U4991 (N_4991,N_3745,N_2765);
nand U4992 (N_4992,N_3111,N_3351);
xnor U4993 (N_4993,N_2936,N_2554);
xor U4994 (N_4994,N_3528,N_3097);
xor U4995 (N_4995,N_3338,N_3667);
or U4996 (N_4996,N_3192,N_3403);
nand U4997 (N_4997,N_2614,N_3516);
nand U4998 (N_4998,N_2670,N_2844);
xor U4999 (N_4999,N_3727,N_2072);
nor U5000 (N_5000,N_3192,N_2350);
or U5001 (N_5001,N_3491,N_2182);
or U5002 (N_5002,N_2941,N_2758);
xnor U5003 (N_5003,N_3647,N_3203);
xor U5004 (N_5004,N_3868,N_2566);
and U5005 (N_5005,N_2124,N_3476);
xnor U5006 (N_5006,N_2092,N_3094);
and U5007 (N_5007,N_3373,N_2468);
or U5008 (N_5008,N_2089,N_3016);
xnor U5009 (N_5009,N_3585,N_3063);
xor U5010 (N_5010,N_2495,N_2924);
and U5011 (N_5011,N_3154,N_3804);
nand U5012 (N_5012,N_3914,N_3556);
and U5013 (N_5013,N_2650,N_3396);
nor U5014 (N_5014,N_3137,N_2876);
or U5015 (N_5015,N_3155,N_3163);
or U5016 (N_5016,N_2996,N_2106);
and U5017 (N_5017,N_2018,N_2788);
or U5018 (N_5018,N_3429,N_3205);
nand U5019 (N_5019,N_2390,N_2084);
or U5020 (N_5020,N_3508,N_2337);
or U5021 (N_5021,N_3708,N_3003);
nand U5022 (N_5022,N_3476,N_3503);
nor U5023 (N_5023,N_3283,N_3318);
and U5024 (N_5024,N_2972,N_3952);
nand U5025 (N_5025,N_3009,N_2363);
or U5026 (N_5026,N_3639,N_2507);
xor U5027 (N_5027,N_2872,N_2898);
and U5028 (N_5028,N_3317,N_2663);
nor U5029 (N_5029,N_3372,N_2923);
and U5030 (N_5030,N_2902,N_3245);
xnor U5031 (N_5031,N_2185,N_2609);
nor U5032 (N_5032,N_2377,N_3478);
and U5033 (N_5033,N_3483,N_2002);
nor U5034 (N_5034,N_3915,N_2201);
nor U5035 (N_5035,N_3842,N_3371);
or U5036 (N_5036,N_3798,N_2118);
or U5037 (N_5037,N_3240,N_2318);
or U5038 (N_5038,N_2906,N_2456);
and U5039 (N_5039,N_3344,N_2734);
xor U5040 (N_5040,N_2034,N_2123);
nand U5041 (N_5041,N_2522,N_2850);
or U5042 (N_5042,N_3722,N_2304);
nand U5043 (N_5043,N_2422,N_2777);
xor U5044 (N_5044,N_2405,N_2763);
nand U5045 (N_5045,N_3261,N_2094);
and U5046 (N_5046,N_2555,N_2188);
nand U5047 (N_5047,N_2004,N_2140);
nor U5048 (N_5048,N_2998,N_2253);
nand U5049 (N_5049,N_3173,N_2777);
or U5050 (N_5050,N_2974,N_3392);
nand U5051 (N_5051,N_2353,N_3491);
xnor U5052 (N_5052,N_3007,N_3287);
xnor U5053 (N_5053,N_2043,N_2217);
xnor U5054 (N_5054,N_2571,N_2681);
or U5055 (N_5055,N_3887,N_2257);
and U5056 (N_5056,N_3837,N_3453);
or U5057 (N_5057,N_2542,N_3177);
nor U5058 (N_5058,N_2658,N_3505);
nor U5059 (N_5059,N_3667,N_3827);
xnor U5060 (N_5060,N_3524,N_3869);
nand U5061 (N_5061,N_2991,N_2748);
xor U5062 (N_5062,N_3664,N_3027);
nor U5063 (N_5063,N_2392,N_3202);
nor U5064 (N_5064,N_2154,N_2499);
or U5065 (N_5065,N_2708,N_2222);
nand U5066 (N_5066,N_2623,N_2333);
and U5067 (N_5067,N_2852,N_2332);
and U5068 (N_5068,N_2999,N_2023);
xnor U5069 (N_5069,N_2676,N_2996);
nor U5070 (N_5070,N_3589,N_3498);
nor U5071 (N_5071,N_2143,N_2914);
xor U5072 (N_5072,N_2490,N_2597);
xnor U5073 (N_5073,N_2027,N_2952);
and U5074 (N_5074,N_2077,N_3589);
nor U5075 (N_5075,N_3448,N_3711);
nor U5076 (N_5076,N_3115,N_3855);
xnor U5077 (N_5077,N_3818,N_2352);
nor U5078 (N_5078,N_3175,N_3522);
and U5079 (N_5079,N_3848,N_2753);
nand U5080 (N_5080,N_2084,N_2293);
and U5081 (N_5081,N_2170,N_2430);
and U5082 (N_5082,N_3971,N_2182);
and U5083 (N_5083,N_3495,N_3009);
nor U5084 (N_5084,N_2108,N_3267);
nor U5085 (N_5085,N_3769,N_2437);
nand U5086 (N_5086,N_2790,N_3968);
nand U5087 (N_5087,N_3780,N_2944);
nor U5088 (N_5088,N_2071,N_3647);
or U5089 (N_5089,N_2536,N_2921);
nor U5090 (N_5090,N_2167,N_3378);
and U5091 (N_5091,N_2850,N_2453);
nand U5092 (N_5092,N_2104,N_3651);
nand U5093 (N_5093,N_3514,N_3004);
or U5094 (N_5094,N_2864,N_3211);
nor U5095 (N_5095,N_3226,N_2383);
nand U5096 (N_5096,N_3962,N_2756);
nor U5097 (N_5097,N_2179,N_2534);
xor U5098 (N_5098,N_2338,N_2073);
nand U5099 (N_5099,N_3413,N_3861);
nand U5100 (N_5100,N_2710,N_2436);
or U5101 (N_5101,N_3908,N_3652);
nand U5102 (N_5102,N_3580,N_2799);
nand U5103 (N_5103,N_2519,N_3282);
nor U5104 (N_5104,N_2375,N_3677);
nand U5105 (N_5105,N_3906,N_2183);
nor U5106 (N_5106,N_2376,N_3403);
nor U5107 (N_5107,N_3459,N_3265);
and U5108 (N_5108,N_3827,N_2751);
nor U5109 (N_5109,N_3508,N_3170);
xnor U5110 (N_5110,N_3973,N_2697);
and U5111 (N_5111,N_3178,N_2314);
or U5112 (N_5112,N_2599,N_3285);
nand U5113 (N_5113,N_3746,N_2479);
xor U5114 (N_5114,N_3631,N_2010);
or U5115 (N_5115,N_3986,N_3668);
and U5116 (N_5116,N_3220,N_3982);
xnor U5117 (N_5117,N_3422,N_3348);
nor U5118 (N_5118,N_2822,N_3875);
and U5119 (N_5119,N_2674,N_2492);
nor U5120 (N_5120,N_3474,N_3948);
nand U5121 (N_5121,N_2315,N_3752);
or U5122 (N_5122,N_3936,N_3915);
nand U5123 (N_5123,N_3626,N_2869);
nand U5124 (N_5124,N_2845,N_2079);
nand U5125 (N_5125,N_3056,N_3986);
xor U5126 (N_5126,N_3130,N_3413);
xnor U5127 (N_5127,N_2762,N_3499);
nor U5128 (N_5128,N_2432,N_2964);
or U5129 (N_5129,N_2607,N_3905);
or U5130 (N_5130,N_3440,N_2900);
nor U5131 (N_5131,N_2605,N_2003);
or U5132 (N_5132,N_3593,N_3617);
nand U5133 (N_5133,N_2329,N_3268);
xnor U5134 (N_5134,N_2742,N_3079);
xor U5135 (N_5135,N_2291,N_2957);
or U5136 (N_5136,N_2704,N_3239);
nand U5137 (N_5137,N_3020,N_3681);
nor U5138 (N_5138,N_2679,N_3843);
nand U5139 (N_5139,N_3420,N_3671);
or U5140 (N_5140,N_3209,N_2822);
and U5141 (N_5141,N_3495,N_2343);
nor U5142 (N_5142,N_3117,N_3440);
and U5143 (N_5143,N_2518,N_3333);
xor U5144 (N_5144,N_2309,N_2536);
xor U5145 (N_5145,N_2180,N_3842);
xor U5146 (N_5146,N_3118,N_2151);
nor U5147 (N_5147,N_2603,N_2856);
xnor U5148 (N_5148,N_2347,N_2047);
nor U5149 (N_5149,N_2943,N_3955);
or U5150 (N_5150,N_2358,N_3597);
nor U5151 (N_5151,N_2827,N_2182);
nor U5152 (N_5152,N_3302,N_2807);
xor U5153 (N_5153,N_3885,N_3380);
or U5154 (N_5154,N_2280,N_2736);
and U5155 (N_5155,N_3191,N_2287);
nor U5156 (N_5156,N_3559,N_2349);
nand U5157 (N_5157,N_3884,N_2733);
nand U5158 (N_5158,N_2044,N_2372);
xor U5159 (N_5159,N_2868,N_3406);
xnor U5160 (N_5160,N_2751,N_3081);
and U5161 (N_5161,N_3891,N_3619);
nand U5162 (N_5162,N_2702,N_3045);
nand U5163 (N_5163,N_3392,N_3562);
nand U5164 (N_5164,N_3559,N_3407);
and U5165 (N_5165,N_3111,N_3006);
nor U5166 (N_5166,N_2390,N_3289);
nand U5167 (N_5167,N_3448,N_2899);
nand U5168 (N_5168,N_2167,N_2322);
nor U5169 (N_5169,N_2484,N_3402);
nand U5170 (N_5170,N_3207,N_3784);
xor U5171 (N_5171,N_2779,N_3547);
xnor U5172 (N_5172,N_2532,N_2466);
nand U5173 (N_5173,N_3633,N_2154);
nand U5174 (N_5174,N_3814,N_2713);
xor U5175 (N_5175,N_3516,N_2766);
nor U5176 (N_5176,N_3307,N_2966);
or U5177 (N_5177,N_2292,N_2444);
and U5178 (N_5178,N_2107,N_3795);
nand U5179 (N_5179,N_3498,N_3378);
nor U5180 (N_5180,N_3782,N_3956);
xnor U5181 (N_5181,N_2853,N_2367);
nand U5182 (N_5182,N_3288,N_2663);
xor U5183 (N_5183,N_2686,N_3876);
nor U5184 (N_5184,N_2724,N_2581);
nand U5185 (N_5185,N_3176,N_3108);
or U5186 (N_5186,N_2286,N_2489);
and U5187 (N_5187,N_3560,N_3020);
xnor U5188 (N_5188,N_3028,N_2661);
or U5189 (N_5189,N_3211,N_2842);
nand U5190 (N_5190,N_2950,N_2361);
and U5191 (N_5191,N_3800,N_2767);
xor U5192 (N_5192,N_2322,N_2546);
nand U5193 (N_5193,N_3367,N_3956);
and U5194 (N_5194,N_3657,N_3287);
or U5195 (N_5195,N_2124,N_2912);
nor U5196 (N_5196,N_3027,N_3022);
nor U5197 (N_5197,N_3144,N_3454);
nand U5198 (N_5198,N_2962,N_3831);
and U5199 (N_5199,N_2832,N_3062);
nand U5200 (N_5200,N_3422,N_3439);
and U5201 (N_5201,N_3020,N_2368);
xor U5202 (N_5202,N_3844,N_3913);
and U5203 (N_5203,N_3537,N_2913);
nor U5204 (N_5204,N_3076,N_3541);
xnor U5205 (N_5205,N_3918,N_3492);
nand U5206 (N_5206,N_2292,N_2367);
nor U5207 (N_5207,N_3761,N_2554);
and U5208 (N_5208,N_3647,N_3992);
xnor U5209 (N_5209,N_3253,N_3033);
or U5210 (N_5210,N_3249,N_3375);
and U5211 (N_5211,N_3826,N_2173);
and U5212 (N_5212,N_2835,N_3026);
nor U5213 (N_5213,N_3396,N_3120);
nor U5214 (N_5214,N_2238,N_3536);
nand U5215 (N_5215,N_3261,N_2757);
or U5216 (N_5216,N_2480,N_3518);
nor U5217 (N_5217,N_2198,N_3249);
or U5218 (N_5218,N_3197,N_2454);
and U5219 (N_5219,N_2180,N_2856);
or U5220 (N_5220,N_2261,N_3603);
or U5221 (N_5221,N_3969,N_3527);
and U5222 (N_5222,N_3048,N_3779);
and U5223 (N_5223,N_2926,N_2944);
and U5224 (N_5224,N_3074,N_3837);
or U5225 (N_5225,N_3108,N_3140);
xnor U5226 (N_5226,N_3261,N_3402);
xor U5227 (N_5227,N_3301,N_2529);
xor U5228 (N_5228,N_2668,N_3270);
or U5229 (N_5229,N_2152,N_2157);
nand U5230 (N_5230,N_3510,N_2423);
nand U5231 (N_5231,N_2400,N_2335);
nor U5232 (N_5232,N_2404,N_3766);
nor U5233 (N_5233,N_2094,N_3877);
xnor U5234 (N_5234,N_3481,N_2873);
nor U5235 (N_5235,N_3612,N_3354);
nand U5236 (N_5236,N_3159,N_2330);
nand U5237 (N_5237,N_3469,N_2424);
nor U5238 (N_5238,N_2856,N_2298);
and U5239 (N_5239,N_3227,N_3179);
xor U5240 (N_5240,N_3234,N_3648);
and U5241 (N_5241,N_3464,N_2282);
and U5242 (N_5242,N_2863,N_3875);
xor U5243 (N_5243,N_3458,N_2982);
nor U5244 (N_5244,N_3257,N_2968);
or U5245 (N_5245,N_2468,N_3363);
and U5246 (N_5246,N_3326,N_2405);
nand U5247 (N_5247,N_2205,N_2122);
xor U5248 (N_5248,N_3589,N_2095);
or U5249 (N_5249,N_2374,N_2166);
nand U5250 (N_5250,N_2196,N_2112);
and U5251 (N_5251,N_2535,N_2063);
and U5252 (N_5252,N_2408,N_2692);
xor U5253 (N_5253,N_3274,N_2469);
nor U5254 (N_5254,N_3211,N_3378);
nand U5255 (N_5255,N_2468,N_2885);
xor U5256 (N_5256,N_2973,N_3531);
and U5257 (N_5257,N_2327,N_3821);
or U5258 (N_5258,N_3300,N_2481);
nor U5259 (N_5259,N_2826,N_2865);
nand U5260 (N_5260,N_3325,N_3934);
nor U5261 (N_5261,N_2346,N_3152);
xor U5262 (N_5262,N_3636,N_3318);
and U5263 (N_5263,N_3290,N_3619);
xor U5264 (N_5264,N_3970,N_3351);
and U5265 (N_5265,N_2666,N_2983);
and U5266 (N_5266,N_3705,N_3435);
and U5267 (N_5267,N_3356,N_2194);
nand U5268 (N_5268,N_3190,N_3543);
nand U5269 (N_5269,N_3137,N_3618);
nand U5270 (N_5270,N_2462,N_3825);
xnor U5271 (N_5271,N_2972,N_2997);
or U5272 (N_5272,N_3916,N_2645);
nor U5273 (N_5273,N_2907,N_2903);
xor U5274 (N_5274,N_2034,N_2745);
nand U5275 (N_5275,N_2033,N_3026);
and U5276 (N_5276,N_2655,N_2424);
nand U5277 (N_5277,N_2264,N_3614);
xor U5278 (N_5278,N_3075,N_3971);
nor U5279 (N_5279,N_2852,N_3386);
nor U5280 (N_5280,N_2760,N_3013);
xnor U5281 (N_5281,N_2680,N_3762);
nand U5282 (N_5282,N_2928,N_3756);
and U5283 (N_5283,N_3706,N_3703);
xor U5284 (N_5284,N_3664,N_2303);
and U5285 (N_5285,N_2802,N_3648);
and U5286 (N_5286,N_2200,N_3390);
nor U5287 (N_5287,N_2824,N_2555);
xor U5288 (N_5288,N_3169,N_3623);
and U5289 (N_5289,N_2337,N_2300);
xnor U5290 (N_5290,N_2843,N_3454);
nor U5291 (N_5291,N_3711,N_3600);
nand U5292 (N_5292,N_2559,N_2252);
and U5293 (N_5293,N_3309,N_2828);
nor U5294 (N_5294,N_2198,N_2977);
or U5295 (N_5295,N_2604,N_2042);
xor U5296 (N_5296,N_3939,N_2383);
xnor U5297 (N_5297,N_3888,N_2334);
xnor U5298 (N_5298,N_3368,N_2117);
and U5299 (N_5299,N_3749,N_3540);
or U5300 (N_5300,N_2599,N_3919);
or U5301 (N_5301,N_2901,N_3101);
and U5302 (N_5302,N_3455,N_2629);
nor U5303 (N_5303,N_3761,N_2551);
or U5304 (N_5304,N_3819,N_3710);
nor U5305 (N_5305,N_3965,N_3878);
nor U5306 (N_5306,N_3161,N_2827);
or U5307 (N_5307,N_2966,N_3138);
nor U5308 (N_5308,N_3989,N_2193);
xnor U5309 (N_5309,N_3123,N_3439);
xnor U5310 (N_5310,N_2475,N_2693);
and U5311 (N_5311,N_3854,N_2527);
or U5312 (N_5312,N_2439,N_3866);
nand U5313 (N_5313,N_2613,N_3719);
xor U5314 (N_5314,N_2604,N_2363);
nand U5315 (N_5315,N_2091,N_3107);
or U5316 (N_5316,N_3706,N_2168);
and U5317 (N_5317,N_3011,N_3893);
or U5318 (N_5318,N_2153,N_3760);
xor U5319 (N_5319,N_3277,N_2836);
nand U5320 (N_5320,N_2028,N_2741);
xor U5321 (N_5321,N_2209,N_3942);
xor U5322 (N_5322,N_2363,N_2058);
nand U5323 (N_5323,N_3294,N_3933);
nand U5324 (N_5324,N_3541,N_2452);
and U5325 (N_5325,N_2588,N_2372);
xnor U5326 (N_5326,N_2451,N_3290);
nand U5327 (N_5327,N_3362,N_2483);
and U5328 (N_5328,N_3931,N_2177);
xnor U5329 (N_5329,N_3189,N_2055);
xnor U5330 (N_5330,N_2093,N_2992);
nand U5331 (N_5331,N_3953,N_3223);
xor U5332 (N_5332,N_2376,N_3755);
xnor U5333 (N_5333,N_2192,N_3643);
nand U5334 (N_5334,N_3690,N_2918);
or U5335 (N_5335,N_3933,N_3403);
and U5336 (N_5336,N_2222,N_3683);
or U5337 (N_5337,N_2451,N_2666);
nor U5338 (N_5338,N_3967,N_3730);
nor U5339 (N_5339,N_3892,N_3545);
nor U5340 (N_5340,N_2894,N_2829);
nand U5341 (N_5341,N_3217,N_3793);
xor U5342 (N_5342,N_3259,N_2021);
xor U5343 (N_5343,N_3934,N_3948);
and U5344 (N_5344,N_2432,N_3134);
xnor U5345 (N_5345,N_2572,N_2436);
and U5346 (N_5346,N_3025,N_3192);
nand U5347 (N_5347,N_3131,N_3099);
nor U5348 (N_5348,N_2235,N_3042);
xor U5349 (N_5349,N_3812,N_3085);
nand U5350 (N_5350,N_2336,N_2011);
nor U5351 (N_5351,N_2776,N_3043);
xor U5352 (N_5352,N_3369,N_3489);
or U5353 (N_5353,N_3836,N_2586);
and U5354 (N_5354,N_3410,N_2953);
nor U5355 (N_5355,N_3228,N_3196);
nand U5356 (N_5356,N_2413,N_3800);
and U5357 (N_5357,N_3641,N_3795);
and U5358 (N_5358,N_2535,N_3449);
nor U5359 (N_5359,N_3803,N_3654);
nand U5360 (N_5360,N_3679,N_2818);
nand U5361 (N_5361,N_3301,N_2369);
nor U5362 (N_5362,N_3211,N_2779);
xnor U5363 (N_5363,N_3761,N_2154);
or U5364 (N_5364,N_2103,N_2501);
xor U5365 (N_5365,N_2273,N_2594);
nand U5366 (N_5366,N_3381,N_2740);
or U5367 (N_5367,N_3460,N_3594);
or U5368 (N_5368,N_2322,N_2076);
and U5369 (N_5369,N_3857,N_2253);
and U5370 (N_5370,N_2878,N_2343);
nand U5371 (N_5371,N_2807,N_2285);
nand U5372 (N_5372,N_2009,N_2530);
nand U5373 (N_5373,N_3472,N_3203);
and U5374 (N_5374,N_3954,N_3566);
nand U5375 (N_5375,N_3931,N_3632);
nand U5376 (N_5376,N_2554,N_3475);
xor U5377 (N_5377,N_3924,N_3601);
and U5378 (N_5378,N_3537,N_2018);
or U5379 (N_5379,N_2614,N_2573);
nor U5380 (N_5380,N_2191,N_2308);
or U5381 (N_5381,N_3780,N_2404);
xnor U5382 (N_5382,N_2787,N_2898);
xnor U5383 (N_5383,N_3816,N_2106);
nor U5384 (N_5384,N_2265,N_2495);
or U5385 (N_5385,N_2442,N_3306);
xor U5386 (N_5386,N_3989,N_3647);
or U5387 (N_5387,N_3213,N_3494);
xnor U5388 (N_5388,N_3052,N_3966);
nand U5389 (N_5389,N_3544,N_2699);
or U5390 (N_5390,N_3823,N_3458);
nand U5391 (N_5391,N_2965,N_3391);
nand U5392 (N_5392,N_3409,N_2959);
nand U5393 (N_5393,N_3929,N_3445);
nand U5394 (N_5394,N_2177,N_3739);
nor U5395 (N_5395,N_2284,N_2676);
nand U5396 (N_5396,N_3660,N_3833);
and U5397 (N_5397,N_3095,N_2113);
nand U5398 (N_5398,N_3545,N_2124);
nand U5399 (N_5399,N_3749,N_3838);
xnor U5400 (N_5400,N_3903,N_3511);
or U5401 (N_5401,N_2015,N_2021);
and U5402 (N_5402,N_3700,N_3899);
or U5403 (N_5403,N_3646,N_2645);
xor U5404 (N_5404,N_2179,N_2503);
and U5405 (N_5405,N_2093,N_2269);
or U5406 (N_5406,N_2160,N_2586);
and U5407 (N_5407,N_2564,N_3331);
nand U5408 (N_5408,N_3007,N_3817);
xor U5409 (N_5409,N_2111,N_3110);
nand U5410 (N_5410,N_3839,N_3690);
nand U5411 (N_5411,N_3067,N_3044);
nor U5412 (N_5412,N_2329,N_3995);
and U5413 (N_5413,N_2776,N_2777);
xnor U5414 (N_5414,N_2687,N_3393);
nor U5415 (N_5415,N_2308,N_2466);
and U5416 (N_5416,N_3516,N_3720);
nor U5417 (N_5417,N_3844,N_3922);
and U5418 (N_5418,N_2858,N_3208);
or U5419 (N_5419,N_2127,N_3012);
and U5420 (N_5420,N_3496,N_3068);
or U5421 (N_5421,N_3281,N_3458);
or U5422 (N_5422,N_3241,N_3006);
or U5423 (N_5423,N_3783,N_3539);
nand U5424 (N_5424,N_3727,N_3161);
or U5425 (N_5425,N_2933,N_3038);
and U5426 (N_5426,N_2278,N_3253);
or U5427 (N_5427,N_2732,N_3443);
or U5428 (N_5428,N_2751,N_3951);
nor U5429 (N_5429,N_2751,N_2703);
and U5430 (N_5430,N_3937,N_2760);
xor U5431 (N_5431,N_3584,N_2081);
or U5432 (N_5432,N_3067,N_3712);
or U5433 (N_5433,N_3985,N_2563);
or U5434 (N_5434,N_2161,N_2914);
nor U5435 (N_5435,N_3320,N_2464);
and U5436 (N_5436,N_3121,N_3684);
and U5437 (N_5437,N_2201,N_2435);
or U5438 (N_5438,N_2619,N_2567);
xnor U5439 (N_5439,N_2092,N_3398);
xnor U5440 (N_5440,N_3175,N_3935);
nor U5441 (N_5441,N_3775,N_2267);
or U5442 (N_5442,N_3047,N_3707);
nand U5443 (N_5443,N_2643,N_2776);
xor U5444 (N_5444,N_2946,N_3977);
nand U5445 (N_5445,N_3743,N_3368);
nor U5446 (N_5446,N_3485,N_2180);
nor U5447 (N_5447,N_3257,N_3443);
nand U5448 (N_5448,N_2877,N_2115);
nor U5449 (N_5449,N_2789,N_2699);
nand U5450 (N_5450,N_3070,N_3670);
and U5451 (N_5451,N_3603,N_3549);
xor U5452 (N_5452,N_2190,N_2216);
xor U5453 (N_5453,N_3079,N_2137);
nand U5454 (N_5454,N_3084,N_2098);
nor U5455 (N_5455,N_3794,N_3700);
nand U5456 (N_5456,N_3326,N_2750);
or U5457 (N_5457,N_3466,N_2395);
and U5458 (N_5458,N_2237,N_2486);
or U5459 (N_5459,N_3931,N_3455);
nand U5460 (N_5460,N_3827,N_2732);
nor U5461 (N_5461,N_2973,N_3091);
xor U5462 (N_5462,N_2596,N_3449);
and U5463 (N_5463,N_3582,N_3029);
and U5464 (N_5464,N_2553,N_2668);
nand U5465 (N_5465,N_3502,N_2993);
nand U5466 (N_5466,N_3218,N_2912);
or U5467 (N_5467,N_3219,N_2895);
xnor U5468 (N_5468,N_2327,N_2812);
or U5469 (N_5469,N_3855,N_3391);
or U5470 (N_5470,N_2913,N_2218);
and U5471 (N_5471,N_2765,N_3068);
and U5472 (N_5472,N_3020,N_3546);
and U5473 (N_5473,N_2638,N_2231);
nand U5474 (N_5474,N_3242,N_2698);
and U5475 (N_5475,N_2702,N_2522);
nand U5476 (N_5476,N_3205,N_2571);
xor U5477 (N_5477,N_3791,N_2483);
nor U5478 (N_5478,N_3174,N_2675);
nor U5479 (N_5479,N_3105,N_2936);
or U5480 (N_5480,N_2109,N_3118);
nand U5481 (N_5481,N_2673,N_3244);
xnor U5482 (N_5482,N_2177,N_2443);
xor U5483 (N_5483,N_3236,N_3064);
nor U5484 (N_5484,N_3420,N_3231);
or U5485 (N_5485,N_3939,N_3147);
xnor U5486 (N_5486,N_2850,N_2250);
xnor U5487 (N_5487,N_2005,N_2178);
and U5488 (N_5488,N_2407,N_3915);
nor U5489 (N_5489,N_2977,N_3593);
xor U5490 (N_5490,N_3754,N_2625);
nor U5491 (N_5491,N_3737,N_2553);
and U5492 (N_5492,N_2876,N_2303);
nand U5493 (N_5493,N_2243,N_3343);
xor U5494 (N_5494,N_3102,N_2709);
and U5495 (N_5495,N_3196,N_2031);
or U5496 (N_5496,N_3013,N_3828);
and U5497 (N_5497,N_2232,N_3207);
or U5498 (N_5498,N_3811,N_3087);
and U5499 (N_5499,N_2571,N_2771);
or U5500 (N_5500,N_2209,N_2976);
nand U5501 (N_5501,N_3369,N_3002);
nor U5502 (N_5502,N_3310,N_2419);
nor U5503 (N_5503,N_3726,N_2341);
nor U5504 (N_5504,N_3299,N_2868);
xor U5505 (N_5505,N_2988,N_3664);
or U5506 (N_5506,N_2717,N_3513);
nand U5507 (N_5507,N_2335,N_3219);
nor U5508 (N_5508,N_2847,N_3531);
nor U5509 (N_5509,N_2416,N_3123);
or U5510 (N_5510,N_2878,N_2029);
nand U5511 (N_5511,N_3093,N_3350);
nand U5512 (N_5512,N_3506,N_2583);
and U5513 (N_5513,N_3061,N_3632);
xnor U5514 (N_5514,N_3947,N_2761);
and U5515 (N_5515,N_3158,N_2834);
and U5516 (N_5516,N_3340,N_2275);
or U5517 (N_5517,N_2049,N_3883);
and U5518 (N_5518,N_2129,N_2330);
nor U5519 (N_5519,N_2623,N_3715);
and U5520 (N_5520,N_2422,N_2187);
xnor U5521 (N_5521,N_2734,N_3909);
xnor U5522 (N_5522,N_2840,N_3290);
and U5523 (N_5523,N_2637,N_3012);
or U5524 (N_5524,N_2156,N_2581);
or U5525 (N_5525,N_2561,N_2103);
or U5526 (N_5526,N_2472,N_3624);
nor U5527 (N_5527,N_3558,N_2543);
and U5528 (N_5528,N_3117,N_2777);
and U5529 (N_5529,N_3448,N_3382);
and U5530 (N_5530,N_2195,N_2492);
or U5531 (N_5531,N_3257,N_2037);
xor U5532 (N_5532,N_3873,N_2820);
nand U5533 (N_5533,N_3051,N_3027);
nand U5534 (N_5534,N_2112,N_2632);
nor U5535 (N_5535,N_2334,N_2372);
and U5536 (N_5536,N_2217,N_2556);
or U5537 (N_5537,N_3579,N_2468);
xor U5538 (N_5538,N_2927,N_2241);
nand U5539 (N_5539,N_2803,N_2992);
nand U5540 (N_5540,N_3020,N_3884);
xnor U5541 (N_5541,N_3776,N_3606);
nor U5542 (N_5542,N_3498,N_2888);
nor U5543 (N_5543,N_3979,N_3672);
nand U5544 (N_5544,N_3547,N_3786);
and U5545 (N_5545,N_2064,N_2346);
or U5546 (N_5546,N_2809,N_2068);
or U5547 (N_5547,N_3110,N_2076);
and U5548 (N_5548,N_2102,N_2334);
nor U5549 (N_5549,N_2926,N_3486);
nand U5550 (N_5550,N_3935,N_3764);
xor U5551 (N_5551,N_3231,N_3045);
and U5552 (N_5552,N_2313,N_2693);
and U5553 (N_5553,N_3465,N_2352);
nor U5554 (N_5554,N_3186,N_2966);
and U5555 (N_5555,N_2133,N_3811);
and U5556 (N_5556,N_3029,N_2346);
nand U5557 (N_5557,N_2481,N_2294);
nand U5558 (N_5558,N_3857,N_3678);
xnor U5559 (N_5559,N_3570,N_2584);
nor U5560 (N_5560,N_3364,N_3359);
and U5561 (N_5561,N_2117,N_2213);
xor U5562 (N_5562,N_2047,N_3156);
nor U5563 (N_5563,N_2930,N_2777);
and U5564 (N_5564,N_3709,N_2195);
xor U5565 (N_5565,N_2132,N_3374);
nor U5566 (N_5566,N_2610,N_3072);
and U5567 (N_5567,N_3321,N_2845);
xor U5568 (N_5568,N_3063,N_2140);
nand U5569 (N_5569,N_2661,N_3506);
and U5570 (N_5570,N_3426,N_3322);
nor U5571 (N_5571,N_2772,N_2304);
or U5572 (N_5572,N_3679,N_2300);
nand U5573 (N_5573,N_3489,N_3954);
and U5574 (N_5574,N_2426,N_3457);
and U5575 (N_5575,N_2622,N_2267);
xor U5576 (N_5576,N_2386,N_2644);
or U5577 (N_5577,N_2610,N_3094);
and U5578 (N_5578,N_3487,N_3011);
nor U5579 (N_5579,N_3678,N_3040);
and U5580 (N_5580,N_3966,N_2372);
xnor U5581 (N_5581,N_2572,N_3995);
nor U5582 (N_5582,N_2346,N_3399);
or U5583 (N_5583,N_2869,N_3094);
and U5584 (N_5584,N_2909,N_3767);
xor U5585 (N_5585,N_3772,N_2158);
or U5586 (N_5586,N_3796,N_3831);
xor U5587 (N_5587,N_3565,N_3378);
nor U5588 (N_5588,N_3714,N_3183);
xor U5589 (N_5589,N_2796,N_2046);
and U5590 (N_5590,N_2368,N_2679);
nor U5591 (N_5591,N_3604,N_3519);
xor U5592 (N_5592,N_3832,N_3264);
nand U5593 (N_5593,N_2488,N_2545);
nand U5594 (N_5594,N_3700,N_3643);
or U5595 (N_5595,N_3193,N_2436);
or U5596 (N_5596,N_2419,N_3843);
or U5597 (N_5597,N_3573,N_2433);
nor U5598 (N_5598,N_3216,N_2563);
xnor U5599 (N_5599,N_2139,N_3930);
or U5600 (N_5600,N_2772,N_3099);
and U5601 (N_5601,N_3836,N_2541);
nor U5602 (N_5602,N_3164,N_3753);
nand U5603 (N_5603,N_2966,N_3449);
and U5604 (N_5604,N_3052,N_3500);
or U5605 (N_5605,N_2895,N_2144);
xnor U5606 (N_5606,N_3035,N_2191);
or U5607 (N_5607,N_2462,N_2187);
xor U5608 (N_5608,N_3670,N_3399);
nor U5609 (N_5609,N_3056,N_2973);
and U5610 (N_5610,N_2609,N_2917);
or U5611 (N_5611,N_2572,N_2868);
and U5612 (N_5612,N_3317,N_3626);
nor U5613 (N_5613,N_2033,N_3884);
nor U5614 (N_5614,N_3668,N_2148);
xnor U5615 (N_5615,N_2888,N_3666);
and U5616 (N_5616,N_3981,N_2175);
xor U5617 (N_5617,N_2030,N_2455);
nand U5618 (N_5618,N_2951,N_2574);
or U5619 (N_5619,N_3499,N_3860);
nand U5620 (N_5620,N_2349,N_3227);
nor U5621 (N_5621,N_3547,N_2868);
xor U5622 (N_5622,N_2834,N_2825);
nor U5623 (N_5623,N_3739,N_3149);
xnor U5624 (N_5624,N_2241,N_3682);
xnor U5625 (N_5625,N_3839,N_2149);
nor U5626 (N_5626,N_2786,N_2533);
xor U5627 (N_5627,N_3374,N_2955);
and U5628 (N_5628,N_2863,N_3314);
xor U5629 (N_5629,N_2618,N_3964);
or U5630 (N_5630,N_2187,N_3390);
nand U5631 (N_5631,N_3540,N_3636);
nor U5632 (N_5632,N_3673,N_3524);
or U5633 (N_5633,N_2336,N_2711);
and U5634 (N_5634,N_3298,N_2264);
or U5635 (N_5635,N_2020,N_3104);
and U5636 (N_5636,N_2969,N_2769);
nand U5637 (N_5637,N_2319,N_2942);
or U5638 (N_5638,N_2064,N_3303);
and U5639 (N_5639,N_2796,N_3643);
nand U5640 (N_5640,N_2635,N_2262);
nor U5641 (N_5641,N_3228,N_3188);
nor U5642 (N_5642,N_2866,N_2619);
or U5643 (N_5643,N_3115,N_2863);
and U5644 (N_5644,N_2770,N_2549);
and U5645 (N_5645,N_3874,N_3453);
xnor U5646 (N_5646,N_2750,N_3320);
nor U5647 (N_5647,N_2205,N_3379);
nor U5648 (N_5648,N_2001,N_2364);
nor U5649 (N_5649,N_3082,N_2080);
or U5650 (N_5650,N_2287,N_3849);
or U5651 (N_5651,N_2287,N_2425);
nor U5652 (N_5652,N_3255,N_2682);
nor U5653 (N_5653,N_2171,N_3761);
xnor U5654 (N_5654,N_3841,N_3291);
nor U5655 (N_5655,N_3901,N_3250);
or U5656 (N_5656,N_2245,N_2424);
and U5657 (N_5657,N_2123,N_2534);
or U5658 (N_5658,N_2393,N_2497);
nand U5659 (N_5659,N_3486,N_3398);
nand U5660 (N_5660,N_3515,N_3160);
xnor U5661 (N_5661,N_2654,N_2708);
nor U5662 (N_5662,N_2135,N_2615);
or U5663 (N_5663,N_3160,N_3867);
nor U5664 (N_5664,N_3236,N_2730);
nor U5665 (N_5665,N_3862,N_3691);
and U5666 (N_5666,N_2608,N_3784);
nand U5667 (N_5667,N_3064,N_3177);
and U5668 (N_5668,N_2794,N_2089);
nor U5669 (N_5669,N_2561,N_2306);
nand U5670 (N_5670,N_3202,N_3331);
nor U5671 (N_5671,N_3296,N_3641);
and U5672 (N_5672,N_2498,N_3659);
and U5673 (N_5673,N_2604,N_3620);
and U5674 (N_5674,N_3157,N_2484);
nand U5675 (N_5675,N_3814,N_2411);
nand U5676 (N_5676,N_2855,N_3011);
and U5677 (N_5677,N_3996,N_3187);
and U5678 (N_5678,N_3327,N_2604);
nor U5679 (N_5679,N_3873,N_2106);
xor U5680 (N_5680,N_2017,N_3598);
nor U5681 (N_5681,N_3368,N_3921);
and U5682 (N_5682,N_2678,N_2338);
nor U5683 (N_5683,N_2568,N_2093);
or U5684 (N_5684,N_3514,N_2577);
nand U5685 (N_5685,N_3086,N_3782);
and U5686 (N_5686,N_3968,N_3664);
and U5687 (N_5687,N_2515,N_3424);
xor U5688 (N_5688,N_3113,N_3393);
and U5689 (N_5689,N_3726,N_2821);
nor U5690 (N_5690,N_3078,N_3990);
xnor U5691 (N_5691,N_2407,N_2235);
xnor U5692 (N_5692,N_3930,N_3902);
and U5693 (N_5693,N_2656,N_3795);
or U5694 (N_5694,N_2299,N_3327);
nor U5695 (N_5695,N_3095,N_3449);
nand U5696 (N_5696,N_3964,N_3479);
and U5697 (N_5697,N_3564,N_3815);
xnor U5698 (N_5698,N_3124,N_2364);
nand U5699 (N_5699,N_3096,N_2400);
or U5700 (N_5700,N_3014,N_3186);
nand U5701 (N_5701,N_3841,N_3591);
and U5702 (N_5702,N_3887,N_2857);
nor U5703 (N_5703,N_2922,N_2091);
xnor U5704 (N_5704,N_2325,N_3178);
nor U5705 (N_5705,N_2550,N_2425);
and U5706 (N_5706,N_3580,N_2990);
or U5707 (N_5707,N_2779,N_2137);
nor U5708 (N_5708,N_3705,N_3047);
nand U5709 (N_5709,N_2504,N_3454);
and U5710 (N_5710,N_3883,N_3943);
nand U5711 (N_5711,N_2190,N_2831);
or U5712 (N_5712,N_2615,N_2160);
and U5713 (N_5713,N_3603,N_3797);
nor U5714 (N_5714,N_3418,N_3898);
nand U5715 (N_5715,N_2993,N_2007);
and U5716 (N_5716,N_2745,N_3038);
nand U5717 (N_5717,N_3001,N_2364);
and U5718 (N_5718,N_2832,N_3519);
nor U5719 (N_5719,N_3264,N_2931);
xor U5720 (N_5720,N_2830,N_2106);
and U5721 (N_5721,N_3530,N_3181);
or U5722 (N_5722,N_2276,N_2839);
nand U5723 (N_5723,N_3990,N_3208);
xnor U5724 (N_5724,N_2408,N_3403);
or U5725 (N_5725,N_3804,N_2550);
and U5726 (N_5726,N_2549,N_3623);
nand U5727 (N_5727,N_2026,N_3552);
or U5728 (N_5728,N_3736,N_3537);
nor U5729 (N_5729,N_2195,N_3251);
nor U5730 (N_5730,N_2182,N_2318);
nor U5731 (N_5731,N_2874,N_3631);
nand U5732 (N_5732,N_3691,N_2495);
xnor U5733 (N_5733,N_3058,N_3390);
nor U5734 (N_5734,N_2705,N_2035);
nor U5735 (N_5735,N_2538,N_2745);
nor U5736 (N_5736,N_2843,N_3228);
nor U5737 (N_5737,N_3714,N_2300);
nand U5738 (N_5738,N_3844,N_2485);
and U5739 (N_5739,N_3774,N_2686);
or U5740 (N_5740,N_3060,N_3868);
nor U5741 (N_5741,N_2264,N_3698);
and U5742 (N_5742,N_3407,N_3536);
or U5743 (N_5743,N_3582,N_3758);
or U5744 (N_5744,N_3044,N_2969);
and U5745 (N_5745,N_3478,N_3465);
xor U5746 (N_5746,N_2189,N_3368);
or U5747 (N_5747,N_3872,N_2766);
nor U5748 (N_5748,N_2672,N_3685);
nor U5749 (N_5749,N_3362,N_2564);
nand U5750 (N_5750,N_3654,N_2228);
xor U5751 (N_5751,N_2920,N_3186);
nand U5752 (N_5752,N_2183,N_3232);
or U5753 (N_5753,N_3918,N_3327);
and U5754 (N_5754,N_3761,N_2189);
nor U5755 (N_5755,N_2024,N_2842);
xor U5756 (N_5756,N_3561,N_3978);
nand U5757 (N_5757,N_3945,N_2891);
and U5758 (N_5758,N_3431,N_3103);
nand U5759 (N_5759,N_2338,N_3108);
or U5760 (N_5760,N_2531,N_2090);
and U5761 (N_5761,N_2961,N_2592);
nor U5762 (N_5762,N_3377,N_2705);
nand U5763 (N_5763,N_3099,N_3744);
or U5764 (N_5764,N_3491,N_3801);
nand U5765 (N_5765,N_2978,N_3243);
nand U5766 (N_5766,N_2779,N_3877);
and U5767 (N_5767,N_3653,N_3868);
and U5768 (N_5768,N_2667,N_2129);
xnor U5769 (N_5769,N_3397,N_3727);
nand U5770 (N_5770,N_2886,N_3976);
and U5771 (N_5771,N_2574,N_2949);
nand U5772 (N_5772,N_3775,N_2868);
nand U5773 (N_5773,N_2449,N_2880);
and U5774 (N_5774,N_3530,N_3001);
nor U5775 (N_5775,N_3920,N_3599);
nand U5776 (N_5776,N_2113,N_3984);
xor U5777 (N_5777,N_3424,N_3250);
and U5778 (N_5778,N_2925,N_2042);
or U5779 (N_5779,N_3780,N_3606);
and U5780 (N_5780,N_2577,N_3354);
or U5781 (N_5781,N_2093,N_2392);
or U5782 (N_5782,N_3543,N_2471);
or U5783 (N_5783,N_3081,N_3936);
or U5784 (N_5784,N_3553,N_2774);
xor U5785 (N_5785,N_2385,N_2045);
nand U5786 (N_5786,N_2166,N_3889);
nand U5787 (N_5787,N_2159,N_2767);
nand U5788 (N_5788,N_2756,N_2555);
xnor U5789 (N_5789,N_3795,N_2349);
nor U5790 (N_5790,N_3109,N_3927);
nand U5791 (N_5791,N_2398,N_3439);
nand U5792 (N_5792,N_3374,N_3389);
xor U5793 (N_5793,N_3032,N_2598);
and U5794 (N_5794,N_2303,N_3232);
nor U5795 (N_5795,N_3576,N_3277);
nor U5796 (N_5796,N_3432,N_3597);
xor U5797 (N_5797,N_3516,N_3938);
xor U5798 (N_5798,N_3279,N_2636);
or U5799 (N_5799,N_3541,N_3676);
xor U5800 (N_5800,N_3459,N_3198);
nor U5801 (N_5801,N_2480,N_3667);
or U5802 (N_5802,N_3439,N_3824);
nand U5803 (N_5803,N_3713,N_2765);
nand U5804 (N_5804,N_2282,N_2691);
and U5805 (N_5805,N_2958,N_2554);
xnor U5806 (N_5806,N_2271,N_3023);
and U5807 (N_5807,N_2441,N_3749);
and U5808 (N_5808,N_2178,N_2281);
or U5809 (N_5809,N_3755,N_3963);
nand U5810 (N_5810,N_3892,N_2864);
xor U5811 (N_5811,N_3715,N_2647);
or U5812 (N_5812,N_3755,N_3057);
xor U5813 (N_5813,N_2371,N_2249);
and U5814 (N_5814,N_2228,N_3162);
xor U5815 (N_5815,N_2182,N_3662);
xnor U5816 (N_5816,N_2197,N_3571);
xnor U5817 (N_5817,N_3522,N_2673);
nor U5818 (N_5818,N_2439,N_3722);
or U5819 (N_5819,N_2259,N_2464);
xor U5820 (N_5820,N_2793,N_2748);
xor U5821 (N_5821,N_3394,N_2337);
and U5822 (N_5822,N_2212,N_2143);
or U5823 (N_5823,N_3624,N_3387);
nor U5824 (N_5824,N_2772,N_3211);
nor U5825 (N_5825,N_3625,N_2992);
xnor U5826 (N_5826,N_3115,N_3014);
nand U5827 (N_5827,N_2136,N_2186);
and U5828 (N_5828,N_2964,N_3857);
xnor U5829 (N_5829,N_2321,N_2804);
xor U5830 (N_5830,N_3163,N_2517);
and U5831 (N_5831,N_2887,N_3526);
nand U5832 (N_5832,N_2374,N_3628);
xnor U5833 (N_5833,N_3939,N_2251);
nand U5834 (N_5834,N_3595,N_3001);
and U5835 (N_5835,N_3519,N_2414);
and U5836 (N_5836,N_2524,N_2384);
or U5837 (N_5837,N_3885,N_3139);
xnor U5838 (N_5838,N_2426,N_2633);
nand U5839 (N_5839,N_3602,N_2501);
nand U5840 (N_5840,N_2036,N_3022);
xnor U5841 (N_5841,N_3665,N_3777);
nand U5842 (N_5842,N_3230,N_2051);
or U5843 (N_5843,N_3372,N_3437);
or U5844 (N_5844,N_2404,N_2167);
nand U5845 (N_5845,N_2014,N_3904);
nand U5846 (N_5846,N_2532,N_3239);
and U5847 (N_5847,N_2058,N_3617);
and U5848 (N_5848,N_3446,N_3280);
nor U5849 (N_5849,N_3171,N_2633);
nor U5850 (N_5850,N_2962,N_2416);
nand U5851 (N_5851,N_3180,N_3616);
nor U5852 (N_5852,N_3387,N_2046);
or U5853 (N_5853,N_2744,N_3052);
or U5854 (N_5854,N_3889,N_3555);
nor U5855 (N_5855,N_3352,N_2124);
or U5856 (N_5856,N_2465,N_2139);
or U5857 (N_5857,N_2471,N_2487);
or U5858 (N_5858,N_2623,N_3161);
xnor U5859 (N_5859,N_3394,N_2344);
nor U5860 (N_5860,N_2194,N_2565);
or U5861 (N_5861,N_2473,N_3816);
or U5862 (N_5862,N_2575,N_3283);
nand U5863 (N_5863,N_2917,N_3950);
nor U5864 (N_5864,N_3582,N_2275);
xor U5865 (N_5865,N_2662,N_3143);
nand U5866 (N_5866,N_2401,N_2599);
or U5867 (N_5867,N_2272,N_3915);
and U5868 (N_5868,N_3555,N_3395);
xnor U5869 (N_5869,N_2920,N_2637);
or U5870 (N_5870,N_2690,N_2409);
or U5871 (N_5871,N_2513,N_2849);
nand U5872 (N_5872,N_3277,N_3508);
xnor U5873 (N_5873,N_3090,N_3533);
nand U5874 (N_5874,N_2581,N_2510);
and U5875 (N_5875,N_2042,N_3604);
nor U5876 (N_5876,N_2837,N_2571);
or U5877 (N_5877,N_2790,N_2488);
or U5878 (N_5878,N_3063,N_2108);
nor U5879 (N_5879,N_3017,N_3502);
nor U5880 (N_5880,N_2233,N_3958);
and U5881 (N_5881,N_2931,N_2082);
or U5882 (N_5882,N_3480,N_3356);
xnor U5883 (N_5883,N_2444,N_2331);
and U5884 (N_5884,N_2163,N_3205);
or U5885 (N_5885,N_2153,N_3566);
and U5886 (N_5886,N_3048,N_3823);
nor U5887 (N_5887,N_3494,N_2949);
nand U5888 (N_5888,N_2547,N_2787);
nand U5889 (N_5889,N_2969,N_3746);
nand U5890 (N_5890,N_2268,N_2471);
nand U5891 (N_5891,N_2580,N_3672);
or U5892 (N_5892,N_3989,N_2423);
and U5893 (N_5893,N_2060,N_2993);
nor U5894 (N_5894,N_3468,N_2678);
xor U5895 (N_5895,N_3789,N_2617);
and U5896 (N_5896,N_2579,N_3463);
or U5897 (N_5897,N_3616,N_3673);
nand U5898 (N_5898,N_2802,N_3304);
or U5899 (N_5899,N_3972,N_3329);
nor U5900 (N_5900,N_3785,N_3439);
xnor U5901 (N_5901,N_2439,N_3055);
nand U5902 (N_5902,N_2659,N_3858);
and U5903 (N_5903,N_2156,N_2459);
or U5904 (N_5904,N_3826,N_3462);
nand U5905 (N_5905,N_2427,N_3157);
nand U5906 (N_5906,N_2961,N_2925);
xnor U5907 (N_5907,N_3275,N_2996);
and U5908 (N_5908,N_3368,N_2688);
nand U5909 (N_5909,N_2683,N_2096);
nor U5910 (N_5910,N_3590,N_3078);
nor U5911 (N_5911,N_2428,N_3735);
nand U5912 (N_5912,N_3856,N_3398);
or U5913 (N_5913,N_2976,N_2662);
xor U5914 (N_5914,N_3983,N_2871);
xor U5915 (N_5915,N_3089,N_3749);
nand U5916 (N_5916,N_2236,N_2857);
nand U5917 (N_5917,N_3266,N_2090);
or U5918 (N_5918,N_3486,N_2524);
and U5919 (N_5919,N_3411,N_2211);
or U5920 (N_5920,N_2060,N_2874);
and U5921 (N_5921,N_3706,N_3981);
nor U5922 (N_5922,N_2400,N_3434);
xor U5923 (N_5923,N_2620,N_2466);
or U5924 (N_5924,N_3450,N_3465);
nand U5925 (N_5925,N_3899,N_2672);
or U5926 (N_5926,N_2833,N_3532);
nor U5927 (N_5927,N_3233,N_3770);
nand U5928 (N_5928,N_3167,N_3696);
nand U5929 (N_5929,N_3203,N_2125);
nand U5930 (N_5930,N_2677,N_3470);
nand U5931 (N_5931,N_2990,N_3189);
xor U5932 (N_5932,N_3905,N_2899);
and U5933 (N_5933,N_3154,N_2821);
nor U5934 (N_5934,N_2354,N_2847);
nand U5935 (N_5935,N_3678,N_3229);
nand U5936 (N_5936,N_2599,N_3322);
xor U5937 (N_5937,N_2962,N_3705);
and U5938 (N_5938,N_2096,N_3614);
nand U5939 (N_5939,N_3045,N_3416);
and U5940 (N_5940,N_3926,N_2255);
or U5941 (N_5941,N_3315,N_3980);
nor U5942 (N_5942,N_3958,N_3064);
xnor U5943 (N_5943,N_2124,N_2101);
or U5944 (N_5944,N_3052,N_3944);
or U5945 (N_5945,N_3257,N_2785);
and U5946 (N_5946,N_2704,N_3851);
nand U5947 (N_5947,N_3562,N_2512);
or U5948 (N_5948,N_2576,N_2621);
and U5949 (N_5949,N_2818,N_3401);
xnor U5950 (N_5950,N_3216,N_3017);
or U5951 (N_5951,N_2897,N_2720);
nor U5952 (N_5952,N_2250,N_2411);
xnor U5953 (N_5953,N_2520,N_3606);
or U5954 (N_5954,N_2862,N_3097);
xor U5955 (N_5955,N_3996,N_2451);
or U5956 (N_5956,N_2875,N_2154);
and U5957 (N_5957,N_3242,N_2451);
nand U5958 (N_5958,N_3941,N_2269);
nand U5959 (N_5959,N_2973,N_2982);
nand U5960 (N_5960,N_3047,N_2068);
or U5961 (N_5961,N_2481,N_2687);
xor U5962 (N_5962,N_2837,N_2601);
xor U5963 (N_5963,N_2294,N_2426);
and U5964 (N_5964,N_3373,N_2587);
xor U5965 (N_5965,N_3315,N_2346);
nor U5966 (N_5966,N_2058,N_3060);
and U5967 (N_5967,N_2544,N_3980);
nand U5968 (N_5968,N_2099,N_2034);
nand U5969 (N_5969,N_2183,N_3105);
and U5970 (N_5970,N_3518,N_3580);
xnor U5971 (N_5971,N_3207,N_3393);
xnor U5972 (N_5972,N_3627,N_3749);
or U5973 (N_5973,N_3527,N_2962);
nor U5974 (N_5974,N_3997,N_3491);
nor U5975 (N_5975,N_2975,N_3720);
or U5976 (N_5976,N_3573,N_3396);
nand U5977 (N_5977,N_2730,N_3497);
xnor U5978 (N_5978,N_2180,N_2937);
or U5979 (N_5979,N_3629,N_3121);
nand U5980 (N_5980,N_2785,N_3026);
and U5981 (N_5981,N_3357,N_2853);
nand U5982 (N_5982,N_2641,N_3203);
xnor U5983 (N_5983,N_2013,N_2856);
or U5984 (N_5984,N_2692,N_3132);
nor U5985 (N_5985,N_2200,N_3150);
nor U5986 (N_5986,N_2035,N_3330);
nand U5987 (N_5987,N_2350,N_2792);
xnor U5988 (N_5988,N_2595,N_3793);
or U5989 (N_5989,N_2949,N_3764);
nor U5990 (N_5990,N_3901,N_3628);
nor U5991 (N_5991,N_2670,N_2005);
nor U5992 (N_5992,N_3425,N_2937);
nand U5993 (N_5993,N_2700,N_2392);
nand U5994 (N_5994,N_2434,N_3429);
or U5995 (N_5995,N_2786,N_2792);
xor U5996 (N_5996,N_2090,N_2283);
xor U5997 (N_5997,N_2122,N_3982);
or U5998 (N_5998,N_2117,N_2321);
nand U5999 (N_5999,N_3311,N_3939);
or U6000 (N_6000,N_4616,N_5429);
xnor U6001 (N_6001,N_4836,N_5189);
and U6002 (N_6002,N_4583,N_5185);
xor U6003 (N_6003,N_5918,N_4303);
or U6004 (N_6004,N_5818,N_4174);
or U6005 (N_6005,N_5486,N_4342);
nand U6006 (N_6006,N_5014,N_5625);
xnor U6007 (N_6007,N_5313,N_5238);
nor U6008 (N_6008,N_4697,N_5096);
or U6009 (N_6009,N_4282,N_4129);
nor U6010 (N_6010,N_5754,N_5536);
or U6011 (N_6011,N_4851,N_4821);
and U6012 (N_6012,N_4216,N_4768);
xnor U6013 (N_6013,N_5632,N_4491);
xor U6014 (N_6014,N_4354,N_5514);
and U6015 (N_6015,N_5959,N_4134);
nand U6016 (N_6016,N_5018,N_4476);
or U6017 (N_6017,N_4399,N_4553);
or U6018 (N_6018,N_5041,N_4034);
nand U6019 (N_6019,N_5676,N_4474);
and U6020 (N_6020,N_4153,N_4818);
and U6021 (N_6021,N_5762,N_4597);
nand U6022 (N_6022,N_5215,N_4906);
nor U6023 (N_6023,N_4338,N_5957);
and U6024 (N_6024,N_4519,N_4205);
nor U6025 (N_6025,N_4409,N_5944);
nand U6026 (N_6026,N_5589,N_5262);
nand U6027 (N_6027,N_4295,N_4899);
or U6028 (N_6028,N_5115,N_4149);
or U6029 (N_6029,N_5023,N_4150);
nand U6030 (N_6030,N_5979,N_5803);
xor U6031 (N_6031,N_5225,N_5424);
and U6032 (N_6032,N_4707,N_5022);
and U6033 (N_6033,N_5922,N_5111);
nand U6034 (N_6034,N_4085,N_4680);
and U6035 (N_6035,N_5091,N_5745);
nor U6036 (N_6036,N_5905,N_4739);
xor U6037 (N_6037,N_4652,N_5743);
nor U6038 (N_6038,N_4865,N_5988);
and U6039 (N_6039,N_5511,N_4656);
nand U6040 (N_6040,N_4179,N_5492);
nor U6041 (N_6041,N_5274,N_5320);
and U6042 (N_6042,N_4459,N_5484);
or U6043 (N_6043,N_4671,N_5688);
or U6044 (N_6044,N_4941,N_4239);
and U6045 (N_6045,N_4943,N_5124);
nand U6046 (N_6046,N_4376,N_4223);
or U6047 (N_6047,N_5611,N_4933);
xnor U6048 (N_6048,N_5706,N_4277);
and U6049 (N_6049,N_4892,N_5002);
or U6050 (N_6050,N_4402,N_5981);
or U6051 (N_6051,N_4250,N_5519);
nand U6052 (N_6052,N_5788,N_4547);
nor U6053 (N_6053,N_4572,N_5744);
and U6054 (N_6054,N_4956,N_5971);
nand U6055 (N_6055,N_4695,N_5452);
or U6056 (N_6056,N_5691,N_4591);
or U6057 (N_6057,N_5107,N_5937);
or U6058 (N_6058,N_4729,N_5212);
and U6059 (N_6059,N_4189,N_4323);
or U6060 (N_6060,N_4646,N_4903);
nor U6061 (N_6061,N_5456,N_5904);
and U6062 (N_6062,N_5213,N_4191);
or U6063 (N_6063,N_4738,N_5813);
or U6064 (N_6064,N_4766,N_5682);
and U6065 (N_6065,N_4214,N_4701);
and U6066 (N_6066,N_4651,N_5100);
nor U6067 (N_6067,N_5701,N_5050);
and U6068 (N_6068,N_4820,N_5928);
xnor U6069 (N_6069,N_4272,N_5074);
or U6070 (N_6070,N_4421,N_5112);
nor U6071 (N_6071,N_4114,N_5304);
or U6072 (N_6072,N_5653,N_5357);
nand U6073 (N_6073,N_5311,N_5787);
xor U6074 (N_6074,N_5325,N_5098);
or U6075 (N_6075,N_5746,N_4942);
nand U6076 (N_6076,N_5872,N_4552);
xnor U6077 (N_6077,N_5224,N_5403);
nand U6078 (N_6078,N_5640,N_5896);
xnor U6079 (N_6079,N_5425,N_4925);
nand U6080 (N_6080,N_5468,N_5533);
xor U6081 (N_6081,N_4884,N_4703);
nor U6082 (N_6082,N_5666,N_4918);
or U6083 (N_6083,N_5055,N_5470);
xnor U6084 (N_6084,N_4046,N_5868);
xor U6085 (N_6085,N_4613,N_5651);
nor U6086 (N_6086,N_4245,N_5817);
or U6087 (N_6087,N_4015,N_5463);
xor U6088 (N_6088,N_4938,N_4507);
or U6089 (N_6089,N_4844,N_4447);
nand U6090 (N_6090,N_4281,N_4091);
or U6091 (N_6091,N_4353,N_5349);
and U6092 (N_6092,N_4193,N_5363);
nand U6093 (N_6093,N_4551,N_5206);
and U6094 (N_6094,N_4914,N_5563);
nand U6095 (N_6095,N_5503,N_4681);
or U6096 (N_6096,N_4894,N_5087);
nand U6097 (N_6097,N_5013,N_4458);
nor U6098 (N_6098,N_4244,N_4582);
nor U6099 (N_6099,N_5732,N_4740);
or U6100 (N_6100,N_5920,N_4708);
or U6101 (N_6101,N_4994,N_5646);
nand U6102 (N_6102,N_5901,N_5370);
nor U6103 (N_6103,N_5030,N_5007);
or U6104 (N_6104,N_4722,N_4158);
xnor U6105 (N_6105,N_4575,N_4518);
nor U6106 (N_6106,N_4837,N_4356);
nor U6107 (N_6107,N_5358,N_4144);
nand U6108 (N_6108,N_4562,N_4784);
nor U6109 (N_6109,N_4104,N_4327);
nor U6110 (N_6110,N_4999,N_5218);
xnor U6111 (N_6111,N_4333,N_5902);
xor U6112 (N_6112,N_4383,N_4684);
nor U6113 (N_6113,N_4287,N_4005);
xor U6114 (N_6114,N_5512,N_4025);
nand U6115 (N_6115,N_5652,N_4991);
nand U6116 (N_6116,N_5941,N_4457);
nor U6117 (N_6117,N_5807,N_4544);
nor U6118 (N_6118,N_4390,N_4247);
nand U6119 (N_6119,N_4389,N_4175);
nor U6120 (N_6120,N_5581,N_4319);
and U6121 (N_6121,N_5889,N_4027);
and U6122 (N_6122,N_5373,N_4312);
or U6123 (N_6123,N_4139,N_4964);
xor U6124 (N_6124,N_5203,N_5708);
nand U6125 (N_6125,N_4464,N_5281);
or U6126 (N_6126,N_4240,N_5942);
xnor U6127 (N_6127,N_4954,N_5140);
nor U6128 (N_6128,N_5862,N_4921);
xnor U6129 (N_6129,N_4569,N_4422);
nor U6130 (N_6130,N_4510,N_5939);
and U6131 (N_6131,N_5010,N_4610);
nand U6132 (N_6132,N_4413,N_4445);
and U6133 (N_6133,N_4886,N_5626);
and U6134 (N_6134,N_4625,N_4828);
and U6135 (N_6135,N_5162,N_4276);
xor U6136 (N_6136,N_4294,N_5873);
xor U6137 (N_6137,N_4461,N_5604);
nor U6138 (N_6138,N_4881,N_4563);
nor U6139 (N_6139,N_5113,N_5638);
nor U6140 (N_6140,N_4463,N_4967);
nand U6141 (N_6141,N_5237,N_4371);
or U6142 (N_6142,N_5431,N_4092);
or U6143 (N_6143,N_5716,N_5481);
nor U6144 (N_6144,N_5459,N_4796);
or U6145 (N_6145,N_4307,N_4643);
nor U6146 (N_6146,N_5852,N_4514);
xnor U6147 (N_6147,N_4133,N_4847);
nand U6148 (N_6148,N_4946,N_5532);
nand U6149 (N_6149,N_4073,N_5850);
nand U6150 (N_6150,N_5956,N_4382);
nor U6151 (N_6151,N_4741,N_5681);
nand U6152 (N_6152,N_5199,N_5061);
nand U6153 (N_6153,N_4854,N_5133);
nand U6154 (N_6154,N_5406,N_4430);
nand U6155 (N_6155,N_5337,N_4958);
nor U6156 (N_6156,N_5547,N_4309);
or U6157 (N_6157,N_5034,N_4649);
nor U6158 (N_6158,N_5141,N_5142);
nor U6159 (N_6159,N_4291,N_5072);
nor U6160 (N_6160,N_4587,N_5953);
nand U6161 (N_6161,N_4455,N_5720);
nand U6162 (N_6162,N_5663,N_5377);
nand U6163 (N_6163,N_4664,N_5837);
or U6164 (N_6164,N_4154,N_4674);
nand U6165 (N_6165,N_5538,N_5594);
and U6166 (N_6166,N_5065,N_4871);
nor U6167 (N_6167,N_5175,N_4485);
or U6168 (N_6168,N_4069,N_5692);
and U6169 (N_6169,N_5321,N_4590);
or U6170 (N_6170,N_5739,N_5925);
or U6171 (N_6171,N_5340,N_5938);
or U6172 (N_6172,N_5378,N_5348);
nor U6173 (N_6173,N_5083,N_5724);
nand U6174 (N_6174,N_4595,N_4217);
xor U6175 (N_6175,N_4059,N_5315);
nand U6176 (N_6176,N_4960,N_5783);
xor U6177 (N_6177,N_4364,N_4384);
and U6178 (N_6178,N_5844,N_5973);
and U6179 (N_6179,N_5610,N_4840);
or U6180 (N_6180,N_4861,N_4718);
nand U6181 (N_6181,N_4834,N_5931);
nand U6182 (N_6182,N_5020,N_4869);
nand U6183 (N_6183,N_4301,N_5801);
nor U6184 (N_6184,N_5564,N_5241);
nand U6185 (N_6185,N_5795,N_4502);
xor U6186 (N_6186,N_4103,N_5996);
nor U6187 (N_6187,N_4254,N_4325);
nand U6188 (N_6188,N_4047,N_4877);
and U6189 (N_6189,N_4265,N_5168);
xor U6190 (N_6190,N_4475,N_5401);
and U6191 (N_6191,N_5549,N_4672);
xnor U6192 (N_6192,N_5280,N_5958);
xnor U6193 (N_6193,N_5462,N_5255);
and U6194 (N_6194,N_5200,N_4581);
and U6195 (N_6195,N_5802,N_5620);
nand U6196 (N_6196,N_4665,N_5725);
and U6197 (N_6197,N_5840,N_5275);
nor U6198 (N_6198,N_4585,N_5123);
nand U6199 (N_6199,N_4100,N_5164);
and U6200 (N_6200,N_4617,N_4067);
xor U6201 (N_6201,N_5407,N_4078);
xor U6202 (N_6202,N_4311,N_5539);
nor U6203 (N_6203,N_4096,N_4101);
or U6204 (N_6204,N_4063,N_5972);
xor U6205 (N_6205,N_5360,N_5223);
xnor U6206 (N_6206,N_5985,N_4119);
nand U6207 (N_6207,N_4839,N_4490);
nor U6208 (N_6208,N_4170,N_4907);
and U6209 (N_6209,N_4996,N_5119);
nand U6210 (N_6210,N_5296,N_4407);
nand U6211 (N_6211,N_4622,N_4833);
nor U6212 (N_6212,N_5201,N_4774);
or U6213 (N_6213,N_5861,N_4509);
nor U6214 (N_6214,N_4166,N_4759);
and U6215 (N_6215,N_4763,N_5530);
and U6216 (N_6216,N_5293,N_5552);
xnor U6217 (N_6217,N_4795,N_5859);
and U6218 (N_6218,N_5219,N_4990);
nand U6219 (N_6219,N_4478,N_5190);
xor U6220 (N_6220,N_4879,N_4630);
nor U6221 (N_6221,N_4670,N_4650);
nor U6222 (N_6222,N_5121,N_4880);
nand U6223 (N_6223,N_4470,N_5232);
nand U6224 (N_6224,N_4456,N_4201);
nand U6225 (N_6225,N_4271,N_5857);
xnor U6226 (N_6226,N_4159,N_5863);
or U6227 (N_6227,N_5039,N_4127);
or U6228 (N_6228,N_4066,N_4976);
xnor U6229 (N_6229,N_4586,N_5440);
xnor U6230 (N_6230,N_4565,N_4488);
or U6231 (N_6231,N_5450,N_4431);
and U6232 (N_6232,N_5242,N_5076);
nand U6233 (N_6233,N_4721,N_5019);
nor U6234 (N_6234,N_5316,N_5374);
nand U6235 (N_6235,N_4980,N_4746);
xor U6236 (N_6236,N_5687,N_5915);
nand U6237 (N_6237,N_5271,N_4762);
and U6238 (N_6238,N_4028,N_4076);
nor U6239 (N_6239,N_5025,N_5409);
or U6240 (N_6240,N_4444,N_4052);
nor U6241 (N_6241,N_4349,N_4760);
or U6242 (N_6242,N_5016,N_4940);
or U6243 (N_6243,N_4711,N_5534);
nor U6244 (N_6244,N_5144,N_5457);
nor U6245 (N_6245,N_5602,N_4038);
or U6246 (N_6246,N_5900,N_5088);
or U6247 (N_6247,N_4298,N_5525);
or U6248 (N_6248,N_4064,N_4360);
or U6249 (N_6249,N_4520,N_5031);
or U6250 (N_6250,N_5864,N_4503);
nor U6251 (N_6251,N_5731,N_5359);
or U6252 (N_6252,N_4511,N_5427);
nor U6253 (N_6253,N_4604,N_4710);
nand U6254 (N_6254,N_5328,N_5839);
nor U6255 (N_6255,N_4831,N_5490);
and U6256 (N_6256,N_4767,N_5299);
nand U6257 (N_6257,N_4468,N_4324);
nor U6258 (N_6258,N_5623,N_4882);
xnor U6259 (N_6259,N_5913,N_5078);
and U6260 (N_6260,N_5656,N_4068);
nor U6261 (N_6261,N_4177,N_5176);
nor U6262 (N_6262,N_5258,N_5765);
nand U6263 (N_6263,N_4607,N_4156);
xnor U6264 (N_6264,N_5584,N_5499);
nor U6265 (N_6265,N_5624,N_4115);
xnor U6266 (N_6266,N_5485,N_4300);
or U6267 (N_6267,N_4788,N_5510);
nand U6268 (N_6268,N_4576,N_4228);
and U6269 (N_6269,N_5609,N_4986);
nor U6270 (N_6270,N_4806,N_4167);
xnor U6271 (N_6271,N_5588,N_4369);
or U6272 (N_6272,N_4623,N_5331);
and U6273 (N_6273,N_5898,N_4326);
xor U6274 (N_6274,N_4013,N_5714);
or U6275 (N_6275,N_5570,N_4124);
xor U6276 (N_6276,N_4184,N_5138);
nand U6277 (N_6277,N_4668,N_4978);
xnor U6278 (N_6278,N_5811,N_4974);
nand U6279 (N_6279,N_4062,N_4698);
and U6280 (N_6280,N_4658,N_5488);
and U6281 (N_6281,N_4805,N_5353);
nor U6282 (N_6282,N_4268,N_4913);
xnor U6283 (N_6283,N_5040,N_4352);
xor U6284 (N_6284,N_4448,N_5382);
nand U6285 (N_6285,N_4341,N_5158);
xor U6286 (N_6286,N_4053,N_4329);
and U6287 (N_6287,N_5848,N_5622);
nor U6288 (N_6288,N_5778,N_5451);
nor U6289 (N_6289,N_5633,N_4036);
nor U6290 (N_6290,N_4594,N_5204);
xnor U6291 (N_6291,N_4009,N_5880);
or U6292 (N_6292,N_5800,N_5887);
xnor U6293 (N_6293,N_5476,N_5289);
and U6294 (N_6294,N_4357,N_5772);
nor U6295 (N_6295,N_5193,N_4952);
xor U6296 (N_6296,N_4497,N_4972);
nand U6297 (N_6297,N_5924,N_5650);
and U6298 (N_6298,N_4346,N_4479);
and U6299 (N_6299,N_4895,N_4056);
or U6300 (N_6300,N_5388,N_4460);
nor U6301 (N_6301,N_4406,N_4819);
xnor U6302 (N_6302,N_4773,N_4602);
or U6303 (N_6303,N_5028,N_4350);
and U6304 (N_6304,N_4532,N_4614);
nand U6305 (N_6305,N_5841,N_4543);
xor U6306 (N_6306,N_4176,N_4285);
or U6307 (N_6307,N_4424,N_5433);
nor U6308 (N_6308,N_4771,N_4809);
or U6309 (N_6309,N_4112,N_4797);
or U6310 (N_6310,N_5208,N_5198);
xor U6311 (N_6311,N_4838,N_5734);
or U6312 (N_6312,N_4012,N_5757);
xnor U6313 (N_6313,N_4225,N_4466);
xnor U6314 (N_6314,N_5128,N_4434);
nand U6315 (N_6315,N_5046,N_5933);
nand U6316 (N_6316,N_5254,N_4322);
nand U6317 (N_6317,N_4130,N_4368);
nand U6318 (N_6318,N_4558,N_5310);
or U6319 (N_6319,N_4070,N_5312);
and U6320 (N_6320,N_4690,N_4930);
nor U6321 (N_6321,N_4142,N_4042);
nor U6322 (N_6322,N_4683,N_5167);
nand U6323 (N_6323,N_4724,N_4403);
and U6324 (N_6324,N_5690,N_5415);
nand U6325 (N_6325,N_4527,N_4450);
and U6326 (N_6326,N_5675,N_4661);
nand U6327 (N_6327,N_4016,N_4637);
nand U6328 (N_6328,N_4535,N_5268);
xnor U6329 (N_6329,N_4253,N_5540);
nor U6330 (N_6330,N_5101,N_5474);
nand U6331 (N_6331,N_4259,N_4523);
nor U6332 (N_6332,N_4014,N_4121);
nand U6333 (N_6333,N_5166,N_4550);
and U6334 (N_6334,N_4187,N_5507);
xnor U6335 (N_6335,N_5600,N_4752);
or U6336 (N_6336,N_4385,N_4775);
xor U6337 (N_6337,N_5053,N_4515);
and U6338 (N_6338,N_5551,N_5644);
nor U6339 (N_6339,N_4920,N_4568);
xor U6340 (N_6340,N_5789,N_4089);
xnor U6341 (N_6341,N_4733,N_5477);
and U6342 (N_6342,N_4084,N_5084);
nand U6343 (N_6343,N_5723,N_4269);
nand U6344 (N_6344,N_4123,N_5194);
nand U6345 (N_6345,N_5393,N_5642);
or U6346 (N_6346,N_5390,N_4079);
xnor U6347 (N_6347,N_4634,N_4388);
nand U6348 (N_6348,N_4693,N_4947);
and U6349 (N_6349,N_4236,N_5195);
and U6350 (N_6350,N_4147,N_4397);
or U6351 (N_6351,N_5444,N_5590);
or U6352 (N_6352,N_5758,N_4010);
xor U6353 (N_6353,N_4919,N_5151);
nor U6354 (N_6354,N_5736,N_5799);
xnor U6355 (N_6355,N_5541,N_5986);
and U6356 (N_6356,N_4218,N_4608);
and U6357 (N_6357,N_4885,N_5773);
nand U6358 (N_6358,N_4692,N_5881);
or U6359 (N_6359,N_5641,N_5580);
nor U6360 (N_6360,N_5361,N_4438);
xor U6361 (N_6361,N_5919,N_5471);
nand U6362 (N_6362,N_5911,N_4802);
and U6363 (N_6363,N_5523,N_4297);
and U6364 (N_6364,N_5914,N_5071);
nand U6365 (N_6365,N_5577,N_4283);
xnor U6366 (N_6366,N_4017,N_4148);
nand U6367 (N_6367,N_4501,N_4332);
xnor U6368 (N_6368,N_5420,N_4564);
nor U6369 (N_6369,N_4874,N_4004);
and U6370 (N_6370,N_4723,N_5099);
and U6371 (N_6371,N_5821,N_4365);
nor U6372 (N_6372,N_5120,N_4286);
xnor U6373 (N_6373,N_5106,N_5759);
or U6374 (N_6374,N_5188,N_4541);
nor U6375 (N_6375,N_5601,N_4657);
or U6376 (N_6376,N_5404,N_5182);
xor U6377 (N_6377,N_5849,N_4971);
or U6378 (N_6378,N_4599,N_5035);
nand U6379 (N_6379,N_5715,N_5793);
nand U6380 (N_6380,N_5702,N_5032);
or U6381 (N_6381,N_4779,N_4086);
nand U6382 (N_6382,N_4561,N_4196);
nor U6383 (N_6383,N_4932,N_4132);
or U6384 (N_6384,N_4419,N_5603);
and U6385 (N_6385,N_4720,N_4975);
nand U6386 (N_6386,N_4486,N_5569);
nand U6387 (N_6387,N_5227,N_5472);
xor U6388 (N_6388,N_4270,N_5077);
xnor U6389 (N_6389,N_5782,N_5389);
xor U6390 (N_6390,N_5465,N_4031);
or U6391 (N_6391,N_4660,N_4669);
nand U6392 (N_6392,N_4798,N_4621);
and U6393 (N_6393,N_4749,N_5748);
xor U6394 (N_6394,N_4453,N_5960);
nand U6395 (N_6395,N_5171,N_5812);
or U6396 (N_6396,N_4030,N_4731);
or U6397 (N_6397,N_5467,N_4629);
and U6398 (N_6398,N_4308,N_5717);
or U6399 (N_6399,N_5598,N_5805);
or U6400 (N_6400,N_5090,N_5308);
and U6401 (N_6401,N_5829,N_5058);
and U6402 (N_6402,N_4417,N_4810);
or U6403 (N_6403,N_5828,N_4367);
nor U6404 (N_6404,N_4530,N_5879);
or U6405 (N_6405,N_4246,N_5545);
or U6406 (N_6406,N_5410,N_4489);
nand U6407 (N_6407,N_5830,N_4612);
xor U6408 (N_6408,N_4973,N_5386);
nor U6409 (N_6409,N_4405,N_4712);
xnor U6410 (N_6410,N_4241,N_4785);
nand U6411 (N_6411,N_5876,N_4605);
nor U6412 (N_6412,N_5946,N_5347);
and U6413 (N_6413,N_5326,N_4647);
nand U6414 (N_6414,N_4203,N_4579);
or U6415 (N_6415,N_5413,N_5356);
nor U6416 (N_6416,N_4686,N_5082);
xor U6417 (N_6417,N_5657,N_5583);
xnor U6418 (N_6418,N_4209,N_5423);
xor U6419 (N_6419,N_4953,N_5033);
nand U6420 (N_6420,N_4548,N_4339);
and U6421 (N_6421,N_5174,N_4116);
nor U6422 (N_6422,N_5582,N_5694);
xor U6423 (N_6423,N_5334,N_5568);
or U6424 (N_6424,N_5085,N_4811);
nor U6425 (N_6425,N_4462,N_5335);
xor U6426 (N_6426,N_5679,N_4955);
xnor U6427 (N_6427,N_4340,N_5907);
and U6428 (N_6428,N_5877,N_4687);
nor U6429 (N_6429,N_4615,N_4813);
nor U6430 (N_6430,N_5612,N_4772);
xor U6431 (N_6431,N_5630,N_5136);
nand U6432 (N_6432,N_5395,N_4135);
xor U6433 (N_6433,N_4870,N_4451);
or U6434 (N_6434,N_4512,N_5235);
nor U6435 (N_6435,N_4896,N_5210);
xor U6436 (N_6436,N_4374,N_4164);
nand U6437 (N_6437,N_4743,N_5069);
nor U6438 (N_6438,N_5963,N_4786);
and U6439 (N_6439,N_5822,N_4559);
nor U6440 (N_6440,N_4105,N_5908);
nor U6441 (N_6441,N_4632,N_5283);
or U6442 (N_6442,N_5381,N_5921);
xor U6443 (N_6443,N_4855,N_4125);
nand U6444 (N_6444,N_4452,N_4446);
nor U6445 (N_6445,N_4578,N_4945);
xnor U6446 (N_6446,N_5780,N_5284);
or U6447 (N_6447,N_4215,N_5196);
xnor U6448 (N_6448,N_5729,N_4765);
and U6449 (N_6449,N_5355,N_5441);
nand U6450 (N_6450,N_5697,N_5464);
xor U6451 (N_6451,N_5376,N_5408);
xnor U6452 (N_6452,N_5804,N_4513);
or U6453 (N_6453,N_5169,N_4824);
nor U6454 (N_6454,N_4727,N_4526);
nand U6455 (N_6455,N_4700,N_5250);
nor U6456 (N_6456,N_4636,N_5737);
and U6457 (N_6457,N_5767,N_5505);
nor U6458 (N_6458,N_5969,N_4904);
or U6459 (N_6459,N_4926,N_5248);
and U6460 (N_6460,N_4626,N_4923);
xnor U6461 (N_6461,N_4747,N_5785);
and U6462 (N_6462,N_4910,N_4715);
or U6463 (N_6463,N_5131,N_4709);
nand U6464 (N_6464,N_4000,N_5665);
nor U6465 (N_6465,N_4094,N_5305);
nand U6466 (N_6466,N_4645,N_5678);
nand U6467 (N_6467,N_5992,N_5947);
xnor U6468 (N_6468,N_4051,N_4682);
nand U6469 (N_6469,N_5669,N_5741);
or U6470 (N_6470,N_4314,N_5556);
nand U6471 (N_6471,N_5005,N_5469);
nand U6472 (N_6472,N_5515,N_4571);
nor U6473 (N_6473,N_5302,N_5202);
xor U6474 (N_6474,N_5860,N_4293);
nor U6475 (N_6475,N_5068,N_5930);
or U6476 (N_6476,N_5266,N_5798);
or U6477 (N_6477,N_4032,N_5984);
or U6478 (N_6478,N_5187,N_4803);
nor U6479 (N_6479,N_5991,N_4480);
xor U6480 (N_6480,N_4931,N_4963);
nand U6481 (N_6481,N_5553,N_4408);
nor U6482 (N_6482,N_5749,N_5836);
nor U6483 (N_6483,N_4126,N_5683);
or U6484 (N_6484,N_4889,N_4495);
nand U6485 (N_6485,N_4140,N_4107);
xnor U6486 (N_6486,N_4057,N_5192);
or U6487 (N_6487,N_4024,N_4172);
or U6488 (N_6488,N_4699,N_4190);
nor U6489 (N_6489,N_4162,N_5894);
nand U6490 (N_6490,N_5064,N_5156);
nand U6491 (N_6491,N_4529,N_4151);
and U6492 (N_6492,N_5180,N_5866);
nor U6493 (N_6493,N_5978,N_5659);
or U6494 (N_6494,N_4420,N_4620);
xnor U6495 (N_6495,N_4908,N_4335);
or U6496 (N_6496,N_4194,N_4165);
nor U6497 (N_6497,N_4929,N_5596);
xnor U6498 (N_6498,N_5605,N_4160);
xor U6499 (N_6499,N_5059,N_5854);
or U6500 (N_6500,N_4860,N_5157);
and U6501 (N_6501,N_4905,N_4542);
xnor U6502 (N_6502,N_5259,N_5502);
and U6503 (N_6503,N_5496,N_5475);
xor U6504 (N_6504,N_4363,N_4593);
nand U6505 (N_6505,N_5339,N_5089);
xor U6506 (N_6506,N_4757,N_5412);
xnor U6507 (N_6507,N_5118,N_5685);
or U6508 (N_6508,N_4536,N_5814);
nand U6509 (N_6509,N_5392,N_4481);
nor U6510 (N_6510,N_5587,N_5566);
and U6511 (N_6511,N_4278,N_5062);
or U6512 (N_6512,N_5267,N_5575);
xor U6513 (N_6513,N_5216,N_5170);
or U6514 (N_6514,N_4428,N_4288);
nor U6515 (N_6515,N_5230,N_4628);
xor U6516 (N_6516,N_5021,N_5455);
nand U6517 (N_6517,N_5796,N_4386);
nand U6518 (N_6518,N_4557,N_5265);
nor U6519 (N_6519,N_5333,N_5442);
and U6520 (N_6520,N_5516,N_4492);
nor U6521 (N_6521,N_5585,N_5686);
and U6522 (N_6522,N_5784,N_5043);
xor U6523 (N_6523,N_4734,N_5827);
and U6524 (N_6524,N_4936,N_4229);
nor U6525 (N_6525,N_5173,N_4022);
and U6526 (N_6526,N_5856,N_5205);
and U6527 (N_6527,N_4618,N_4742);
nand U6528 (N_6528,N_4168,N_5178);
nor U6529 (N_6529,N_5819,N_4890);
and U6530 (N_6530,N_5048,N_4783);
nand U6531 (N_6531,N_5012,N_5292);
nand U6532 (N_6532,N_4750,N_4186);
nand U6533 (N_6533,N_5369,N_4867);
nor U6534 (N_6534,N_5497,N_4212);
nor U6535 (N_6535,N_5029,N_5695);
and U6536 (N_6536,N_4609,N_4292);
nand U6537 (N_6537,N_5365,N_4853);
xor U6538 (N_6538,N_4318,N_5649);
and U6539 (N_6539,N_5260,N_5400);
or U6540 (N_6540,N_4496,N_5269);
or U6541 (N_6541,N_5593,N_5352);
and U6542 (N_6542,N_4872,N_5186);
nor U6543 (N_6543,N_4782,N_4827);
and U6544 (N_6544,N_4355,N_5222);
nand U6545 (N_6545,N_4415,N_4573);
nor U6546 (N_6546,N_4849,N_4095);
xor U6547 (N_6547,N_5057,N_5177);
or U6548 (N_6548,N_5705,N_4816);
xor U6549 (N_6549,N_5661,N_5146);
or U6550 (N_6550,N_5820,N_5671);
nand U6551 (N_6551,N_4145,N_4380);
xor U6552 (N_6552,N_4429,N_4898);
nor U6553 (N_6553,N_4745,N_5648);
nor U6554 (N_6554,N_4396,N_5249);
nand U6555 (N_6555,N_4442,N_4235);
xor U6556 (N_6556,N_5226,N_4862);
xor U6557 (N_6557,N_5912,N_4021);
xor U6558 (N_6558,N_5943,N_5161);
nor U6559 (N_6559,N_5247,N_4373);
nand U6560 (N_6560,N_4673,N_4987);
nand U6561 (N_6561,N_5508,N_4231);
nor U6562 (N_6562,N_5832,N_5742);
nand U6563 (N_6563,N_4321,N_5940);
or U6564 (N_6564,N_5917,N_5207);
or U6565 (N_6565,N_5478,N_5135);
nor U6566 (N_6566,N_5892,N_5752);
xor U6567 (N_6567,N_5015,N_5562);
nor U6568 (N_6568,N_5243,N_5923);
xor U6569 (N_6569,N_4815,N_4970);
nor U6570 (N_6570,N_4029,N_5493);
or U6571 (N_6571,N_5372,N_5454);
or U6572 (N_6572,N_4997,N_5883);
nor U6573 (N_6573,N_4120,N_4640);
nor U6574 (N_6574,N_4065,N_5961);
and U6575 (N_6575,N_5183,N_5037);
nor U6576 (N_6576,N_4546,N_5527);
nor U6577 (N_6577,N_4304,N_4441);
or U6578 (N_6578,N_4678,N_5346);
nand U6579 (N_6579,N_4830,N_5461);
nand U6580 (N_6580,N_4185,N_5636);
xnor U6581 (N_6581,N_5700,N_4226);
or U6582 (N_6582,N_5264,N_5052);
or U6583 (N_6583,N_4054,N_5619);
or U6584 (N_6584,N_4887,N_4846);
xnor U6585 (N_6585,N_4751,N_5009);
or U6586 (N_6586,N_4398,N_4644);
nor U6587 (N_6587,N_4726,N_4391);
or U6588 (N_6588,N_4345,N_5764);
xor U6589 (N_6589,N_4655,N_5647);
nand U6590 (N_6590,N_5774,N_4188);
and U6591 (N_6591,N_5179,N_4804);
or U6592 (N_6592,N_5416,N_5093);
nand U6593 (N_6593,N_4208,N_4498);
nor U6594 (N_6594,N_5405,N_4211);
nand U6595 (N_6595,N_5835,N_5330);
and U6596 (N_6596,N_4728,N_4764);
xor U6597 (N_6597,N_4676,N_4714);
nand U6598 (N_6598,N_4588,N_5834);
and U6599 (N_6599,N_5422,N_4969);
nor U6600 (N_6600,N_4006,N_5419);
nand U6601 (N_6601,N_5214,N_4968);
xnor U6602 (N_6602,N_4716,N_5414);
nand U6603 (N_6603,N_4989,N_5965);
nand U6604 (N_6604,N_5149,N_5038);
or U6605 (N_6605,N_4344,N_4928);
nand U6606 (N_6606,N_5797,N_4560);
xnor U6607 (N_6607,N_4487,N_5129);
nor U6608 (N_6608,N_5542,N_4290);
nor U6609 (N_6609,N_4110,N_4171);
nand U6610 (N_6610,N_5066,N_4252);
or U6611 (N_6611,N_4136,N_4310);
or U6612 (N_6612,N_5263,N_5329);
nand U6613 (N_6613,N_4090,N_4949);
nand U6614 (N_6614,N_4822,N_4210);
and U6615 (N_6615,N_5003,N_5777);
nand U6616 (N_6616,N_4493,N_4873);
and U6617 (N_6617,N_4808,N_4893);
or U6618 (N_6618,N_4891,N_5086);
nor U6619 (N_6619,N_4275,N_5831);
xor U6620 (N_6620,N_4814,N_4580);
and U6621 (N_6621,N_5816,N_5535);
xnor U6622 (N_6622,N_4917,N_4641);
or U6623 (N_6623,N_4688,N_5890);
nor U6624 (N_6624,N_5635,N_5998);
or U6625 (N_6625,N_4122,N_5060);
and U6626 (N_6626,N_4848,N_5824);
nand U6627 (N_6627,N_4506,N_4099);
nor U6628 (N_6628,N_4048,N_5261);
nor U6629 (N_6629,N_5270,N_4260);
and U6630 (N_6630,N_4394,N_5870);
xor U6631 (N_6631,N_4793,N_5049);
and U6632 (N_6632,N_4230,N_5935);
or U6633 (N_6633,N_4237,N_5761);
or U6634 (N_6634,N_5092,N_5768);
nand U6635 (N_6635,N_5974,N_4060);
and U6636 (N_6636,N_5122,N_4256);
xnor U6637 (N_6637,N_5980,N_4912);
or U6638 (N_6638,N_4961,N_4412);
or U6639 (N_6639,N_4525,N_4702);
and U6640 (N_6640,N_5109,N_4018);
or U6641 (N_6641,N_4689,N_5806);
nand U6642 (N_6642,N_5521,N_4473);
nor U6643 (N_6643,N_5501,N_4856);
nor U6644 (N_6644,N_4982,N_5239);
nor U6645 (N_6645,N_4411,N_5234);
nor U6646 (N_6646,N_5397,N_5664);
or U6647 (N_6647,N_4372,N_5285);
or U6648 (N_6648,N_4744,N_4705);
or U6649 (N_6649,N_4534,N_5721);
xnor U6650 (N_6650,N_5906,N_4439);
xor U6651 (N_6651,N_4315,N_4888);
or U6652 (N_6652,N_4538,N_4251);
and U6653 (N_6653,N_4414,N_4823);
xnor U6654 (N_6654,N_5660,N_4058);
and U6655 (N_6655,N_4337,N_5236);
nor U6656 (N_6656,N_5703,N_5290);
or U6657 (N_6657,N_5081,N_4979);
and U6658 (N_6658,N_4426,N_4909);
and U6659 (N_6659,N_5989,N_4331);
nor U6660 (N_6660,N_5287,N_4280);
or U6661 (N_6661,N_5006,N_5555);
nand U6662 (N_6662,N_4336,N_4317);
nand U6663 (N_6663,N_4071,N_4375);
and U6664 (N_6664,N_4654,N_4736);
and U6665 (N_6665,N_5786,N_5448);
nor U6666 (N_6666,N_4966,N_5680);
or U6667 (N_6667,N_5253,N_5815);
or U6668 (N_6668,N_4704,N_5853);
nor U6669 (N_6669,N_4540,N_4423);
xnor U6670 (N_6670,N_4787,N_5755);
nand U6671 (N_6671,N_5617,N_4249);
and U6672 (N_6672,N_5327,N_4984);
or U6673 (N_6673,N_4662,N_5878);
and U6674 (N_6674,N_4379,N_5160);
xor U6675 (N_6675,N_4792,N_5114);
nand U6676 (N_6676,N_4200,N_5398);
xnor U6677 (N_6677,N_4566,N_5572);
nand U6678 (N_6678,N_4570,N_4934);
xnor U6679 (N_6679,N_5338,N_4624);
or U6680 (N_6680,N_5282,N_5674);
xnor U6681 (N_6681,N_5567,N_5418);
nand U6682 (N_6682,N_5771,N_5738);
or U6683 (N_6683,N_5874,N_4433);
and U6684 (N_6684,N_5368,N_5826);
nor U6685 (N_6685,N_5067,N_4378);
nand U6686 (N_6686,N_4255,N_4131);
nor U6687 (N_6687,N_4238,N_4469);
nor U6688 (N_6688,N_5495,N_4901);
and U6689 (N_6689,N_5385,N_5181);
nor U6690 (N_6690,N_4264,N_5273);
nand U6691 (N_6691,N_4801,N_5888);
nor U6692 (N_6692,N_5323,N_5673);
xnor U6693 (N_6693,N_4220,N_4659);
and U6694 (N_6694,N_5350,N_5576);
nor U6695 (N_6695,N_5528,N_5148);
nor U6696 (N_6696,N_4875,N_5482);
and U6697 (N_6697,N_5753,N_5903);
xnor U6698 (N_6698,N_5544,N_5150);
nor U6699 (N_6699,N_4852,N_4596);
or U6700 (N_6700,N_5145,N_4927);
and U6701 (N_6701,N_5364,N_5317);
and U6702 (N_6702,N_4531,N_5865);
and U6703 (N_6703,N_5833,N_4761);
nand U6704 (N_6704,N_4178,N_4007);
nand U6705 (N_6705,N_4584,N_5301);
or U6706 (N_6706,N_5134,N_4524);
or U6707 (N_6707,N_4505,N_5718);
and U6708 (N_6708,N_4778,N_4508);
or U6709 (N_6709,N_4083,N_5051);
and U6710 (N_6710,N_4799,N_5432);
or U6711 (N_6711,N_5104,N_4242);
nor U6712 (N_6712,N_5054,N_4108);
nand U6713 (N_6713,N_5948,N_4404);
xor U6714 (N_6714,N_4395,N_5847);
and U6715 (N_6715,N_5045,N_4416);
and U6716 (N_6716,N_4500,N_5102);
xnor U6717 (N_6717,N_4735,N_4868);
or U6718 (N_6718,N_5080,N_4663);
nand U6719 (N_6719,N_5698,N_5108);
nand U6720 (N_6720,N_5779,N_4035);
or U6721 (N_6721,N_4935,N_4850);
and U6722 (N_6722,N_4437,N_5693);
nor U6723 (N_6723,N_4677,N_5909);
and U6724 (N_6724,N_4109,N_4305);
nand U6725 (N_6725,N_5047,N_5056);
nor U6726 (N_6726,N_5628,N_5561);
nor U6727 (N_6727,N_5875,N_4528);
xnor U6728 (N_6728,N_4163,N_4182);
xnor U6729 (N_6729,N_5970,N_5899);
nand U6730 (N_6730,N_5103,N_4939);
or U6731 (N_6731,N_4289,N_4195);
or U6732 (N_6732,N_5079,N_5845);
and U6733 (N_6733,N_4082,N_4574);
nand U6734 (N_6734,N_5117,N_5319);
xnor U6735 (N_6735,N_5375,N_5402);
nand U6736 (N_6736,N_4995,N_4224);
nor U6737 (N_6737,N_4227,N_4717);
nor U6738 (N_6738,N_5885,N_4981);
and U6739 (N_6739,N_5858,N_4521);
or U6740 (N_6740,N_4098,N_4627);
and U6741 (N_6741,N_5211,N_5954);
nand U6742 (N_6742,N_5341,N_4983);
nand U6743 (N_6743,N_5172,N_4467);
nor U6744 (N_6744,N_4204,N_5309);
nand U6745 (N_6745,N_5426,N_4213);
nor U6746 (N_6746,N_5163,N_5522);
nor U6747 (N_6747,N_5391,N_4435);
or U6748 (N_6748,N_5524,N_5949);
nor U6749 (N_6749,N_4033,N_4351);
and U6750 (N_6750,N_5286,N_4299);
nand U6751 (N_6751,N_4998,N_4008);
and U6752 (N_6752,N_5345,N_4440);
nor U6753 (N_6753,N_4088,N_5983);
or U6754 (N_6754,N_5677,N_5443);
xnor U6755 (N_6755,N_5897,N_4222);
or U6756 (N_6756,N_5436,N_4471);
xor U6757 (N_6757,N_5318,N_4039);
nand U6758 (N_6758,N_5513,N_5143);
and U6759 (N_6759,N_5244,N_4756);
and U6760 (N_6760,N_5362,N_4192);
or U6761 (N_6761,N_5518,N_5449);
and U6762 (N_6762,N_4754,N_5645);
nand U6763 (N_6763,N_5322,N_5565);
and U6764 (N_6764,N_5277,N_4876);
nor U6765 (N_6765,N_5613,N_5306);
nand U6766 (N_6766,N_5396,N_4482);
nand U6767 (N_6767,N_5197,N_4841);
xnor U6768 (N_6768,N_5891,N_5982);
nand U6769 (N_6769,N_4472,N_4685);
or U6770 (N_6770,N_4730,N_4858);
nand U6771 (N_6771,N_5517,N_5351);
nor U6772 (N_6772,N_5344,N_4050);
nand U6773 (N_6773,N_5662,N_5229);
nor U6774 (N_6774,N_4679,N_5479);
and U6775 (N_6775,N_4306,N_5434);
or U6776 (N_6776,N_5869,N_4043);
and U6777 (N_6777,N_5592,N_4302);
or U6778 (N_6778,N_4019,N_5838);
nor U6779 (N_6779,N_4902,N_5473);
or U6780 (N_6780,N_4328,N_4758);
and U6781 (N_6781,N_5842,N_5766);
nand U6782 (N_6782,N_4780,N_5668);
nor U6783 (N_6783,N_5955,N_4504);
or U6784 (N_6784,N_5579,N_4567);
and U6785 (N_6785,N_5851,N_5256);
xor U6786 (N_6786,N_4951,N_5294);
nand U6787 (N_6787,N_4274,N_5231);
or U6788 (N_6788,N_4002,N_4001);
nand U6789 (N_6789,N_4924,N_4706);
nor U6790 (N_6790,N_4358,N_4857);
and U6791 (N_6791,N_4737,N_4638);
nor U6792 (N_6792,N_5466,N_5105);
and U6793 (N_6793,N_4549,N_5615);
nand U6794 (N_6794,N_5491,N_4725);
xnor U6795 (N_6795,N_5926,N_4791);
nand U6796 (N_6796,N_4937,N_4418);
nand U6797 (N_6797,N_5095,N_5159);
xor U6798 (N_6798,N_4755,N_5453);
xor U6799 (N_6799,N_4102,N_4533);
nor U6800 (N_6800,N_4359,N_5483);
xor U6801 (N_6801,N_4362,N_4117);
and U6802 (N_6802,N_5722,N_4781);
or U6803 (N_6803,N_5438,N_4183);
or U6804 (N_6804,N_4589,N_5127);
xor U6805 (N_6805,N_5910,N_4077);
nand U6806 (N_6806,N_4393,N_5559);
nand U6807 (N_6807,N_4944,N_4366);
and U6808 (N_6808,N_5042,N_4261);
nand U6809 (N_6809,N_5945,N_5094);
nand U6810 (N_6810,N_4377,N_4207);
nand U6811 (N_6811,N_4807,N_4800);
nor U6812 (N_6812,N_5747,N_5008);
nor U6813 (N_6813,N_5629,N_4667);
and U6814 (N_6814,N_4897,N_5537);
xnor U6815 (N_6815,N_4049,N_5684);
nor U6816 (N_6816,N_4267,N_5987);
nand U6817 (N_6817,N_5756,N_5489);
nand U6818 (N_6818,N_4499,N_4266);
or U6819 (N_6819,N_4826,N_5509);
nand U6820 (N_6820,N_4248,N_4545);
and U6821 (N_6821,N_5704,N_4221);
and U6822 (N_6822,N_4219,N_5548);
nor U6823 (N_6823,N_5809,N_4436);
nor U6824 (N_6824,N_5712,N_4864);
and U6825 (N_6825,N_4600,N_5578);
nand U6826 (N_6826,N_5927,N_5571);
and U6827 (N_6827,N_5733,N_5546);
and U6828 (N_6828,N_5994,N_5504);
or U6829 (N_6829,N_5599,N_5606);
nand U6830 (N_6830,N_5300,N_4284);
xnor U6831 (N_6831,N_4258,N_4648);
nand U6832 (N_6832,N_5618,N_4619);
nand U6833 (N_6833,N_4592,N_4138);
xnor U6834 (N_6834,N_5643,N_5279);
xor U6835 (N_6835,N_4128,N_4606);
nor U6836 (N_6836,N_5689,N_5116);
or U6837 (N_6837,N_5990,N_5932);
xor U6838 (N_6838,N_4633,N_5480);
or U6839 (N_6839,N_5027,N_5916);
nor U6840 (N_6840,N_4330,N_5550);
and U6841 (N_6841,N_4770,N_4922);
nand U6842 (N_6842,N_5670,N_4233);
xnor U6843 (N_6843,N_5366,N_5882);
xor U6844 (N_6844,N_4106,N_4465);
or U6845 (N_6845,N_5500,N_4263);
or U6846 (N_6846,N_5977,N_5735);
or U6847 (N_6847,N_5276,N_5614);
nor U6848 (N_6848,N_4962,N_4157);
nor U6849 (N_6849,N_4878,N_4348);
nand U6850 (N_6850,N_4173,N_4769);
and U6851 (N_6851,N_4859,N_4320);
xnor U6852 (N_6852,N_4691,N_4370);
nor U6853 (N_6853,N_4143,N_4957);
nand U6854 (N_6854,N_5968,N_5769);
and U6855 (N_6855,N_5278,N_5929);
xnor U6856 (N_6856,N_5574,N_5867);
nor U6857 (N_6857,N_4777,N_4198);
nor U6858 (N_6858,N_5775,N_4539);
and U6859 (N_6859,N_4087,N_5655);
xor U6860 (N_6860,N_4296,N_4832);
and U6861 (N_6861,N_5964,N_5367);
and U6862 (N_6862,N_4081,N_4400);
nand U6863 (N_6863,N_4011,N_5557);
nor U6864 (N_6864,N_5531,N_5740);
nand U6865 (N_6865,N_4845,N_4197);
xnor U6866 (N_6866,N_5130,N_4812);
xnor U6867 (N_6867,N_5417,N_4169);
or U6868 (N_6868,N_5586,N_5233);
and U6869 (N_6869,N_4516,N_4842);
nand U6870 (N_6870,N_5855,N_5132);
and U6871 (N_6871,N_4603,N_4993);
and U6872 (N_6872,N_5558,N_4273);
nand U6873 (N_6873,N_4794,N_5962);
or U6874 (N_6874,N_4577,N_5137);
nand U6875 (N_6875,N_4387,N_4675);
nand U6876 (N_6876,N_5097,N_4427);
nand U6877 (N_6877,N_5976,N_4137);
or U6878 (N_6878,N_5139,N_5936);
nand U6879 (N_6879,N_5760,N_5446);
xor U6880 (N_6880,N_4916,N_4883);
xor U6881 (N_6881,N_5995,N_4753);
nor U6882 (N_6882,N_4023,N_5790);
or U6883 (N_6883,N_5428,N_5125);
or U6884 (N_6884,N_5750,N_4045);
or U6885 (N_6885,N_5952,N_4537);
or U6886 (N_6886,N_5707,N_5295);
nand U6887 (N_6887,N_5399,N_5713);
and U6888 (N_6888,N_4948,N_4141);
and U6889 (N_6889,N_4181,N_5437);
and U6890 (N_6890,N_4055,N_5073);
nor U6891 (N_6891,N_5336,N_5825);
nor U6892 (N_6892,N_5526,N_4522);
xnor U6893 (N_6893,N_5637,N_4425);
or U6894 (N_6894,N_4666,N_5554);
xnor U6895 (N_6895,N_5631,N_5217);
or U6896 (N_6896,N_5658,N_5147);
or U6897 (N_6897,N_5000,N_4361);
or U6898 (N_6898,N_5063,N_4093);
or U6899 (N_6899,N_4432,N_5460);
xnor U6900 (N_6900,N_5999,N_5719);
or U6901 (N_6901,N_4313,N_4555);
or U6902 (N_6902,N_5993,N_4642);
xnor U6903 (N_6903,N_4316,N_5291);
nor U6904 (N_6904,N_4155,N_5153);
nor U6905 (N_6905,N_5950,N_4080);
nor U6906 (N_6906,N_5627,N_4020);
nand U6907 (N_6907,N_4243,N_4040);
or U6908 (N_6908,N_5298,N_4985);
and U6909 (N_6909,N_4517,N_4074);
nand U6910 (N_6910,N_5573,N_5044);
or U6911 (N_6911,N_5257,N_5871);
or U6912 (N_6912,N_4343,N_5506);
nand U6913 (N_6913,N_5154,N_5228);
or U6914 (N_6914,N_5240,N_5529);
nand U6915 (N_6915,N_5371,N_5314);
xnor U6916 (N_6916,N_5075,N_5699);
and U6917 (N_6917,N_4748,N_4037);
and U6918 (N_6918,N_4180,N_4992);
and U6919 (N_6919,N_5297,N_5781);
nor U6920 (N_6920,N_5763,N_4003);
nor U6921 (N_6921,N_5272,N_4825);
nor U6922 (N_6922,N_5246,N_4866);
xor U6923 (N_6923,N_5727,N_5220);
or U6924 (N_6924,N_4911,N_4449);
nand U6925 (N_6925,N_4146,N_4863);
xor U6926 (N_6926,N_5591,N_5893);
xnor U6927 (N_6927,N_5997,N_4601);
nand U6928 (N_6928,N_4111,N_4334);
nor U6929 (N_6929,N_5595,N_5810);
nand U6930 (N_6930,N_5934,N_5696);
or U6931 (N_6931,N_4965,N_4279);
nand U6932 (N_6932,N_5421,N_4113);
nor U6933 (N_6933,N_4199,N_4694);
nor U6934 (N_6934,N_5001,N_5494);
and U6935 (N_6935,N_4061,N_4977);
xor U6936 (N_6936,N_5324,N_5792);
xnor U6937 (N_6937,N_4988,N_5639);
and U6938 (N_6938,N_4631,N_4900);
or U6939 (N_6939,N_5445,N_4044);
nand U6940 (N_6940,N_5447,N_5191);
nor U6941 (N_6941,N_5967,N_5884);
nand U6942 (N_6942,N_4262,N_4611);
and U6943 (N_6943,N_4732,N_4232);
nand U6944 (N_6944,N_5794,N_5394);
nand U6945 (N_6945,N_5387,N_5070);
and U6946 (N_6946,N_5384,N_5951);
nand U6947 (N_6947,N_4696,N_5152);
nand U6948 (N_6948,N_5770,N_5251);
or U6949 (N_6949,N_5332,N_5411);
nand U6950 (N_6950,N_4484,N_4206);
nand U6951 (N_6951,N_5975,N_5026);
or U6952 (N_6952,N_4494,N_5634);
nand U6953 (N_6953,N_5487,N_5498);
xor U6954 (N_6954,N_4443,N_4401);
or U6955 (N_6955,N_4598,N_5024);
and U6956 (N_6956,N_5379,N_4202);
nor U6957 (N_6957,N_5342,N_5711);
or U6958 (N_6958,N_4915,N_5165);
and U6959 (N_6959,N_5607,N_5380);
nand U6960 (N_6960,N_5307,N_4959);
or U6961 (N_6961,N_4639,N_4257);
and U6962 (N_6962,N_5616,N_4829);
nor U6963 (N_6963,N_4713,N_5709);
nor U6964 (N_6964,N_5036,N_5966);
or U6965 (N_6965,N_5011,N_5155);
and U6966 (N_6966,N_4454,N_5843);
and U6967 (N_6967,N_4477,N_5288);
nor U6968 (N_6968,N_4161,N_5430);
nand U6969 (N_6969,N_4835,N_5895);
xnor U6970 (N_6970,N_4392,N_5667);
xor U6971 (N_6971,N_5110,N_4072);
xor U6972 (N_6972,N_5608,N_5808);
xor U6973 (N_6973,N_5560,N_5245);
nand U6974 (N_6974,N_5710,N_5621);
or U6975 (N_6975,N_5209,N_4843);
nor U6976 (N_6976,N_4483,N_4041);
or U6977 (N_6977,N_5435,N_5654);
or U6978 (N_6978,N_5354,N_5791);
and U6979 (N_6979,N_4097,N_4789);
or U6980 (N_6980,N_4554,N_5846);
or U6981 (N_6981,N_5672,N_4234);
or U6982 (N_6982,N_4075,N_4556);
and U6983 (N_6983,N_4410,N_5126);
nand U6984 (N_6984,N_5343,N_4635);
nand U6985 (N_6985,N_4026,N_4950);
nor U6986 (N_6986,N_5184,N_4381);
or U6987 (N_6987,N_4152,N_5221);
xor U6988 (N_6988,N_5728,N_5383);
and U6989 (N_6989,N_5520,N_5823);
and U6990 (N_6990,N_5303,N_5776);
or U6991 (N_6991,N_5004,N_5543);
nor U6992 (N_6992,N_4776,N_5252);
or U6993 (N_6993,N_5730,N_5439);
and U6994 (N_6994,N_5726,N_4719);
xor U6995 (N_6995,N_5597,N_5751);
xor U6996 (N_6996,N_5886,N_4118);
xnor U6997 (N_6997,N_5017,N_5458);
nand U6998 (N_6998,N_4653,N_4817);
xnor U6999 (N_6999,N_4790,N_4347);
nor U7000 (N_7000,N_5100,N_5967);
nand U7001 (N_7001,N_5650,N_4997);
or U7002 (N_7002,N_5142,N_4652);
nand U7003 (N_7003,N_4518,N_4986);
xor U7004 (N_7004,N_4889,N_4800);
or U7005 (N_7005,N_4745,N_5512);
xor U7006 (N_7006,N_5828,N_5795);
or U7007 (N_7007,N_4943,N_4620);
xor U7008 (N_7008,N_5543,N_4335);
nand U7009 (N_7009,N_5603,N_4269);
and U7010 (N_7010,N_5440,N_5157);
or U7011 (N_7011,N_5373,N_5097);
nand U7012 (N_7012,N_4745,N_4307);
xnor U7013 (N_7013,N_4392,N_5918);
and U7014 (N_7014,N_5855,N_4128);
nand U7015 (N_7015,N_4213,N_5810);
nand U7016 (N_7016,N_5013,N_4606);
and U7017 (N_7017,N_4151,N_5059);
xnor U7018 (N_7018,N_4117,N_5578);
xor U7019 (N_7019,N_4478,N_5636);
nand U7020 (N_7020,N_5962,N_4943);
or U7021 (N_7021,N_5267,N_5689);
nor U7022 (N_7022,N_5130,N_5508);
xor U7023 (N_7023,N_4569,N_4210);
xnor U7024 (N_7024,N_5155,N_5496);
nand U7025 (N_7025,N_5630,N_5328);
xnor U7026 (N_7026,N_4286,N_5818);
nand U7027 (N_7027,N_5297,N_4410);
and U7028 (N_7028,N_4765,N_4547);
or U7029 (N_7029,N_4086,N_4614);
and U7030 (N_7030,N_4027,N_4170);
nor U7031 (N_7031,N_4091,N_5176);
xnor U7032 (N_7032,N_5486,N_5900);
nor U7033 (N_7033,N_4915,N_5655);
and U7034 (N_7034,N_5839,N_4322);
nand U7035 (N_7035,N_5246,N_4515);
and U7036 (N_7036,N_4332,N_4098);
xor U7037 (N_7037,N_4265,N_5916);
nor U7038 (N_7038,N_5544,N_5280);
or U7039 (N_7039,N_5575,N_5562);
and U7040 (N_7040,N_4858,N_4932);
nor U7041 (N_7041,N_4145,N_5044);
or U7042 (N_7042,N_4793,N_5499);
nor U7043 (N_7043,N_4162,N_5727);
nand U7044 (N_7044,N_4334,N_4262);
xnor U7045 (N_7045,N_4164,N_5791);
nand U7046 (N_7046,N_5808,N_5511);
nor U7047 (N_7047,N_4721,N_5530);
xor U7048 (N_7048,N_4915,N_5860);
xor U7049 (N_7049,N_4938,N_4712);
or U7050 (N_7050,N_5922,N_4398);
nor U7051 (N_7051,N_4385,N_5239);
nand U7052 (N_7052,N_5750,N_4801);
nor U7053 (N_7053,N_5786,N_4286);
and U7054 (N_7054,N_5469,N_4365);
xor U7055 (N_7055,N_5896,N_5401);
or U7056 (N_7056,N_4251,N_4983);
and U7057 (N_7057,N_4053,N_4182);
nand U7058 (N_7058,N_5567,N_4371);
nand U7059 (N_7059,N_5921,N_4611);
nand U7060 (N_7060,N_5091,N_4818);
nand U7061 (N_7061,N_5077,N_5159);
and U7062 (N_7062,N_4745,N_5933);
and U7063 (N_7063,N_5484,N_4385);
or U7064 (N_7064,N_5229,N_5563);
and U7065 (N_7065,N_4510,N_5214);
and U7066 (N_7066,N_5180,N_4194);
xnor U7067 (N_7067,N_5560,N_4423);
xnor U7068 (N_7068,N_5049,N_4024);
nand U7069 (N_7069,N_5709,N_4604);
and U7070 (N_7070,N_5801,N_5821);
and U7071 (N_7071,N_5458,N_4063);
or U7072 (N_7072,N_4949,N_5419);
or U7073 (N_7073,N_4519,N_5089);
xnor U7074 (N_7074,N_5068,N_4978);
and U7075 (N_7075,N_5975,N_5724);
and U7076 (N_7076,N_5162,N_4468);
or U7077 (N_7077,N_4961,N_4138);
nor U7078 (N_7078,N_5307,N_5189);
or U7079 (N_7079,N_5275,N_5046);
and U7080 (N_7080,N_4339,N_4264);
and U7081 (N_7081,N_5646,N_4480);
and U7082 (N_7082,N_4953,N_4422);
nor U7083 (N_7083,N_5869,N_4972);
or U7084 (N_7084,N_5698,N_5154);
nor U7085 (N_7085,N_5396,N_5185);
nor U7086 (N_7086,N_5114,N_5463);
nand U7087 (N_7087,N_4821,N_4960);
nand U7088 (N_7088,N_5446,N_4796);
or U7089 (N_7089,N_5575,N_4547);
nor U7090 (N_7090,N_4444,N_5337);
nand U7091 (N_7091,N_4868,N_5924);
xnor U7092 (N_7092,N_4069,N_4131);
and U7093 (N_7093,N_5453,N_5861);
nor U7094 (N_7094,N_5219,N_4554);
nor U7095 (N_7095,N_5809,N_4499);
or U7096 (N_7096,N_4827,N_4414);
nand U7097 (N_7097,N_4808,N_4394);
and U7098 (N_7098,N_4460,N_5459);
or U7099 (N_7099,N_4384,N_4297);
and U7100 (N_7100,N_4548,N_4161);
nor U7101 (N_7101,N_4777,N_5088);
nand U7102 (N_7102,N_5035,N_4256);
nand U7103 (N_7103,N_4703,N_4228);
xor U7104 (N_7104,N_4290,N_4723);
nor U7105 (N_7105,N_5917,N_4489);
nand U7106 (N_7106,N_4195,N_5771);
or U7107 (N_7107,N_4652,N_4379);
nand U7108 (N_7108,N_4056,N_4216);
and U7109 (N_7109,N_4597,N_4186);
nand U7110 (N_7110,N_4282,N_4476);
or U7111 (N_7111,N_4451,N_4443);
or U7112 (N_7112,N_5973,N_5740);
and U7113 (N_7113,N_4037,N_4801);
nand U7114 (N_7114,N_4197,N_4776);
nor U7115 (N_7115,N_4908,N_4229);
or U7116 (N_7116,N_4348,N_5937);
xnor U7117 (N_7117,N_4503,N_5153);
xor U7118 (N_7118,N_5123,N_4842);
nor U7119 (N_7119,N_4878,N_4625);
xor U7120 (N_7120,N_4719,N_4103);
nor U7121 (N_7121,N_4522,N_5309);
or U7122 (N_7122,N_5143,N_5066);
and U7123 (N_7123,N_5554,N_4351);
nor U7124 (N_7124,N_5099,N_5349);
or U7125 (N_7125,N_4732,N_4198);
nor U7126 (N_7126,N_5347,N_4016);
or U7127 (N_7127,N_4105,N_4646);
or U7128 (N_7128,N_4704,N_5671);
xor U7129 (N_7129,N_5963,N_5853);
or U7130 (N_7130,N_4669,N_5142);
nand U7131 (N_7131,N_5316,N_5548);
nand U7132 (N_7132,N_4044,N_5569);
xor U7133 (N_7133,N_4001,N_5116);
and U7134 (N_7134,N_5451,N_4403);
and U7135 (N_7135,N_5269,N_4788);
or U7136 (N_7136,N_4521,N_5954);
nand U7137 (N_7137,N_5424,N_4998);
xnor U7138 (N_7138,N_5966,N_4600);
nand U7139 (N_7139,N_4186,N_5440);
nor U7140 (N_7140,N_5204,N_5246);
nor U7141 (N_7141,N_5455,N_5478);
nor U7142 (N_7142,N_5030,N_5031);
nand U7143 (N_7143,N_5387,N_4777);
nor U7144 (N_7144,N_5437,N_4834);
nand U7145 (N_7145,N_5538,N_5966);
nor U7146 (N_7146,N_4279,N_5335);
nor U7147 (N_7147,N_5686,N_5099);
xnor U7148 (N_7148,N_4830,N_4070);
xor U7149 (N_7149,N_5019,N_5183);
xor U7150 (N_7150,N_4799,N_4766);
nand U7151 (N_7151,N_5001,N_5406);
nand U7152 (N_7152,N_5304,N_5065);
nor U7153 (N_7153,N_4309,N_5831);
nor U7154 (N_7154,N_4129,N_4893);
nor U7155 (N_7155,N_5979,N_4154);
nand U7156 (N_7156,N_5552,N_4808);
xnor U7157 (N_7157,N_4318,N_4495);
and U7158 (N_7158,N_4048,N_5797);
or U7159 (N_7159,N_5384,N_4123);
xor U7160 (N_7160,N_5896,N_5347);
and U7161 (N_7161,N_5987,N_5877);
and U7162 (N_7162,N_5660,N_4995);
xor U7163 (N_7163,N_4650,N_5424);
and U7164 (N_7164,N_4756,N_5020);
xor U7165 (N_7165,N_5246,N_5049);
and U7166 (N_7166,N_4900,N_4127);
nor U7167 (N_7167,N_4327,N_5440);
or U7168 (N_7168,N_4895,N_5785);
or U7169 (N_7169,N_5307,N_5744);
nand U7170 (N_7170,N_4418,N_4533);
xor U7171 (N_7171,N_4757,N_5875);
and U7172 (N_7172,N_4445,N_4065);
nor U7173 (N_7173,N_5132,N_4753);
nor U7174 (N_7174,N_5635,N_5195);
and U7175 (N_7175,N_4436,N_4557);
and U7176 (N_7176,N_5140,N_4557);
nor U7177 (N_7177,N_5037,N_4396);
and U7178 (N_7178,N_5508,N_4479);
nand U7179 (N_7179,N_5622,N_5139);
nand U7180 (N_7180,N_4308,N_5118);
nand U7181 (N_7181,N_5624,N_4205);
xnor U7182 (N_7182,N_4923,N_5481);
or U7183 (N_7183,N_4267,N_4472);
or U7184 (N_7184,N_5189,N_4907);
or U7185 (N_7185,N_5548,N_4912);
and U7186 (N_7186,N_4427,N_5453);
and U7187 (N_7187,N_4874,N_5724);
and U7188 (N_7188,N_5949,N_5731);
nor U7189 (N_7189,N_4761,N_5666);
or U7190 (N_7190,N_4424,N_5723);
nand U7191 (N_7191,N_4184,N_4880);
nor U7192 (N_7192,N_5987,N_4812);
and U7193 (N_7193,N_4063,N_5118);
and U7194 (N_7194,N_5461,N_5583);
xor U7195 (N_7195,N_4048,N_5174);
and U7196 (N_7196,N_4148,N_4561);
nor U7197 (N_7197,N_4965,N_5291);
nor U7198 (N_7198,N_5009,N_4165);
and U7199 (N_7199,N_4348,N_5680);
nand U7200 (N_7200,N_4773,N_4801);
and U7201 (N_7201,N_5098,N_4347);
or U7202 (N_7202,N_5126,N_5311);
and U7203 (N_7203,N_4667,N_5667);
nand U7204 (N_7204,N_5161,N_5253);
or U7205 (N_7205,N_4322,N_5127);
and U7206 (N_7206,N_4164,N_5175);
and U7207 (N_7207,N_5199,N_5163);
and U7208 (N_7208,N_4088,N_5840);
and U7209 (N_7209,N_4081,N_4255);
xnor U7210 (N_7210,N_4640,N_5690);
nor U7211 (N_7211,N_4563,N_4986);
nand U7212 (N_7212,N_4253,N_5806);
xor U7213 (N_7213,N_5239,N_4052);
or U7214 (N_7214,N_5851,N_5893);
or U7215 (N_7215,N_5274,N_4485);
and U7216 (N_7216,N_4256,N_4865);
xnor U7217 (N_7217,N_4870,N_4599);
nand U7218 (N_7218,N_5518,N_4285);
nand U7219 (N_7219,N_5780,N_4355);
xnor U7220 (N_7220,N_5751,N_5528);
nor U7221 (N_7221,N_5639,N_5528);
and U7222 (N_7222,N_4037,N_5575);
nand U7223 (N_7223,N_5593,N_5270);
nor U7224 (N_7224,N_4886,N_5044);
nand U7225 (N_7225,N_4023,N_5471);
nor U7226 (N_7226,N_5888,N_5558);
and U7227 (N_7227,N_5931,N_4395);
xor U7228 (N_7228,N_4664,N_4280);
nor U7229 (N_7229,N_4913,N_4612);
xor U7230 (N_7230,N_4206,N_5236);
or U7231 (N_7231,N_5966,N_4731);
nand U7232 (N_7232,N_5460,N_4455);
xor U7233 (N_7233,N_4410,N_4560);
and U7234 (N_7234,N_5411,N_5530);
or U7235 (N_7235,N_5899,N_4112);
and U7236 (N_7236,N_4818,N_5382);
nor U7237 (N_7237,N_5604,N_5676);
nor U7238 (N_7238,N_5995,N_5621);
xnor U7239 (N_7239,N_4952,N_4480);
and U7240 (N_7240,N_4039,N_4962);
xnor U7241 (N_7241,N_5870,N_5365);
or U7242 (N_7242,N_5978,N_4928);
xnor U7243 (N_7243,N_4882,N_4632);
or U7244 (N_7244,N_5872,N_5060);
nor U7245 (N_7245,N_5776,N_4466);
or U7246 (N_7246,N_4032,N_5637);
xnor U7247 (N_7247,N_5354,N_4264);
and U7248 (N_7248,N_4464,N_4106);
and U7249 (N_7249,N_4635,N_4876);
nand U7250 (N_7250,N_5085,N_4003);
and U7251 (N_7251,N_4509,N_5027);
and U7252 (N_7252,N_4691,N_4399);
nand U7253 (N_7253,N_5621,N_4733);
xnor U7254 (N_7254,N_5157,N_5364);
xor U7255 (N_7255,N_4567,N_4173);
nor U7256 (N_7256,N_5331,N_5447);
nand U7257 (N_7257,N_5306,N_5147);
xor U7258 (N_7258,N_4452,N_4333);
or U7259 (N_7259,N_4403,N_5358);
xnor U7260 (N_7260,N_5973,N_4793);
xor U7261 (N_7261,N_4566,N_4424);
or U7262 (N_7262,N_5497,N_5016);
or U7263 (N_7263,N_4142,N_5342);
xor U7264 (N_7264,N_4441,N_4111);
nand U7265 (N_7265,N_4067,N_4358);
nor U7266 (N_7266,N_5618,N_5249);
nand U7267 (N_7267,N_4368,N_5225);
and U7268 (N_7268,N_4735,N_4946);
and U7269 (N_7269,N_4018,N_5725);
nand U7270 (N_7270,N_5672,N_5010);
nand U7271 (N_7271,N_4573,N_4524);
nor U7272 (N_7272,N_4842,N_4155);
or U7273 (N_7273,N_4844,N_4038);
xnor U7274 (N_7274,N_4795,N_5810);
xor U7275 (N_7275,N_4128,N_4860);
or U7276 (N_7276,N_4340,N_5911);
xnor U7277 (N_7277,N_5273,N_4306);
xor U7278 (N_7278,N_5510,N_5938);
and U7279 (N_7279,N_4926,N_5864);
or U7280 (N_7280,N_4648,N_5481);
nand U7281 (N_7281,N_4578,N_5313);
nor U7282 (N_7282,N_4031,N_4687);
nor U7283 (N_7283,N_4578,N_4971);
and U7284 (N_7284,N_4090,N_4393);
nor U7285 (N_7285,N_4781,N_5469);
or U7286 (N_7286,N_5540,N_4439);
or U7287 (N_7287,N_5511,N_4915);
or U7288 (N_7288,N_4040,N_5641);
xnor U7289 (N_7289,N_5709,N_5411);
xnor U7290 (N_7290,N_5924,N_5532);
and U7291 (N_7291,N_5092,N_4004);
and U7292 (N_7292,N_4140,N_4265);
nand U7293 (N_7293,N_5239,N_4963);
nor U7294 (N_7294,N_5454,N_5545);
and U7295 (N_7295,N_5704,N_4509);
or U7296 (N_7296,N_4423,N_4418);
nor U7297 (N_7297,N_4311,N_4616);
or U7298 (N_7298,N_4779,N_4586);
nor U7299 (N_7299,N_5533,N_5365);
nand U7300 (N_7300,N_5115,N_5766);
nand U7301 (N_7301,N_4067,N_4039);
nand U7302 (N_7302,N_5518,N_4464);
nand U7303 (N_7303,N_5704,N_5672);
nand U7304 (N_7304,N_4614,N_5584);
nor U7305 (N_7305,N_4358,N_5291);
nor U7306 (N_7306,N_4346,N_5352);
or U7307 (N_7307,N_4797,N_5105);
xor U7308 (N_7308,N_4509,N_5376);
and U7309 (N_7309,N_5244,N_4796);
and U7310 (N_7310,N_5801,N_4589);
and U7311 (N_7311,N_4601,N_5161);
xor U7312 (N_7312,N_4740,N_5424);
xor U7313 (N_7313,N_4855,N_4052);
nand U7314 (N_7314,N_5947,N_5441);
or U7315 (N_7315,N_4514,N_4975);
and U7316 (N_7316,N_5645,N_5475);
or U7317 (N_7317,N_4230,N_4619);
xnor U7318 (N_7318,N_5351,N_4572);
nand U7319 (N_7319,N_4460,N_4228);
nand U7320 (N_7320,N_5953,N_5877);
and U7321 (N_7321,N_5823,N_5949);
nand U7322 (N_7322,N_5933,N_5055);
or U7323 (N_7323,N_5101,N_4898);
xor U7324 (N_7324,N_4521,N_4649);
or U7325 (N_7325,N_4424,N_5155);
and U7326 (N_7326,N_5160,N_4356);
and U7327 (N_7327,N_5482,N_5489);
nor U7328 (N_7328,N_4686,N_5299);
and U7329 (N_7329,N_5212,N_4777);
and U7330 (N_7330,N_5811,N_4587);
xnor U7331 (N_7331,N_4924,N_4034);
and U7332 (N_7332,N_4195,N_4502);
nor U7333 (N_7333,N_5886,N_4343);
xnor U7334 (N_7334,N_5745,N_4317);
xor U7335 (N_7335,N_4752,N_5087);
and U7336 (N_7336,N_5949,N_4272);
and U7337 (N_7337,N_5875,N_5796);
nand U7338 (N_7338,N_5426,N_4733);
or U7339 (N_7339,N_5457,N_5176);
nand U7340 (N_7340,N_5799,N_5929);
nor U7341 (N_7341,N_4327,N_4018);
xor U7342 (N_7342,N_4595,N_4277);
nor U7343 (N_7343,N_4167,N_4144);
xor U7344 (N_7344,N_5351,N_5191);
and U7345 (N_7345,N_5193,N_4486);
or U7346 (N_7346,N_5121,N_5245);
or U7347 (N_7347,N_4352,N_4722);
nor U7348 (N_7348,N_4738,N_5771);
or U7349 (N_7349,N_4299,N_5873);
or U7350 (N_7350,N_4106,N_4154);
nor U7351 (N_7351,N_4561,N_5509);
xor U7352 (N_7352,N_5430,N_5736);
and U7353 (N_7353,N_4556,N_5668);
xnor U7354 (N_7354,N_5615,N_4647);
xnor U7355 (N_7355,N_5230,N_4466);
nor U7356 (N_7356,N_5512,N_4604);
nand U7357 (N_7357,N_4432,N_5950);
or U7358 (N_7358,N_4936,N_5707);
nor U7359 (N_7359,N_5012,N_5513);
xnor U7360 (N_7360,N_5593,N_5946);
xor U7361 (N_7361,N_4572,N_5662);
nand U7362 (N_7362,N_4653,N_4503);
nand U7363 (N_7363,N_5568,N_5119);
nor U7364 (N_7364,N_4013,N_5177);
or U7365 (N_7365,N_5956,N_4268);
xnor U7366 (N_7366,N_4716,N_4804);
nand U7367 (N_7367,N_4349,N_5303);
and U7368 (N_7368,N_5422,N_4011);
and U7369 (N_7369,N_5675,N_4102);
nand U7370 (N_7370,N_5014,N_4541);
and U7371 (N_7371,N_4431,N_4365);
xnor U7372 (N_7372,N_5881,N_4576);
or U7373 (N_7373,N_5526,N_5513);
xor U7374 (N_7374,N_5679,N_5903);
and U7375 (N_7375,N_5479,N_4430);
or U7376 (N_7376,N_4910,N_5701);
xor U7377 (N_7377,N_5254,N_4490);
or U7378 (N_7378,N_4396,N_4493);
and U7379 (N_7379,N_4420,N_5606);
or U7380 (N_7380,N_4178,N_4481);
and U7381 (N_7381,N_5415,N_5510);
nor U7382 (N_7382,N_5288,N_5419);
nand U7383 (N_7383,N_4191,N_5951);
nor U7384 (N_7384,N_4419,N_4771);
nor U7385 (N_7385,N_4839,N_5263);
or U7386 (N_7386,N_4036,N_4821);
xor U7387 (N_7387,N_5073,N_4917);
xnor U7388 (N_7388,N_5039,N_5441);
and U7389 (N_7389,N_4901,N_4894);
nand U7390 (N_7390,N_5745,N_5896);
nand U7391 (N_7391,N_5726,N_4097);
nand U7392 (N_7392,N_4287,N_5268);
and U7393 (N_7393,N_4400,N_4600);
or U7394 (N_7394,N_5252,N_4722);
nand U7395 (N_7395,N_5064,N_4664);
nor U7396 (N_7396,N_4213,N_5248);
xnor U7397 (N_7397,N_4492,N_4859);
xnor U7398 (N_7398,N_4670,N_4597);
or U7399 (N_7399,N_4332,N_4851);
nor U7400 (N_7400,N_4017,N_4032);
xor U7401 (N_7401,N_5751,N_5272);
nor U7402 (N_7402,N_5447,N_4064);
and U7403 (N_7403,N_4538,N_5460);
xor U7404 (N_7404,N_5672,N_5953);
nand U7405 (N_7405,N_5823,N_4061);
xnor U7406 (N_7406,N_4002,N_5714);
and U7407 (N_7407,N_5403,N_4589);
and U7408 (N_7408,N_5989,N_5450);
xnor U7409 (N_7409,N_4372,N_5484);
xor U7410 (N_7410,N_5456,N_5052);
or U7411 (N_7411,N_4911,N_5544);
or U7412 (N_7412,N_4799,N_5393);
nand U7413 (N_7413,N_5343,N_4993);
nand U7414 (N_7414,N_5342,N_5385);
xor U7415 (N_7415,N_5526,N_4912);
nor U7416 (N_7416,N_5896,N_4623);
and U7417 (N_7417,N_4333,N_4658);
xnor U7418 (N_7418,N_4857,N_4926);
nor U7419 (N_7419,N_5044,N_4489);
and U7420 (N_7420,N_4073,N_5872);
and U7421 (N_7421,N_4767,N_5938);
nor U7422 (N_7422,N_4111,N_4697);
nor U7423 (N_7423,N_4458,N_5407);
xnor U7424 (N_7424,N_5192,N_5453);
and U7425 (N_7425,N_4258,N_4059);
xnor U7426 (N_7426,N_4386,N_4921);
nand U7427 (N_7427,N_5203,N_4811);
nor U7428 (N_7428,N_4554,N_5570);
or U7429 (N_7429,N_4051,N_4698);
and U7430 (N_7430,N_5941,N_4803);
nand U7431 (N_7431,N_4811,N_4541);
and U7432 (N_7432,N_5604,N_4863);
nor U7433 (N_7433,N_5305,N_5835);
or U7434 (N_7434,N_4812,N_4595);
and U7435 (N_7435,N_4775,N_5668);
nand U7436 (N_7436,N_5062,N_4331);
nand U7437 (N_7437,N_4101,N_5288);
nor U7438 (N_7438,N_5422,N_5996);
or U7439 (N_7439,N_5244,N_4059);
and U7440 (N_7440,N_5717,N_4817);
nor U7441 (N_7441,N_4153,N_4598);
and U7442 (N_7442,N_5338,N_4007);
nand U7443 (N_7443,N_4695,N_4097);
nand U7444 (N_7444,N_5866,N_4121);
or U7445 (N_7445,N_4114,N_4110);
nor U7446 (N_7446,N_4901,N_5697);
and U7447 (N_7447,N_4585,N_5499);
nor U7448 (N_7448,N_5029,N_5484);
nand U7449 (N_7449,N_5382,N_5900);
nor U7450 (N_7450,N_4952,N_4455);
xor U7451 (N_7451,N_5520,N_5121);
and U7452 (N_7452,N_4397,N_5662);
xor U7453 (N_7453,N_4936,N_5360);
nor U7454 (N_7454,N_5239,N_5474);
nor U7455 (N_7455,N_5871,N_4150);
nand U7456 (N_7456,N_5128,N_4661);
or U7457 (N_7457,N_4535,N_4007);
nand U7458 (N_7458,N_4718,N_4027);
and U7459 (N_7459,N_5652,N_4628);
and U7460 (N_7460,N_5395,N_5681);
or U7461 (N_7461,N_5382,N_5826);
nor U7462 (N_7462,N_4491,N_4969);
and U7463 (N_7463,N_4230,N_5834);
xnor U7464 (N_7464,N_5673,N_5098);
and U7465 (N_7465,N_4205,N_4830);
xor U7466 (N_7466,N_5261,N_4850);
and U7467 (N_7467,N_5270,N_5347);
xnor U7468 (N_7468,N_4212,N_4144);
xor U7469 (N_7469,N_4161,N_4816);
xor U7470 (N_7470,N_4936,N_5343);
and U7471 (N_7471,N_5747,N_5714);
xor U7472 (N_7472,N_4303,N_5725);
and U7473 (N_7473,N_5407,N_5733);
nor U7474 (N_7474,N_5889,N_4763);
or U7475 (N_7475,N_4019,N_5921);
xor U7476 (N_7476,N_4362,N_4701);
nand U7477 (N_7477,N_4985,N_5848);
xor U7478 (N_7478,N_5723,N_4255);
nor U7479 (N_7479,N_4398,N_5987);
or U7480 (N_7480,N_4073,N_4844);
nor U7481 (N_7481,N_4311,N_4943);
and U7482 (N_7482,N_4944,N_4882);
and U7483 (N_7483,N_4812,N_4774);
or U7484 (N_7484,N_4471,N_5416);
xnor U7485 (N_7485,N_4709,N_4003);
nand U7486 (N_7486,N_5599,N_4470);
nand U7487 (N_7487,N_4917,N_4624);
xnor U7488 (N_7488,N_5207,N_5530);
nand U7489 (N_7489,N_5759,N_5119);
nor U7490 (N_7490,N_5078,N_4200);
or U7491 (N_7491,N_5405,N_5029);
nor U7492 (N_7492,N_5565,N_4130);
xor U7493 (N_7493,N_5357,N_5680);
and U7494 (N_7494,N_4666,N_5315);
xnor U7495 (N_7495,N_5906,N_5717);
nand U7496 (N_7496,N_5594,N_4283);
or U7497 (N_7497,N_4139,N_4923);
xnor U7498 (N_7498,N_4145,N_4132);
and U7499 (N_7499,N_4573,N_5278);
xnor U7500 (N_7500,N_4966,N_5405);
and U7501 (N_7501,N_5107,N_4390);
nand U7502 (N_7502,N_4543,N_5365);
nor U7503 (N_7503,N_4108,N_5693);
xnor U7504 (N_7504,N_4535,N_4849);
nor U7505 (N_7505,N_5380,N_4512);
or U7506 (N_7506,N_4788,N_4813);
xnor U7507 (N_7507,N_4844,N_5832);
or U7508 (N_7508,N_4886,N_4624);
xnor U7509 (N_7509,N_4189,N_4754);
nor U7510 (N_7510,N_5510,N_5656);
nand U7511 (N_7511,N_4530,N_4337);
and U7512 (N_7512,N_4676,N_4235);
nand U7513 (N_7513,N_4774,N_5173);
and U7514 (N_7514,N_4421,N_5434);
xor U7515 (N_7515,N_4713,N_4926);
and U7516 (N_7516,N_4140,N_4387);
or U7517 (N_7517,N_4256,N_5356);
or U7518 (N_7518,N_5751,N_5425);
nor U7519 (N_7519,N_4099,N_4631);
or U7520 (N_7520,N_4962,N_5553);
or U7521 (N_7521,N_4529,N_4807);
xnor U7522 (N_7522,N_5575,N_5821);
nand U7523 (N_7523,N_5390,N_4499);
and U7524 (N_7524,N_5170,N_5908);
nand U7525 (N_7525,N_4389,N_5966);
nor U7526 (N_7526,N_4466,N_5490);
nor U7527 (N_7527,N_4033,N_5291);
xor U7528 (N_7528,N_4338,N_5935);
xor U7529 (N_7529,N_5226,N_5728);
xnor U7530 (N_7530,N_4770,N_5180);
nand U7531 (N_7531,N_5831,N_5294);
or U7532 (N_7532,N_5165,N_4896);
or U7533 (N_7533,N_4730,N_4128);
or U7534 (N_7534,N_4171,N_5254);
xnor U7535 (N_7535,N_5435,N_5489);
and U7536 (N_7536,N_4472,N_4300);
xnor U7537 (N_7537,N_4182,N_4094);
xnor U7538 (N_7538,N_5282,N_4006);
or U7539 (N_7539,N_4129,N_4662);
xor U7540 (N_7540,N_4332,N_4285);
and U7541 (N_7541,N_4777,N_5126);
nand U7542 (N_7542,N_5158,N_4231);
or U7543 (N_7543,N_5777,N_4406);
nand U7544 (N_7544,N_4203,N_4431);
nand U7545 (N_7545,N_4589,N_4553);
nor U7546 (N_7546,N_4260,N_5833);
or U7547 (N_7547,N_5525,N_4637);
nand U7548 (N_7548,N_5447,N_4195);
nor U7549 (N_7549,N_4718,N_5532);
xor U7550 (N_7550,N_5514,N_5678);
xnor U7551 (N_7551,N_4178,N_4959);
nand U7552 (N_7552,N_4205,N_5371);
nor U7553 (N_7553,N_5503,N_4071);
nand U7554 (N_7554,N_4786,N_5768);
nand U7555 (N_7555,N_5199,N_5207);
xnor U7556 (N_7556,N_5777,N_5863);
xor U7557 (N_7557,N_4388,N_4382);
and U7558 (N_7558,N_5972,N_4844);
xnor U7559 (N_7559,N_4565,N_4200);
or U7560 (N_7560,N_5743,N_5176);
nand U7561 (N_7561,N_4912,N_4913);
and U7562 (N_7562,N_4780,N_5395);
nand U7563 (N_7563,N_5424,N_5590);
or U7564 (N_7564,N_4579,N_4307);
or U7565 (N_7565,N_4029,N_5646);
nand U7566 (N_7566,N_4811,N_5195);
or U7567 (N_7567,N_4808,N_4663);
and U7568 (N_7568,N_5845,N_5559);
xnor U7569 (N_7569,N_5974,N_4007);
or U7570 (N_7570,N_4921,N_4765);
nand U7571 (N_7571,N_5222,N_5162);
nand U7572 (N_7572,N_5782,N_4607);
nor U7573 (N_7573,N_4408,N_4124);
or U7574 (N_7574,N_4117,N_4657);
nand U7575 (N_7575,N_5629,N_4528);
nand U7576 (N_7576,N_4376,N_4476);
nor U7577 (N_7577,N_4710,N_5446);
nor U7578 (N_7578,N_4371,N_5991);
and U7579 (N_7579,N_4391,N_5204);
and U7580 (N_7580,N_5088,N_4455);
xnor U7581 (N_7581,N_5168,N_5304);
nor U7582 (N_7582,N_4213,N_4050);
nand U7583 (N_7583,N_5696,N_5052);
nor U7584 (N_7584,N_4071,N_5808);
or U7585 (N_7585,N_4153,N_5350);
nor U7586 (N_7586,N_5190,N_4365);
and U7587 (N_7587,N_4338,N_4572);
nand U7588 (N_7588,N_4242,N_4500);
xor U7589 (N_7589,N_4257,N_5011);
or U7590 (N_7590,N_4765,N_5829);
or U7591 (N_7591,N_4073,N_4782);
xnor U7592 (N_7592,N_5901,N_5168);
xor U7593 (N_7593,N_4260,N_5424);
xor U7594 (N_7594,N_4932,N_4171);
and U7595 (N_7595,N_5618,N_4443);
or U7596 (N_7596,N_4804,N_5090);
and U7597 (N_7597,N_5502,N_4211);
and U7598 (N_7598,N_4674,N_5784);
nand U7599 (N_7599,N_5347,N_4540);
and U7600 (N_7600,N_5941,N_4223);
nor U7601 (N_7601,N_5936,N_4260);
nand U7602 (N_7602,N_5443,N_5217);
and U7603 (N_7603,N_4327,N_4472);
xor U7604 (N_7604,N_4555,N_4961);
xor U7605 (N_7605,N_4572,N_4304);
and U7606 (N_7606,N_4539,N_5824);
nand U7607 (N_7607,N_4314,N_4716);
nor U7608 (N_7608,N_5694,N_5467);
nor U7609 (N_7609,N_4187,N_4933);
xnor U7610 (N_7610,N_4077,N_4363);
nand U7611 (N_7611,N_4444,N_5027);
xor U7612 (N_7612,N_4508,N_5706);
nor U7613 (N_7613,N_5021,N_5764);
nor U7614 (N_7614,N_4004,N_5024);
or U7615 (N_7615,N_5345,N_4195);
or U7616 (N_7616,N_5465,N_5036);
nand U7617 (N_7617,N_4414,N_4078);
nor U7618 (N_7618,N_5642,N_4691);
or U7619 (N_7619,N_5724,N_4858);
nor U7620 (N_7620,N_5017,N_5046);
xor U7621 (N_7621,N_5048,N_5549);
xor U7622 (N_7622,N_4350,N_5057);
xnor U7623 (N_7623,N_5759,N_4147);
nand U7624 (N_7624,N_5706,N_5901);
xor U7625 (N_7625,N_4867,N_4800);
nor U7626 (N_7626,N_5153,N_5424);
and U7627 (N_7627,N_5916,N_5474);
nand U7628 (N_7628,N_5129,N_4658);
nor U7629 (N_7629,N_5711,N_5167);
or U7630 (N_7630,N_5505,N_5496);
nand U7631 (N_7631,N_4379,N_4114);
nand U7632 (N_7632,N_5450,N_5401);
or U7633 (N_7633,N_5377,N_5806);
nand U7634 (N_7634,N_5165,N_4194);
xnor U7635 (N_7635,N_5288,N_4842);
nand U7636 (N_7636,N_5239,N_4653);
and U7637 (N_7637,N_4648,N_4840);
nand U7638 (N_7638,N_5945,N_4780);
and U7639 (N_7639,N_4767,N_5812);
nor U7640 (N_7640,N_4324,N_4910);
xnor U7641 (N_7641,N_5605,N_4657);
nand U7642 (N_7642,N_5333,N_4983);
nor U7643 (N_7643,N_5115,N_4386);
xnor U7644 (N_7644,N_5496,N_5047);
or U7645 (N_7645,N_5983,N_4060);
nor U7646 (N_7646,N_5235,N_4848);
nor U7647 (N_7647,N_4652,N_4998);
or U7648 (N_7648,N_5186,N_5658);
and U7649 (N_7649,N_4503,N_5175);
xor U7650 (N_7650,N_5911,N_4287);
or U7651 (N_7651,N_5151,N_4023);
xnor U7652 (N_7652,N_4536,N_4606);
or U7653 (N_7653,N_5225,N_4436);
nand U7654 (N_7654,N_5685,N_5793);
nor U7655 (N_7655,N_5967,N_5045);
and U7656 (N_7656,N_5295,N_5711);
and U7657 (N_7657,N_5238,N_5096);
nor U7658 (N_7658,N_5235,N_5053);
and U7659 (N_7659,N_4778,N_4916);
nor U7660 (N_7660,N_4439,N_5807);
or U7661 (N_7661,N_4373,N_4525);
or U7662 (N_7662,N_4108,N_5577);
nand U7663 (N_7663,N_5126,N_5676);
nor U7664 (N_7664,N_4859,N_5165);
xor U7665 (N_7665,N_4096,N_4810);
xor U7666 (N_7666,N_4516,N_4233);
xnor U7667 (N_7667,N_5224,N_5963);
and U7668 (N_7668,N_4509,N_4698);
and U7669 (N_7669,N_5927,N_5588);
xnor U7670 (N_7670,N_5035,N_4656);
nand U7671 (N_7671,N_5056,N_5866);
xor U7672 (N_7672,N_5352,N_5675);
and U7673 (N_7673,N_4102,N_5888);
nand U7674 (N_7674,N_5125,N_5054);
nand U7675 (N_7675,N_5199,N_4920);
xnor U7676 (N_7676,N_4906,N_4010);
or U7677 (N_7677,N_4676,N_4154);
and U7678 (N_7678,N_4405,N_4494);
and U7679 (N_7679,N_4247,N_4331);
nor U7680 (N_7680,N_5027,N_5920);
nand U7681 (N_7681,N_5071,N_5915);
nor U7682 (N_7682,N_4948,N_4556);
xnor U7683 (N_7683,N_5068,N_5980);
xor U7684 (N_7684,N_4019,N_5962);
nand U7685 (N_7685,N_4821,N_4292);
xnor U7686 (N_7686,N_4970,N_4337);
or U7687 (N_7687,N_5654,N_4451);
or U7688 (N_7688,N_5828,N_5688);
xor U7689 (N_7689,N_5985,N_4135);
xnor U7690 (N_7690,N_5285,N_4438);
or U7691 (N_7691,N_5125,N_4102);
nor U7692 (N_7692,N_4148,N_4790);
nor U7693 (N_7693,N_4133,N_5214);
nand U7694 (N_7694,N_4376,N_4883);
nand U7695 (N_7695,N_5129,N_4271);
and U7696 (N_7696,N_5267,N_5214);
nor U7697 (N_7697,N_5355,N_5164);
or U7698 (N_7698,N_5307,N_4471);
xnor U7699 (N_7699,N_4154,N_4684);
and U7700 (N_7700,N_4601,N_5590);
nand U7701 (N_7701,N_4992,N_5180);
or U7702 (N_7702,N_4307,N_5029);
xnor U7703 (N_7703,N_4203,N_5245);
xnor U7704 (N_7704,N_4701,N_5085);
or U7705 (N_7705,N_4414,N_5940);
and U7706 (N_7706,N_5791,N_4654);
nand U7707 (N_7707,N_4662,N_4101);
nand U7708 (N_7708,N_5212,N_5972);
nand U7709 (N_7709,N_5984,N_5295);
nand U7710 (N_7710,N_4316,N_5106);
xor U7711 (N_7711,N_5462,N_4113);
or U7712 (N_7712,N_4787,N_4212);
xor U7713 (N_7713,N_4493,N_4500);
nor U7714 (N_7714,N_4121,N_4758);
or U7715 (N_7715,N_5824,N_4197);
nand U7716 (N_7716,N_4653,N_4369);
and U7717 (N_7717,N_4660,N_4616);
nor U7718 (N_7718,N_5933,N_5560);
and U7719 (N_7719,N_4579,N_5886);
xor U7720 (N_7720,N_4020,N_5850);
and U7721 (N_7721,N_5984,N_4934);
xor U7722 (N_7722,N_4197,N_5831);
and U7723 (N_7723,N_4224,N_4784);
nand U7724 (N_7724,N_4612,N_5238);
or U7725 (N_7725,N_4775,N_4116);
xor U7726 (N_7726,N_4334,N_5676);
xor U7727 (N_7727,N_5890,N_5990);
or U7728 (N_7728,N_4098,N_5943);
nand U7729 (N_7729,N_4143,N_4474);
nand U7730 (N_7730,N_4283,N_4012);
and U7731 (N_7731,N_4335,N_5237);
xnor U7732 (N_7732,N_5242,N_5405);
or U7733 (N_7733,N_4652,N_5927);
and U7734 (N_7734,N_4818,N_4420);
xor U7735 (N_7735,N_4565,N_5798);
or U7736 (N_7736,N_5452,N_4278);
xnor U7737 (N_7737,N_4852,N_4631);
and U7738 (N_7738,N_4051,N_4949);
xnor U7739 (N_7739,N_4542,N_5616);
nor U7740 (N_7740,N_4338,N_5621);
or U7741 (N_7741,N_4381,N_4704);
xnor U7742 (N_7742,N_5681,N_4704);
and U7743 (N_7743,N_4558,N_4764);
and U7744 (N_7744,N_4599,N_5530);
and U7745 (N_7745,N_4842,N_5057);
or U7746 (N_7746,N_4442,N_5712);
nand U7747 (N_7747,N_4796,N_5944);
nor U7748 (N_7748,N_5528,N_5437);
and U7749 (N_7749,N_5382,N_4554);
or U7750 (N_7750,N_5852,N_4951);
or U7751 (N_7751,N_4414,N_4437);
and U7752 (N_7752,N_4804,N_4026);
or U7753 (N_7753,N_4690,N_5566);
nor U7754 (N_7754,N_5235,N_5352);
nor U7755 (N_7755,N_4656,N_4556);
and U7756 (N_7756,N_5004,N_4453);
xor U7757 (N_7757,N_4570,N_4866);
nor U7758 (N_7758,N_5532,N_4077);
nor U7759 (N_7759,N_4483,N_5941);
nand U7760 (N_7760,N_4390,N_5186);
nand U7761 (N_7761,N_5094,N_5063);
nor U7762 (N_7762,N_4857,N_4809);
nand U7763 (N_7763,N_5832,N_5669);
nand U7764 (N_7764,N_4263,N_5796);
nor U7765 (N_7765,N_5793,N_4582);
and U7766 (N_7766,N_4796,N_5803);
nor U7767 (N_7767,N_4248,N_5660);
nor U7768 (N_7768,N_5930,N_4169);
nor U7769 (N_7769,N_4902,N_5735);
or U7770 (N_7770,N_4768,N_5555);
nor U7771 (N_7771,N_5533,N_5377);
or U7772 (N_7772,N_5397,N_4464);
xor U7773 (N_7773,N_4751,N_5559);
nand U7774 (N_7774,N_5038,N_5826);
or U7775 (N_7775,N_5794,N_5362);
and U7776 (N_7776,N_5421,N_4740);
and U7777 (N_7777,N_4594,N_4608);
nor U7778 (N_7778,N_5817,N_5672);
nand U7779 (N_7779,N_5658,N_5678);
nand U7780 (N_7780,N_5246,N_5668);
xnor U7781 (N_7781,N_4848,N_4850);
or U7782 (N_7782,N_5980,N_4997);
nand U7783 (N_7783,N_4794,N_5612);
or U7784 (N_7784,N_4175,N_4246);
nand U7785 (N_7785,N_5473,N_4768);
and U7786 (N_7786,N_4950,N_5676);
nor U7787 (N_7787,N_5224,N_5644);
or U7788 (N_7788,N_5252,N_5919);
nor U7789 (N_7789,N_5850,N_5096);
nor U7790 (N_7790,N_5058,N_4919);
nand U7791 (N_7791,N_4797,N_4764);
nor U7792 (N_7792,N_5025,N_4969);
xor U7793 (N_7793,N_5923,N_4745);
nand U7794 (N_7794,N_4131,N_5806);
nand U7795 (N_7795,N_5350,N_4239);
xnor U7796 (N_7796,N_5131,N_4708);
or U7797 (N_7797,N_4601,N_4431);
nand U7798 (N_7798,N_5947,N_5627);
nor U7799 (N_7799,N_4465,N_5983);
xor U7800 (N_7800,N_4607,N_4594);
xor U7801 (N_7801,N_4983,N_5149);
xnor U7802 (N_7802,N_5579,N_5019);
nand U7803 (N_7803,N_4608,N_4564);
nand U7804 (N_7804,N_5261,N_4387);
or U7805 (N_7805,N_5623,N_5909);
and U7806 (N_7806,N_5164,N_4563);
and U7807 (N_7807,N_4813,N_5583);
xor U7808 (N_7808,N_5498,N_5067);
xor U7809 (N_7809,N_4266,N_5383);
nand U7810 (N_7810,N_4555,N_4067);
nand U7811 (N_7811,N_5555,N_5135);
nor U7812 (N_7812,N_4635,N_5067);
and U7813 (N_7813,N_4456,N_5945);
or U7814 (N_7814,N_5209,N_5660);
xor U7815 (N_7815,N_5383,N_4864);
and U7816 (N_7816,N_4867,N_4900);
nand U7817 (N_7817,N_5009,N_4130);
nor U7818 (N_7818,N_4493,N_5722);
nand U7819 (N_7819,N_4083,N_5215);
nor U7820 (N_7820,N_5501,N_5962);
or U7821 (N_7821,N_5020,N_5540);
xnor U7822 (N_7822,N_4951,N_5141);
nor U7823 (N_7823,N_4905,N_4969);
xor U7824 (N_7824,N_4603,N_5938);
nor U7825 (N_7825,N_4046,N_5850);
nor U7826 (N_7826,N_4853,N_5363);
xnor U7827 (N_7827,N_5408,N_4679);
nor U7828 (N_7828,N_4961,N_5589);
and U7829 (N_7829,N_5892,N_4384);
xnor U7830 (N_7830,N_4870,N_5637);
or U7831 (N_7831,N_4529,N_5599);
or U7832 (N_7832,N_4569,N_5764);
and U7833 (N_7833,N_4458,N_5720);
or U7834 (N_7834,N_4476,N_4751);
xnor U7835 (N_7835,N_5398,N_4495);
xnor U7836 (N_7836,N_4915,N_5919);
xor U7837 (N_7837,N_4788,N_5462);
and U7838 (N_7838,N_5565,N_5138);
xor U7839 (N_7839,N_5437,N_4195);
or U7840 (N_7840,N_4887,N_5975);
nand U7841 (N_7841,N_5848,N_4272);
nor U7842 (N_7842,N_5187,N_5695);
nand U7843 (N_7843,N_4661,N_4974);
or U7844 (N_7844,N_5551,N_4460);
or U7845 (N_7845,N_5020,N_4794);
xor U7846 (N_7846,N_5556,N_4612);
nor U7847 (N_7847,N_4061,N_4270);
and U7848 (N_7848,N_4737,N_4729);
or U7849 (N_7849,N_4996,N_5211);
nand U7850 (N_7850,N_5446,N_4938);
or U7851 (N_7851,N_5794,N_4574);
nand U7852 (N_7852,N_4103,N_5843);
and U7853 (N_7853,N_5406,N_4805);
nand U7854 (N_7854,N_5577,N_5223);
and U7855 (N_7855,N_4376,N_5995);
and U7856 (N_7856,N_5748,N_5331);
nor U7857 (N_7857,N_5978,N_5060);
nor U7858 (N_7858,N_5397,N_4040);
nand U7859 (N_7859,N_4790,N_5920);
or U7860 (N_7860,N_4357,N_5624);
nand U7861 (N_7861,N_4539,N_5579);
xor U7862 (N_7862,N_4289,N_5474);
xor U7863 (N_7863,N_4621,N_4853);
nand U7864 (N_7864,N_5858,N_4497);
or U7865 (N_7865,N_5959,N_4903);
xnor U7866 (N_7866,N_5528,N_4367);
nand U7867 (N_7867,N_4323,N_5592);
nor U7868 (N_7868,N_4623,N_4143);
and U7869 (N_7869,N_5125,N_5954);
and U7870 (N_7870,N_5840,N_4496);
or U7871 (N_7871,N_4319,N_5266);
xor U7872 (N_7872,N_5955,N_5115);
nor U7873 (N_7873,N_5203,N_4782);
or U7874 (N_7874,N_4479,N_5262);
nand U7875 (N_7875,N_4812,N_4067);
nand U7876 (N_7876,N_5984,N_5321);
xnor U7877 (N_7877,N_4056,N_5009);
or U7878 (N_7878,N_4572,N_5525);
or U7879 (N_7879,N_5732,N_5546);
nor U7880 (N_7880,N_4877,N_5811);
and U7881 (N_7881,N_5023,N_5324);
and U7882 (N_7882,N_4681,N_4080);
xnor U7883 (N_7883,N_4305,N_5198);
or U7884 (N_7884,N_5832,N_5615);
xnor U7885 (N_7885,N_4959,N_5891);
xnor U7886 (N_7886,N_5424,N_5871);
and U7887 (N_7887,N_5886,N_5999);
nand U7888 (N_7888,N_5547,N_5116);
nor U7889 (N_7889,N_5185,N_5038);
and U7890 (N_7890,N_4887,N_4893);
nor U7891 (N_7891,N_5359,N_4050);
nand U7892 (N_7892,N_4432,N_5711);
nor U7893 (N_7893,N_5797,N_4509);
or U7894 (N_7894,N_5740,N_4231);
nand U7895 (N_7895,N_4560,N_5588);
nand U7896 (N_7896,N_5915,N_5495);
or U7897 (N_7897,N_4617,N_5667);
nand U7898 (N_7898,N_5433,N_5683);
nor U7899 (N_7899,N_4538,N_5636);
and U7900 (N_7900,N_4493,N_5332);
or U7901 (N_7901,N_5448,N_4749);
xnor U7902 (N_7902,N_5465,N_5444);
or U7903 (N_7903,N_5650,N_4600);
xor U7904 (N_7904,N_4389,N_4017);
or U7905 (N_7905,N_5734,N_5852);
and U7906 (N_7906,N_5958,N_5297);
and U7907 (N_7907,N_5162,N_5463);
nand U7908 (N_7908,N_4166,N_5068);
or U7909 (N_7909,N_5021,N_5010);
or U7910 (N_7910,N_5322,N_4238);
xor U7911 (N_7911,N_5780,N_4310);
or U7912 (N_7912,N_5062,N_4986);
or U7913 (N_7913,N_4890,N_4799);
and U7914 (N_7914,N_5509,N_4370);
or U7915 (N_7915,N_4095,N_4411);
xor U7916 (N_7916,N_5702,N_4603);
or U7917 (N_7917,N_4400,N_5138);
nor U7918 (N_7918,N_5406,N_4173);
and U7919 (N_7919,N_4505,N_4153);
and U7920 (N_7920,N_5845,N_5606);
and U7921 (N_7921,N_4798,N_5796);
xnor U7922 (N_7922,N_5428,N_4456);
and U7923 (N_7923,N_5259,N_5997);
xor U7924 (N_7924,N_4394,N_4759);
nor U7925 (N_7925,N_4524,N_4136);
nand U7926 (N_7926,N_5145,N_5959);
nand U7927 (N_7927,N_4239,N_4556);
nor U7928 (N_7928,N_5471,N_5818);
nor U7929 (N_7929,N_5006,N_4920);
nand U7930 (N_7930,N_4748,N_5363);
nor U7931 (N_7931,N_5316,N_5758);
and U7932 (N_7932,N_4709,N_5582);
or U7933 (N_7933,N_5792,N_5634);
and U7934 (N_7934,N_5122,N_5784);
xor U7935 (N_7935,N_5850,N_4885);
and U7936 (N_7936,N_4181,N_5661);
or U7937 (N_7937,N_4619,N_4668);
or U7938 (N_7938,N_4456,N_5563);
and U7939 (N_7939,N_4778,N_5186);
and U7940 (N_7940,N_4200,N_4954);
or U7941 (N_7941,N_4637,N_5126);
nor U7942 (N_7942,N_4883,N_5353);
nand U7943 (N_7943,N_4707,N_5424);
or U7944 (N_7944,N_5902,N_5577);
xor U7945 (N_7945,N_4262,N_5606);
nand U7946 (N_7946,N_4433,N_4998);
and U7947 (N_7947,N_5514,N_5694);
or U7948 (N_7948,N_5346,N_4441);
xnor U7949 (N_7949,N_4770,N_5063);
nor U7950 (N_7950,N_5276,N_5697);
nand U7951 (N_7951,N_5000,N_4930);
and U7952 (N_7952,N_4189,N_5319);
xnor U7953 (N_7953,N_5790,N_5311);
nor U7954 (N_7954,N_4142,N_4429);
or U7955 (N_7955,N_4542,N_5327);
xor U7956 (N_7956,N_5264,N_4051);
and U7957 (N_7957,N_4237,N_5700);
nor U7958 (N_7958,N_4378,N_5895);
nand U7959 (N_7959,N_4764,N_5923);
and U7960 (N_7960,N_5194,N_4688);
or U7961 (N_7961,N_5215,N_5325);
nand U7962 (N_7962,N_5000,N_5185);
nor U7963 (N_7963,N_5641,N_5604);
nand U7964 (N_7964,N_4309,N_5273);
nand U7965 (N_7965,N_5619,N_5587);
nor U7966 (N_7966,N_5558,N_4614);
and U7967 (N_7967,N_5456,N_5588);
and U7968 (N_7968,N_4543,N_5442);
nand U7969 (N_7969,N_4048,N_4927);
nand U7970 (N_7970,N_5753,N_4975);
xor U7971 (N_7971,N_4116,N_5540);
xor U7972 (N_7972,N_5567,N_4106);
xor U7973 (N_7973,N_4929,N_5456);
and U7974 (N_7974,N_4044,N_4820);
xor U7975 (N_7975,N_4956,N_5832);
nand U7976 (N_7976,N_5075,N_5755);
and U7977 (N_7977,N_5762,N_4243);
nor U7978 (N_7978,N_4789,N_5342);
nand U7979 (N_7979,N_4425,N_5942);
nor U7980 (N_7980,N_5099,N_5551);
nor U7981 (N_7981,N_4389,N_5390);
nand U7982 (N_7982,N_5772,N_4042);
nand U7983 (N_7983,N_5985,N_5025);
or U7984 (N_7984,N_4406,N_4670);
xnor U7985 (N_7985,N_5505,N_5663);
and U7986 (N_7986,N_4201,N_5559);
nand U7987 (N_7987,N_5930,N_5222);
nor U7988 (N_7988,N_4985,N_4783);
nor U7989 (N_7989,N_4186,N_4690);
and U7990 (N_7990,N_5474,N_5301);
nor U7991 (N_7991,N_4744,N_5290);
and U7992 (N_7992,N_5025,N_5446);
nand U7993 (N_7993,N_5443,N_5469);
nand U7994 (N_7994,N_4557,N_5261);
and U7995 (N_7995,N_4600,N_5699);
nand U7996 (N_7996,N_5478,N_4550);
or U7997 (N_7997,N_5037,N_5320);
or U7998 (N_7998,N_4010,N_5924);
or U7999 (N_7999,N_4060,N_4135);
xor U8000 (N_8000,N_6048,N_6254);
nand U8001 (N_8001,N_6098,N_6531);
and U8002 (N_8002,N_7364,N_7946);
or U8003 (N_8003,N_6508,N_7753);
nor U8004 (N_8004,N_6660,N_6308);
or U8005 (N_8005,N_7503,N_6776);
or U8006 (N_8006,N_7093,N_6699);
nor U8007 (N_8007,N_6831,N_7211);
or U8008 (N_8008,N_7852,N_7583);
xnor U8009 (N_8009,N_6779,N_7670);
and U8010 (N_8010,N_7728,N_7194);
xnor U8011 (N_8011,N_7202,N_7723);
and U8012 (N_8012,N_7338,N_6970);
nand U8013 (N_8013,N_6681,N_7128);
and U8014 (N_8014,N_6386,N_6871);
nand U8015 (N_8015,N_6244,N_7132);
nor U8016 (N_8016,N_6041,N_6951);
or U8017 (N_8017,N_6542,N_6469);
nand U8018 (N_8018,N_7501,N_7185);
nor U8019 (N_8019,N_7810,N_6275);
nand U8020 (N_8020,N_6309,N_6290);
xnor U8021 (N_8021,N_7689,N_7551);
or U8022 (N_8022,N_6197,N_7507);
xor U8023 (N_8023,N_6642,N_7573);
and U8024 (N_8024,N_6927,N_7001);
and U8025 (N_8025,N_7319,N_7172);
xnor U8026 (N_8026,N_6421,N_6032);
nor U8027 (N_8027,N_6043,N_7578);
or U8028 (N_8028,N_7966,N_6511);
xor U8029 (N_8029,N_7391,N_7531);
xor U8030 (N_8030,N_7295,N_6196);
and U8031 (N_8031,N_6759,N_7030);
nand U8032 (N_8032,N_6109,N_6390);
xnor U8033 (N_8033,N_6065,N_6519);
and U8034 (N_8034,N_6572,N_6015);
or U8035 (N_8035,N_7726,N_6441);
or U8036 (N_8036,N_7053,N_6600);
and U8037 (N_8037,N_7239,N_7684);
nor U8038 (N_8038,N_6371,N_6123);
nor U8039 (N_8039,N_7699,N_6412);
nor U8040 (N_8040,N_6881,N_7894);
nor U8041 (N_8041,N_6500,N_6852);
nor U8042 (N_8042,N_6712,N_7910);
nand U8043 (N_8043,N_6543,N_6935);
or U8044 (N_8044,N_6506,N_7525);
xor U8045 (N_8045,N_6557,N_7557);
and U8046 (N_8046,N_7809,N_7443);
and U8047 (N_8047,N_6992,N_6804);
or U8048 (N_8048,N_6830,N_7237);
or U8049 (N_8049,N_6757,N_7885);
or U8050 (N_8050,N_7775,N_7886);
nor U8051 (N_8051,N_7906,N_6171);
xor U8052 (N_8052,N_7440,N_7213);
and U8053 (N_8053,N_7203,N_6916);
nand U8054 (N_8054,N_6991,N_7609);
xor U8055 (N_8055,N_6869,N_6429);
or U8056 (N_8056,N_6633,N_6424);
nand U8057 (N_8057,N_6799,N_7173);
nor U8058 (N_8058,N_7368,N_7312);
xnor U8059 (N_8059,N_7511,N_7439);
and U8060 (N_8060,N_7066,N_7581);
xnor U8061 (N_8061,N_6083,N_6444);
nor U8062 (N_8062,N_6632,N_7940);
or U8063 (N_8063,N_7673,N_6057);
or U8064 (N_8064,N_7600,N_6217);
and U8065 (N_8065,N_7328,N_6369);
xnor U8066 (N_8066,N_7158,N_7057);
nor U8067 (N_8067,N_7624,N_6399);
nor U8068 (N_8068,N_7959,N_6184);
xor U8069 (N_8069,N_7831,N_7956);
nand U8070 (N_8070,N_7605,N_6857);
xor U8071 (N_8071,N_6661,N_6241);
and U8072 (N_8072,N_6853,N_7941);
xnor U8073 (N_8073,N_6398,N_6593);
nand U8074 (N_8074,N_7614,N_7550);
xnor U8075 (N_8075,N_7303,N_7954);
xor U8076 (N_8076,N_7655,N_7606);
nand U8077 (N_8077,N_6018,N_6204);
nor U8078 (N_8078,N_6476,N_6082);
and U8079 (N_8079,N_6218,N_6652);
xor U8080 (N_8080,N_6163,N_6605);
or U8081 (N_8081,N_6708,N_6868);
or U8082 (N_8082,N_7949,N_6368);
or U8083 (N_8083,N_7871,N_6775);
nor U8084 (N_8084,N_6351,N_7226);
or U8085 (N_8085,N_7963,N_6953);
nor U8086 (N_8086,N_7702,N_7496);
and U8087 (N_8087,N_7672,N_7932);
nor U8088 (N_8088,N_6603,N_6932);
xor U8089 (N_8089,N_6581,N_6122);
nand U8090 (N_8090,N_7739,N_7322);
and U8091 (N_8091,N_7462,N_7141);
xnor U8092 (N_8092,N_7031,N_7647);
and U8093 (N_8093,N_7039,N_7412);
nor U8094 (N_8094,N_6730,N_7792);
and U8095 (N_8095,N_6484,N_6293);
nor U8096 (N_8096,N_6934,N_6240);
nor U8097 (N_8097,N_6433,N_6694);
xnor U8098 (N_8098,N_6627,N_7323);
or U8099 (N_8099,N_7235,N_7341);
nor U8100 (N_8100,N_6099,N_6906);
and U8101 (N_8101,N_6613,N_6058);
or U8102 (N_8102,N_6013,N_7730);
nand U8103 (N_8103,N_7184,N_6489);
and U8104 (N_8104,N_6022,N_6522);
nand U8105 (N_8105,N_6372,N_6439);
and U8106 (N_8106,N_7196,N_7055);
nand U8107 (N_8107,N_6789,N_6588);
and U8108 (N_8108,N_7659,N_7408);
and U8109 (N_8109,N_7216,N_7283);
xnor U8110 (N_8110,N_7414,N_7528);
or U8111 (N_8111,N_7482,N_6385);
nand U8112 (N_8112,N_7160,N_6523);
xnor U8113 (N_8113,N_7253,N_6253);
nand U8114 (N_8114,N_6237,N_6216);
nor U8115 (N_8115,N_6527,N_7373);
nand U8116 (N_8116,N_7153,N_6479);
and U8117 (N_8117,N_6014,N_6987);
or U8118 (N_8118,N_6250,N_6135);
nor U8119 (N_8119,N_6639,N_7703);
nand U8120 (N_8120,N_7931,N_7288);
and U8121 (N_8121,N_7856,N_6400);
or U8122 (N_8122,N_6541,N_6726);
nand U8123 (N_8123,N_6635,N_7523);
or U8124 (N_8124,N_6822,N_7631);
or U8125 (N_8125,N_7428,N_6981);
nor U8126 (N_8126,N_6931,N_7526);
or U8127 (N_8127,N_7823,N_6446);
nor U8128 (N_8128,N_7637,N_6884);
nor U8129 (N_8129,N_6112,N_6379);
xor U8130 (N_8130,N_7367,N_6702);
or U8131 (N_8131,N_6282,N_7580);
xor U8132 (N_8132,N_7109,N_6644);
xnor U8133 (N_8133,N_6006,N_6791);
nor U8134 (N_8134,N_6937,N_7765);
or U8135 (N_8135,N_6658,N_7891);
xor U8136 (N_8136,N_6411,N_6289);
or U8137 (N_8137,N_6715,N_6454);
and U8138 (N_8138,N_6897,N_7467);
or U8139 (N_8139,N_7527,N_7760);
nand U8140 (N_8140,N_7603,N_6679);
or U8141 (N_8141,N_7187,N_7882);
and U8142 (N_8142,N_6481,N_6036);
nand U8143 (N_8143,N_7078,N_7320);
nand U8144 (N_8144,N_6363,N_7063);
and U8145 (N_8145,N_7261,N_7189);
xnor U8146 (N_8146,N_7192,N_6425);
xor U8147 (N_8147,N_6815,N_6521);
xor U8148 (N_8148,N_7926,N_6969);
nand U8149 (N_8149,N_7370,N_6885);
or U8150 (N_8150,N_7299,N_6374);
nor U8151 (N_8151,N_6535,N_7399);
or U8152 (N_8152,N_7460,N_6909);
nand U8153 (N_8153,N_7033,N_6315);
nor U8154 (N_8154,N_6248,N_6938);
or U8155 (N_8155,N_6066,N_6219);
or U8156 (N_8156,N_6895,N_6144);
and U8157 (N_8157,N_6553,N_7686);
xnor U8158 (N_8158,N_7964,N_7669);
nand U8159 (N_8159,N_7329,N_7282);
or U8160 (N_8160,N_7372,N_7738);
nor U8161 (N_8161,N_6415,N_7755);
nand U8162 (N_8162,N_7385,N_7072);
and U8163 (N_8163,N_6276,N_6138);
nand U8164 (N_8164,N_6811,N_7490);
nor U8165 (N_8165,N_6963,N_6306);
nor U8166 (N_8166,N_7150,N_7500);
and U8167 (N_8167,N_7445,N_6516);
nor U8168 (N_8168,N_7734,N_7131);
nor U8169 (N_8169,N_6222,N_7678);
nor U8170 (N_8170,N_6643,N_6915);
or U8171 (N_8171,N_7390,N_7756);
or U8172 (N_8172,N_6071,N_7725);
and U8173 (N_8173,N_7543,N_6806);
nand U8174 (N_8174,N_7514,N_6845);
or U8175 (N_8175,N_7137,N_7361);
nor U8176 (N_8176,N_7970,N_7575);
nor U8177 (N_8177,N_7204,N_7987);
xnor U8178 (N_8178,N_7444,N_6312);
nand U8179 (N_8179,N_7068,N_6837);
nand U8180 (N_8180,N_6698,N_6536);
nor U8181 (N_8181,N_6558,N_6188);
nor U8182 (N_8182,N_6512,N_7418);
and U8183 (N_8183,N_6227,N_6790);
nor U8184 (N_8184,N_7942,N_6157);
or U8185 (N_8185,N_7974,N_6550);
or U8186 (N_8186,N_6983,N_6338);
nand U8187 (N_8187,N_7263,N_6136);
or U8188 (N_8188,N_7981,N_7342);
or U8189 (N_8189,N_6464,N_6149);
and U8190 (N_8190,N_6105,N_7768);
or U8191 (N_8191,N_6313,N_7144);
or U8192 (N_8192,N_7247,N_6801);
or U8193 (N_8193,N_6703,N_7447);
or U8194 (N_8194,N_7667,N_6078);
or U8195 (N_8195,N_7294,N_6011);
nor U8196 (N_8196,N_6202,N_7973);
xnor U8197 (N_8197,N_7084,N_6753);
nor U8198 (N_8198,N_7876,N_6754);
nand U8199 (N_8199,N_7569,N_7874);
nand U8200 (N_8200,N_6731,N_7777);
or U8201 (N_8201,N_7957,N_7736);
xor U8202 (N_8202,N_7909,N_7661);
xnor U8203 (N_8203,N_7198,N_6445);
xnor U8204 (N_8204,N_6861,N_7094);
xor U8205 (N_8205,N_7555,N_6206);
nand U8206 (N_8206,N_7912,N_6628);
nor U8207 (N_8207,N_6354,N_7148);
and U8208 (N_8208,N_7893,N_6463);
nand U8209 (N_8209,N_6843,N_6169);
xnor U8210 (N_8210,N_6183,N_6957);
nand U8211 (N_8211,N_6457,N_7817);
xnor U8212 (N_8212,N_6346,N_6328);
and U8213 (N_8213,N_6540,N_6785);
nand U8214 (N_8214,N_7415,N_7748);
nor U8215 (N_8215,N_6323,N_7218);
or U8216 (N_8216,N_7830,N_6580);
nand U8217 (N_8217,N_6020,N_7025);
nor U8218 (N_8218,N_6209,N_7592);
and U8219 (N_8219,N_7091,N_7233);
xor U8220 (N_8220,N_7758,N_6419);
or U8221 (N_8221,N_7967,N_6849);
nor U8222 (N_8222,N_6740,N_6034);
nor U8223 (N_8223,N_7348,N_7197);
nor U8224 (N_8224,N_6033,N_7166);
or U8225 (N_8225,N_6575,N_7420);
xor U8226 (N_8226,N_6586,N_7664);
xnor U8227 (N_8227,N_6496,N_6824);
nand U8228 (N_8228,N_6195,N_7545);
nor U8229 (N_8229,N_6220,N_6173);
xor U8230 (N_8230,N_6159,N_7992);
nor U8231 (N_8231,N_7300,N_6504);
nor U8232 (N_8232,N_7163,N_7993);
or U8233 (N_8233,N_6755,N_6142);
or U8234 (N_8234,N_7741,N_7688);
nand U8235 (N_8235,N_7552,N_7200);
or U8236 (N_8236,N_7922,N_6859);
nand U8237 (N_8237,N_6744,N_7746);
or U8238 (N_8238,N_7847,N_6686);
or U8239 (N_8239,N_7881,N_7147);
xnor U8240 (N_8240,N_6554,N_6207);
xor U8241 (N_8241,N_6009,N_6460);
or U8242 (N_8242,N_7888,N_6391);
or U8243 (N_8243,N_6499,N_6345);
nor U8244 (N_8244,N_6274,N_7086);
or U8245 (N_8245,N_7654,N_6748);
xnor U8246 (N_8246,N_7138,N_6666);
or U8247 (N_8247,N_7921,N_7269);
nand U8248 (N_8248,N_7599,N_7409);
nor U8249 (N_8249,N_7617,N_6321);
and U8250 (N_8250,N_7896,N_6280);
or U8251 (N_8251,N_6692,N_7316);
nor U8252 (N_8252,N_6455,N_7508);
nor U8253 (N_8253,N_6729,N_6548);
xor U8254 (N_8254,N_7014,N_6839);
nor U8255 (N_8255,N_7230,N_7900);
and U8256 (N_8256,N_6080,N_7277);
xor U8257 (N_8257,N_6174,N_7690);
or U8258 (N_8258,N_7308,N_6828);
or U8259 (N_8259,N_7548,N_6711);
nor U8260 (N_8260,N_6515,N_6294);
nand U8261 (N_8261,N_6710,N_6816);
xnor U8262 (N_8262,N_7105,N_6084);
and U8263 (N_8263,N_7143,N_7584);
and U8264 (N_8264,N_6721,N_6514);
nand U8265 (N_8265,N_6150,N_6827);
and U8266 (N_8266,N_7972,N_6784);
nor U8267 (N_8267,N_6905,N_6417);
nand U8268 (N_8268,N_6212,N_7424);
nand U8269 (N_8269,N_7676,N_6055);
nor U8270 (N_8270,N_7089,N_7767);
nand U8271 (N_8271,N_7274,N_6768);
xnor U8272 (N_8272,N_6251,N_6292);
nor U8273 (N_8273,N_7707,N_6579);
and U8274 (N_8274,N_7793,N_7953);
nor U8275 (N_8275,N_7464,N_6560);
xnor U8276 (N_8276,N_6611,N_6162);
xnor U8277 (N_8277,N_6846,N_6085);
and U8278 (N_8278,N_6994,N_6304);
and U8279 (N_8279,N_6539,N_6555);
nor U8280 (N_8280,N_7556,N_6490);
xor U8281 (N_8281,N_6175,N_7701);
xnor U8282 (N_8282,N_7626,N_7924);
nand U8283 (N_8283,N_7687,N_7286);
nand U8284 (N_8284,N_7733,N_6273);
or U8285 (N_8285,N_6912,N_6279);
and U8286 (N_8286,N_6471,N_6623);
or U8287 (N_8287,N_7928,N_7165);
nor U8288 (N_8288,N_7457,N_7727);
xnor U8289 (N_8289,N_7589,N_6001);
nor U8290 (N_8290,N_7950,N_6567);
or U8291 (N_8291,N_7436,N_6630);
xor U8292 (N_8292,N_6876,N_6185);
and U8293 (N_8293,N_7630,N_6782);
nand U8294 (N_8294,N_6718,N_7759);
and U8295 (N_8295,N_7167,N_7877);
and U8296 (N_8296,N_6189,N_6622);
nand U8297 (N_8297,N_7821,N_7287);
nor U8298 (N_8298,N_7860,N_6862);
nand U8299 (N_8299,N_7280,N_6302);
nand U8300 (N_8300,N_7958,N_6821);
nand U8301 (N_8301,N_6311,N_6146);
or U8302 (N_8302,N_6355,N_6303);
nor U8303 (N_8303,N_6342,N_6920);
xor U8304 (N_8304,N_6589,N_6520);
xnor U8305 (N_8305,N_7404,N_7634);
xor U8306 (N_8306,N_6650,N_6160);
and U8307 (N_8307,N_7681,N_7351);
nand U8308 (N_8308,N_7773,N_6509);
nand U8309 (N_8309,N_7214,N_7657);
nor U8310 (N_8310,N_7506,N_7849);
or U8311 (N_8311,N_7547,N_6074);
nor U8312 (N_8312,N_6148,N_6077);
xnor U8313 (N_8313,N_7538,N_6413);
nor U8314 (N_8314,N_6025,N_7903);
xor U8315 (N_8315,N_6239,N_7383);
nor U8316 (N_8316,N_6724,N_6349);
nand U8317 (N_8317,N_7417,N_6854);
nor U8318 (N_8318,N_6187,N_7859);
and U8319 (N_8319,N_7176,N_7222);
nand U8320 (N_8320,N_6118,N_6676);
xnor U8321 (N_8321,N_6996,N_7021);
and U8322 (N_8322,N_7292,N_7721);
nand U8323 (N_8323,N_6813,N_6335);
and U8324 (N_8324,N_7996,N_7816);
or U8325 (N_8325,N_7246,N_6477);
nand U8326 (N_8326,N_7455,N_6752);
nor U8327 (N_8327,N_6941,N_6794);
nor U8328 (N_8328,N_6127,N_7095);
and U8329 (N_8329,N_6634,N_7757);
or U8330 (N_8330,N_7593,N_7016);
or U8331 (N_8331,N_6761,N_7199);
nand U8332 (N_8332,N_7825,N_6738);
or U8333 (N_8333,N_7154,N_6551);
nor U8334 (N_8334,N_6917,N_7914);
and U8335 (N_8335,N_7771,N_7435);
or U8336 (N_8336,N_6975,N_6964);
or U8337 (N_8337,N_7518,N_7375);
nor U8338 (N_8338,N_6422,N_7930);
nand U8339 (N_8339,N_6384,N_6673);
xor U8340 (N_8340,N_7056,N_7358);
nand U8341 (N_8341,N_6322,N_7245);
and U8342 (N_8342,N_6326,N_6448);
xor U8343 (N_8343,N_6111,N_6832);
nor U8344 (N_8344,N_6904,N_7179);
nand U8345 (N_8345,N_7427,N_6907);
or U8346 (N_8346,N_7011,N_7118);
and U8347 (N_8347,N_7708,N_7713);
or U8348 (N_8348,N_6672,N_6119);
xor U8349 (N_8349,N_6818,N_7010);
and U8350 (N_8350,N_6267,N_7944);
nor U8351 (N_8351,N_7836,N_6974);
nor U8352 (N_8352,N_7868,N_6662);
or U8353 (N_8353,N_6224,N_7359);
and U8354 (N_8354,N_6392,N_7662);
nand U8355 (N_8355,N_6780,N_7763);
and U8356 (N_8356,N_6924,N_7977);
nand U8357 (N_8357,N_6106,N_6751);
or U8358 (N_8358,N_6973,N_6362);
xnor U8359 (N_8359,N_7971,N_6493);
and U8360 (N_8360,N_7572,N_6552);
nor U8361 (N_8361,N_7613,N_6898);
xnor U8362 (N_8362,N_6121,N_6353);
nand U8363 (N_8363,N_6747,N_7934);
xnor U8364 (N_8364,N_6668,N_6430);
nand U8365 (N_8365,N_7933,N_6366);
nand U8366 (N_8366,N_6327,N_6096);
nor U8367 (N_8367,N_6378,N_6796);
or U8368 (N_8368,N_7157,N_6023);
or U8369 (N_8369,N_6468,N_7054);
xnor U8370 (N_8370,N_7382,N_6842);
xor U8371 (N_8371,N_6962,N_6295);
or U8372 (N_8372,N_6826,N_6598);
nand U8373 (N_8373,N_7558,N_7422);
and U8374 (N_8374,N_7486,N_7048);
and U8375 (N_8375,N_6235,N_7706);
xor U8376 (N_8376,N_6793,N_6069);
and U8377 (N_8377,N_6246,N_6005);
nand U8378 (N_8378,N_7497,N_6918);
xor U8379 (N_8379,N_7622,N_7652);
and U8380 (N_8380,N_6654,N_6638);
nor U8381 (N_8381,N_6670,N_7908);
or U8382 (N_8382,N_6517,N_6976);
nor U8383 (N_8383,N_6781,N_6788);
nand U8384 (N_8384,N_7369,N_7715);
or U8385 (N_8385,N_6381,N_6997);
and U8386 (N_8386,N_6172,N_7310);
or U8387 (N_8387,N_6875,N_7272);
xor U8388 (N_8388,N_7752,N_6812);
and U8389 (N_8389,N_7178,N_7059);
nand U8390 (N_8390,N_7978,N_6902);
or U8391 (N_8391,N_6263,N_7695);
nand U8392 (N_8392,N_7587,N_6000);
and U8393 (N_8393,N_7394,N_7772);
xnor U8394 (N_8394,N_7122,N_6010);
xnor U8395 (N_8395,N_7850,N_7018);
nand U8396 (N_8396,N_6954,N_6961);
nor U8397 (N_8397,N_6134,N_6525);
nor U8398 (N_8398,N_6467,N_7350);
nand U8399 (N_8399,N_7719,N_7110);
xor U8400 (N_8400,N_6442,N_6595);
nand U8401 (N_8401,N_7330,N_7162);
and U8402 (N_8402,N_7883,N_7190);
or U8403 (N_8403,N_7549,N_6193);
nand U8404 (N_8404,N_7139,N_7212);
xnor U8405 (N_8405,N_7510,N_7857);
nor U8406 (N_8406,N_7623,N_7466);
nor U8407 (N_8407,N_7660,N_7803);
nor U8408 (N_8408,N_7535,N_6984);
nand U8409 (N_8409,N_7618,N_7374);
xor U8410 (N_8410,N_6361,N_7854);
and U8411 (N_8411,N_6538,N_6110);
nand U8412 (N_8412,N_6200,N_6310);
or U8413 (N_8413,N_7480,N_7539);
xor U8414 (N_8414,N_7743,N_7749);
nor U8415 (N_8415,N_7419,N_7872);
or U8416 (N_8416,N_6225,N_7136);
nor U8417 (N_8417,N_7125,N_7402);
xnor U8418 (N_8418,N_6044,N_7515);
xor U8419 (N_8419,N_7103,N_7430);
and U8420 (N_8420,N_7516,N_7468);
nor U8421 (N_8421,N_6408,N_7306);
xnor U8422 (N_8422,N_7629,N_6039);
xor U8423 (N_8423,N_6230,N_6395);
xor U8424 (N_8424,N_6810,N_6233);
or U8425 (N_8425,N_7357,N_7437);
xnor U8426 (N_8426,N_6440,N_6647);
nand U8427 (N_8427,N_6943,N_6696);
and U8428 (N_8428,N_6375,N_7834);
xnor U8429 (N_8429,N_7380,N_7285);
nor U8430 (N_8430,N_7879,N_6436);
nor U8431 (N_8431,N_6456,N_7149);
xnor U8432 (N_8432,N_7858,N_6277);
nor U8433 (N_8433,N_6985,N_7791);
nand U8434 (N_8434,N_7754,N_6305);
nor U8435 (N_8435,N_6617,N_7298);
and U8436 (N_8436,N_7193,N_6107);
nand U8437 (N_8437,N_6850,N_6719);
or U8438 (N_8438,N_6571,N_6940);
nor U8439 (N_8439,N_7229,N_6566);
or U8440 (N_8440,N_6215,N_7258);
nand U8441 (N_8441,N_7938,N_7015);
nor U8442 (N_8442,N_6689,N_7887);
nor U8443 (N_8443,N_7260,N_7164);
xnor U8444 (N_8444,N_7223,N_6618);
or U8445 (N_8445,N_6671,N_7371);
xnor U8446 (N_8446,N_7123,N_7766);
and U8447 (N_8447,N_6234,N_7619);
nor U8448 (N_8448,N_7340,N_7249);
xnor U8449 (N_8449,N_7902,N_7898);
and U8450 (N_8450,N_6021,N_6108);
or U8451 (N_8451,N_6097,N_6663);
or U8452 (N_8452,N_6872,N_6620);
nand U8453 (N_8453,N_7512,N_6347);
or U8454 (N_8454,N_7919,N_6129);
nor U8455 (N_8455,N_6942,N_7379);
and U8456 (N_8456,N_6046,N_6388);
xnor U8457 (N_8457,N_6578,N_6995);
and U8458 (N_8458,N_6367,N_7504);
and U8459 (N_8459,N_6948,N_6067);
xor U8460 (N_8460,N_6704,N_6319);
or U8461 (N_8461,N_7234,N_7724);
and U8462 (N_8462,N_7566,N_7776);
and U8463 (N_8463,N_6356,N_6405);
nor U8464 (N_8464,N_6194,N_7171);
or U8465 (N_8465,N_7916,N_7597);
xnor U8466 (N_8466,N_6570,N_7406);
nor U8467 (N_8467,N_7281,N_7215);
xor U8468 (N_8468,N_7737,N_7029);
xor U8469 (N_8469,N_7041,N_6092);
and U8470 (N_8470,N_6858,N_6573);
nand U8471 (N_8471,N_6133,N_6452);
and U8472 (N_8472,N_7080,N_6051);
nand U8473 (N_8473,N_7668,N_7636);
or U8474 (N_8474,N_7022,N_7352);
nor U8475 (N_8475,N_7180,N_7458);
nand U8476 (N_8476,N_7806,N_6547);
and U8477 (N_8477,N_6063,N_6762);
xnor U8478 (N_8478,N_6177,N_7135);
xnor U8479 (N_8479,N_7905,N_6528);
nor U8480 (N_8480,N_7666,N_6585);
nand U8481 (N_8481,N_7889,N_7241);
xnor U8482 (N_8482,N_6393,N_7311);
nand U8483 (N_8483,N_7988,N_7704);
nand U8484 (N_8484,N_7851,N_7610);
nor U8485 (N_8485,N_7307,N_6583);
nand U8486 (N_8486,N_7665,N_6896);
xor U8487 (N_8487,N_6431,N_7360);
or U8488 (N_8488,N_6377,N_6409);
and U8489 (N_8489,N_7778,N_6829);
nand U8490 (N_8490,N_6178,N_6923);
nand U8491 (N_8491,N_7291,N_6114);
or U8492 (N_8492,N_6736,N_6590);
or U8493 (N_8493,N_7807,N_6803);
xnor U8494 (N_8494,N_7431,N_6944);
and U8495 (N_8495,N_7265,N_6714);
and U8496 (N_8496,N_6153,N_6472);
nor U8497 (N_8497,N_7864,N_7519);
or U8498 (N_8498,N_6154,N_6814);
nand U8499 (N_8499,N_6383,N_6268);
and U8500 (N_8500,N_7602,N_6285);
nor U8501 (N_8501,N_7451,N_6126);
xor U8502 (N_8502,N_6317,N_7867);
nand U8503 (N_8503,N_7590,N_6680);
xnor U8504 (N_8504,N_7009,N_6802);
or U8505 (N_8505,N_7301,N_7786);
nor U8506 (N_8506,N_6038,N_6836);
or U8507 (N_8507,N_6394,N_6257);
xnor U8508 (N_8508,N_6914,N_6059);
xnor U8509 (N_8509,N_7477,N_7546);
or U8510 (N_8510,N_6339,N_7070);
xnor U8511 (N_8511,N_6825,N_6298);
nor U8512 (N_8512,N_7835,N_6908);
nand U8513 (N_8513,N_7465,N_7663);
xor U8514 (N_8514,N_7049,N_6877);
and U8515 (N_8515,N_6002,N_6086);
or U8516 (N_8516,N_7483,N_7815);
nor U8517 (N_8517,N_6518,N_6229);
nand U8518 (N_8518,N_6743,N_7248);
nand U8519 (N_8519,N_6820,N_6320);
xor U8520 (N_8520,N_7985,N_7327);
and U8521 (N_8521,N_6161,N_7146);
nand U8522 (N_8522,N_7052,N_7188);
or U8523 (N_8523,N_6494,N_6631);
and U8524 (N_8524,N_6420,N_6988);
and U8525 (N_8525,N_6270,N_6259);
nand U8526 (N_8526,N_6855,N_7114);
and U8527 (N_8527,N_7750,N_7717);
nand U8528 (N_8528,N_6769,N_7762);
nand U8529 (N_8529,N_6636,N_6949);
or U8530 (N_8530,N_7043,N_7986);
xnor U8531 (N_8531,N_7452,N_7220);
and U8532 (N_8532,N_7264,N_6664);
or U8533 (N_8533,N_7680,N_6928);
and U8534 (N_8534,N_7521,N_7096);
and U8535 (N_8535,N_7073,N_7488);
or U8536 (N_8536,N_7120,N_6221);
and U8537 (N_8537,N_6749,N_7062);
xnor U8538 (N_8538,N_7820,N_6507);
and U8539 (N_8539,N_7788,N_6199);
or U8540 (N_8540,N_6333,N_7082);
or U8541 (N_8541,N_7983,N_7632);
and U8542 (N_8542,N_6596,N_6348);
xnor U8543 (N_8543,N_7487,N_7064);
nor U8544 (N_8544,N_7611,N_6616);
xor U8545 (N_8545,N_6584,N_6675);
and U8546 (N_8546,N_6370,N_6795);
or U8547 (N_8547,N_7897,N_7008);
nand U8548 (N_8548,N_6739,N_6307);
and U8549 (N_8549,N_6458,N_7804);
nor U8550 (N_8550,N_7648,N_7875);
xor U8551 (N_8551,N_6637,N_7601);
nor U8552 (N_8552,N_6690,N_6880);
nor U8553 (N_8553,N_7712,N_6903);
nor U8554 (N_8554,N_6296,N_7892);
nor U8555 (N_8555,N_6054,N_6343);
nor U8556 (N_8556,N_6669,N_7494);
xor U8557 (N_8557,N_6863,N_6756);
xor U8558 (N_8558,N_6407,N_6688);
nand U8559 (N_8559,N_6532,N_6324);
or U8560 (N_8560,N_6745,N_7042);
or U8561 (N_8561,N_6856,N_6255);
or U8562 (N_8562,N_7051,N_6443);
and U8563 (N_8563,N_7939,N_6640);
nand U8564 (N_8564,N_6545,N_7735);
nor U8565 (N_8565,N_7396,N_7517);
xor U8566 (N_8566,N_7522,N_7585);
and U8567 (N_8567,N_7976,N_7720);
or U8568 (N_8568,N_6029,N_7305);
nor U8569 (N_8569,N_6592,N_6723);
nand U8570 (N_8570,N_7076,N_7947);
nor U8571 (N_8571,N_6428,N_7671);
or U8572 (N_8572,N_7377,N_6337);
or U8573 (N_8573,N_6765,N_7034);
and U8574 (N_8574,N_6607,N_6291);
nand U8575 (N_8575,N_6297,N_6451);
xor U8576 (N_8576,N_7498,N_7353);
nor U8577 (N_8577,N_6152,N_7331);
and U8578 (N_8578,N_7644,N_7782);
nor U8579 (N_8579,N_6722,N_7012);
and U8580 (N_8580,N_6040,N_7313);
nor U8581 (N_8581,N_7191,N_6807);
nor U8582 (N_8582,N_6725,N_7115);
xor U8583 (N_8583,N_7975,N_6380);
and U8584 (N_8584,N_7255,N_7347);
xor U8585 (N_8585,N_7221,N_7795);
or U8586 (N_8586,N_7832,N_7675);
and U8587 (N_8587,N_7783,N_7819);
xnor U8588 (N_8588,N_6890,N_7266);
nor U8589 (N_8589,N_7761,N_6288);
or U8590 (N_8590,N_7927,N_6261);
nand U8591 (N_8591,N_7175,N_7079);
or U8592 (N_8592,N_6564,N_6485);
xor U8593 (N_8593,N_7530,N_6659);
xor U8594 (N_8594,N_6042,N_6252);
and U8595 (N_8595,N_6396,N_7426);
xnor U8596 (N_8596,N_6565,N_7037);
nand U8597 (N_8597,N_6882,N_7254);
xnor U8598 (N_8598,N_6950,N_7334);
xor U8599 (N_8599,N_6266,N_7582);
nor U8600 (N_8600,N_6960,N_7764);
and U8601 (N_8601,N_7344,N_6534);
or U8602 (N_8602,N_7002,N_6750);
nand U8603 (N_8603,N_7709,N_7491);
nor U8604 (N_8604,N_6655,N_7965);
nor U8605 (N_8605,N_7813,N_7398);
nand U8606 (N_8606,N_7024,N_7088);
xnor U8607 (N_8607,N_6687,N_6783);
nor U8608 (N_8608,N_7047,N_6674);
nand U8609 (N_8609,N_6733,N_6648);
xnor U8610 (N_8610,N_6678,N_7509);
nand U8611 (N_8611,N_7895,N_6474);
and U8612 (N_8612,N_7290,N_7421);
and U8613 (N_8613,N_6502,N_7060);
and U8614 (N_8614,N_6569,N_6283);
xnor U8615 (N_8615,N_6382,N_7799);
or U8616 (N_8616,N_7607,N_6488);
or U8617 (N_8617,N_6300,N_7354);
or U8618 (N_8618,N_6088,N_7827);
nand U8619 (N_8619,N_6562,N_7107);
or U8620 (N_8620,N_6478,N_7499);
or U8621 (N_8621,N_7092,N_6865);
nand U8622 (N_8622,N_6281,N_6264);
and U8623 (N_8623,N_6475,N_6693);
xor U8624 (N_8624,N_6213,N_6125);
nand U8625 (N_8625,N_7729,N_7805);
xnor U8626 (N_8626,N_7217,N_7744);
xor U8627 (N_8627,N_7917,N_6864);
nor U8628 (N_8628,N_6075,N_7711);
xor U8629 (N_8629,N_7638,N_7411);
or U8630 (N_8630,N_7273,N_7007);
nand U8631 (N_8631,N_6977,N_7325);
xnor U8632 (N_8632,N_6945,N_7410);
and U8633 (N_8633,N_6624,N_6758);
or U8634 (N_8634,N_7270,N_7124);
or U8635 (N_8635,N_6007,N_7127);
or U8636 (N_8636,N_7085,N_7450);
and U8637 (N_8637,N_6851,N_6685);
nor U8638 (N_8638,N_7461,N_6402);
nand U8639 (N_8639,N_6103,N_7997);
nor U8640 (N_8640,N_7802,N_6434);
nand U8641 (N_8641,N_7979,N_7685);
nor U8642 (N_8642,N_7446,N_7075);
xor U8643 (N_8643,N_6120,N_7873);
nor U8644 (N_8644,N_6410,N_7478);
nor U8645 (N_8645,N_7126,N_7279);
and U8646 (N_8646,N_7740,N_6272);
xor U8647 (N_8647,N_7918,N_6269);
nand U8648 (N_8648,N_6979,N_7769);
or U8649 (N_8649,N_7284,N_6094);
nor U8650 (N_8650,N_7633,N_6993);
nand U8651 (N_8651,N_6626,N_6510);
or U8652 (N_8652,N_7395,N_7824);
nor U8653 (N_8653,N_7505,N_6012);
nor U8654 (N_8654,N_6887,N_6093);
nand U8655 (N_8655,N_6284,N_7537);
xnor U8656 (N_8656,N_6615,N_6968);
nand U8657 (N_8657,N_6764,N_7534);
xnor U8658 (N_8658,N_7159,N_7393);
xnor U8659 (N_8659,N_6141,N_7563);
or U8660 (N_8660,N_6767,N_6697);
and U8661 (N_8661,N_6318,N_7745);
xor U8662 (N_8662,N_7969,N_6683);
and U8663 (N_8663,N_6840,N_6608);
and U8664 (N_8664,N_7065,N_7948);
and U8665 (N_8665,N_7700,N_7968);
or U8666 (N_8666,N_6665,N_6364);
nor U8667 (N_8667,N_7425,N_7524);
xnor U8668 (N_8668,N_7787,N_7318);
and U8669 (N_8669,N_7267,N_6530);
nor U8670 (N_8670,N_7111,N_7692);
nand U8671 (N_8671,N_7335,N_7219);
and U8672 (N_8672,N_6910,N_6205);
xor U8673 (N_8673,N_7628,N_7026);
or U8674 (N_8674,N_6947,N_7116);
or U8675 (N_8675,N_7208,N_7870);
nor U8676 (N_8676,N_7275,N_7920);
and U8677 (N_8677,N_6190,N_6492);
nor U8678 (N_8678,N_6728,N_6889);
and U8679 (N_8679,N_6331,N_6359);
xor U8680 (N_8680,N_7625,N_6024);
nand U8681 (N_8681,N_6486,N_7168);
or U8682 (N_8682,N_6437,N_6705);
nor U8683 (N_8683,N_6893,N_6878);
or U8684 (N_8684,N_7271,N_6980);
xor U8685 (N_8685,N_6867,N_7564);
xor U8686 (N_8686,N_7540,N_7077);
xor U8687 (N_8687,N_6913,N_7098);
and U8688 (N_8688,N_7243,N_6168);
nor U8689 (N_8689,N_7794,N_7035);
nand U8690 (N_8690,N_7841,N_7598);
nor U8691 (N_8691,N_7710,N_6062);
or U8692 (N_8692,N_6900,N_6208);
or U8693 (N_8693,N_7321,N_7826);
or U8694 (N_8694,N_6971,N_6805);
and U8695 (N_8695,N_6577,N_6432);
xor U8696 (N_8696,N_7784,N_6834);
nand U8697 (N_8697,N_6329,N_6952);
nor U8698 (N_8698,N_7183,N_6866);
nand U8699 (N_8699,N_6053,N_7554);
or U8700 (N_8700,N_7134,N_7454);
or U8701 (N_8701,N_7800,N_6888);
and U8702 (N_8702,N_6770,N_6008);
nor U8703 (N_8703,N_6130,N_7475);
nand U8704 (N_8704,N_6495,N_7129);
and U8705 (N_8705,N_6344,N_7541);
xor U8706 (N_8706,N_6621,N_7389);
xor U8707 (N_8707,N_6503,N_7502);
xnor U8708 (N_8708,N_7653,N_7586);
or U8709 (N_8709,N_7960,N_6373);
or U8710 (N_8710,N_6186,N_6035);
and U8711 (N_8711,N_6165,N_7346);
and U8712 (N_8712,N_6145,N_7570);
xor U8713 (N_8713,N_6223,N_6143);
or U8714 (N_8714,N_7268,N_6226);
nand U8715 (N_8715,N_7317,N_7493);
nor U8716 (N_8716,N_6079,N_7403);
xor U8717 (N_8717,N_7544,N_7438);
and U8718 (N_8718,N_6480,N_6965);
nor U8719 (N_8719,N_6073,N_6271);
and U8720 (N_8720,N_7961,N_7413);
nand U8721 (N_8721,N_7036,N_6247);
nor U8722 (N_8722,N_7209,N_7441);
nor U8723 (N_8723,N_6966,N_7182);
xnor U8724 (N_8724,N_7365,N_6823);
nor U8725 (N_8725,N_6017,N_7595);
or U8726 (N_8726,N_7067,N_7170);
nor U8727 (N_8727,N_6228,N_7145);
and U8728 (N_8728,N_6181,N_6706);
nor U8729 (N_8729,N_7995,N_6684);
nor U8730 (N_8730,N_7913,N_6883);
xor U8731 (N_8731,N_7696,N_6591);
and U8732 (N_8732,N_6449,N_7206);
nor U8733 (N_8733,N_6929,N_6990);
or U8734 (N_8734,N_7100,N_6537);
nand U8735 (N_8735,N_7574,N_6314);
xnor U8736 (N_8736,N_7463,N_7651);
nand U8737 (N_8737,N_7032,N_7207);
or U8738 (N_8738,N_6606,N_7152);
or U8739 (N_8739,N_7829,N_6334);
and U8740 (N_8740,N_7174,N_6068);
and U8741 (N_8741,N_7416,N_6482);
nand U8742 (N_8742,N_7257,N_6462);
or U8743 (N_8743,N_6604,N_6989);
or U8744 (N_8744,N_6848,N_6700);
nor U8745 (N_8745,N_6104,N_6653);
or U8746 (N_8746,N_6056,N_6091);
or U8747 (N_8747,N_7492,N_7104);
or U8748 (N_8748,N_7484,N_6438);
xor U8749 (N_8749,N_7658,N_7345);
nand U8750 (N_8750,N_7945,N_7117);
xnor U8751 (N_8751,N_7231,N_7576);
or U8752 (N_8752,N_6265,N_7381);
nand U8753 (N_8753,N_6179,N_7615);
nand U8754 (N_8754,N_7040,N_6967);
nand U8755 (N_8755,N_6360,N_7151);
xnor U8756 (N_8756,N_6180,N_6198);
or U8757 (N_8757,N_7336,N_7225);
and U8758 (N_8758,N_6132,N_7101);
nor U8759 (N_8759,N_7013,N_7113);
nand U8760 (N_8760,N_7865,N_7181);
and U8761 (N_8761,N_7855,N_6365);
or U8762 (N_8762,N_7304,N_7674);
nand U8763 (N_8763,N_7050,N_7027);
nand U8764 (N_8764,N_6958,N_7201);
nor U8765 (N_8765,N_6115,N_6026);
and U8766 (N_8766,N_6427,N_6879);
or U8767 (N_8767,N_6513,N_6524);
nor U8768 (N_8768,N_6899,N_6497);
nand U8769 (N_8769,N_7627,N_7228);
and U8770 (N_8770,N_6030,N_7384);
nor U8771 (N_8771,N_6072,N_6844);
and U8772 (N_8772,N_7513,N_6657);
nor U8773 (N_8773,N_6833,N_7560);
nor U8774 (N_8774,N_6336,N_6397);
and U8775 (N_8775,N_6746,N_6972);
or U8776 (N_8776,N_7161,N_6860);
nand U8777 (N_8777,N_7293,N_7878);
xor U8778 (N_8778,N_7639,N_7133);
xor U8779 (N_8779,N_6211,N_6325);
or U8780 (N_8780,N_7520,N_7751);
or U8781 (N_8781,N_6619,N_6352);
xnor U8782 (N_8782,N_7332,N_7276);
xor U8783 (N_8783,N_6771,N_6978);
nand U8784 (N_8784,N_7980,N_6709);
nor U8785 (N_8785,N_7612,N_7789);
nor U8786 (N_8786,N_7326,N_7044);
xnor U8787 (N_8787,N_7747,N_7296);
xor U8788 (N_8788,N_7904,N_6610);
xnor U8789 (N_8789,N_6599,N_6921);
xnor U8790 (N_8790,N_7577,N_7087);
or U8791 (N_8791,N_6919,N_6695);
xnor U8792 (N_8792,N_7697,N_7366);
and U8793 (N_8793,N_7349,N_6090);
nand U8794 (N_8794,N_7797,N_7814);
or U8795 (N_8795,N_6742,N_7923);
nand U8796 (N_8796,N_7387,N_6629);
xnor U8797 (N_8797,N_7474,N_6016);
nand U8798 (N_8798,N_6498,N_7679);
xor U8799 (N_8799,N_7568,N_6156);
nor U8800 (N_8800,N_6933,N_7236);
or U8801 (N_8801,N_6278,N_6050);
nor U8802 (N_8802,N_7925,N_6332);
nand U8803 (N_8803,N_7620,N_6113);
nand U8804 (N_8804,N_6998,N_6691);
nor U8805 (N_8805,N_7000,N_7102);
nor U8806 (N_8806,N_7432,N_7837);
xor U8807 (N_8807,N_7845,N_7650);
and U8808 (N_8808,N_7407,N_7028);
and U8809 (N_8809,N_6260,N_7691);
nor U8810 (N_8810,N_6701,N_7884);
nor U8811 (N_8811,N_6625,N_7473);
xnor U8812 (N_8812,N_6299,N_7812);
nand U8813 (N_8813,N_6004,N_6151);
xor U8814 (N_8814,N_7297,N_6101);
or U8815 (N_8815,N_7869,N_7459);
nand U8816 (N_8816,N_6649,N_6819);
nor U8817 (N_8817,N_6238,N_7561);
or U8818 (N_8818,N_7588,N_6798);
nor U8819 (N_8819,N_7469,N_6124);
xnor U8820 (N_8820,N_7019,N_6602);
nor U8821 (N_8821,N_6231,N_7861);
xnor U8822 (N_8822,N_7955,N_6414);
nand U8823 (N_8823,N_6614,N_6838);
nor U8824 (N_8824,N_6242,N_7429);
xnor U8825 (N_8825,N_7911,N_6473);
nand U8826 (N_8826,N_7880,N_7991);
and U8827 (N_8827,N_7808,N_6045);
xor U8828 (N_8828,N_6835,N_7994);
nand U8829 (N_8829,N_7640,N_7565);
xnor U8830 (N_8830,N_7324,N_7256);
nor U8831 (N_8831,N_7694,N_7259);
nor U8832 (N_8832,N_7476,N_7643);
nor U8833 (N_8833,N_6609,N_7846);
nor U8834 (N_8834,N_6594,N_7250);
and U8835 (N_8835,N_7343,N_7943);
xor U8836 (N_8836,N_7984,N_6483);
xnor U8837 (N_8837,N_7315,N_7240);
and U8838 (N_8838,N_6936,N_6601);
and U8839 (N_8839,N_6792,N_6894);
nand U8840 (N_8840,N_7621,N_6809);
nand U8841 (N_8841,N_7656,N_7844);
nor U8842 (N_8842,N_7990,N_6716);
and U8843 (N_8843,N_6028,N_6727);
xor U8844 (N_8844,N_7907,N_7596);
nand U8845 (N_8845,N_6060,N_7646);
nand U8846 (N_8846,N_6982,N_6236);
or U8847 (N_8847,N_6137,N_6357);
xor U8848 (N_8848,N_7489,N_6167);
nor U8849 (N_8849,N_7378,N_6243);
nor U8850 (N_8850,N_6656,N_7935);
and U8851 (N_8851,N_6019,N_7251);
or U8852 (N_8852,N_7392,N_7616);
nand U8853 (N_8853,N_7142,N_7929);
or U8854 (N_8854,N_6102,N_6713);
xnor U8855 (N_8855,N_7705,N_7038);
or U8856 (N_8856,N_7532,N_7989);
and U8857 (N_8857,N_7481,N_6286);
or U8858 (N_8858,N_6561,N_6301);
or U8859 (N_8859,N_6453,N_7641);
xor U8860 (N_8860,N_7722,N_6930);
nand U8861 (N_8861,N_7156,N_6891);
nand U8862 (N_8862,N_6797,N_6946);
or U8863 (N_8863,N_7005,N_7401);
xnor U8864 (N_8864,N_6808,N_6574);
or U8865 (N_8865,N_6466,N_7244);
or U8866 (N_8866,N_6450,N_6027);
nand U8867 (N_8867,N_6358,N_7355);
xor U8868 (N_8868,N_7314,N_7058);
nor U8869 (N_8869,N_7309,N_6182);
nor U8870 (N_8870,N_7853,N_6646);
nor U8871 (N_8871,N_7901,N_6340);
nor U8872 (N_8872,N_6901,N_7252);
xor U8873 (N_8873,N_6651,N_6459);
nor U8874 (N_8874,N_7423,N_7732);
and U8875 (N_8875,N_7362,N_6389);
and U8876 (N_8876,N_7693,N_6999);
and U8877 (N_8877,N_7649,N_6210);
xor U8878 (N_8878,N_6128,N_7017);
nand U8879 (N_8879,N_7542,N_7045);
or U8880 (N_8880,N_7397,N_6533);
and U8881 (N_8881,N_6052,N_7798);
nor U8882 (N_8882,N_7004,N_6116);
nor U8883 (N_8883,N_7456,N_6911);
and U8884 (N_8884,N_6732,N_7069);
nor U8885 (N_8885,N_7774,N_7951);
xor U8886 (N_8886,N_7731,N_7470);
or U8887 (N_8887,N_7224,N_6049);
nand U8888 (N_8888,N_6376,N_6582);
or U8889 (N_8889,N_7262,N_6003);
nor U8890 (N_8890,N_7177,N_7848);
nor U8891 (N_8891,N_6203,N_7169);
xnor U8892 (N_8892,N_6418,N_7186);
nor U8893 (N_8893,N_6772,N_6847);
and U8894 (N_8894,N_7376,N_6387);
nor U8895 (N_8895,N_6505,N_7962);
nor U8896 (N_8896,N_7388,N_6155);
or U8897 (N_8897,N_6563,N_6874);
and U8898 (N_8898,N_7781,N_7232);
nand U8899 (N_8899,N_7130,N_7119);
or U8900 (N_8900,N_7472,N_6529);
xnor U8901 (N_8901,N_7363,N_6095);
and U8902 (N_8902,N_6766,N_6737);
and U8903 (N_8903,N_7433,N_6191);
and U8904 (N_8904,N_6956,N_6147);
and U8905 (N_8905,N_6070,N_6139);
and U8906 (N_8906,N_7842,N_6546);
or U8907 (N_8907,N_7790,N_7604);
and U8908 (N_8908,N_6249,N_6192);
nor U8909 (N_8909,N_6677,N_7562);
and U8910 (N_8910,N_6986,N_6667);
or U8911 (N_8911,N_6597,N_6645);
nand U8912 (N_8912,N_7714,N_6892);
xor U8913 (N_8913,N_6786,N_6461);
nand U8914 (N_8914,N_6087,N_6841);
nor U8915 (N_8915,N_7594,N_7121);
or U8916 (N_8916,N_7242,N_6491);
xor U8917 (N_8917,N_7061,N_6741);
nor U8918 (N_8918,N_6089,N_6287);
nor U8919 (N_8919,N_7112,N_6262);
or U8920 (N_8920,N_7339,N_6773);
or U8921 (N_8921,N_7155,N_7046);
or U8922 (N_8922,N_6164,N_7780);
nor U8923 (N_8923,N_6447,N_7099);
nand U8924 (N_8924,N_7811,N_7936);
nor U8925 (N_8925,N_6870,N_6559);
or U8926 (N_8926,N_7083,N_7559);
xnor U8927 (N_8927,N_7471,N_6487);
or U8928 (N_8928,N_7796,N_7999);
and U8929 (N_8929,N_7081,N_7553);
and U8930 (N_8930,N_7097,N_7899);
xor U8931 (N_8931,N_6612,N_7140);
nand U8932 (N_8932,N_7536,N_7434);
or U8933 (N_8933,N_6925,N_7998);
or U8934 (N_8934,N_6404,N_7863);
or U8935 (N_8935,N_7442,N_7210);
nor U8936 (N_8936,N_6100,N_7205);
nand U8937 (N_8937,N_6717,N_6470);
xor U8938 (N_8938,N_7838,N_7533);
or U8939 (N_8939,N_6682,N_7866);
or U8940 (N_8940,N_7822,N_6117);
nor U8941 (N_8941,N_7529,N_7495);
and U8942 (N_8942,N_6131,N_6031);
nor U8943 (N_8943,N_7106,N_7333);
or U8944 (N_8944,N_6047,N_6140);
or U8945 (N_8945,N_7023,N_6403);
nor U8946 (N_8946,N_7238,N_6416);
nor U8947 (N_8947,N_6245,N_7915);
or U8948 (N_8948,N_6037,N_6316);
and U8949 (N_8949,N_6176,N_7833);
xor U8950 (N_8950,N_6544,N_6926);
nand U8951 (N_8951,N_6465,N_6330);
and U8952 (N_8952,N_7645,N_7890);
xor U8953 (N_8953,N_6787,N_7642);
or U8954 (N_8954,N_6922,N_6760);
or U8955 (N_8955,N_7448,N_7952);
xor U8956 (N_8956,N_6061,N_7405);
and U8957 (N_8957,N_7337,N_7591);
or U8958 (N_8958,N_7071,N_6401);
and U8959 (N_8959,N_6800,N_6556);
or U8960 (N_8960,N_7278,N_6886);
and U8961 (N_8961,N_7227,N_6170);
nor U8962 (N_8962,N_7006,N_7449);
or U8963 (N_8963,N_7608,N_6064);
nand U8964 (N_8964,N_7698,N_7090);
nand U8965 (N_8965,N_6735,N_6763);
xnor U8966 (N_8966,N_7683,N_6214);
nand U8967 (N_8967,N_7020,N_6081);
and U8968 (N_8968,N_7716,N_6587);
nand U8969 (N_8969,N_7937,N_6707);
or U8970 (N_8970,N_7195,N_6873);
and U8971 (N_8971,N_7356,N_6166);
xor U8972 (N_8972,N_7289,N_6076);
nand U8973 (N_8973,N_6955,N_7074);
or U8974 (N_8974,N_7843,N_7453);
nor U8975 (N_8975,N_6258,N_6720);
or U8976 (N_8976,N_6939,N_6501);
or U8977 (N_8977,N_7801,N_7635);
nand U8978 (N_8978,N_7108,N_7485);
nor U8979 (N_8979,N_7479,N_6817);
nor U8980 (N_8980,N_7567,N_7003);
and U8981 (N_8981,N_7840,N_7718);
nand U8982 (N_8982,N_6423,N_7400);
xor U8983 (N_8983,N_6959,N_7818);
or U8984 (N_8984,N_6777,N_7386);
or U8985 (N_8985,N_7579,N_7682);
xnor U8986 (N_8986,N_6549,N_6158);
nor U8987 (N_8987,N_6734,N_6256);
xnor U8988 (N_8988,N_6350,N_6774);
xnor U8989 (N_8989,N_7677,N_7785);
nand U8990 (N_8990,N_7571,N_6426);
or U8991 (N_8991,N_6232,N_7779);
or U8992 (N_8992,N_7828,N_7302);
or U8993 (N_8993,N_7982,N_6568);
nor U8994 (N_8994,N_6341,N_6406);
and U8995 (N_8995,N_6778,N_6576);
or U8996 (N_8996,N_6526,N_7839);
xnor U8997 (N_8997,N_7770,N_6435);
nor U8998 (N_8998,N_6201,N_7862);
and U8999 (N_8999,N_7742,N_6641);
or U9000 (N_9000,N_7899,N_7005);
nor U9001 (N_9001,N_7592,N_7195);
nand U9002 (N_9002,N_6985,N_6251);
nand U9003 (N_9003,N_6271,N_7968);
nor U9004 (N_9004,N_7077,N_7789);
nand U9005 (N_9005,N_6299,N_6856);
nand U9006 (N_9006,N_6320,N_6013);
and U9007 (N_9007,N_7452,N_7582);
nand U9008 (N_9008,N_6879,N_6236);
xor U9009 (N_9009,N_6995,N_7152);
xnor U9010 (N_9010,N_6514,N_7654);
xor U9011 (N_9011,N_6848,N_7127);
or U9012 (N_9012,N_7386,N_6699);
xnor U9013 (N_9013,N_6457,N_7980);
and U9014 (N_9014,N_6569,N_7363);
xnor U9015 (N_9015,N_7836,N_7209);
xnor U9016 (N_9016,N_7578,N_6014);
nand U9017 (N_9017,N_6193,N_6282);
and U9018 (N_9018,N_7350,N_6826);
and U9019 (N_9019,N_7176,N_6149);
nor U9020 (N_9020,N_6416,N_6962);
or U9021 (N_9021,N_6556,N_7115);
and U9022 (N_9022,N_6649,N_6084);
and U9023 (N_9023,N_6963,N_6090);
nor U9024 (N_9024,N_6473,N_6643);
nand U9025 (N_9025,N_7738,N_6666);
xor U9026 (N_9026,N_6303,N_6174);
xor U9027 (N_9027,N_7894,N_6964);
nand U9028 (N_9028,N_6897,N_6889);
nor U9029 (N_9029,N_6378,N_6998);
or U9030 (N_9030,N_6992,N_7938);
xor U9031 (N_9031,N_7794,N_7171);
xor U9032 (N_9032,N_7363,N_7185);
xor U9033 (N_9033,N_7444,N_6577);
or U9034 (N_9034,N_6210,N_7656);
or U9035 (N_9035,N_6192,N_7818);
nand U9036 (N_9036,N_6784,N_6464);
xnor U9037 (N_9037,N_6325,N_7508);
nand U9038 (N_9038,N_7162,N_7238);
xnor U9039 (N_9039,N_6534,N_7063);
xnor U9040 (N_9040,N_6411,N_6924);
nand U9041 (N_9041,N_6525,N_6575);
and U9042 (N_9042,N_6214,N_6309);
nor U9043 (N_9043,N_6077,N_6856);
or U9044 (N_9044,N_6965,N_6790);
nor U9045 (N_9045,N_7531,N_6400);
xor U9046 (N_9046,N_7828,N_6929);
xor U9047 (N_9047,N_6956,N_6575);
xnor U9048 (N_9048,N_7803,N_7813);
or U9049 (N_9049,N_6390,N_6331);
nand U9050 (N_9050,N_6269,N_6548);
or U9051 (N_9051,N_6908,N_7232);
nand U9052 (N_9052,N_6109,N_7030);
or U9053 (N_9053,N_6648,N_7039);
nand U9054 (N_9054,N_6309,N_6907);
or U9055 (N_9055,N_7552,N_7761);
xnor U9056 (N_9056,N_7284,N_6710);
xor U9057 (N_9057,N_6379,N_6772);
xnor U9058 (N_9058,N_7653,N_7443);
nand U9059 (N_9059,N_7603,N_6554);
xnor U9060 (N_9060,N_7652,N_7633);
nor U9061 (N_9061,N_6170,N_7382);
and U9062 (N_9062,N_6424,N_6636);
xor U9063 (N_9063,N_7941,N_6129);
or U9064 (N_9064,N_6046,N_7259);
xor U9065 (N_9065,N_6357,N_6021);
and U9066 (N_9066,N_6549,N_6127);
xor U9067 (N_9067,N_6653,N_7753);
xnor U9068 (N_9068,N_6848,N_7650);
nand U9069 (N_9069,N_7742,N_6859);
nor U9070 (N_9070,N_6383,N_6361);
xnor U9071 (N_9071,N_6421,N_6332);
xor U9072 (N_9072,N_7506,N_6920);
nand U9073 (N_9073,N_7453,N_7842);
and U9074 (N_9074,N_6293,N_7198);
xor U9075 (N_9075,N_6034,N_6721);
xor U9076 (N_9076,N_7211,N_7794);
nand U9077 (N_9077,N_6217,N_7453);
nor U9078 (N_9078,N_7274,N_7771);
nor U9079 (N_9079,N_6395,N_7015);
nor U9080 (N_9080,N_6922,N_6951);
nor U9081 (N_9081,N_7273,N_6300);
and U9082 (N_9082,N_7400,N_6758);
nand U9083 (N_9083,N_6108,N_6675);
and U9084 (N_9084,N_6340,N_7590);
nor U9085 (N_9085,N_7990,N_7766);
or U9086 (N_9086,N_6854,N_6709);
or U9087 (N_9087,N_6862,N_7852);
or U9088 (N_9088,N_7735,N_6093);
nor U9089 (N_9089,N_7266,N_6289);
nor U9090 (N_9090,N_7916,N_6756);
and U9091 (N_9091,N_6057,N_7060);
nand U9092 (N_9092,N_6510,N_7194);
or U9093 (N_9093,N_7282,N_7664);
and U9094 (N_9094,N_7632,N_7230);
nor U9095 (N_9095,N_6314,N_6927);
nor U9096 (N_9096,N_6756,N_6482);
nand U9097 (N_9097,N_7797,N_7194);
and U9098 (N_9098,N_7228,N_7149);
and U9099 (N_9099,N_6771,N_7564);
and U9100 (N_9100,N_6438,N_7935);
or U9101 (N_9101,N_6741,N_7158);
and U9102 (N_9102,N_6802,N_6165);
and U9103 (N_9103,N_6399,N_6424);
and U9104 (N_9104,N_6271,N_6434);
xor U9105 (N_9105,N_7431,N_7935);
nor U9106 (N_9106,N_6481,N_7786);
nor U9107 (N_9107,N_7806,N_6563);
xor U9108 (N_9108,N_7861,N_7526);
nand U9109 (N_9109,N_7539,N_7882);
and U9110 (N_9110,N_6307,N_6985);
nor U9111 (N_9111,N_6395,N_7193);
and U9112 (N_9112,N_6890,N_7284);
nor U9113 (N_9113,N_7083,N_7943);
nand U9114 (N_9114,N_6135,N_7315);
or U9115 (N_9115,N_6339,N_7339);
and U9116 (N_9116,N_7223,N_6531);
nor U9117 (N_9117,N_6764,N_7978);
nor U9118 (N_9118,N_7872,N_7024);
nand U9119 (N_9119,N_6636,N_6443);
and U9120 (N_9120,N_6304,N_7544);
and U9121 (N_9121,N_7107,N_6010);
or U9122 (N_9122,N_7640,N_6260);
nand U9123 (N_9123,N_7910,N_6805);
xnor U9124 (N_9124,N_7752,N_6144);
nand U9125 (N_9125,N_6075,N_6222);
or U9126 (N_9126,N_7422,N_7670);
xor U9127 (N_9127,N_6562,N_7990);
and U9128 (N_9128,N_7350,N_7839);
and U9129 (N_9129,N_6859,N_7348);
or U9130 (N_9130,N_6177,N_6082);
nand U9131 (N_9131,N_7400,N_7504);
nor U9132 (N_9132,N_6410,N_7126);
and U9133 (N_9133,N_7964,N_7711);
nor U9134 (N_9134,N_7045,N_7065);
xnor U9135 (N_9135,N_6005,N_6309);
or U9136 (N_9136,N_7634,N_7440);
nor U9137 (N_9137,N_7602,N_6137);
or U9138 (N_9138,N_7510,N_6496);
nor U9139 (N_9139,N_7224,N_7798);
nand U9140 (N_9140,N_7878,N_6601);
xor U9141 (N_9141,N_6468,N_6605);
or U9142 (N_9142,N_7851,N_7639);
nand U9143 (N_9143,N_7156,N_6047);
xor U9144 (N_9144,N_7596,N_7148);
xnor U9145 (N_9145,N_7187,N_7836);
and U9146 (N_9146,N_7836,N_7834);
xor U9147 (N_9147,N_6244,N_6611);
or U9148 (N_9148,N_6810,N_7874);
or U9149 (N_9149,N_6928,N_6201);
and U9150 (N_9150,N_6510,N_6937);
or U9151 (N_9151,N_7887,N_6555);
xnor U9152 (N_9152,N_7144,N_6484);
xnor U9153 (N_9153,N_6803,N_6684);
and U9154 (N_9154,N_7235,N_6260);
or U9155 (N_9155,N_7020,N_7369);
xnor U9156 (N_9156,N_6734,N_7958);
nand U9157 (N_9157,N_6733,N_7881);
and U9158 (N_9158,N_7294,N_6966);
or U9159 (N_9159,N_6062,N_7265);
nand U9160 (N_9160,N_7940,N_6778);
nand U9161 (N_9161,N_7182,N_7988);
xor U9162 (N_9162,N_6952,N_6766);
xnor U9163 (N_9163,N_7471,N_7564);
and U9164 (N_9164,N_7647,N_7918);
nor U9165 (N_9165,N_7749,N_6166);
nand U9166 (N_9166,N_6529,N_6494);
and U9167 (N_9167,N_7317,N_6664);
nor U9168 (N_9168,N_6320,N_6509);
xnor U9169 (N_9169,N_7612,N_7012);
or U9170 (N_9170,N_7360,N_7884);
or U9171 (N_9171,N_7261,N_7756);
or U9172 (N_9172,N_6944,N_7905);
xnor U9173 (N_9173,N_7892,N_6665);
nand U9174 (N_9174,N_7079,N_7980);
or U9175 (N_9175,N_7925,N_6137);
nand U9176 (N_9176,N_6349,N_6677);
and U9177 (N_9177,N_6844,N_7949);
xnor U9178 (N_9178,N_7083,N_6742);
xnor U9179 (N_9179,N_7722,N_7640);
or U9180 (N_9180,N_6174,N_6150);
or U9181 (N_9181,N_7116,N_6064);
nand U9182 (N_9182,N_7701,N_7981);
nand U9183 (N_9183,N_6615,N_6704);
xor U9184 (N_9184,N_7131,N_6741);
xor U9185 (N_9185,N_6375,N_6320);
xor U9186 (N_9186,N_6426,N_7540);
xnor U9187 (N_9187,N_7710,N_6911);
xor U9188 (N_9188,N_7783,N_7747);
xor U9189 (N_9189,N_6019,N_7054);
xnor U9190 (N_9190,N_6936,N_6249);
and U9191 (N_9191,N_7809,N_6794);
and U9192 (N_9192,N_6174,N_6867);
xor U9193 (N_9193,N_7104,N_7466);
and U9194 (N_9194,N_6061,N_6891);
nand U9195 (N_9195,N_6308,N_6849);
nor U9196 (N_9196,N_7271,N_7902);
or U9197 (N_9197,N_6919,N_6456);
xor U9198 (N_9198,N_6284,N_7256);
nor U9199 (N_9199,N_6292,N_6758);
xor U9200 (N_9200,N_6238,N_7990);
and U9201 (N_9201,N_7608,N_7650);
or U9202 (N_9202,N_7738,N_6568);
xor U9203 (N_9203,N_6745,N_6353);
nand U9204 (N_9204,N_6707,N_6667);
nor U9205 (N_9205,N_6069,N_7431);
xnor U9206 (N_9206,N_6489,N_6914);
and U9207 (N_9207,N_7553,N_7697);
nand U9208 (N_9208,N_7750,N_6215);
xor U9209 (N_9209,N_7091,N_6109);
and U9210 (N_9210,N_7567,N_7082);
and U9211 (N_9211,N_6581,N_7811);
and U9212 (N_9212,N_6560,N_7210);
nor U9213 (N_9213,N_7624,N_6293);
nand U9214 (N_9214,N_7233,N_6587);
and U9215 (N_9215,N_7828,N_6152);
nor U9216 (N_9216,N_6377,N_6493);
nor U9217 (N_9217,N_7548,N_7919);
nand U9218 (N_9218,N_6034,N_6330);
xnor U9219 (N_9219,N_6816,N_6607);
and U9220 (N_9220,N_7360,N_7350);
and U9221 (N_9221,N_6678,N_7251);
nor U9222 (N_9222,N_6541,N_7641);
xnor U9223 (N_9223,N_7558,N_6535);
and U9224 (N_9224,N_6883,N_7599);
xor U9225 (N_9225,N_6184,N_6179);
nor U9226 (N_9226,N_6241,N_7003);
xor U9227 (N_9227,N_6021,N_6586);
and U9228 (N_9228,N_6147,N_7261);
or U9229 (N_9229,N_6329,N_6755);
nor U9230 (N_9230,N_6956,N_6817);
nor U9231 (N_9231,N_6842,N_7209);
and U9232 (N_9232,N_7114,N_6566);
and U9233 (N_9233,N_6679,N_7474);
and U9234 (N_9234,N_7308,N_6366);
xnor U9235 (N_9235,N_6560,N_6086);
nand U9236 (N_9236,N_6241,N_6322);
nand U9237 (N_9237,N_6458,N_6015);
nor U9238 (N_9238,N_7741,N_7181);
xnor U9239 (N_9239,N_7689,N_7096);
or U9240 (N_9240,N_7983,N_6648);
nand U9241 (N_9241,N_7161,N_6936);
or U9242 (N_9242,N_7667,N_7937);
and U9243 (N_9243,N_6473,N_7582);
or U9244 (N_9244,N_7483,N_6595);
nand U9245 (N_9245,N_7399,N_7500);
nor U9246 (N_9246,N_7984,N_7035);
nor U9247 (N_9247,N_7841,N_7189);
xor U9248 (N_9248,N_6595,N_6408);
xor U9249 (N_9249,N_6946,N_7518);
and U9250 (N_9250,N_7377,N_7197);
and U9251 (N_9251,N_7919,N_6691);
nand U9252 (N_9252,N_7046,N_7028);
nor U9253 (N_9253,N_6470,N_6574);
nor U9254 (N_9254,N_7295,N_7168);
or U9255 (N_9255,N_7430,N_7621);
nand U9256 (N_9256,N_6256,N_7815);
nand U9257 (N_9257,N_7341,N_6518);
or U9258 (N_9258,N_7702,N_7464);
nor U9259 (N_9259,N_6003,N_6417);
xor U9260 (N_9260,N_7366,N_6208);
xor U9261 (N_9261,N_7554,N_6015);
and U9262 (N_9262,N_6975,N_7399);
nand U9263 (N_9263,N_7091,N_6434);
nor U9264 (N_9264,N_6823,N_6897);
nand U9265 (N_9265,N_7789,N_6083);
xnor U9266 (N_9266,N_6742,N_7956);
xor U9267 (N_9267,N_6638,N_6412);
or U9268 (N_9268,N_6863,N_7241);
xor U9269 (N_9269,N_6935,N_6852);
xnor U9270 (N_9270,N_7639,N_7292);
nand U9271 (N_9271,N_6059,N_7257);
or U9272 (N_9272,N_6077,N_6943);
nor U9273 (N_9273,N_7203,N_7924);
and U9274 (N_9274,N_6994,N_7980);
and U9275 (N_9275,N_7541,N_6381);
or U9276 (N_9276,N_6909,N_7337);
and U9277 (N_9277,N_7007,N_7823);
nand U9278 (N_9278,N_7731,N_6775);
or U9279 (N_9279,N_7230,N_6638);
and U9280 (N_9280,N_6608,N_6193);
and U9281 (N_9281,N_7522,N_6216);
or U9282 (N_9282,N_6572,N_6780);
nor U9283 (N_9283,N_6402,N_7994);
nand U9284 (N_9284,N_7791,N_7849);
xor U9285 (N_9285,N_6389,N_6785);
or U9286 (N_9286,N_7317,N_7131);
or U9287 (N_9287,N_7992,N_6939);
nand U9288 (N_9288,N_6799,N_7159);
nand U9289 (N_9289,N_6715,N_7394);
xnor U9290 (N_9290,N_7352,N_7149);
nor U9291 (N_9291,N_7543,N_7137);
xnor U9292 (N_9292,N_6777,N_7353);
nor U9293 (N_9293,N_7937,N_7154);
xor U9294 (N_9294,N_6818,N_6842);
nor U9295 (N_9295,N_7204,N_6487);
nand U9296 (N_9296,N_6888,N_7632);
or U9297 (N_9297,N_6938,N_6676);
or U9298 (N_9298,N_6356,N_6739);
xnor U9299 (N_9299,N_6348,N_7475);
or U9300 (N_9300,N_7288,N_7727);
and U9301 (N_9301,N_6156,N_6757);
and U9302 (N_9302,N_7464,N_7075);
nand U9303 (N_9303,N_6243,N_6059);
or U9304 (N_9304,N_6126,N_6540);
or U9305 (N_9305,N_7476,N_7929);
and U9306 (N_9306,N_6118,N_6882);
nor U9307 (N_9307,N_6500,N_6181);
or U9308 (N_9308,N_6496,N_7791);
nand U9309 (N_9309,N_6787,N_7558);
and U9310 (N_9310,N_6685,N_7328);
xnor U9311 (N_9311,N_7072,N_6998);
nand U9312 (N_9312,N_6317,N_7623);
and U9313 (N_9313,N_6258,N_7949);
nor U9314 (N_9314,N_7307,N_7777);
xor U9315 (N_9315,N_7657,N_6727);
and U9316 (N_9316,N_6608,N_6227);
or U9317 (N_9317,N_6499,N_6240);
nand U9318 (N_9318,N_6095,N_7255);
and U9319 (N_9319,N_6651,N_7047);
or U9320 (N_9320,N_7719,N_7119);
and U9321 (N_9321,N_7909,N_7328);
or U9322 (N_9322,N_7557,N_6307);
nor U9323 (N_9323,N_7945,N_6037);
nand U9324 (N_9324,N_6893,N_7418);
nand U9325 (N_9325,N_6871,N_6999);
and U9326 (N_9326,N_6811,N_6826);
xnor U9327 (N_9327,N_7591,N_6636);
and U9328 (N_9328,N_7996,N_7875);
or U9329 (N_9329,N_6348,N_7480);
nand U9330 (N_9330,N_6061,N_6486);
nand U9331 (N_9331,N_6145,N_7160);
and U9332 (N_9332,N_6178,N_7978);
xnor U9333 (N_9333,N_7983,N_7929);
or U9334 (N_9334,N_7646,N_7219);
or U9335 (N_9335,N_6580,N_7153);
nand U9336 (N_9336,N_6169,N_6895);
and U9337 (N_9337,N_7092,N_7615);
nand U9338 (N_9338,N_6552,N_7472);
or U9339 (N_9339,N_7398,N_6048);
or U9340 (N_9340,N_7124,N_7301);
nor U9341 (N_9341,N_6498,N_7526);
or U9342 (N_9342,N_6511,N_6253);
nor U9343 (N_9343,N_7500,N_7341);
and U9344 (N_9344,N_7877,N_6453);
nor U9345 (N_9345,N_7363,N_7979);
nor U9346 (N_9346,N_6079,N_7099);
nor U9347 (N_9347,N_7187,N_6805);
nand U9348 (N_9348,N_6180,N_7815);
or U9349 (N_9349,N_7588,N_7711);
nand U9350 (N_9350,N_6341,N_7489);
nor U9351 (N_9351,N_7077,N_6814);
nor U9352 (N_9352,N_7634,N_7276);
nand U9353 (N_9353,N_7203,N_6274);
or U9354 (N_9354,N_6480,N_7692);
xnor U9355 (N_9355,N_7937,N_6029);
nor U9356 (N_9356,N_7610,N_7950);
and U9357 (N_9357,N_6885,N_6758);
nand U9358 (N_9358,N_6335,N_7477);
xnor U9359 (N_9359,N_6563,N_7964);
nor U9360 (N_9360,N_6237,N_6348);
and U9361 (N_9361,N_6825,N_7892);
nand U9362 (N_9362,N_7421,N_7575);
and U9363 (N_9363,N_6722,N_6525);
and U9364 (N_9364,N_7180,N_7741);
nand U9365 (N_9365,N_6698,N_7183);
nand U9366 (N_9366,N_7049,N_6690);
and U9367 (N_9367,N_7719,N_6033);
and U9368 (N_9368,N_6174,N_7083);
nor U9369 (N_9369,N_7458,N_7460);
or U9370 (N_9370,N_6381,N_7031);
nand U9371 (N_9371,N_6667,N_6937);
nor U9372 (N_9372,N_7810,N_7271);
or U9373 (N_9373,N_7960,N_7593);
nor U9374 (N_9374,N_7496,N_6875);
and U9375 (N_9375,N_6401,N_6405);
xnor U9376 (N_9376,N_7362,N_7200);
nand U9377 (N_9377,N_7902,N_7363);
and U9378 (N_9378,N_7109,N_6464);
nand U9379 (N_9379,N_7126,N_6534);
and U9380 (N_9380,N_7792,N_6825);
or U9381 (N_9381,N_7458,N_6398);
xor U9382 (N_9382,N_7182,N_6682);
nor U9383 (N_9383,N_7949,N_7007);
nor U9384 (N_9384,N_7279,N_6811);
or U9385 (N_9385,N_6277,N_7541);
nand U9386 (N_9386,N_6157,N_6796);
or U9387 (N_9387,N_7066,N_6185);
and U9388 (N_9388,N_6978,N_6737);
nand U9389 (N_9389,N_6942,N_6720);
nand U9390 (N_9390,N_7186,N_7593);
and U9391 (N_9391,N_6014,N_6341);
or U9392 (N_9392,N_6914,N_6182);
or U9393 (N_9393,N_7583,N_7486);
nand U9394 (N_9394,N_6168,N_7648);
and U9395 (N_9395,N_6086,N_6175);
nor U9396 (N_9396,N_7278,N_6703);
nor U9397 (N_9397,N_7980,N_6158);
or U9398 (N_9398,N_6192,N_7651);
and U9399 (N_9399,N_7036,N_7701);
and U9400 (N_9400,N_7567,N_6308);
and U9401 (N_9401,N_6601,N_7564);
nand U9402 (N_9402,N_6759,N_6813);
nand U9403 (N_9403,N_6522,N_6334);
xnor U9404 (N_9404,N_7579,N_6498);
nor U9405 (N_9405,N_6799,N_7617);
nor U9406 (N_9406,N_7249,N_6226);
and U9407 (N_9407,N_7332,N_7336);
xnor U9408 (N_9408,N_7471,N_6673);
and U9409 (N_9409,N_6043,N_6845);
or U9410 (N_9410,N_6615,N_6588);
xnor U9411 (N_9411,N_6959,N_6606);
and U9412 (N_9412,N_7969,N_7006);
or U9413 (N_9413,N_6785,N_7245);
and U9414 (N_9414,N_6590,N_6433);
nor U9415 (N_9415,N_7987,N_7201);
or U9416 (N_9416,N_7457,N_6702);
nand U9417 (N_9417,N_7873,N_7354);
nor U9418 (N_9418,N_7690,N_7495);
nand U9419 (N_9419,N_6284,N_7550);
or U9420 (N_9420,N_6077,N_7472);
and U9421 (N_9421,N_7090,N_7827);
xor U9422 (N_9422,N_6234,N_7030);
xnor U9423 (N_9423,N_6842,N_7426);
nor U9424 (N_9424,N_6531,N_6839);
xnor U9425 (N_9425,N_6644,N_6887);
xnor U9426 (N_9426,N_6653,N_7396);
or U9427 (N_9427,N_7967,N_7297);
or U9428 (N_9428,N_6075,N_7670);
nand U9429 (N_9429,N_7076,N_6355);
or U9430 (N_9430,N_7742,N_7381);
nand U9431 (N_9431,N_6898,N_6695);
xnor U9432 (N_9432,N_6298,N_6896);
and U9433 (N_9433,N_6373,N_6885);
nor U9434 (N_9434,N_6779,N_6060);
nor U9435 (N_9435,N_6793,N_6103);
and U9436 (N_9436,N_6021,N_6131);
and U9437 (N_9437,N_7456,N_7503);
nand U9438 (N_9438,N_7418,N_7968);
xnor U9439 (N_9439,N_7802,N_7560);
nand U9440 (N_9440,N_6867,N_6795);
xor U9441 (N_9441,N_6508,N_7611);
xnor U9442 (N_9442,N_7328,N_7848);
and U9443 (N_9443,N_7251,N_7872);
and U9444 (N_9444,N_6878,N_7658);
and U9445 (N_9445,N_6746,N_6000);
and U9446 (N_9446,N_6613,N_7927);
and U9447 (N_9447,N_6608,N_6818);
and U9448 (N_9448,N_7728,N_6929);
xor U9449 (N_9449,N_7284,N_6661);
xor U9450 (N_9450,N_6691,N_7843);
or U9451 (N_9451,N_6345,N_7303);
nand U9452 (N_9452,N_7362,N_7879);
or U9453 (N_9453,N_7740,N_6446);
or U9454 (N_9454,N_6341,N_6567);
or U9455 (N_9455,N_6057,N_6955);
and U9456 (N_9456,N_7161,N_7659);
nor U9457 (N_9457,N_6001,N_7616);
and U9458 (N_9458,N_6870,N_6847);
nor U9459 (N_9459,N_6870,N_6184);
nor U9460 (N_9460,N_6110,N_6537);
nand U9461 (N_9461,N_6397,N_6219);
nor U9462 (N_9462,N_7977,N_7829);
nand U9463 (N_9463,N_6918,N_7112);
nand U9464 (N_9464,N_6309,N_7597);
nor U9465 (N_9465,N_7520,N_6230);
or U9466 (N_9466,N_7989,N_7512);
xnor U9467 (N_9467,N_7539,N_6569);
nor U9468 (N_9468,N_6456,N_6995);
nand U9469 (N_9469,N_6485,N_6788);
nor U9470 (N_9470,N_7899,N_6124);
nor U9471 (N_9471,N_6054,N_6158);
xnor U9472 (N_9472,N_6786,N_7066);
xnor U9473 (N_9473,N_7218,N_6213);
nand U9474 (N_9474,N_7886,N_6706);
and U9475 (N_9475,N_7768,N_6041);
or U9476 (N_9476,N_7474,N_6389);
nor U9477 (N_9477,N_7070,N_7037);
nor U9478 (N_9478,N_6855,N_6824);
nor U9479 (N_9479,N_6211,N_6688);
and U9480 (N_9480,N_6816,N_6933);
nor U9481 (N_9481,N_6485,N_6635);
or U9482 (N_9482,N_7053,N_7216);
nand U9483 (N_9483,N_6900,N_6323);
nand U9484 (N_9484,N_6276,N_7952);
and U9485 (N_9485,N_7383,N_7000);
or U9486 (N_9486,N_7129,N_7429);
nand U9487 (N_9487,N_6334,N_6949);
and U9488 (N_9488,N_7253,N_6257);
and U9489 (N_9489,N_7303,N_7915);
nand U9490 (N_9490,N_6631,N_7788);
nand U9491 (N_9491,N_7382,N_7218);
and U9492 (N_9492,N_6392,N_7498);
xnor U9493 (N_9493,N_6251,N_7227);
nand U9494 (N_9494,N_6368,N_7629);
xor U9495 (N_9495,N_7230,N_7466);
xor U9496 (N_9496,N_6736,N_6109);
nor U9497 (N_9497,N_6004,N_7254);
nor U9498 (N_9498,N_6866,N_6008);
nor U9499 (N_9499,N_7768,N_7782);
and U9500 (N_9500,N_7670,N_6128);
or U9501 (N_9501,N_7549,N_7248);
nand U9502 (N_9502,N_7391,N_6166);
or U9503 (N_9503,N_6746,N_7286);
nor U9504 (N_9504,N_7424,N_6058);
or U9505 (N_9505,N_7097,N_6435);
nand U9506 (N_9506,N_6315,N_7801);
nand U9507 (N_9507,N_7048,N_6796);
nand U9508 (N_9508,N_7959,N_6674);
xor U9509 (N_9509,N_7752,N_6529);
xnor U9510 (N_9510,N_6720,N_6395);
and U9511 (N_9511,N_7305,N_7025);
nor U9512 (N_9512,N_6233,N_6026);
and U9513 (N_9513,N_7087,N_7301);
xor U9514 (N_9514,N_7192,N_6114);
and U9515 (N_9515,N_6116,N_6339);
nand U9516 (N_9516,N_6664,N_7316);
and U9517 (N_9517,N_7163,N_6489);
nor U9518 (N_9518,N_6479,N_6593);
xnor U9519 (N_9519,N_6410,N_7594);
nand U9520 (N_9520,N_7460,N_6805);
nor U9521 (N_9521,N_6656,N_6856);
xor U9522 (N_9522,N_7609,N_7680);
and U9523 (N_9523,N_6852,N_6707);
nand U9524 (N_9524,N_6714,N_6210);
or U9525 (N_9525,N_6898,N_6288);
or U9526 (N_9526,N_7220,N_6157);
xor U9527 (N_9527,N_6465,N_7899);
nand U9528 (N_9528,N_7256,N_7287);
xor U9529 (N_9529,N_6706,N_6119);
nor U9530 (N_9530,N_7521,N_6651);
and U9531 (N_9531,N_7718,N_7110);
nor U9532 (N_9532,N_7126,N_7781);
and U9533 (N_9533,N_7657,N_7914);
and U9534 (N_9534,N_6355,N_7835);
nor U9535 (N_9535,N_6594,N_7555);
xnor U9536 (N_9536,N_6924,N_6705);
nor U9537 (N_9537,N_7729,N_6040);
xor U9538 (N_9538,N_6795,N_7250);
xnor U9539 (N_9539,N_7768,N_6233);
nand U9540 (N_9540,N_7272,N_7713);
xnor U9541 (N_9541,N_7213,N_6499);
xnor U9542 (N_9542,N_7623,N_6421);
nor U9543 (N_9543,N_6186,N_7905);
nand U9544 (N_9544,N_7251,N_6170);
or U9545 (N_9545,N_6815,N_7960);
and U9546 (N_9546,N_7757,N_7143);
nor U9547 (N_9547,N_6335,N_7299);
nand U9548 (N_9548,N_7559,N_6563);
xnor U9549 (N_9549,N_6598,N_7569);
and U9550 (N_9550,N_6249,N_7961);
nor U9551 (N_9551,N_7603,N_7404);
nand U9552 (N_9552,N_6251,N_7188);
or U9553 (N_9553,N_7654,N_7290);
nand U9554 (N_9554,N_6659,N_7460);
and U9555 (N_9555,N_7174,N_6161);
nand U9556 (N_9556,N_6294,N_7099);
nand U9557 (N_9557,N_6377,N_6787);
xor U9558 (N_9558,N_6504,N_7995);
nand U9559 (N_9559,N_6841,N_6818);
xnor U9560 (N_9560,N_6896,N_6017);
nor U9561 (N_9561,N_7034,N_6306);
nand U9562 (N_9562,N_7952,N_7233);
nand U9563 (N_9563,N_6467,N_7663);
nand U9564 (N_9564,N_6361,N_6064);
nand U9565 (N_9565,N_6798,N_6873);
nor U9566 (N_9566,N_7796,N_6616);
and U9567 (N_9567,N_6872,N_6537);
xor U9568 (N_9568,N_7928,N_7892);
nand U9569 (N_9569,N_6155,N_7202);
nor U9570 (N_9570,N_7180,N_6523);
and U9571 (N_9571,N_7954,N_7445);
nor U9572 (N_9572,N_6990,N_6596);
or U9573 (N_9573,N_7632,N_7755);
or U9574 (N_9574,N_7206,N_6769);
nor U9575 (N_9575,N_6047,N_6905);
and U9576 (N_9576,N_6402,N_7303);
nand U9577 (N_9577,N_6453,N_6281);
or U9578 (N_9578,N_6618,N_7243);
and U9579 (N_9579,N_6753,N_6340);
xnor U9580 (N_9580,N_6515,N_7210);
xor U9581 (N_9581,N_7677,N_7185);
and U9582 (N_9582,N_7745,N_6775);
xnor U9583 (N_9583,N_6158,N_6282);
nand U9584 (N_9584,N_6254,N_6108);
nor U9585 (N_9585,N_6248,N_7789);
nand U9586 (N_9586,N_6179,N_7889);
nand U9587 (N_9587,N_7838,N_7231);
nand U9588 (N_9588,N_7101,N_7920);
or U9589 (N_9589,N_7878,N_7495);
nor U9590 (N_9590,N_6869,N_7094);
and U9591 (N_9591,N_6035,N_7474);
or U9592 (N_9592,N_6717,N_7605);
or U9593 (N_9593,N_6888,N_6897);
xor U9594 (N_9594,N_6120,N_7843);
nand U9595 (N_9595,N_6482,N_7040);
or U9596 (N_9596,N_7864,N_7223);
nor U9597 (N_9597,N_7319,N_7455);
nand U9598 (N_9598,N_6597,N_6172);
nor U9599 (N_9599,N_6016,N_6779);
or U9600 (N_9600,N_6499,N_6060);
and U9601 (N_9601,N_6413,N_7045);
nand U9602 (N_9602,N_6120,N_7414);
xnor U9603 (N_9603,N_7165,N_6934);
xor U9604 (N_9604,N_6259,N_7703);
xor U9605 (N_9605,N_7605,N_6854);
and U9606 (N_9606,N_7989,N_7747);
or U9607 (N_9607,N_7074,N_7763);
xor U9608 (N_9608,N_6267,N_6142);
or U9609 (N_9609,N_7018,N_7711);
nand U9610 (N_9610,N_7285,N_6900);
and U9611 (N_9611,N_6825,N_6655);
and U9612 (N_9612,N_7265,N_7151);
nand U9613 (N_9613,N_6307,N_6904);
and U9614 (N_9614,N_7004,N_6747);
nor U9615 (N_9615,N_6737,N_6083);
xor U9616 (N_9616,N_7014,N_7027);
xnor U9617 (N_9617,N_7294,N_6598);
nand U9618 (N_9618,N_7767,N_6610);
xnor U9619 (N_9619,N_6614,N_7951);
or U9620 (N_9620,N_7297,N_6282);
and U9621 (N_9621,N_6416,N_6942);
nor U9622 (N_9622,N_7670,N_6529);
xnor U9623 (N_9623,N_6995,N_6142);
nand U9624 (N_9624,N_7453,N_7263);
and U9625 (N_9625,N_6185,N_6631);
nand U9626 (N_9626,N_7894,N_7035);
xor U9627 (N_9627,N_7111,N_6985);
and U9628 (N_9628,N_7704,N_7304);
and U9629 (N_9629,N_6877,N_7970);
nand U9630 (N_9630,N_6404,N_7616);
and U9631 (N_9631,N_7326,N_6350);
nor U9632 (N_9632,N_6276,N_7710);
or U9633 (N_9633,N_7052,N_7174);
or U9634 (N_9634,N_6468,N_6544);
nand U9635 (N_9635,N_6189,N_6928);
and U9636 (N_9636,N_6007,N_7859);
and U9637 (N_9637,N_7471,N_7395);
or U9638 (N_9638,N_7033,N_7580);
and U9639 (N_9639,N_6500,N_6331);
and U9640 (N_9640,N_6605,N_6689);
nand U9641 (N_9641,N_6237,N_6955);
xnor U9642 (N_9642,N_6309,N_6154);
nor U9643 (N_9643,N_6151,N_7816);
xor U9644 (N_9644,N_6719,N_6485);
or U9645 (N_9645,N_7603,N_6181);
or U9646 (N_9646,N_6071,N_6853);
nor U9647 (N_9647,N_7478,N_7595);
xnor U9648 (N_9648,N_7959,N_6884);
nor U9649 (N_9649,N_6016,N_6174);
nor U9650 (N_9650,N_6215,N_6759);
and U9651 (N_9651,N_6466,N_7433);
xor U9652 (N_9652,N_6738,N_6592);
xnor U9653 (N_9653,N_7198,N_6026);
xor U9654 (N_9654,N_6818,N_6487);
nor U9655 (N_9655,N_7479,N_7678);
and U9656 (N_9656,N_6464,N_6115);
nor U9657 (N_9657,N_6702,N_6148);
nand U9658 (N_9658,N_7517,N_6372);
nand U9659 (N_9659,N_6458,N_7386);
and U9660 (N_9660,N_6192,N_6320);
and U9661 (N_9661,N_6043,N_7891);
nand U9662 (N_9662,N_6224,N_6594);
nor U9663 (N_9663,N_7900,N_7402);
nor U9664 (N_9664,N_6415,N_7731);
nor U9665 (N_9665,N_6033,N_6839);
xnor U9666 (N_9666,N_7993,N_7834);
and U9667 (N_9667,N_6626,N_6386);
nor U9668 (N_9668,N_6270,N_7913);
xor U9669 (N_9669,N_6252,N_7229);
or U9670 (N_9670,N_6913,N_7432);
nand U9671 (N_9671,N_6931,N_6625);
or U9672 (N_9672,N_6561,N_6881);
xor U9673 (N_9673,N_6843,N_7494);
and U9674 (N_9674,N_7634,N_6802);
or U9675 (N_9675,N_6319,N_6568);
and U9676 (N_9676,N_6067,N_6704);
or U9677 (N_9677,N_7740,N_6311);
nand U9678 (N_9678,N_6800,N_7334);
and U9679 (N_9679,N_6933,N_6325);
nor U9680 (N_9680,N_6027,N_7729);
nor U9681 (N_9681,N_7670,N_6298);
nor U9682 (N_9682,N_6409,N_7367);
nor U9683 (N_9683,N_6415,N_6848);
nor U9684 (N_9684,N_7218,N_7423);
nand U9685 (N_9685,N_7429,N_7727);
or U9686 (N_9686,N_7396,N_7028);
nor U9687 (N_9687,N_7763,N_7962);
xor U9688 (N_9688,N_6077,N_6448);
xor U9689 (N_9689,N_6996,N_7976);
nor U9690 (N_9690,N_7985,N_7461);
nand U9691 (N_9691,N_6995,N_6239);
xnor U9692 (N_9692,N_6359,N_7266);
or U9693 (N_9693,N_6068,N_6795);
xor U9694 (N_9694,N_7639,N_6799);
and U9695 (N_9695,N_6150,N_7533);
nand U9696 (N_9696,N_6144,N_6156);
nor U9697 (N_9697,N_6166,N_6369);
xnor U9698 (N_9698,N_7768,N_6422);
xor U9699 (N_9699,N_6093,N_7815);
xor U9700 (N_9700,N_6446,N_7045);
and U9701 (N_9701,N_6029,N_7098);
nor U9702 (N_9702,N_6059,N_6108);
and U9703 (N_9703,N_6490,N_6779);
or U9704 (N_9704,N_7396,N_6697);
and U9705 (N_9705,N_6157,N_7499);
or U9706 (N_9706,N_6875,N_7452);
nand U9707 (N_9707,N_6927,N_6555);
nor U9708 (N_9708,N_6160,N_6304);
nor U9709 (N_9709,N_6005,N_6835);
and U9710 (N_9710,N_6915,N_7024);
and U9711 (N_9711,N_7256,N_6487);
nor U9712 (N_9712,N_6097,N_6706);
nand U9713 (N_9713,N_6126,N_7520);
and U9714 (N_9714,N_7455,N_6603);
nor U9715 (N_9715,N_7805,N_6807);
and U9716 (N_9716,N_7262,N_6701);
nor U9717 (N_9717,N_7412,N_7849);
nand U9718 (N_9718,N_6319,N_6304);
and U9719 (N_9719,N_7127,N_7461);
and U9720 (N_9720,N_7200,N_7752);
and U9721 (N_9721,N_7785,N_6975);
nor U9722 (N_9722,N_7541,N_6193);
nand U9723 (N_9723,N_7650,N_6744);
nand U9724 (N_9724,N_6288,N_6316);
and U9725 (N_9725,N_6922,N_7944);
nand U9726 (N_9726,N_7443,N_6280);
nand U9727 (N_9727,N_7850,N_6706);
nor U9728 (N_9728,N_6207,N_7025);
xor U9729 (N_9729,N_7453,N_6147);
and U9730 (N_9730,N_6796,N_6568);
or U9731 (N_9731,N_7636,N_7538);
nand U9732 (N_9732,N_6605,N_6408);
and U9733 (N_9733,N_6927,N_6622);
and U9734 (N_9734,N_6700,N_7108);
or U9735 (N_9735,N_7060,N_6016);
or U9736 (N_9736,N_6401,N_7175);
xor U9737 (N_9737,N_7364,N_7657);
and U9738 (N_9738,N_6083,N_7748);
and U9739 (N_9739,N_6601,N_6253);
nand U9740 (N_9740,N_7288,N_6154);
or U9741 (N_9741,N_6931,N_6120);
and U9742 (N_9742,N_6152,N_7618);
nand U9743 (N_9743,N_6006,N_6373);
xor U9744 (N_9744,N_6717,N_7526);
xnor U9745 (N_9745,N_6781,N_6413);
or U9746 (N_9746,N_7294,N_6403);
nand U9747 (N_9747,N_7046,N_7461);
nand U9748 (N_9748,N_7338,N_6589);
and U9749 (N_9749,N_6616,N_7671);
or U9750 (N_9750,N_7113,N_6345);
and U9751 (N_9751,N_7838,N_7227);
or U9752 (N_9752,N_7288,N_7594);
xor U9753 (N_9753,N_6894,N_7159);
and U9754 (N_9754,N_7651,N_6334);
nor U9755 (N_9755,N_6527,N_7667);
nand U9756 (N_9756,N_7148,N_6879);
nand U9757 (N_9757,N_6699,N_7868);
nand U9758 (N_9758,N_7335,N_7373);
or U9759 (N_9759,N_6662,N_6293);
or U9760 (N_9760,N_7615,N_6256);
nor U9761 (N_9761,N_7268,N_7269);
xnor U9762 (N_9762,N_6238,N_7417);
nor U9763 (N_9763,N_6389,N_7920);
and U9764 (N_9764,N_7136,N_7599);
and U9765 (N_9765,N_6894,N_7115);
nand U9766 (N_9766,N_7132,N_6259);
or U9767 (N_9767,N_7543,N_7363);
and U9768 (N_9768,N_6220,N_7498);
nand U9769 (N_9769,N_7972,N_6727);
nor U9770 (N_9770,N_6862,N_7194);
xnor U9771 (N_9771,N_6507,N_6375);
nand U9772 (N_9772,N_6739,N_6836);
xor U9773 (N_9773,N_7296,N_7425);
nor U9774 (N_9774,N_7358,N_6014);
xor U9775 (N_9775,N_6801,N_6079);
nand U9776 (N_9776,N_7306,N_7574);
xor U9777 (N_9777,N_6549,N_6544);
xor U9778 (N_9778,N_7454,N_6212);
and U9779 (N_9779,N_6451,N_6056);
and U9780 (N_9780,N_7901,N_6462);
nor U9781 (N_9781,N_6506,N_7425);
nor U9782 (N_9782,N_6052,N_7685);
and U9783 (N_9783,N_6960,N_7755);
nand U9784 (N_9784,N_7897,N_7392);
or U9785 (N_9785,N_7755,N_7454);
or U9786 (N_9786,N_6927,N_6175);
and U9787 (N_9787,N_7678,N_7077);
and U9788 (N_9788,N_7165,N_6459);
or U9789 (N_9789,N_6472,N_6872);
xnor U9790 (N_9790,N_7716,N_7931);
or U9791 (N_9791,N_7018,N_6106);
nand U9792 (N_9792,N_7289,N_6158);
xnor U9793 (N_9793,N_6484,N_7092);
nor U9794 (N_9794,N_7603,N_7502);
or U9795 (N_9795,N_7839,N_7300);
nor U9796 (N_9796,N_7092,N_6145);
nor U9797 (N_9797,N_7807,N_6425);
or U9798 (N_9798,N_7788,N_7317);
xnor U9799 (N_9799,N_7976,N_7132);
or U9800 (N_9800,N_7879,N_6622);
nor U9801 (N_9801,N_7276,N_7407);
nand U9802 (N_9802,N_7548,N_7173);
nand U9803 (N_9803,N_7004,N_7566);
or U9804 (N_9804,N_6006,N_7842);
nor U9805 (N_9805,N_7071,N_6287);
or U9806 (N_9806,N_6510,N_7845);
and U9807 (N_9807,N_6490,N_6770);
nand U9808 (N_9808,N_6289,N_6150);
nor U9809 (N_9809,N_6999,N_7623);
or U9810 (N_9810,N_6670,N_6493);
and U9811 (N_9811,N_7503,N_6073);
nand U9812 (N_9812,N_6985,N_6712);
xor U9813 (N_9813,N_7008,N_6871);
xor U9814 (N_9814,N_6843,N_7859);
xor U9815 (N_9815,N_7844,N_7380);
nor U9816 (N_9816,N_7984,N_7931);
and U9817 (N_9817,N_6554,N_6971);
and U9818 (N_9818,N_6281,N_6967);
and U9819 (N_9819,N_7027,N_7186);
or U9820 (N_9820,N_6453,N_7125);
and U9821 (N_9821,N_6778,N_7262);
xor U9822 (N_9822,N_6876,N_6267);
nand U9823 (N_9823,N_7713,N_6731);
and U9824 (N_9824,N_7632,N_6168);
or U9825 (N_9825,N_6293,N_7423);
nor U9826 (N_9826,N_6763,N_7264);
nand U9827 (N_9827,N_6871,N_6424);
nand U9828 (N_9828,N_6196,N_6522);
nor U9829 (N_9829,N_6398,N_7211);
and U9830 (N_9830,N_6730,N_7414);
nor U9831 (N_9831,N_7850,N_6929);
and U9832 (N_9832,N_6148,N_7080);
or U9833 (N_9833,N_6303,N_6503);
nand U9834 (N_9834,N_7626,N_7599);
nand U9835 (N_9835,N_7626,N_6280);
or U9836 (N_9836,N_7712,N_7228);
nor U9837 (N_9837,N_7283,N_7557);
nor U9838 (N_9838,N_7575,N_6353);
nor U9839 (N_9839,N_7711,N_7429);
or U9840 (N_9840,N_6613,N_7821);
or U9841 (N_9841,N_6462,N_6500);
and U9842 (N_9842,N_6809,N_6107);
and U9843 (N_9843,N_7048,N_6513);
xnor U9844 (N_9844,N_6225,N_7121);
and U9845 (N_9845,N_7661,N_7927);
nand U9846 (N_9846,N_7832,N_6528);
and U9847 (N_9847,N_7436,N_7644);
and U9848 (N_9848,N_7584,N_7021);
xnor U9849 (N_9849,N_7830,N_7429);
nand U9850 (N_9850,N_6020,N_7662);
xnor U9851 (N_9851,N_7006,N_7066);
xor U9852 (N_9852,N_7666,N_7298);
nand U9853 (N_9853,N_7402,N_6564);
nor U9854 (N_9854,N_6912,N_7834);
and U9855 (N_9855,N_6555,N_6824);
nand U9856 (N_9856,N_6492,N_7196);
and U9857 (N_9857,N_6222,N_6393);
and U9858 (N_9858,N_6650,N_7057);
and U9859 (N_9859,N_6416,N_6652);
xnor U9860 (N_9860,N_6464,N_7720);
nor U9861 (N_9861,N_6891,N_7176);
xnor U9862 (N_9862,N_6917,N_6632);
and U9863 (N_9863,N_6776,N_6757);
xnor U9864 (N_9864,N_6362,N_7200);
and U9865 (N_9865,N_7294,N_7714);
nand U9866 (N_9866,N_7073,N_7601);
nor U9867 (N_9867,N_6017,N_6433);
or U9868 (N_9868,N_7620,N_7236);
xnor U9869 (N_9869,N_7877,N_6494);
or U9870 (N_9870,N_7823,N_6402);
or U9871 (N_9871,N_7688,N_7710);
nand U9872 (N_9872,N_6640,N_6139);
or U9873 (N_9873,N_6864,N_7815);
nor U9874 (N_9874,N_7117,N_7947);
or U9875 (N_9875,N_6246,N_7810);
or U9876 (N_9876,N_7965,N_7890);
nand U9877 (N_9877,N_6987,N_7574);
nor U9878 (N_9878,N_6954,N_7134);
and U9879 (N_9879,N_7148,N_6090);
or U9880 (N_9880,N_6328,N_6344);
xnor U9881 (N_9881,N_7039,N_6400);
nand U9882 (N_9882,N_6245,N_6275);
nand U9883 (N_9883,N_7349,N_6555);
nand U9884 (N_9884,N_7300,N_7171);
or U9885 (N_9885,N_6365,N_6306);
nand U9886 (N_9886,N_7716,N_6893);
or U9887 (N_9887,N_7971,N_7406);
xor U9888 (N_9888,N_7561,N_6726);
xor U9889 (N_9889,N_7630,N_7204);
and U9890 (N_9890,N_7535,N_6323);
nand U9891 (N_9891,N_7807,N_7075);
nand U9892 (N_9892,N_7918,N_6051);
xor U9893 (N_9893,N_6941,N_6118);
and U9894 (N_9894,N_7133,N_6884);
or U9895 (N_9895,N_7307,N_6894);
and U9896 (N_9896,N_7276,N_6641);
and U9897 (N_9897,N_7137,N_6467);
xor U9898 (N_9898,N_6433,N_6159);
and U9899 (N_9899,N_6165,N_7305);
or U9900 (N_9900,N_7686,N_6529);
and U9901 (N_9901,N_6823,N_6297);
and U9902 (N_9902,N_6912,N_7242);
nor U9903 (N_9903,N_6278,N_6318);
nor U9904 (N_9904,N_7950,N_7049);
nand U9905 (N_9905,N_7628,N_6511);
nand U9906 (N_9906,N_7075,N_6326);
xnor U9907 (N_9907,N_7140,N_7804);
nor U9908 (N_9908,N_6976,N_6691);
or U9909 (N_9909,N_7893,N_7312);
and U9910 (N_9910,N_6272,N_6845);
nand U9911 (N_9911,N_6737,N_7683);
or U9912 (N_9912,N_7440,N_6153);
nor U9913 (N_9913,N_7383,N_7352);
nor U9914 (N_9914,N_6775,N_7889);
or U9915 (N_9915,N_6910,N_7257);
and U9916 (N_9916,N_6923,N_6308);
xnor U9917 (N_9917,N_6270,N_7673);
xor U9918 (N_9918,N_7452,N_6772);
or U9919 (N_9919,N_7924,N_7700);
nor U9920 (N_9920,N_7212,N_6071);
nor U9921 (N_9921,N_6250,N_6496);
nand U9922 (N_9922,N_7154,N_7507);
or U9923 (N_9923,N_6773,N_7130);
xnor U9924 (N_9924,N_6293,N_7006);
and U9925 (N_9925,N_7736,N_7592);
and U9926 (N_9926,N_6021,N_6711);
and U9927 (N_9927,N_6977,N_7553);
nor U9928 (N_9928,N_6631,N_6971);
or U9929 (N_9929,N_6754,N_6532);
nor U9930 (N_9930,N_6330,N_7521);
nand U9931 (N_9931,N_7117,N_6525);
and U9932 (N_9932,N_6937,N_7580);
xnor U9933 (N_9933,N_6523,N_6501);
nand U9934 (N_9934,N_6019,N_7086);
xnor U9935 (N_9935,N_7877,N_7026);
or U9936 (N_9936,N_7230,N_7341);
nor U9937 (N_9937,N_6059,N_6662);
and U9938 (N_9938,N_7158,N_7612);
and U9939 (N_9939,N_7168,N_7960);
or U9940 (N_9940,N_7418,N_6794);
nor U9941 (N_9941,N_6527,N_7949);
xnor U9942 (N_9942,N_6494,N_6764);
nand U9943 (N_9943,N_7405,N_7254);
nor U9944 (N_9944,N_7122,N_6716);
and U9945 (N_9945,N_6315,N_7715);
xnor U9946 (N_9946,N_6106,N_6635);
nand U9947 (N_9947,N_7078,N_6937);
and U9948 (N_9948,N_6093,N_7947);
nor U9949 (N_9949,N_7707,N_7575);
or U9950 (N_9950,N_7753,N_7072);
nor U9951 (N_9951,N_6436,N_7650);
nand U9952 (N_9952,N_7538,N_7872);
or U9953 (N_9953,N_6715,N_6841);
xnor U9954 (N_9954,N_7345,N_7232);
or U9955 (N_9955,N_6050,N_7816);
or U9956 (N_9956,N_7219,N_7913);
xor U9957 (N_9957,N_6012,N_6521);
and U9958 (N_9958,N_7127,N_6504);
nor U9959 (N_9959,N_6223,N_7598);
nand U9960 (N_9960,N_6755,N_6305);
xnor U9961 (N_9961,N_7904,N_6172);
and U9962 (N_9962,N_7683,N_6236);
nor U9963 (N_9963,N_7838,N_7979);
and U9964 (N_9964,N_6711,N_7951);
nand U9965 (N_9965,N_7199,N_6298);
nand U9966 (N_9966,N_7350,N_7018);
xor U9967 (N_9967,N_7293,N_7553);
and U9968 (N_9968,N_6491,N_6025);
and U9969 (N_9969,N_6218,N_6450);
or U9970 (N_9970,N_7667,N_7197);
or U9971 (N_9971,N_6420,N_7233);
and U9972 (N_9972,N_7483,N_7793);
and U9973 (N_9973,N_7324,N_6713);
or U9974 (N_9974,N_6603,N_6567);
and U9975 (N_9975,N_7385,N_6983);
nor U9976 (N_9976,N_6809,N_6079);
nand U9977 (N_9977,N_7553,N_7060);
and U9978 (N_9978,N_6783,N_6229);
nor U9979 (N_9979,N_6777,N_6431);
xor U9980 (N_9980,N_6355,N_6177);
xor U9981 (N_9981,N_7932,N_7767);
nor U9982 (N_9982,N_7662,N_6740);
nor U9983 (N_9983,N_6459,N_7284);
nor U9984 (N_9984,N_7711,N_6826);
nor U9985 (N_9985,N_6013,N_6230);
or U9986 (N_9986,N_7239,N_6156);
and U9987 (N_9987,N_7234,N_6622);
xnor U9988 (N_9988,N_7616,N_7556);
nor U9989 (N_9989,N_7738,N_7491);
nor U9990 (N_9990,N_7715,N_7278);
nor U9991 (N_9991,N_7113,N_7773);
and U9992 (N_9992,N_6889,N_6234);
nor U9993 (N_9993,N_6294,N_7072);
nor U9994 (N_9994,N_7828,N_7776);
or U9995 (N_9995,N_6650,N_7677);
nand U9996 (N_9996,N_7258,N_7365);
xor U9997 (N_9997,N_7183,N_6372);
xor U9998 (N_9998,N_7612,N_6127);
nor U9999 (N_9999,N_6841,N_7001);
and U10000 (N_10000,N_9787,N_9517);
and U10001 (N_10001,N_9217,N_8683);
and U10002 (N_10002,N_9982,N_8153);
xor U10003 (N_10003,N_9620,N_8528);
or U10004 (N_10004,N_8500,N_9151);
nor U10005 (N_10005,N_9014,N_8251);
nand U10006 (N_10006,N_9247,N_8167);
or U10007 (N_10007,N_8940,N_9958);
xor U10008 (N_10008,N_9715,N_9726);
and U10009 (N_10009,N_9945,N_8836);
nor U10010 (N_10010,N_8618,N_8448);
nor U10011 (N_10011,N_8177,N_9834);
or U10012 (N_10012,N_8484,N_9328);
and U10013 (N_10013,N_8865,N_9667);
and U10014 (N_10014,N_9510,N_8914);
xnor U10015 (N_10015,N_8267,N_9224);
nand U10016 (N_10016,N_8330,N_9680);
xor U10017 (N_10017,N_8212,N_9756);
nor U10018 (N_10018,N_8762,N_8269);
nand U10019 (N_10019,N_8975,N_8272);
or U10020 (N_10020,N_8199,N_8846);
nor U10021 (N_10021,N_8591,N_8634);
nor U10022 (N_10022,N_9216,N_9229);
nor U10023 (N_10023,N_9366,N_9985);
nor U10024 (N_10024,N_8687,N_9287);
xnor U10025 (N_10025,N_9896,N_8410);
or U10026 (N_10026,N_9949,N_8315);
and U10027 (N_10027,N_8635,N_9649);
nor U10028 (N_10028,N_8572,N_9969);
nand U10029 (N_10029,N_9874,N_8690);
and U10030 (N_10030,N_9955,N_9487);
or U10031 (N_10031,N_8653,N_9137);
nor U10032 (N_10032,N_9314,N_9181);
or U10033 (N_10033,N_8499,N_9763);
and U10034 (N_10034,N_9677,N_9850);
nor U10035 (N_10035,N_9994,N_9920);
or U10036 (N_10036,N_9263,N_8682);
nand U10037 (N_10037,N_8501,N_9389);
nor U10038 (N_10038,N_9662,N_9999);
and U10039 (N_10039,N_9924,N_8818);
nor U10040 (N_10040,N_8884,N_8899);
and U10041 (N_10041,N_9296,N_9978);
or U10042 (N_10042,N_8761,N_9555);
xnor U10043 (N_10043,N_9436,N_8502);
and U10044 (N_10044,N_9091,N_9722);
nor U10045 (N_10045,N_9461,N_8915);
nand U10046 (N_10046,N_8783,N_8360);
nand U10047 (N_10047,N_8446,N_8142);
and U10048 (N_10048,N_9133,N_8790);
nor U10049 (N_10049,N_8489,N_8747);
and U10050 (N_10050,N_9377,N_9940);
nand U10051 (N_10051,N_9149,N_8609);
or U10052 (N_10052,N_9718,N_9541);
and U10053 (N_10053,N_9212,N_8912);
or U10054 (N_10054,N_9188,N_9866);
or U10055 (N_10055,N_8900,N_9488);
xnor U10056 (N_10056,N_9663,N_9456);
or U10057 (N_10057,N_9672,N_8325);
xor U10058 (N_10058,N_8978,N_9753);
and U10059 (N_10059,N_9141,N_9407);
xnor U10060 (N_10060,N_9466,N_8195);
or U10061 (N_10061,N_8028,N_8281);
nand U10062 (N_10062,N_8359,N_9597);
nor U10063 (N_10063,N_9150,N_9077);
nand U10064 (N_10064,N_9975,N_9085);
or U10065 (N_10065,N_8666,N_8808);
nor U10066 (N_10066,N_8479,N_8172);
and U10067 (N_10067,N_9401,N_8292);
or U10068 (N_10068,N_8497,N_8873);
or U10069 (N_10069,N_8010,N_9479);
nand U10070 (N_10070,N_8972,N_8693);
nand U10071 (N_10071,N_8245,N_8045);
or U10072 (N_10072,N_9725,N_9180);
nor U10073 (N_10073,N_8749,N_9024);
or U10074 (N_10074,N_9724,N_9897);
nor U10075 (N_10075,N_8151,N_9552);
xnor U10076 (N_10076,N_9121,N_9509);
nand U10077 (N_10077,N_9804,N_9573);
nor U10078 (N_10078,N_9334,N_8671);
xor U10079 (N_10079,N_8897,N_9194);
or U10080 (N_10080,N_9757,N_9255);
nand U10081 (N_10081,N_9749,N_8525);
xnor U10082 (N_10082,N_8119,N_9010);
or U10083 (N_10083,N_8435,N_8011);
and U10084 (N_10084,N_8298,N_8816);
xnor U10085 (N_10085,N_8833,N_8530);
and U10086 (N_10086,N_9388,N_9412);
and U10087 (N_10087,N_9415,N_8120);
xnor U10088 (N_10088,N_8539,N_9950);
xor U10089 (N_10089,N_9343,N_8411);
and U10090 (N_10090,N_9326,N_8799);
and U10091 (N_10091,N_8506,N_8349);
or U10092 (N_10092,N_9965,N_9571);
xnor U10093 (N_10093,N_8146,N_8291);
nand U10094 (N_10094,N_9867,N_8161);
and U10095 (N_10095,N_9111,N_9125);
nor U10096 (N_10096,N_8384,N_9136);
and U10097 (N_10097,N_9530,N_8989);
nor U10098 (N_10098,N_8089,N_8728);
xor U10099 (N_10099,N_8218,N_8821);
nand U10100 (N_10100,N_8961,N_9475);
or U10101 (N_10101,N_9392,N_9972);
nand U10102 (N_10102,N_9645,N_9173);
or U10103 (N_10103,N_8936,N_8234);
or U10104 (N_10104,N_8434,N_9878);
and U10105 (N_10105,N_9235,N_8594);
nand U10106 (N_10106,N_9183,N_8152);
xnor U10107 (N_10107,N_9588,N_9813);
nand U10108 (N_10108,N_9886,N_8565);
and U10109 (N_10109,N_9685,N_8829);
or U10110 (N_10110,N_8731,N_8741);
nand U10111 (N_10111,N_9175,N_8176);
xor U10112 (N_10112,N_8187,N_8573);
and U10113 (N_10113,N_9448,N_8304);
and U10114 (N_10114,N_9186,N_8110);
nor U10115 (N_10115,N_8454,N_9058);
nand U10116 (N_10116,N_8886,N_9963);
and U10117 (N_10117,N_9852,N_8283);
or U10118 (N_10118,N_8824,N_9786);
xnor U10119 (N_10119,N_9554,N_8381);
nand U10120 (N_10120,N_8813,N_8612);
or U10121 (N_10121,N_8297,N_8826);
nand U10122 (N_10122,N_9210,N_8467);
nand U10123 (N_10123,N_8070,N_9073);
xor U10124 (N_10124,N_9933,N_8585);
nor U10125 (N_10125,N_8405,N_9634);
and U10126 (N_10126,N_8705,N_9642);
nor U10127 (N_10127,N_9030,N_9257);
nor U10128 (N_10128,N_9550,N_8703);
or U10129 (N_10129,N_9286,N_9721);
nand U10130 (N_10130,N_8850,N_9489);
nor U10131 (N_10131,N_9609,N_9581);
nor U10132 (N_10132,N_9013,N_8803);
and U10133 (N_10133,N_9311,N_8845);
nand U10134 (N_10134,N_8536,N_9900);
xnor U10135 (N_10135,N_8382,N_9616);
xnor U10136 (N_10136,N_9157,N_8748);
xor U10137 (N_10137,N_8664,N_9790);
and U10138 (N_10138,N_9929,N_9665);
xnor U10139 (N_10139,N_9386,N_9692);
and U10140 (N_10140,N_9041,N_8809);
and U10141 (N_10141,N_9840,N_9054);
nand U10142 (N_10142,N_8582,N_8510);
nand U10143 (N_10143,N_8851,N_8593);
and U10144 (N_10144,N_9827,N_8495);
or U10145 (N_10145,N_8346,N_8812);
nor U10146 (N_10146,N_9538,N_9486);
xnor U10147 (N_10147,N_8050,N_9460);
nand U10148 (N_10148,N_9281,N_8383);
or U10149 (N_10149,N_9223,N_8995);
xnor U10150 (N_10150,N_8576,N_8229);
or U10151 (N_10151,N_9577,N_9791);
nor U10152 (N_10152,N_8196,N_9087);
or U10153 (N_10153,N_9274,N_9893);
xnor U10154 (N_10154,N_9008,N_8137);
nor U10155 (N_10155,N_9711,N_8008);
and U10156 (N_10156,N_8774,N_9331);
nand U10157 (N_10157,N_8546,N_8772);
and U10158 (N_10158,N_9011,N_8643);
nor U10159 (N_10159,N_9469,N_8859);
nand U10160 (N_10160,N_8994,N_8586);
nand U10161 (N_10161,N_8584,N_9098);
nand U10162 (N_10162,N_9355,N_8885);
nor U10163 (N_10163,N_8159,N_9807);
nand U10164 (N_10164,N_9953,N_8621);
nor U10165 (N_10165,N_8453,N_9862);
xnor U10166 (N_10166,N_9822,N_9587);
nand U10167 (N_10167,N_8680,N_8337);
and U10168 (N_10168,N_9864,N_9444);
nor U10169 (N_10169,N_9164,N_9214);
nand U10170 (N_10170,N_9481,N_9272);
nand U10171 (N_10171,N_8108,N_9092);
or U10172 (N_10172,N_8001,N_8751);
or U10173 (N_10173,N_8615,N_8314);
or U10174 (N_10174,N_9176,N_9567);
nor U10175 (N_10175,N_8352,N_9513);
or U10176 (N_10176,N_8319,N_9131);
xnor U10177 (N_10177,N_9166,N_8601);
and U10178 (N_10178,N_9047,N_8758);
and U10179 (N_10179,N_8939,N_8475);
or U10180 (N_10180,N_9764,N_9076);
xnor U10181 (N_10181,N_9037,N_8165);
nand U10182 (N_10182,N_8563,N_9310);
or U10183 (N_10183,N_8396,N_9584);
xnor U10184 (N_10184,N_8947,N_8745);
nor U10185 (N_10185,N_9171,N_8872);
and U10186 (N_10186,N_9497,N_9745);
xor U10187 (N_10187,N_8227,N_9391);
nand U10188 (N_10188,N_8347,N_8583);
or U10189 (N_10189,N_8681,N_8131);
or U10190 (N_10190,N_9796,N_8060);
xnor U10191 (N_10191,N_9032,N_8094);
or U10192 (N_10192,N_9514,N_8350);
or U10193 (N_10193,N_9371,N_8778);
or U10194 (N_10194,N_8037,N_9678);
or U10195 (N_10195,N_8169,N_8869);
and U10196 (N_10196,N_8400,N_8521);
xor U10197 (N_10197,N_8672,N_9633);
nand U10198 (N_10198,N_9707,N_9907);
or U10199 (N_10199,N_8775,N_8397);
and U10200 (N_10200,N_9873,N_9516);
xor U10201 (N_10201,N_8605,N_9580);
nand U10202 (N_10202,N_8898,N_8160);
nor U10203 (N_10203,N_9204,N_8852);
nor U10204 (N_10204,N_9789,N_8374);
and U10205 (N_10205,N_8787,N_9779);
nor U10206 (N_10206,N_9101,N_8599);
nand U10207 (N_10207,N_9705,N_9062);
xor U10208 (N_10208,N_9113,N_9781);
nor U10209 (N_10209,N_8014,N_8266);
nor U10210 (N_10210,N_9921,N_8607);
nor U10211 (N_10211,N_9848,N_8064);
and U10212 (N_10212,N_9433,N_9851);
or U10213 (N_10213,N_8622,N_9653);
and U10214 (N_10214,N_9492,N_8999);
and U10215 (N_10215,N_8162,N_9123);
xor U10216 (N_10216,N_8181,N_9983);
xnor U10217 (N_10217,N_8923,N_9564);
xor U10218 (N_10218,N_9413,N_9241);
nor U10219 (N_10219,N_9674,N_8318);
and U10220 (N_10220,N_8966,N_9358);
and U10221 (N_10221,N_8560,N_9376);
and U10222 (N_10222,N_8823,N_8922);
and U10223 (N_10223,N_8764,N_8219);
nor U10224 (N_10224,N_9209,N_9624);
and U10225 (N_10225,N_9467,N_8825);
nand U10226 (N_10226,N_9626,N_9454);
nand U10227 (N_10227,N_9539,N_9484);
nor U10228 (N_10228,N_8600,N_9312);
xor U10229 (N_10229,N_8633,N_8112);
xor U10230 (N_10230,N_8684,N_9816);
xnor U10231 (N_10231,N_8240,N_9207);
or U10232 (N_10232,N_8048,N_9061);
nor U10233 (N_10233,N_9892,N_9941);
or U10234 (N_10234,N_9198,N_9040);
and U10235 (N_10235,N_9419,N_9035);
nand U10236 (N_10236,N_8876,N_9687);
or U10237 (N_10237,N_8306,N_8953);
nor U10238 (N_10238,N_9315,N_8930);
or U10239 (N_10239,N_9938,N_8678);
or U10240 (N_10240,N_8648,N_8597);
and U10241 (N_10241,N_9547,N_8675);
nand U10242 (N_10242,N_9503,N_8193);
xor U10243 (N_10243,N_9915,N_9110);
nand U10244 (N_10244,N_8494,N_8676);
nor U10245 (N_10245,N_9797,N_9522);
nand U10246 (N_10246,N_8450,N_8777);
xor U10247 (N_10247,N_9540,N_8598);
nand U10248 (N_10248,N_8355,N_8614);
xor U10249 (N_10249,N_8083,N_8403);
xnor U10250 (N_10250,N_8230,N_9440);
and U10251 (N_10251,N_9285,N_9325);
or U10252 (N_10252,N_9846,N_9890);
or U10253 (N_10253,N_9382,N_8716);
xnor U10254 (N_10254,N_9277,N_9565);
nor U10255 (N_10255,N_9868,N_9189);
or U10256 (N_10256,N_8638,N_9364);
nor U10257 (N_10257,N_8562,N_9424);
or U10258 (N_10258,N_8882,N_9780);
nor U10259 (N_10259,N_9954,N_9278);
nor U10260 (N_10260,N_8039,N_8099);
xor U10261 (N_10261,N_9105,N_9420);
nor U10262 (N_10262,N_9720,N_8895);
or U10263 (N_10263,N_8575,N_8093);
xnor U10264 (N_10264,N_9772,N_9283);
nor U10265 (N_10265,N_9346,N_9269);
nand U10266 (N_10266,N_8458,N_8340);
or U10267 (N_10267,N_8144,N_9462);
xor U10268 (N_10268,N_8984,N_8461);
nor U10269 (N_10269,N_8451,N_9069);
nand U10270 (N_10270,N_9345,N_8333);
xor U10271 (N_10271,N_8721,N_9174);
and U10272 (N_10272,N_8848,N_8827);
nor U10273 (N_10273,N_8373,N_8545);
xor U10274 (N_10274,N_8116,N_9821);
nor U10275 (N_10275,N_9396,N_9882);
nor U10276 (N_10276,N_9064,N_9519);
and U10277 (N_10277,N_8431,N_9908);
nor U10278 (N_10278,N_8619,N_8854);
nand U10279 (N_10279,N_9059,N_9876);
nand U10280 (N_10280,N_8233,N_8965);
xnor U10281 (N_10281,N_9323,N_9844);
nand U10282 (N_10282,N_9022,N_8077);
nand U10283 (N_10283,N_9195,N_8316);
xor U10284 (N_10284,N_9544,N_9952);
and U10285 (N_10285,N_9421,N_9585);
nor U10286 (N_10286,N_9109,N_9880);
xor U10287 (N_10287,N_8955,N_8471);
nand U10288 (N_10288,N_9794,N_8921);
xor U10289 (N_10289,N_9701,N_9613);
nor U10290 (N_10290,N_9398,N_9528);
and U10291 (N_10291,N_8202,N_9534);
nor U10292 (N_10292,N_8727,N_8910);
nor U10293 (N_10293,N_8058,N_9138);
or U10294 (N_10294,N_8017,N_8065);
xnor U10295 (N_10295,N_8868,N_8265);
and U10296 (N_10296,N_9365,N_8071);
xor U10297 (N_10297,N_8136,N_8487);
or U10298 (N_10298,N_8725,N_8069);
or U10299 (N_10299,N_9055,N_9853);
or U10300 (N_10300,N_8127,N_9504);
nand U10301 (N_10301,N_8481,N_9622);
nor U10302 (N_10302,N_9230,N_9535);
nor U10303 (N_10303,N_9548,N_8656);
and U10304 (N_10304,N_9934,N_9858);
nor U10305 (N_10305,N_9993,N_9758);
xnor U10306 (N_10306,N_8553,N_8279);
nand U10307 (N_10307,N_9927,N_8857);
xor U10308 (N_10308,N_8205,N_8581);
or U10309 (N_10309,N_9192,N_9379);
nand U10310 (N_10310,N_9911,N_8055);
nand U10311 (N_10311,N_8505,N_8709);
nor U10312 (N_10312,N_8754,N_8466);
nor U10313 (N_10313,N_9784,N_8990);
nor U10314 (N_10314,N_9148,N_8765);
or U10315 (N_10315,N_9575,N_8858);
or U10316 (N_10316,N_8263,N_9308);
xnor U10317 (N_10317,N_8192,N_9464);
nor U10318 (N_10318,N_8012,N_9637);
and U10319 (N_10319,N_9956,N_8490);
nor U10320 (N_10320,N_9778,N_8423);
nor U10321 (N_10321,N_8225,N_9818);
nor U10322 (N_10322,N_8832,N_8928);
or U10323 (N_10323,N_9276,N_9349);
xor U10324 (N_10324,N_9191,N_9727);
or U10325 (N_10325,N_8356,N_8773);
or U10326 (N_10326,N_8704,N_9165);
nand U10327 (N_10327,N_9002,N_9754);
nor U10328 (N_10328,N_9671,N_8617);
and U10329 (N_10329,N_8051,N_8323);
nor U10330 (N_10330,N_9177,N_8086);
or U10331 (N_10331,N_8085,N_9390);
and U10332 (N_10332,N_8209,N_9144);
and U10333 (N_10333,N_8201,N_9158);
nor U10334 (N_10334,N_8548,N_9583);
nand U10335 (N_10335,N_9700,N_9748);
or U10336 (N_10336,N_9704,N_9747);
or U10337 (N_10337,N_8157,N_8270);
nor U10338 (N_10338,N_8753,N_9658);
xor U10339 (N_10339,N_9211,N_9738);
xnor U10340 (N_10340,N_9869,N_9118);
nor U10341 (N_10341,N_8075,N_8061);
nand U10342 (N_10342,N_9805,N_8103);
xnor U10343 (N_10343,N_8444,N_9036);
and U10344 (N_10344,N_9028,N_8968);
xnor U10345 (N_10345,N_8128,N_9072);
and U10346 (N_10346,N_8519,N_9561);
or U10347 (N_10347,N_8188,N_8121);
xnor U10348 (N_10348,N_9162,N_8026);
xnor U10349 (N_10349,N_8996,N_9708);
nor U10350 (N_10350,N_9712,N_9317);
and U10351 (N_10351,N_9339,N_8511);
or U10352 (N_10352,N_8880,N_9361);
and U10353 (N_10353,N_8300,N_9341);
xnor U10354 (N_10354,N_8973,N_8543);
nand U10355 (N_10355,N_8566,N_8784);
xor U10356 (N_10356,N_8210,N_8134);
nor U10357 (N_10357,N_8630,N_8529);
or U10358 (N_10358,N_9843,N_8637);
or U10359 (N_10359,N_8054,N_9429);
nand U10360 (N_10360,N_9053,N_9643);
or U10361 (N_10361,N_8062,N_9065);
nand U10362 (N_10362,N_8059,N_8290);
xor U10363 (N_10363,N_9473,N_8455);
xor U10364 (N_10364,N_8864,N_8009);
xnor U10365 (N_10365,N_9861,N_8805);
and U10366 (N_10366,N_8387,N_8567);
and U10367 (N_10367,N_9447,N_8485);
xnor U10368 (N_10368,N_9208,N_8792);
nand U10369 (N_10369,N_8712,N_8433);
nand U10370 (N_10370,N_9572,N_8399);
and U10371 (N_10371,N_8655,N_9172);
nor U10372 (N_10372,N_8372,N_9380);
nand U10373 (N_10373,N_9000,N_8236);
xor U10374 (N_10374,N_9696,N_8508);
or U10375 (N_10375,N_9351,N_8221);
nor U10376 (N_10376,N_8022,N_8215);
nand U10377 (N_10377,N_8688,N_9134);
xor U10378 (N_10378,N_9179,N_9515);
and U10379 (N_10379,N_8322,N_8421);
or U10380 (N_10380,N_8424,N_9847);
nor U10381 (N_10381,N_9236,N_9342);
or U10382 (N_10382,N_9320,N_8393);
or U10383 (N_10383,N_9114,N_9266);
or U10384 (N_10384,N_9332,N_8742);
nor U10385 (N_10385,N_9683,N_9819);
and U10386 (N_10386,N_8053,N_9012);
nor U10387 (N_10387,N_8154,N_9648);
and U10388 (N_10388,N_9883,N_8997);
nor U10389 (N_10389,N_8420,N_8588);
nand U10390 (N_10390,N_9742,N_8960);
nand U10391 (N_10391,N_8534,N_8568);
nand U10392 (N_10392,N_8354,N_8538);
or U10393 (N_10393,N_9291,N_9080);
and U10394 (N_10394,N_8235,N_8875);
nand U10395 (N_10395,N_9001,N_9056);
and U10396 (N_10396,N_9576,N_8697);
nand U10397 (N_10397,N_8685,N_9679);
or U10398 (N_10398,N_8324,N_9566);
xnor U10399 (N_10399,N_8604,N_8043);
nand U10400 (N_10400,N_8478,N_8906);
and U10401 (N_10401,N_8213,N_9295);
or U10402 (N_10402,N_9673,N_8351);
or U10403 (N_10403,N_8925,N_9232);
or U10404 (N_10404,N_9508,N_8677);
xor U10405 (N_10405,N_8124,N_9218);
nand U10406 (N_10406,N_8920,N_9803);
xnor U10407 (N_10407,N_9124,N_9330);
or U10408 (N_10408,N_8927,N_8312);
nand U10409 (N_10409,N_8719,N_9525);
or U10410 (N_10410,N_8881,N_8830);
and U10411 (N_10411,N_8770,N_8517);
nor U10412 (N_10412,N_9155,N_9045);
and U10413 (N_10413,N_8610,N_9130);
nor U10414 (N_10414,N_8156,N_8038);
nor U10415 (N_10415,N_9455,N_9215);
or U10416 (N_10416,N_8867,N_9226);
xor U10417 (N_10417,N_8004,N_8926);
nor U10418 (N_10418,N_9855,N_9783);
or U10419 (N_10419,N_9106,N_8133);
nand U10420 (N_10420,N_9182,N_9833);
or U10421 (N_10421,N_8722,N_9914);
xor U10422 (N_10422,N_8559,N_9605);
or U10423 (N_10423,N_9842,N_9926);
or U10424 (N_10424,N_8334,N_9556);
nand U10425 (N_10425,N_8815,N_8198);
xor U10426 (N_10426,N_9568,N_8577);
nand U10427 (N_10427,N_8244,N_9777);
nor U10428 (N_10428,N_8348,N_9636);
nand U10429 (N_10429,N_9931,N_8358);
or U10430 (N_10430,N_9289,N_9660);
xor U10431 (N_10431,N_9169,N_8862);
xnor U10432 (N_10432,N_8616,N_8047);
or U10433 (N_10433,N_8493,N_9774);
or U10434 (N_10434,N_9478,N_9128);
nand U10435 (N_10435,N_9126,N_8394);
and U10436 (N_10436,N_9249,N_9093);
and U10437 (N_10437,N_9728,N_8877);
xnor U10438 (N_10438,N_8231,N_9531);
nor U10439 (N_10439,N_8307,N_8757);
and U10440 (N_10440,N_8706,N_8948);
nor U10441 (N_10441,N_9919,N_8952);
and U10442 (N_10442,N_9115,N_8067);
xnor U10443 (N_10443,N_9253,N_8555);
nor U10444 (N_10444,N_8179,N_9075);
nand U10445 (N_10445,N_9203,N_8465);
nand U10446 (N_10446,N_8056,N_9664);
nor U10447 (N_10447,N_9078,N_9494);
and U10448 (N_10448,N_9116,N_8800);
or U10449 (N_10449,N_9425,N_8224);
nor U10450 (N_10450,N_8442,N_8313);
nor U10451 (N_10451,N_9817,N_8535);
nor U10452 (N_10452,N_9889,N_9690);
nor U10453 (N_10453,N_8416,N_9741);
xnor U10454 (N_10454,N_8284,N_9007);
nand U10455 (N_10455,N_9029,N_8407);
xnor U10456 (N_10456,N_9928,N_8401);
nand U10457 (N_10457,N_8285,N_9823);
and U10458 (N_10458,N_8962,N_9418);
xor U10459 (N_10459,N_8336,N_8367);
and U10460 (N_10460,N_9839,N_8668);
and U10461 (N_10461,N_8993,N_8802);
nand U10462 (N_10462,N_8733,N_8640);
nand U10463 (N_10463,N_9381,N_8804);
or U10464 (N_10464,N_9074,N_9459);
or U10465 (N_10465,N_8512,N_9290);
nor U10466 (N_10466,N_9545,N_8311);
xor U10467 (N_10467,N_9019,N_8247);
xnor U10468 (N_10468,N_8700,N_8532);
nor U10469 (N_10469,N_9338,N_8752);
xnor U10470 (N_10470,N_8068,N_9608);
xnor U10471 (N_10471,N_8755,N_8273);
and U10472 (N_10472,N_9592,N_8115);
and U10473 (N_10473,N_9601,N_8472);
and U10474 (N_10474,N_9904,N_8456);
and U10475 (N_10475,N_9097,N_9152);
xnor U10476 (N_10476,N_8908,N_8717);
nand U10477 (N_10477,N_8486,N_8933);
nor U10478 (N_10478,N_8606,N_8105);
and U10479 (N_10479,N_9483,N_9385);
or U10480 (N_10480,N_9520,N_9930);
and U10481 (N_10481,N_9132,N_8977);
or U10482 (N_10482,N_8907,N_8217);
nor U10483 (N_10483,N_8811,N_8987);
nand U10484 (N_10484,N_8780,N_8141);
or U10485 (N_10485,N_8701,N_9693);
and U10486 (N_10486,N_9759,N_8847);
xor U10487 (N_10487,N_9582,N_8463);
or U10488 (N_10488,N_9242,N_9405);
and U10489 (N_10489,N_9676,N_8005);
or U10490 (N_10490,N_8743,N_8321);
or U10491 (N_10491,N_8449,N_9820);
and U10492 (N_10492,N_9775,N_8750);
nand U10493 (N_10493,N_8018,N_9652);
nand U10494 (N_10494,N_9694,N_9802);
and U10495 (N_10495,N_8166,N_8969);
nor U10496 (N_10496,N_9913,N_9127);
and U10497 (N_10497,N_8919,N_8835);
and U10498 (N_10498,N_8628,N_8738);
nor U10499 (N_10499,N_8714,N_8260);
and U10500 (N_10500,N_9606,N_9406);
and U10501 (N_10501,N_9614,N_8513);
xnor U10502 (N_10502,N_9060,N_9895);
and U10503 (N_10503,N_8208,N_8531);
xor U10504 (N_10504,N_9668,N_9905);
nand U10505 (N_10505,N_8797,N_8896);
and U10506 (N_10506,N_8791,N_8006);
nand U10507 (N_10507,N_9602,N_9200);
and U10508 (N_10508,N_8232,N_9899);
nor U10509 (N_10509,N_9306,N_9416);
and U10510 (N_10510,N_9108,N_8092);
and U10511 (N_10511,N_8418,N_8934);
nor U10512 (N_10512,N_8184,N_9630);
xor U10513 (N_10513,N_8698,N_8129);
or U10514 (N_10514,N_9675,N_9410);
xnor U10515 (N_10515,N_9273,N_9735);
xor U10516 (N_10516,N_9350,N_9768);
or U10517 (N_10517,N_8730,N_9340);
or U10518 (N_10518,N_9279,N_8533);
or U10519 (N_10519,N_9096,N_8175);
and U10520 (N_10520,N_9238,N_9558);
or U10521 (N_10521,N_9767,N_8197);
nor U10522 (N_10522,N_8164,N_9603);
xor U10523 (N_10523,N_8020,N_9423);
and U10524 (N_10524,N_9439,N_8967);
or U10525 (N_10525,N_9832,N_8667);
nor U10526 (N_10526,N_8945,N_8707);
and U10527 (N_10527,N_9574,N_8708);
xor U10528 (N_10528,N_9856,N_9303);
nor U10529 (N_10529,N_9335,N_9875);
nor U10530 (N_10530,N_9301,N_9968);
and U10531 (N_10531,N_8946,N_9884);
nor U10532 (N_10532,N_9329,N_9815);
and U10533 (N_10533,N_9048,N_9944);
xor U10534 (N_10534,N_8287,N_9996);
and U10535 (N_10535,N_9607,N_9219);
or U10536 (N_10536,N_8327,N_9743);
nor U10537 (N_10537,N_9463,N_9161);
xor U10538 (N_10538,N_8427,N_8520);
nand U10539 (N_10539,N_9051,N_8839);
xor U10540 (N_10540,N_8557,N_8243);
and U10541 (N_10541,N_8148,N_9831);
xnor U10542 (N_10542,N_8296,N_8744);
or U10543 (N_10543,N_9563,N_9559);
xnor U10544 (N_10544,N_9083,N_8781);
and U10545 (N_10545,N_8391,N_9570);
nor U10546 (N_10546,N_8104,N_8226);
or U10547 (N_10547,N_8271,N_9666);
and U10548 (N_10548,N_9316,N_9877);
xnor U10549 (N_10549,N_8032,N_9154);
and U10550 (N_10550,N_9688,N_8956);
and U10551 (N_10551,N_9619,N_8817);
or U10552 (N_10552,N_8834,N_8090);
nand U10553 (N_10553,N_9631,N_8674);
and U10554 (N_10554,N_8949,N_9297);
or U10555 (N_10555,N_9246,N_8140);
or U10556 (N_10556,N_9639,N_9168);
xor U10557 (N_10557,N_9901,N_8091);
nor U10558 (N_10558,N_8883,N_9482);
or U10559 (N_10559,N_8718,N_8558);
or U10560 (N_10560,N_8439,N_9635);
xor U10561 (N_10561,N_9984,N_8679);
and U10562 (N_10562,N_8288,N_8097);
nor U10563 (N_10563,N_9404,N_8970);
nor U10564 (N_10564,N_8255,N_8739);
nor U10565 (N_10565,N_8190,N_9146);
xor U10566 (N_10566,N_9129,N_8641);
nor U10567 (N_10567,N_8066,N_8789);
xnor U10568 (N_10568,N_8918,N_9015);
and U10569 (N_10569,N_8866,N_9006);
and U10570 (N_10570,N_8204,N_8076);
and U10571 (N_10571,N_8042,N_8702);
and U10572 (N_10572,N_8353,N_8904);
nor U10573 (N_10573,N_9809,N_8983);
or U10574 (N_10574,N_8483,N_8556);
and U10575 (N_10575,N_9120,N_9546);
xor U10576 (N_10576,N_8696,N_8779);
and U10577 (N_10577,N_9104,N_9801);
nand U10578 (N_10578,N_8145,N_9845);
nand U10579 (N_10579,N_8096,N_9213);
or U10580 (N_10580,N_8669,N_8763);
nand U10581 (N_10581,N_8878,N_8903);
and U10582 (N_10582,N_8759,N_8735);
or U10583 (N_10583,N_8686,N_8438);
xor U10584 (N_10584,N_9026,N_8178);
nor U10585 (N_10585,N_9733,N_9009);
xnor U10586 (N_10586,N_9414,N_9650);
nor U10587 (N_10587,N_8238,N_9684);
nor U10588 (N_10588,N_9551,N_8771);
and U10589 (N_10589,N_9646,N_9387);
xor U10590 (N_10590,N_9770,N_8909);
nor U10591 (N_10591,N_8734,N_8732);
and U10592 (N_10592,N_8301,N_9156);
nand U10593 (N_10593,N_8642,N_8214);
nand U10594 (N_10594,N_8149,N_8979);
nor U10595 (N_10595,N_9995,N_9512);
nand U10596 (N_10596,N_9593,N_9739);
and U10597 (N_10597,N_9039,N_8016);
xnor U10598 (N_10598,N_9324,N_9962);
nand U10599 (N_10599,N_8756,N_8482);
and U10600 (N_10600,N_8692,N_9378);
or U10601 (N_10601,N_8856,N_8503);
or U10602 (N_10602,N_8087,N_9971);
nand U10603 (N_10603,N_8395,N_9830);
or U10604 (N_10604,N_8469,N_8363);
nand U10605 (N_10605,N_9088,N_8954);
nand U10606 (N_10606,N_9989,N_8222);
xor U10607 (N_10607,N_8646,N_9227);
nor U10608 (N_10608,N_9067,N_8516);
nand U10609 (N_10609,N_8130,N_9640);
and U10610 (N_10610,N_9233,N_8710);
xnor U10611 (N_10611,N_8415,N_8474);
and U10612 (N_10612,N_9935,N_9081);
nor U10613 (N_10613,N_9723,N_8305);
xnor U10614 (N_10614,N_8944,N_8766);
and U10615 (N_10615,N_9399,N_9443);
or U10616 (N_10616,N_9990,N_8262);
or U10617 (N_10617,N_9347,N_8033);
nor U10618 (N_10618,N_8404,N_9808);
xnor U10619 (N_10619,N_9403,N_8673);
and U10620 (N_10620,N_9579,N_9348);
nand U10621 (N_10621,N_9369,N_9305);
or U10622 (N_10622,N_9501,N_9254);
or U10623 (N_10623,N_9267,N_8689);
nand U10624 (N_10624,N_9259,N_8985);
or U10625 (N_10625,N_9234,N_8951);
xnor U10626 (N_10626,N_9449,N_8189);
or U10627 (N_10627,N_8282,N_8526);
and U10628 (N_10628,N_9442,N_8796);
xnor U10629 (N_10629,N_8988,N_9957);
xor U10630 (N_10630,N_8798,N_8932);
and U10631 (N_10631,N_9942,N_8303);
or U10632 (N_10632,N_9885,N_8711);
nand U10633 (N_10633,N_9760,N_8000);
xor U10634 (N_10634,N_9966,N_9744);
or U10635 (N_10635,N_9411,N_8113);
nor U10636 (N_10636,N_9980,N_9402);
nor U10637 (N_10637,N_9647,N_9562);
nand U10638 (N_10638,N_8595,N_9140);
or U10639 (N_10639,N_9313,N_9586);
nor U10640 (N_10640,N_9569,N_9903);
nand U10641 (N_10641,N_9618,N_8302);
nand U10642 (N_10642,N_9135,N_9422);
and U10643 (N_10643,N_9170,N_9505);
nand U10644 (N_10644,N_9793,N_8436);
nor U10645 (N_10645,N_8542,N_9557);
and U10646 (N_10646,N_8504,N_9145);
or U10647 (N_10647,N_8013,N_8242);
xor U10648 (N_10648,N_9644,N_9292);
nand U10649 (N_10649,N_8554,N_8107);
xnor U10650 (N_10650,N_9438,N_8842);
xnor U10651 (N_10651,N_9997,N_8078);
nor U10652 (N_10652,N_8432,N_9245);
and U10653 (N_10653,N_9967,N_9709);
nor U10654 (N_10654,N_8991,N_8524);
and U10655 (N_10655,N_9524,N_9841);
and U10656 (N_10656,N_8894,N_8561);
nand U10657 (N_10657,N_8429,N_8863);
xor U10658 (N_10658,N_8843,N_9909);
nor U10659 (N_10659,N_8207,N_9322);
and U10660 (N_10660,N_9491,N_8916);
xnor U10661 (N_10661,N_9632,N_8019);
or U10662 (N_10662,N_8203,N_9333);
or U10663 (N_10663,N_8720,N_8760);
or U10664 (N_10664,N_8540,N_9496);
xnor U10665 (N_10665,N_8343,N_8841);
nor U10666 (N_10666,N_9495,N_8206);
xnor U10667 (N_10667,N_9485,N_9190);
nand U10668 (N_10668,N_9184,N_9506);
nor U10669 (N_10669,N_8943,N_9871);
nand U10670 (N_10670,N_8662,N_9860);
or U10671 (N_10671,N_8462,N_9409);
or U10672 (N_10672,N_8589,N_8613);
xnor U10673 (N_10673,N_8344,N_8376);
and U10674 (N_10674,N_8030,N_8241);
nand U10675 (N_10675,N_8807,N_8249);
nor U10676 (N_10676,N_8620,N_9307);
or U10677 (N_10677,N_8740,N_8981);
nand U10678 (N_10678,N_8855,N_9457);
and U10679 (N_10679,N_8392,N_8377);
or U10680 (N_10680,N_9799,N_8541);
xnor U10681 (N_10681,N_8035,N_8182);
nand U10682 (N_10682,N_9974,N_8509);
and U10683 (N_10683,N_9084,N_8623);
or U10684 (N_10684,N_8044,N_8125);
or U10685 (N_10685,N_8414,N_9532);
xor U10686 (N_10686,N_8098,N_8040);
and U10687 (N_10687,N_9625,N_9695);
xor U10688 (N_10688,N_9916,N_8111);
or U10689 (N_10689,N_9627,N_9502);
nor U10690 (N_10690,N_8665,N_8527);
xor U10691 (N_10691,N_8729,N_8139);
nor U10692 (N_10692,N_8117,N_9681);
and U10693 (N_10693,N_9669,N_9309);
and U10694 (N_10694,N_8082,N_8457);
nand U10695 (N_10695,N_8651,N_8254);
and U10696 (N_10696,N_8723,N_8072);
nor U10697 (N_10697,N_9493,N_9736);
nand U10698 (N_10698,N_8036,N_8699);
nor U10699 (N_10699,N_8737,N_9197);
or U10700 (N_10700,N_8194,N_9621);
xnor U10701 (N_10701,N_8938,N_8724);
and U10702 (N_10702,N_8476,N_9139);
xor U10703 (N_10703,N_8366,N_9477);
and U10704 (N_10704,N_9275,N_8031);
nor U10705 (N_10705,N_9068,N_9271);
nor U10706 (N_10706,N_9902,N_8408);
and U10707 (N_10707,N_9446,N_9806);
nand U10708 (N_10708,N_8186,N_8552);
or U10709 (N_10709,N_8849,N_8295);
xnor U10710 (N_10710,N_8695,N_9082);
or U10711 (N_10711,N_8445,N_8652);
and U10712 (N_10712,N_8216,N_8422);
nand U10713 (N_10713,N_8286,N_8890);
nor U10714 (N_10714,N_8660,N_9452);
or U10715 (N_10715,N_9435,N_8041);
xnor U10716 (N_10716,N_9353,N_9589);
nor U10717 (N_10717,N_8371,N_8892);
nand U10718 (N_10718,N_8782,N_9231);
or U10719 (N_10719,N_8021,N_9167);
or U10720 (N_10720,N_8046,N_8338);
nand U10721 (N_10721,N_9792,N_8237);
or U10722 (N_10722,N_9368,N_8931);
or U10723 (N_10723,N_8498,N_9395);
xor U10724 (N_10724,N_9810,N_9450);
and U10725 (N_10725,N_8518,N_9005);
and U10726 (N_10726,N_9417,N_9731);
nor U10727 (N_10727,N_9252,N_8950);
and U10728 (N_10728,N_8507,N_8258);
and U10729 (N_10729,N_9829,N_8957);
nor U10730 (N_10730,N_8649,N_8248);
xnor U10731 (N_10731,N_9887,N_8132);
nand U10732 (N_10732,N_8631,N_9049);
or U10733 (N_10733,N_8523,N_8844);
nor U10734 (N_10734,N_9925,N_9536);
nor U10735 (N_10735,N_9891,N_9798);
or U10736 (N_10736,N_9159,N_9713);
and U10737 (N_10737,N_9337,N_9367);
and U10738 (N_10738,N_9740,N_9598);
xnor U10739 (N_10739,N_8073,N_8901);
nand U10740 (N_10740,N_9202,N_8409);
nor U10741 (N_10741,N_9703,N_8034);
nand U10742 (N_10742,N_8084,N_8715);
or U10743 (N_10743,N_8309,N_9431);
and U10744 (N_10744,N_9752,N_9499);
and U10745 (N_10745,N_8691,N_8264);
xnor U10746 (N_10746,N_9811,N_9018);
or U10747 (N_10747,N_8592,N_8929);
nor U10748 (N_10748,N_9470,N_9163);
and U10749 (N_10749,N_8101,N_9336);
nor U10750 (N_10750,N_8982,N_8417);
nor U10751 (N_10751,N_8935,N_9221);
nor U10752 (N_10752,N_9595,N_9776);
and U10753 (N_10753,N_9393,N_8428);
or U10754 (N_10754,N_9578,N_8122);
nand U10755 (N_10755,N_8971,N_9782);
xor U10756 (N_10756,N_9611,N_9527);
xor U10757 (N_10757,N_8806,N_8937);
nor U10758 (N_10758,N_8171,N_8831);
nand U10759 (N_10759,N_8126,N_8580);
or U10760 (N_10760,N_8211,N_8871);
xnor U10761 (N_10761,N_9363,N_9617);
or U10762 (N_10762,N_8389,N_9795);
or U10763 (N_10763,N_9560,N_9261);
and U10764 (N_10764,N_8173,N_9826);
nor U10765 (N_10765,N_8425,N_8370);
or U10766 (N_10766,N_9122,N_8549);
nand U10767 (N_10767,N_8180,N_8339);
xor U10768 (N_10768,N_9042,N_9523);
xnor U10769 (N_10769,N_8277,N_9991);
nor U10770 (N_10770,N_9063,N_8341);
or U10771 (N_10771,N_8964,N_9879);
xor U10772 (N_10772,N_9356,N_9397);
nor U10773 (N_10773,N_8632,N_8905);
and U10774 (N_10774,N_9755,N_9716);
nand U10775 (N_10775,N_9244,N_9732);
nor U10776 (N_10776,N_8624,N_9641);
nand U10777 (N_10777,N_9698,N_9766);
nor U10778 (N_10778,N_9142,N_8941);
and U10779 (N_10779,N_8658,N_9686);
and U10780 (N_10780,N_9288,N_8603);
nor U10781 (N_10781,N_8123,N_9100);
xor U10782 (N_10782,N_8861,N_8276);
nand U10783 (N_10783,N_9691,N_8959);
nor U10784 (N_10784,N_8645,N_9025);
xor U10785 (N_10785,N_9835,N_9294);
and U10786 (N_10786,N_9251,N_9979);
xor U10787 (N_10787,N_9066,N_9769);
xnor U10788 (N_10788,N_8174,N_9521);
nand U10789 (N_10789,N_9814,N_9360);
nor U10790 (N_10790,N_8135,N_8289);
and U10791 (N_10791,N_8608,N_8870);
nand U10792 (N_10792,N_8822,N_9490);
and U10793 (N_10793,N_9543,N_8657);
and U10794 (N_10794,N_9143,N_8891);
or U10795 (N_10795,N_9304,N_8185);
nor U10796 (N_10796,N_9222,N_9220);
nand U10797 (N_10797,N_8810,N_9689);
and U10798 (N_10798,N_9825,N_8769);
xnor U10799 (N_10799,N_9265,N_8261);
nor U10800 (N_10800,N_9280,N_9629);
and U10801 (N_10801,N_9031,N_9697);
xor U10802 (N_10802,N_9327,N_9661);
nor U10803 (N_10803,N_9434,N_9591);
nor U10804 (N_10804,N_9153,N_9160);
nor U10805 (N_10805,N_9243,N_9670);
or U10806 (N_10806,N_8081,N_9453);
nor U10807 (N_10807,N_9437,N_8362);
xnor U10808 (N_10808,N_8694,N_9016);
nor U10809 (N_10809,N_8879,N_8986);
xnor U10810 (N_10810,N_9946,N_9432);
nor U10811 (N_10811,N_9187,N_9863);
or U10812 (N_10812,N_8147,N_8611);
xor U10813 (N_10813,N_9373,N_8413);
or U10814 (N_10814,N_9500,N_8426);
nor U10815 (N_10815,N_9003,N_9734);
nand U10816 (N_10816,N_9960,N_8647);
nand U10817 (N_10817,N_9293,N_8480);
xor U10818 (N_10818,N_8650,N_9988);
or U10819 (N_10819,N_9837,N_9824);
xnor U10820 (N_10820,N_8659,N_9612);
or U10821 (N_10821,N_8911,N_9714);
or U10822 (N_10822,N_8496,N_8488);
and U10823 (N_10823,N_8602,N_9103);
and U10824 (N_10824,N_8578,N_8063);
xnor U10825 (N_10825,N_8223,N_9451);
or U10826 (N_10826,N_8515,N_9228);
nor U10827 (N_10827,N_9981,N_9746);
nand U10828 (N_10828,N_8644,N_8357);
nor U10829 (N_10829,N_8768,N_9428);
nand U10830 (N_10830,N_9970,N_8163);
xor U10831 (N_10831,N_8551,N_8049);
nand U10832 (N_10832,N_8002,N_9737);
nor U10833 (N_10833,N_8025,N_9964);
and U10834 (N_10834,N_8440,N_8143);
or U10835 (N_10835,N_9465,N_9836);
nand U10836 (N_10836,N_8310,N_8329);
nor U10837 (N_10837,N_9445,N_8388);
nand U10838 (N_10838,N_9986,N_8331);
nor U10839 (N_10839,N_9936,N_9017);
nand U10840 (N_10840,N_9961,N_8958);
xor U10841 (N_10841,N_8003,N_9344);
xor U10842 (N_10842,N_9383,N_9788);
or U10843 (N_10843,N_8402,N_9471);
and U10844 (N_10844,N_8443,N_9057);
xnor U10845 (N_10845,N_8776,N_8579);
xnor U10846 (N_10846,N_9537,N_9881);
nor U10847 (N_10847,N_9717,N_8239);
nand U10848 (N_10848,N_9912,N_8365);
nand U10849 (N_10849,N_9638,N_9319);
nor U10850 (N_10850,N_9937,N_9533);
and U10851 (N_10851,N_8293,N_9302);
or U10852 (N_10852,N_9426,N_8342);
and U10853 (N_10853,N_9800,N_8057);
or U10854 (N_10854,N_9932,N_9604);
or U10855 (N_10855,N_9699,N_8250);
xor U10856 (N_10856,N_9657,N_8569);
nor U10857 (N_10857,N_8278,N_9761);
xnor U10858 (N_10858,N_9384,N_9549);
or U10859 (N_10859,N_8913,N_9372);
and U10860 (N_10860,N_9038,N_9859);
nand U10861 (N_10861,N_8795,N_8029);
and U10862 (N_10862,N_8477,N_8118);
or U10863 (N_10863,N_9615,N_9476);
and U10864 (N_10864,N_9923,N_9702);
nor U10865 (N_10865,N_9854,N_8364);
and U10866 (N_10866,N_8976,N_8155);
or U10867 (N_10867,N_8887,N_9656);
xor U10868 (N_10868,N_8629,N_8838);
nand U10869 (N_10869,N_8345,N_8636);
nor U10870 (N_10870,N_8980,N_8138);
nor U10871 (N_10871,N_8746,N_9730);
xnor U10872 (N_10872,N_8626,N_9710);
and U10873 (N_10873,N_8379,N_9043);
and U10874 (N_10874,N_8544,N_8088);
nor U10875 (N_10875,N_8590,N_8820);
nor U10876 (N_10876,N_9394,N_8441);
or U10877 (N_10877,N_8998,N_9948);
nand U10878 (N_10878,N_9090,N_8814);
nor U10879 (N_10879,N_9865,N_9659);
xor U10880 (N_10880,N_8491,N_9771);
nand U10881 (N_10881,N_9441,N_8419);
and U10882 (N_10882,N_9046,N_8663);
nor U10883 (N_10883,N_8080,N_8473);
or U10884 (N_10884,N_9828,N_8259);
nor U10885 (N_10885,N_9529,N_9298);
and U10886 (N_10886,N_8257,N_9511);
xnor U10887 (N_10887,N_9201,N_9610);
or U10888 (N_10888,N_9033,N_8378);
nand U10889 (N_10889,N_9193,N_9590);
nand U10890 (N_10890,N_9225,N_9374);
or U10891 (N_10891,N_9785,N_9951);
nor U10892 (N_10892,N_9260,N_9468);
and U10893 (N_10893,N_9268,N_9973);
or U10894 (N_10894,N_9270,N_9427);
or U10895 (N_10895,N_9052,N_8390);
xor U10896 (N_10896,N_9112,N_8514);
nor U10897 (N_10897,N_9044,N_8785);
nor U10898 (N_10898,N_8537,N_9628);
or U10899 (N_10899,N_8406,N_9894);
or U10900 (N_10900,N_9719,N_8074);
and U10901 (N_10901,N_8437,N_9256);
or U10902 (N_10902,N_8468,N_8942);
xnor U10903 (N_10903,N_9872,N_8786);
xnor U10904 (N_10904,N_8299,N_9910);
nand U10905 (N_10905,N_9838,N_8550);
nor U10906 (N_10906,N_9248,N_9870);
or U10907 (N_10907,N_9375,N_8853);
nand U10908 (N_10908,N_9359,N_9498);
nor U10909 (N_10909,N_8924,N_9812);
or U10910 (N_10910,N_8220,N_8670);
xnor U10911 (N_10911,N_9094,N_8430);
nor U10912 (N_10912,N_9655,N_9408);
nand U10913 (N_10913,N_9773,N_9474);
and U10914 (N_10914,N_9262,N_9206);
and U10915 (N_10915,N_9264,N_8574);
nand U10916 (N_10916,N_8024,N_9021);
or U10917 (N_10917,N_9762,N_8819);
xnor U10918 (N_10918,N_8587,N_8992);
nand U10919 (N_10919,N_8228,N_8840);
or U10920 (N_10920,N_8547,N_9318);
nor U10921 (N_10921,N_9050,N_9357);
or U10922 (N_10922,N_8794,N_9472);
and U10923 (N_10923,N_8015,N_8079);
or U10924 (N_10924,N_9300,N_9099);
and U10925 (N_10925,N_9237,N_8837);
or U10926 (N_10926,N_9354,N_8492);
or U10927 (N_10927,N_8386,N_9599);
nand U10928 (N_10928,N_8200,N_8726);
and U10929 (N_10929,N_9906,N_8447);
nor U10930 (N_10930,N_8109,N_9765);
nor U10931 (N_10931,N_9370,N_9917);
nor U10932 (N_10932,N_8828,N_9507);
or U10933 (N_10933,N_8412,N_8654);
or U10934 (N_10934,N_9071,N_8889);
xor U10935 (N_10935,N_8252,N_8902);
or U10936 (N_10936,N_9939,N_9352);
and U10937 (N_10937,N_9086,N_8158);
nor U10938 (N_10938,N_9239,N_8308);
nor U10939 (N_10939,N_9518,N_8571);
nor U10940 (N_10940,N_9070,N_8570);
nor U10941 (N_10941,N_8974,N_9987);
nand U10942 (N_10942,N_8452,N_8368);
nor U10943 (N_10943,N_9147,N_8793);
and U10944 (N_10944,N_9959,N_9542);
nand U10945 (N_10945,N_8150,N_9729);
nor U10946 (N_10946,N_8326,N_8361);
or U10947 (N_10947,N_9023,N_9117);
or U10948 (N_10948,N_9849,N_8320);
nand U10949 (N_10949,N_8639,N_9706);
or U10950 (N_10950,N_8460,N_8917);
nor U10951 (N_10951,N_8596,N_9888);
xnor U10952 (N_10952,N_9857,N_9922);
nand U10953 (N_10953,N_8625,N_8522);
or U10954 (N_10954,N_9480,N_8268);
nor U10955 (N_10955,N_9553,N_8100);
nand U10956 (N_10956,N_8256,N_9898);
and U10957 (N_10957,N_9089,N_8191);
and U10958 (N_10958,N_9976,N_9321);
and U10959 (N_10959,N_9654,N_9258);
nand U10960 (N_10960,N_8102,N_8168);
and U10961 (N_10961,N_8627,N_8963);
xnor U10962 (N_10962,N_8767,N_9947);
or U10963 (N_10963,N_9027,N_8470);
xor U10964 (N_10964,N_9282,N_8398);
or U10965 (N_10965,N_9178,N_9185);
nand U10966 (N_10966,N_8253,N_9458);
or U10967 (N_10967,N_8888,N_9750);
nand U10968 (N_10968,N_8661,N_8317);
or U10969 (N_10969,N_8801,N_8332);
xnor U10970 (N_10970,N_9119,N_9034);
xnor U10971 (N_10971,N_8788,N_8027);
nor U10972 (N_10972,N_9596,N_9682);
and U10973 (N_10973,N_8335,N_8380);
or U10974 (N_10974,N_9526,N_9199);
nor U10975 (N_10975,N_9020,N_9004);
nand U10976 (N_10976,N_9943,N_8459);
nor U10977 (N_10977,N_9400,N_9430);
nand U10978 (N_10978,N_9250,N_9102);
or U10979 (N_10979,N_9977,N_9751);
nand U10980 (N_10980,N_9918,N_9299);
or U10981 (N_10981,N_9362,N_9095);
and U10982 (N_10982,N_8170,N_9998);
nor U10983 (N_10983,N_8375,N_8246);
or U10984 (N_10984,N_8713,N_8007);
xor U10985 (N_10985,N_8183,N_9600);
xnor U10986 (N_10986,N_8274,N_8106);
nor U10987 (N_10987,N_8275,N_8095);
xor U10988 (N_10988,N_9594,N_9107);
nor U10989 (N_10989,N_8564,N_8114);
or U10990 (N_10990,N_9196,N_9240);
nand U10991 (N_10991,N_8385,N_8280);
nor U10992 (N_10992,N_9205,N_8023);
nand U10993 (N_10993,N_9284,N_8369);
nand U10994 (N_10994,N_9623,N_9651);
nand U10995 (N_10995,N_8874,N_8328);
or U10996 (N_10996,N_8893,N_9992);
nand U10997 (N_10997,N_8294,N_8736);
nor U10998 (N_10998,N_9079,N_8860);
nor U10999 (N_10999,N_8052,N_8464);
and U11000 (N_11000,N_8896,N_8530);
nand U11001 (N_11001,N_9025,N_9414);
and U11002 (N_11002,N_8227,N_9297);
xnor U11003 (N_11003,N_9774,N_8756);
xnor U11004 (N_11004,N_8619,N_8252);
nand U11005 (N_11005,N_8906,N_8489);
nand U11006 (N_11006,N_8270,N_8526);
and U11007 (N_11007,N_8856,N_8611);
or U11008 (N_11008,N_8889,N_8385);
nand U11009 (N_11009,N_9787,N_9969);
xnor U11010 (N_11010,N_9007,N_9411);
and U11011 (N_11011,N_9172,N_9477);
nor U11012 (N_11012,N_9406,N_8940);
or U11013 (N_11013,N_8601,N_8317);
or U11014 (N_11014,N_8613,N_9160);
nor U11015 (N_11015,N_8750,N_9487);
nor U11016 (N_11016,N_9710,N_8473);
nand U11017 (N_11017,N_9520,N_8469);
and U11018 (N_11018,N_9327,N_9057);
and U11019 (N_11019,N_9209,N_8072);
nand U11020 (N_11020,N_9904,N_9542);
nor U11021 (N_11021,N_8706,N_8148);
or U11022 (N_11022,N_9532,N_9892);
nor U11023 (N_11023,N_8319,N_9369);
and U11024 (N_11024,N_9496,N_8715);
nand U11025 (N_11025,N_9764,N_8025);
and U11026 (N_11026,N_8068,N_8730);
and U11027 (N_11027,N_8028,N_8569);
xor U11028 (N_11028,N_8409,N_8888);
and U11029 (N_11029,N_8610,N_9569);
nand U11030 (N_11030,N_8860,N_8208);
xor U11031 (N_11031,N_9956,N_8355);
or U11032 (N_11032,N_9915,N_9271);
nand U11033 (N_11033,N_8538,N_9202);
and U11034 (N_11034,N_9648,N_9170);
or U11035 (N_11035,N_9122,N_9973);
and U11036 (N_11036,N_8596,N_9536);
nand U11037 (N_11037,N_8532,N_8604);
or U11038 (N_11038,N_9098,N_8380);
and U11039 (N_11039,N_8822,N_9034);
or U11040 (N_11040,N_9380,N_8627);
xor U11041 (N_11041,N_9555,N_8019);
nand U11042 (N_11042,N_9279,N_9144);
nor U11043 (N_11043,N_8854,N_9720);
and U11044 (N_11044,N_8301,N_9654);
or U11045 (N_11045,N_9532,N_8745);
xnor U11046 (N_11046,N_9383,N_8306);
and U11047 (N_11047,N_9526,N_9952);
and U11048 (N_11048,N_8172,N_9037);
xnor U11049 (N_11049,N_8368,N_8838);
nor U11050 (N_11050,N_9610,N_8811);
or U11051 (N_11051,N_9272,N_9164);
nand U11052 (N_11052,N_8710,N_9047);
xor U11053 (N_11053,N_9384,N_8727);
or U11054 (N_11054,N_9008,N_8015);
or U11055 (N_11055,N_8734,N_9305);
or U11056 (N_11056,N_9782,N_8966);
xor U11057 (N_11057,N_8050,N_9865);
nand U11058 (N_11058,N_9865,N_9721);
and U11059 (N_11059,N_9930,N_8323);
xnor U11060 (N_11060,N_9166,N_8930);
nor U11061 (N_11061,N_9310,N_9128);
nor U11062 (N_11062,N_8218,N_8778);
nor U11063 (N_11063,N_9808,N_9458);
and U11064 (N_11064,N_9749,N_9443);
xnor U11065 (N_11065,N_8039,N_8096);
nor U11066 (N_11066,N_8842,N_8095);
and U11067 (N_11067,N_8519,N_8573);
nor U11068 (N_11068,N_8670,N_8693);
or U11069 (N_11069,N_8844,N_9534);
and U11070 (N_11070,N_8639,N_8694);
and U11071 (N_11071,N_9785,N_8890);
and U11072 (N_11072,N_9433,N_8299);
nor U11073 (N_11073,N_8164,N_9903);
nor U11074 (N_11074,N_9202,N_8946);
nor U11075 (N_11075,N_8744,N_9430);
and U11076 (N_11076,N_9990,N_9619);
nand U11077 (N_11077,N_8362,N_8905);
xor U11078 (N_11078,N_8754,N_8362);
and U11079 (N_11079,N_8330,N_9876);
or U11080 (N_11080,N_8217,N_9629);
nor U11081 (N_11081,N_8739,N_9265);
nor U11082 (N_11082,N_8849,N_8123);
or U11083 (N_11083,N_9851,N_9301);
nand U11084 (N_11084,N_9510,N_9069);
xnor U11085 (N_11085,N_8249,N_9337);
nand U11086 (N_11086,N_9876,N_9412);
xor U11087 (N_11087,N_8960,N_8277);
xor U11088 (N_11088,N_8388,N_9489);
xnor U11089 (N_11089,N_9522,N_8996);
xnor U11090 (N_11090,N_9936,N_8482);
xor U11091 (N_11091,N_9938,N_9362);
or U11092 (N_11092,N_9992,N_9751);
and U11093 (N_11093,N_9572,N_8249);
nand U11094 (N_11094,N_8979,N_9741);
and U11095 (N_11095,N_9014,N_9917);
and U11096 (N_11096,N_8046,N_9140);
or U11097 (N_11097,N_8189,N_9158);
and U11098 (N_11098,N_9367,N_8871);
nor U11099 (N_11099,N_8599,N_9017);
nor U11100 (N_11100,N_9432,N_9152);
xnor U11101 (N_11101,N_9609,N_9348);
nand U11102 (N_11102,N_9013,N_8498);
and U11103 (N_11103,N_9002,N_9195);
nand U11104 (N_11104,N_9015,N_9933);
xor U11105 (N_11105,N_8907,N_9983);
or U11106 (N_11106,N_9197,N_9045);
or U11107 (N_11107,N_9562,N_9710);
and U11108 (N_11108,N_9636,N_8731);
or U11109 (N_11109,N_9037,N_9220);
and U11110 (N_11110,N_8201,N_8077);
xor U11111 (N_11111,N_8699,N_8731);
and U11112 (N_11112,N_9652,N_8712);
nor U11113 (N_11113,N_9521,N_9990);
nand U11114 (N_11114,N_9265,N_8197);
and U11115 (N_11115,N_9658,N_8195);
and U11116 (N_11116,N_8935,N_8800);
or U11117 (N_11117,N_9238,N_8314);
nand U11118 (N_11118,N_8041,N_9397);
nand U11119 (N_11119,N_8414,N_9876);
or U11120 (N_11120,N_9041,N_8915);
or U11121 (N_11121,N_8243,N_8854);
nand U11122 (N_11122,N_8094,N_9624);
xnor U11123 (N_11123,N_9256,N_8012);
and U11124 (N_11124,N_9055,N_8872);
and U11125 (N_11125,N_8483,N_9259);
and U11126 (N_11126,N_9351,N_9111);
and U11127 (N_11127,N_8897,N_8740);
nand U11128 (N_11128,N_9259,N_8197);
and U11129 (N_11129,N_9595,N_8821);
nand U11130 (N_11130,N_8945,N_9095);
nand U11131 (N_11131,N_9170,N_8929);
nand U11132 (N_11132,N_9234,N_8989);
xnor U11133 (N_11133,N_8865,N_8018);
and U11134 (N_11134,N_8902,N_9414);
nand U11135 (N_11135,N_9645,N_9361);
or U11136 (N_11136,N_8211,N_8455);
and U11137 (N_11137,N_9891,N_8028);
xor U11138 (N_11138,N_9973,N_9316);
xor U11139 (N_11139,N_8689,N_9634);
nand U11140 (N_11140,N_8213,N_9580);
or U11141 (N_11141,N_8908,N_8863);
xor U11142 (N_11142,N_8414,N_8245);
xor U11143 (N_11143,N_9308,N_9831);
or U11144 (N_11144,N_9777,N_8008);
nor U11145 (N_11145,N_8306,N_8602);
and U11146 (N_11146,N_8323,N_8619);
xor U11147 (N_11147,N_9360,N_9670);
xor U11148 (N_11148,N_9187,N_8835);
or U11149 (N_11149,N_9253,N_8453);
xnor U11150 (N_11150,N_9409,N_9940);
or U11151 (N_11151,N_8376,N_9735);
nand U11152 (N_11152,N_8786,N_9451);
or U11153 (N_11153,N_9409,N_9095);
or U11154 (N_11154,N_9896,N_8566);
xnor U11155 (N_11155,N_9817,N_9769);
and U11156 (N_11156,N_8144,N_9888);
nand U11157 (N_11157,N_8276,N_8990);
and U11158 (N_11158,N_8032,N_8427);
nor U11159 (N_11159,N_8108,N_8637);
xor U11160 (N_11160,N_9331,N_8071);
nor U11161 (N_11161,N_9798,N_8743);
nor U11162 (N_11162,N_8507,N_8859);
and U11163 (N_11163,N_8878,N_9734);
nand U11164 (N_11164,N_9391,N_9150);
xor U11165 (N_11165,N_8880,N_9710);
xnor U11166 (N_11166,N_8702,N_8599);
or U11167 (N_11167,N_9918,N_9181);
nand U11168 (N_11168,N_9653,N_9600);
nand U11169 (N_11169,N_9858,N_8864);
nand U11170 (N_11170,N_8947,N_9051);
and U11171 (N_11171,N_8480,N_9775);
nor U11172 (N_11172,N_9631,N_9134);
and U11173 (N_11173,N_8196,N_8018);
and U11174 (N_11174,N_9685,N_9221);
nor U11175 (N_11175,N_9479,N_8683);
xor U11176 (N_11176,N_9885,N_8309);
nor U11177 (N_11177,N_8467,N_9349);
and U11178 (N_11178,N_9754,N_8813);
nor U11179 (N_11179,N_8518,N_9032);
or U11180 (N_11180,N_8845,N_8571);
nand U11181 (N_11181,N_8038,N_8371);
or U11182 (N_11182,N_9310,N_8808);
nor U11183 (N_11183,N_9619,N_9520);
nor U11184 (N_11184,N_9626,N_9854);
and U11185 (N_11185,N_8498,N_9652);
and U11186 (N_11186,N_8449,N_9784);
nor U11187 (N_11187,N_9835,N_9067);
or U11188 (N_11188,N_8770,N_8999);
nand U11189 (N_11189,N_8335,N_9545);
or U11190 (N_11190,N_9438,N_8185);
or U11191 (N_11191,N_9779,N_8231);
xor U11192 (N_11192,N_9597,N_8598);
nand U11193 (N_11193,N_9130,N_8538);
xor U11194 (N_11194,N_8443,N_9890);
nand U11195 (N_11195,N_9142,N_8105);
and U11196 (N_11196,N_8094,N_9891);
nor U11197 (N_11197,N_9672,N_8743);
or U11198 (N_11198,N_9349,N_8920);
or U11199 (N_11199,N_8800,N_9702);
nor U11200 (N_11200,N_8944,N_9556);
or U11201 (N_11201,N_8755,N_8694);
xnor U11202 (N_11202,N_9229,N_8009);
xor U11203 (N_11203,N_9513,N_9697);
nand U11204 (N_11204,N_9620,N_8159);
nor U11205 (N_11205,N_9507,N_9853);
and U11206 (N_11206,N_8637,N_9708);
nor U11207 (N_11207,N_9616,N_9400);
and U11208 (N_11208,N_9797,N_8282);
xor U11209 (N_11209,N_9933,N_8796);
or U11210 (N_11210,N_9906,N_9593);
or U11211 (N_11211,N_9965,N_8290);
nand U11212 (N_11212,N_9068,N_8963);
xnor U11213 (N_11213,N_9508,N_8558);
or U11214 (N_11214,N_9136,N_8080);
nor U11215 (N_11215,N_8555,N_8392);
or U11216 (N_11216,N_9786,N_9543);
nor U11217 (N_11217,N_8734,N_9435);
nor U11218 (N_11218,N_8487,N_9179);
nor U11219 (N_11219,N_9891,N_8337);
nor U11220 (N_11220,N_8996,N_8775);
nor U11221 (N_11221,N_9561,N_8172);
nor U11222 (N_11222,N_8319,N_8361);
and U11223 (N_11223,N_9865,N_9561);
xnor U11224 (N_11224,N_8595,N_9731);
xnor U11225 (N_11225,N_9121,N_9928);
xor U11226 (N_11226,N_8666,N_8267);
xor U11227 (N_11227,N_8219,N_8532);
nor U11228 (N_11228,N_8406,N_8955);
xor U11229 (N_11229,N_9332,N_8490);
and U11230 (N_11230,N_8658,N_9784);
nor U11231 (N_11231,N_9149,N_9392);
or U11232 (N_11232,N_9819,N_9492);
nand U11233 (N_11233,N_9731,N_9160);
or U11234 (N_11234,N_9808,N_8442);
and U11235 (N_11235,N_9173,N_8431);
or U11236 (N_11236,N_9136,N_9591);
nor U11237 (N_11237,N_9833,N_9643);
and U11238 (N_11238,N_9839,N_9593);
nor U11239 (N_11239,N_8009,N_9314);
nor U11240 (N_11240,N_9604,N_8045);
nor U11241 (N_11241,N_8671,N_9849);
nor U11242 (N_11242,N_8604,N_9968);
xnor U11243 (N_11243,N_9042,N_8987);
nor U11244 (N_11244,N_8915,N_8219);
nor U11245 (N_11245,N_9710,N_8575);
or U11246 (N_11246,N_8389,N_9090);
nand U11247 (N_11247,N_8523,N_8554);
nor U11248 (N_11248,N_8687,N_9426);
nor U11249 (N_11249,N_8411,N_8817);
or U11250 (N_11250,N_8929,N_9477);
nor U11251 (N_11251,N_8121,N_9547);
or U11252 (N_11252,N_8212,N_8648);
or U11253 (N_11253,N_8436,N_9686);
nor U11254 (N_11254,N_8190,N_9152);
nor U11255 (N_11255,N_8217,N_8656);
xnor U11256 (N_11256,N_9623,N_9010);
and U11257 (N_11257,N_8732,N_8041);
xor U11258 (N_11258,N_9839,N_9831);
nor U11259 (N_11259,N_9765,N_8355);
or U11260 (N_11260,N_9969,N_9629);
and U11261 (N_11261,N_8538,N_9617);
nand U11262 (N_11262,N_8048,N_8832);
nor U11263 (N_11263,N_9194,N_9322);
nor U11264 (N_11264,N_9056,N_8766);
xnor U11265 (N_11265,N_9386,N_8249);
and U11266 (N_11266,N_8805,N_8507);
and U11267 (N_11267,N_9790,N_9818);
nand U11268 (N_11268,N_8602,N_9793);
nor U11269 (N_11269,N_8188,N_9963);
nor U11270 (N_11270,N_9819,N_9031);
or U11271 (N_11271,N_9891,N_9633);
and U11272 (N_11272,N_9958,N_8621);
xor U11273 (N_11273,N_9972,N_9704);
nor U11274 (N_11274,N_8050,N_9702);
and U11275 (N_11275,N_8884,N_9606);
xnor U11276 (N_11276,N_9765,N_8435);
nand U11277 (N_11277,N_8060,N_8702);
xor U11278 (N_11278,N_8773,N_9693);
or U11279 (N_11279,N_9219,N_8833);
nand U11280 (N_11280,N_8033,N_8138);
nand U11281 (N_11281,N_8227,N_9910);
xor U11282 (N_11282,N_8393,N_9353);
nor U11283 (N_11283,N_9103,N_8771);
nand U11284 (N_11284,N_8124,N_8873);
and U11285 (N_11285,N_9519,N_9263);
nor U11286 (N_11286,N_9651,N_8236);
and U11287 (N_11287,N_8225,N_8369);
xnor U11288 (N_11288,N_9765,N_9267);
nor U11289 (N_11289,N_8972,N_9016);
and U11290 (N_11290,N_9094,N_8883);
and U11291 (N_11291,N_9370,N_8313);
xor U11292 (N_11292,N_9739,N_8663);
nand U11293 (N_11293,N_9168,N_9003);
and U11294 (N_11294,N_8295,N_8911);
nor U11295 (N_11295,N_9142,N_9912);
nor U11296 (N_11296,N_9922,N_8660);
or U11297 (N_11297,N_8328,N_8061);
and U11298 (N_11298,N_8925,N_8412);
nand U11299 (N_11299,N_9049,N_9666);
nand U11300 (N_11300,N_8228,N_8936);
nor U11301 (N_11301,N_8507,N_9352);
nand U11302 (N_11302,N_9955,N_9177);
and U11303 (N_11303,N_8298,N_9735);
nand U11304 (N_11304,N_9453,N_9851);
nor U11305 (N_11305,N_9833,N_8196);
and U11306 (N_11306,N_9985,N_9540);
xor U11307 (N_11307,N_8355,N_9665);
nor U11308 (N_11308,N_8620,N_8855);
and U11309 (N_11309,N_9211,N_9733);
xor U11310 (N_11310,N_8235,N_9792);
nor U11311 (N_11311,N_8831,N_9681);
xor U11312 (N_11312,N_9393,N_8481);
xnor U11313 (N_11313,N_9108,N_9703);
xor U11314 (N_11314,N_9068,N_9479);
nor U11315 (N_11315,N_8821,N_9214);
nand U11316 (N_11316,N_8278,N_8939);
nand U11317 (N_11317,N_9253,N_8974);
and U11318 (N_11318,N_9557,N_8575);
nor U11319 (N_11319,N_8699,N_9447);
xor U11320 (N_11320,N_8395,N_9824);
xnor U11321 (N_11321,N_8713,N_9512);
nor U11322 (N_11322,N_8328,N_8461);
nand U11323 (N_11323,N_9469,N_8534);
nor U11324 (N_11324,N_9022,N_8254);
or U11325 (N_11325,N_9517,N_9086);
nand U11326 (N_11326,N_8784,N_8793);
or U11327 (N_11327,N_9814,N_9752);
and U11328 (N_11328,N_8631,N_8451);
and U11329 (N_11329,N_9873,N_8254);
and U11330 (N_11330,N_8112,N_9282);
or U11331 (N_11331,N_8571,N_8088);
xor U11332 (N_11332,N_9867,N_8740);
nand U11333 (N_11333,N_9120,N_9984);
or U11334 (N_11334,N_9201,N_8251);
xor U11335 (N_11335,N_9058,N_8348);
and U11336 (N_11336,N_8546,N_9841);
or U11337 (N_11337,N_8694,N_8875);
xnor U11338 (N_11338,N_9598,N_9212);
or U11339 (N_11339,N_9073,N_9221);
or U11340 (N_11340,N_8684,N_8768);
xor U11341 (N_11341,N_8562,N_8862);
xnor U11342 (N_11342,N_9095,N_8657);
nor U11343 (N_11343,N_9777,N_9435);
xnor U11344 (N_11344,N_8839,N_9927);
and U11345 (N_11345,N_9697,N_8538);
nor U11346 (N_11346,N_9776,N_8590);
nor U11347 (N_11347,N_9058,N_9867);
nor U11348 (N_11348,N_8111,N_8245);
nand U11349 (N_11349,N_8419,N_9599);
and U11350 (N_11350,N_8690,N_9046);
xnor U11351 (N_11351,N_9305,N_9059);
xor U11352 (N_11352,N_8769,N_8424);
or U11353 (N_11353,N_8057,N_8447);
nor U11354 (N_11354,N_8071,N_9909);
nor U11355 (N_11355,N_9450,N_8764);
nand U11356 (N_11356,N_8513,N_9484);
xnor U11357 (N_11357,N_8503,N_8394);
xnor U11358 (N_11358,N_9919,N_9154);
nand U11359 (N_11359,N_9621,N_8090);
or U11360 (N_11360,N_9738,N_9553);
and U11361 (N_11361,N_8129,N_9937);
nor U11362 (N_11362,N_8136,N_9651);
or U11363 (N_11363,N_9936,N_8258);
xnor U11364 (N_11364,N_9350,N_9732);
or U11365 (N_11365,N_9024,N_9369);
nand U11366 (N_11366,N_8247,N_8787);
or U11367 (N_11367,N_9407,N_8138);
xor U11368 (N_11368,N_9951,N_8405);
xor U11369 (N_11369,N_8314,N_8838);
nor U11370 (N_11370,N_9371,N_8641);
nor U11371 (N_11371,N_9992,N_9190);
nand U11372 (N_11372,N_8124,N_9255);
nand U11373 (N_11373,N_9590,N_9120);
xnor U11374 (N_11374,N_9766,N_9720);
and U11375 (N_11375,N_8216,N_8071);
or U11376 (N_11376,N_8270,N_9184);
nand U11377 (N_11377,N_9853,N_8405);
xor U11378 (N_11378,N_8320,N_9085);
xnor U11379 (N_11379,N_8211,N_8237);
nand U11380 (N_11380,N_8899,N_8090);
xor U11381 (N_11381,N_9141,N_9228);
nand U11382 (N_11382,N_8479,N_8495);
xnor U11383 (N_11383,N_9755,N_9965);
and U11384 (N_11384,N_9437,N_9055);
xor U11385 (N_11385,N_8810,N_9899);
nand U11386 (N_11386,N_8715,N_9126);
and U11387 (N_11387,N_8493,N_9257);
nor U11388 (N_11388,N_9180,N_8068);
and U11389 (N_11389,N_9651,N_8073);
xnor U11390 (N_11390,N_8646,N_9079);
xor U11391 (N_11391,N_9726,N_9462);
nand U11392 (N_11392,N_9566,N_9935);
nor U11393 (N_11393,N_8934,N_9949);
xor U11394 (N_11394,N_9805,N_8344);
xnor U11395 (N_11395,N_9741,N_8196);
nand U11396 (N_11396,N_9218,N_8613);
nand U11397 (N_11397,N_8073,N_9142);
and U11398 (N_11398,N_9533,N_8727);
and U11399 (N_11399,N_8752,N_9200);
and U11400 (N_11400,N_8640,N_9963);
or U11401 (N_11401,N_8320,N_8326);
nor U11402 (N_11402,N_9658,N_8892);
xnor U11403 (N_11403,N_9187,N_9990);
nand U11404 (N_11404,N_9832,N_8190);
nor U11405 (N_11405,N_9400,N_8552);
xnor U11406 (N_11406,N_8304,N_8614);
or U11407 (N_11407,N_8381,N_9137);
or U11408 (N_11408,N_9648,N_9212);
and U11409 (N_11409,N_9758,N_8430);
nor U11410 (N_11410,N_9424,N_8983);
nand U11411 (N_11411,N_9130,N_8287);
nand U11412 (N_11412,N_8928,N_8276);
nand U11413 (N_11413,N_8684,N_9122);
nor U11414 (N_11414,N_8592,N_9395);
and U11415 (N_11415,N_8628,N_8176);
or U11416 (N_11416,N_9805,N_9641);
and U11417 (N_11417,N_8357,N_8917);
or U11418 (N_11418,N_9321,N_9948);
and U11419 (N_11419,N_9586,N_9868);
and U11420 (N_11420,N_8184,N_8897);
nand U11421 (N_11421,N_8384,N_8394);
or U11422 (N_11422,N_9975,N_9417);
nand U11423 (N_11423,N_8999,N_9790);
nand U11424 (N_11424,N_9372,N_9091);
nand U11425 (N_11425,N_9603,N_8441);
or U11426 (N_11426,N_8325,N_8835);
and U11427 (N_11427,N_8858,N_9623);
and U11428 (N_11428,N_8258,N_8208);
or U11429 (N_11429,N_8641,N_8995);
and U11430 (N_11430,N_9093,N_9448);
nor U11431 (N_11431,N_8746,N_9866);
xor U11432 (N_11432,N_9158,N_9728);
and U11433 (N_11433,N_8391,N_8087);
nor U11434 (N_11434,N_8638,N_8132);
or U11435 (N_11435,N_9830,N_9864);
nand U11436 (N_11436,N_9498,N_8073);
nor U11437 (N_11437,N_9922,N_9459);
nor U11438 (N_11438,N_9652,N_9807);
xor U11439 (N_11439,N_8481,N_9033);
nand U11440 (N_11440,N_8583,N_9414);
nand U11441 (N_11441,N_9342,N_9140);
and U11442 (N_11442,N_9885,N_8449);
or U11443 (N_11443,N_9077,N_8127);
nand U11444 (N_11444,N_8764,N_8584);
xor U11445 (N_11445,N_8681,N_9860);
xor U11446 (N_11446,N_9483,N_8541);
nand U11447 (N_11447,N_8985,N_9571);
xnor U11448 (N_11448,N_8301,N_8448);
nand U11449 (N_11449,N_8993,N_8252);
xnor U11450 (N_11450,N_9486,N_9313);
or U11451 (N_11451,N_8361,N_8430);
or U11452 (N_11452,N_8753,N_8692);
nand U11453 (N_11453,N_8954,N_8895);
nand U11454 (N_11454,N_8781,N_9275);
nor U11455 (N_11455,N_9346,N_8051);
xnor U11456 (N_11456,N_8700,N_9977);
xnor U11457 (N_11457,N_9856,N_9213);
xor U11458 (N_11458,N_8982,N_9292);
xor U11459 (N_11459,N_8868,N_8327);
nor U11460 (N_11460,N_8668,N_9330);
or U11461 (N_11461,N_9172,N_8627);
xnor U11462 (N_11462,N_9036,N_8596);
xor U11463 (N_11463,N_8842,N_9601);
nor U11464 (N_11464,N_8554,N_8703);
xnor U11465 (N_11465,N_9170,N_9875);
and U11466 (N_11466,N_9081,N_9645);
or U11467 (N_11467,N_8417,N_8380);
or U11468 (N_11468,N_8619,N_9574);
and U11469 (N_11469,N_8041,N_9194);
nor U11470 (N_11470,N_9971,N_8330);
nor U11471 (N_11471,N_8427,N_8597);
and U11472 (N_11472,N_9248,N_8056);
nor U11473 (N_11473,N_8445,N_9611);
nand U11474 (N_11474,N_9133,N_8704);
nor U11475 (N_11475,N_8761,N_9922);
and U11476 (N_11476,N_8651,N_8445);
and U11477 (N_11477,N_8611,N_9970);
or U11478 (N_11478,N_9632,N_8467);
nor U11479 (N_11479,N_8702,N_9295);
nor U11480 (N_11480,N_9785,N_8023);
and U11481 (N_11481,N_8787,N_9732);
nand U11482 (N_11482,N_8511,N_8174);
xor U11483 (N_11483,N_9813,N_8758);
and U11484 (N_11484,N_8648,N_8216);
or U11485 (N_11485,N_9757,N_8763);
nand U11486 (N_11486,N_8880,N_8256);
xnor U11487 (N_11487,N_8914,N_9455);
and U11488 (N_11488,N_9308,N_9340);
and U11489 (N_11489,N_9860,N_9168);
nand U11490 (N_11490,N_8182,N_8096);
or U11491 (N_11491,N_9871,N_9962);
or U11492 (N_11492,N_8485,N_9791);
nand U11493 (N_11493,N_9348,N_8068);
xor U11494 (N_11494,N_9020,N_8073);
or U11495 (N_11495,N_8273,N_8666);
nand U11496 (N_11496,N_9152,N_8829);
or U11497 (N_11497,N_9869,N_9800);
nand U11498 (N_11498,N_8301,N_8509);
nand U11499 (N_11499,N_9155,N_8506);
or U11500 (N_11500,N_9425,N_9300);
nand U11501 (N_11501,N_9512,N_8482);
nor U11502 (N_11502,N_8667,N_9858);
xor U11503 (N_11503,N_9785,N_8487);
xor U11504 (N_11504,N_8474,N_8064);
or U11505 (N_11505,N_8959,N_8008);
or U11506 (N_11506,N_8947,N_8219);
nand U11507 (N_11507,N_8861,N_8042);
nand U11508 (N_11508,N_9206,N_9958);
xnor U11509 (N_11509,N_9109,N_9845);
xor U11510 (N_11510,N_8985,N_9305);
or U11511 (N_11511,N_9331,N_9455);
nand U11512 (N_11512,N_9526,N_8021);
nand U11513 (N_11513,N_8947,N_8070);
nand U11514 (N_11514,N_8954,N_8678);
and U11515 (N_11515,N_8906,N_8416);
xor U11516 (N_11516,N_8541,N_8563);
or U11517 (N_11517,N_8217,N_9306);
or U11518 (N_11518,N_9554,N_8495);
xor U11519 (N_11519,N_8033,N_8106);
or U11520 (N_11520,N_9456,N_8328);
nand U11521 (N_11521,N_9930,N_9366);
nor U11522 (N_11522,N_8489,N_9181);
and U11523 (N_11523,N_9001,N_8241);
or U11524 (N_11524,N_8899,N_8474);
nor U11525 (N_11525,N_9973,N_9200);
or U11526 (N_11526,N_9868,N_8164);
nor U11527 (N_11527,N_9896,N_9109);
and U11528 (N_11528,N_9422,N_9032);
and U11529 (N_11529,N_9059,N_9546);
nand U11530 (N_11530,N_8278,N_9818);
or U11531 (N_11531,N_9909,N_9263);
nor U11532 (N_11532,N_8217,N_9833);
and U11533 (N_11533,N_9726,N_8897);
nand U11534 (N_11534,N_8556,N_8015);
or U11535 (N_11535,N_9127,N_8464);
nand U11536 (N_11536,N_9163,N_9051);
and U11537 (N_11537,N_8067,N_8834);
or U11538 (N_11538,N_8153,N_9006);
xnor U11539 (N_11539,N_9170,N_9185);
xor U11540 (N_11540,N_8460,N_8718);
or U11541 (N_11541,N_9270,N_8825);
or U11542 (N_11542,N_8695,N_8267);
or U11543 (N_11543,N_8933,N_9923);
nor U11544 (N_11544,N_8602,N_9829);
and U11545 (N_11545,N_9523,N_8605);
nand U11546 (N_11546,N_9232,N_8742);
xor U11547 (N_11547,N_8036,N_9768);
nor U11548 (N_11548,N_9628,N_8111);
or U11549 (N_11549,N_9112,N_8498);
nand U11550 (N_11550,N_8498,N_9914);
or U11551 (N_11551,N_8103,N_8702);
xor U11552 (N_11552,N_9681,N_9115);
xnor U11553 (N_11553,N_8991,N_9862);
nand U11554 (N_11554,N_8656,N_8355);
and U11555 (N_11555,N_9568,N_9223);
nand U11556 (N_11556,N_8225,N_8077);
nand U11557 (N_11557,N_8603,N_8956);
and U11558 (N_11558,N_8425,N_9413);
nand U11559 (N_11559,N_9437,N_8693);
nor U11560 (N_11560,N_9048,N_8985);
xor U11561 (N_11561,N_9715,N_9858);
nor U11562 (N_11562,N_8084,N_8318);
xnor U11563 (N_11563,N_8635,N_8281);
xnor U11564 (N_11564,N_9280,N_8274);
or U11565 (N_11565,N_8875,N_8080);
or U11566 (N_11566,N_9194,N_8173);
and U11567 (N_11567,N_9590,N_8046);
nand U11568 (N_11568,N_8493,N_8628);
or U11569 (N_11569,N_8131,N_9614);
nor U11570 (N_11570,N_9174,N_8466);
nor U11571 (N_11571,N_9940,N_9601);
nor U11572 (N_11572,N_9462,N_8294);
nor U11573 (N_11573,N_8119,N_8749);
or U11574 (N_11574,N_9657,N_9858);
and U11575 (N_11575,N_8590,N_9570);
xor U11576 (N_11576,N_9794,N_8473);
and U11577 (N_11577,N_9438,N_8124);
or U11578 (N_11578,N_8731,N_9968);
nand U11579 (N_11579,N_9392,N_9463);
nand U11580 (N_11580,N_9129,N_9635);
xor U11581 (N_11581,N_9216,N_8645);
and U11582 (N_11582,N_8946,N_9626);
nor U11583 (N_11583,N_9477,N_8923);
and U11584 (N_11584,N_8554,N_9419);
and U11585 (N_11585,N_9542,N_8585);
and U11586 (N_11586,N_9296,N_9062);
or U11587 (N_11587,N_8833,N_8524);
or U11588 (N_11588,N_8060,N_9060);
and U11589 (N_11589,N_8105,N_9773);
xor U11590 (N_11590,N_9400,N_9344);
nor U11591 (N_11591,N_8264,N_8690);
nor U11592 (N_11592,N_8949,N_8890);
xnor U11593 (N_11593,N_8969,N_8170);
and U11594 (N_11594,N_8582,N_8031);
nand U11595 (N_11595,N_9896,N_8904);
nor U11596 (N_11596,N_9399,N_9874);
nor U11597 (N_11597,N_9954,N_9788);
and U11598 (N_11598,N_8252,N_8352);
and U11599 (N_11599,N_8124,N_8821);
and U11600 (N_11600,N_9375,N_8617);
or U11601 (N_11601,N_8900,N_8550);
nand U11602 (N_11602,N_9007,N_9325);
xnor U11603 (N_11603,N_8348,N_9350);
nand U11604 (N_11604,N_8936,N_9895);
nor U11605 (N_11605,N_9655,N_8674);
or U11606 (N_11606,N_9548,N_8383);
xor U11607 (N_11607,N_9563,N_9330);
nand U11608 (N_11608,N_9028,N_9251);
and U11609 (N_11609,N_9023,N_8326);
nor U11610 (N_11610,N_9990,N_8273);
nor U11611 (N_11611,N_9335,N_9510);
xor U11612 (N_11612,N_9552,N_8590);
nor U11613 (N_11613,N_8285,N_9756);
and U11614 (N_11614,N_8116,N_8139);
xor U11615 (N_11615,N_8476,N_9428);
and U11616 (N_11616,N_8126,N_8827);
nand U11617 (N_11617,N_8380,N_9492);
xor U11618 (N_11618,N_9652,N_8769);
nor U11619 (N_11619,N_9988,N_9202);
nor U11620 (N_11620,N_9927,N_8246);
nor U11621 (N_11621,N_8602,N_9532);
nand U11622 (N_11622,N_8399,N_9088);
or U11623 (N_11623,N_9247,N_9276);
or U11624 (N_11624,N_9843,N_9614);
xnor U11625 (N_11625,N_9004,N_9830);
nand U11626 (N_11626,N_9686,N_8751);
nor U11627 (N_11627,N_9096,N_8067);
nand U11628 (N_11628,N_8433,N_9149);
or U11629 (N_11629,N_8420,N_8601);
nand U11630 (N_11630,N_9624,N_9144);
and U11631 (N_11631,N_8714,N_9204);
xor U11632 (N_11632,N_9135,N_8817);
nand U11633 (N_11633,N_8216,N_8123);
and U11634 (N_11634,N_9037,N_8738);
nand U11635 (N_11635,N_8841,N_9078);
xor U11636 (N_11636,N_9508,N_9171);
nor U11637 (N_11637,N_8636,N_9380);
or U11638 (N_11638,N_9533,N_9262);
nand U11639 (N_11639,N_9527,N_9438);
and U11640 (N_11640,N_9271,N_9756);
nand U11641 (N_11641,N_9241,N_8740);
nor U11642 (N_11642,N_9027,N_8416);
nand U11643 (N_11643,N_9885,N_8263);
and U11644 (N_11644,N_8692,N_8477);
or U11645 (N_11645,N_9962,N_9881);
and U11646 (N_11646,N_9637,N_8453);
nand U11647 (N_11647,N_9761,N_9132);
nor U11648 (N_11648,N_8089,N_9863);
and U11649 (N_11649,N_8436,N_9030);
nor U11650 (N_11650,N_9411,N_8196);
or U11651 (N_11651,N_8068,N_8012);
or U11652 (N_11652,N_9679,N_8020);
nor U11653 (N_11653,N_9447,N_9867);
xnor U11654 (N_11654,N_8355,N_9550);
nor U11655 (N_11655,N_9938,N_8326);
xnor U11656 (N_11656,N_9120,N_9089);
nand U11657 (N_11657,N_8141,N_8288);
or U11658 (N_11658,N_8811,N_9745);
or U11659 (N_11659,N_9573,N_8365);
nor U11660 (N_11660,N_9346,N_8777);
xnor U11661 (N_11661,N_8759,N_8212);
xnor U11662 (N_11662,N_8659,N_9927);
nand U11663 (N_11663,N_8585,N_9539);
or U11664 (N_11664,N_9069,N_8133);
or U11665 (N_11665,N_8227,N_8953);
nand U11666 (N_11666,N_9603,N_9667);
and U11667 (N_11667,N_8968,N_8982);
or U11668 (N_11668,N_8388,N_8894);
or U11669 (N_11669,N_8972,N_9169);
nand U11670 (N_11670,N_9560,N_8199);
nand U11671 (N_11671,N_8070,N_9689);
xnor U11672 (N_11672,N_9878,N_8260);
or U11673 (N_11673,N_9116,N_8424);
nand U11674 (N_11674,N_8057,N_9981);
xor U11675 (N_11675,N_9289,N_9483);
nor U11676 (N_11676,N_8360,N_9531);
and U11677 (N_11677,N_9988,N_8522);
nor U11678 (N_11678,N_8354,N_9095);
xnor U11679 (N_11679,N_9609,N_8665);
or U11680 (N_11680,N_9802,N_9817);
or U11681 (N_11681,N_8175,N_8408);
nand U11682 (N_11682,N_8493,N_8587);
xor U11683 (N_11683,N_9525,N_9320);
xor U11684 (N_11684,N_9526,N_9392);
nor U11685 (N_11685,N_8632,N_8819);
xor U11686 (N_11686,N_8050,N_9090);
and U11687 (N_11687,N_8839,N_8538);
or U11688 (N_11688,N_9645,N_9432);
and U11689 (N_11689,N_9843,N_8590);
or U11690 (N_11690,N_9994,N_9252);
or U11691 (N_11691,N_8668,N_9064);
and U11692 (N_11692,N_8548,N_8986);
xor U11693 (N_11693,N_8010,N_9708);
or U11694 (N_11694,N_9193,N_9992);
nor U11695 (N_11695,N_9250,N_8536);
or U11696 (N_11696,N_9341,N_9598);
xnor U11697 (N_11697,N_8290,N_8435);
and U11698 (N_11698,N_9793,N_8788);
xor U11699 (N_11699,N_9073,N_9330);
nand U11700 (N_11700,N_8741,N_8408);
xor U11701 (N_11701,N_8114,N_9637);
nor U11702 (N_11702,N_8423,N_8911);
nand U11703 (N_11703,N_8593,N_9513);
or U11704 (N_11704,N_8729,N_9167);
nor U11705 (N_11705,N_8515,N_9876);
or U11706 (N_11706,N_8363,N_9501);
xor U11707 (N_11707,N_9468,N_9378);
and U11708 (N_11708,N_9005,N_9104);
nand U11709 (N_11709,N_8227,N_8486);
nor U11710 (N_11710,N_9223,N_9772);
nor U11711 (N_11711,N_8700,N_9014);
nand U11712 (N_11712,N_8820,N_9800);
and U11713 (N_11713,N_8753,N_8926);
nor U11714 (N_11714,N_9375,N_8466);
and U11715 (N_11715,N_8647,N_8786);
or U11716 (N_11716,N_8974,N_9082);
nand U11717 (N_11717,N_8402,N_9085);
nor U11718 (N_11718,N_8449,N_8391);
nand U11719 (N_11719,N_8223,N_9871);
nand U11720 (N_11720,N_9270,N_8887);
xnor U11721 (N_11721,N_9563,N_8541);
xnor U11722 (N_11722,N_8539,N_9031);
nand U11723 (N_11723,N_9931,N_9716);
nor U11724 (N_11724,N_8408,N_8446);
and U11725 (N_11725,N_9640,N_9265);
nor U11726 (N_11726,N_8644,N_9126);
or U11727 (N_11727,N_8961,N_9245);
and U11728 (N_11728,N_9373,N_9408);
or U11729 (N_11729,N_9216,N_9006);
xor U11730 (N_11730,N_8931,N_9980);
xnor U11731 (N_11731,N_9359,N_9778);
xor U11732 (N_11732,N_8440,N_9615);
and U11733 (N_11733,N_8593,N_9978);
nor U11734 (N_11734,N_9052,N_8316);
nor U11735 (N_11735,N_9585,N_8256);
xnor U11736 (N_11736,N_8205,N_8319);
xnor U11737 (N_11737,N_8029,N_8564);
and U11738 (N_11738,N_9708,N_8442);
nor U11739 (N_11739,N_8918,N_9253);
nor U11740 (N_11740,N_9406,N_8699);
xor U11741 (N_11741,N_9524,N_8900);
xnor U11742 (N_11742,N_9223,N_9800);
nor U11743 (N_11743,N_8549,N_8186);
nand U11744 (N_11744,N_9350,N_9014);
or U11745 (N_11745,N_9756,N_9096);
or U11746 (N_11746,N_8075,N_9000);
nand U11747 (N_11747,N_9108,N_9180);
or U11748 (N_11748,N_8787,N_9997);
and U11749 (N_11749,N_9721,N_9257);
or U11750 (N_11750,N_9808,N_9494);
nor U11751 (N_11751,N_9467,N_8543);
or U11752 (N_11752,N_9907,N_8500);
xor U11753 (N_11753,N_8617,N_9515);
or U11754 (N_11754,N_9892,N_9096);
or U11755 (N_11755,N_9478,N_9625);
or U11756 (N_11756,N_9540,N_8896);
xor U11757 (N_11757,N_9278,N_8737);
or U11758 (N_11758,N_9027,N_9263);
and U11759 (N_11759,N_8314,N_9547);
nand U11760 (N_11760,N_9653,N_9127);
xor U11761 (N_11761,N_9565,N_9717);
nand U11762 (N_11762,N_8855,N_9058);
xnor U11763 (N_11763,N_9469,N_8345);
nor U11764 (N_11764,N_9042,N_9338);
nand U11765 (N_11765,N_8046,N_8584);
nor U11766 (N_11766,N_9202,N_9186);
xnor U11767 (N_11767,N_9264,N_8014);
xor U11768 (N_11768,N_8059,N_9743);
xnor U11769 (N_11769,N_8623,N_8121);
or U11770 (N_11770,N_9383,N_9211);
nor U11771 (N_11771,N_9468,N_9064);
nand U11772 (N_11772,N_8922,N_8021);
or U11773 (N_11773,N_8820,N_8215);
xnor U11774 (N_11774,N_9818,N_9149);
nand U11775 (N_11775,N_8759,N_9211);
nor U11776 (N_11776,N_8442,N_9368);
nand U11777 (N_11777,N_9828,N_9321);
xnor U11778 (N_11778,N_9923,N_9921);
nand U11779 (N_11779,N_8465,N_9916);
xor U11780 (N_11780,N_8999,N_9242);
nand U11781 (N_11781,N_9784,N_8920);
nor U11782 (N_11782,N_9886,N_9857);
or U11783 (N_11783,N_9612,N_8052);
and U11784 (N_11784,N_8146,N_8000);
or U11785 (N_11785,N_8420,N_8708);
nor U11786 (N_11786,N_9736,N_8951);
and U11787 (N_11787,N_9727,N_8853);
nor U11788 (N_11788,N_9865,N_8239);
or U11789 (N_11789,N_9602,N_8611);
nand U11790 (N_11790,N_9407,N_8523);
and U11791 (N_11791,N_9050,N_9341);
and U11792 (N_11792,N_8774,N_9974);
nor U11793 (N_11793,N_9777,N_9173);
xnor U11794 (N_11794,N_9866,N_9049);
nor U11795 (N_11795,N_9064,N_9255);
nand U11796 (N_11796,N_8431,N_9051);
xnor U11797 (N_11797,N_9105,N_8025);
nand U11798 (N_11798,N_9287,N_8139);
and U11799 (N_11799,N_9776,N_8416);
or U11800 (N_11800,N_9064,N_8890);
nand U11801 (N_11801,N_8661,N_9717);
nand U11802 (N_11802,N_9143,N_8115);
nor U11803 (N_11803,N_9245,N_8462);
and U11804 (N_11804,N_9337,N_9782);
or U11805 (N_11805,N_8750,N_8253);
and U11806 (N_11806,N_9778,N_9597);
nand U11807 (N_11807,N_9928,N_8460);
nor U11808 (N_11808,N_9037,N_9650);
and U11809 (N_11809,N_9432,N_8223);
xor U11810 (N_11810,N_8469,N_9599);
or U11811 (N_11811,N_9559,N_9052);
nor U11812 (N_11812,N_8470,N_9354);
xnor U11813 (N_11813,N_8426,N_9889);
nor U11814 (N_11814,N_8888,N_8867);
or U11815 (N_11815,N_9577,N_9330);
xnor U11816 (N_11816,N_9619,N_8164);
nor U11817 (N_11817,N_8328,N_9959);
nand U11818 (N_11818,N_8429,N_8491);
or U11819 (N_11819,N_8452,N_9913);
or U11820 (N_11820,N_9595,N_8053);
and U11821 (N_11821,N_8874,N_8125);
xnor U11822 (N_11822,N_9541,N_8930);
and U11823 (N_11823,N_9225,N_9653);
nand U11824 (N_11824,N_8526,N_9651);
nand U11825 (N_11825,N_9457,N_8464);
or U11826 (N_11826,N_9528,N_9245);
or U11827 (N_11827,N_9248,N_8896);
nand U11828 (N_11828,N_9018,N_8593);
nor U11829 (N_11829,N_9941,N_9815);
or U11830 (N_11830,N_8374,N_9243);
nand U11831 (N_11831,N_8299,N_9907);
xnor U11832 (N_11832,N_9214,N_8508);
xnor U11833 (N_11833,N_8188,N_9943);
and U11834 (N_11834,N_9423,N_9834);
xnor U11835 (N_11835,N_8394,N_8758);
nor U11836 (N_11836,N_9475,N_9964);
nand U11837 (N_11837,N_9430,N_8114);
xor U11838 (N_11838,N_9319,N_9182);
nor U11839 (N_11839,N_9673,N_9905);
or U11840 (N_11840,N_9325,N_9223);
and U11841 (N_11841,N_9248,N_9745);
or U11842 (N_11842,N_8810,N_9686);
nand U11843 (N_11843,N_9442,N_9600);
nor U11844 (N_11844,N_8718,N_9359);
and U11845 (N_11845,N_9782,N_9880);
and U11846 (N_11846,N_8744,N_8701);
nand U11847 (N_11847,N_9051,N_8798);
and U11848 (N_11848,N_9324,N_8649);
or U11849 (N_11849,N_8729,N_9316);
xnor U11850 (N_11850,N_9127,N_9844);
nor U11851 (N_11851,N_9723,N_9860);
and U11852 (N_11852,N_9768,N_8100);
or U11853 (N_11853,N_8388,N_8979);
and U11854 (N_11854,N_9033,N_9944);
or U11855 (N_11855,N_8305,N_9961);
and U11856 (N_11856,N_9967,N_9224);
nand U11857 (N_11857,N_9439,N_8530);
nand U11858 (N_11858,N_8470,N_8170);
nand U11859 (N_11859,N_8372,N_9776);
nor U11860 (N_11860,N_8087,N_8225);
or U11861 (N_11861,N_8277,N_9313);
nor U11862 (N_11862,N_9065,N_9255);
and U11863 (N_11863,N_9602,N_8483);
and U11864 (N_11864,N_8125,N_9189);
and U11865 (N_11865,N_8368,N_9403);
and U11866 (N_11866,N_8897,N_8042);
nand U11867 (N_11867,N_9133,N_9374);
xnor U11868 (N_11868,N_8579,N_9971);
nor U11869 (N_11869,N_8623,N_9414);
and U11870 (N_11870,N_9653,N_9237);
or U11871 (N_11871,N_8393,N_9859);
nor U11872 (N_11872,N_8498,N_8637);
xor U11873 (N_11873,N_9239,N_8638);
nor U11874 (N_11874,N_9643,N_9647);
or U11875 (N_11875,N_9540,N_8564);
and U11876 (N_11876,N_9844,N_9706);
nor U11877 (N_11877,N_8644,N_9236);
and U11878 (N_11878,N_9602,N_8729);
xnor U11879 (N_11879,N_8861,N_8954);
nor U11880 (N_11880,N_8135,N_9180);
and U11881 (N_11881,N_9882,N_9721);
xnor U11882 (N_11882,N_8706,N_8519);
nand U11883 (N_11883,N_9077,N_8251);
nor U11884 (N_11884,N_9600,N_8917);
and U11885 (N_11885,N_8732,N_8694);
or U11886 (N_11886,N_8435,N_8661);
and U11887 (N_11887,N_9620,N_8267);
nor U11888 (N_11888,N_9458,N_8805);
or U11889 (N_11889,N_8253,N_9309);
nand U11890 (N_11890,N_9598,N_9012);
nand U11891 (N_11891,N_8542,N_8070);
nor U11892 (N_11892,N_8694,N_8505);
xnor U11893 (N_11893,N_8586,N_8062);
nand U11894 (N_11894,N_9027,N_8352);
or U11895 (N_11895,N_8115,N_8224);
xor U11896 (N_11896,N_9503,N_8296);
or U11897 (N_11897,N_8227,N_8945);
and U11898 (N_11898,N_8454,N_9398);
nand U11899 (N_11899,N_9910,N_8106);
nor U11900 (N_11900,N_8040,N_8946);
nor U11901 (N_11901,N_8004,N_8078);
xnor U11902 (N_11902,N_8495,N_8542);
and U11903 (N_11903,N_8390,N_9717);
xor U11904 (N_11904,N_8351,N_9839);
nor U11905 (N_11905,N_9925,N_9722);
nor U11906 (N_11906,N_9901,N_8970);
or U11907 (N_11907,N_8583,N_8187);
and U11908 (N_11908,N_9322,N_9443);
nor U11909 (N_11909,N_8729,N_8830);
xor U11910 (N_11910,N_9858,N_8299);
or U11911 (N_11911,N_9031,N_8049);
nand U11912 (N_11912,N_8120,N_9645);
nand U11913 (N_11913,N_8099,N_8429);
or U11914 (N_11914,N_9234,N_8451);
and U11915 (N_11915,N_8288,N_9689);
nand U11916 (N_11916,N_8086,N_9191);
or U11917 (N_11917,N_8326,N_8526);
and U11918 (N_11918,N_9746,N_8518);
and U11919 (N_11919,N_9753,N_9764);
xor U11920 (N_11920,N_8531,N_8658);
or U11921 (N_11921,N_8771,N_9865);
or U11922 (N_11922,N_8307,N_8629);
and U11923 (N_11923,N_9138,N_9020);
or U11924 (N_11924,N_8257,N_9881);
nor U11925 (N_11925,N_9607,N_9624);
and U11926 (N_11926,N_8716,N_9459);
nand U11927 (N_11927,N_9861,N_9357);
nand U11928 (N_11928,N_8924,N_9561);
xnor U11929 (N_11929,N_8285,N_8155);
or U11930 (N_11930,N_9234,N_8937);
and U11931 (N_11931,N_9002,N_8159);
and U11932 (N_11932,N_8698,N_9407);
or U11933 (N_11933,N_8143,N_8976);
nand U11934 (N_11934,N_9769,N_8609);
nor U11935 (N_11935,N_8651,N_8437);
and U11936 (N_11936,N_8960,N_8521);
nor U11937 (N_11937,N_9408,N_9406);
or U11938 (N_11938,N_8153,N_8259);
or U11939 (N_11939,N_9029,N_9314);
xnor U11940 (N_11940,N_8442,N_8439);
or U11941 (N_11941,N_9097,N_9935);
xor U11942 (N_11942,N_8562,N_9007);
nand U11943 (N_11943,N_9549,N_8149);
xor U11944 (N_11944,N_8505,N_8760);
or U11945 (N_11945,N_8656,N_8361);
xnor U11946 (N_11946,N_9885,N_9866);
or U11947 (N_11947,N_9009,N_9709);
xnor U11948 (N_11948,N_9164,N_8894);
xnor U11949 (N_11949,N_9038,N_8428);
nand U11950 (N_11950,N_8788,N_9959);
and U11951 (N_11951,N_8713,N_8985);
xnor U11952 (N_11952,N_8504,N_8617);
xnor U11953 (N_11953,N_9990,N_9861);
and U11954 (N_11954,N_8650,N_8535);
xnor U11955 (N_11955,N_9230,N_8023);
or U11956 (N_11956,N_8711,N_9174);
or U11957 (N_11957,N_9420,N_9877);
nor U11958 (N_11958,N_8489,N_9546);
or U11959 (N_11959,N_9930,N_9544);
xor U11960 (N_11960,N_8382,N_9183);
nand U11961 (N_11961,N_8048,N_8187);
xnor U11962 (N_11962,N_9046,N_8283);
nor U11963 (N_11963,N_9266,N_9164);
and U11964 (N_11964,N_9500,N_8568);
nand U11965 (N_11965,N_8905,N_8893);
xor U11966 (N_11966,N_8793,N_8417);
xnor U11967 (N_11967,N_8633,N_8831);
nand U11968 (N_11968,N_9376,N_8698);
nor U11969 (N_11969,N_9240,N_8471);
xnor U11970 (N_11970,N_8858,N_9725);
nand U11971 (N_11971,N_9176,N_9765);
or U11972 (N_11972,N_8473,N_8208);
and U11973 (N_11973,N_9822,N_8067);
nor U11974 (N_11974,N_9721,N_9609);
or U11975 (N_11975,N_9045,N_8184);
nor U11976 (N_11976,N_9492,N_9949);
nor U11977 (N_11977,N_8246,N_9766);
nor U11978 (N_11978,N_9024,N_8300);
or U11979 (N_11979,N_8786,N_8760);
nand U11980 (N_11980,N_8605,N_8912);
or U11981 (N_11981,N_9494,N_9622);
nor U11982 (N_11982,N_9235,N_9232);
and U11983 (N_11983,N_8365,N_9098);
or U11984 (N_11984,N_9405,N_8523);
and U11985 (N_11985,N_8512,N_8085);
nand U11986 (N_11986,N_8274,N_9026);
or U11987 (N_11987,N_9858,N_9767);
or U11988 (N_11988,N_9252,N_8446);
or U11989 (N_11989,N_9290,N_8764);
or U11990 (N_11990,N_9844,N_9449);
nor U11991 (N_11991,N_8237,N_9901);
nor U11992 (N_11992,N_8614,N_9248);
or U11993 (N_11993,N_9616,N_8559);
or U11994 (N_11994,N_9818,N_9646);
and U11995 (N_11995,N_8695,N_9603);
or U11996 (N_11996,N_9264,N_9380);
or U11997 (N_11997,N_9706,N_8958);
nand U11998 (N_11998,N_9326,N_8983);
xnor U11999 (N_11999,N_8007,N_9922);
nor U12000 (N_12000,N_11246,N_11463);
nor U12001 (N_12001,N_10209,N_11789);
nor U12002 (N_12002,N_10824,N_10275);
nand U12003 (N_12003,N_10413,N_10897);
xnor U12004 (N_12004,N_11747,N_10126);
xor U12005 (N_12005,N_11744,N_10959);
or U12006 (N_12006,N_10798,N_10327);
and U12007 (N_12007,N_11259,N_11501);
nand U12008 (N_12008,N_11739,N_10859);
nor U12009 (N_12009,N_10265,N_11908);
xnor U12010 (N_12010,N_11869,N_10412);
or U12011 (N_12011,N_10768,N_10567);
nand U12012 (N_12012,N_10869,N_10669);
xor U12013 (N_12013,N_10432,N_11576);
or U12014 (N_12014,N_10460,N_10703);
nor U12015 (N_12015,N_11765,N_11482);
nor U12016 (N_12016,N_10304,N_11552);
nor U12017 (N_12017,N_10563,N_11047);
nand U12018 (N_12018,N_10407,N_10343);
xnor U12019 (N_12019,N_11484,N_10402);
and U12020 (N_12020,N_11123,N_11052);
xnor U12021 (N_12021,N_10152,N_10328);
and U12022 (N_12022,N_10499,N_11396);
nor U12023 (N_12023,N_11451,N_11168);
xor U12024 (N_12024,N_10292,N_11797);
or U12025 (N_12025,N_10438,N_11000);
xor U12026 (N_12026,N_11836,N_10347);
or U12027 (N_12027,N_11679,N_11401);
xnor U12028 (N_12028,N_11476,N_11738);
xnor U12029 (N_12029,N_10713,N_10358);
nor U12030 (N_12030,N_11068,N_10093);
nor U12031 (N_12031,N_10106,N_10382);
and U12032 (N_12032,N_10542,N_10877);
nand U12033 (N_12033,N_11080,N_10102);
xor U12034 (N_12034,N_10365,N_11550);
nand U12035 (N_12035,N_10040,N_10788);
nand U12036 (N_12036,N_10643,N_11289);
and U12037 (N_12037,N_11745,N_10251);
and U12038 (N_12038,N_10188,N_10868);
nand U12039 (N_12039,N_11641,N_11192);
or U12040 (N_12040,N_11893,N_10145);
nor U12041 (N_12041,N_11147,N_10659);
xor U12042 (N_12042,N_10144,N_11555);
xnor U12043 (N_12043,N_11479,N_11701);
nor U12044 (N_12044,N_11616,N_11464);
nand U12045 (N_12045,N_10689,N_11607);
nand U12046 (N_12046,N_10712,N_11545);
or U12047 (N_12047,N_11390,N_11413);
nand U12048 (N_12048,N_11216,N_11339);
nand U12049 (N_12049,N_10172,N_10325);
nand U12050 (N_12050,N_11500,N_11353);
or U12051 (N_12051,N_10790,N_10520);
nor U12052 (N_12052,N_11245,N_11958);
nor U12053 (N_12053,N_10758,N_10021);
nor U12054 (N_12054,N_11720,N_10577);
nand U12055 (N_12055,N_10383,N_11508);
xnor U12056 (N_12056,N_10227,N_10738);
nand U12057 (N_12057,N_10146,N_11428);
and U12058 (N_12058,N_11157,N_10905);
and U12059 (N_12059,N_10470,N_10579);
nand U12060 (N_12060,N_10571,N_11170);
or U12061 (N_12061,N_10418,N_10472);
nand U12062 (N_12062,N_11549,N_11467);
xnor U12063 (N_12063,N_11193,N_10084);
nand U12064 (N_12064,N_11427,N_10160);
or U12065 (N_12065,N_11696,N_10456);
nor U12066 (N_12066,N_10881,N_11323);
xnor U12067 (N_12067,N_11936,N_10598);
nor U12068 (N_12068,N_11595,N_11814);
xnor U12069 (N_12069,N_10119,N_10932);
and U12070 (N_12070,N_10071,N_11272);
and U12071 (N_12071,N_11802,N_10606);
nor U12072 (N_12072,N_11169,N_11079);
xnor U12073 (N_12073,N_11882,N_10746);
nor U12074 (N_12074,N_11903,N_10331);
nand U12075 (N_12075,N_11307,N_10849);
nor U12076 (N_12076,N_11022,N_10078);
or U12077 (N_12077,N_10793,N_11602);
xnor U12078 (N_12078,N_10170,N_10872);
and U12079 (N_12079,N_10642,N_10756);
nand U12080 (N_12080,N_11481,N_10914);
xor U12081 (N_12081,N_10506,N_11369);
and U12082 (N_12082,N_10297,N_10596);
xor U12083 (N_12083,N_11407,N_10926);
or U12084 (N_12084,N_10433,N_11772);
nand U12085 (N_12085,N_11559,N_11448);
xor U12086 (N_12086,N_10922,N_11061);
xnor U12087 (N_12087,N_11579,N_10896);
xnor U12088 (N_12088,N_10162,N_10471);
and U12089 (N_12089,N_11122,N_10175);
or U12090 (N_12090,N_11431,N_11255);
nand U12091 (N_12091,N_10018,N_11506);
nor U12092 (N_12092,N_11857,N_11196);
or U12093 (N_12093,N_10819,N_10857);
and U12094 (N_12094,N_11257,N_10385);
xor U12095 (N_12095,N_10785,N_10330);
or U12096 (N_12096,N_11241,N_11537);
and U12097 (N_12097,N_11212,N_11455);
or U12098 (N_12098,N_11891,N_10879);
xor U12099 (N_12099,N_10234,N_11194);
nand U12100 (N_12100,N_11996,N_10865);
xnor U12101 (N_12101,N_10833,N_11791);
nand U12102 (N_12102,N_11190,N_11724);
nand U12103 (N_12103,N_11689,N_10960);
nor U12104 (N_12104,N_11266,N_10646);
nand U12105 (N_12105,N_10769,N_11183);
and U12106 (N_12106,N_10120,N_11864);
or U12107 (N_12107,N_10786,N_11906);
xnor U12108 (N_12108,N_10381,N_10201);
and U12109 (N_12109,N_11648,N_10714);
or U12110 (N_12110,N_11449,N_11094);
or U12111 (N_12111,N_10233,N_10452);
nor U12112 (N_12112,N_10090,N_10741);
xor U12113 (N_12113,N_11415,N_11297);
nand U12114 (N_12114,N_10259,N_11767);
or U12115 (N_12115,N_11828,N_11851);
or U12116 (N_12116,N_11106,N_10086);
nand U12117 (N_12117,N_11182,N_11362);
nand U12118 (N_12118,N_10094,N_11329);
or U12119 (N_12119,N_11005,N_11944);
or U12120 (N_12120,N_11780,N_11581);
or U12121 (N_12121,N_11280,N_10183);
xnor U12122 (N_12122,N_10522,N_11900);
and U12123 (N_12123,N_11139,N_10332);
xnor U12124 (N_12124,N_11217,N_11790);
or U12125 (N_12125,N_10489,N_10414);
or U12126 (N_12126,N_11447,N_11554);
or U12127 (N_12127,N_10361,N_10197);
and U12128 (N_12128,N_11404,N_11543);
and U12129 (N_12129,N_11824,N_10444);
and U12130 (N_12130,N_10931,N_10295);
or U12131 (N_12131,N_10067,N_10009);
or U12132 (N_12132,N_10037,N_10864);
or U12133 (N_12133,N_11349,N_10687);
xor U12134 (N_12134,N_11165,N_10129);
nand U12135 (N_12135,N_10561,N_10633);
nor U12136 (N_12136,N_10566,N_10799);
nor U12137 (N_12137,N_11760,N_10097);
xnor U12138 (N_12138,N_10987,N_11435);
nor U12139 (N_12139,N_10620,N_11995);
xor U12140 (N_12140,N_10813,N_10436);
nor U12141 (N_12141,N_11303,N_11888);
or U12142 (N_12142,N_10440,N_10986);
nand U12143 (N_12143,N_10509,N_11116);
xor U12144 (N_12144,N_11728,N_11854);
xor U12145 (N_12145,N_11606,N_10462);
nand U12146 (N_12146,N_11432,N_10848);
and U12147 (N_12147,N_11074,N_11174);
or U12148 (N_12148,N_10716,N_11810);
nor U12149 (N_12149,N_11110,N_10366);
or U12150 (N_12150,N_10230,N_10928);
nand U12151 (N_12151,N_11541,N_10280);
nor U12152 (N_12152,N_11097,N_10692);
nor U12153 (N_12153,N_10377,N_10762);
xor U12154 (N_12154,N_10116,N_11643);
or U12155 (N_12155,N_11815,N_10903);
and U12156 (N_12156,N_10518,N_11918);
or U12157 (N_12157,N_11914,N_10150);
xor U12158 (N_12158,N_10795,N_11222);
xnor U12159 (N_12159,N_10764,N_11997);
or U12160 (N_12160,N_11151,N_11529);
and U12161 (N_12161,N_11633,N_10809);
nand U12162 (N_12162,N_10752,N_11593);
or U12163 (N_12163,N_10161,N_11951);
xor U12164 (N_12164,N_11285,N_10484);
xor U12165 (N_12165,N_11667,N_10323);
nor U12166 (N_12166,N_11710,N_10973);
xnor U12167 (N_12167,N_11743,N_11355);
nor U12168 (N_12168,N_10006,N_10671);
and U12169 (N_12169,N_10469,N_10238);
nand U12170 (N_12170,N_11370,N_10613);
or U12171 (N_12171,N_11034,N_10783);
xor U12172 (N_12172,N_11262,N_11597);
and U12173 (N_12173,N_11322,N_10027);
and U12174 (N_12174,N_11265,N_10655);
xnor U12175 (N_12175,N_10013,N_10396);
and U12176 (N_12176,N_10668,N_11298);
or U12177 (N_12177,N_10417,N_10709);
nor U12178 (N_12178,N_10774,N_11735);
or U12179 (N_12179,N_11820,N_11316);
or U12180 (N_12180,N_10455,N_10157);
nand U12181 (N_12181,N_10254,N_11440);
xnor U12182 (N_12182,N_11998,N_11220);
and U12183 (N_12183,N_10476,N_11081);
or U12184 (N_12184,N_10354,N_11395);
and U12185 (N_12185,N_10371,N_11938);
and U12186 (N_12186,N_11675,N_11125);
nor U12187 (N_12187,N_10125,N_10490);
and U12188 (N_12188,N_10012,N_10014);
nand U12189 (N_12189,N_10723,N_11837);
nand U12190 (N_12190,N_10461,N_10908);
or U12191 (N_12191,N_10832,N_10672);
or U12192 (N_12192,N_10039,N_11055);
nor U12193 (N_12193,N_11637,N_10670);
nand U12194 (N_12194,N_11546,N_11293);
nand U12195 (N_12195,N_10486,N_11184);
xnor U12196 (N_12196,N_11060,N_11892);
nand U12197 (N_12197,N_10581,N_10171);
nand U12198 (N_12198,N_10511,N_11776);
nand U12199 (N_12199,N_10543,N_11325);
nor U12200 (N_12200,N_11713,N_10590);
and U12201 (N_12201,N_11987,N_10838);
nand U12202 (N_12202,N_11371,N_10165);
or U12203 (N_12203,N_10674,N_11126);
nand U12204 (N_12204,N_11750,N_10473);
nor U12205 (N_12205,N_10258,N_10728);
or U12206 (N_12206,N_10825,N_10479);
and U12207 (N_12207,N_11487,N_11964);
nor U12208 (N_12208,N_11982,N_11173);
or U12209 (N_12209,N_11567,N_10141);
xnor U12210 (N_12210,N_11980,N_10302);
nand U12211 (N_12211,N_11528,N_11947);
or U12212 (N_12212,N_10963,N_10441);
nor U12213 (N_12213,N_11916,N_11089);
xnor U12214 (N_12214,N_10336,N_11650);
xnor U12215 (N_12215,N_11140,N_11494);
or U12216 (N_12216,N_11294,N_11300);
nand U12217 (N_12217,N_11187,N_11002);
nand U12218 (N_12218,N_11681,N_10187);
nor U12219 (N_12219,N_10337,N_10420);
or U12220 (N_12220,N_11013,N_10095);
xor U12221 (N_12221,N_10537,N_10691);
xnor U12222 (N_12222,N_10025,N_10059);
and U12223 (N_12223,N_11418,N_10992);
nor U12224 (N_12224,N_11990,N_11066);
xor U12225 (N_12225,N_11093,N_10777);
xnor U12226 (N_12226,N_10058,N_10404);
xor U12227 (N_12227,N_11269,N_11845);
nand U12228 (N_12228,N_10195,N_11970);
xnor U12229 (N_12229,N_10164,N_11751);
and U12230 (N_12230,N_11993,N_11831);
nor U12231 (N_12231,N_11346,N_11913);
and U12232 (N_12232,N_10154,N_11770);
xnor U12233 (N_12233,N_11178,N_10508);
nor U12234 (N_12234,N_11364,N_11227);
and U12235 (N_12235,N_11589,N_11514);
xor U12236 (N_12236,N_10005,N_10271);
nand U12237 (N_12237,N_11497,N_10463);
or U12238 (N_12238,N_10350,N_10378);
and U12239 (N_12239,N_11261,N_11665);
and U12240 (N_12240,N_11977,N_10285);
xnor U12241 (N_12241,N_11965,N_11969);
xnor U12242 (N_12242,N_11087,N_11839);
or U12243 (N_12243,N_10887,N_10589);
nand U12244 (N_12244,N_10065,N_10950);
and U12245 (N_12245,N_10697,N_11287);
xnor U12246 (N_12246,N_10784,N_11522);
and U12247 (N_12247,N_11305,N_11012);
or U12248 (N_12248,N_10423,N_10092);
or U12249 (N_12249,N_11561,N_10351);
or U12250 (N_12250,N_11832,N_11741);
and U12251 (N_12251,N_10446,N_10226);
xnor U12252 (N_12252,N_10079,N_10624);
or U12253 (N_12253,N_11657,N_10000);
nor U12254 (N_12254,N_10720,N_10657);
nor U12255 (N_12255,N_11161,N_11356);
nand U12256 (N_12256,N_10411,N_11368);
and U12257 (N_12257,N_10996,N_10569);
xor U12258 (N_12258,N_11644,N_10046);
xor U12259 (N_12259,N_11748,N_11692);
and U12260 (N_12260,N_11250,N_11100);
and U12261 (N_12261,N_10318,N_10442);
xor U12262 (N_12262,N_11258,N_11450);
or U12263 (N_12263,N_10649,N_11027);
xnor U12264 (N_12264,N_10826,N_10866);
and U12265 (N_12265,N_11510,N_10211);
nor U12266 (N_12266,N_11185,N_11758);
and U12267 (N_12267,N_11134,N_10246);
nand U12268 (N_12268,N_11578,N_11408);
nand U12269 (N_12269,N_10317,N_11434);
xor U12270 (N_12270,N_11822,N_11752);
nor U12271 (N_12271,N_10443,N_11984);
and U12272 (N_12272,N_11830,N_11700);
and U12273 (N_12273,N_11483,N_11131);
xnor U12274 (N_12274,N_11694,N_11721);
and U12275 (N_12275,N_11896,N_11053);
nor U12276 (N_12276,N_11623,N_10507);
or U12277 (N_12277,N_10780,N_10754);
and U12278 (N_12278,N_10816,N_11605);
xor U12279 (N_12279,N_10368,N_10883);
nand U12280 (N_12280,N_11782,N_10426);
xnor U12281 (N_12281,N_10514,N_11507);
and U12282 (N_12282,N_11073,N_10525);
xor U12283 (N_12283,N_11237,N_11551);
nor U12284 (N_12284,N_11345,N_10629);
and U12285 (N_12285,N_10699,N_10829);
nor U12286 (N_12286,N_10736,N_11860);
nor U12287 (N_12287,N_11117,N_11105);
and U12288 (N_12288,N_10193,N_10186);
or U12289 (N_12289,N_10863,N_11474);
or U12290 (N_12290,N_11453,N_11684);
nor U12291 (N_12291,N_11024,N_11344);
and U12292 (N_12292,N_10968,N_11175);
xnor U12293 (N_12293,N_11712,N_10345);
xnor U12294 (N_12294,N_11273,N_11711);
or U12295 (N_12295,N_10818,N_10431);
nand U12296 (N_12296,N_11583,N_11264);
or U12297 (N_12297,N_11804,N_10437);
nor U12298 (N_12298,N_10972,N_11624);
nand U12299 (N_12299,N_11978,N_10177);
and U12300 (N_12300,N_10132,N_11441);
nand U12301 (N_12301,N_10815,N_11314);
nor U12302 (N_12302,N_10453,N_10936);
or U12303 (N_12303,N_10004,N_10555);
or U12304 (N_12304,N_11382,N_11668);
or U12305 (N_12305,N_11600,N_10406);
or U12306 (N_12306,N_10121,N_11871);
nor U12307 (N_12307,N_10978,N_10134);
nor U12308 (N_12308,N_11331,N_11392);
nand U12309 (N_12309,N_11366,N_10158);
xor U12310 (N_12310,N_10107,N_10306);
nor U12311 (N_12311,N_11211,N_10273);
xor U12312 (N_12312,N_10386,N_10237);
and U12313 (N_12313,N_10850,N_10862);
or U12314 (N_12314,N_10007,N_10390);
or U12315 (N_12315,N_11321,N_10895);
and U12316 (N_12316,N_11564,N_11516);
and U12317 (N_12317,N_10278,N_11278);
and U12318 (N_12318,N_10966,N_10847);
nor U12319 (N_12319,N_10958,N_10787);
or U12320 (N_12320,N_10951,N_11729);
or U12321 (N_12321,N_10684,N_11253);
nand U12322 (N_12322,N_10459,N_11863);
xnor U12323 (N_12323,N_10900,N_10047);
or U12324 (N_12324,N_10889,N_11957);
xor U12325 (N_12325,N_10844,N_11788);
nor U12326 (N_12326,N_11717,N_10512);
nand U12327 (N_12327,N_11685,N_11638);
xor U12328 (N_12328,N_10261,N_10010);
xor U12329 (N_12329,N_10051,N_10289);
nor U12330 (N_12330,N_10155,N_10944);
and U12331 (N_12331,N_11778,N_11517);
nand U12332 (N_12332,N_10989,N_11023);
and U12333 (N_12333,N_11381,N_11697);
xor U12334 (N_12334,N_11092,N_10398);
and U12335 (N_12335,N_10458,N_11631);
nor U12336 (N_12336,N_11628,N_11911);
xnor U12337 (N_12337,N_10220,N_10856);
and U12338 (N_12338,N_11994,N_10885);
nand U12339 (N_12339,N_11932,N_11242);
nand U12340 (N_12340,N_10749,N_11688);
and U12341 (N_12341,N_10319,N_11838);
xor U12342 (N_12342,N_11847,N_10400);
nor U12343 (N_12343,N_11252,N_11239);
nand U12344 (N_12344,N_10792,N_10673);
nor U12345 (N_12345,N_11313,N_10503);
and U12346 (N_12346,N_10878,N_10370);
nor U12347 (N_12347,N_11466,N_11210);
nand U12348 (N_12348,N_11843,N_10759);
nor U12349 (N_12349,N_10029,N_11787);
nor U12350 (N_12350,N_10820,N_11099);
nor U12351 (N_12351,N_11730,N_10266);
xnor U12352 (N_12352,N_11683,N_10800);
nor U12353 (N_12353,N_10449,N_10487);
or U12354 (N_12354,N_11894,N_10257);
and U12355 (N_12355,N_10312,N_11332);
nor U12356 (N_12356,N_10727,N_11586);
or U12357 (N_12357,N_11416,N_11063);
and U12358 (N_12358,N_11887,N_11340);
and U12359 (N_12359,N_11394,N_11146);
nand U12360 (N_12360,N_11458,N_11009);
xnor U12361 (N_12361,N_10946,N_10239);
nor U12362 (N_12362,N_11764,N_10942);
xnor U12363 (N_12363,N_10218,N_11723);
xnor U12364 (N_12364,N_11251,N_11925);
xnor U12365 (N_12365,N_11477,N_11571);
nor U12366 (N_12366,N_10696,N_10056);
nand U12367 (N_12367,N_10305,N_10212);
or U12368 (N_12368,N_11619,N_10801);
nand U12369 (N_12369,N_10464,N_11542);
xor U12370 (N_12370,N_11872,N_10299);
or U12371 (N_12371,N_11138,N_10105);
and U12372 (N_12372,N_10262,N_11766);
nand U12373 (N_12373,N_11438,N_10976);
nand U12374 (N_12374,N_11704,N_11403);
nand U12375 (N_12375,N_11703,N_11335);
nor U12376 (N_12376,N_11493,N_10185);
xnor U12377 (N_12377,N_11284,N_10538);
or U12378 (N_12378,N_11682,N_11103);
xnor U12379 (N_12379,N_11402,N_11164);
xnor U12380 (N_12380,N_10990,N_11861);
or U12381 (N_12381,N_10477,N_11221);
nand U12382 (N_12382,N_10810,N_10772);
and U12383 (N_12383,N_10982,N_11195);
xnor U12384 (N_12384,N_10085,N_10584);
nand U12385 (N_12385,N_10861,N_10724);
xor U12386 (N_12386,N_11560,N_11823);
nor U12387 (N_12387,N_11565,N_11557);
or U12388 (N_12388,N_10704,N_11933);
or U12389 (N_12389,N_10711,N_11727);
nand U12390 (N_12390,N_10307,N_10880);
or U12391 (N_12391,N_11498,N_10991);
nor U12392 (N_12392,N_11538,N_10910);
xnor U12393 (N_12393,N_10544,N_10702);
nor U12394 (N_12394,N_10855,N_10448);
xor U12395 (N_12395,N_10834,N_11071);
or U12396 (N_12396,N_10811,N_10353);
nor U12397 (N_12397,N_11150,N_11746);
nand U12398 (N_12398,N_10781,N_11393);
nor U12399 (N_12399,N_11422,N_11875);
nand U12400 (N_12400,N_10214,N_10002);
or U12401 (N_12401,N_10725,N_11862);
nand U12402 (N_12402,N_11291,N_11330);
and U12403 (N_12403,N_11952,N_11599);
nand U12404 (N_12404,N_10372,N_10148);
xor U12405 (N_12405,N_11879,N_10405);
nor U12406 (N_12406,N_10267,N_10531);
xor U12407 (N_12407,N_11274,N_10279);
nand U12408 (N_12408,N_11189,N_11378);
nor U12409 (N_12409,N_11399,N_10957);
or U12410 (N_12410,N_11234,N_11950);
and U12411 (N_12411,N_10817,N_10902);
xor U12412 (N_12412,N_10778,N_11032);
and U12413 (N_12413,N_10779,N_10964);
or U12414 (N_12414,N_10574,N_10159);
and U12415 (N_12415,N_10970,N_10551);
and U12416 (N_12416,N_11243,N_10424);
nor U12417 (N_12417,N_10054,N_11342);
xnor U12418 (N_12418,N_11256,N_10562);
nand U12419 (N_12419,N_10814,N_11975);
xor U12420 (N_12420,N_11136,N_10871);
and U12421 (N_12421,N_11124,N_11905);
or U12422 (N_12422,N_11634,N_10595);
and U12423 (N_12423,N_11031,N_10938);
or U12424 (N_12424,N_10314,N_10594);
xor U12425 (N_12425,N_10494,N_11373);
nor U12426 (N_12426,N_11144,N_10203);
or U12427 (N_12427,N_10073,N_11065);
nand U12428 (N_12428,N_10168,N_11142);
nor U12429 (N_12429,N_10099,N_11304);
xor U12430 (N_12430,N_10705,N_11375);
xor U12431 (N_12431,N_11445,N_10231);
xor U12432 (N_12432,N_11611,N_10533);
xor U12433 (N_12433,N_11948,N_10342);
nor U12434 (N_12434,N_11041,N_11354);
nor U12435 (N_12435,N_11229,N_11632);
or U12436 (N_12436,N_10894,N_11755);
nor U12437 (N_12437,N_10393,N_11763);
or U12438 (N_12438,N_10835,N_11020);
and U12439 (N_12439,N_10008,N_10096);
and U12440 (N_12440,N_10204,N_10173);
nand U12441 (N_12441,N_10425,N_10925);
and U12442 (N_12442,N_11320,N_11591);
nand U12443 (N_12443,N_10287,N_11946);
and U12444 (N_12444,N_10416,N_10650);
and U12445 (N_12445,N_11495,N_10283);
and U12446 (N_12446,N_10961,N_11885);
and U12447 (N_12447,N_11945,N_10252);
and U12448 (N_12448,N_11676,N_10632);
nand U12449 (N_12449,N_10929,N_11646);
nand U12450 (N_12450,N_11505,N_11430);
and U12451 (N_12451,N_10049,N_11014);
nand U12452 (N_12452,N_11942,N_10721);
or U12453 (N_12453,N_10242,N_10174);
or U12454 (N_12454,N_11577,N_11459);
xor U12455 (N_12455,N_11405,N_10391);
nand U12456 (N_12456,N_11460,N_11365);
xnor U12457 (N_12457,N_11825,N_10955);
or U12458 (N_12458,N_10591,N_11328);
nand U12459 (N_12459,N_11301,N_10851);
or U12460 (N_12460,N_10344,N_11640);
xor U12461 (N_12461,N_10726,N_10118);
and U12462 (N_12462,N_10110,N_10136);
or U12463 (N_12463,N_10559,N_11028);
and U12464 (N_12464,N_10886,N_11203);
nand U12465 (N_12465,N_10535,N_10549);
or U12466 (N_12466,N_10645,N_11732);
nor U12467 (N_12467,N_10526,N_10628);
nor U12468 (N_12468,N_11171,N_11806);
or U12469 (N_12469,N_10715,N_10748);
and U12470 (N_12470,N_11197,N_10546);
xnor U12471 (N_12471,N_10677,N_10042);
nor U12472 (N_12472,N_11469,N_11004);
xnor U12473 (N_12473,N_10892,N_11604);
and U12474 (N_12474,N_10899,N_11930);
nand U12475 (N_12475,N_11671,N_10087);
nand U12476 (N_12476,N_10623,N_10468);
nand U12477 (N_12477,N_10256,N_11818);
nor U12478 (N_12478,N_10064,N_10495);
nor U12479 (N_12479,N_11708,N_11215);
nand U12480 (N_12480,N_11343,N_10355);
nand U12481 (N_12481,N_11058,N_11919);
nor U12482 (N_12482,N_11488,N_11846);
or U12483 (N_12483,N_11442,N_11902);
or U12484 (N_12484,N_10497,N_10918);
and U12485 (N_12485,N_10969,N_10683);
or U12486 (N_12486,N_11127,N_11113);
xor U12487 (N_12487,N_11254,N_11992);
and U12488 (N_12488,N_11691,N_10196);
and U12489 (N_12489,N_11275,N_10131);
nor U12490 (N_12490,N_11615,N_11426);
xnor U12491 (N_12491,N_11201,N_10352);
and U12492 (N_12492,N_11090,N_11793);
nor U12493 (N_12493,N_10182,N_10066);
nor U12494 (N_12494,N_10482,N_11535);
nand U12495 (N_12495,N_10023,N_10399);
or U12496 (N_12496,N_11033,N_11709);
nor U12497 (N_12497,N_10644,N_10744);
xor U12498 (N_12498,N_10180,N_11974);
nand U12499 (N_12499,N_10891,N_11928);
or U12500 (N_12500,N_11104,N_10707);
xor U12501 (N_12501,N_10374,N_10167);
xnor U12502 (N_12502,N_11636,N_11207);
and U12503 (N_12503,N_10339,N_11799);
and U12504 (N_12504,N_10791,N_10088);
nand U12505 (N_12505,N_10206,N_10367);
xor U12506 (N_12506,N_11686,N_11901);
or U12507 (N_12507,N_10913,N_11412);
nor U12508 (N_12508,N_11645,N_10260);
nor U12509 (N_12509,N_11475,N_11943);
or U12510 (N_12510,N_10422,N_11042);
nor U12511 (N_12511,N_11054,N_11608);
or U12512 (N_12512,N_11398,N_11177);
nor U12513 (N_12513,N_10451,N_10030);
nor U12514 (N_12514,N_10755,N_11209);
or U12515 (N_12515,N_10101,N_10600);
xnor U12516 (N_12516,N_10994,N_11695);
xor U12517 (N_12517,N_10445,N_11417);
xnor U12518 (N_12518,N_11898,N_11573);
xnor U12519 (N_12519,N_11937,N_11228);
nor U12520 (N_12520,N_11098,N_10293);
or U12521 (N_12521,N_11006,N_10583);
and U12522 (N_12522,N_11045,N_11470);
nor U12523 (N_12523,N_11961,N_11397);
nor U12524 (N_12524,N_11036,N_10114);
or U12525 (N_12525,N_10607,N_10698);
nand U12526 (N_12526,N_11276,N_10225);
or U12527 (N_12527,N_10357,N_10191);
nor U12528 (N_12528,N_10139,N_10622);
or U12529 (N_12529,N_11967,N_10428);
or U12530 (N_12530,N_10708,N_11421);
xnor U12531 (N_12531,N_11621,N_11226);
or U12532 (N_12532,N_10060,N_11248);
and U12533 (N_12533,N_11603,N_11075);
or U12534 (N_12534,N_10338,N_11102);
nand U12535 (N_12535,N_11333,N_11912);
nand U12536 (N_12536,N_11076,N_10286);
nor U12537 (N_12537,N_10019,N_10024);
nand U12538 (N_12538,N_11794,N_11046);
nor U12539 (N_12539,N_11518,N_10117);
or U12540 (N_12540,N_10682,N_11069);
and U12541 (N_12541,N_11654,N_10830);
and U12542 (N_12542,N_11889,N_11829);
xor U12543 (N_12543,N_11468,N_11674);
nor U12544 (N_12544,N_10893,N_11338);
xnor U12545 (N_12545,N_11897,N_10200);
nand U12546 (N_12546,N_10717,N_11048);
nor U12547 (N_12547,N_11181,N_10128);
and U12548 (N_12548,N_11205,N_10143);
and U12549 (N_12549,N_10465,N_11377);
nand U12550 (N_12550,N_10403,N_10450);
nor U12551 (N_12551,N_11761,N_10586);
xnor U12552 (N_12552,N_10032,N_10072);
or U12553 (N_12553,N_10770,N_11267);
or U12554 (N_12554,N_10408,N_10733);
or U12555 (N_12555,N_11706,N_11472);
and U12556 (N_12556,N_10983,N_11334);
nor U12557 (N_12557,N_11374,N_10732);
or U12558 (N_12558,N_10205,N_11480);
nor U12559 (N_12559,N_10812,N_10977);
and U12560 (N_12560,N_10631,N_11319);
nand U12561 (N_12561,N_10492,N_10035);
or U12562 (N_12562,N_10701,N_10565);
or U12563 (N_12563,N_10311,N_11792);
nand U12564 (N_12564,N_10324,N_11580);
nand U12565 (N_12565,N_10521,N_11379);
or U12566 (N_12566,N_10656,N_10127);
nand U12567 (N_12567,N_10827,N_10653);
or U12568 (N_12568,N_11533,N_11292);
and U12569 (N_12569,N_10028,N_11176);
xor U12570 (N_12570,N_10467,N_11086);
and U12571 (N_12571,N_10041,N_10553);
xnor U12572 (N_12572,N_11849,N_10975);
or U12573 (N_12573,N_10580,N_11224);
and U12574 (N_12574,N_10907,N_11812);
or U12575 (N_12575,N_10916,N_10498);
and U12576 (N_12576,N_11740,N_11909);
xor U12577 (N_12577,N_11341,N_10410);
xor U12578 (N_12578,N_10548,N_10055);
nor U12579 (N_12579,N_11114,N_10303);
xor U12580 (N_12580,N_10447,N_10466);
xor U12581 (N_12581,N_11437,N_11163);
nand U12582 (N_12582,N_11295,N_11841);
nand U12583 (N_12583,N_10906,N_11568);
and U12584 (N_12584,N_11852,N_10300);
nand U12585 (N_12585,N_10076,N_10612);
or U12586 (N_12586,N_10034,N_10272);
or U12587 (N_12587,N_11762,N_10547);
xor U12588 (N_12588,N_11935,N_11547);
nor U12589 (N_12589,N_11673,N_10089);
or U12590 (N_12590,N_11154,N_10380);
nor U12591 (N_12591,N_11072,N_10967);
nor U12592 (N_12592,N_10516,N_10648);
xnor U12593 (N_12593,N_11652,N_11376);
nor U12594 (N_12594,N_10217,N_10409);
nor U12595 (N_12595,N_10585,N_10316);
and U12596 (N_12596,N_11091,N_10228);
xnor U12597 (N_12597,N_11202,N_11283);
nand U12598 (N_12598,N_10340,N_10038);
nand U12599 (N_12599,N_11553,N_10806);
or U12600 (N_12600,N_10757,N_11499);
nand U12601 (N_12601,N_10943,N_10888);
or U12602 (N_12602,N_11927,N_11452);
xnor U12603 (N_12603,N_11312,N_11409);
xor U12604 (N_12604,N_11380,N_11191);
xnor U12605 (N_12605,N_10510,N_11954);
xor U12606 (N_12606,N_10288,N_10582);
xnor U12607 (N_12607,N_10322,N_10681);
and U12608 (N_12608,N_11742,N_10082);
or U12609 (N_12609,N_10387,N_11238);
nor U12610 (N_12610,N_11083,N_11813);
or U12611 (N_12611,N_11647,N_11214);
nand U12612 (N_12612,N_11981,N_11953);
or U12613 (N_12613,N_10805,N_10541);
or U12614 (N_12614,N_11698,N_10232);
nor U12615 (N_12615,N_10676,N_10001);
nor U12616 (N_12616,N_11218,N_11800);
or U12617 (N_12617,N_11859,N_11240);
nor U12618 (N_12618,N_10636,N_10142);
nand U12619 (N_12619,N_10807,N_11347);
and U12620 (N_12620,N_10773,N_10839);
and U12621 (N_12621,N_11955,N_10822);
nand U12622 (N_12622,N_10276,N_11156);
xor U12623 (N_12623,N_10363,N_10695);
xnor U12624 (N_12624,N_11419,N_11811);
xnor U12625 (N_12625,N_10349,N_11360);
nand U12626 (N_12626,N_11590,N_10763);
nor U12627 (N_12627,N_11922,N_11425);
nand U12628 (N_12628,N_10053,N_10528);
nand U12629 (N_12629,N_10937,N_11388);
nand U12630 (N_12630,N_10255,N_10882);
or U12631 (N_12631,N_11574,N_11050);
or U12632 (N_12632,N_10123,N_11318);
nand U12633 (N_12633,N_11309,N_10923);
and U12634 (N_12634,N_11456,N_11223);
nand U12635 (N_12635,N_10294,N_11135);
and U12636 (N_12636,N_11337,N_10026);
or U12637 (N_12637,N_11021,N_10326);
xor U12638 (N_12638,N_11722,N_11629);
xnor U12639 (N_12639,N_11921,N_11786);
or U12640 (N_12640,N_11876,N_11690);
nor U12641 (N_12641,N_11523,N_10022);
xnor U12642 (N_12642,N_11798,N_10854);
xnor U12643 (N_12643,N_11999,N_11311);
nor U12644 (N_12644,N_10240,N_10475);
nor U12645 (N_12645,N_11705,N_11907);
and U12646 (N_12646,N_10803,N_10804);
and U12647 (N_12647,N_10052,N_11129);
nand U12648 (N_12648,N_10320,N_11734);
and U12649 (N_12649,N_11988,N_10999);
nor U12650 (N_12650,N_11400,N_10103);
xnor U12651 (N_12651,N_11513,N_10480);
xor U12652 (N_12652,N_10971,N_10842);
xnor U12653 (N_12653,N_10179,N_11886);
xor U12654 (N_12654,N_11454,N_10917);
xor U12655 (N_12655,N_11527,N_11569);
and U12656 (N_12656,N_10213,N_10904);
nor U12657 (N_12657,N_11043,N_10223);
nor U12658 (N_12658,N_10927,N_11049);
xor U12659 (N_12659,N_10135,N_11917);
and U12660 (N_12660,N_11856,N_11233);
xor U12661 (N_12661,N_10641,N_11598);
nor U12662 (N_12662,N_10578,N_10069);
or U12663 (N_12663,N_11317,N_11231);
or U12664 (N_12664,N_10678,N_11971);
or U12665 (N_12665,N_11348,N_11358);
xnor U12666 (N_12666,N_10635,N_11120);
or U12667 (N_12667,N_10153,N_11923);
or U12668 (N_12668,N_10074,N_10930);
xor U12669 (N_12669,N_10245,N_10313);
nand U12670 (N_12670,N_11044,N_11617);
nand U12671 (N_12671,N_10694,N_10729);
nor U12672 (N_12672,N_11659,N_10933);
or U12673 (N_12673,N_11920,N_11130);
xnor U12674 (N_12674,N_10647,N_11084);
nand U12675 (N_12675,N_11834,N_10427);
xor U12676 (N_12676,N_10282,N_10109);
nand U12677 (N_12677,N_11244,N_11848);
xnor U12678 (N_12678,N_11433,N_10831);
xor U12679 (N_12679,N_11627,N_10767);
nor U12680 (N_12680,N_10199,N_10524);
or U12681 (N_12681,N_10771,N_11635);
nor U12682 (N_12682,N_10823,N_11736);
or U12683 (N_12683,N_10356,N_10224);
or U12684 (N_12684,N_11384,N_10667);
and U12685 (N_12685,N_10921,N_10952);
nor U12686 (N_12686,N_11485,N_11357);
nand U12687 (N_12687,N_10333,N_11962);
and U12688 (N_12688,N_10710,N_11979);
and U12689 (N_12689,N_11367,N_11152);
nor U12690 (N_12690,N_11436,N_10236);
nand U12691 (N_12691,N_11067,N_11282);
nand U12692 (N_12692,N_11017,N_11059);
and U12693 (N_12693,N_10080,N_10794);
xor U12694 (N_12694,N_10250,N_11056);
or U12695 (N_12695,N_11471,N_11853);
or U12696 (N_12696,N_11754,N_11949);
or U12697 (N_12697,N_11610,N_10296);
or U12698 (N_12698,N_11940,N_11062);
and U12699 (N_12699,N_11959,N_10614);
nand U12700 (N_12700,N_10853,N_11963);
or U12701 (N_12701,N_11878,N_10965);
xnor U12702 (N_12702,N_11016,N_11145);
nand U12703 (N_12703,N_10836,N_10602);
xor U12704 (N_12704,N_10775,N_11026);
nand U12705 (N_12705,N_11784,N_11768);
nand U12706 (N_12706,N_11842,N_10821);
nor U12707 (N_12707,N_11934,N_10947);
nor U12708 (N_12708,N_11263,N_10540);
xnor U12709 (N_12709,N_11363,N_10530);
or U12710 (N_12710,N_10750,N_11614);
xor U12711 (N_12711,N_11389,N_10321);
or U12712 (N_12712,N_10169,N_11410);
and U12713 (N_12713,N_11286,N_11350);
nor U12714 (N_12714,N_11661,N_11926);
nor U12715 (N_12715,N_10315,N_10846);
nand U12716 (N_12716,N_10401,N_10760);
and U12717 (N_12717,N_10638,N_11383);
or U12718 (N_12718,N_10015,N_11230);
xor U12719 (N_12719,N_10140,N_11167);
xnor U12720 (N_12720,N_11877,N_11530);
and U12721 (N_12721,N_11796,N_10940);
nand U12722 (N_12722,N_10115,N_10216);
nor U12723 (N_12723,N_10501,N_11411);
and U12724 (N_12724,N_10301,N_11502);
nand U12725 (N_12725,N_11236,N_11594);
nand U12726 (N_12726,N_11121,N_11159);
nor U12727 (N_12727,N_11670,N_11805);
and U12728 (N_12728,N_10690,N_10277);
xnor U12729 (N_12729,N_11656,N_11521);
nor U12730 (N_12730,N_11771,N_11153);
nand U12731 (N_12731,N_10291,N_10840);
nand U12732 (N_12732,N_11874,N_10189);
and U12733 (N_12733,N_10124,N_10176);
or U12734 (N_12734,N_10050,N_11520);
nand U12735 (N_12735,N_11816,N_11277);
nand U12736 (N_12736,N_11155,N_10112);
xnor U12737 (N_12737,N_11001,N_10219);
xor U12738 (N_12738,N_10981,N_10379);
xnor U12739 (N_12739,N_11111,N_10415);
and U12740 (N_12740,N_10309,N_10660);
xor U12741 (N_12741,N_10202,N_10138);
xnor U12742 (N_12742,N_11570,N_10984);
or U12743 (N_12743,N_10588,N_11037);
nand U12744 (N_12744,N_11664,N_10573);
nor U12745 (N_12745,N_11288,N_11956);
nand U12746 (N_12746,N_11162,N_11715);
and U12747 (N_12747,N_10734,N_10639);
and U12748 (N_12748,N_11931,N_10700);
xnor U12749 (N_12749,N_10873,N_11461);
nand U12750 (N_12750,N_11840,N_11821);
nor U12751 (N_12751,N_11562,N_11336);
and U12752 (N_12752,N_11504,N_10797);
nand U12753 (N_12753,N_11429,N_11989);
nor U12754 (N_12754,N_11509,N_10550);
xor U12755 (N_12755,N_11777,N_11858);
nor U12756 (N_12756,N_10979,N_11180);
nor U12757 (N_12757,N_11833,N_11915);
nor U12758 (N_12758,N_11473,N_11612);
nand U12759 (N_12759,N_10747,N_10545);
nor U12760 (N_12760,N_10651,N_10192);
xor U12761 (N_12761,N_10664,N_10693);
nand U12762 (N_12762,N_10539,N_10515);
nand U12763 (N_12763,N_10229,N_10828);
or U12764 (N_12764,N_11785,N_11677);
nor U12765 (N_12765,N_10104,N_11939);
xor U12766 (N_12766,N_11783,N_10151);
nand U12767 (N_12767,N_10953,N_10284);
nand U12768 (N_12768,N_10335,N_10264);
nand U12769 (N_12769,N_11779,N_10083);
and U12770 (N_12770,N_11983,N_10375);
or U12771 (N_12771,N_11057,N_11119);
xnor U12772 (N_12772,N_10091,N_11781);
or U12773 (N_12773,N_10100,N_10348);
or U12774 (N_12774,N_11718,N_11247);
and U12775 (N_12775,N_11490,N_11775);
nand U12776 (N_12776,N_11587,N_11687);
and U12777 (N_12777,N_10576,N_11148);
xor U12778 (N_12778,N_11563,N_11819);
nor U12779 (N_12779,N_10505,N_11749);
or U12780 (N_12780,N_10098,N_10743);
and U12781 (N_12781,N_10529,N_10184);
xnor U12782 (N_12782,N_10430,N_10919);
and U12783 (N_12783,N_11149,N_11572);
nor U12784 (N_12784,N_11078,N_11759);
xor U12785 (N_12785,N_10113,N_10061);
nand U12786 (N_12786,N_11385,N_10243);
and U12787 (N_12787,N_11973,N_11801);
and U12788 (N_12788,N_10935,N_10346);
nor U12789 (N_12789,N_10634,N_10527);
and U12790 (N_12790,N_11850,N_11968);
xnor U12791 (N_12791,N_10156,N_11660);
nand U12792 (N_12792,N_10178,N_11359);
and U12793 (N_12793,N_10075,N_11007);
nor U12794 (N_12794,N_10198,N_11731);
or U12795 (N_12795,N_11439,N_11826);
or U12796 (N_12796,N_10557,N_10985);
xnor U12797 (N_12797,N_10247,N_10640);
and U12798 (N_12798,N_11880,N_10534);
nand U12799 (N_12799,N_10845,N_10194);
nor U12800 (N_12800,N_10373,N_10137);
or U12801 (N_12801,N_11531,N_10841);
and U12802 (N_12802,N_11503,N_10993);
or U12803 (N_12803,N_11306,N_11064);
nand U12804 (N_12804,N_10761,N_11025);
nor U12805 (N_12805,N_10263,N_11038);
xor U12806 (N_12806,N_10081,N_11324);
nor U12807 (N_12807,N_10274,N_11910);
nor U12808 (N_12808,N_11558,N_11029);
xnor U12809 (N_12809,N_10997,N_11986);
nand U12810 (N_12810,N_10751,N_10491);
xor U12811 (N_12811,N_10685,N_11219);
and U12812 (N_12812,N_10627,N_10592);
nand U12813 (N_12813,N_10523,N_11018);
or U12814 (N_12814,N_11976,N_11302);
nand U12815 (N_12815,N_10554,N_11352);
nand U12816 (N_12816,N_10478,N_11719);
nand U12817 (N_12817,N_10434,N_10556);
xor U12818 (N_12818,N_10630,N_10875);
nand U12819 (N_12819,N_11444,N_11372);
nand U12820 (N_12820,N_10901,N_10766);
and U12821 (N_12821,N_11406,N_11003);
nand U12822 (N_12822,N_11200,N_11625);
nor U12823 (N_12823,N_10858,N_11669);
and U12824 (N_12824,N_11584,N_10974);
nand U12825 (N_12825,N_10962,N_11077);
or U12826 (N_12826,N_11544,N_11249);
xor U12827 (N_12827,N_10735,N_10031);
and U12828 (N_12828,N_10662,N_10044);
nor U12829 (N_12829,N_10016,N_10939);
xnor U12830 (N_12830,N_11186,N_11807);
nor U12831 (N_12831,N_11299,N_10389);
nand U12832 (N_12832,N_11725,N_11160);
xnor U12833 (N_12833,N_10111,N_11540);
or U12834 (N_12834,N_10679,N_10248);
nand U12835 (N_12835,N_11179,N_11492);
or U12836 (N_12836,N_11085,N_11260);
nor U12837 (N_12837,N_11678,N_11213);
and U12838 (N_12838,N_11310,N_11737);
and U12839 (N_12839,N_10909,N_10298);
and U12840 (N_12840,N_10362,N_10782);
and U12841 (N_12841,N_10587,N_11512);
nor U12842 (N_12842,N_10730,N_10063);
xor U12843 (N_12843,N_11575,N_10617);
xor U12844 (N_12844,N_11662,N_10920);
nand U12845 (N_12845,N_10253,N_11884);
nand U12846 (N_12846,N_10163,N_10439);
and U12847 (N_12847,N_10686,N_10241);
xnor U12848 (N_12848,N_10474,N_11941);
xor U12849 (N_12849,N_11361,N_11666);
and U12850 (N_12850,N_10207,N_11511);
and U12851 (N_12851,N_11532,N_10570);
nand U12852 (N_12852,N_10680,N_10956);
or U12853 (N_12853,N_11536,N_10269);
or U12854 (N_12854,N_11486,N_10934);
or U12855 (N_12855,N_10740,N_10334);
xor U12856 (N_12856,N_11524,N_11109);
nor U12857 (N_12857,N_10500,N_10376);
nor U12858 (N_12858,N_11082,N_11095);
nor U12859 (N_12859,N_10457,N_11855);
nor U12860 (N_12860,N_11835,N_11753);
xnor U12861 (N_12861,N_11188,N_11143);
nand U12862 (N_12862,N_10517,N_10941);
nor U12863 (N_12863,N_10616,N_10419);
nor U12864 (N_12864,N_11817,N_10737);
xnor U12865 (N_12865,N_11827,N_11108);
and U12866 (N_12866,N_10181,N_11716);
or U12867 (N_12867,N_11653,N_11132);
or U12868 (N_12868,N_11866,N_10808);
or U12869 (N_12869,N_11271,N_11290);
xnor U12870 (N_12870,N_11868,N_10619);
nand U12871 (N_12871,N_10745,N_10122);
and U12872 (N_12872,N_11204,N_11270);
xor U12873 (N_12873,N_11387,N_11649);
nor U12874 (N_12874,N_11769,N_10597);
and U12875 (N_12875,N_11663,N_11515);
nor U12876 (N_12876,N_10388,N_10658);
and U12877 (N_12877,N_10395,N_11865);
xor U12878 (N_12878,N_10564,N_10945);
xor U12879 (N_12879,N_11895,N_11809);
nor U12880 (N_12880,N_10860,N_10036);
xor U12881 (N_12881,N_10599,N_11496);
xnor U12882 (N_12882,N_10625,N_11890);
and U12883 (N_12883,N_10397,N_11088);
and U12884 (N_12884,N_11118,N_11881);
nor U12885 (N_12885,N_10488,N_10867);
xnor U12886 (N_12886,N_10731,N_10609);
and U12887 (N_12887,N_11478,N_10244);
or U12888 (N_12888,N_10359,N_11235);
nand U12889 (N_12889,N_11519,N_10603);
or U12890 (N_12890,N_10222,N_11991);
or U12891 (N_12891,N_11774,N_10133);
xor U12892 (N_12892,N_11158,N_11924);
nor U12893 (N_12893,N_10483,N_10870);
or U12894 (N_12894,N_10341,N_10949);
or U12895 (N_12895,N_11327,N_10874);
xor U12896 (N_12896,N_11225,N_11808);
nor U12897 (N_12897,N_11035,N_11773);
and U12898 (N_12898,N_10011,N_10663);
xor U12899 (N_12899,N_11929,N_10837);
nand U12900 (N_12900,N_10915,N_10739);
or U12901 (N_12901,N_11208,N_11443);
xor U12902 (N_12902,N_10722,N_11566);
and U12903 (N_12903,N_11609,N_10924);
or U12904 (N_12904,N_11870,N_10481);
or U12905 (N_12905,N_11757,N_11707);
or U12906 (N_12906,N_10615,N_11548);
nand U12907 (N_12907,N_11883,N_10666);
or U12908 (N_12908,N_10575,N_11051);
or U12909 (N_12909,N_11112,N_10496);
and U12910 (N_12910,N_10604,N_10718);
xnor U12911 (N_12911,N_11844,N_11714);
and U12912 (N_12912,N_11128,N_10948);
nor U12913 (N_12913,N_10043,N_10048);
nor U12914 (N_12914,N_10077,N_11658);
nor U12915 (N_12915,N_11462,N_10249);
nand U12916 (N_12916,N_11526,N_10045);
nor U12917 (N_12917,N_11101,N_11596);
nor U12918 (N_12918,N_10621,N_11030);
nand U12919 (N_12919,N_10290,N_11423);
or U12920 (N_12920,N_10601,N_10268);
or U12921 (N_12921,N_10688,N_11019);
and U12922 (N_12922,N_10719,N_11489);
and U12923 (N_12923,N_11070,N_10190);
xor U12924 (N_12924,N_10329,N_10884);
nand U12925 (N_12925,N_11904,N_11639);
and U12926 (N_12926,N_10147,N_10270);
and U12927 (N_12927,N_11414,N_10998);
xor U12928 (N_12928,N_11556,N_10068);
xor U12929 (N_12929,N_10149,N_10611);
nand U12930 (N_12930,N_10070,N_10843);
nand U12931 (N_12931,N_11008,N_11296);
nor U12932 (N_12932,N_11420,N_11351);
and U12933 (N_12933,N_10988,N_10485);
or U12934 (N_12934,N_10166,N_11588);
xor U12935 (N_12935,N_11651,N_11613);
nor U12936 (N_12936,N_11040,N_10753);
xor U12937 (N_12937,N_11315,N_10493);
and U12938 (N_12938,N_10513,N_11391);
or U12939 (N_12939,N_10560,N_11096);
nand U12940 (N_12940,N_10980,N_10235);
nor U12941 (N_12941,N_10890,N_10802);
or U12942 (N_12942,N_11141,N_11386);
xor U12943 (N_12943,N_11733,N_10706);
nor U12944 (N_12944,N_11534,N_10665);
xor U12945 (N_12945,N_10898,N_11726);
xnor U12946 (N_12946,N_11137,N_10912);
nand U12947 (N_12947,N_10454,N_11539);
and U12948 (N_12948,N_10742,N_11424);
nor U12949 (N_12949,N_10995,N_11867);
nand U12950 (N_12950,N_11582,N_10654);
xnor U12951 (N_12951,N_10776,N_10394);
and U12952 (N_12952,N_10675,N_11491);
and U12953 (N_12953,N_11672,N_10637);
and U12954 (N_12954,N_11601,N_11457);
nand U12955 (N_12955,N_11166,N_11232);
nand U12956 (N_12956,N_11960,N_11693);
nor U12957 (N_12957,N_10532,N_10652);
nand U12958 (N_12958,N_11206,N_11115);
or U12959 (N_12959,N_10130,N_11326);
xnor U12960 (N_12960,N_11172,N_10369);
or U12961 (N_12961,N_10392,N_11622);
or U12962 (N_12962,N_10310,N_11107);
and U12963 (N_12963,N_11308,N_11985);
nor U12964 (N_12964,N_10504,N_11655);
and U12965 (N_12965,N_10876,N_11199);
or U12966 (N_12966,N_10852,N_10502);
nand U12967 (N_12967,N_11620,N_10221);
nand U12968 (N_12968,N_11592,N_11972);
or U12969 (N_12969,N_11680,N_11279);
nand U12970 (N_12970,N_11446,N_10429);
nand U12971 (N_12971,N_10572,N_10057);
nor U12972 (N_12972,N_10558,N_10364);
and U12973 (N_12973,N_10435,N_10610);
or U12974 (N_12974,N_10062,N_11015);
nor U12975 (N_12975,N_10552,N_10360);
or U12976 (N_12976,N_11702,N_11281);
nand U12977 (N_12977,N_11010,N_10789);
and U12978 (N_12978,N_10605,N_10765);
xor U12979 (N_12979,N_11795,N_10421);
nor U12980 (N_12980,N_10208,N_10954);
or U12981 (N_12981,N_11011,N_11899);
or U12982 (N_12982,N_11756,N_10210);
xnor U12983 (N_12983,N_10215,N_10911);
nor U12984 (N_12984,N_10796,N_10593);
nand U12985 (N_12985,N_10568,N_10618);
or U12986 (N_12986,N_11133,N_11268);
nor U12987 (N_12987,N_11465,N_11873);
nand U12988 (N_12988,N_10626,N_10017);
nand U12989 (N_12989,N_10536,N_10108);
and U12990 (N_12990,N_10033,N_10519);
nand U12991 (N_12991,N_10003,N_11198);
nand U12992 (N_12992,N_10661,N_11039);
xor U12993 (N_12993,N_11803,N_11630);
and U12994 (N_12994,N_11699,N_10608);
xnor U12995 (N_12995,N_11966,N_10020);
or U12996 (N_12996,N_11642,N_11525);
and U12997 (N_12997,N_10281,N_11626);
and U12998 (N_12998,N_11585,N_10384);
nand U12999 (N_12999,N_11618,N_10308);
or U13000 (N_13000,N_10873,N_11906);
nand U13001 (N_13001,N_10430,N_10536);
xor U13002 (N_13002,N_11237,N_10657);
xnor U13003 (N_13003,N_11973,N_10308);
or U13004 (N_13004,N_10080,N_10593);
nand U13005 (N_13005,N_10686,N_10883);
and U13006 (N_13006,N_10099,N_11398);
nor U13007 (N_13007,N_11170,N_11767);
xnor U13008 (N_13008,N_11537,N_10686);
nand U13009 (N_13009,N_11608,N_10474);
and U13010 (N_13010,N_10355,N_11505);
nand U13011 (N_13011,N_11355,N_10107);
nand U13012 (N_13012,N_10141,N_11466);
xnor U13013 (N_13013,N_10619,N_10416);
xor U13014 (N_13014,N_11418,N_10690);
nand U13015 (N_13015,N_11485,N_10233);
xor U13016 (N_13016,N_11190,N_10432);
nor U13017 (N_13017,N_10974,N_10000);
xnor U13018 (N_13018,N_10276,N_10256);
xnor U13019 (N_13019,N_11736,N_10404);
and U13020 (N_13020,N_10123,N_10764);
nor U13021 (N_13021,N_11638,N_11129);
nor U13022 (N_13022,N_11108,N_11482);
xnor U13023 (N_13023,N_11089,N_10933);
nand U13024 (N_13024,N_11575,N_11989);
nand U13025 (N_13025,N_11403,N_11173);
xor U13026 (N_13026,N_10314,N_10352);
nor U13027 (N_13027,N_11149,N_11950);
or U13028 (N_13028,N_11608,N_10435);
xnor U13029 (N_13029,N_11334,N_11501);
and U13030 (N_13030,N_11837,N_10708);
nor U13031 (N_13031,N_11555,N_10660);
nand U13032 (N_13032,N_10519,N_10715);
nor U13033 (N_13033,N_11971,N_11921);
nor U13034 (N_13034,N_11911,N_10863);
or U13035 (N_13035,N_10093,N_11287);
nand U13036 (N_13036,N_11666,N_11068);
xnor U13037 (N_13037,N_10727,N_11762);
nand U13038 (N_13038,N_11034,N_10018);
and U13039 (N_13039,N_11182,N_10264);
xor U13040 (N_13040,N_11571,N_11948);
nor U13041 (N_13041,N_10453,N_10908);
or U13042 (N_13042,N_10552,N_11016);
nor U13043 (N_13043,N_11832,N_10527);
nand U13044 (N_13044,N_11628,N_11776);
xnor U13045 (N_13045,N_10870,N_11364);
nor U13046 (N_13046,N_10495,N_10918);
xor U13047 (N_13047,N_10322,N_10496);
or U13048 (N_13048,N_11853,N_11239);
nor U13049 (N_13049,N_10468,N_11658);
or U13050 (N_13050,N_10222,N_11622);
nand U13051 (N_13051,N_10700,N_11705);
and U13052 (N_13052,N_10550,N_11563);
nand U13053 (N_13053,N_10120,N_11491);
and U13054 (N_13054,N_11514,N_11074);
or U13055 (N_13055,N_10674,N_11031);
and U13056 (N_13056,N_10757,N_10493);
nor U13057 (N_13057,N_10456,N_11713);
xnor U13058 (N_13058,N_11850,N_11407);
xor U13059 (N_13059,N_10679,N_10041);
nor U13060 (N_13060,N_10613,N_10367);
xnor U13061 (N_13061,N_10968,N_11384);
nor U13062 (N_13062,N_10667,N_11461);
or U13063 (N_13063,N_11638,N_10586);
and U13064 (N_13064,N_10207,N_10894);
or U13065 (N_13065,N_10258,N_11519);
xnor U13066 (N_13066,N_11527,N_10822);
xnor U13067 (N_13067,N_10029,N_10049);
nand U13068 (N_13068,N_11965,N_11075);
and U13069 (N_13069,N_10554,N_10750);
nand U13070 (N_13070,N_10241,N_11503);
nor U13071 (N_13071,N_11947,N_11715);
nand U13072 (N_13072,N_10472,N_11662);
nand U13073 (N_13073,N_11719,N_10527);
nand U13074 (N_13074,N_10143,N_10331);
nor U13075 (N_13075,N_11416,N_10242);
or U13076 (N_13076,N_10051,N_10347);
xnor U13077 (N_13077,N_10214,N_11507);
nand U13078 (N_13078,N_11325,N_10600);
and U13079 (N_13079,N_11333,N_11183);
or U13080 (N_13080,N_10997,N_10826);
xnor U13081 (N_13081,N_11072,N_11960);
or U13082 (N_13082,N_11681,N_10414);
or U13083 (N_13083,N_10510,N_10177);
nand U13084 (N_13084,N_10549,N_10369);
or U13085 (N_13085,N_10996,N_11756);
xor U13086 (N_13086,N_10415,N_10062);
nor U13087 (N_13087,N_10994,N_11434);
and U13088 (N_13088,N_11576,N_11359);
nand U13089 (N_13089,N_11154,N_10917);
nand U13090 (N_13090,N_11603,N_10043);
nand U13091 (N_13091,N_10132,N_10384);
xor U13092 (N_13092,N_10664,N_10733);
xnor U13093 (N_13093,N_10288,N_10996);
nor U13094 (N_13094,N_10818,N_10069);
nor U13095 (N_13095,N_11169,N_10763);
or U13096 (N_13096,N_10924,N_11199);
and U13097 (N_13097,N_10563,N_11433);
nor U13098 (N_13098,N_10734,N_10153);
nor U13099 (N_13099,N_10666,N_11968);
nor U13100 (N_13100,N_11611,N_10513);
and U13101 (N_13101,N_10186,N_11781);
nor U13102 (N_13102,N_11075,N_10739);
or U13103 (N_13103,N_10111,N_11078);
nor U13104 (N_13104,N_10805,N_11790);
or U13105 (N_13105,N_11550,N_10614);
and U13106 (N_13106,N_10918,N_11922);
xor U13107 (N_13107,N_11764,N_11583);
xnor U13108 (N_13108,N_11425,N_11986);
nor U13109 (N_13109,N_11662,N_11897);
or U13110 (N_13110,N_10121,N_10917);
and U13111 (N_13111,N_10672,N_10576);
xnor U13112 (N_13112,N_11400,N_10627);
nor U13113 (N_13113,N_10221,N_11641);
nor U13114 (N_13114,N_11248,N_11256);
nand U13115 (N_13115,N_10269,N_10582);
or U13116 (N_13116,N_11132,N_11231);
and U13117 (N_13117,N_10964,N_11099);
or U13118 (N_13118,N_10683,N_11830);
xnor U13119 (N_13119,N_11927,N_10756);
xnor U13120 (N_13120,N_10404,N_10126);
xnor U13121 (N_13121,N_10057,N_10299);
nor U13122 (N_13122,N_10994,N_10809);
xnor U13123 (N_13123,N_11173,N_11766);
and U13124 (N_13124,N_10367,N_10418);
or U13125 (N_13125,N_10832,N_11568);
or U13126 (N_13126,N_10390,N_11924);
or U13127 (N_13127,N_10979,N_10423);
and U13128 (N_13128,N_10683,N_10194);
nand U13129 (N_13129,N_10765,N_11798);
nand U13130 (N_13130,N_10624,N_11281);
or U13131 (N_13131,N_10258,N_10360);
or U13132 (N_13132,N_10624,N_11913);
xor U13133 (N_13133,N_10164,N_11924);
xnor U13134 (N_13134,N_10134,N_10512);
nor U13135 (N_13135,N_10793,N_11506);
xor U13136 (N_13136,N_11642,N_10331);
xor U13137 (N_13137,N_10898,N_10688);
nand U13138 (N_13138,N_11473,N_10625);
xor U13139 (N_13139,N_10575,N_11264);
xnor U13140 (N_13140,N_11251,N_10163);
nor U13141 (N_13141,N_11555,N_11410);
nor U13142 (N_13142,N_11343,N_11950);
nand U13143 (N_13143,N_10288,N_11135);
nor U13144 (N_13144,N_11170,N_10034);
xor U13145 (N_13145,N_10012,N_10380);
or U13146 (N_13146,N_10135,N_11235);
or U13147 (N_13147,N_11866,N_11958);
nor U13148 (N_13148,N_10517,N_11571);
xor U13149 (N_13149,N_10520,N_10043);
nor U13150 (N_13150,N_10682,N_10693);
xor U13151 (N_13151,N_10196,N_11316);
or U13152 (N_13152,N_11785,N_11559);
nand U13153 (N_13153,N_10070,N_10847);
and U13154 (N_13154,N_10550,N_11923);
nor U13155 (N_13155,N_11942,N_11013);
nor U13156 (N_13156,N_10225,N_11952);
nand U13157 (N_13157,N_11191,N_11857);
nand U13158 (N_13158,N_10898,N_10199);
or U13159 (N_13159,N_11849,N_10150);
xor U13160 (N_13160,N_10417,N_11921);
xor U13161 (N_13161,N_11946,N_11284);
or U13162 (N_13162,N_11888,N_10107);
xnor U13163 (N_13163,N_11975,N_10354);
and U13164 (N_13164,N_11775,N_11239);
or U13165 (N_13165,N_10407,N_10599);
xnor U13166 (N_13166,N_11491,N_10943);
or U13167 (N_13167,N_11451,N_10386);
nor U13168 (N_13168,N_11482,N_11647);
and U13169 (N_13169,N_10677,N_10054);
nor U13170 (N_13170,N_10778,N_11221);
xor U13171 (N_13171,N_11406,N_11832);
or U13172 (N_13172,N_10771,N_10334);
and U13173 (N_13173,N_10789,N_10968);
nor U13174 (N_13174,N_10867,N_11238);
xnor U13175 (N_13175,N_10740,N_11723);
or U13176 (N_13176,N_11628,N_11764);
nand U13177 (N_13177,N_11900,N_11677);
or U13178 (N_13178,N_11501,N_11632);
nand U13179 (N_13179,N_11962,N_11546);
xnor U13180 (N_13180,N_11808,N_10567);
and U13181 (N_13181,N_10547,N_11056);
nor U13182 (N_13182,N_10505,N_10412);
or U13183 (N_13183,N_10096,N_11670);
or U13184 (N_13184,N_10178,N_11728);
xnor U13185 (N_13185,N_11712,N_11980);
and U13186 (N_13186,N_10407,N_10587);
or U13187 (N_13187,N_11457,N_11050);
xor U13188 (N_13188,N_10425,N_11389);
nand U13189 (N_13189,N_10687,N_10334);
nor U13190 (N_13190,N_11256,N_10194);
nand U13191 (N_13191,N_11124,N_11887);
nand U13192 (N_13192,N_11681,N_11821);
nand U13193 (N_13193,N_10533,N_11111);
and U13194 (N_13194,N_10596,N_10714);
and U13195 (N_13195,N_11958,N_10263);
nand U13196 (N_13196,N_10310,N_10820);
or U13197 (N_13197,N_10589,N_10829);
nand U13198 (N_13198,N_10887,N_10327);
nand U13199 (N_13199,N_10840,N_10256);
nand U13200 (N_13200,N_11216,N_10496);
xnor U13201 (N_13201,N_11020,N_11213);
and U13202 (N_13202,N_10990,N_10328);
nor U13203 (N_13203,N_10439,N_10471);
and U13204 (N_13204,N_10943,N_10825);
nand U13205 (N_13205,N_11658,N_10381);
nor U13206 (N_13206,N_10389,N_10363);
xor U13207 (N_13207,N_10562,N_11473);
or U13208 (N_13208,N_10812,N_10024);
nand U13209 (N_13209,N_10701,N_10982);
or U13210 (N_13210,N_11784,N_10798);
xor U13211 (N_13211,N_11638,N_10688);
nand U13212 (N_13212,N_11220,N_10424);
xnor U13213 (N_13213,N_11862,N_10269);
nor U13214 (N_13214,N_11466,N_11044);
and U13215 (N_13215,N_11593,N_11944);
and U13216 (N_13216,N_10348,N_10478);
xor U13217 (N_13217,N_10747,N_11212);
nand U13218 (N_13218,N_10764,N_10099);
nor U13219 (N_13219,N_10356,N_11734);
nor U13220 (N_13220,N_10610,N_10163);
nor U13221 (N_13221,N_11779,N_11597);
or U13222 (N_13222,N_11853,N_10624);
nand U13223 (N_13223,N_10740,N_11746);
nor U13224 (N_13224,N_10381,N_10726);
and U13225 (N_13225,N_10856,N_11739);
and U13226 (N_13226,N_11848,N_11221);
and U13227 (N_13227,N_10096,N_10047);
or U13228 (N_13228,N_10012,N_11651);
xor U13229 (N_13229,N_11969,N_10560);
and U13230 (N_13230,N_11437,N_10930);
and U13231 (N_13231,N_10129,N_10131);
xnor U13232 (N_13232,N_11612,N_11462);
and U13233 (N_13233,N_11833,N_11505);
and U13234 (N_13234,N_11456,N_10983);
nand U13235 (N_13235,N_10459,N_10173);
nand U13236 (N_13236,N_10071,N_10972);
or U13237 (N_13237,N_11687,N_10820);
or U13238 (N_13238,N_10826,N_10077);
xor U13239 (N_13239,N_10299,N_10655);
or U13240 (N_13240,N_11773,N_11870);
nor U13241 (N_13241,N_11679,N_10242);
nor U13242 (N_13242,N_11044,N_10398);
or U13243 (N_13243,N_10935,N_11436);
xnor U13244 (N_13244,N_11303,N_10766);
and U13245 (N_13245,N_10016,N_10295);
nor U13246 (N_13246,N_11693,N_10473);
and U13247 (N_13247,N_11254,N_10647);
xnor U13248 (N_13248,N_10680,N_10987);
nor U13249 (N_13249,N_10264,N_10163);
nand U13250 (N_13250,N_11637,N_11263);
and U13251 (N_13251,N_11696,N_11863);
xor U13252 (N_13252,N_10897,N_10308);
xor U13253 (N_13253,N_10220,N_10877);
nor U13254 (N_13254,N_11899,N_11321);
and U13255 (N_13255,N_11462,N_10018);
nor U13256 (N_13256,N_10945,N_11567);
nor U13257 (N_13257,N_11325,N_10592);
nand U13258 (N_13258,N_10801,N_10742);
nor U13259 (N_13259,N_10851,N_10114);
nand U13260 (N_13260,N_11726,N_11429);
nor U13261 (N_13261,N_10510,N_11362);
and U13262 (N_13262,N_10292,N_10675);
or U13263 (N_13263,N_10444,N_11167);
and U13264 (N_13264,N_10512,N_11802);
and U13265 (N_13265,N_10527,N_11119);
xor U13266 (N_13266,N_11574,N_11538);
or U13267 (N_13267,N_11982,N_11842);
nor U13268 (N_13268,N_10931,N_11650);
nand U13269 (N_13269,N_10247,N_11407);
nor U13270 (N_13270,N_10192,N_10636);
and U13271 (N_13271,N_10127,N_10784);
or U13272 (N_13272,N_10592,N_10147);
nand U13273 (N_13273,N_11570,N_10353);
nand U13274 (N_13274,N_10418,N_10215);
and U13275 (N_13275,N_11989,N_11041);
nand U13276 (N_13276,N_11511,N_10088);
nand U13277 (N_13277,N_11812,N_10847);
and U13278 (N_13278,N_10287,N_11253);
and U13279 (N_13279,N_10995,N_11064);
xnor U13280 (N_13280,N_10211,N_10394);
xnor U13281 (N_13281,N_10600,N_11575);
and U13282 (N_13282,N_11622,N_10225);
xnor U13283 (N_13283,N_11923,N_10880);
or U13284 (N_13284,N_11778,N_10573);
and U13285 (N_13285,N_11898,N_10593);
nor U13286 (N_13286,N_10842,N_11049);
or U13287 (N_13287,N_11196,N_11652);
and U13288 (N_13288,N_10808,N_10651);
nor U13289 (N_13289,N_11401,N_10368);
xnor U13290 (N_13290,N_11753,N_10173);
xor U13291 (N_13291,N_10891,N_10614);
nor U13292 (N_13292,N_11508,N_10238);
nor U13293 (N_13293,N_10378,N_10272);
and U13294 (N_13294,N_11436,N_10597);
or U13295 (N_13295,N_11419,N_10174);
nor U13296 (N_13296,N_10623,N_11621);
nor U13297 (N_13297,N_11956,N_10599);
nor U13298 (N_13298,N_11307,N_10665);
or U13299 (N_13299,N_10339,N_10947);
and U13300 (N_13300,N_11051,N_10365);
nor U13301 (N_13301,N_11586,N_10880);
xor U13302 (N_13302,N_10580,N_10118);
nor U13303 (N_13303,N_11244,N_11592);
and U13304 (N_13304,N_10537,N_11366);
and U13305 (N_13305,N_11949,N_11618);
nor U13306 (N_13306,N_11786,N_11336);
xnor U13307 (N_13307,N_10051,N_11412);
xnor U13308 (N_13308,N_11602,N_11119);
nor U13309 (N_13309,N_10262,N_11971);
and U13310 (N_13310,N_11545,N_11343);
nor U13311 (N_13311,N_11092,N_11283);
or U13312 (N_13312,N_11500,N_11580);
xnor U13313 (N_13313,N_10431,N_10871);
and U13314 (N_13314,N_10519,N_10522);
or U13315 (N_13315,N_10560,N_10405);
nor U13316 (N_13316,N_10624,N_10582);
xor U13317 (N_13317,N_10996,N_10465);
nand U13318 (N_13318,N_11878,N_11658);
nand U13319 (N_13319,N_11887,N_11475);
nor U13320 (N_13320,N_11248,N_10444);
or U13321 (N_13321,N_10875,N_11142);
nor U13322 (N_13322,N_10107,N_11791);
or U13323 (N_13323,N_10759,N_10370);
and U13324 (N_13324,N_10875,N_11276);
xor U13325 (N_13325,N_10105,N_11434);
nor U13326 (N_13326,N_11220,N_10490);
xnor U13327 (N_13327,N_11776,N_10207);
or U13328 (N_13328,N_11148,N_10269);
nor U13329 (N_13329,N_11981,N_10365);
and U13330 (N_13330,N_11308,N_10040);
nor U13331 (N_13331,N_10401,N_10281);
or U13332 (N_13332,N_11216,N_10770);
or U13333 (N_13333,N_10838,N_10635);
xnor U13334 (N_13334,N_10197,N_10088);
or U13335 (N_13335,N_11925,N_10982);
nor U13336 (N_13336,N_11115,N_10958);
xor U13337 (N_13337,N_11629,N_11980);
nand U13338 (N_13338,N_10691,N_11990);
xor U13339 (N_13339,N_10708,N_11208);
or U13340 (N_13340,N_11525,N_10515);
nand U13341 (N_13341,N_11590,N_10891);
and U13342 (N_13342,N_10555,N_11139);
nand U13343 (N_13343,N_11030,N_11239);
and U13344 (N_13344,N_10945,N_10758);
xor U13345 (N_13345,N_11382,N_10963);
nor U13346 (N_13346,N_11190,N_10905);
and U13347 (N_13347,N_10635,N_10931);
nor U13348 (N_13348,N_11164,N_10597);
and U13349 (N_13349,N_11237,N_11851);
and U13350 (N_13350,N_10426,N_10614);
nand U13351 (N_13351,N_10138,N_10495);
nand U13352 (N_13352,N_11819,N_10996);
nor U13353 (N_13353,N_10681,N_10648);
nand U13354 (N_13354,N_10823,N_10963);
nor U13355 (N_13355,N_11836,N_10793);
and U13356 (N_13356,N_11744,N_10050);
xor U13357 (N_13357,N_11642,N_11448);
nor U13358 (N_13358,N_10807,N_10675);
and U13359 (N_13359,N_11237,N_10926);
nor U13360 (N_13360,N_11077,N_11776);
xor U13361 (N_13361,N_11251,N_11645);
and U13362 (N_13362,N_10090,N_11543);
xor U13363 (N_13363,N_11327,N_10363);
nand U13364 (N_13364,N_11946,N_10353);
nand U13365 (N_13365,N_10478,N_11166);
xnor U13366 (N_13366,N_11202,N_10391);
or U13367 (N_13367,N_11767,N_11333);
nand U13368 (N_13368,N_11803,N_10357);
and U13369 (N_13369,N_11815,N_10208);
xor U13370 (N_13370,N_11270,N_11450);
nor U13371 (N_13371,N_10127,N_11844);
nand U13372 (N_13372,N_11568,N_10765);
nand U13373 (N_13373,N_10384,N_11924);
and U13374 (N_13374,N_11495,N_10112);
nor U13375 (N_13375,N_11559,N_11662);
nand U13376 (N_13376,N_11194,N_10187);
xnor U13377 (N_13377,N_10974,N_11947);
xnor U13378 (N_13378,N_11837,N_11230);
and U13379 (N_13379,N_11449,N_10757);
or U13380 (N_13380,N_11616,N_10517);
xor U13381 (N_13381,N_11680,N_10242);
xor U13382 (N_13382,N_10201,N_10642);
nor U13383 (N_13383,N_10973,N_10819);
nor U13384 (N_13384,N_11350,N_10461);
nor U13385 (N_13385,N_10092,N_11545);
nor U13386 (N_13386,N_10584,N_11678);
and U13387 (N_13387,N_11093,N_10364);
and U13388 (N_13388,N_10819,N_11978);
or U13389 (N_13389,N_10785,N_10668);
or U13390 (N_13390,N_10633,N_11513);
and U13391 (N_13391,N_10806,N_11396);
and U13392 (N_13392,N_10948,N_10211);
or U13393 (N_13393,N_11440,N_11171);
xor U13394 (N_13394,N_10022,N_10921);
xor U13395 (N_13395,N_11359,N_11343);
xor U13396 (N_13396,N_10213,N_11917);
nand U13397 (N_13397,N_11521,N_11069);
or U13398 (N_13398,N_11360,N_11896);
or U13399 (N_13399,N_11949,N_10312);
and U13400 (N_13400,N_10266,N_11713);
nand U13401 (N_13401,N_10023,N_11974);
nand U13402 (N_13402,N_11721,N_10438);
nand U13403 (N_13403,N_11682,N_11498);
and U13404 (N_13404,N_10093,N_11775);
or U13405 (N_13405,N_10245,N_10325);
xor U13406 (N_13406,N_11810,N_10530);
and U13407 (N_13407,N_11692,N_11569);
nand U13408 (N_13408,N_11836,N_10256);
and U13409 (N_13409,N_10051,N_11248);
nand U13410 (N_13410,N_10192,N_11585);
and U13411 (N_13411,N_10022,N_10843);
nand U13412 (N_13412,N_10796,N_10821);
xnor U13413 (N_13413,N_11495,N_11236);
xnor U13414 (N_13414,N_11117,N_11073);
xor U13415 (N_13415,N_10596,N_11942);
xor U13416 (N_13416,N_11606,N_10985);
nor U13417 (N_13417,N_11109,N_11974);
nor U13418 (N_13418,N_10079,N_11391);
nand U13419 (N_13419,N_10963,N_11142);
and U13420 (N_13420,N_11220,N_11939);
nand U13421 (N_13421,N_10427,N_11558);
and U13422 (N_13422,N_11406,N_11962);
and U13423 (N_13423,N_11695,N_11500);
xor U13424 (N_13424,N_10862,N_11886);
and U13425 (N_13425,N_11819,N_10319);
or U13426 (N_13426,N_11989,N_11490);
or U13427 (N_13427,N_10153,N_10319);
nor U13428 (N_13428,N_10251,N_11599);
nor U13429 (N_13429,N_11151,N_10339);
nand U13430 (N_13430,N_10742,N_10563);
nand U13431 (N_13431,N_10319,N_10307);
and U13432 (N_13432,N_11010,N_10274);
and U13433 (N_13433,N_11896,N_11902);
xnor U13434 (N_13434,N_11171,N_11442);
or U13435 (N_13435,N_11043,N_11117);
nand U13436 (N_13436,N_11091,N_10037);
or U13437 (N_13437,N_11867,N_11886);
nor U13438 (N_13438,N_10984,N_11928);
or U13439 (N_13439,N_11018,N_11685);
or U13440 (N_13440,N_11114,N_10258);
and U13441 (N_13441,N_10639,N_11628);
and U13442 (N_13442,N_11768,N_10705);
or U13443 (N_13443,N_10876,N_11735);
nor U13444 (N_13444,N_11811,N_10125);
nor U13445 (N_13445,N_11704,N_11528);
nand U13446 (N_13446,N_10085,N_10136);
or U13447 (N_13447,N_10846,N_11111);
nand U13448 (N_13448,N_11184,N_10336);
xnor U13449 (N_13449,N_10847,N_11658);
nand U13450 (N_13450,N_11310,N_10631);
nor U13451 (N_13451,N_11132,N_10975);
or U13452 (N_13452,N_11193,N_11308);
nand U13453 (N_13453,N_11126,N_11752);
or U13454 (N_13454,N_10114,N_10261);
and U13455 (N_13455,N_10522,N_10247);
nand U13456 (N_13456,N_10726,N_10657);
nor U13457 (N_13457,N_10431,N_10288);
nand U13458 (N_13458,N_10622,N_10758);
nor U13459 (N_13459,N_11816,N_10354);
and U13460 (N_13460,N_10170,N_11780);
or U13461 (N_13461,N_11406,N_10295);
xor U13462 (N_13462,N_11503,N_10893);
xor U13463 (N_13463,N_11659,N_10601);
and U13464 (N_13464,N_11341,N_10973);
nand U13465 (N_13465,N_10656,N_10055);
nand U13466 (N_13466,N_11955,N_10328);
and U13467 (N_13467,N_11045,N_10876);
and U13468 (N_13468,N_11349,N_11714);
nand U13469 (N_13469,N_11761,N_10226);
nor U13470 (N_13470,N_10929,N_11129);
nor U13471 (N_13471,N_10943,N_11268);
and U13472 (N_13472,N_10574,N_11029);
and U13473 (N_13473,N_10982,N_10402);
nand U13474 (N_13474,N_10387,N_10373);
nand U13475 (N_13475,N_11057,N_10202);
or U13476 (N_13476,N_10424,N_10723);
nor U13477 (N_13477,N_11337,N_11006);
nand U13478 (N_13478,N_11086,N_11348);
nor U13479 (N_13479,N_10538,N_11023);
nor U13480 (N_13480,N_10304,N_11436);
xor U13481 (N_13481,N_10099,N_10312);
and U13482 (N_13482,N_10611,N_10929);
or U13483 (N_13483,N_10847,N_11383);
nand U13484 (N_13484,N_11199,N_11610);
xor U13485 (N_13485,N_11915,N_11438);
or U13486 (N_13486,N_10072,N_11134);
xnor U13487 (N_13487,N_11158,N_10556);
nand U13488 (N_13488,N_11490,N_11113);
or U13489 (N_13489,N_11145,N_10489);
nand U13490 (N_13490,N_11963,N_10876);
and U13491 (N_13491,N_11048,N_10373);
or U13492 (N_13492,N_11432,N_11458);
xnor U13493 (N_13493,N_11356,N_10200);
or U13494 (N_13494,N_11243,N_11933);
nor U13495 (N_13495,N_11455,N_10671);
xor U13496 (N_13496,N_10693,N_10829);
nor U13497 (N_13497,N_11997,N_11014);
nor U13498 (N_13498,N_10233,N_10716);
xnor U13499 (N_13499,N_10431,N_10799);
nand U13500 (N_13500,N_11914,N_10508);
nor U13501 (N_13501,N_10533,N_11583);
xor U13502 (N_13502,N_11999,N_11194);
and U13503 (N_13503,N_10703,N_10170);
nand U13504 (N_13504,N_11935,N_11617);
and U13505 (N_13505,N_11566,N_10224);
nand U13506 (N_13506,N_11023,N_11736);
and U13507 (N_13507,N_10170,N_10053);
nor U13508 (N_13508,N_11864,N_11195);
or U13509 (N_13509,N_10069,N_11665);
and U13510 (N_13510,N_10705,N_10219);
xnor U13511 (N_13511,N_11599,N_11408);
nand U13512 (N_13512,N_10606,N_10989);
or U13513 (N_13513,N_10347,N_10188);
xnor U13514 (N_13514,N_10849,N_10423);
nor U13515 (N_13515,N_11337,N_10965);
nand U13516 (N_13516,N_10288,N_10110);
xnor U13517 (N_13517,N_11531,N_11650);
nand U13518 (N_13518,N_10549,N_11417);
xor U13519 (N_13519,N_11678,N_10957);
xor U13520 (N_13520,N_11982,N_11635);
xor U13521 (N_13521,N_10171,N_10934);
nand U13522 (N_13522,N_11841,N_10030);
nand U13523 (N_13523,N_10964,N_10778);
or U13524 (N_13524,N_11409,N_10810);
or U13525 (N_13525,N_10229,N_11777);
nor U13526 (N_13526,N_11124,N_11784);
or U13527 (N_13527,N_11434,N_11123);
or U13528 (N_13528,N_10589,N_11950);
or U13529 (N_13529,N_11689,N_10480);
xor U13530 (N_13530,N_10953,N_10069);
nor U13531 (N_13531,N_10184,N_10669);
xor U13532 (N_13532,N_10850,N_10766);
xnor U13533 (N_13533,N_11059,N_11494);
or U13534 (N_13534,N_11182,N_10438);
or U13535 (N_13535,N_11606,N_11904);
or U13536 (N_13536,N_10696,N_10377);
nand U13537 (N_13537,N_11596,N_10344);
and U13538 (N_13538,N_11771,N_10610);
and U13539 (N_13539,N_10009,N_11532);
xnor U13540 (N_13540,N_11180,N_11770);
xor U13541 (N_13541,N_11305,N_11968);
nor U13542 (N_13542,N_11544,N_10521);
nor U13543 (N_13543,N_10534,N_11981);
nand U13544 (N_13544,N_10757,N_11600);
nor U13545 (N_13545,N_11794,N_11899);
nor U13546 (N_13546,N_10451,N_11715);
or U13547 (N_13547,N_10431,N_11504);
or U13548 (N_13548,N_11951,N_11176);
or U13549 (N_13549,N_10446,N_10439);
nand U13550 (N_13550,N_10308,N_11251);
xnor U13551 (N_13551,N_11656,N_10521);
or U13552 (N_13552,N_10344,N_10990);
nor U13553 (N_13553,N_11447,N_11571);
and U13554 (N_13554,N_11726,N_10597);
xor U13555 (N_13555,N_10272,N_11557);
nor U13556 (N_13556,N_10028,N_11859);
or U13557 (N_13557,N_11194,N_11842);
nor U13558 (N_13558,N_10797,N_11605);
and U13559 (N_13559,N_10800,N_10230);
xor U13560 (N_13560,N_11536,N_11527);
xor U13561 (N_13561,N_11516,N_11790);
nor U13562 (N_13562,N_10759,N_11377);
nand U13563 (N_13563,N_11632,N_11966);
xor U13564 (N_13564,N_10626,N_11592);
nand U13565 (N_13565,N_10145,N_11144);
xor U13566 (N_13566,N_10141,N_11467);
nor U13567 (N_13567,N_10316,N_11146);
nor U13568 (N_13568,N_10516,N_10692);
nor U13569 (N_13569,N_11238,N_11031);
or U13570 (N_13570,N_10835,N_11314);
xnor U13571 (N_13571,N_11980,N_11748);
and U13572 (N_13572,N_10805,N_10019);
nand U13573 (N_13573,N_10634,N_11976);
nor U13574 (N_13574,N_11542,N_11948);
or U13575 (N_13575,N_10190,N_11754);
xor U13576 (N_13576,N_11441,N_10708);
nand U13577 (N_13577,N_11921,N_10866);
or U13578 (N_13578,N_11425,N_11154);
and U13579 (N_13579,N_10143,N_10237);
nand U13580 (N_13580,N_10414,N_10446);
or U13581 (N_13581,N_10369,N_11637);
nand U13582 (N_13582,N_10003,N_11486);
and U13583 (N_13583,N_11187,N_10464);
nand U13584 (N_13584,N_10163,N_10137);
nand U13585 (N_13585,N_10964,N_11636);
xnor U13586 (N_13586,N_10760,N_11058);
and U13587 (N_13587,N_11532,N_11323);
nor U13588 (N_13588,N_11560,N_11406);
xnor U13589 (N_13589,N_11508,N_10386);
nor U13590 (N_13590,N_10429,N_10102);
and U13591 (N_13591,N_11860,N_11958);
nand U13592 (N_13592,N_10236,N_11491);
and U13593 (N_13593,N_10399,N_11732);
nand U13594 (N_13594,N_10175,N_11278);
xor U13595 (N_13595,N_11202,N_10079);
nor U13596 (N_13596,N_10200,N_10438);
xnor U13597 (N_13597,N_10167,N_11700);
nand U13598 (N_13598,N_11741,N_10529);
nand U13599 (N_13599,N_11031,N_10612);
xnor U13600 (N_13600,N_10382,N_11491);
or U13601 (N_13601,N_11226,N_10273);
nand U13602 (N_13602,N_11672,N_11270);
or U13603 (N_13603,N_11016,N_11834);
nor U13604 (N_13604,N_10152,N_11907);
nand U13605 (N_13605,N_10757,N_11296);
xnor U13606 (N_13606,N_10383,N_10581);
nor U13607 (N_13607,N_11345,N_11215);
nor U13608 (N_13608,N_10421,N_10381);
or U13609 (N_13609,N_11252,N_11795);
and U13610 (N_13610,N_11290,N_10802);
nand U13611 (N_13611,N_11736,N_10582);
and U13612 (N_13612,N_11861,N_11297);
xor U13613 (N_13613,N_11152,N_10897);
and U13614 (N_13614,N_10896,N_10451);
or U13615 (N_13615,N_11904,N_11805);
nand U13616 (N_13616,N_10676,N_11242);
nand U13617 (N_13617,N_10174,N_10386);
nor U13618 (N_13618,N_11898,N_11665);
or U13619 (N_13619,N_10167,N_11090);
xor U13620 (N_13620,N_10437,N_10873);
or U13621 (N_13621,N_11066,N_10059);
nor U13622 (N_13622,N_10477,N_11518);
xnor U13623 (N_13623,N_10913,N_10615);
nor U13624 (N_13624,N_10607,N_11605);
and U13625 (N_13625,N_11908,N_11759);
or U13626 (N_13626,N_11478,N_10503);
nor U13627 (N_13627,N_10216,N_10277);
xor U13628 (N_13628,N_11900,N_11226);
nand U13629 (N_13629,N_10186,N_11101);
nand U13630 (N_13630,N_10174,N_11560);
nand U13631 (N_13631,N_11225,N_10905);
nand U13632 (N_13632,N_11162,N_10999);
nand U13633 (N_13633,N_10744,N_10656);
xnor U13634 (N_13634,N_10694,N_11397);
nor U13635 (N_13635,N_11384,N_10469);
nor U13636 (N_13636,N_11272,N_11408);
nor U13637 (N_13637,N_11553,N_11499);
and U13638 (N_13638,N_10076,N_11791);
nand U13639 (N_13639,N_11210,N_10263);
or U13640 (N_13640,N_10545,N_10632);
nor U13641 (N_13641,N_10220,N_10828);
nor U13642 (N_13642,N_10395,N_10207);
nand U13643 (N_13643,N_11421,N_11761);
nor U13644 (N_13644,N_10500,N_11625);
and U13645 (N_13645,N_10760,N_11397);
nor U13646 (N_13646,N_10241,N_11194);
xnor U13647 (N_13647,N_11081,N_10300);
or U13648 (N_13648,N_10189,N_11822);
xor U13649 (N_13649,N_10922,N_11031);
xor U13650 (N_13650,N_11659,N_10302);
or U13651 (N_13651,N_10125,N_10665);
and U13652 (N_13652,N_10265,N_11429);
or U13653 (N_13653,N_11353,N_11659);
and U13654 (N_13654,N_10574,N_11592);
nand U13655 (N_13655,N_10556,N_11138);
or U13656 (N_13656,N_10760,N_11098);
or U13657 (N_13657,N_11736,N_10515);
or U13658 (N_13658,N_11391,N_10165);
or U13659 (N_13659,N_11185,N_11719);
nand U13660 (N_13660,N_11626,N_10253);
nor U13661 (N_13661,N_11303,N_10858);
and U13662 (N_13662,N_10248,N_10090);
nor U13663 (N_13663,N_11190,N_11907);
and U13664 (N_13664,N_10988,N_10932);
nor U13665 (N_13665,N_10406,N_10450);
nand U13666 (N_13666,N_11436,N_11674);
or U13667 (N_13667,N_10615,N_10252);
or U13668 (N_13668,N_11850,N_10487);
and U13669 (N_13669,N_11988,N_10453);
nor U13670 (N_13670,N_11986,N_10915);
xor U13671 (N_13671,N_11029,N_10158);
nor U13672 (N_13672,N_10033,N_10180);
xor U13673 (N_13673,N_11727,N_10898);
and U13674 (N_13674,N_11119,N_10263);
nand U13675 (N_13675,N_11549,N_10009);
nand U13676 (N_13676,N_11827,N_10521);
xnor U13677 (N_13677,N_11360,N_11969);
nor U13678 (N_13678,N_10385,N_11906);
and U13679 (N_13679,N_10930,N_11218);
xor U13680 (N_13680,N_11838,N_11903);
xnor U13681 (N_13681,N_11237,N_10350);
xnor U13682 (N_13682,N_11972,N_11470);
nand U13683 (N_13683,N_11851,N_11988);
and U13684 (N_13684,N_11190,N_11372);
or U13685 (N_13685,N_10634,N_11933);
xor U13686 (N_13686,N_11887,N_10769);
and U13687 (N_13687,N_10059,N_10731);
nor U13688 (N_13688,N_11788,N_11188);
or U13689 (N_13689,N_10238,N_11613);
and U13690 (N_13690,N_10903,N_11080);
xor U13691 (N_13691,N_11125,N_11457);
nor U13692 (N_13692,N_10855,N_11558);
nand U13693 (N_13693,N_11352,N_10779);
or U13694 (N_13694,N_10179,N_11719);
or U13695 (N_13695,N_11193,N_11939);
xnor U13696 (N_13696,N_10903,N_10364);
or U13697 (N_13697,N_11492,N_11791);
nand U13698 (N_13698,N_11180,N_10871);
xor U13699 (N_13699,N_11715,N_10531);
nor U13700 (N_13700,N_10647,N_10841);
or U13701 (N_13701,N_11183,N_11509);
nand U13702 (N_13702,N_10460,N_11786);
nor U13703 (N_13703,N_10429,N_11871);
nor U13704 (N_13704,N_10550,N_10326);
nor U13705 (N_13705,N_10076,N_10482);
xnor U13706 (N_13706,N_10348,N_10483);
nor U13707 (N_13707,N_11169,N_10943);
nor U13708 (N_13708,N_10346,N_10276);
nand U13709 (N_13709,N_11868,N_10858);
and U13710 (N_13710,N_11720,N_10407);
or U13711 (N_13711,N_11824,N_11766);
xnor U13712 (N_13712,N_11704,N_11039);
xnor U13713 (N_13713,N_11000,N_10689);
nor U13714 (N_13714,N_10040,N_11955);
xnor U13715 (N_13715,N_11955,N_10613);
xor U13716 (N_13716,N_11029,N_11682);
nor U13717 (N_13717,N_11676,N_10814);
nand U13718 (N_13718,N_11521,N_10363);
xnor U13719 (N_13719,N_10467,N_11665);
nor U13720 (N_13720,N_11239,N_11161);
nor U13721 (N_13721,N_10953,N_10971);
and U13722 (N_13722,N_11055,N_10914);
nand U13723 (N_13723,N_11872,N_11306);
xnor U13724 (N_13724,N_10187,N_11403);
nor U13725 (N_13725,N_10491,N_11076);
or U13726 (N_13726,N_11335,N_11983);
nand U13727 (N_13727,N_10423,N_10611);
nand U13728 (N_13728,N_11160,N_11340);
nand U13729 (N_13729,N_11887,N_11884);
and U13730 (N_13730,N_11417,N_10966);
and U13731 (N_13731,N_10624,N_10271);
nand U13732 (N_13732,N_10681,N_10206);
nand U13733 (N_13733,N_11030,N_11262);
xor U13734 (N_13734,N_10498,N_11354);
xor U13735 (N_13735,N_10666,N_10965);
or U13736 (N_13736,N_11927,N_10294);
nor U13737 (N_13737,N_10470,N_10729);
or U13738 (N_13738,N_11396,N_10027);
and U13739 (N_13739,N_11361,N_10662);
nand U13740 (N_13740,N_11942,N_11000);
xor U13741 (N_13741,N_11922,N_10856);
nand U13742 (N_13742,N_10206,N_10656);
nor U13743 (N_13743,N_10422,N_10927);
nor U13744 (N_13744,N_11305,N_11055);
nor U13745 (N_13745,N_10774,N_10193);
nor U13746 (N_13746,N_10081,N_10401);
and U13747 (N_13747,N_11025,N_11669);
and U13748 (N_13748,N_10447,N_11431);
nand U13749 (N_13749,N_10241,N_11963);
nor U13750 (N_13750,N_11066,N_10443);
and U13751 (N_13751,N_10580,N_10428);
nand U13752 (N_13752,N_11036,N_11856);
nand U13753 (N_13753,N_10788,N_11443);
and U13754 (N_13754,N_10000,N_10171);
nand U13755 (N_13755,N_10643,N_11009);
xor U13756 (N_13756,N_11036,N_11829);
nor U13757 (N_13757,N_10454,N_10270);
nor U13758 (N_13758,N_10428,N_11676);
or U13759 (N_13759,N_10053,N_11126);
and U13760 (N_13760,N_10684,N_11003);
xnor U13761 (N_13761,N_10132,N_10487);
and U13762 (N_13762,N_10417,N_11342);
nand U13763 (N_13763,N_11233,N_10803);
and U13764 (N_13764,N_11071,N_10050);
and U13765 (N_13765,N_10715,N_11364);
nand U13766 (N_13766,N_10531,N_10946);
and U13767 (N_13767,N_10625,N_10367);
nand U13768 (N_13768,N_10817,N_11872);
nor U13769 (N_13769,N_11732,N_10579);
xnor U13770 (N_13770,N_10106,N_10128);
xnor U13771 (N_13771,N_11670,N_11331);
nand U13772 (N_13772,N_11752,N_11056);
or U13773 (N_13773,N_10914,N_11991);
or U13774 (N_13774,N_10659,N_11138);
nor U13775 (N_13775,N_10408,N_11083);
nor U13776 (N_13776,N_10448,N_11552);
or U13777 (N_13777,N_10183,N_10754);
nand U13778 (N_13778,N_10615,N_10660);
xnor U13779 (N_13779,N_11817,N_10591);
or U13780 (N_13780,N_11972,N_11398);
nand U13781 (N_13781,N_10947,N_11530);
xor U13782 (N_13782,N_11480,N_10785);
or U13783 (N_13783,N_11460,N_11414);
nor U13784 (N_13784,N_10484,N_11449);
and U13785 (N_13785,N_10503,N_10157);
or U13786 (N_13786,N_10374,N_11672);
nor U13787 (N_13787,N_11729,N_11938);
xnor U13788 (N_13788,N_11381,N_10681);
and U13789 (N_13789,N_10887,N_11229);
or U13790 (N_13790,N_11495,N_11527);
or U13791 (N_13791,N_11167,N_10586);
and U13792 (N_13792,N_10545,N_11033);
xor U13793 (N_13793,N_11773,N_10675);
nand U13794 (N_13794,N_10910,N_10135);
nor U13795 (N_13795,N_11841,N_10669);
xor U13796 (N_13796,N_10773,N_10249);
xnor U13797 (N_13797,N_10002,N_11897);
nor U13798 (N_13798,N_11851,N_11631);
xnor U13799 (N_13799,N_11836,N_11181);
nand U13800 (N_13800,N_10365,N_10415);
xor U13801 (N_13801,N_10306,N_10895);
nand U13802 (N_13802,N_10871,N_11418);
nand U13803 (N_13803,N_11313,N_10847);
or U13804 (N_13804,N_11539,N_11604);
and U13805 (N_13805,N_10952,N_10584);
nand U13806 (N_13806,N_10133,N_10863);
and U13807 (N_13807,N_11527,N_11702);
or U13808 (N_13808,N_10368,N_11611);
nand U13809 (N_13809,N_10168,N_10433);
or U13810 (N_13810,N_11964,N_10165);
xnor U13811 (N_13811,N_10438,N_11811);
nand U13812 (N_13812,N_10255,N_11128);
or U13813 (N_13813,N_10064,N_10033);
nand U13814 (N_13814,N_10398,N_11643);
nand U13815 (N_13815,N_10348,N_10938);
nand U13816 (N_13816,N_10888,N_11773);
or U13817 (N_13817,N_11008,N_11994);
and U13818 (N_13818,N_11281,N_11005);
nor U13819 (N_13819,N_11031,N_11795);
nand U13820 (N_13820,N_11362,N_10190);
or U13821 (N_13821,N_10406,N_10888);
nand U13822 (N_13822,N_11388,N_11154);
xnor U13823 (N_13823,N_10403,N_11842);
or U13824 (N_13824,N_10669,N_11859);
nor U13825 (N_13825,N_10902,N_10534);
or U13826 (N_13826,N_11549,N_10587);
nor U13827 (N_13827,N_10825,N_10707);
or U13828 (N_13828,N_10165,N_10666);
and U13829 (N_13829,N_10536,N_11168);
nand U13830 (N_13830,N_10829,N_11403);
xnor U13831 (N_13831,N_10190,N_11395);
nor U13832 (N_13832,N_11979,N_11405);
xnor U13833 (N_13833,N_10915,N_10202);
nand U13834 (N_13834,N_11565,N_11540);
xnor U13835 (N_13835,N_10149,N_10730);
nor U13836 (N_13836,N_10084,N_11061);
nor U13837 (N_13837,N_10872,N_10983);
nand U13838 (N_13838,N_11122,N_10253);
xor U13839 (N_13839,N_10003,N_11044);
and U13840 (N_13840,N_11503,N_10028);
nor U13841 (N_13841,N_10282,N_10956);
and U13842 (N_13842,N_10696,N_10755);
nor U13843 (N_13843,N_11926,N_10831);
nor U13844 (N_13844,N_11503,N_11498);
nand U13845 (N_13845,N_11693,N_11235);
or U13846 (N_13846,N_11568,N_10932);
xnor U13847 (N_13847,N_11471,N_11683);
and U13848 (N_13848,N_11461,N_11080);
xnor U13849 (N_13849,N_11242,N_11034);
nor U13850 (N_13850,N_10895,N_11758);
nand U13851 (N_13851,N_11570,N_10812);
nand U13852 (N_13852,N_10038,N_10727);
nor U13853 (N_13853,N_10541,N_10808);
xnor U13854 (N_13854,N_11522,N_10555);
xor U13855 (N_13855,N_10300,N_10928);
or U13856 (N_13856,N_11933,N_10787);
xor U13857 (N_13857,N_11058,N_11841);
nand U13858 (N_13858,N_10948,N_10742);
nand U13859 (N_13859,N_11023,N_10566);
nand U13860 (N_13860,N_10063,N_10907);
nand U13861 (N_13861,N_11517,N_11988);
xnor U13862 (N_13862,N_10112,N_11156);
xor U13863 (N_13863,N_11316,N_10655);
and U13864 (N_13864,N_11011,N_11301);
nand U13865 (N_13865,N_11837,N_10865);
and U13866 (N_13866,N_11210,N_10798);
nor U13867 (N_13867,N_10102,N_11872);
or U13868 (N_13868,N_11922,N_11148);
xor U13869 (N_13869,N_11417,N_10538);
nor U13870 (N_13870,N_11449,N_11765);
or U13871 (N_13871,N_10180,N_10938);
nand U13872 (N_13872,N_10241,N_11318);
xor U13873 (N_13873,N_10245,N_11568);
nand U13874 (N_13874,N_10700,N_11574);
nand U13875 (N_13875,N_10488,N_11568);
xnor U13876 (N_13876,N_11155,N_10674);
or U13877 (N_13877,N_10060,N_10479);
and U13878 (N_13878,N_10302,N_11177);
nand U13879 (N_13879,N_11713,N_10881);
and U13880 (N_13880,N_11034,N_11981);
and U13881 (N_13881,N_10581,N_10388);
or U13882 (N_13882,N_11327,N_11531);
and U13883 (N_13883,N_11499,N_10842);
xnor U13884 (N_13884,N_10824,N_10424);
and U13885 (N_13885,N_11054,N_11114);
xor U13886 (N_13886,N_11324,N_11771);
nand U13887 (N_13887,N_11507,N_10368);
or U13888 (N_13888,N_11784,N_10354);
or U13889 (N_13889,N_11135,N_11664);
or U13890 (N_13890,N_10733,N_10368);
nor U13891 (N_13891,N_10429,N_11841);
nand U13892 (N_13892,N_11554,N_11498);
xnor U13893 (N_13893,N_10789,N_10377);
nand U13894 (N_13894,N_11684,N_11373);
nor U13895 (N_13895,N_10516,N_11219);
nand U13896 (N_13896,N_11917,N_11536);
nor U13897 (N_13897,N_11310,N_10060);
xnor U13898 (N_13898,N_10292,N_10588);
xor U13899 (N_13899,N_11995,N_10637);
and U13900 (N_13900,N_11483,N_11441);
xnor U13901 (N_13901,N_10768,N_10828);
xor U13902 (N_13902,N_10895,N_11506);
or U13903 (N_13903,N_11605,N_11615);
xor U13904 (N_13904,N_10369,N_11584);
nor U13905 (N_13905,N_10164,N_10064);
or U13906 (N_13906,N_10771,N_11761);
or U13907 (N_13907,N_11605,N_11922);
nor U13908 (N_13908,N_11756,N_10755);
xnor U13909 (N_13909,N_11210,N_10942);
and U13910 (N_13910,N_10527,N_11226);
and U13911 (N_13911,N_10729,N_10605);
nor U13912 (N_13912,N_11048,N_11504);
or U13913 (N_13913,N_11129,N_10622);
xnor U13914 (N_13914,N_11615,N_10287);
or U13915 (N_13915,N_10090,N_10808);
xor U13916 (N_13916,N_10865,N_10211);
nor U13917 (N_13917,N_10532,N_11571);
nand U13918 (N_13918,N_11293,N_10122);
nand U13919 (N_13919,N_11016,N_11580);
xor U13920 (N_13920,N_10553,N_10256);
xnor U13921 (N_13921,N_10883,N_11885);
or U13922 (N_13922,N_10346,N_10874);
xnor U13923 (N_13923,N_10734,N_10885);
nand U13924 (N_13924,N_10457,N_10824);
and U13925 (N_13925,N_10681,N_11666);
or U13926 (N_13926,N_11859,N_10463);
nand U13927 (N_13927,N_11995,N_11376);
nand U13928 (N_13928,N_10396,N_11177);
nor U13929 (N_13929,N_10305,N_11498);
nor U13930 (N_13930,N_11590,N_10175);
and U13931 (N_13931,N_11552,N_10549);
nand U13932 (N_13932,N_11249,N_11241);
nor U13933 (N_13933,N_11814,N_10316);
nand U13934 (N_13934,N_11319,N_11188);
nand U13935 (N_13935,N_10493,N_10330);
and U13936 (N_13936,N_10374,N_10995);
nor U13937 (N_13937,N_10071,N_11606);
or U13938 (N_13938,N_10308,N_10361);
nor U13939 (N_13939,N_11985,N_10903);
or U13940 (N_13940,N_10480,N_10483);
and U13941 (N_13941,N_11932,N_11785);
and U13942 (N_13942,N_11747,N_10922);
and U13943 (N_13943,N_11982,N_11485);
nor U13944 (N_13944,N_11502,N_10431);
xnor U13945 (N_13945,N_11840,N_11405);
or U13946 (N_13946,N_11866,N_10638);
xnor U13947 (N_13947,N_11838,N_11579);
nand U13948 (N_13948,N_10944,N_10294);
or U13949 (N_13949,N_10942,N_10815);
or U13950 (N_13950,N_11963,N_11463);
and U13951 (N_13951,N_10042,N_10530);
nor U13952 (N_13952,N_10338,N_11253);
xnor U13953 (N_13953,N_11834,N_10781);
xor U13954 (N_13954,N_10303,N_10489);
or U13955 (N_13955,N_10031,N_10904);
nor U13956 (N_13956,N_11677,N_10902);
and U13957 (N_13957,N_10769,N_11205);
nor U13958 (N_13958,N_11639,N_10289);
nor U13959 (N_13959,N_10042,N_11191);
nand U13960 (N_13960,N_10017,N_11614);
or U13961 (N_13961,N_10358,N_10065);
nand U13962 (N_13962,N_10491,N_11319);
nor U13963 (N_13963,N_10480,N_10540);
xor U13964 (N_13964,N_11839,N_10383);
nand U13965 (N_13965,N_11923,N_11060);
nor U13966 (N_13966,N_11077,N_10360);
or U13967 (N_13967,N_11984,N_10472);
and U13968 (N_13968,N_11198,N_11028);
xnor U13969 (N_13969,N_11289,N_10960);
nor U13970 (N_13970,N_11712,N_11136);
or U13971 (N_13971,N_10597,N_10849);
and U13972 (N_13972,N_11527,N_10481);
nand U13973 (N_13973,N_10538,N_11698);
nand U13974 (N_13974,N_10289,N_11960);
or U13975 (N_13975,N_11646,N_10458);
nor U13976 (N_13976,N_10643,N_10546);
xor U13977 (N_13977,N_10285,N_10801);
nor U13978 (N_13978,N_11649,N_11670);
nand U13979 (N_13979,N_10299,N_11157);
or U13980 (N_13980,N_10748,N_10873);
xor U13981 (N_13981,N_11589,N_10443);
xor U13982 (N_13982,N_10816,N_11470);
nor U13983 (N_13983,N_10403,N_11423);
nor U13984 (N_13984,N_10491,N_10383);
and U13985 (N_13985,N_10793,N_11088);
nor U13986 (N_13986,N_10450,N_11416);
nor U13987 (N_13987,N_10001,N_10455);
xor U13988 (N_13988,N_11592,N_10864);
nor U13989 (N_13989,N_11279,N_10380);
nor U13990 (N_13990,N_11450,N_10121);
xor U13991 (N_13991,N_11426,N_10345);
or U13992 (N_13992,N_10014,N_10537);
nor U13993 (N_13993,N_11811,N_11111);
nor U13994 (N_13994,N_10305,N_11659);
nand U13995 (N_13995,N_11627,N_10835);
or U13996 (N_13996,N_11356,N_10468);
nor U13997 (N_13997,N_11482,N_11742);
nor U13998 (N_13998,N_10218,N_10424);
nand U13999 (N_13999,N_11862,N_10938);
nand U14000 (N_14000,N_13242,N_13139);
nor U14001 (N_14001,N_12946,N_12341);
nor U14002 (N_14002,N_13959,N_13106);
nor U14003 (N_14003,N_12949,N_12947);
and U14004 (N_14004,N_12011,N_12756);
or U14005 (N_14005,N_13868,N_13880);
nor U14006 (N_14006,N_12176,N_13903);
nor U14007 (N_14007,N_13526,N_13873);
or U14008 (N_14008,N_12021,N_13252);
nand U14009 (N_14009,N_13041,N_13766);
or U14010 (N_14010,N_13324,N_12244);
xor U14011 (N_14011,N_12932,N_12173);
nor U14012 (N_14012,N_12207,N_13897);
or U14013 (N_14013,N_13973,N_12983);
nand U14014 (N_14014,N_13877,N_12823);
or U14015 (N_14015,N_13121,N_13616);
nand U14016 (N_14016,N_12449,N_13478);
or U14017 (N_14017,N_13112,N_13827);
nand U14018 (N_14018,N_13376,N_12027);
and U14019 (N_14019,N_12772,N_12688);
xnor U14020 (N_14020,N_12632,N_13931);
or U14021 (N_14021,N_12258,N_12738);
or U14022 (N_14022,N_13605,N_13489);
nor U14023 (N_14023,N_12408,N_12092);
nand U14024 (N_14024,N_13234,N_12369);
xor U14025 (N_14025,N_13350,N_13800);
xor U14026 (N_14026,N_13179,N_12787);
nor U14027 (N_14027,N_13963,N_12054);
and U14028 (N_14028,N_13365,N_13983);
and U14029 (N_14029,N_13803,N_12733);
or U14030 (N_14030,N_13673,N_12612);
nor U14031 (N_14031,N_13322,N_13101);
nor U14032 (N_14032,N_12046,N_12058);
xor U14033 (N_14033,N_13011,N_12421);
or U14034 (N_14034,N_12468,N_13721);
nor U14035 (N_14035,N_13355,N_12479);
nand U14036 (N_14036,N_12981,N_12559);
or U14037 (N_14037,N_13163,N_13074);
nand U14038 (N_14038,N_13127,N_12890);
and U14039 (N_14039,N_13028,N_12859);
or U14040 (N_14040,N_12610,N_12619);
nand U14041 (N_14041,N_12144,N_12695);
nor U14042 (N_14042,N_13644,N_12831);
and U14043 (N_14043,N_13250,N_13681);
nor U14044 (N_14044,N_13889,N_12305);
and U14045 (N_14045,N_12069,N_12972);
and U14046 (N_14046,N_13772,N_12065);
or U14047 (N_14047,N_13885,N_12237);
and U14048 (N_14048,N_12243,N_13842);
nor U14049 (N_14049,N_13439,N_12259);
or U14050 (N_14050,N_12709,N_12793);
xnor U14051 (N_14051,N_13913,N_12440);
xnor U14052 (N_14052,N_13709,N_13178);
nand U14053 (N_14053,N_13937,N_13536);
nor U14054 (N_14054,N_12541,N_13302);
xnor U14055 (N_14055,N_12804,N_13735);
and U14056 (N_14056,N_13646,N_12416);
or U14057 (N_14057,N_13342,N_12002);
nand U14058 (N_14058,N_12893,N_13136);
nand U14059 (N_14059,N_13490,N_13484);
and U14060 (N_14060,N_13278,N_13154);
xor U14061 (N_14061,N_13327,N_13148);
and U14062 (N_14062,N_12669,N_12064);
and U14063 (N_14063,N_12912,N_13155);
nand U14064 (N_14064,N_13883,N_13660);
xor U14065 (N_14065,N_12419,N_13864);
nor U14066 (N_14066,N_12097,N_12781);
xnor U14067 (N_14067,N_12013,N_12569);
and U14068 (N_14068,N_13259,N_12673);
xnor U14069 (N_14069,N_12750,N_13021);
or U14070 (N_14070,N_12825,N_13576);
or U14071 (N_14071,N_12889,N_12677);
xnor U14072 (N_14072,N_12216,N_13131);
xnor U14073 (N_14073,N_13916,N_13182);
or U14074 (N_14074,N_12422,N_13509);
nor U14075 (N_14075,N_12347,N_13346);
and U14076 (N_14076,N_13780,N_12114);
nor U14077 (N_14077,N_13831,N_13216);
and U14078 (N_14078,N_13549,N_12463);
or U14079 (N_14079,N_13239,N_13656);
and U14080 (N_14080,N_13450,N_13675);
nor U14081 (N_14081,N_13991,N_13690);
and U14082 (N_14082,N_12155,N_12183);
xnor U14083 (N_14083,N_12840,N_13017);
xnor U14084 (N_14084,N_13285,N_12068);
xor U14085 (N_14085,N_13705,N_12799);
xnor U14086 (N_14086,N_12521,N_12314);
nand U14087 (N_14087,N_12138,N_13826);
xor U14088 (N_14088,N_13953,N_13020);
and U14089 (N_14089,N_12993,N_12194);
or U14090 (N_14090,N_13980,N_13366);
or U14091 (N_14091,N_12077,N_12676);
nand U14092 (N_14092,N_12289,N_12435);
and U14093 (N_14093,N_12844,N_12407);
and U14094 (N_14094,N_13978,N_13714);
or U14095 (N_14095,N_13144,N_13098);
xnor U14096 (N_14096,N_13201,N_13624);
or U14097 (N_14097,N_13898,N_12806);
nand U14098 (N_14098,N_13422,N_12248);
or U14099 (N_14099,N_12241,N_12641);
nor U14100 (N_14100,N_12420,N_12556);
and U14101 (N_14101,N_13486,N_12461);
nor U14102 (N_14102,N_13974,N_13005);
nor U14103 (N_14103,N_12627,N_13400);
or U14104 (N_14104,N_12494,N_12220);
nor U14105 (N_14105,N_13286,N_13798);
or U14106 (N_14106,N_12953,N_12024);
and U14107 (N_14107,N_12557,N_13156);
nor U14108 (N_14108,N_13396,N_12158);
and U14109 (N_14109,N_12417,N_12121);
and U14110 (N_14110,N_13501,N_12473);
and U14111 (N_14111,N_13844,N_12734);
nor U14112 (N_14112,N_13961,N_13134);
nand U14113 (N_14113,N_12376,N_12814);
nand U14114 (N_14114,N_12399,N_12218);
and U14115 (N_14115,N_13778,N_13640);
xor U14116 (N_14116,N_13702,N_13494);
xor U14117 (N_14117,N_13226,N_12919);
and U14118 (N_14118,N_12916,N_13861);
nand U14119 (N_14119,N_13001,N_12066);
and U14120 (N_14120,N_12096,N_13792);
and U14121 (N_14121,N_13858,N_12899);
nand U14122 (N_14122,N_12712,N_13161);
xor U14123 (N_14123,N_12251,N_12987);
nand U14124 (N_14124,N_12204,N_12699);
and U14125 (N_14125,N_12434,N_12043);
nor U14126 (N_14126,N_12892,N_13756);
xor U14127 (N_14127,N_12458,N_13957);
or U14128 (N_14128,N_13905,N_12891);
and U14129 (N_14129,N_13232,N_13398);
nor U14130 (N_14130,N_12165,N_12731);
nor U14131 (N_14131,N_13231,N_13520);
nand U14132 (N_14132,N_13693,N_13661);
nand U14133 (N_14133,N_12273,N_13678);
and U14134 (N_14134,N_12265,N_13901);
xnor U14135 (N_14135,N_12585,N_12256);
or U14136 (N_14136,N_13689,N_12506);
nor U14137 (N_14137,N_12701,N_12741);
or U14138 (N_14138,N_12328,N_13846);
or U14139 (N_14139,N_13888,N_13513);
nand U14140 (N_14140,N_12430,N_12360);
nor U14141 (N_14141,N_12729,N_12877);
or U14142 (N_14142,N_12812,N_12615);
xnor U14143 (N_14143,N_13863,N_13191);
and U14144 (N_14144,N_12446,N_12854);
nand U14145 (N_14145,N_12540,N_13908);
nor U14146 (N_14146,N_13315,N_12000);
and U14147 (N_14147,N_12147,N_13288);
or U14148 (N_14148,N_13395,N_12425);
nor U14149 (N_14149,N_13171,N_13012);
nand U14150 (N_14150,N_13471,N_12211);
nor U14151 (N_14151,N_12965,N_12785);
xor U14152 (N_14152,N_13024,N_13596);
nand U14153 (N_14153,N_12941,N_12480);
or U14154 (N_14154,N_12390,N_13264);
nor U14155 (N_14155,N_13409,N_13195);
or U14156 (N_14156,N_12040,N_13577);
and U14157 (N_14157,N_12386,N_12606);
nor U14158 (N_14158,N_13502,N_12613);
nand U14159 (N_14159,N_13696,N_12291);
xor U14160 (N_14160,N_12548,N_12990);
and U14161 (N_14161,N_12022,N_12570);
and U14162 (N_14162,N_12295,N_13951);
xor U14163 (N_14163,N_12576,N_12202);
or U14164 (N_14164,N_12842,N_13639);
or U14165 (N_14165,N_13956,N_12514);
and U14166 (N_14166,N_12490,N_12682);
or U14167 (N_14167,N_13022,N_12736);
nor U14168 (N_14168,N_12751,N_13432);
and U14169 (N_14169,N_12924,N_12552);
and U14170 (N_14170,N_12937,N_13924);
nand U14171 (N_14171,N_12284,N_13850);
nor U14172 (N_14172,N_12384,N_13891);
nand U14173 (N_14173,N_13051,N_13741);
xnor U14174 (N_14174,N_13500,N_13782);
nand U14175 (N_14175,N_12107,N_12604);
or U14176 (N_14176,N_12979,N_12443);
nand U14177 (N_14177,N_12456,N_12658);
nor U14178 (N_14178,N_12796,N_12162);
and U14179 (N_14179,N_12670,N_13065);
xnor U14180 (N_14180,N_13033,N_12830);
and U14181 (N_14181,N_12603,N_13375);
nor U14182 (N_14182,N_13541,N_12190);
and U14183 (N_14183,N_12780,N_13097);
xor U14184 (N_14184,N_13575,N_13706);
nand U14185 (N_14185,N_12774,N_13755);
nor U14186 (N_14186,N_12678,N_13967);
xor U14187 (N_14187,N_12856,N_12039);
or U14188 (N_14188,N_12227,N_12119);
xor U14189 (N_14189,N_12511,N_13157);
nand U14190 (N_14190,N_12336,N_12389);
and U14191 (N_14191,N_12685,N_12622);
or U14192 (N_14192,N_13902,N_12404);
and U14193 (N_14193,N_13305,N_13926);
nor U14194 (N_14194,N_13124,N_12187);
nor U14195 (N_14195,N_13110,N_13445);
and U14196 (N_14196,N_13413,N_13146);
nand U14197 (N_14197,N_13194,N_13421);
nand U14198 (N_14198,N_13614,N_12030);
nor U14199 (N_14199,N_12084,N_12483);
or U14200 (N_14200,N_13184,N_12869);
and U14201 (N_14201,N_12795,N_12075);
nor U14202 (N_14202,N_12359,N_12116);
and U14203 (N_14203,N_13254,N_12574);
xnor U14204 (N_14204,N_12459,N_13518);
or U14205 (N_14205,N_13204,N_13274);
nor U14206 (N_14206,N_12992,N_13562);
or U14207 (N_14207,N_13372,N_13567);
nor U14208 (N_14208,N_12356,N_12624);
and U14209 (N_14209,N_13406,N_13572);
or U14210 (N_14210,N_12105,N_13843);
xor U14211 (N_14211,N_12402,N_13103);
nand U14212 (N_14212,N_12855,N_13467);
nor U14213 (N_14213,N_12783,N_12128);
or U14214 (N_14214,N_13440,N_13728);
nand U14215 (N_14215,N_12059,N_13986);
and U14216 (N_14216,N_12395,N_12179);
nand U14217 (N_14217,N_13802,N_12807);
xnor U14218 (N_14218,N_12154,N_13433);
and U14219 (N_14219,N_12631,N_13952);
or U14220 (N_14220,N_12055,N_12224);
nor U14221 (N_14221,N_13817,N_13424);
nand U14222 (N_14222,N_13828,N_13739);
nor U14223 (N_14223,N_12522,N_12726);
nor U14224 (N_14224,N_12076,N_13860);
xnor U14225 (N_14225,N_13192,N_13308);
xor U14226 (N_14226,N_13448,N_12275);
nor U14227 (N_14227,N_13708,N_12429);
nand U14228 (N_14228,N_12927,N_13167);
nor U14229 (N_14229,N_13746,N_13466);
and U14230 (N_14230,N_13634,N_13046);
nor U14231 (N_14231,N_12464,N_12038);
or U14232 (N_14232,N_12482,N_13933);
xnor U14233 (N_14233,N_12755,N_12888);
xnor U14234 (N_14234,N_12820,N_13687);
nor U14235 (N_14235,N_13267,N_12809);
xor U14236 (N_14236,N_12801,N_13998);
nand U14237 (N_14237,N_13193,N_12880);
nand U14238 (N_14238,N_13674,N_12135);
nor U14239 (N_14239,N_13283,N_12597);
xnor U14240 (N_14240,N_13840,N_12846);
xnor U14241 (N_14241,N_13205,N_13699);
xnor U14242 (N_14242,N_12383,N_12872);
or U14243 (N_14243,N_12088,N_13886);
nor U14244 (N_14244,N_12991,N_13944);
and U14245 (N_14245,N_13629,N_12438);
or U14246 (N_14246,N_13377,N_12231);
xor U14247 (N_14247,N_12832,N_13474);
and U14248 (N_14248,N_12486,N_12431);
xnor U14249 (N_14249,N_13909,N_13071);
nand U14250 (N_14250,N_13233,N_12454);
xnor U14251 (N_14251,N_12499,N_13558);
nand U14252 (N_14252,N_12197,N_13632);
nand U14253 (N_14253,N_13092,N_12131);
xor U14254 (N_14254,N_13790,N_13982);
and U14255 (N_14255,N_12943,N_12042);
or U14256 (N_14256,N_12942,N_12873);
nor U14257 (N_14257,N_12394,N_12562);
and U14258 (N_14258,N_13943,N_12436);
or U14259 (N_14259,N_12954,N_13105);
or U14260 (N_14260,N_12193,N_13807);
and U14261 (N_14261,N_12591,N_12598);
xor U14262 (N_14262,N_12381,N_13525);
or U14263 (N_14263,N_13565,N_12827);
or U14264 (N_14264,N_13715,N_12730);
and U14265 (N_14265,N_12245,N_13397);
or U14266 (N_14266,N_12644,N_13934);
and U14267 (N_14267,N_13896,N_13202);
nor U14268 (N_14268,N_13227,N_12026);
and U14269 (N_14269,N_13096,N_13691);
xor U14270 (N_14270,N_13971,N_13917);
and U14271 (N_14271,N_12593,N_13206);
nor U14272 (N_14272,N_12509,N_12062);
and U14273 (N_14273,N_13857,N_13253);
and U14274 (N_14274,N_13418,N_12023);
or U14275 (N_14275,N_13160,N_12998);
or U14276 (N_14276,N_12818,N_12634);
nand U14277 (N_14277,N_13704,N_13527);
xnor U14278 (N_14278,N_13540,N_12952);
nor U14279 (N_14279,N_13488,N_12922);
xor U14280 (N_14280,N_13208,N_12274);
nand U14281 (N_14281,N_13138,N_12684);
or U14282 (N_14282,N_12415,N_12721);
xor U14283 (N_14283,N_12316,N_13373);
nor U14284 (N_14284,N_12614,N_12448);
nand U14285 (N_14285,N_13276,N_12142);
xnor U14286 (N_14286,N_12255,N_13764);
or U14287 (N_14287,N_12852,N_13805);
and U14288 (N_14288,N_13351,N_13894);
and U14289 (N_14289,N_13218,N_13023);
xnor U14290 (N_14290,N_12073,N_12323);
or U14291 (N_14291,N_13085,N_12784);
or U14292 (N_14292,N_13415,N_12348);
and U14293 (N_14293,N_12764,N_13465);
or U14294 (N_14294,N_12516,N_12298);
nor U14295 (N_14295,N_12626,N_13052);
or U14296 (N_14296,N_13174,N_12029);
xnor U14297 (N_14297,N_12413,N_12303);
or U14298 (N_14298,N_12513,N_13859);
xnor U14299 (N_14299,N_13650,N_12582);
or U14300 (N_14300,N_12287,N_12045);
nand U14301 (N_14301,N_13940,N_12321);
nor U14302 (N_14302,N_12260,N_13316);
nand U14303 (N_14303,N_13137,N_13468);
and U14304 (N_14304,N_12329,N_12087);
or U14305 (N_14305,N_12571,N_12444);
nor U14306 (N_14306,N_12178,N_13716);
or U14307 (N_14307,N_12004,N_13410);
and U14308 (N_14308,N_13722,N_13679);
nand U14309 (N_14309,N_13523,N_13635);
xnor U14310 (N_14310,N_13811,N_13820);
nor U14311 (N_14311,N_12645,N_13662);
nor U14312 (N_14312,N_13969,N_13119);
nand U14313 (N_14313,N_12938,N_13356);
nor U14314 (N_14314,N_13126,N_12277);
or U14315 (N_14315,N_12581,N_13919);
and U14316 (N_14316,N_12379,N_12308);
or U14317 (N_14317,N_13993,N_12080);
and U14318 (N_14318,N_13870,N_12286);
and U14319 (N_14319,N_12501,N_13947);
nand U14320 (N_14320,N_13628,N_12910);
and U14321 (N_14321,N_12654,N_12884);
or U14322 (N_14322,N_12980,N_13570);
nand U14323 (N_14323,N_13214,N_13834);
or U14324 (N_14324,N_13698,N_13677);
nand U14325 (N_14325,N_13701,N_13884);
nor U14326 (N_14326,N_12355,N_13994);
nand U14327 (N_14327,N_13469,N_12428);
nand U14328 (N_14328,N_13580,N_12519);
nor U14329 (N_14329,N_13149,N_13318);
nor U14330 (N_14330,N_13479,N_13970);
nor U14331 (N_14331,N_12391,N_13882);
xor U14332 (N_14332,N_13747,N_12725);
nor U14333 (N_14333,N_13289,N_12380);
or U14334 (N_14334,N_12285,N_12534);
or U14335 (N_14335,N_12607,N_13434);
and U14336 (N_14336,N_12166,N_12007);
and U14337 (N_14337,N_12748,N_13918);
nor U14338 (N_14338,N_12403,N_13881);
xnor U14339 (N_14339,N_12471,N_13320);
nor U14340 (N_14340,N_13791,N_13784);
or U14341 (N_14341,N_13522,N_13564);
xor U14342 (N_14342,N_13744,N_12469);
and U14343 (N_14343,N_13364,N_12957);
nor U14344 (N_14344,N_12169,N_12909);
or U14345 (N_14345,N_12765,N_13925);
xor U14346 (N_14346,N_12281,N_13977);
xnor U14347 (N_14347,N_13050,N_13006);
nor U14348 (N_14348,N_13865,N_12487);
nor U14349 (N_14349,N_13874,N_13477);
xor U14350 (N_14350,N_13555,N_13142);
nand U14351 (N_14351,N_13554,N_13293);
nor U14352 (N_14352,N_13987,N_12112);
nand U14353 (N_14353,N_12319,N_12962);
nor U14354 (N_14354,N_13326,N_12775);
nand U14355 (N_14355,N_12815,N_12526);
nor U14356 (N_14356,N_13695,N_12186);
xnor U14357 (N_14357,N_13072,N_12249);
nand U14358 (N_14358,N_13426,N_12406);
or U14359 (N_14359,N_13945,N_13626);
and U14360 (N_14360,N_13579,N_13030);
nor U14361 (N_14361,N_13476,N_12271);
xor U14362 (N_14362,N_13496,N_12609);
nand U14363 (N_14363,N_12090,N_13962);
and U14364 (N_14364,N_12450,N_13453);
and U14365 (N_14365,N_12817,N_12517);
or U14366 (N_14366,N_12498,N_13009);
nor U14367 (N_14367,N_13700,N_12344);
or U14368 (N_14368,N_13775,N_13323);
or U14369 (N_14369,N_13258,N_12834);
nor U14370 (N_14370,N_12020,N_13852);
xor U14371 (N_14371,N_12697,N_12761);
and U14372 (N_14372,N_13984,N_12867);
xor U14373 (N_14373,N_13370,N_12675);
nor U14374 (N_14374,N_12887,N_13303);
nor U14375 (N_14375,N_13382,N_13212);
and U14376 (N_14376,N_13759,N_13284);
and U14377 (N_14377,N_13543,N_13334);
nor U14378 (N_14378,N_12172,N_12340);
or U14379 (N_14379,N_13016,N_12951);
or U14380 (N_14380,N_13654,N_12970);
and U14381 (N_14381,N_12717,N_13153);
and U14382 (N_14382,N_12320,N_13597);
and U14383 (N_14383,N_13330,N_12550);
or U14384 (N_14384,N_13581,N_12595);
nand U14385 (N_14385,N_12306,N_12948);
nand U14386 (N_14386,N_12520,N_13102);
nor U14387 (N_14387,N_12779,N_12367);
and U14388 (N_14388,N_12010,N_13599);
and U14389 (N_14389,N_12374,N_13277);
or U14390 (N_14390,N_13717,N_13649);
nor U14391 (N_14391,N_13095,N_13412);
xnor U14392 (N_14392,N_12442,N_13093);
and U14393 (N_14393,N_13813,N_13246);
nand U14394 (N_14394,N_13228,N_13292);
xnor U14395 (N_14395,N_12182,N_12836);
xor U14396 (N_14396,N_12460,N_13055);
nor U14397 (N_14397,N_12518,N_12918);
xor U14398 (N_14398,N_12657,N_12439);
nor U14399 (N_14399,N_12125,N_13796);
xnor U14400 (N_14400,N_12588,N_12085);
and U14401 (N_14401,N_12120,N_12681);
xnor U14402 (N_14402,N_12876,N_12578);
and U14403 (N_14403,N_12542,N_12537);
xor U14404 (N_14404,N_13298,N_12648);
xor U14405 (N_14405,N_13053,N_13388);
xnor U14406 (N_14406,N_12544,N_13595);
nor U14407 (N_14407,N_13306,N_13657);
nor U14408 (N_14408,N_13109,N_12156);
and U14409 (N_14409,N_13912,N_13039);
xnor U14410 (N_14410,N_12914,N_13879);
nand U14411 (N_14411,N_12358,N_12372);
or U14412 (N_14412,N_12200,N_12475);
or U14413 (N_14413,N_12203,N_12385);
nand U14414 (N_14414,N_12565,N_12504);
or U14415 (N_14415,N_13872,N_12773);
or U14416 (N_14416,N_13740,N_12145);
nor U14417 (N_14417,N_13773,N_13210);
nor U14418 (N_14418,N_12174,N_13645);
and U14419 (N_14419,N_12920,N_12976);
or U14420 (N_14420,N_13235,N_12950);
nor U14421 (N_14421,N_12524,N_12944);
and U14422 (N_14422,N_13829,N_13019);
nor U14423 (N_14423,N_12651,N_12387);
or U14424 (N_14424,N_13435,N_13026);
xor U14425 (N_14425,N_13383,N_13979);
or U14426 (N_14426,N_13942,N_13213);
nor U14427 (N_14427,N_13738,N_12491);
nor U14428 (N_14428,N_13187,N_12445);
and U14429 (N_14429,N_12343,N_13615);
xnor U14430 (N_14430,N_13553,N_13753);
and U14431 (N_14431,N_13578,N_13394);
xor U14432 (N_14432,N_13362,N_12051);
xor U14433 (N_14433,N_13186,N_12232);
nand U14434 (N_14434,N_12126,N_13869);
xnor U14435 (N_14435,N_12288,N_12017);
or U14436 (N_14436,N_12310,N_13841);
or U14437 (N_14437,N_13180,N_12364);
or U14438 (N_14438,N_12098,N_13655);
or U14439 (N_14439,N_13168,N_13610);
nor U14440 (N_14440,N_12961,N_12102);
and U14441 (N_14441,N_12307,N_12740);
nand U14442 (N_14442,N_13013,N_12997);
or U14443 (N_14443,N_13367,N_13524);
nor U14444 (N_14444,N_12882,N_13256);
or U14445 (N_14445,N_13499,N_12269);
nand U14446 (N_14446,N_13911,N_12579);
nor U14447 (N_14447,N_13401,N_12837);
xor U14448 (N_14448,N_13236,N_12535);
nand U14449 (N_14449,N_13594,N_12122);
or U14450 (N_14450,N_12056,N_12759);
nor U14451 (N_14451,N_13456,N_13748);
xnor U14452 (N_14452,N_12163,N_13958);
or U14453 (N_14453,N_12841,N_13262);
xor U14454 (N_14454,N_13459,N_13862);
xor U14455 (N_14455,N_13839,N_13243);
or U14456 (N_14456,N_12283,N_13783);
xor U14457 (N_14457,N_13516,N_12149);
nand U14458 (N_14458,N_12235,N_13244);
nand U14459 (N_14459,N_12130,N_13141);
nor U14460 (N_14460,N_12412,N_13732);
and U14461 (N_14461,N_12140,N_13932);
and U14462 (N_14462,N_13613,N_12318);
nand U14463 (N_14463,N_13871,N_12838);
and U14464 (N_14464,N_13018,N_13084);
or U14465 (N_14465,N_13344,N_13530);
and U14466 (N_14466,N_12636,N_12667);
nor U14467 (N_14467,N_12382,N_12188);
and U14468 (N_14468,N_12123,N_12396);
nand U14469 (N_14469,N_13703,N_12555);
nand U14470 (N_14470,N_12037,N_13671);
nor U14471 (N_14471,N_13920,N_13606);
xnor U14472 (N_14472,N_13164,N_12354);
and U14473 (N_14473,N_12050,N_13392);
and U14474 (N_14474,N_13463,N_13057);
nor U14475 (N_14475,N_12349,N_13140);
or U14476 (N_14476,N_13769,N_13574);
and U14477 (N_14477,N_12324,N_13710);
nand U14478 (N_14478,N_13222,N_12956);
nand U14479 (N_14479,N_13545,N_13321);
nand U14480 (N_14480,N_12782,N_13789);
or U14481 (N_14481,N_13079,N_13379);
nand U14482 (N_14482,N_13548,N_13785);
or U14483 (N_14483,N_12679,N_13151);
nor U14484 (N_14484,N_12536,N_12587);
nor U14485 (N_14485,N_12008,N_13825);
nand U14486 (N_14486,N_12530,N_13539);
nor U14487 (N_14487,N_13751,N_13712);
nor U14488 (N_14488,N_13313,N_13960);
and U14489 (N_14489,N_12019,N_13713);
nand U14490 (N_14490,N_12230,N_13295);
and U14491 (N_14491,N_12628,N_12527);
nand U14492 (N_14492,N_12048,N_13669);
or U14493 (N_14493,N_13135,N_12655);
nor U14494 (N_14494,N_13358,N_12294);
nand U14495 (N_14495,N_13128,N_13642);
or U14496 (N_14496,N_12934,N_13240);
xor U14497 (N_14497,N_13866,N_12723);
and U14498 (N_14498,N_12053,N_12226);
xor U14499 (N_14499,N_12794,N_13310);
and U14500 (N_14500,N_12160,N_12564);
or U14501 (N_14501,N_12014,N_12739);
or U14502 (N_14502,N_13380,N_13014);
or U14503 (N_14503,N_13427,N_13988);
and U14504 (N_14504,N_13799,N_12637);
nand U14505 (N_14505,N_13291,N_12963);
xnor U14506 (N_14506,N_12242,N_13263);
nand U14507 (N_14507,N_12653,N_13172);
nand U14508 (N_14508,N_12339,N_12713);
or U14509 (N_14509,N_12629,N_13685);
or U14510 (N_14510,N_12333,N_13795);
or U14511 (N_14511,N_13008,N_12700);
nor U14512 (N_14512,N_13972,N_12605);
and U14513 (N_14513,N_13215,N_12378);
and U14514 (N_14514,N_12665,N_12647);
and U14515 (N_14515,N_12508,N_13776);
nor U14516 (N_14516,N_12999,N_12862);
and U14517 (N_14517,N_12254,N_12638);
nand U14518 (N_14518,N_13521,N_12489);
nand U14519 (N_14519,N_13374,N_13651);
xnor U14520 (N_14520,N_12091,N_12505);
nor U14521 (N_14521,N_13823,N_12497);
nand U14522 (N_14522,N_12219,N_12272);
nor U14523 (N_14523,N_12594,N_13935);
xnor U14524 (N_14524,N_12345,N_13617);
xor U14525 (N_14525,N_12845,N_12928);
xor U14526 (N_14526,N_13419,N_12371);
nand U14527 (N_14527,N_12006,N_12586);
and U14528 (N_14528,N_12763,N_13810);
nand U14529 (N_14529,N_13907,N_13338);
nand U14530 (N_14530,N_12315,N_13637);
nor U14531 (N_14531,N_13551,N_12968);
xnor U14532 (N_14532,N_12032,N_12223);
xnor U14533 (N_14533,N_13152,N_13498);
nand U14534 (N_14534,N_12083,N_12363);
nand U14535 (N_14535,N_12955,N_12268);
or U14536 (N_14536,N_13718,N_13335);
nand U14537 (N_14537,N_12279,N_13493);
or U14538 (N_14538,N_13771,N_12561);
nor U14539 (N_14539,N_13665,N_12301);
and U14540 (N_14540,N_13584,N_12789);
nor U14541 (N_14541,N_13528,N_13217);
nor U14542 (N_14542,N_13462,N_12874);
or U14543 (N_14543,N_12485,N_13515);
or U14544 (N_14544,N_13169,N_12640);
nand U14545 (N_14545,N_12253,N_13837);
or U14546 (N_14546,N_13504,N_13762);
nor U14547 (N_14547,N_12635,N_13088);
xor U14548 (N_14548,N_13573,N_12826);
and U14549 (N_14549,N_12798,N_13078);
nand U14550 (N_14550,N_13353,N_13280);
nor U14551 (N_14551,N_12805,N_12964);
nor U14552 (N_14552,N_13354,N_12863);
nor U14553 (N_14553,N_13441,N_12225);
or U14554 (N_14554,N_13587,N_13929);
or U14555 (N_14555,N_12554,N_13765);
nand U14556 (N_14556,N_13995,N_12690);
or U14557 (N_14557,N_13070,N_13165);
xor U14558 (N_14558,N_13768,N_12282);
nor U14559 (N_14559,N_13633,N_13992);
and U14560 (N_14560,N_12545,N_13900);
nand U14561 (N_14561,N_13430,N_13720);
xor U14562 (N_14562,N_12878,N_13534);
or U14563 (N_14563,N_13757,N_12317);
and U14564 (N_14564,N_12332,N_13038);
nor U14565 (N_14565,N_12671,N_12896);
and U14566 (N_14566,N_12760,N_13801);
or U14567 (N_14567,N_13120,N_12322);
nand U14568 (N_14568,N_12134,N_12861);
and U14569 (N_14569,N_12706,N_12477);
and U14570 (N_14570,N_12558,N_13927);
and U14571 (N_14571,N_13188,N_12745);
nand U14572 (N_14572,N_12935,N_12642);
and U14573 (N_14573,N_12813,N_12860);
or U14574 (N_14574,N_12239,N_12931);
xor U14575 (N_14575,N_13269,N_13438);
xor U14576 (N_14576,N_13627,N_12099);
or U14577 (N_14577,N_13517,N_13473);
and U14578 (N_14578,N_13505,N_12865);
nand U14579 (N_14579,N_12462,N_12252);
xor U14580 (N_14580,N_12724,N_13118);
or U14581 (N_14581,N_13936,N_13048);
and U14582 (N_14582,N_13794,N_13428);
nand U14583 (N_14583,N_12549,N_12365);
nand U14584 (N_14584,N_12103,N_13608);
nand U14585 (N_14585,N_13510,N_13123);
nand U14586 (N_14586,N_13423,N_12646);
or U14587 (N_14587,N_12580,N_12596);
nor U14588 (N_14588,N_12885,N_12111);
nand U14589 (N_14589,N_13390,N_13175);
xor U14590 (N_14590,N_13111,N_13414);
and U14591 (N_14591,N_12432,N_12143);
or U14592 (N_14592,N_12299,N_12672);
or U14593 (N_14593,N_13196,N_12280);
nor U14594 (N_14594,N_12958,N_13219);
xnor U14595 (N_14595,N_12177,N_13878);
or U14596 (N_14596,N_13170,N_12447);
xor U14597 (N_14597,N_13268,N_12094);
or U14598 (N_14598,N_12515,N_13058);
or U14599 (N_14599,N_12455,N_12680);
or U14600 (N_14600,N_12264,N_12735);
nand U14601 (N_14601,N_12849,N_13686);
nor U14602 (N_14602,N_12864,N_12484);
nand U14603 (N_14603,N_13002,N_13117);
or U14604 (N_14604,N_13047,N_13601);
and U14605 (N_14605,N_12208,N_13381);
nor U14606 (N_14606,N_12664,N_12791);
nand U14607 (N_14607,N_13384,N_13847);
nand U14608 (N_14608,N_13833,N_13560);
nand U14609 (N_14609,N_13029,N_12153);
xor U14610 (N_14610,N_12662,N_13806);
xor U14611 (N_14611,N_12719,N_13402);
xor U14612 (N_14612,N_13603,N_13814);
and U14613 (N_14613,N_13856,N_13664);
xor U14614 (N_14614,N_13368,N_13189);
xnor U14615 (N_14615,N_12572,N_13083);
xnor U14616 (N_14616,N_13750,N_13075);
nand U14617 (N_14617,N_12829,N_13638);
and U14618 (N_14618,N_12959,N_12659);
nor U14619 (N_14619,N_12883,N_12705);
and U14620 (N_14620,N_12222,N_12441);
or U14621 (N_14621,N_12016,N_13533);
or U14622 (N_14622,N_12159,N_12426);
or U14623 (N_14623,N_13257,N_13725);
xnor U14624 (N_14624,N_13835,N_12293);
and U14625 (N_14625,N_12727,N_12493);
and U14626 (N_14626,N_13514,N_13042);
and U14627 (N_14627,N_13483,N_12263);
xnor U14628 (N_14628,N_12311,N_12335);
and U14629 (N_14629,N_12737,N_13955);
nand U14630 (N_14630,N_12966,N_13255);
xor U14631 (N_14631,N_12451,N_12971);
xnor U14632 (N_14632,N_12656,N_13273);
or U14633 (N_14633,N_12539,N_12330);
nand U14634 (N_14634,N_12601,N_12304);
nand U14635 (N_14635,N_13890,N_13352);
or U14636 (N_14636,N_12900,N_12346);
nand U14637 (N_14637,N_12392,N_12009);
nand U14638 (N_14638,N_12049,N_13636);
and U14639 (N_14639,N_13485,N_13343);
or U14640 (N_14640,N_13547,N_13275);
xor U14641 (N_14641,N_13290,N_12960);
or U14642 (N_14642,N_13224,N_12977);
nor U14643 (N_14643,N_13495,N_13754);
xor U14644 (N_14644,N_13647,N_12808);
and U14645 (N_14645,N_12547,N_12691);
nand U14646 (N_14646,N_13177,N_12067);
xor U14647 (N_14647,N_13260,N_13190);
nand U14648 (N_14648,N_13619,N_13369);
xnor U14649 (N_14649,N_12577,N_13220);
and U14650 (N_14650,N_12151,N_12625);
nand U14651 (N_14651,N_13569,N_13309);
and U14652 (N_14652,N_13779,N_13938);
nand U14653 (N_14653,N_13266,N_13887);
nand U14654 (N_14654,N_13125,N_13271);
and U14655 (N_14655,N_12573,N_12375);
and U14656 (N_14656,N_12109,N_13081);
nand U14657 (N_14657,N_13332,N_12728);
xor U14658 (N_14658,N_12261,N_12742);
and U14659 (N_14659,N_13104,N_13845);
nor U14660 (N_14660,N_13836,N_12985);
or U14661 (N_14661,N_12905,N_13666);
xor U14662 (N_14662,N_12566,N_13416);
nor U14663 (N_14663,N_12754,N_13325);
and U14664 (N_14664,N_13663,N_12028);
or U14665 (N_14665,N_13631,N_12969);
nor U14666 (N_14666,N_12769,N_13067);
nor U14667 (N_14667,N_13519,N_12035);
nand U14668 (N_14668,N_13552,N_12136);
xnor U14669 (N_14669,N_12835,N_12044);
and U14670 (N_14670,N_12921,N_12195);
or U14671 (N_14671,N_13145,N_12811);
xnor U14672 (N_14672,N_13064,N_13975);
nor U14673 (N_14673,N_12692,N_13797);
nor U14674 (N_14674,N_12238,N_13407);
and U14675 (N_14675,N_12989,N_12106);
xor U14676 (N_14676,N_12689,N_12749);
or U14677 (N_14677,N_13248,N_13598);
and U14678 (N_14678,N_13251,N_13066);
or U14679 (N_14679,N_13470,N_12437);
nand U14680 (N_14680,N_12478,N_12467);
nand U14681 (N_14681,N_12907,N_13749);
nor U14682 (N_14682,N_12746,N_13329);
nor U14683 (N_14683,N_13559,N_12777);
and U14684 (N_14684,N_12168,N_12296);
nand U14685 (N_14685,N_13680,N_12752);
nand U14686 (N_14686,N_13939,N_12152);
nor U14687 (N_14687,N_13312,N_12133);
or U14688 (N_14688,N_12936,N_12538);
or U14689 (N_14689,N_12481,N_13830);
xnor U14690 (N_14690,N_13099,N_12262);
nor U14691 (N_14691,N_12788,N_13761);
nand U14692 (N_14692,N_13045,N_12803);
xor U14693 (N_14693,N_13623,N_13612);
or U14694 (N_14694,N_13063,N_13568);
xnor U14695 (N_14695,N_13230,N_12474);
and U14696 (N_14696,N_13948,N_12503);
nand U14697 (N_14697,N_12060,N_12453);
nand U14698 (N_14698,N_12031,N_12089);
and U14699 (N_14699,N_13853,N_13659);
nand U14700 (N_14700,N_13094,N_13361);
and U14701 (N_14701,N_12424,N_13319);
nor U14702 (N_14702,N_12072,N_13311);
xor U14703 (N_14703,N_13503,N_12618);
nand U14704 (N_14704,N_13076,N_13821);
nor U14705 (N_14705,N_13043,N_13386);
nand U14706 (N_14706,N_13089,N_13892);
nor U14707 (N_14707,N_12543,N_12778);
and U14708 (N_14708,N_12247,N_13116);
xnor U14709 (N_14709,N_13770,N_12234);
or U14710 (N_14710,N_13207,N_12124);
xnor U14711 (N_14711,N_12366,N_13996);
xor U14712 (N_14712,N_12828,N_12047);
nor U14713 (N_14713,N_12800,N_12897);
xnor U14714 (N_14714,N_13393,N_12995);
or U14715 (N_14715,N_12563,N_13281);
and U14716 (N_14716,N_13571,N_12326);
nor U14717 (N_14717,N_13752,N_12078);
nand U14718 (N_14718,N_13914,N_13550);
xor U14719 (N_14719,N_13385,N_12553);
nand U14720 (N_14720,N_12821,N_13600);
xor U14721 (N_14721,N_12411,N_13360);
or U14722 (N_14722,N_13985,N_13199);
and U14723 (N_14723,N_13694,N_12686);
nand U14724 (N_14724,N_13954,N_13300);
nor U14725 (N_14725,N_13760,N_12753);
or U14726 (N_14726,N_12276,N_13007);
nand U14727 (N_14727,N_12660,N_13183);
nand U14728 (N_14728,N_13229,N_13147);
nand U14729 (N_14729,N_13399,N_12589);
or U14730 (N_14730,N_12974,N_12161);
nor U14731 (N_14731,N_12776,N_13452);
nor U14732 (N_14732,N_13781,N_13363);
nor U14733 (N_14733,N_13542,N_13621);
xor U14734 (N_14734,N_12649,N_13724);
xor U14735 (N_14735,N_13777,N_13025);
and U14736 (N_14736,N_13697,N_12528);
nor U14737 (N_14737,N_13855,N_13707);
xor U14738 (N_14738,N_13895,N_12472);
and U14739 (N_14739,N_12599,N_12221);
nor U14740 (N_14740,N_13150,N_13491);
nand U14741 (N_14741,N_12270,N_13108);
or U14742 (N_14742,N_13347,N_13537);
nor U14743 (N_14743,N_13221,N_12418);
nand U14744 (N_14744,N_12502,N_12213);
nor U14745 (N_14745,N_13113,N_13245);
and U14746 (N_14746,N_12257,N_12405);
xor U14747 (N_14747,N_13069,N_12012);
xor U14748 (N_14748,N_13086,N_13340);
nand U14749 (N_14749,N_12703,N_13475);
and U14750 (N_14750,N_12476,N_12694);
nand U14751 (N_14751,N_13875,N_13851);
nand U14752 (N_14752,N_12137,N_12246);
or U14753 (N_14753,N_12822,N_12157);
or U14754 (N_14754,N_12410,N_12714);
or U14755 (N_14755,N_13511,N_12762);
nand U14756 (N_14756,N_12005,N_12868);
or U14757 (N_14757,N_12802,N_12915);
nor U14758 (N_14758,N_13711,N_13408);
or U14759 (N_14759,N_13652,N_12325);
xor U14760 (N_14760,N_12081,N_12357);
or U14761 (N_14761,N_12233,N_13173);
xnor U14762 (N_14762,N_13037,N_12427);
nand U14763 (N_14763,N_13941,N_13625);
xor U14764 (N_14764,N_13786,N_13604);
nor U14765 (N_14765,N_13307,N_12933);
and U14766 (N_14766,N_12250,N_13010);
xor U14767 (N_14767,N_12074,N_12945);
and U14768 (N_14768,N_12620,N_12978);
and U14769 (N_14769,N_13436,N_12093);
nor U14770 (N_14770,N_13449,N_12911);
xnor U14771 (N_14771,N_13417,N_13371);
nor U14772 (N_14772,N_13563,N_12452);
nor U14773 (N_14773,N_13060,N_12086);
and U14774 (N_14774,N_12704,N_13667);
or U14775 (N_14775,N_13223,N_13129);
nand U14776 (N_14776,N_12940,N_12767);
nor U14777 (N_14777,N_13592,N_12870);
xor U14778 (N_14778,N_13556,N_13349);
and U14779 (N_14779,N_12393,N_13087);
or U14780 (N_14780,N_13668,N_12908);
or U14781 (N_14781,N_12507,N_13734);
and U14782 (N_14782,N_12858,N_12104);
xnor U14783 (N_14783,N_13653,N_12214);
and U14784 (N_14784,N_13027,N_12770);
nand U14785 (N_14785,N_12929,N_13054);
xor U14786 (N_14786,N_12913,N_13593);
and U14787 (N_14787,N_13774,N_12015);
nand U14788 (N_14788,N_12710,N_13727);
xor U14789 (N_14789,N_13357,N_13387);
and U14790 (N_14790,N_13339,N_12850);
or U14791 (N_14791,N_12095,N_13997);
or U14792 (N_14792,N_13457,N_12551);
nor U14793 (N_14793,N_12674,N_13100);
and U14794 (N_14794,N_12926,N_12623);
or U14795 (N_14795,N_12061,N_13176);
nor U14796 (N_14796,N_12766,N_13061);
xnor U14797 (N_14797,N_12988,N_12292);
and U14798 (N_14798,N_12297,N_12533);
nand U14799 (N_14799,N_13676,N_12792);
nor U14800 (N_14800,N_12602,N_12063);
or U14801 (N_14801,N_12639,N_13809);
xnor U14802 (N_14802,N_13672,N_12621);
nand U14803 (N_14803,N_13249,N_12082);
and U14804 (N_14804,N_12362,N_12146);
or U14805 (N_14805,N_12398,N_12696);
nor U14806 (N_14806,N_12266,N_13000);
nand U14807 (N_14807,N_12189,N_13461);
or U14808 (N_14808,N_13059,N_13159);
or U14809 (N_14809,N_13301,N_12209);
or U14810 (N_14810,N_12758,N_13736);
xor U14811 (N_14811,N_13238,N_12267);
or U14812 (N_14812,N_12744,N_13586);
nor U14813 (N_14813,N_13981,N_13282);
nor U14814 (N_14814,N_12584,N_13460);
and U14815 (N_14815,N_12747,N_13004);
and U14816 (N_14816,N_13876,N_12824);
and U14817 (N_14817,N_12720,N_13429);
or U14818 (N_14818,N_12698,N_13949);
xor U14819 (N_14819,N_12170,N_13923);
xor U14820 (N_14820,N_13824,N_13730);
nor U14821 (N_14821,N_13607,N_12633);
xor U14822 (N_14822,N_13348,N_13733);
nor U14823 (N_14823,N_12898,N_12906);
or U14824 (N_14824,N_13299,N_12523);
or U14825 (N_14825,N_13082,N_13359);
and U14826 (N_14826,N_12199,N_12071);
xor U14827 (N_14827,N_12895,N_13964);
xor U14828 (N_14828,N_12848,N_13966);
xnor U14829 (N_14829,N_12857,N_12994);
or U14830 (N_14830,N_13788,N_13849);
or U14831 (N_14831,N_12930,N_12901);
xor U14832 (N_14832,N_12470,N_12903);
nor U14833 (N_14833,N_12768,N_12331);
nor U14834 (N_14834,N_13731,N_13532);
or U14835 (N_14835,N_13723,N_12018);
nand U14836 (N_14836,N_12185,N_13294);
nand U14837 (N_14837,N_13968,N_13804);
or U14838 (N_14838,N_13487,N_13062);
nor U14839 (N_14839,N_12433,N_12025);
xor U14840 (N_14840,N_12875,N_13812);
or U14841 (N_14841,N_12495,N_12525);
xnor U14842 (N_14842,N_13787,N_12351);
xnor U14843 (N_14843,N_12973,N_13389);
nor U14844 (N_14844,N_13077,N_13132);
xor U14845 (N_14845,N_12967,N_12600);
xor U14846 (N_14846,N_12003,N_13056);
xor U14847 (N_14847,N_12057,N_13976);
nor U14848 (N_14848,N_12167,N_12722);
and U14849 (N_14849,N_12217,N_13643);
and U14850 (N_14850,N_13297,N_13990);
and U14851 (N_14851,N_13130,N_13437);
nand U14852 (N_14852,N_12309,N_12715);
and U14853 (N_14853,N_13122,N_13333);
or U14854 (N_14854,N_13166,N_12300);
nor U14855 (N_14855,N_12388,N_13622);
nor U14856 (N_14856,N_12902,N_13472);
nor U14857 (N_14857,N_13492,N_12666);
and U14858 (N_14858,N_12716,N_13068);
nand U14859 (N_14859,N_13893,N_12708);
or U14860 (N_14860,N_12984,N_12663);
xnor U14861 (N_14861,N_12373,N_12650);
xnor U14862 (N_14862,N_12560,N_12117);
and U14863 (N_14863,N_12370,N_12210);
nand U14864 (N_14864,N_13209,N_12771);
and U14865 (N_14865,N_12290,N_12041);
and U14866 (N_14866,N_13451,N_13454);
nand U14867 (N_14867,N_12401,N_13688);
nor U14868 (N_14868,N_13296,N_13443);
and U14869 (N_14869,N_13036,N_13589);
xor U14870 (N_14870,N_12871,N_12198);
xor U14871 (N_14871,N_13411,N_12457);
and U14872 (N_14872,N_12036,N_13561);
nor U14873 (N_14873,N_12608,N_12113);
xor U14874 (N_14874,N_13641,N_13272);
nand U14875 (N_14875,N_13848,N_12847);
and U14876 (N_14876,N_13915,N_13203);
nand U14877 (N_14877,N_13767,N_13819);
or U14878 (N_14878,N_12939,N_12205);
xor U14879 (N_14879,N_13591,N_13758);
nand U14880 (N_14880,N_12643,N_12590);
nor U14881 (N_14881,N_13049,N_12492);
nor U14882 (N_14882,N_12101,N_13630);
xnor U14883 (N_14883,N_13742,N_12583);
or U14884 (N_14884,N_13261,N_13158);
or U14885 (N_14885,N_12568,N_13115);
nor U14886 (N_14886,N_13265,N_13420);
nand U14887 (N_14887,N_13950,N_12175);
and U14888 (N_14888,N_12361,N_13838);
nand U14889 (N_14889,N_13609,N_13034);
nor U14890 (N_14890,N_12496,N_12079);
and U14891 (N_14891,N_12313,N_12711);
xnor U14892 (N_14892,N_13822,N_13032);
nand U14893 (N_14893,N_13854,N_12368);
and U14894 (N_14894,N_13442,N_13031);
xnor U14895 (N_14895,N_13247,N_12687);
nor U14896 (N_14896,N_12923,N_13684);
nand U14897 (N_14897,N_12757,N_12229);
and U14898 (N_14898,N_12118,N_13620);
nor U14899 (N_14899,N_12034,N_13425);
xnor U14900 (N_14900,N_12683,N_13458);
xor U14901 (N_14901,N_12488,N_13546);
nor U14902 (N_14902,N_12567,N_12512);
nand U14903 (N_14903,N_12810,N_12129);
or U14904 (N_14904,N_12409,N_13241);
xnor U14905 (N_14905,N_12312,N_12342);
xor U14906 (N_14906,N_12833,N_13682);
nand U14907 (N_14907,N_13538,N_12397);
and U14908 (N_14908,N_13602,N_12148);
and U14909 (N_14909,N_12466,N_13566);
nor U14910 (N_14910,N_12732,N_13431);
and U14911 (N_14911,N_12851,N_13531);
xor U14912 (N_14912,N_13133,N_13583);
and U14913 (N_14913,N_12652,N_13481);
nor U14914 (N_14914,N_12894,N_13403);
nand U14915 (N_14915,N_13225,N_13590);
nand U14916 (N_14916,N_12853,N_13906);
xor U14917 (N_14917,N_13405,N_13946);
and U14918 (N_14918,N_12215,N_13073);
xor U14919 (N_14919,N_13683,N_13162);
xor U14920 (N_14920,N_13930,N_13198);
and U14921 (N_14921,N_13582,N_13197);
nor U14922 (N_14922,N_12127,N_12414);
and U14923 (N_14923,N_12191,N_13237);
nor U14924 (N_14924,N_13726,N_12141);
nor U14925 (N_14925,N_12423,N_13867);
and U14926 (N_14926,N_13114,N_13091);
or U14927 (N_14927,N_13080,N_12797);
or U14928 (N_14928,N_12400,N_13181);
nand U14929 (N_14929,N_13304,N_13818);
nor U14930 (N_14930,N_13090,N_13480);
and U14931 (N_14931,N_12278,N_13928);
nand U14932 (N_14932,N_13482,N_13107);
nor U14933 (N_14933,N_12707,N_12100);
nor U14934 (N_14934,N_12510,N_12001);
or U14935 (N_14935,N_12206,N_13507);
or U14936 (N_14936,N_13497,N_12352);
nor U14937 (N_14937,N_12070,N_12617);
or U14938 (N_14938,N_12500,N_13535);
nor U14939 (N_14939,N_12110,N_12529);
and U14940 (N_14940,N_13391,N_12996);
or U14941 (N_14941,N_12139,N_13270);
or U14942 (N_14942,N_13745,N_12592);
and U14943 (N_14943,N_12546,N_13003);
xnor U14944 (N_14944,N_12843,N_12975);
nor U14945 (N_14945,N_12236,N_12917);
nand U14946 (N_14946,N_13444,N_12115);
and U14947 (N_14947,N_13035,N_13314);
nor U14948 (N_14948,N_13512,N_12201);
or U14949 (N_14949,N_13832,N_13044);
xor U14950 (N_14950,N_12465,N_13446);
nand U14951 (N_14951,N_13921,N_13506);
xor U14952 (N_14952,N_13336,N_13508);
xnor U14953 (N_14953,N_12150,N_13763);
nor U14954 (N_14954,N_13585,N_13922);
nor U14955 (N_14955,N_12377,N_12718);
or U14956 (N_14956,N_13464,N_13337);
nand U14957 (N_14957,N_13378,N_12886);
xor U14958 (N_14958,N_12668,N_13557);
nand U14959 (N_14959,N_12353,N_13544);
xnor U14960 (N_14960,N_12819,N_12228);
or U14961 (N_14961,N_13345,N_12879);
nand U14962 (N_14962,N_12839,N_12212);
nand U14963 (N_14963,N_13211,N_13529);
xor U14964 (N_14964,N_12052,N_13719);
nor U14965 (N_14965,N_13692,N_12196);
nor U14966 (N_14966,N_12132,N_12033);
nor U14967 (N_14967,N_12661,N_13455);
nor U14968 (N_14968,N_12337,N_13331);
xnor U14969 (N_14969,N_13670,N_12790);
nand U14970 (N_14970,N_12816,N_12866);
and U14971 (N_14971,N_13999,N_13279);
and U14972 (N_14972,N_13793,N_13287);
nand U14973 (N_14973,N_13317,N_12532);
nand U14974 (N_14974,N_12925,N_13015);
xor U14975 (N_14975,N_13965,N_13404);
nand U14976 (N_14976,N_12702,N_12184);
and U14977 (N_14977,N_12327,N_12334);
xnor U14978 (N_14978,N_13447,N_12743);
or U14979 (N_14979,N_13611,N_12616);
nand U14980 (N_14980,N_12350,N_12693);
nand U14981 (N_14981,N_12904,N_12986);
and U14982 (N_14982,N_13989,N_13185);
or U14983 (N_14983,N_13200,N_12181);
xnor U14984 (N_14984,N_13143,N_13588);
nand U14985 (N_14985,N_12302,N_12164);
xnor U14986 (N_14986,N_12611,N_13808);
nand U14987 (N_14987,N_13904,N_12630);
nor U14988 (N_14988,N_13648,N_13341);
and U14989 (N_14989,N_12982,N_12192);
and U14990 (N_14990,N_12338,N_13618);
nor U14991 (N_14991,N_12180,N_12575);
nand U14992 (N_14992,N_12171,N_13899);
and U14993 (N_14993,N_13729,N_12108);
nand U14994 (N_14994,N_13743,N_13737);
or U14995 (N_14995,N_13328,N_12240);
nand U14996 (N_14996,N_13815,N_13658);
nor U14997 (N_14997,N_13816,N_13040);
nand U14998 (N_14998,N_12531,N_13910);
or U14999 (N_14999,N_12786,N_12881);
or U15000 (N_15000,N_13783,N_12476);
xor U15001 (N_15001,N_13392,N_13040);
and U15002 (N_15002,N_13158,N_13464);
and U15003 (N_15003,N_12042,N_13437);
and U15004 (N_15004,N_12632,N_12839);
or U15005 (N_15005,N_12602,N_12090);
xnor U15006 (N_15006,N_12627,N_12078);
xnor U15007 (N_15007,N_12040,N_13803);
and U15008 (N_15008,N_13293,N_13236);
nor U15009 (N_15009,N_13170,N_12652);
and U15010 (N_15010,N_13753,N_12304);
nor U15011 (N_15011,N_12700,N_12241);
nand U15012 (N_15012,N_13293,N_12575);
and U15013 (N_15013,N_13041,N_13331);
and U15014 (N_15014,N_13777,N_12516);
nand U15015 (N_15015,N_12213,N_13507);
nand U15016 (N_15016,N_13825,N_12836);
or U15017 (N_15017,N_13190,N_13176);
xor U15018 (N_15018,N_12080,N_13061);
and U15019 (N_15019,N_12791,N_12278);
nand U15020 (N_15020,N_13168,N_12199);
nor U15021 (N_15021,N_12652,N_13962);
nand U15022 (N_15022,N_12418,N_12071);
or U15023 (N_15023,N_12183,N_12728);
and U15024 (N_15024,N_12642,N_12366);
xor U15025 (N_15025,N_13585,N_12541);
xnor U15026 (N_15026,N_12939,N_13397);
xnor U15027 (N_15027,N_13573,N_13764);
nor U15028 (N_15028,N_13097,N_13974);
nand U15029 (N_15029,N_12627,N_13331);
xor U15030 (N_15030,N_13052,N_13967);
and U15031 (N_15031,N_13163,N_12422);
xor U15032 (N_15032,N_13990,N_13790);
or U15033 (N_15033,N_13028,N_12642);
and U15034 (N_15034,N_13772,N_13257);
nand U15035 (N_15035,N_12866,N_13680);
nand U15036 (N_15036,N_12892,N_13102);
nor U15037 (N_15037,N_12692,N_13973);
nor U15038 (N_15038,N_13594,N_12648);
or U15039 (N_15039,N_12178,N_13268);
nor U15040 (N_15040,N_12346,N_12497);
nor U15041 (N_15041,N_12790,N_12864);
or U15042 (N_15042,N_13042,N_12743);
xor U15043 (N_15043,N_13587,N_13066);
nand U15044 (N_15044,N_13746,N_12187);
xnor U15045 (N_15045,N_13755,N_13348);
nand U15046 (N_15046,N_12130,N_12029);
xnor U15047 (N_15047,N_13207,N_13215);
nor U15048 (N_15048,N_12401,N_12144);
or U15049 (N_15049,N_13214,N_12759);
xor U15050 (N_15050,N_12418,N_12345);
or U15051 (N_15051,N_12940,N_12942);
xnor U15052 (N_15052,N_13711,N_13494);
nand U15053 (N_15053,N_13242,N_12042);
nor U15054 (N_15054,N_13295,N_12095);
nor U15055 (N_15055,N_13843,N_12185);
xnor U15056 (N_15056,N_12105,N_13974);
xor U15057 (N_15057,N_12580,N_12024);
nor U15058 (N_15058,N_13485,N_13078);
nand U15059 (N_15059,N_12306,N_12974);
nand U15060 (N_15060,N_12150,N_12977);
nand U15061 (N_15061,N_13082,N_13583);
and U15062 (N_15062,N_13069,N_13668);
nor U15063 (N_15063,N_13409,N_13267);
nor U15064 (N_15064,N_12045,N_13213);
or U15065 (N_15065,N_13814,N_13010);
or U15066 (N_15066,N_13675,N_12047);
nor U15067 (N_15067,N_13423,N_13895);
xnor U15068 (N_15068,N_13898,N_13418);
or U15069 (N_15069,N_13546,N_12436);
or U15070 (N_15070,N_13072,N_13629);
and U15071 (N_15071,N_13172,N_13823);
nand U15072 (N_15072,N_13700,N_12394);
and U15073 (N_15073,N_12448,N_12128);
and U15074 (N_15074,N_13731,N_13163);
or U15075 (N_15075,N_13196,N_12091);
nor U15076 (N_15076,N_12169,N_12518);
nand U15077 (N_15077,N_12025,N_12620);
and U15078 (N_15078,N_12164,N_12993);
nand U15079 (N_15079,N_13442,N_12878);
nor U15080 (N_15080,N_12725,N_13100);
and U15081 (N_15081,N_12379,N_12694);
xnor U15082 (N_15082,N_12446,N_13844);
and U15083 (N_15083,N_13796,N_12782);
and U15084 (N_15084,N_12091,N_12848);
xor U15085 (N_15085,N_13353,N_12523);
nor U15086 (N_15086,N_12978,N_13420);
nor U15087 (N_15087,N_12886,N_12402);
and U15088 (N_15088,N_12289,N_12926);
nand U15089 (N_15089,N_12256,N_12538);
nand U15090 (N_15090,N_12086,N_13497);
xnor U15091 (N_15091,N_12127,N_12276);
nand U15092 (N_15092,N_12954,N_12096);
or U15093 (N_15093,N_12280,N_13338);
nand U15094 (N_15094,N_12143,N_13241);
and U15095 (N_15095,N_13650,N_13659);
nand U15096 (N_15096,N_12371,N_12205);
xor U15097 (N_15097,N_12156,N_13386);
nor U15098 (N_15098,N_13930,N_13065);
xor U15099 (N_15099,N_13766,N_13380);
nand U15100 (N_15100,N_13357,N_13814);
nor U15101 (N_15101,N_12744,N_12394);
nand U15102 (N_15102,N_12161,N_13801);
xnor U15103 (N_15103,N_12765,N_13268);
or U15104 (N_15104,N_12706,N_12397);
xnor U15105 (N_15105,N_13260,N_12629);
nand U15106 (N_15106,N_13251,N_12202);
and U15107 (N_15107,N_12135,N_12957);
xnor U15108 (N_15108,N_13120,N_13839);
and U15109 (N_15109,N_12994,N_12044);
nand U15110 (N_15110,N_13484,N_13228);
xnor U15111 (N_15111,N_12615,N_13401);
or U15112 (N_15112,N_13267,N_13519);
nor U15113 (N_15113,N_12886,N_13415);
or U15114 (N_15114,N_13573,N_13599);
nor U15115 (N_15115,N_12033,N_13959);
xnor U15116 (N_15116,N_13183,N_12849);
nand U15117 (N_15117,N_12946,N_12065);
nand U15118 (N_15118,N_12051,N_12102);
nor U15119 (N_15119,N_13940,N_13320);
nor U15120 (N_15120,N_13321,N_12220);
nor U15121 (N_15121,N_12966,N_12914);
and U15122 (N_15122,N_13053,N_12439);
and U15123 (N_15123,N_12613,N_13118);
xor U15124 (N_15124,N_13313,N_12991);
and U15125 (N_15125,N_13973,N_12506);
and U15126 (N_15126,N_12878,N_13944);
nor U15127 (N_15127,N_12826,N_12478);
nor U15128 (N_15128,N_12952,N_13507);
and U15129 (N_15129,N_13317,N_12437);
xor U15130 (N_15130,N_12602,N_13349);
xor U15131 (N_15131,N_12362,N_12928);
and U15132 (N_15132,N_12314,N_12762);
nand U15133 (N_15133,N_12940,N_12615);
nor U15134 (N_15134,N_13080,N_13689);
and U15135 (N_15135,N_13972,N_12303);
nor U15136 (N_15136,N_13075,N_12234);
and U15137 (N_15137,N_13689,N_12880);
xor U15138 (N_15138,N_12631,N_12200);
nor U15139 (N_15139,N_13284,N_12467);
xor U15140 (N_15140,N_13556,N_12712);
or U15141 (N_15141,N_13399,N_12277);
nor U15142 (N_15142,N_13352,N_12669);
nor U15143 (N_15143,N_12853,N_13567);
nand U15144 (N_15144,N_12714,N_12417);
and U15145 (N_15145,N_12767,N_13629);
or U15146 (N_15146,N_13921,N_12019);
xnor U15147 (N_15147,N_13780,N_13152);
nand U15148 (N_15148,N_13038,N_12843);
or U15149 (N_15149,N_13043,N_12570);
nand U15150 (N_15150,N_12944,N_13570);
and U15151 (N_15151,N_12440,N_13491);
and U15152 (N_15152,N_13238,N_12843);
nand U15153 (N_15153,N_12751,N_12534);
nand U15154 (N_15154,N_12927,N_12783);
xnor U15155 (N_15155,N_13463,N_13417);
or U15156 (N_15156,N_13933,N_12680);
and U15157 (N_15157,N_12736,N_12883);
nand U15158 (N_15158,N_12886,N_13386);
nor U15159 (N_15159,N_13274,N_12669);
or U15160 (N_15160,N_12292,N_13664);
or U15161 (N_15161,N_12133,N_13337);
or U15162 (N_15162,N_12406,N_13344);
nor U15163 (N_15163,N_13163,N_13634);
and U15164 (N_15164,N_13560,N_12649);
or U15165 (N_15165,N_13105,N_13286);
nor U15166 (N_15166,N_12476,N_13705);
or U15167 (N_15167,N_12296,N_12929);
nand U15168 (N_15168,N_12809,N_13918);
nor U15169 (N_15169,N_13432,N_12163);
xor U15170 (N_15170,N_12962,N_12997);
or U15171 (N_15171,N_12917,N_12528);
or U15172 (N_15172,N_13663,N_13093);
nor U15173 (N_15173,N_13164,N_12473);
nand U15174 (N_15174,N_13342,N_12669);
xor U15175 (N_15175,N_12106,N_12844);
and U15176 (N_15176,N_12995,N_12021);
nand U15177 (N_15177,N_13508,N_12623);
nand U15178 (N_15178,N_13729,N_13816);
or U15179 (N_15179,N_13686,N_12268);
or U15180 (N_15180,N_13883,N_13235);
nand U15181 (N_15181,N_13056,N_13287);
nor U15182 (N_15182,N_13171,N_12980);
xnor U15183 (N_15183,N_13164,N_13379);
xor U15184 (N_15184,N_12825,N_12715);
and U15185 (N_15185,N_13425,N_12097);
xnor U15186 (N_15186,N_12460,N_13512);
and U15187 (N_15187,N_13631,N_12277);
xnor U15188 (N_15188,N_12442,N_12659);
nor U15189 (N_15189,N_13901,N_12373);
nor U15190 (N_15190,N_12705,N_13199);
xor U15191 (N_15191,N_13800,N_13815);
xor U15192 (N_15192,N_12717,N_13819);
and U15193 (N_15193,N_13873,N_12750);
nand U15194 (N_15194,N_12269,N_12435);
xnor U15195 (N_15195,N_12602,N_12263);
nand U15196 (N_15196,N_13320,N_13411);
nand U15197 (N_15197,N_12557,N_13346);
nand U15198 (N_15198,N_12693,N_12566);
xnor U15199 (N_15199,N_12328,N_12190);
nand U15200 (N_15200,N_13258,N_12419);
xor U15201 (N_15201,N_13869,N_13452);
or U15202 (N_15202,N_13816,N_12710);
and U15203 (N_15203,N_13621,N_12593);
or U15204 (N_15204,N_13933,N_12945);
or U15205 (N_15205,N_12509,N_12103);
nor U15206 (N_15206,N_13476,N_13503);
and U15207 (N_15207,N_13061,N_13914);
xor U15208 (N_15208,N_12143,N_12257);
and U15209 (N_15209,N_13358,N_12925);
nand U15210 (N_15210,N_12211,N_12255);
nand U15211 (N_15211,N_12321,N_13789);
and U15212 (N_15212,N_13249,N_12937);
or U15213 (N_15213,N_12657,N_13995);
or U15214 (N_15214,N_12144,N_13798);
nand U15215 (N_15215,N_13529,N_12768);
nand U15216 (N_15216,N_13817,N_12243);
nor U15217 (N_15217,N_12381,N_12925);
nand U15218 (N_15218,N_12640,N_13566);
or U15219 (N_15219,N_13602,N_13941);
nand U15220 (N_15220,N_12719,N_12317);
and U15221 (N_15221,N_13743,N_12747);
nand U15222 (N_15222,N_13022,N_13334);
nor U15223 (N_15223,N_13985,N_12296);
nor U15224 (N_15224,N_12758,N_13856);
xnor U15225 (N_15225,N_12462,N_13637);
nor U15226 (N_15226,N_12963,N_13498);
or U15227 (N_15227,N_12184,N_12354);
and U15228 (N_15228,N_12728,N_12537);
nand U15229 (N_15229,N_12057,N_12413);
and U15230 (N_15230,N_12682,N_13283);
nor U15231 (N_15231,N_13826,N_12903);
xor U15232 (N_15232,N_12881,N_12013);
nand U15233 (N_15233,N_12022,N_12709);
or U15234 (N_15234,N_13856,N_12284);
xnor U15235 (N_15235,N_13075,N_13668);
nor U15236 (N_15236,N_13389,N_12953);
nand U15237 (N_15237,N_12165,N_13959);
or U15238 (N_15238,N_13950,N_12909);
or U15239 (N_15239,N_13159,N_13275);
and U15240 (N_15240,N_12791,N_12957);
nor U15241 (N_15241,N_13349,N_12803);
xnor U15242 (N_15242,N_12054,N_12582);
nand U15243 (N_15243,N_12308,N_13649);
and U15244 (N_15244,N_12984,N_12554);
nor U15245 (N_15245,N_12323,N_12566);
xnor U15246 (N_15246,N_12417,N_13263);
xnor U15247 (N_15247,N_12883,N_13028);
and U15248 (N_15248,N_13454,N_12799);
xor U15249 (N_15249,N_12089,N_12767);
or U15250 (N_15250,N_13064,N_12243);
or U15251 (N_15251,N_13451,N_12514);
nor U15252 (N_15252,N_13765,N_12170);
or U15253 (N_15253,N_13397,N_13411);
nand U15254 (N_15254,N_13255,N_12990);
and U15255 (N_15255,N_13130,N_13560);
nand U15256 (N_15256,N_13173,N_12653);
or U15257 (N_15257,N_13726,N_12959);
xnor U15258 (N_15258,N_12203,N_12069);
nand U15259 (N_15259,N_13933,N_13842);
and U15260 (N_15260,N_12897,N_12491);
nor U15261 (N_15261,N_13721,N_13773);
nand U15262 (N_15262,N_13242,N_13381);
and U15263 (N_15263,N_13989,N_13378);
nand U15264 (N_15264,N_12770,N_13713);
and U15265 (N_15265,N_13977,N_13179);
nand U15266 (N_15266,N_12059,N_12408);
xor U15267 (N_15267,N_12856,N_12994);
and U15268 (N_15268,N_12304,N_13224);
and U15269 (N_15269,N_13149,N_13780);
or U15270 (N_15270,N_13030,N_12859);
nor U15271 (N_15271,N_12824,N_13602);
nor U15272 (N_15272,N_12027,N_13472);
and U15273 (N_15273,N_13061,N_13036);
xor U15274 (N_15274,N_13585,N_13171);
nor U15275 (N_15275,N_12004,N_13725);
or U15276 (N_15276,N_13996,N_12922);
and U15277 (N_15277,N_12648,N_13465);
xor U15278 (N_15278,N_13356,N_12792);
and U15279 (N_15279,N_12979,N_12557);
nor U15280 (N_15280,N_13335,N_13531);
or U15281 (N_15281,N_13914,N_12814);
nor U15282 (N_15282,N_13798,N_12504);
and U15283 (N_15283,N_12339,N_12164);
nand U15284 (N_15284,N_13068,N_12999);
nor U15285 (N_15285,N_12166,N_12985);
and U15286 (N_15286,N_13832,N_12899);
xnor U15287 (N_15287,N_13684,N_13680);
nand U15288 (N_15288,N_13180,N_13499);
and U15289 (N_15289,N_13256,N_12597);
xor U15290 (N_15290,N_13226,N_12946);
xnor U15291 (N_15291,N_13814,N_13311);
or U15292 (N_15292,N_13198,N_12796);
nor U15293 (N_15293,N_13770,N_13672);
nor U15294 (N_15294,N_13196,N_12636);
xor U15295 (N_15295,N_13041,N_13360);
nor U15296 (N_15296,N_13123,N_13325);
nor U15297 (N_15297,N_12642,N_13735);
xnor U15298 (N_15298,N_13624,N_12995);
xnor U15299 (N_15299,N_13834,N_12259);
xnor U15300 (N_15300,N_13346,N_12723);
nor U15301 (N_15301,N_12333,N_13665);
xor U15302 (N_15302,N_13496,N_13936);
nand U15303 (N_15303,N_13556,N_12561);
and U15304 (N_15304,N_13393,N_12749);
nor U15305 (N_15305,N_12848,N_12027);
nor U15306 (N_15306,N_12884,N_13984);
and U15307 (N_15307,N_13017,N_13301);
and U15308 (N_15308,N_13402,N_12240);
and U15309 (N_15309,N_12920,N_12704);
nor U15310 (N_15310,N_13794,N_12807);
nand U15311 (N_15311,N_12510,N_13470);
and U15312 (N_15312,N_13278,N_12533);
and U15313 (N_15313,N_13194,N_12070);
or U15314 (N_15314,N_13396,N_12386);
or U15315 (N_15315,N_13256,N_13753);
nand U15316 (N_15316,N_12499,N_12595);
xor U15317 (N_15317,N_13250,N_12610);
xnor U15318 (N_15318,N_13918,N_12862);
xnor U15319 (N_15319,N_13108,N_12370);
nand U15320 (N_15320,N_13884,N_12478);
nor U15321 (N_15321,N_13835,N_12055);
nand U15322 (N_15322,N_12718,N_13936);
nor U15323 (N_15323,N_12760,N_13040);
xnor U15324 (N_15324,N_12186,N_13595);
xor U15325 (N_15325,N_13882,N_12345);
and U15326 (N_15326,N_13281,N_12592);
nor U15327 (N_15327,N_12701,N_12178);
nor U15328 (N_15328,N_13703,N_13331);
or U15329 (N_15329,N_12712,N_13690);
nor U15330 (N_15330,N_13140,N_13774);
or U15331 (N_15331,N_12881,N_13893);
nor U15332 (N_15332,N_13620,N_13017);
and U15333 (N_15333,N_13375,N_12197);
and U15334 (N_15334,N_12949,N_12759);
xnor U15335 (N_15335,N_12247,N_13261);
xor U15336 (N_15336,N_13158,N_13996);
nand U15337 (N_15337,N_12181,N_12478);
nand U15338 (N_15338,N_12376,N_12531);
or U15339 (N_15339,N_12637,N_13315);
or U15340 (N_15340,N_12035,N_13030);
nand U15341 (N_15341,N_13503,N_12761);
nor U15342 (N_15342,N_12727,N_13515);
or U15343 (N_15343,N_13093,N_13732);
and U15344 (N_15344,N_13346,N_12716);
nor U15345 (N_15345,N_13529,N_12821);
and U15346 (N_15346,N_12675,N_12692);
xor U15347 (N_15347,N_13837,N_13509);
xor U15348 (N_15348,N_13649,N_13086);
nor U15349 (N_15349,N_13329,N_12014);
nand U15350 (N_15350,N_13756,N_12175);
nor U15351 (N_15351,N_12660,N_12451);
xor U15352 (N_15352,N_13512,N_12071);
xnor U15353 (N_15353,N_12534,N_13793);
or U15354 (N_15354,N_12090,N_13889);
xnor U15355 (N_15355,N_13596,N_13180);
nand U15356 (N_15356,N_13936,N_13998);
or U15357 (N_15357,N_12592,N_13153);
nor U15358 (N_15358,N_12640,N_12838);
nand U15359 (N_15359,N_12452,N_13571);
nand U15360 (N_15360,N_12119,N_12273);
nor U15361 (N_15361,N_12102,N_13658);
and U15362 (N_15362,N_13888,N_13858);
nor U15363 (N_15363,N_12125,N_13743);
and U15364 (N_15364,N_12483,N_12260);
and U15365 (N_15365,N_12254,N_12214);
xnor U15366 (N_15366,N_13752,N_13210);
nor U15367 (N_15367,N_12427,N_12866);
xnor U15368 (N_15368,N_13789,N_12255);
nor U15369 (N_15369,N_12755,N_13617);
nand U15370 (N_15370,N_12470,N_13620);
and U15371 (N_15371,N_12559,N_12259);
xnor U15372 (N_15372,N_13669,N_13787);
or U15373 (N_15373,N_12264,N_12145);
nand U15374 (N_15374,N_13552,N_13490);
or U15375 (N_15375,N_13844,N_13188);
and U15376 (N_15376,N_12737,N_13416);
and U15377 (N_15377,N_12997,N_12037);
nor U15378 (N_15378,N_13050,N_13313);
and U15379 (N_15379,N_12085,N_13775);
or U15380 (N_15380,N_13809,N_12026);
and U15381 (N_15381,N_12388,N_13275);
or U15382 (N_15382,N_13200,N_13594);
and U15383 (N_15383,N_13308,N_12671);
xor U15384 (N_15384,N_13795,N_12241);
and U15385 (N_15385,N_13407,N_12492);
nor U15386 (N_15386,N_13926,N_13352);
and U15387 (N_15387,N_12241,N_12077);
nor U15388 (N_15388,N_12434,N_13004);
and U15389 (N_15389,N_12937,N_13429);
or U15390 (N_15390,N_13711,N_12943);
or U15391 (N_15391,N_13232,N_13169);
xnor U15392 (N_15392,N_12720,N_12978);
or U15393 (N_15393,N_12797,N_13089);
nor U15394 (N_15394,N_12508,N_13344);
nand U15395 (N_15395,N_13314,N_12151);
xor U15396 (N_15396,N_12275,N_13647);
nor U15397 (N_15397,N_12295,N_12545);
and U15398 (N_15398,N_12087,N_12043);
nand U15399 (N_15399,N_13919,N_12074);
xnor U15400 (N_15400,N_12397,N_13164);
nand U15401 (N_15401,N_12878,N_12496);
or U15402 (N_15402,N_13117,N_13339);
and U15403 (N_15403,N_13772,N_13153);
or U15404 (N_15404,N_12980,N_13204);
xnor U15405 (N_15405,N_13289,N_12124);
and U15406 (N_15406,N_12529,N_13291);
nor U15407 (N_15407,N_13793,N_12208);
xnor U15408 (N_15408,N_13886,N_12480);
or U15409 (N_15409,N_13672,N_13495);
and U15410 (N_15410,N_12226,N_13427);
or U15411 (N_15411,N_12316,N_13828);
xor U15412 (N_15412,N_13093,N_13443);
or U15413 (N_15413,N_13232,N_13793);
nor U15414 (N_15414,N_13843,N_13790);
or U15415 (N_15415,N_12453,N_12999);
or U15416 (N_15416,N_13047,N_13705);
or U15417 (N_15417,N_13175,N_12856);
and U15418 (N_15418,N_13733,N_13597);
and U15419 (N_15419,N_13800,N_12303);
or U15420 (N_15420,N_13627,N_13832);
or U15421 (N_15421,N_13922,N_12298);
xnor U15422 (N_15422,N_13998,N_13121);
nand U15423 (N_15423,N_12372,N_13647);
nor U15424 (N_15424,N_13944,N_12840);
nand U15425 (N_15425,N_12283,N_12724);
nand U15426 (N_15426,N_13334,N_13161);
nand U15427 (N_15427,N_12758,N_13674);
or U15428 (N_15428,N_12414,N_12483);
xor U15429 (N_15429,N_12869,N_13562);
nor U15430 (N_15430,N_13428,N_13349);
xnor U15431 (N_15431,N_13593,N_12795);
nor U15432 (N_15432,N_12687,N_12230);
or U15433 (N_15433,N_13987,N_13469);
xnor U15434 (N_15434,N_12708,N_12169);
or U15435 (N_15435,N_13589,N_12626);
and U15436 (N_15436,N_12971,N_13087);
xor U15437 (N_15437,N_12517,N_12658);
and U15438 (N_15438,N_13839,N_12588);
nor U15439 (N_15439,N_12263,N_13952);
nand U15440 (N_15440,N_13693,N_13298);
and U15441 (N_15441,N_13894,N_12779);
nand U15442 (N_15442,N_12125,N_13058);
and U15443 (N_15443,N_12386,N_12184);
or U15444 (N_15444,N_13014,N_12468);
or U15445 (N_15445,N_12396,N_13588);
nand U15446 (N_15446,N_12528,N_12665);
and U15447 (N_15447,N_12904,N_13951);
xor U15448 (N_15448,N_12183,N_12755);
nand U15449 (N_15449,N_12821,N_12105);
or U15450 (N_15450,N_13266,N_13530);
nand U15451 (N_15451,N_13728,N_12713);
nor U15452 (N_15452,N_12265,N_13281);
and U15453 (N_15453,N_12004,N_13324);
nand U15454 (N_15454,N_13342,N_12400);
nand U15455 (N_15455,N_13268,N_12474);
xnor U15456 (N_15456,N_13109,N_13612);
nand U15457 (N_15457,N_13463,N_13884);
or U15458 (N_15458,N_13966,N_12931);
nand U15459 (N_15459,N_12474,N_12981);
nand U15460 (N_15460,N_12164,N_12945);
or U15461 (N_15461,N_13272,N_12356);
and U15462 (N_15462,N_13580,N_13339);
or U15463 (N_15463,N_12149,N_13579);
xor U15464 (N_15464,N_13101,N_13059);
or U15465 (N_15465,N_13454,N_12703);
xor U15466 (N_15466,N_12889,N_12284);
nand U15467 (N_15467,N_13268,N_13729);
xnor U15468 (N_15468,N_12007,N_13642);
nor U15469 (N_15469,N_12224,N_13096);
or U15470 (N_15470,N_13185,N_12762);
or U15471 (N_15471,N_13660,N_13526);
nor U15472 (N_15472,N_13093,N_12739);
nand U15473 (N_15473,N_13940,N_12862);
xnor U15474 (N_15474,N_12170,N_12010);
xor U15475 (N_15475,N_12797,N_12954);
or U15476 (N_15476,N_12876,N_13854);
nor U15477 (N_15477,N_12468,N_12278);
and U15478 (N_15478,N_13474,N_12142);
and U15479 (N_15479,N_13254,N_13830);
or U15480 (N_15480,N_12680,N_12459);
xnor U15481 (N_15481,N_12039,N_13858);
nor U15482 (N_15482,N_13098,N_12902);
nand U15483 (N_15483,N_13911,N_12391);
xor U15484 (N_15484,N_12203,N_13411);
and U15485 (N_15485,N_13251,N_12058);
xor U15486 (N_15486,N_13733,N_13383);
or U15487 (N_15487,N_12913,N_13252);
nor U15488 (N_15488,N_12749,N_13817);
and U15489 (N_15489,N_12393,N_13503);
xnor U15490 (N_15490,N_12537,N_13773);
xnor U15491 (N_15491,N_13161,N_13396);
nand U15492 (N_15492,N_13963,N_13888);
xnor U15493 (N_15493,N_13237,N_12192);
and U15494 (N_15494,N_13365,N_12609);
xor U15495 (N_15495,N_12707,N_13438);
and U15496 (N_15496,N_13272,N_13263);
nor U15497 (N_15497,N_12938,N_13162);
xor U15498 (N_15498,N_13367,N_13214);
and U15499 (N_15499,N_13198,N_12493);
xnor U15500 (N_15500,N_12170,N_13397);
nor U15501 (N_15501,N_13242,N_13448);
nand U15502 (N_15502,N_12998,N_13976);
and U15503 (N_15503,N_13490,N_13844);
xnor U15504 (N_15504,N_13377,N_13305);
and U15505 (N_15505,N_13644,N_13010);
or U15506 (N_15506,N_12818,N_13141);
xor U15507 (N_15507,N_12003,N_13065);
nor U15508 (N_15508,N_13217,N_12319);
xor U15509 (N_15509,N_13669,N_13177);
or U15510 (N_15510,N_13271,N_13619);
and U15511 (N_15511,N_12560,N_12502);
and U15512 (N_15512,N_13503,N_13691);
and U15513 (N_15513,N_13059,N_13707);
or U15514 (N_15514,N_12478,N_12315);
xor U15515 (N_15515,N_12646,N_13011);
nor U15516 (N_15516,N_13361,N_12125);
and U15517 (N_15517,N_13851,N_12826);
nand U15518 (N_15518,N_12291,N_13594);
nor U15519 (N_15519,N_13559,N_12350);
or U15520 (N_15520,N_12380,N_13536);
or U15521 (N_15521,N_13295,N_12173);
nor U15522 (N_15522,N_13816,N_12007);
and U15523 (N_15523,N_12618,N_12431);
xnor U15524 (N_15524,N_12397,N_12646);
and U15525 (N_15525,N_13010,N_12988);
xnor U15526 (N_15526,N_13396,N_12160);
nand U15527 (N_15527,N_12805,N_13891);
nand U15528 (N_15528,N_12986,N_13495);
xnor U15529 (N_15529,N_13372,N_13248);
nand U15530 (N_15530,N_12737,N_12791);
or U15531 (N_15531,N_13067,N_12187);
nand U15532 (N_15532,N_12957,N_13788);
or U15533 (N_15533,N_13494,N_12589);
nand U15534 (N_15534,N_12255,N_13485);
nand U15535 (N_15535,N_12939,N_13289);
and U15536 (N_15536,N_12386,N_13430);
and U15537 (N_15537,N_12793,N_12548);
xnor U15538 (N_15538,N_12360,N_12063);
nand U15539 (N_15539,N_13385,N_13211);
or U15540 (N_15540,N_13531,N_12834);
nor U15541 (N_15541,N_13482,N_12808);
nand U15542 (N_15542,N_12701,N_13126);
and U15543 (N_15543,N_13249,N_12946);
or U15544 (N_15544,N_12752,N_12413);
nand U15545 (N_15545,N_12387,N_12461);
or U15546 (N_15546,N_13650,N_13739);
xor U15547 (N_15547,N_13972,N_12408);
nor U15548 (N_15548,N_13543,N_12032);
or U15549 (N_15549,N_13610,N_12188);
and U15550 (N_15550,N_13110,N_13606);
nand U15551 (N_15551,N_12541,N_13550);
xnor U15552 (N_15552,N_13993,N_13692);
and U15553 (N_15553,N_13045,N_12639);
and U15554 (N_15554,N_13096,N_12998);
nor U15555 (N_15555,N_13587,N_13952);
or U15556 (N_15556,N_12265,N_13154);
nand U15557 (N_15557,N_12678,N_13825);
nor U15558 (N_15558,N_13768,N_12098);
or U15559 (N_15559,N_12382,N_12757);
xnor U15560 (N_15560,N_13835,N_13129);
nand U15561 (N_15561,N_12474,N_12138);
nand U15562 (N_15562,N_12909,N_12933);
nor U15563 (N_15563,N_13244,N_13725);
nor U15564 (N_15564,N_13004,N_13349);
or U15565 (N_15565,N_13325,N_12959);
or U15566 (N_15566,N_12179,N_13851);
xor U15567 (N_15567,N_13796,N_13810);
xnor U15568 (N_15568,N_13134,N_13245);
nand U15569 (N_15569,N_13539,N_12075);
nor U15570 (N_15570,N_13874,N_13121);
and U15571 (N_15571,N_13403,N_13052);
or U15572 (N_15572,N_12564,N_12465);
or U15573 (N_15573,N_13975,N_13784);
nand U15574 (N_15574,N_12405,N_12444);
and U15575 (N_15575,N_12638,N_13643);
nor U15576 (N_15576,N_13377,N_12024);
or U15577 (N_15577,N_13358,N_13323);
or U15578 (N_15578,N_13668,N_12828);
nor U15579 (N_15579,N_13978,N_13285);
nand U15580 (N_15580,N_12739,N_13714);
xor U15581 (N_15581,N_13067,N_12693);
nor U15582 (N_15582,N_13416,N_12939);
xor U15583 (N_15583,N_13250,N_13615);
nor U15584 (N_15584,N_12035,N_13989);
nand U15585 (N_15585,N_12133,N_12180);
or U15586 (N_15586,N_12576,N_12153);
nand U15587 (N_15587,N_13420,N_12788);
and U15588 (N_15588,N_13882,N_13508);
nand U15589 (N_15589,N_12171,N_13152);
or U15590 (N_15590,N_13287,N_12269);
nand U15591 (N_15591,N_12709,N_13383);
nor U15592 (N_15592,N_12957,N_12470);
nor U15593 (N_15593,N_13208,N_12209);
xnor U15594 (N_15594,N_12650,N_12826);
xnor U15595 (N_15595,N_13054,N_13076);
and U15596 (N_15596,N_12128,N_13063);
and U15597 (N_15597,N_13821,N_13709);
nand U15598 (N_15598,N_12676,N_12476);
and U15599 (N_15599,N_13554,N_12761);
xor U15600 (N_15600,N_12932,N_12953);
nand U15601 (N_15601,N_12009,N_13688);
nand U15602 (N_15602,N_13132,N_13761);
or U15603 (N_15603,N_12296,N_12056);
or U15604 (N_15604,N_13556,N_13164);
xnor U15605 (N_15605,N_12695,N_12812);
and U15606 (N_15606,N_12153,N_12132);
and U15607 (N_15607,N_12965,N_13215);
and U15608 (N_15608,N_12920,N_13582);
nor U15609 (N_15609,N_12592,N_13664);
or U15610 (N_15610,N_12201,N_12164);
nor U15611 (N_15611,N_12013,N_12059);
nand U15612 (N_15612,N_12818,N_12755);
or U15613 (N_15613,N_12410,N_13022);
nand U15614 (N_15614,N_12324,N_12533);
or U15615 (N_15615,N_13312,N_13861);
xnor U15616 (N_15616,N_13213,N_13969);
and U15617 (N_15617,N_12265,N_13813);
or U15618 (N_15618,N_13043,N_13993);
nor U15619 (N_15619,N_12335,N_13541);
nand U15620 (N_15620,N_13237,N_13256);
nor U15621 (N_15621,N_13996,N_12236);
or U15622 (N_15622,N_13189,N_12641);
nor U15623 (N_15623,N_12346,N_12128);
and U15624 (N_15624,N_13867,N_12890);
nor U15625 (N_15625,N_13349,N_13913);
nand U15626 (N_15626,N_12356,N_13705);
nor U15627 (N_15627,N_13682,N_13815);
xnor U15628 (N_15628,N_13470,N_13406);
nand U15629 (N_15629,N_12692,N_13376);
nand U15630 (N_15630,N_13506,N_13965);
and U15631 (N_15631,N_13507,N_12079);
or U15632 (N_15632,N_12804,N_13444);
nand U15633 (N_15633,N_12731,N_13962);
nand U15634 (N_15634,N_13243,N_12471);
nor U15635 (N_15635,N_13606,N_12039);
or U15636 (N_15636,N_13027,N_12746);
nand U15637 (N_15637,N_12749,N_13550);
xnor U15638 (N_15638,N_12961,N_12847);
nand U15639 (N_15639,N_12169,N_12171);
nand U15640 (N_15640,N_13277,N_12989);
and U15641 (N_15641,N_13830,N_13421);
or U15642 (N_15642,N_12837,N_13506);
or U15643 (N_15643,N_13744,N_12564);
and U15644 (N_15644,N_12159,N_13224);
nor U15645 (N_15645,N_12840,N_12932);
nor U15646 (N_15646,N_13309,N_13112);
nor U15647 (N_15647,N_12717,N_12459);
nand U15648 (N_15648,N_12839,N_13956);
or U15649 (N_15649,N_12568,N_12494);
nor U15650 (N_15650,N_13182,N_12941);
and U15651 (N_15651,N_13849,N_12056);
nand U15652 (N_15652,N_12921,N_13133);
nor U15653 (N_15653,N_13739,N_13168);
nor U15654 (N_15654,N_13907,N_13072);
xnor U15655 (N_15655,N_13277,N_13370);
nand U15656 (N_15656,N_13678,N_12204);
and U15657 (N_15657,N_13391,N_13244);
nand U15658 (N_15658,N_13530,N_13441);
or U15659 (N_15659,N_12813,N_13414);
and U15660 (N_15660,N_12969,N_12286);
nor U15661 (N_15661,N_12409,N_12338);
nand U15662 (N_15662,N_12228,N_12140);
nor U15663 (N_15663,N_13195,N_12285);
or U15664 (N_15664,N_13742,N_13032);
nor U15665 (N_15665,N_12182,N_13503);
and U15666 (N_15666,N_13084,N_13059);
nand U15667 (N_15667,N_13379,N_12034);
xnor U15668 (N_15668,N_13524,N_12945);
nand U15669 (N_15669,N_12513,N_13631);
nor U15670 (N_15670,N_12524,N_13760);
xor U15671 (N_15671,N_13270,N_13002);
and U15672 (N_15672,N_13965,N_13699);
or U15673 (N_15673,N_13866,N_13823);
nor U15674 (N_15674,N_13732,N_13904);
and U15675 (N_15675,N_13077,N_12427);
and U15676 (N_15676,N_13100,N_13879);
nand U15677 (N_15677,N_13874,N_12166);
or U15678 (N_15678,N_12620,N_13114);
or U15679 (N_15679,N_13863,N_13206);
or U15680 (N_15680,N_12162,N_13317);
or U15681 (N_15681,N_12425,N_12590);
xor U15682 (N_15682,N_12988,N_12595);
nor U15683 (N_15683,N_13891,N_12763);
and U15684 (N_15684,N_12904,N_12733);
nand U15685 (N_15685,N_13854,N_13141);
xnor U15686 (N_15686,N_12345,N_13203);
or U15687 (N_15687,N_12698,N_12321);
and U15688 (N_15688,N_13929,N_12267);
or U15689 (N_15689,N_12253,N_13022);
nor U15690 (N_15690,N_13632,N_13741);
xnor U15691 (N_15691,N_13776,N_12936);
nand U15692 (N_15692,N_12653,N_12165);
nor U15693 (N_15693,N_13395,N_12861);
and U15694 (N_15694,N_12371,N_12432);
nand U15695 (N_15695,N_13014,N_12769);
nand U15696 (N_15696,N_12826,N_13037);
xor U15697 (N_15697,N_13076,N_12408);
and U15698 (N_15698,N_12268,N_12723);
nand U15699 (N_15699,N_12029,N_13584);
xnor U15700 (N_15700,N_13783,N_13604);
nand U15701 (N_15701,N_13402,N_13717);
xnor U15702 (N_15702,N_13922,N_12650);
nor U15703 (N_15703,N_13807,N_13280);
nand U15704 (N_15704,N_12307,N_13868);
nor U15705 (N_15705,N_13787,N_13068);
nor U15706 (N_15706,N_12557,N_12037);
nand U15707 (N_15707,N_13065,N_13887);
xor U15708 (N_15708,N_13715,N_13677);
nand U15709 (N_15709,N_12049,N_12874);
nand U15710 (N_15710,N_12304,N_12522);
and U15711 (N_15711,N_12543,N_12167);
or U15712 (N_15712,N_13192,N_13008);
or U15713 (N_15713,N_13223,N_13930);
nand U15714 (N_15714,N_12036,N_12042);
nor U15715 (N_15715,N_13949,N_13866);
xnor U15716 (N_15716,N_13626,N_12981);
or U15717 (N_15717,N_13096,N_13462);
xnor U15718 (N_15718,N_13575,N_13884);
and U15719 (N_15719,N_12903,N_12914);
nand U15720 (N_15720,N_13935,N_12672);
nand U15721 (N_15721,N_13473,N_12317);
or U15722 (N_15722,N_13441,N_13820);
xor U15723 (N_15723,N_12265,N_12046);
nor U15724 (N_15724,N_12787,N_13677);
nand U15725 (N_15725,N_13857,N_13068);
nor U15726 (N_15726,N_13545,N_12189);
xor U15727 (N_15727,N_13299,N_12928);
and U15728 (N_15728,N_13620,N_13128);
nor U15729 (N_15729,N_12574,N_12494);
nand U15730 (N_15730,N_13590,N_12306);
xor U15731 (N_15731,N_12188,N_12132);
nand U15732 (N_15732,N_12527,N_13492);
or U15733 (N_15733,N_12843,N_13402);
xnor U15734 (N_15734,N_12955,N_12152);
nand U15735 (N_15735,N_13792,N_13345);
nand U15736 (N_15736,N_12650,N_13082);
nand U15737 (N_15737,N_12286,N_12545);
xnor U15738 (N_15738,N_12178,N_12972);
nor U15739 (N_15739,N_12377,N_12481);
nor U15740 (N_15740,N_12684,N_12250);
nor U15741 (N_15741,N_13239,N_12062);
xnor U15742 (N_15742,N_13533,N_12435);
nor U15743 (N_15743,N_13245,N_13168);
nor U15744 (N_15744,N_12243,N_13011);
or U15745 (N_15745,N_12293,N_12612);
and U15746 (N_15746,N_12139,N_13674);
or U15747 (N_15747,N_12322,N_13588);
xnor U15748 (N_15748,N_13444,N_12665);
nor U15749 (N_15749,N_13829,N_12737);
nor U15750 (N_15750,N_13807,N_13222);
and U15751 (N_15751,N_13509,N_12331);
and U15752 (N_15752,N_12237,N_12065);
nor U15753 (N_15753,N_13585,N_12087);
xnor U15754 (N_15754,N_12132,N_12669);
nor U15755 (N_15755,N_12977,N_12302);
xnor U15756 (N_15756,N_13273,N_12870);
nand U15757 (N_15757,N_12555,N_12519);
or U15758 (N_15758,N_12996,N_12052);
nand U15759 (N_15759,N_12714,N_13415);
nand U15760 (N_15760,N_13332,N_13042);
or U15761 (N_15761,N_13625,N_12756);
nor U15762 (N_15762,N_13322,N_13416);
nor U15763 (N_15763,N_13814,N_12290);
nor U15764 (N_15764,N_13866,N_13531);
and U15765 (N_15765,N_12802,N_13927);
or U15766 (N_15766,N_13199,N_13589);
nand U15767 (N_15767,N_12590,N_13660);
and U15768 (N_15768,N_13328,N_12695);
and U15769 (N_15769,N_13244,N_12867);
or U15770 (N_15770,N_12767,N_13885);
nor U15771 (N_15771,N_12130,N_13647);
or U15772 (N_15772,N_12696,N_12562);
nor U15773 (N_15773,N_12194,N_12235);
xor U15774 (N_15774,N_13193,N_13523);
xnor U15775 (N_15775,N_13130,N_13772);
nor U15776 (N_15776,N_13438,N_13195);
xor U15777 (N_15777,N_12212,N_12443);
nor U15778 (N_15778,N_12711,N_13719);
or U15779 (N_15779,N_12306,N_13918);
nor U15780 (N_15780,N_13401,N_13310);
xor U15781 (N_15781,N_12013,N_12915);
and U15782 (N_15782,N_12466,N_13659);
and U15783 (N_15783,N_13841,N_13705);
nand U15784 (N_15784,N_13689,N_12986);
nand U15785 (N_15785,N_12563,N_13987);
xnor U15786 (N_15786,N_12730,N_12216);
or U15787 (N_15787,N_12714,N_12657);
and U15788 (N_15788,N_12125,N_12531);
or U15789 (N_15789,N_13441,N_12548);
nor U15790 (N_15790,N_12855,N_12021);
and U15791 (N_15791,N_12158,N_12312);
nor U15792 (N_15792,N_12127,N_13968);
nor U15793 (N_15793,N_12708,N_12798);
nor U15794 (N_15794,N_13007,N_12185);
nor U15795 (N_15795,N_12093,N_13504);
and U15796 (N_15796,N_13772,N_13867);
nor U15797 (N_15797,N_12538,N_13797);
xnor U15798 (N_15798,N_13327,N_13993);
or U15799 (N_15799,N_12456,N_12316);
nand U15800 (N_15800,N_13763,N_13401);
and U15801 (N_15801,N_13495,N_12707);
and U15802 (N_15802,N_13980,N_12908);
xnor U15803 (N_15803,N_12227,N_12722);
nand U15804 (N_15804,N_12865,N_12875);
or U15805 (N_15805,N_13777,N_13398);
nor U15806 (N_15806,N_13015,N_12796);
nor U15807 (N_15807,N_13649,N_12950);
xnor U15808 (N_15808,N_13638,N_13331);
xnor U15809 (N_15809,N_13496,N_13398);
xnor U15810 (N_15810,N_13883,N_12138);
xor U15811 (N_15811,N_12354,N_12558);
nand U15812 (N_15812,N_13817,N_12618);
and U15813 (N_15813,N_12746,N_12441);
and U15814 (N_15814,N_12536,N_13999);
and U15815 (N_15815,N_13043,N_12567);
nand U15816 (N_15816,N_12925,N_12257);
and U15817 (N_15817,N_13827,N_13015);
nand U15818 (N_15818,N_13073,N_12877);
and U15819 (N_15819,N_13196,N_13750);
xnor U15820 (N_15820,N_12012,N_13762);
or U15821 (N_15821,N_13252,N_12239);
xnor U15822 (N_15822,N_12626,N_13161);
or U15823 (N_15823,N_12534,N_12512);
xnor U15824 (N_15824,N_13969,N_13050);
nand U15825 (N_15825,N_13741,N_13943);
nand U15826 (N_15826,N_13624,N_12476);
or U15827 (N_15827,N_12506,N_12708);
nor U15828 (N_15828,N_13948,N_13897);
nand U15829 (N_15829,N_12829,N_12353);
xor U15830 (N_15830,N_13691,N_12851);
or U15831 (N_15831,N_13862,N_13429);
nand U15832 (N_15832,N_13784,N_12776);
and U15833 (N_15833,N_13968,N_13162);
nor U15834 (N_15834,N_13533,N_12858);
xnor U15835 (N_15835,N_12949,N_12316);
nand U15836 (N_15836,N_13198,N_12708);
and U15837 (N_15837,N_12284,N_12435);
nor U15838 (N_15838,N_12165,N_12094);
xor U15839 (N_15839,N_12355,N_12242);
nand U15840 (N_15840,N_12723,N_13133);
nor U15841 (N_15841,N_12754,N_13638);
nand U15842 (N_15842,N_13803,N_12132);
and U15843 (N_15843,N_12629,N_12468);
nand U15844 (N_15844,N_12788,N_13067);
nor U15845 (N_15845,N_13554,N_13291);
nor U15846 (N_15846,N_13377,N_12570);
xnor U15847 (N_15847,N_13007,N_12031);
nand U15848 (N_15848,N_12128,N_12070);
xor U15849 (N_15849,N_12102,N_12328);
nor U15850 (N_15850,N_13199,N_13677);
xor U15851 (N_15851,N_13432,N_13920);
or U15852 (N_15852,N_12113,N_13285);
or U15853 (N_15853,N_12265,N_12369);
xor U15854 (N_15854,N_13500,N_12519);
xor U15855 (N_15855,N_13872,N_12419);
nor U15856 (N_15856,N_13064,N_12519);
and U15857 (N_15857,N_12945,N_13398);
nor U15858 (N_15858,N_12079,N_13446);
nor U15859 (N_15859,N_13884,N_12214);
nor U15860 (N_15860,N_12105,N_13730);
nor U15861 (N_15861,N_12669,N_12154);
nand U15862 (N_15862,N_13772,N_12110);
and U15863 (N_15863,N_12597,N_13697);
xor U15864 (N_15864,N_13677,N_13324);
nand U15865 (N_15865,N_12983,N_12698);
and U15866 (N_15866,N_12330,N_12233);
nand U15867 (N_15867,N_12950,N_13121);
and U15868 (N_15868,N_13908,N_13407);
xnor U15869 (N_15869,N_13562,N_13988);
nor U15870 (N_15870,N_13776,N_13743);
or U15871 (N_15871,N_13206,N_13655);
or U15872 (N_15872,N_12625,N_13604);
nand U15873 (N_15873,N_12469,N_12965);
nor U15874 (N_15874,N_12968,N_12077);
nor U15875 (N_15875,N_12728,N_12057);
or U15876 (N_15876,N_12024,N_12738);
nand U15877 (N_15877,N_13079,N_13225);
and U15878 (N_15878,N_13052,N_13767);
xnor U15879 (N_15879,N_12735,N_12526);
or U15880 (N_15880,N_12119,N_13615);
and U15881 (N_15881,N_12022,N_12179);
nor U15882 (N_15882,N_13556,N_12518);
nand U15883 (N_15883,N_13103,N_12498);
nand U15884 (N_15884,N_12587,N_13350);
xor U15885 (N_15885,N_13042,N_12627);
nor U15886 (N_15886,N_12590,N_12602);
and U15887 (N_15887,N_13364,N_12539);
nand U15888 (N_15888,N_13415,N_13474);
nor U15889 (N_15889,N_12186,N_13577);
or U15890 (N_15890,N_12911,N_13542);
and U15891 (N_15891,N_12666,N_12681);
nand U15892 (N_15892,N_12783,N_12435);
and U15893 (N_15893,N_13504,N_12815);
nand U15894 (N_15894,N_12401,N_12057);
and U15895 (N_15895,N_13931,N_12486);
nand U15896 (N_15896,N_13583,N_12825);
nand U15897 (N_15897,N_12552,N_13397);
xor U15898 (N_15898,N_12643,N_12779);
and U15899 (N_15899,N_12680,N_12693);
xor U15900 (N_15900,N_12351,N_12799);
and U15901 (N_15901,N_12822,N_13173);
nand U15902 (N_15902,N_13731,N_13819);
or U15903 (N_15903,N_13397,N_12456);
nand U15904 (N_15904,N_12608,N_13513);
xnor U15905 (N_15905,N_12853,N_12056);
xnor U15906 (N_15906,N_12711,N_13008);
or U15907 (N_15907,N_13296,N_13740);
and U15908 (N_15908,N_12474,N_12021);
nand U15909 (N_15909,N_13996,N_13310);
nand U15910 (N_15910,N_13472,N_13349);
and U15911 (N_15911,N_13959,N_12616);
nor U15912 (N_15912,N_13208,N_12843);
or U15913 (N_15913,N_13536,N_12842);
nor U15914 (N_15914,N_12045,N_12504);
nand U15915 (N_15915,N_12307,N_13692);
and U15916 (N_15916,N_13666,N_12548);
xor U15917 (N_15917,N_13845,N_12245);
xnor U15918 (N_15918,N_12420,N_13685);
or U15919 (N_15919,N_13514,N_12522);
nor U15920 (N_15920,N_12283,N_12742);
or U15921 (N_15921,N_13303,N_13000);
nor U15922 (N_15922,N_13774,N_12240);
xor U15923 (N_15923,N_12110,N_12198);
nand U15924 (N_15924,N_13088,N_12897);
and U15925 (N_15925,N_13367,N_13753);
nand U15926 (N_15926,N_12706,N_12595);
nor U15927 (N_15927,N_12184,N_12498);
nor U15928 (N_15928,N_12049,N_13264);
xnor U15929 (N_15929,N_12274,N_12424);
nor U15930 (N_15930,N_13948,N_12350);
nand U15931 (N_15931,N_12221,N_12888);
nor U15932 (N_15932,N_13374,N_12592);
and U15933 (N_15933,N_13794,N_13545);
nand U15934 (N_15934,N_12158,N_13167);
and U15935 (N_15935,N_13835,N_13055);
xor U15936 (N_15936,N_13842,N_12922);
and U15937 (N_15937,N_13468,N_13395);
xor U15938 (N_15938,N_12407,N_12442);
xor U15939 (N_15939,N_13230,N_12707);
nor U15940 (N_15940,N_12015,N_13604);
nand U15941 (N_15941,N_12920,N_12148);
and U15942 (N_15942,N_12663,N_13760);
nand U15943 (N_15943,N_13376,N_12050);
or U15944 (N_15944,N_13368,N_13103);
nor U15945 (N_15945,N_12740,N_13773);
or U15946 (N_15946,N_13065,N_12014);
nand U15947 (N_15947,N_13812,N_12140);
nand U15948 (N_15948,N_13429,N_12369);
nor U15949 (N_15949,N_12153,N_12992);
xnor U15950 (N_15950,N_12220,N_12398);
xnor U15951 (N_15951,N_13010,N_13008);
or U15952 (N_15952,N_13865,N_12346);
nor U15953 (N_15953,N_13581,N_12727);
xor U15954 (N_15954,N_12171,N_12298);
nand U15955 (N_15955,N_12714,N_13027);
or U15956 (N_15956,N_13573,N_12515);
nor U15957 (N_15957,N_13116,N_13381);
nor U15958 (N_15958,N_12121,N_13769);
nor U15959 (N_15959,N_13242,N_12420);
and U15960 (N_15960,N_13141,N_13859);
or U15961 (N_15961,N_13117,N_13111);
nand U15962 (N_15962,N_13896,N_13431);
nand U15963 (N_15963,N_12637,N_12599);
or U15964 (N_15964,N_13285,N_13980);
or U15965 (N_15965,N_12375,N_13905);
or U15966 (N_15966,N_12220,N_12333);
xnor U15967 (N_15967,N_13604,N_12120);
and U15968 (N_15968,N_12248,N_12486);
nand U15969 (N_15969,N_13227,N_13331);
nand U15970 (N_15970,N_12637,N_12018);
nand U15971 (N_15971,N_13812,N_12482);
and U15972 (N_15972,N_13840,N_13203);
or U15973 (N_15973,N_13066,N_12318);
nor U15974 (N_15974,N_13282,N_13448);
nand U15975 (N_15975,N_13248,N_12458);
nand U15976 (N_15976,N_13557,N_12714);
xnor U15977 (N_15977,N_13002,N_12131);
and U15978 (N_15978,N_12816,N_12900);
nor U15979 (N_15979,N_13052,N_12556);
nand U15980 (N_15980,N_12101,N_13220);
xor U15981 (N_15981,N_13276,N_13236);
xor U15982 (N_15982,N_12116,N_13780);
or U15983 (N_15983,N_13776,N_13186);
xor U15984 (N_15984,N_13179,N_13047);
nor U15985 (N_15985,N_12770,N_13540);
and U15986 (N_15986,N_12775,N_13368);
nor U15987 (N_15987,N_12433,N_12883);
and U15988 (N_15988,N_13147,N_12659);
xnor U15989 (N_15989,N_12021,N_13495);
nand U15990 (N_15990,N_12591,N_12365);
xor U15991 (N_15991,N_13995,N_13186);
or U15992 (N_15992,N_12911,N_13154);
nand U15993 (N_15993,N_12868,N_12588);
xnor U15994 (N_15994,N_13129,N_13701);
and U15995 (N_15995,N_13904,N_12325);
and U15996 (N_15996,N_13544,N_12957);
or U15997 (N_15997,N_12333,N_12211);
or U15998 (N_15998,N_12658,N_12467);
or U15999 (N_15999,N_13998,N_12708);
xor U16000 (N_16000,N_14725,N_15394);
nor U16001 (N_16001,N_14329,N_14043);
nand U16002 (N_16002,N_14560,N_14228);
nand U16003 (N_16003,N_15588,N_15555);
nor U16004 (N_16004,N_14480,N_15808);
nor U16005 (N_16005,N_15744,N_15146);
xnor U16006 (N_16006,N_15391,N_14941);
nand U16007 (N_16007,N_14619,N_15540);
and U16008 (N_16008,N_15234,N_14240);
nor U16009 (N_16009,N_15210,N_14924);
and U16010 (N_16010,N_15503,N_15524);
or U16011 (N_16011,N_14889,N_15439);
or U16012 (N_16012,N_15088,N_14973);
or U16013 (N_16013,N_14007,N_14584);
or U16014 (N_16014,N_14113,N_15519);
and U16015 (N_16015,N_14188,N_14731);
nand U16016 (N_16016,N_15792,N_14376);
nor U16017 (N_16017,N_15732,N_15125);
and U16018 (N_16018,N_15919,N_15991);
nand U16019 (N_16019,N_14651,N_15355);
nor U16020 (N_16020,N_14611,N_15186);
nand U16021 (N_16021,N_14243,N_15859);
or U16022 (N_16022,N_15675,N_15518);
xor U16023 (N_16023,N_15830,N_15111);
and U16024 (N_16024,N_15143,N_14710);
or U16025 (N_16025,N_14729,N_15052);
or U16026 (N_16026,N_15305,N_15538);
xor U16027 (N_16027,N_14919,N_14750);
or U16028 (N_16028,N_14896,N_14749);
nor U16029 (N_16029,N_14022,N_15688);
xnor U16030 (N_16030,N_15451,N_14878);
nor U16031 (N_16031,N_15119,N_15846);
or U16032 (N_16032,N_14829,N_15331);
xor U16033 (N_16033,N_15168,N_15662);
nor U16034 (N_16034,N_14492,N_14106);
nand U16035 (N_16035,N_14988,N_14014);
or U16036 (N_16036,N_14332,N_15083);
xor U16037 (N_16037,N_15115,N_14039);
or U16038 (N_16038,N_14002,N_14618);
nand U16039 (N_16039,N_15800,N_14672);
xor U16040 (N_16040,N_14516,N_15110);
and U16041 (N_16041,N_15340,N_14679);
and U16042 (N_16042,N_15856,N_15383);
and U16043 (N_16043,N_14925,N_15736);
and U16044 (N_16044,N_14174,N_15342);
and U16045 (N_16045,N_14377,N_14649);
xor U16046 (N_16046,N_14169,N_15109);
or U16047 (N_16047,N_14694,N_15063);
and U16048 (N_16048,N_14975,N_14459);
nor U16049 (N_16049,N_15563,N_15657);
nand U16050 (N_16050,N_15378,N_15287);
nand U16051 (N_16051,N_14762,N_15698);
xnor U16052 (N_16052,N_14860,N_15703);
nand U16053 (N_16053,N_15395,N_15087);
xnor U16054 (N_16054,N_15733,N_15105);
or U16055 (N_16055,N_15084,N_14264);
nor U16056 (N_16056,N_14470,N_15386);
or U16057 (N_16057,N_15623,N_15481);
nor U16058 (N_16058,N_15738,N_15285);
or U16059 (N_16059,N_15334,N_15018);
xor U16060 (N_16060,N_14094,N_15248);
or U16061 (N_16061,N_15631,N_15136);
nor U16062 (N_16062,N_14872,N_14382);
xnor U16063 (N_16063,N_15909,N_15674);
nor U16064 (N_16064,N_15174,N_14756);
nand U16065 (N_16065,N_15825,N_14708);
and U16066 (N_16066,N_14876,N_15075);
nor U16067 (N_16067,N_15527,N_15372);
nor U16068 (N_16068,N_14780,N_15145);
nand U16069 (N_16069,N_14139,N_15769);
nand U16070 (N_16070,N_15155,N_14657);
or U16071 (N_16071,N_14206,N_14531);
or U16072 (N_16072,N_15892,N_14341);
or U16073 (N_16073,N_14912,N_14783);
nor U16074 (N_16074,N_14099,N_15150);
nor U16075 (N_16075,N_15534,N_15323);
and U16076 (N_16076,N_15508,N_15878);
xor U16077 (N_16077,N_15941,N_14349);
or U16078 (N_16078,N_14478,N_14449);
xor U16079 (N_16079,N_15795,N_15224);
nor U16080 (N_16080,N_14504,N_15643);
and U16081 (N_16081,N_14309,N_14236);
or U16082 (N_16082,N_15123,N_14251);
xnor U16083 (N_16083,N_14929,N_15341);
nand U16084 (N_16084,N_15200,N_15290);
nand U16085 (N_16085,N_15138,N_14882);
nor U16086 (N_16086,N_14322,N_14127);
xnor U16087 (N_16087,N_14056,N_15868);
or U16088 (N_16088,N_14899,N_14763);
nand U16089 (N_16089,N_14086,N_14301);
xnor U16090 (N_16090,N_14442,N_14947);
nand U16091 (N_16091,N_15324,N_15203);
xor U16092 (N_16092,N_15057,N_14408);
or U16093 (N_16093,N_14418,N_15494);
and U16094 (N_16094,N_15515,N_15983);
nand U16095 (N_16095,N_14663,N_15361);
nand U16096 (N_16096,N_15724,N_15132);
xnor U16097 (N_16097,N_15484,N_15205);
xor U16098 (N_16098,N_14686,N_14913);
nand U16099 (N_16099,N_15928,N_15887);
nand U16100 (N_16100,N_15992,N_14304);
nor U16101 (N_16101,N_14898,N_15262);
nand U16102 (N_16102,N_14930,N_15626);
xor U16103 (N_16103,N_14253,N_14211);
or U16104 (N_16104,N_15961,N_15398);
nor U16105 (N_16105,N_15625,N_15103);
nand U16106 (N_16106,N_15986,N_15901);
xnor U16107 (N_16107,N_14968,N_15010);
nand U16108 (N_16108,N_15475,N_15836);
nor U16109 (N_16109,N_14137,N_15875);
or U16110 (N_16110,N_15078,N_14074);
and U16111 (N_16111,N_15801,N_14786);
and U16112 (N_16112,N_15865,N_15573);
nand U16113 (N_16113,N_14939,N_14358);
nand U16114 (N_16114,N_15905,N_15434);
nor U16115 (N_16115,N_15419,N_15029);
or U16116 (N_16116,N_15762,N_14916);
nand U16117 (N_16117,N_14688,N_14055);
nor U16118 (N_16118,N_14932,N_14668);
or U16119 (N_16119,N_14928,N_15824);
and U16120 (N_16120,N_14095,N_14892);
and U16121 (N_16121,N_15635,N_14967);
nor U16122 (N_16122,N_14573,N_14460);
nor U16123 (N_16123,N_14483,N_14202);
nand U16124 (N_16124,N_15943,N_15760);
nor U16125 (N_16125,N_14414,N_14096);
and U16126 (N_16126,N_14515,N_15788);
or U16127 (N_16127,N_15741,N_15908);
xnor U16128 (N_16128,N_15665,N_15554);
or U16129 (N_16129,N_15007,N_14751);
nand U16130 (N_16130,N_15432,N_15407);
or U16131 (N_16131,N_15458,N_14764);
and U16132 (N_16132,N_14294,N_14360);
and U16133 (N_16133,N_14656,N_15498);
xnor U16134 (N_16134,N_14394,N_15188);
nand U16135 (N_16135,N_15086,N_15929);
or U16136 (N_16136,N_14286,N_14436);
and U16137 (N_16137,N_14716,N_15178);
or U16138 (N_16138,N_14557,N_15707);
or U16139 (N_16139,N_15809,N_14718);
or U16140 (N_16140,N_15373,N_14072);
and U16141 (N_16141,N_15768,N_15402);
nor U16142 (N_16142,N_14844,N_15972);
nand U16143 (N_16143,N_15076,N_15443);
and U16144 (N_16144,N_15399,N_14960);
or U16145 (N_16145,N_15776,N_15172);
xor U16146 (N_16146,N_14849,N_14000);
or U16147 (N_16147,N_14157,N_15604);
or U16148 (N_16148,N_15023,N_15032);
nand U16149 (N_16149,N_14571,N_15851);
and U16150 (N_16150,N_15026,N_15356);
nor U16151 (N_16151,N_14662,N_14295);
xor U16152 (N_16152,N_14276,N_15506);
nor U16153 (N_16153,N_14509,N_15797);
xnor U16154 (N_16154,N_15617,N_15006);
nor U16155 (N_16155,N_14902,N_14108);
or U16156 (N_16156,N_15435,N_14468);
nor U16157 (N_16157,N_15676,N_14175);
or U16158 (N_16158,N_14877,N_15814);
nand U16159 (N_16159,N_15339,N_14392);
nand U16160 (N_16160,N_15579,N_15216);
xnor U16161 (N_16161,N_14566,N_15229);
and U16162 (N_16162,N_14365,N_14350);
nor U16163 (N_16163,N_14858,N_14904);
or U16164 (N_16164,N_15144,N_15864);
and U16165 (N_16165,N_14397,N_15169);
nand U16166 (N_16166,N_15751,N_14146);
xor U16167 (N_16167,N_14634,N_15935);
xor U16168 (N_16168,N_15615,N_14541);
nor U16169 (N_16169,N_15608,N_14704);
and U16170 (N_16170,N_15377,N_15357);
or U16171 (N_16171,N_15039,N_15156);
xor U16172 (N_16172,N_15263,N_14693);
nor U16173 (N_16173,N_14777,N_14069);
or U16174 (N_16174,N_15124,N_14230);
xnor U16175 (N_16175,N_14768,N_14315);
or U16176 (N_16176,N_15525,N_15912);
and U16177 (N_16177,N_14031,N_14035);
and U16178 (N_16178,N_15596,N_14125);
or U16179 (N_16179,N_15055,N_15737);
or U16180 (N_16180,N_14773,N_14111);
nor U16181 (N_16181,N_14555,N_15096);
xor U16182 (N_16182,N_15592,N_14626);
and U16183 (N_16183,N_15478,N_14303);
or U16184 (N_16184,N_14907,N_14241);
or U16185 (N_16185,N_15690,N_15723);
nor U16186 (N_16186,N_15022,N_14739);
nor U16187 (N_16187,N_15107,N_15148);
and U16188 (N_16188,N_14989,N_14451);
or U16189 (N_16189,N_14330,N_14724);
nand U16190 (N_16190,N_15822,N_15677);
nand U16191 (N_16191,N_15058,N_14730);
xnor U16192 (N_16192,N_15456,N_14698);
xnor U16193 (N_16193,N_14354,N_15922);
or U16194 (N_16194,N_15500,N_15896);
or U16195 (N_16195,N_15713,N_14864);
nor U16196 (N_16196,N_14592,N_14713);
nor U16197 (N_16197,N_14009,N_14869);
nor U16198 (N_16198,N_14894,N_14300);
and U16199 (N_16199,N_15535,N_15763);
and U16200 (N_16200,N_14816,N_14542);
nand U16201 (N_16201,N_15872,N_14275);
and U16202 (N_16202,N_14806,N_14824);
or U16203 (N_16203,N_14413,N_14888);
and U16204 (N_16204,N_15359,N_15265);
xnor U16205 (N_16205,N_14424,N_14937);
xor U16206 (N_16206,N_15687,N_14732);
or U16207 (N_16207,N_14855,N_14999);
nor U16208 (N_16208,N_15080,N_14165);
or U16209 (N_16209,N_14905,N_15658);
or U16210 (N_16210,N_15311,N_14701);
and U16211 (N_16211,N_14525,N_14487);
xor U16212 (N_16212,N_14520,N_14800);
and U16213 (N_16213,N_15684,N_15951);
xnor U16214 (N_16214,N_14795,N_15636);
or U16215 (N_16215,N_15979,N_15988);
or U16216 (N_16216,N_14945,N_14471);
nor U16217 (N_16217,N_15947,N_14970);
nor U16218 (N_16218,N_14637,N_14116);
xnor U16219 (N_16219,N_15139,N_14472);
xor U16220 (N_16220,N_14852,N_14802);
xnor U16221 (N_16221,N_14742,N_14847);
or U16222 (N_16222,N_15195,N_15523);
xor U16223 (N_16223,N_15517,N_14521);
or U16224 (N_16224,N_14700,N_14370);
or U16225 (N_16225,N_14420,N_15335);
xnor U16226 (N_16226,N_14643,N_14384);
xor U16227 (N_16227,N_14790,N_14308);
and U16228 (N_16228,N_14311,N_14998);
xor U16229 (N_16229,N_14798,N_14580);
and U16230 (N_16230,N_15421,N_15620);
and U16231 (N_16231,N_15696,N_14058);
nor U16232 (N_16232,N_14636,N_15302);
or U16233 (N_16233,N_14317,N_14235);
nand U16234 (N_16234,N_14543,N_14918);
nand U16235 (N_16235,N_15807,N_14959);
nand U16236 (N_16236,N_15918,N_15247);
nand U16237 (N_16237,N_15996,N_15940);
xnor U16238 (N_16238,N_14517,N_14687);
nor U16239 (N_16239,N_14302,N_14117);
nor U16240 (N_16240,N_14473,N_14121);
and U16241 (N_16241,N_15306,N_15097);
xor U16242 (N_16242,N_14513,N_14278);
nand U16243 (N_16243,N_14208,N_15253);
nor U16244 (N_16244,N_15975,N_14463);
nand U16245 (N_16245,N_15845,N_15780);
xnor U16246 (N_16246,N_15606,N_15766);
nand U16247 (N_16247,N_14164,N_14952);
and U16248 (N_16248,N_15993,N_14401);
nand U16249 (N_16249,N_14920,N_14461);
xnor U16250 (N_16250,N_14604,N_15582);
nor U16251 (N_16251,N_14362,N_14273);
nand U16252 (N_16252,N_15921,N_14128);
nand U16253 (N_16253,N_14771,N_14444);
and U16254 (N_16254,N_15101,N_15962);
nor U16255 (N_16255,N_15298,N_15051);
xor U16256 (N_16256,N_15584,N_14671);
xor U16257 (N_16257,N_14135,N_14267);
and U16258 (N_16258,N_14505,N_15938);
nor U16259 (N_16259,N_15388,N_14083);
xnor U16260 (N_16260,N_14428,N_14971);
or U16261 (N_16261,N_14992,N_14781);
and U16262 (N_16262,N_14310,N_15379);
nor U16263 (N_16263,N_14715,N_14091);
or U16264 (N_16264,N_14827,N_14066);
or U16265 (N_16265,N_14143,N_14222);
or U16266 (N_16266,N_14775,N_15771);
xnor U16267 (N_16267,N_15542,N_14029);
or U16268 (N_16268,N_15318,N_14486);
and U16269 (N_16269,N_15448,N_15678);
nor U16270 (N_16270,N_15572,N_15995);
xnor U16271 (N_16271,N_14032,N_15672);
xnor U16272 (N_16272,N_14062,N_15702);
nand U16273 (N_16273,N_14050,N_14421);
or U16274 (N_16274,N_15597,N_14110);
and U16275 (N_16275,N_15550,N_14484);
nand U16276 (N_16276,N_14176,N_15589);
nand U16277 (N_16277,N_15042,N_15296);
nor U16278 (N_16278,N_14425,N_14283);
nand U16279 (N_16279,N_14813,N_14102);
and U16280 (N_16280,N_14187,N_15842);
and U16281 (N_16281,N_14677,N_14950);
and U16282 (N_16282,N_14448,N_14796);
nor U16283 (N_16283,N_14522,N_15833);
and U16284 (N_16284,N_14644,N_15189);
nand U16285 (N_16285,N_14978,N_15765);
nand U16286 (N_16286,N_15867,N_15396);
xnor U16287 (N_16287,N_15154,N_15219);
and U16288 (N_16288,N_14841,N_15313);
nand U16289 (N_16289,N_15805,N_15066);
nand U16290 (N_16290,N_14389,N_14528);
nand U16291 (N_16291,N_14572,N_14467);
or U16292 (N_16292,N_15497,N_14450);
and U16293 (N_16293,N_15072,N_15014);
xor U16294 (N_16294,N_15045,N_15436);
xor U16295 (N_16295,N_15561,N_15954);
nor U16296 (N_16296,N_15012,N_15495);
xor U16297 (N_16297,N_14647,N_14366);
or U16298 (N_16298,N_15952,N_15873);
nor U16299 (N_16299,N_14455,N_15404);
and U16300 (N_16300,N_15591,N_14639);
xnor U16301 (N_16301,N_15021,N_15222);
nand U16302 (N_16302,N_14182,N_14621);
nor U16303 (N_16303,N_14983,N_14949);
nand U16304 (N_16304,N_15276,N_14874);
nor U16305 (N_16305,N_14443,N_15358);
nor U16306 (N_16306,N_14538,N_15511);
xnor U16307 (N_16307,N_15441,N_15166);
nor U16308 (N_16308,N_14030,N_14326);
nand U16309 (N_16309,N_14897,N_14047);
nor U16310 (N_16310,N_15966,N_14409);
or U16311 (N_16311,N_15041,N_15259);
nor U16312 (N_16312,N_14770,N_14969);
nor U16313 (N_16313,N_15199,N_15440);
and U16314 (N_16314,N_15899,N_15003);
and U16315 (N_16315,N_15114,N_14990);
nor U16316 (N_16316,N_15605,N_15317);
nand U16317 (N_16317,N_14586,N_14296);
xor U16318 (N_16318,N_14840,N_14142);
xor U16319 (N_16319,N_15712,N_14943);
xnor U16320 (N_16320,N_14851,N_15906);
and U16321 (N_16321,N_14689,N_15037);
nand U16322 (N_16322,N_15433,N_14292);
nor U16323 (N_16323,N_15242,N_15418);
or U16324 (N_16324,N_14242,N_14833);
and U16325 (N_16325,N_15997,N_14122);
nor U16326 (N_16326,N_14861,N_14539);
and U16327 (N_16327,N_15813,N_15669);
nand U16328 (N_16328,N_14475,N_15649);
and U16329 (N_16329,N_15140,N_14746);
nand U16330 (N_16330,N_15719,N_15025);
nor U16331 (N_16331,N_15225,N_15465);
xnor U16332 (N_16332,N_14526,N_15239);
or U16333 (N_16333,N_15034,N_14741);
and U16334 (N_16334,N_15161,N_14422);
or U16335 (N_16335,N_15194,N_15350);
and U16336 (N_16336,N_15348,N_15420);
and U16337 (N_16337,N_14962,N_14821);
nor U16338 (N_16338,N_14591,N_14524);
nor U16339 (N_16339,N_14817,N_14645);
xnor U16340 (N_16340,N_15141,N_15193);
nor U16341 (N_16341,N_15330,N_15241);
or U16342 (N_16342,N_14423,N_15834);
and U16343 (N_16343,N_15202,N_14447);
or U16344 (N_16344,N_15730,N_14799);
nor U16345 (N_16345,N_15627,N_14021);
and U16346 (N_16346,N_15321,N_15445);
nor U16347 (N_16347,N_14500,N_15240);
nand U16348 (N_16348,N_15223,N_14221);
or U16349 (N_16349,N_14431,N_14673);
or U16350 (N_16350,N_15005,N_15638);
xnor U16351 (N_16351,N_14545,N_15482);
nand U16352 (N_16352,N_14666,N_14426);
nand U16353 (N_16353,N_14774,N_14130);
and U16354 (N_16354,N_14991,N_15671);
xor U16355 (N_16355,N_15183,N_15071);
nor U16356 (N_16356,N_14336,N_14218);
or U16357 (N_16357,N_14017,N_15228);
or U16358 (N_16358,N_15299,N_14926);
xnor U16359 (N_16359,N_14723,N_15187);
nor U16360 (N_16360,N_14140,N_14659);
nor U16361 (N_16361,N_15070,N_15819);
and U16362 (N_16362,N_14857,N_15163);
nand U16363 (N_16363,N_14785,N_14103);
and U16364 (N_16364,N_15470,N_14665);
xnor U16365 (N_16365,N_15270,N_14274);
nand U16366 (N_16366,N_14068,N_14138);
nor U16367 (N_16367,N_14766,N_15955);
nand U16368 (N_16368,N_14205,N_14265);
xor U16369 (N_16369,N_14340,N_15307);
and U16370 (N_16370,N_14458,N_15984);
xor U16371 (N_16371,N_15118,N_14642);
or U16372 (N_16372,N_14627,N_15466);
or U16373 (N_16373,N_15634,N_15587);
and U16374 (N_16374,N_14699,N_15959);
and U16375 (N_16375,N_14410,N_15706);
xor U16376 (N_16376,N_15725,N_15268);
and U16377 (N_16377,N_14527,N_15642);
nand U16378 (N_16378,N_14951,N_14323);
xor U16379 (N_16379,N_14779,N_15499);
or U16380 (N_16380,N_14588,N_15227);
nand U16381 (N_16381,N_14263,N_15858);
or U16382 (N_16382,N_14597,N_14044);
and U16383 (N_16383,N_14610,N_14153);
or U16384 (N_16384,N_14832,N_14129);
and U16385 (N_16385,N_15539,N_15329);
xor U16386 (N_16386,N_15245,N_15142);
nand U16387 (N_16387,N_15213,N_14733);
xor U16388 (N_16388,N_15192,N_14269);
and U16389 (N_16389,N_15779,N_15177);
xor U16390 (N_16390,N_15457,N_15944);
or U16391 (N_16391,N_14064,N_15739);
and U16392 (N_16392,N_14433,N_15060);
nand U16393 (N_16393,N_15660,N_14946);
and U16394 (N_16394,N_14297,N_14041);
nor U16395 (N_16395,N_15272,N_15826);
or U16396 (N_16396,N_15345,N_14982);
xnor U16397 (N_16397,N_15697,N_15368);
nand U16398 (N_16398,N_14976,N_14015);
nand U16399 (N_16399,N_15516,N_15747);
or U16400 (N_16400,N_14465,N_14147);
or U16401 (N_16401,N_15009,N_14984);
and U16402 (N_16402,N_15548,N_14987);
nor U16403 (N_16403,N_14880,N_15271);
xnor U16404 (N_16404,N_15693,N_15197);
nor U16405 (N_16405,N_15479,N_14214);
nand U16406 (N_16406,N_14477,N_15231);
nor U16407 (N_16407,N_15729,N_14788);
or U16408 (N_16408,N_14071,N_14590);
nand U16409 (N_16409,N_15289,N_14281);
nand U16410 (N_16410,N_15126,N_15031);
xnor U16411 (N_16411,N_15673,N_15266);
nand U16412 (N_16412,N_15184,N_15260);
and U16413 (N_16413,N_14974,N_14356);
nand U16414 (N_16414,N_15734,N_14507);
or U16415 (N_16415,N_15716,N_15077);
and U16416 (N_16416,N_15870,N_14197);
xor U16417 (N_16417,N_14810,N_14705);
and U16418 (N_16418,N_15206,N_15425);
xor U16419 (N_16419,N_14556,N_14997);
nor U16420 (N_16420,N_15492,N_15728);
and U16421 (N_16421,N_14386,N_14885);
and U16422 (N_16422,N_15755,N_15752);
nor U16423 (N_16423,N_15044,N_15871);
or U16424 (N_16424,N_14609,N_15910);
nand U16425 (N_16425,N_15939,N_14432);
nand U16426 (N_16426,N_14061,N_15898);
nand U16427 (N_16427,N_14868,N_14227);
and U16428 (N_16428,N_14028,N_14181);
nor U16429 (N_16429,N_15783,N_14403);
xor U16430 (N_16430,N_15108,N_14453);
xor U16431 (N_16431,N_15855,N_14282);
and U16432 (N_16432,N_15700,N_15679);
xor U16433 (N_16433,N_15969,N_15881);
xor U16434 (N_16434,N_15090,N_14853);
xnor U16435 (N_16435,N_15459,N_14194);
or U16436 (N_16436,N_14720,N_14481);
xnor U16437 (N_16437,N_14107,N_14098);
or U16438 (N_16438,N_14883,N_14011);
and U16439 (N_16439,N_14321,N_14334);
nand U16440 (N_16440,N_14126,N_14753);
or U16441 (N_16441,N_14502,N_15735);
and U16442 (N_16442,N_15973,N_14910);
xor U16443 (N_16443,N_14229,N_14254);
nand U16444 (N_16444,N_14830,N_14381);
nand U16445 (N_16445,N_14752,N_15159);
or U16446 (N_16446,N_15600,N_14523);
nand U16447 (N_16447,N_15284,N_14641);
or U16448 (N_16448,N_15411,N_14248);
nor U16449 (N_16449,N_15128,N_14661);
or U16450 (N_16450,N_15094,N_14284);
and U16451 (N_16451,N_15269,N_15742);
and U16452 (N_16452,N_14942,N_14550);
nand U16453 (N_16453,N_14676,N_14812);
xnor U16454 (N_16454,N_14100,N_14772);
nand U16455 (N_16455,N_15167,N_14023);
or U16456 (N_16456,N_14244,N_14906);
nand U16457 (N_16457,N_14915,N_14854);
nand U16458 (N_16458,N_14818,N_15656);
and U16459 (N_16459,N_14511,N_14090);
and U16460 (N_16460,N_15030,N_15532);
nand U16461 (N_16461,N_15121,N_15863);
nor U16462 (N_16462,N_14530,N_14291);
and U16463 (N_16463,N_15303,N_15980);
and U16464 (N_16464,N_15816,N_14371);
nand U16465 (N_16465,N_15116,N_15438);
nand U16466 (N_16466,N_14012,N_14748);
nand U16467 (N_16467,N_14161,N_15526);
nand U16468 (N_16468,N_15894,N_14359);
nand U16469 (N_16469,N_15246,N_15637);
nand U16470 (N_16470,N_15027,N_14060);
or U16471 (N_16471,N_14119,N_15460);
and U16472 (N_16472,N_15252,N_14089);
nand U16473 (N_16473,N_15661,N_14933);
nor U16474 (N_16474,N_14931,N_15695);
nor U16475 (N_16475,N_15546,N_14178);
or U16476 (N_16476,N_15452,N_15085);
xor U16477 (N_16477,N_15603,N_14615);
nand U16478 (N_16478,N_14681,N_15727);
and U16479 (N_16479,N_14391,N_15884);
or U16480 (N_16480,N_15461,N_15232);
or U16481 (N_16481,N_15521,N_15337);
or U16482 (N_16482,N_15405,N_14602);
xnor U16483 (N_16483,N_14886,N_15580);
xnor U16484 (N_16484,N_15886,N_14268);
nor U16485 (N_16485,N_15844,N_15098);
and U16486 (N_16486,N_14935,N_14293);
nor U16487 (N_16487,N_14057,N_14166);
nor U16488 (N_16488,N_15731,N_14368);
xnor U16489 (N_16489,N_15489,N_14373);
or U16490 (N_16490,N_14503,N_14819);
and U16491 (N_16491,N_15571,N_15593);
nand U16492 (N_16492,N_14184,N_15237);
or U16493 (N_16493,N_14456,N_15152);
nand U16494 (N_16494,N_15283,N_14549);
nand U16495 (N_16495,N_15857,N_15048);
or U16496 (N_16496,N_15416,N_15803);
and U16497 (N_16497,N_14379,N_15653);
and U16498 (N_16498,N_15531,N_15621);
and U16499 (N_16499,N_14875,N_14797);
and U16500 (N_16500,N_15948,N_15170);
xor U16501 (N_16501,N_15300,N_14469);
and U16502 (N_16502,N_15574,N_15490);
nor U16503 (N_16503,N_14049,N_14136);
and U16504 (N_16504,N_15715,N_15230);
xnor U16505 (N_16505,N_14514,N_14402);
nor U16506 (N_16506,N_15565,N_14613);
and U16507 (N_16507,N_15073,N_15074);
xor U16508 (N_16508,N_14353,N_14630);
or U16509 (N_16509,N_14717,N_14979);
or U16510 (N_16510,N_14020,N_15286);
xor U16511 (N_16511,N_15277,N_14496);
nor U16512 (N_16512,N_15282,N_14909);
nor U16513 (N_16513,N_15162,N_14375);
nor U16514 (N_16514,N_14115,N_15352);
nand U16515 (N_16515,N_15746,N_14850);
or U16516 (N_16516,N_14518,N_15774);
nand U16517 (N_16517,N_14279,N_15920);
or U16518 (N_16518,N_14338,N_14430);
xor U16519 (N_16519,N_14216,N_15454);
nor U16520 (N_16520,N_14400,N_14319);
xnor U16521 (N_16521,N_15889,N_15385);
nor U16522 (N_16522,N_15782,N_14684);
nor U16523 (N_16523,N_14081,N_15380);
nor U16524 (N_16524,N_15778,N_14171);
nand U16525 (N_16525,N_14650,N_14711);
nor U16526 (N_16526,N_14873,N_15562);
xnor U16527 (N_16527,N_15488,N_14325);
and U16528 (N_16528,N_14554,N_14348);
or U16529 (N_16529,N_14288,N_14258);
or U16530 (N_16530,N_14261,N_14568);
nor U16531 (N_16531,N_14005,N_15869);
xor U16532 (N_16532,N_15510,N_15829);
nand U16533 (N_16533,N_15839,N_14343);
nand U16534 (N_16534,N_14491,N_14249);
xnor U16535 (N_16535,N_14203,N_15437);
or U16536 (N_16536,N_14277,N_14995);
nand U16537 (N_16537,N_15201,N_15309);
and U16538 (N_16538,N_14025,N_15926);
nand U16539 (N_16539,N_15911,N_14820);
nand U16540 (N_16540,N_14793,N_14034);
nand U16541 (N_16541,N_15624,N_15528);
or U16542 (N_16542,N_15610,N_15958);
xnor U16543 (N_16543,N_15209,N_14290);
nor U16544 (N_16544,N_15151,N_15828);
nand U16545 (N_16545,N_14957,N_15522);
nand U16546 (N_16546,N_14654,N_15477);
nor U16547 (N_16547,N_15831,N_15160);
xor U16548 (N_16548,N_14464,N_15985);
and U16549 (N_16549,N_14607,N_14944);
and U16550 (N_16550,N_15147,N_14124);
or U16551 (N_16551,N_14546,N_14048);
and U16552 (N_16552,N_15647,N_14390);
and U16553 (N_16553,N_15840,N_15907);
nor U16554 (N_16554,N_14964,N_15349);
nor U16555 (N_16555,N_14577,N_15564);
or U16556 (N_16556,N_14598,N_15513);
and U16557 (N_16557,N_15332,N_14593);
and U16558 (N_16558,N_14544,N_15749);
nor U16559 (N_16559,N_14887,N_14393);
nand U16560 (N_16560,N_15750,N_15664);
or U16561 (N_16561,N_15644,N_15471);
xnor U16562 (N_16562,N_15389,N_14594);
xor U16563 (N_16563,N_14245,N_15364);
nand U16564 (N_16564,N_14200,N_14435);
and U16565 (N_16565,N_15835,N_15374);
nand U16566 (N_16566,N_14339,N_15632);
xor U16567 (N_16567,N_14150,N_15171);
or U16568 (N_16568,N_15949,N_15409);
nor U16569 (N_16569,N_14986,N_15261);
nand U16570 (N_16570,N_14347,N_15382);
nand U16571 (N_16571,N_14201,N_15717);
xor U16572 (N_16572,N_15965,N_14314);
and U16573 (N_16573,N_15447,N_14151);
xor U16574 (N_16574,N_14977,N_15990);
or U16575 (N_16575,N_14956,N_14862);
and U16576 (N_16576,N_15304,N_14019);
nand U16577 (N_16577,N_14073,N_14232);
nand U16578 (N_16578,N_14709,N_14457);
nor U16579 (N_16579,N_14728,N_14569);
or U16580 (N_16580,N_14316,N_15509);
nand U16581 (N_16581,N_14051,N_14189);
xnor U16582 (N_16582,N_14063,N_15937);
or U16583 (N_16583,N_14682,N_15453);
xor U16584 (N_16584,N_15280,N_14123);
nor U16585 (N_16585,N_15613,N_15267);
and U16586 (N_16586,N_15536,N_14210);
or U16587 (N_16587,N_15618,N_15180);
nor U16588 (N_16588,N_15757,N_14209);
nor U16589 (N_16589,N_15811,N_15175);
nor U16590 (N_16590,N_14648,N_15320);
nor U16591 (N_16591,N_15761,N_14163);
xnor U16592 (N_16592,N_14287,N_15862);
nor U16593 (N_16593,N_14036,N_15847);
nand U16594 (N_16594,N_15876,N_15711);
xnor U16595 (N_16595,N_14561,N_14001);
nand U16596 (N_16596,N_14411,N_15308);
nor U16597 (N_16597,N_14871,N_14631);
or U16598 (N_16598,N_14914,N_15173);
or U16599 (N_16599,N_15850,N_14234);
nor U16600 (N_16600,N_14087,N_15472);
and U16601 (N_16601,N_15567,N_15467);
or U16602 (N_16602,N_15326,N_14808);
xnor U16603 (N_16603,N_14162,N_15040);
or U16604 (N_16604,N_14805,N_14204);
nor U16605 (N_16605,N_14540,N_15879);
xnor U16606 (N_16606,N_14608,N_14831);
nand U16607 (N_16607,N_15585,N_14738);
and U16608 (N_16608,N_15428,N_14938);
nor U16609 (N_16609,N_14038,N_14378);
xnor U16610 (N_16610,N_14054,N_14298);
or U16611 (N_16611,N_15288,N_15366);
and U16612 (N_16612,N_14658,N_15218);
xor U16613 (N_16613,N_15628,N_14614);
or U16614 (N_16614,N_14369,N_15061);
xor U16615 (N_16615,N_15945,N_14548);
nand U16616 (N_16616,N_15417,N_14131);
xnor U16617 (N_16617,N_15158,N_14712);
or U16618 (N_16618,N_14565,N_15338);
xor U16619 (N_16619,N_15583,N_14822);
nand U16620 (N_16620,N_15982,N_15449);
or U16621 (N_16621,N_14299,N_14534);
xor U16622 (N_16622,N_14807,N_15641);
and U16623 (N_16623,N_14623,N_14842);
or U16624 (N_16624,N_14445,N_15233);
xor U16625 (N_16625,N_14881,N_15971);
nor U16626 (N_16626,N_15226,N_15065);
nor U16627 (N_16627,N_15810,N_15390);
and U16628 (N_16628,N_14600,N_14579);
or U16629 (N_16629,N_15843,N_15273);
and U16630 (N_16630,N_14512,N_14042);
nand U16631 (N_16631,N_14160,N_14417);
nand U16632 (N_16632,N_14231,N_14884);
xor U16633 (N_16633,N_15559,N_14387);
nand U16634 (N_16634,N_14782,N_14903);
and U16635 (N_16635,N_15257,N_15764);
or U16636 (N_16636,N_15256,N_14616);
or U16637 (N_16637,N_14564,N_14870);
xnor U16638 (N_16638,N_14452,N_15264);
nor U16639 (N_16639,N_14628,N_15994);
or U16640 (N_16640,N_15343,N_14846);
nand U16641 (N_16641,N_14776,N_14917);
xor U16642 (N_16642,N_15013,N_14215);
or U16643 (N_16643,N_14836,N_14065);
nor U16644 (N_16644,N_14535,N_14865);
and U16645 (N_16645,N_14156,N_15251);
nand U16646 (N_16646,N_15691,N_14533);
nor U16647 (N_16647,N_14667,N_14053);
or U16648 (N_16648,N_15685,N_15989);
nor U16649 (N_16649,N_14803,N_15612);
or U16650 (N_16650,N_15602,N_15181);
xnor U16651 (N_16651,N_15429,N_14179);
nor U16652 (N_16652,N_15714,N_14374);
or U16653 (N_16653,N_14508,N_14207);
nand U16654 (N_16654,N_15244,N_14837);
and U16655 (N_16655,N_14778,N_15934);
nand U16656 (N_16656,N_14529,N_15999);
or U16657 (N_16657,N_15551,N_14490);
xor U16658 (N_16658,N_15890,N_14495);
xnor U16659 (N_16659,N_15785,N_14828);
nand U16660 (N_16660,N_15430,N_14259);
nor U16661 (N_16661,N_14494,N_14266);
nand U16662 (N_16662,N_15403,N_15004);
or U16663 (N_16663,N_14271,N_15576);
xnor U16664 (N_16664,N_14547,N_15474);
and U16665 (N_16665,N_14437,N_14612);
xnor U16666 (N_16666,N_15915,N_15279);
and U16667 (N_16667,N_15258,N_14767);
xnor U16668 (N_16668,N_14759,N_15179);
or U16669 (N_16669,N_15046,N_14558);
or U16670 (N_16670,N_15520,N_15221);
nor U16671 (N_16671,N_15473,N_14177);
and U16672 (N_16672,N_15553,N_15914);
or U16673 (N_16673,N_15838,N_15392);
or U16674 (N_16674,N_15541,N_15533);
or U16675 (N_16675,N_15794,N_15415);
xor U16676 (N_16676,N_14419,N_15106);
nor U16677 (N_16677,N_14758,N_14405);
or U16678 (N_16678,N_15547,N_14335);
and U16679 (N_16679,N_15292,N_14333);
or U16680 (N_16680,N_14791,N_14327);
nand U16681 (N_16681,N_14395,N_15455);
and U16682 (N_16682,N_15566,N_15250);
xnor U16683 (N_16683,N_15655,N_14404);
and U16684 (N_16684,N_14736,N_14578);
and U16685 (N_16685,N_14190,N_14199);
nor U16686 (N_16686,N_15799,N_15000);
and U16687 (N_16687,N_14575,N_14342);
or U16688 (N_16688,N_14719,N_14801);
or U16689 (N_16689,N_15601,N_14617);
and U16690 (N_16690,N_14345,N_14622);
nor U16691 (N_16691,N_14954,N_14536);
or U16692 (N_16692,N_15501,N_15787);
and U16693 (N_16693,N_14280,N_14388);
and U16694 (N_16694,N_14707,N_14070);
or U16695 (N_16695,N_14936,N_15064);
nand U16696 (N_16696,N_15577,N_15883);
nand U16697 (N_16697,N_14867,N_15748);
nand U16698 (N_16698,N_14252,N_15293);
nand U16699 (N_16699,N_15081,N_14109);
or U16700 (N_16700,N_15998,N_14446);
or U16701 (N_16701,N_14606,N_14922);
and U16702 (N_16702,N_14257,N_14794);
xor U16703 (N_16703,N_14429,N_15594);
xor U16704 (N_16704,N_15630,N_14112);
or U16705 (N_16705,N_15689,N_15900);
xnor U16706 (N_16706,N_15016,N_14233);
and U16707 (N_16707,N_15720,N_15931);
xnor U16708 (N_16708,N_14678,N_14958);
and U16709 (N_16709,N_14256,N_15823);
nor U16710 (N_16710,N_14476,N_15569);
xnor U16711 (N_16711,N_15784,N_14438);
nand U16712 (N_16712,N_15699,N_15275);
xnor U16713 (N_16713,N_15082,N_15424);
nand U16714 (N_16714,N_15376,N_15483);
and U16715 (N_16715,N_15038,N_15590);
nand U16716 (N_16716,N_15705,N_15895);
nand U16717 (N_16717,N_15854,N_14908);
nand U16718 (N_16718,N_15848,N_14351);
and U16719 (N_16719,N_15217,N_15505);
nor U16720 (N_16720,N_14013,N_15770);
xor U16721 (N_16721,N_14196,N_15923);
xor U16722 (N_16722,N_15681,N_14185);
nor U16723 (N_16723,N_14193,N_14843);
nand U16724 (N_16724,N_15827,N_14601);
xnor U16725 (N_16725,N_14921,N_14552);
xnor U16726 (N_16726,N_15011,N_15806);
xnor U16727 (N_16727,N_15759,N_15861);
nand U16728 (N_16728,N_15537,N_14105);
and U16729 (N_16729,N_14085,N_14953);
nor U16730 (N_16730,N_15726,N_14219);
xnor U16731 (N_16731,N_14895,N_14963);
and U16732 (N_16732,N_15120,N_15942);
nand U16733 (N_16733,N_14879,N_15019);
and U16734 (N_16734,N_14337,N_15129);
or U16735 (N_16735,N_15598,N_15775);
nand U16736 (N_16736,N_14220,N_15668);
nor U16737 (N_16737,N_15491,N_14900);
or U16738 (N_16738,N_15319,N_14427);
nand U16739 (N_16739,N_14144,N_14003);
and U16740 (N_16740,N_14440,N_15740);
xor U16741 (N_16741,N_15607,N_14040);
or U16742 (N_16742,N_14792,N_14289);
xor U16743 (N_16743,N_14839,N_15650);
xnor U16744 (N_16744,N_14238,N_15360);
or U16745 (N_16745,N_15301,N_15487);
nand U16746 (N_16746,N_15190,N_14740);
xor U16747 (N_16747,N_14474,N_15427);
or U16748 (N_16748,N_15866,N_14784);
nand U16749 (N_16749,N_15957,N_14702);
xnor U16750 (N_16750,N_15410,N_14052);
and U16751 (N_16751,N_15033,N_14154);
or U16752 (N_16752,N_14891,N_15328);
nor U16753 (N_16753,N_15860,N_14239);
nand U16754 (N_16754,N_15315,N_15369);
or U16755 (N_16755,N_14159,N_14312);
nand U16756 (N_16756,N_15422,N_14823);
nand U16757 (N_16757,N_15970,N_14620);
nand U16758 (N_16758,N_15933,N_15874);
nor U16759 (N_16759,N_14845,N_15493);
xor U16760 (N_16760,N_15413,N_15131);
nor U16761 (N_16761,N_14695,N_14092);
and U16762 (N_16762,N_14004,N_14407);
xnor U16763 (N_16763,N_15557,N_15370);
xor U16764 (N_16764,N_14149,N_15397);
and U16765 (N_16765,N_15558,N_15614);
xor U16766 (N_16766,N_14814,N_15804);
or U16767 (N_16767,N_15897,N_14213);
xor U16768 (N_16768,N_15375,N_15595);
xnor U16769 (N_16769,N_14075,N_14383);
nor U16770 (N_16770,N_14223,N_14361);
nor U16771 (N_16771,N_14835,N_14226);
or U16772 (N_16772,N_15832,N_14180);
and U16773 (N_16773,N_15406,N_15444);
xor U16774 (N_16774,N_15893,N_15314);
nor U16775 (N_16775,N_14078,N_14994);
nor U16776 (N_16776,N_14670,N_14307);
and U16777 (N_16777,N_14890,N_14815);
xnor U16778 (N_16778,N_14743,N_15575);
nand U16779 (N_16779,N_14077,N_14955);
nor U16780 (N_16780,N_14589,N_14640);
nand U16781 (N_16781,N_15692,N_14646);
nand U16782 (N_16782,N_14965,N_15837);
xnor U16783 (N_16783,N_14562,N_15431);
xor U16784 (N_16784,N_14532,N_14583);
nor U16785 (N_16785,N_15903,N_14744);
or U16786 (N_16786,N_14183,N_14696);
xnor U16787 (N_16787,N_15333,N_15099);
nand U16788 (N_16788,N_14198,N_15351);
nand U16789 (N_16789,N_15122,N_14479);
or U16790 (N_16790,N_15310,N_15701);
nand U16791 (N_16791,N_14118,N_14985);
and U16792 (N_16792,N_14080,N_14826);
nand U16793 (N_16793,N_14225,N_15987);
nor U16794 (N_16794,N_14859,N_15578);
xor U16795 (N_16795,N_15891,N_15924);
or U16796 (N_16796,N_14809,N_14595);
nor U16797 (N_16797,N_15414,N_15462);
nand U16798 (N_16798,N_15786,N_14367);
or U16799 (N_16799,N_14320,N_15753);
xor U16800 (N_16800,N_15667,N_15682);
xnor U16801 (N_16801,N_15756,N_15611);
and U16802 (N_16802,N_14653,N_15249);
and U16803 (N_16803,N_15960,N_15790);
nor U16804 (N_16804,N_15238,N_14493);
xnor U16805 (N_16805,N_14683,N_14993);
or U16806 (N_16806,N_15464,N_14416);
xnor U16807 (N_16807,N_15426,N_14141);
xnor U16808 (N_16808,N_15545,N_15925);
nand U16809 (N_16809,N_14510,N_14585);
nor U16810 (N_16810,N_14901,N_15963);
xnor U16811 (N_16811,N_15581,N_14217);
or U16812 (N_16812,N_14940,N_14519);
and U16813 (N_16813,N_15946,N_15294);
nand U16814 (N_16814,N_14441,N_15968);
and U16815 (N_16815,N_14285,N_14581);
xor U16816 (N_16816,N_15327,N_15821);
and U16817 (N_16817,N_14482,N_14097);
xnor U16818 (N_16818,N_14331,N_15412);
and U16819 (N_16819,N_14787,N_15974);
or U16820 (N_16820,N_14246,N_15164);
xor U16821 (N_16821,N_15215,N_15666);
or U16822 (N_16822,N_15916,N_15708);
nand U16823 (N_16823,N_14856,N_14825);
nand U16824 (N_16824,N_14703,N_15176);
nand U16825 (N_16825,N_15964,N_14996);
and U16826 (N_16826,N_15387,N_14660);
and U16827 (N_16827,N_15586,N_14838);
xor U16828 (N_16828,N_14567,N_15182);
nand U16829 (N_16829,N_15543,N_15486);
or U16830 (N_16830,N_14247,N_14024);
or U16831 (N_16831,N_14272,N_14167);
nor U16832 (N_16832,N_15367,N_15568);
nor U16833 (N_16833,N_15514,N_15095);
nor U16834 (N_16834,N_15640,N_15281);
and U16835 (N_16835,N_15852,N_15400);
nor U16836 (N_16836,N_14170,N_15344);
or U16837 (N_16837,N_15646,N_15633);
xnor U16838 (N_16838,N_14722,N_15512);
or U16839 (N_16839,N_15645,N_15841);
or U16840 (N_16840,N_15020,N_15902);
or U16841 (N_16841,N_14489,N_15680);
and U16842 (N_16842,N_14576,N_14675);
and U16843 (N_16843,N_15927,N_15117);
or U16844 (N_16844,N_15191,N_14084);
nor U16845 (N_16845,N_15371,N_14363);
and U16846 (N_16846,N_14498,N_15185);
xor U16847 (N_16847,N_14385,N_14434);
nor U16848 (N_16848,N_15137,N_14398);
nand U16849 (N_16849,N_14132,N_14737);
nor U16850 (N_16850,N_14760,N_14761);
nand U16851 (N_16851,N_15149,N_15743);
xor U16852 (N_16852,N_15812,N_14735);
or U16853 (N_16853,N_15049,N_15616);
and U16854 (N_16854,N_14755,N_14664);
and U16855 (N_16855,N_15104,N_15930);
xor U16856 (N_16856,N_14506,N_14158);
nand U16857 (N_16857,N_15767,N_15853);
nand U16858 (N_16858,N_14313,N_14497);
and U16859 (N_16859,N_15325,N_14563);
or U16860 (N_16860,N_15704,N_14006);
or U16861 (N_16861,N_14318,N_14848);
and U16862 (N_16862,N_15353,N_14212);
nor U16863 (N_16863,N_14324,N_15709);
nor U16864 (N_16864,N_14439,N_14026);
and U16865 (N_16865,N_15502,N_15291);
nor U16866 (N_16866,N_14344,N_14559);
nand U16867 (N_16867,N_15059,N_14357);
and U16868 (N_16868,N_15710,N_15967);
nor U16869 (N_16869,N_15204,N_14893);
nand U16870 (N_16870,N_15401,N_14380);
and U16871 (N_16871,N_14037,N_15659);
xor U16872 (N_16872,N_15754,N_14173);
and U16873 (N_16873,N_15198,N_14079);
and U16874 (N_16874,N_15278,N_15297);
nor U16875 (N_16875,N_14192,N_14045);
nand U16876 (N_16876,N_15100,N_14027);
and U16877 (N_16877,N_14655,N_15093);
or U16878 (N_16878,N_14863,N_15207);
nand U16879 (N_16879,N_14669,N_14104);
nor U16880 (N_16880,N_14134,N_15648);
nor U16881 (N_16881,N_15880,N_15789);
nor U16882 (N_16882,N_14372,N_15062);
nand U16883 (N_16883,N_15507,N_15888);
nand U16884 (N_16884,N_14697,N_15496);
nor U16885 (N_16885,N_14152,N_15781);
nand U16886 (N_16886,N_14067,N_15718);
nor U16887 (N_16887,N_15347,N_15504);
or U16888 (N_16888,N_14972,N_15092);
xnor U16889 (N_16889,N_15570,N_14927);
xnor U16890 (N_16890,N_15745,N_15556);
and U16891 (N_16891,N_14961,N_15043);
nor U16892 (N_16892,N_15346,N_14691);
xnor U16893 (N_16893,N_15135,N_15365);
nand U16894 (N_16894,N_15599,N_15196);
or U16895 (N_16895,N_14195,N_14757);
xor U16896 (N_16896,N_15552,N_15208);
nand U16897 (N_16897,N_15384,N_14237);
or U16898 (N_16898,N_15956,N_15694);
nand U16899 (N_16899,N_14172,N_15978);
or U16900 (N_16900,N_15243,N_15913);
xnor U16901 (N_16901,N_14328,N_14804);
or U16902 (N_16902,N_15214,N_15028);
nor U16903 (N_16903,N_14346,N_15654);
xnor U16904 (N_16904,N_15408,N_14008);
and U16905 (N_16905,N_14406,N_14685);
xnor U16906 (N_16906,N_15017,N_14250);
xor U16907 (N_16907,N_14033,N_15354);
xnor U16908 (N_16908,N_15312,N_15932);
and U16909 (N_16909,N_15818,N_15362);
xor U16910 (N_16910,N_14186,N_15849);
nand U16911 (N_16911,N_14765,N_14834);
xnor U16912 (N_16912,N_15274,N_15663);
nor U16913 (N_16913,N_14570,N_15904);
and U16914 (N_16914,N_15560,N_14016);
nand U16915 (N_16915,N_14255,N_14674);
nand U16916 (N_16916,N_14754,N_14553);
nor U16917 (N_16917,N_15469,N_15050);
and U16918 (N_16918,N_15721,N_14355);
nor U16919 (N_16919,N_15544,N_15468);
xnor U16920 (N_16920,N_15054,N_15917);
or U16921 (N_16921,N_14155,N_14625);
xnor U16922 (N_16922,N_14101,N_15885);
nand U16923 (N_16923,N_15446,N_15683);
and U16924 (N_16924,N_14587,N_14599);
xnor U16925 (N_16925,N_15442,N_15134);
xor U16926 (N_16926,N_15981,N_14605);
and U16927 (N_16927,N_14270,N_14260);
xor U16928 (N_16928,N_14399,N_14305);
nor U16929 (N_16929,N_14629,N_14537);
or U16930 (N_16930,N_14551,N_15652);
xnor U16931 (N_16931,N_14747,N_15235);
and U16932 (N_16932,N_14680,N_15008);
and U16933 (N_16933,N_15067,N_14415);
or U16934 (N_16934,N_15001,N_14145);
and U16935 (N_16935,N_14652,N_15069);
nand U16936 (N_16936,N_15056,N_14721);
or U16937 (N_16937,N_14632,N_14635);
nand U16938 (N_16938,N_15295,N_14934);
nand U16939 (N_16939,N_15529,N_14980);
nor U16940 (N_16940,N_14488,N_14010);
or U16941 (N_16941,N_14501,N_14582);
nand U16942 (N_16942,N_15530,N_15549);
nor U16943 (N_16943,N_15336,N_15212);
nand U16944 (N_16944,N_15423,N_15113);
xor U16945 (N_16945,N_15053,N_15882);
nor U16946 (N_16946,N_15089,N_15363);
nor U16947 (N_16947,N_14866,N_15112);
or U16948 (N_16948,N_14093,N_15316);
nand U16949 (N_16949,N_14734,N_14789);
or U16950 (N_16950,N_15236,N_14690);
and U16951 (N_16951,N_14120,N_14574);
nor U16952 (N_16952,N_15220,N_15211);
nor U16953 (N_16953,N_14306,N_15133);
nand U16954 (N_16954,N_15802,N_15485);
and U16955 (N_16955,N_14148,N_15976);
or U16956 (N_16956,N_15254,N_15793);
and U16957 (N_16957,N_14462,N_14018);
or U16958 (N_16958,N_15670,N_15798);
xor U16959 (N_16959,N_15877,N_15777);
and U16960 (N_16960,N_14633,N_14948);
and U16961 (N_16961,N_14624,N_15015);
or U16962 (N_16962,N_14396,N_15480);
nor U16963 (N_16963,N_14485,N_14638);
xor U16964 (N_16964,N_15102,N_15619);
and U16965 (N_16965,N_14727,N_15950);
xnor U16966 (N_16966,N_14911,N_14059);
nand U16967 (N_16967,N_15651,N_15820);
xor U16968 (N_16968,N_14769,N_15036);
xnor U16969 (N_16969,N_14224,N_15758);
xnor U16970 (N_16970,N_14706,N_15977);
and U16971 (N_16971,N_14454,N_15772);
xnor U16972 (N_16972,N_14726,N_14168);
or U16973 (N_16973,N_14603,N_15153);
and U16974 (N_16974,N_15393,N_15002);
xor U16975 (N_16975,N_15130,N_15815);
or U16976 (N_16976,N_15686,N_15322);
and U16977 (N_16977,N_14076,N_14352);
xnor U16978 (N_16978,N_14133,N_14364);
nand U16979 (N_16979,N_15936,N_14046);
xor U16980 (N_16980,N_14412,N_15796);
or U16981 (N_16981,N_15629,N_15047);
and U16982 (N_16982,N_14981,N_14114);
xor U16983 (N_16983,N_15609,N_15165);
or U16984 (N_16984,N_14088,N_15722);
and U16985 (N_16985,N_15639,N_14596);
xor U16986 (N_16986,N_15773,N_15450);
and U16987 (N_16987,N_14262,N_15079);
xnor U16988 (N_16988,N_14499,N_15024);
nor U16989 (N_16989,N_14082,N_14466);
nor U16990 (N_16990,N_15255,N_15476);
nand U16991 (N_16991,N_14714,N_14966);
nor U16992 (N_16992,N_14692,N_14923);
xnor U16993 (N_16993,N_15157,N_14745);
or U16994 (N_16994,N_15463,N_15953);
or U16995 (N_16995,N_15817,N_14811);
xor U16996 (N_16996,N_15035,N_15091);
nor U16997 (N_16997,N_15791,N_15068);
nand U16998 (N_16998,N_15127,N_15622);
and U16999 (N_16999,N_14191,N_15381);
and U17000 (N_17000,N_15971,N_14868);
or U17001 (N_17001,N_15346,N_15610);
xor U17002 (N_17002,N_15624,N_15960);
and U17003 (N_17003,N_15291,N_14204);
or U17004 (N_17004,N_15851,N_15943);
nand U17005 (N_17005,N_14528,N_14556);
nand U17006 (N_17006,N_14591,N_15591);
and U17007 (N_17007,N_15406,N_15563);
nand U17008 (N_17008,N_15057,N_14032);
nor U17009 (N_17009,N_14142,N_15129);
and U17010 (N_17010,N_15801,N_14289);
or U17011 (N_17011,N_14056,N_14764);
xnor U17012 (N_17012,N_15743,N_15511);
nor U17013 (N_17013,N_15948,N_15877);
xor U17014 (N_17014,N_14620,N_15971);
nand U17015 (N_17015,N_14677,N_14134);
and U17016 (N_17016,N_14904,N_14830);
or U17017 (N_17017,N_15098,N_15864);
and U17018 (N_17018,N_15680,N_15352);
nor U17019 (N_17019,N_15344,N_15765);
xor U17020 (N_17020,N_15870,N_14950);
nand U17021 (N_17021,N_15977,N_15299);
xnor U17022 (N_17022,N_14961,N_14729);
nor U17023 (N_17023,N_15254,N_14197);
nor U17024 (N_17024,N_15291,N_14368);
nand U17025 (N_17025,N_14267,N_14795);
or U17026 (N_17026,N_15689,N_15373);
nand U17027 (N_17027,N_15204,N_14114);
nor U17028 (N_17028,N_15289,N_15341);
nor U17029 (N_17029,N_14157,N_15165);
or U17030 (N_17030,N_15571,N_14112);
nor U17031 (N_17031,N_15723,N_14615);
nor U17032 (N_17032,N_14360,N_15428);
xor U17033 (N_17033,N_15290,N_14558);
nor U17034 (N_17034,N_15180,N_15062);
xor U17035 (N_17035,N_14435,N_14199);
nand U17036 (N_17036,N_14434,N_14334);
or U17037 (N_17037,N_14781,N_14186);
xor U17038 (N_17038,N_14231,N_15195);
nor U17039 (N_17039,N_15934,N_15698);
nand U17040 (N_17040,N_15315,N_15725);
nand U17041 (N_17041,N_14552,N_14781);
and U17042 (N_17042,N_15669,N_15816);
or U17043 (N_17043,N_14115,N_14162);
or U17044 (N_17044,N_15835,N_15590);
and U17045 (N_17045,N_15392,N_14323);
nand U17046 (N_17046,N_15833,N_14820);
and U17047 (N_17047,N_14683,N_15687);
and U17048 (N_17048,N_14868,N_14858);
xnor U17049 (N_17049,N_15483,N_14234);
and U17050 (N_17050,N_14717,N_15520);
or U17051 (N_17051,N_14716,N_14182);
nor U17052 (N_17052,N_14953,N_14962);
and U17053 (N_17053,N_15711,N_15749);
nor U17054 (N_17054,N_14330,N_14226);
nor U17055 (N_17055,N_15923,N_14388);
nor U17056 (N_17056,N_15338,N_14085);
nand U17057 (N_17057,N_14311,N_15957);
nor U17058 (N_17058,N_15804,N_14800);
xor U17059 (N_17059,N_14660,N_15692);
and U17060 (N_17060,N_14560,N_15961);
and U17061 (N_17061,N_15334,N_15841);
xnor U17062 (N_17062,N_15157,N_15801);
and U17063 (N_17063,N_15775,N_15390);
or U17064 (N_17064,N_14691,N_14585);
xor U17065 (N_17065,N_14640,N_15692);
or U17066 (N_17066,N_14725,N_14385);
and U17067 (N_17067,N_15131,N_14257);
and U17068 (N_17068,N_15514,N_15429);
nand U17069 (N_17069,N_14220,N_14491);
xor U17070 (N_17070,N_14779,N_14882);
nor U17071 (N_17071,N_15423,N_14439);
xor U17072 (N_17072,N_14275,N_14287);
and U17073 (N_17073,N_14421,N_14338);
nand U17074 (N_17074,N_15967,N_14238);
xnor U17075 (N_17075,N_14889,N_15347);
nor U17076 (N_17076,N_14176,N_14551);
or U17077 (N_17077,N_14131,N_14294);
or U17078 (N_17078,N_14893,N_14234);
or U17079 (N_17079,N_14454,N_15627);
nand U17080 (N_17080,N_15713,N_14617);
or U17081 (N_17081,N_15026,N_15513);
nor U17082 (N_17082,N_15885,N_15169);
nor U17083 (N_17083,N_15180,N_15603);
nand U17084 (N_17084,N_15021,N_14219);
xor U17085 (N_17085,N_14060,N_15695);
or U17086 (N_17086,N_14808,N_15792);
xnor U17087 (N_17087,N_15633,N_14402);
or U17088 (N_17088,N_14640,N_15647);
nor U17089 (N_17089,N_15325,N_14855);
or U17090 (N_17090,N_14724,N_15734);
and U17091 (N_17091,N_14884,N_14875);
xor U17092 (N_17092,N_14391,N_14532);
or U17093 (N_17093,N_14532,N_14181);
and U17094 (N_17094,N_15970,N_14004);
or U17095 (N_17095,N_14282,N_14411);
or U17096 (N_17096,N_15978,N_15211);
or U17097 (N_17097,N_14404,N_15966);
nand U17098 (N_17098,N_15162,N_14356);
xor U17099 (N_17099,N_14128,N_14605);
xor U17100 (N_17100,N_14270,N_15423);
xor U17101 (N_17101,N_14667,N_14744);
xor U17102 (N_17102,N_14927,N_14269);
xnor U17103 (N_17103,N_15871,N_15389);
or U17104 (N_17104,N_14244,N_14411);
nor U17105 (N_17105,N_15309,N_14979);
and U17106 (N_17106,N_15230,N_14634);
nor U17107 (N_17107,N_14838,N_14562);
or U17108 (N_17108,N_15729,N_15060);
xor U17109 (N_17109,N_14606,N_14030);
or U17110 (N_17110,N_15927,N_15057);
or U17111 (N_17111,N_15279,N_15191);
and U17112 (N_17112,N_15766,N_14898);
nor U17113 (N_17113,N_14306,N_14784);
nor U17114 (N_17114,N_15538,N_15308);
nor U17115 (N_17115,N_15323,N_14543);
or U17116 (N_17116,N_14669,N_15240);
or U17117 (N_17117,N_15519,N_15698);
nand U17118 (N_17118,N_14870,N_14459);
nor U17119 (N_17119,N_14696,N_14326);
nor U17120 (N_17120,N_15236,N_15223);
nor U17121 (N_17121,N_14557,N_15377);
or U17122 (N_17122,N_15103,N_14528);
nand U17123 (N_17123,N_15892,N_15685);
xnor U17124 (N_17124,N_14728,N_14230);
nand U17125 (N_17125,N_15802,N_15241);
or U17126 (N_17126,N_14686,N_15284);
or U17127 (N_17127,N_15864,N_14654);
xnor U17128 (N_17128,N_14000,N_14365);
and U17129 (N_17129,N_15826,N_15695);
or U17130 (N_17130,N_15835,N_15381);
or U17131 (N_17131,N_14515,N_14571);
or U17132 (N_17132,N_15111,N_14756);
nor U17133 (N_17133,N_15379,N_14549);
xor U17134 (N_17134,N_14339,N_14449);
and U17135 (N_17135,N_14552,N_14114);
xor U17136 (N_17136,N_15973,N_15620);
and U17137 (N_17137,N_15064,N_14521);
and U17138 (N_17138,N_15540,N_14898);
nand U17139 (N_17139,N_14838,N_14040);
and U17140 (N_17140,N_15667,N_14318);
nand U17141 (N_17141,N_14269,N_15563);
xnor U17142 (N_17142,N_14258,N_14226);
nand U17143 (N_17143,N_15304,N_15044);
and U17144 (N_17144,N_14991,N_15678);
nor U17145 (N_17145,N_14165,N_15760);
nor U17146 (N_17146,N_15232,N_15836);
nand U17147 (N_17147,N_15152,N_15096);
nand U17148 (N_17148,N_15538,N_14129);
xnor U17149 (N_17149,N_14032,N_15107);
or U17150 (N_17150,N_14816,N_15962);
xnor U17151 (N_17151,N_14987,N_15814);
nand U17152 (N_17152,N_15815,N_14693);
nor U17153 (N_17153,N_15077,N_14234);
and U17154 (N_17154,N_15015,N_15211);
and U17155 (N_17155,N_14085,N_14476);
nand U17156 (N_17156,N_14456,N_15805);
xnor U17157 (N_17157,N_14576,N_14326);
nor U17158 (N_17158,N_14360,N_14019);
or U17159 (N_17159,N_14058,N_15555);
nor U17160 (N_17160,N_14174,N_15550);
nor U17161 (N_17161,N_14674,N_14354);
and U17162 (N_17162,N_14234,N_15175);
nand U17163 (N_17163,N_15336,N_15260);
or U17164 (N_17164,N_14742,N_14406);
or U17165 (N_17165,N_14604,N_15984);
or U17166 (N_17166,N_15458,N_14156);
xor U17167 (N_17167,N_15107,N_14625);
nand U17168 (N_17168,N_14048,N_15090);
and U17169 (N_17169,N_14325,N_14886);
or U17170 (N_17170,N_15202,N_14160);
or U17171 (N_17171,N_14285,N_14465);
xor U17172 (N_17172,N_14541,N_14583);
nand U17173 (N_17173,N_14001,N_14804);
and U17174 (N_17174,N_14302,N_15119);
nor U17175 (N_17175,N_15521,N_14088);
xnor U17176 (N_17176,N_15832,N_14434);
nor U17177 (N_17177,N_15772,N_15940);
nor U17178 (N_17178,N_14648,N_14179);
and U17179 (N_17179,N_14822,N_15280);
and U17180 (N_17180,N_14272,N_14157);
or U17181 (N_17181,N_15473,N_15981);
or U17182 (N_17182,N_15220,N_14417);
or U17183 (N_17183,N_15871,N_15898);
xnor U17184 (N_17184,N_15539,N_15535);
or U17185 (N_17185,N_15535,N_14447);
nor U17186 (N_17186,N_14106,N_14840);
and U17187 (N_17187,N_15135,N_14387);
nor U17188 (N_17188,N_15657,N_14142);
and U17189 (N_17189,N_14564,N_15526);
and U17190 (N_17190,N_15602,N_14442);
and U17191 (N_17191,N_15818,N_15946);
nand U17192 (N_17192,N_14014,N_15921);
nand U17193 (N_17193,N_14558,N_14337);
xor U17194 (N_17194,N_15595,N_14603);
xnor U17195 (N_17195,N_14302,N_15495);
xnor U17196 (N_17196,N_15914,N_14155);
nor U17197 (N_17197,N_14192,N_15268);
xnor U17198 (N_17198,N_15055,N_15024);
xor U17199 (N_17199,N_14565,N_14018);
and U17200 (N_17200,N_14034,N_14789);
xnor U17201 (N_17201,N_15141,N_14053);
and U17202 (N_17202,N_14124,N_14575);
xor U17203 (N_17203,N_15729,N_15220);
nor U17204 (N_17204,N_15799,N_15482);
or U17205 (N_17205,N_15583,N_14767);
or U17206 (N_17206,N_14727,N_14255);
nor U17207 (N_17207,N_14125,N_14768);
and U17208 (N_17208,N_15482,N_15021);
nand U17209 (N_17209,N_14341,N_15943);
and U17210 (N_17210,N_14097,N_15264);
and U17211 (N_17211,N_14649,N_14650);
nor U17212 (N_17212,N_15679,N_15337);
and U17213 (N_17213,N_14779,N_14820);
and U17214 (N_17214,N_15513,N_15011);
xnor U17215 (N_17215,N_14462,N_15927);
nor U17216 (N_17216,N_14759,N_15765);
or U17217 (N_17217,N_15542,N_15201);
or U17218 (N_17218,N_14120,N_14920);
or U17219 (N_17219,N_15851,N_15778);
xor U17220 (N_17220,N_15056,N_15876);
nor U17221 (N_17221,N_15828,N_15456);
and U17222 (N_17222,N_14860,N_15842);
or U17223 (N_17223,N_14124,N_15199);
and U17224 (N_17224,N_15590,N_15087);
xnor U17225 (N_17225,N_15408,N_15337);
xor U17226 (N_17226,N_15801,N_15400);
and U17227 (N_17227,N_15329,N_14464);
and U17228 (N_17228,N_15772,N_14548);
and U17229 (N_17229,N_14255,N_15430);
or U17230 (N_17230,N_14506,N_15265);
xnor U17231 (N_17231,N_14279,N_14827);
nand U17232 (N_17232,N_14343,N_15308);
xnor U17233 (N_17233,N_15076,N_15821);
xor U17234 (N_17234,N_14928,N_14498);
nor U17235 (N_17235,N_14752,N_15059);
or U17236 (N_17236,N_15641,N_14061);
nand U17237 (N_17237,N_15220,N_15074);
nor U17238 (N_17238,N_15369,N_15966);
nand U17239 (N_17239,N_15675,N_15762);
nand U17240 (N_17240,N_14880,N_15060);
or U17241 (N_17241,N_15107,N_14060);
nor U17242 (N_17242,N_14532,N_15215);
nand U17243 (N_17243,N_15280,N_15434);
nor U17244 (N_17244,N_15664,N_15059);
and U17245 (N_17245,N_15841,N_14367);
xnor U17246 (N_17246,N_15150,N_14409);
xnor U17247 (N_17247,N_15108,N_15922);
and U17248 (N_17248,N_15563,N_15356);
nand U17249 (N_17249,N_14285,N_14801);
xor U17250 (N_17250,N_15066,N_15544);
or U17251 (N_17251,N_14274,N_15217);
xor U17252 (N_17252,N_15886,N_14848);
nor U17253 (N_17253,N_14125,N_15121);
xnor U17254 (N_17254,N_15218,N_14825);
nor U17255 (N_17255,N_14281,N_15724);
xor U17256 (N_17256,N_14082,N_14439);
and U17257 (N_17257,N_14325,N_15460);
and U17258 (N_17258,N_14632,N_15116);
and U17259 (N_17259,N_14462,N_15151);
nand U17260 (N_17260,N_14717,N_14547);
nand U17261 (N_17261,N_14383,N_14060);
xor U17262 (N_17262,N_15982,N_14542);
and U17263 (N_17263,N_15136,N_14036);
nand U17264 (N_17264,N_15928,N_14406);
xnor U17265 (N_17265,N_14176,N_15034);
or U17266 (N_17266,N_14947,N_14439);
and U17267 (N_17267,N_15464,N_14299);
and U17268 (N_17268,N_15231,N_14823);
xor U17269 (N_17269,N_14085,N_15348);
or U17270 (N_17270,N_14504,N_14088);
nand U17271 (N_17271,N_14941,N_15301);
xor U17272 (N_17272,N_15515,N_15052);
or U17273 (N_17273,N_15964,N_14173);
or U17274 (N_17274,N_14597,N_15651);
nand U17275 (N_17275,N_15253,N_15440);
and U17276 (N_17276,N_15126,N_14047);
and U17277 (N_17277,N_15035,N_15609);
and U17278 (N_17278,N_15706,N_15435);
nand U17279 (N_17279,N_14738,N_15441);
nand U17280 (N_17280,N_14548,N_15571);
nor U17281 (N_17281,N_15601,N_14445);
and U17282 (N_17282,N_15271,N_15770);
or U17283 (N_17283,N_14754,N_14136);
nor U17284 (N_17284,N_14813,N_14506);
and U17285 (N_17285,N_15557,N_14660);
xor U17286 (N_17286,N_14102,N_14698);
and U17287 (N_17287,N_14125,N_15634);
xor U17288 (N_17288,N_15708,N_14014);
or U17289 (N_17289,N_14088,N_14401);
or U17290 (N_17290,N_15832,N_14021);
nor U17291 (N_17291,N_15499,N_14894);
and U17292 (N_17292,N_15592,N_15588);
nor U17293 (N_17293,N_15421,N_14724);
nand U17294 (N_17294,N_15967,N_14327);
nand U17295 (N_17295,N_14804,N_15915);
xor U17296 (N_17296,N_15214,N_15804);
nand U17297 (N_17297,N_15823,N_14531);
nand U17298 (N_17298,N_15162,N_14278);
or U17299 (N_17299,N_15719,N_15510);
nand U17300 (N_17300,N_14194,N_15947);
or U17301 (N_17301,N_15961,N_15630);
or U17302 (N_17302,N_15800,N_14207);
nor U17303 (N_17303,N_14524,N_14955);
xor U17304 (N_17304,N_14542,N_15545);
nand U17305 (N_17305,N_14719,N_15390);
nand U17306 (N_17306,N_14916,N_14266);
and U17307 (N_17307,N_15119,N_14087);
and U17308 (N_17308,N_15995,N_15148);
nor U17309 (N_17309,N_14807,N_15578);
or U17310 (N_17310,N_14238,N_14101);
nor U17311 (N_17311,N_15258,N_15438);
xnor U17312 (N_17312,N_14479,N_15231);
nand U17313 (N_17313,N_15989,N_15877);
and U17314 (N_17314,N_15709,N_15852);
and U17315 (N_17315,N_14489,N_15503);
or U17316 (N_17316,N_15409,N_14525);
and U17317 (N_17317,N_14363,N_15954);
nor U17318 (N_17318,N_15539,N_15668);
and U17319 (N_17319,N_14008,N_14448);
xnor U17320 (N_17320,N_14919,N_15609);
and U17321 (N_17321,N_14312,N_14768);
xnor U17322 (N_17322,N_15119,N_14137);
or U17323 (N_17323,N_14109,N_15128);
xnor U17324 (N_17324,N_14960,N_14806);
and U17325 (N_17325,N_14994,N_14196);
nor U17326 (N_17326,N_14920,N_15919);
or U17327 (N_17327,N_14521,N_14214);
or U17328 (N_17328,N_14038,N_15078);
nand U17329 (N_17329,N_15294,N_14451);
and U17330 (N_17330,N_14275,N_15709);
nand U17331 (N_17331,N_15700,N_15826);
or U17332 (N_17332,N_14867,N_15148);
xor U17333 (N_17333,N_15191,N_15669);
nor U17334 (N_17334,N_14534,N_14972);
nor U17335 (N_17335,N_14415,N_14615);
xnor U17336 (N_17336,N_15825,N_14158);
and U17337 (N_17337,N_15661,N_15402);
xnor U17338 (N_17338,N_15250,N_15400);
nor U17339 (N_17339,N_14362,N_15939);
nor U17340 (N_17340,N_14789,N_15563);
and U17341 (N_17341,N_14246,N_15655);
or U17342 (N_17342,N_15495,N_14687);
or U17343 (N_17343,N_14219,N_14556);
or U17344 (N_17344,N_15903,N_14972);
xor U17345 (N_17345,N_14557,N_14564);
xnor U17346 (N_17346,N_14444,N_14303);
nor U17347 (N_17347,N_15253,N_15508);
xnor U17348 (N_17348,N_15648,N_14276);
xor U17349 (N_17349,N_14961,N_14339);
and U17350 (N_17350,N_14218,N_15761);
nand U17351 (N_17351,N_14956,N_15836);
xor U17352 (N_17352,N_15655,N_14436);
nand U17353 (N_17353,N_15120,N_14943);
or U17354 (N_17354,N_14828,N_14753);
nor U17355 (N_17355,N_14405,N_14908);
and U17356 (N_17356,N_15931,N_15640);
xor U17357 (N_17357,N_14052,N_14773);
nand U17358 (N_17358,N_14538,N_14806);
nand U17359 (N_17359,N_15657,N_15803);
and U17360 (N_17360,N_15026,N_15620);
nor U17361 (N_17361,N_15499,N_15701);
nor U17362 (N_17362,N_15701,N_14244);
nand U17363 (N_17363,N_14752,N_14342);
and U17364 (N_17364,N_15459,N_14042);
and U17365 (N_17365,N_15050,N_15448);
or U17366 (N_17366,N_15680,N_15791);
xor U17367 (N_17367,N_15769,N_14167);
nand U17368 (N_17368,N_14345,N_15818);
and U17369 (N_17369,N_15362,N_15951);
and U17370 (N_17370,N_14304,N_15463);
and U17371 (N_17371,N_14966,N_14118);
nand U17372 (N_17372,N_14781,N_14605);
or U17373 (N_17373,N_14372,N_15609);
nor U17374 (N_17374,N_15653,N_14316);
xor U17375 (N_17375,N_14356,N_14844);
or U17376 (N_17376,N_14532,N_15452);
xnor U17377 (N_17377,N_15017,N_14065);
xnor U17378 (N_17378,N_15304,N_15654);
and U17379 (N_17379,N_15854,N_14049);
xor U17380 (N_17380,N_14813,N_14474);
xor U17381 (N_17381,N_14019,N_14809);
and U17382 (N_17382,N_15888,N_14608);
or U17383 (N_17383,N_14943,N_15134);
xnor U17384 (N_17384,N_14986,N_14736);
nand U17385 (N_17385,N_15693,N_14830);
or U17386 (N_17386,N_14252,N_15530);
nand U17387 (N_17387,N_15627,N_15229);
nor U17388 (N_17388,N_14149,N_14807);
or U17389 (N_17389,N_14728,N_15167);
xnor U17390 (N_17390,N_14644,N_14203);
nand U17391 (N_17391,N_14556,N_15399);
and U17392 (N_17392,N_14689,N_15115);
or U17393 (N_17393,N_15420,N_14682);
and U17394 (N_17394,N_15104,N_15836);
and U17395 (N_17395,N_14434,N_14129);
or U17396 (N_17396,N_14404,N_14264);
nor U17397 (N_17397,N_14436,N_14989);
nor U17398 (N_17398,N_15710,N_15242);
xnor U17399 (N_17399,N_14521,N_15622);
nand U17400 (N_17400,N_15983,N_15828);
nand U17401 (N_17401,N_14210,N_14197);
and U17402 (N_17402,N_14508,N_15271);
and U17403 (N_17403,N_14421,N_15586);
or U17404 (N_17404,N_15183,N_14860);
nor U17405 (N_17405,N_15235,N_15192);
or U17406 (N_17406,N_15179,N_14971);
nor U17407 (N_17407,N_15737,N_14428);
xnor U17408 (N_17408,N_15244,N_14437);
and U17409 (N_17409,N_15623,N_14074);
and U17410 (N_17410,N_15995,N_14942);
nand U17411 (N_17411,N_14725,N_15503);
xnor U17412 (N_17412,N_15328,N_15365);
or U17413 (N_17413,N_14574,N_15766);
nand U17414 (N_17414,N_14082,N_15090);
or U17415 (N_17415,N_14401,N_15620);
or U17416 (N_17416,N_15725,N_14950);
nor U17417 (N_17417,N_14297,N_15987);
xnor U17418 (N_17418,N_14768,N_14155);
xor U17419 (N_17419,N_15900,N_15569);
nor U17420 (N_17420,N_14694,N_14049);
nor U17421 (N_17421,N_15564,N_15471);
and U17422 (N_17422,N_15342,N_14043);
or U17423 (N_17423,N_14723,N_15021);
or U17424 (N_17424,N_14356,N_15779);
and U17425 (N_17425,N_14173,N_15374);
xor U17426 (N_17426,N_15050,N_15457);
xor U17427 (N_17427,N_14332,N_15303);
nand U17428 (N_17428,N_15943,N_15462);
and U17429 (N_17429,N_15766,N_14906);
xor U17430 (N_17430,N_14537,N_14425);
xor U17431 (N_17431,N_14476,N_15941);
nor U17432 (N_17432,N_14008,N_14348);
nand U17433 (N_17433,N_14526,N_15704);
nand U17434 (N_17434,N_15516,N_15547);
or U17435 (N_17435,N_14141,N_14959);
xor U17436 (N_17436,N_14356,N_15359);
and U17437 (N_17437,N_15542,N_14658);
nand U17438 (N_17438,N_14960,N_14813);
and U17439 (N_17439,N_15959,N_15109);
nor U17440 (N_17440,N_14480,N_14951);
or U17441 (N_17441,N_15332,N_14614);
and U17442 (N_17442,N_15557,N_14250);
and U17443 (N_17443,N_14752,N_15671);
or U17444 (N_17444,N_14092,N_14697);
xor U17445 (N_17445,N_14928,N_14663);
nand U17446 (N_17446,N_15823,N_15689);
and U17447 (N_17447,N_15187,N_15882);
nor U17448 (N_17448,N_15842,N_14792);
xnor U17449 (N_17449,N_15532,N_15862);
xnor U17450 (N_17450,N_15329,N_15533);
nor U17451 (N_17451,N_14191,N_15344);
xnor U17452 (N_17452,N_14499,N_14080);
nand U17453 (N_17453,N_15266,N_14163);
or U17454 (N_17454,N_15419,N_15336);
nand U17455 (N_17455,N_14217,N_14905);
and U17456 (N_17456,N_14427,N_15373);
xnor U17457 (N_17457,N_14473,N_15059);
nand U17458 (N_17458,N_14137,N_14788);
xor U17459 (N_17459,N_15313,N_14154);
or U17460 (N_17460,N_14907,N_14027);
and U17461 (N_17461,N_14115,N_14525);
nand U17462 (N_17462,N_14537,N_14328);
or U17463 (N_17463,N_14329,N_14381);
nor U17464 (N_17464,N_15476,N_14744);
and U17465 (N_17465,N_14407,N_15198);
xor U17466 (N_17466,N_14079,N_14044);
or U17467 (N_17467,N_15923,N_15405);
or U17468 (N_17468,N_14137,N_15771);
nand U17469 (N_17469,N_15788,N_15777);
nor U17470 (N_17470,N_15397,N_15936);
and U17471 (N_17471,N_14468,N_15699);
or U17472 (N_17472,N_15583,N_14552);
xnor U17473 (N_17473,N_14137,N_14155);
xnor U17474 (N_17474,N_14375,N_14392);
nor U17475 (N_17475,N_15076,N_14620);
xor U17476 (N_17476,N_15543,N_15917);
and U17477 (N_17477,N_14349,N_14927);
or U17478 (N_17478,N_15785,N_14233);
xnor U17479 (N_17479,N_15961,N_15329);
xnor U17480 (N_17480,N_14584,N_14673);
xnor U17481 (N_17481,N_15209,N_15100);
nand U17482 (N_17482,N_14595,N_15371);
or U17483 (N_17483,N_14245,N_15688);
or U17484 (N_17484,N_14380,N_15813);
or U17485 (N_17485,N_15799,N_14681);
and U17486 (N_17486,N_14834,N_14194);
nor U17487 (N_17487,N_15894,N_15147);
or U17488 (N_17488,N_15186,N_14331);
or U17489 (N_17489,N_15824,N_15372);
nand U17490 (N_17490,N_15823,N_15424);
nor U17491 (N_17491,N_14666,N_15731);
or U17492 (N_17492,N_14294,N_14960);
xnor U17493 (N_17493,N_15442,N_14877);
nor U17494 (N_17494,N_15537,N_14049);
nor U17495 (N_17495,N_15911,N_14348);
nand U17496 (N_17496,N_15195,N_14691);
or U17497 (N_17497,N_15787,N_14259);
nor U17498 (N_17498,N_15618,N_14359);
or U17499 (N_17499,N_15452,N_15680);
or U17500 (N_17500,N_15035,N_14388);
xnor U17501 (N_17501,N_14041,N_14650);
or U17502 (N_17502,N_14459,N_15425);
and U17503 (N_17503,N_14882,N_15498);
or U17504 (N_17504,N_14263,N_15206);
xor U17505 (N_17505,N_14987,N_15614);
and U17506 (N_17506,N_15759,N_14728);
and U17507 (N_17507,N_15958,N_15010);
nor U17508 (N_17508,N_15754,N_15220);
nor U17509 (N_17509,N_15161,N_14787);
and U17510 (N_17510,N_15213,N_14893);
or U17511 (N_17511,N_15916,N_15709);
and U17512 (N_17512,N_14753,N_15493);
nor U17513 (N_17513,N_15326,N_14273);
or U17514 (N_17514,N_14913,N_14493);
or U17515 (N_17515,N_14697,N_15333);
or U17516 (N_17516,N_15973,N_14781);
xor U17517 (N_17517,N_14773,N_14711);
nor U17518 (N_17518,N_15943,N_15101);
xor U17519 (N_17519,N_14264,N_14373);
xnor U17520 (N_17520,N_14378,N_14081);
nor U17521 (N_17521,N_15486,N_14592);
xnor U17522 (N_17522,N_15846,N_14537);
or U17523 (N_17523,N_14986,N_14299);
and U17524 (N_17524,N_14983,N_15252);
or U17525 (N_17525,N_15928,N_15314);
nor U17526 (N_17526,N_14019,N_14025);
nor U17527 (N_17527,N_15752,N_15732);
nor U17528 (N_17528,N_14023,N_15720);
nand U17529 (N_17529,N_15051,N_14971);
nor U17530 (N_17530,N_14438,N_14611);
xnor U17531 (N_17531,N_15829,N_14014);
nor U17532 (N_17532,N_14447,N_15071);
nor U17533 (N_17533,N_15866,N_15789);
and U17534 (N_17534,N_14820,N_15734);
and U17535 (N_17535,N_15941,N_15462);
xnor U17536 (N_17536,N_14116,N_15173);
and U17537 (N_17537,N_14184,N_15299);
and U17538 (N_17538,N_15726,N_15533);
nand U17539 (N_17539,N_14286,N_14018);
nand U17540 (N_17540,N_15580,N_14602);
nand U17541 (N_17541,N_14530,N_14428);
and U17542 (N_17542,N_15551,N_15047);
xnor U17543 (N_17543,N_15132,N_15568);
and U17544 (N_17544,N_14505,N_14044);
or U17545 (N_17545,N_15802,N_15754);
nor U17546 (N_17546,N_14879,N_14674);
or U17547 (N_17547,N_15448,N_15301);
and U17548 (N_17548,N_15414,N_14607);
xnor U17549 (N_17549,N_14022,N_15205);
nor U17550 (N_17550,N_15354,N_14440);
nor U17551 (N_17551,N_14801,N_15518);
nor U17552 (N_17552,N_14546,N_14364);
xnor U17553 (N_17553,N_14084,N_14856);
nor U17554 (N_17554,N_15902,N_14294);
xor U17555 (N_17555,N_15105,N_14188);
xnor U17556 (N_17556,N_14962,N_15810);
xnor U17557 (N_17557,N_15165,N_15586);
and U17558 (N_17558,N_15699,N_15849);
xor U17559 (N_17559,N_15506,N_15546);
or U17560 (N_17560,N_15266,N_15743);
nand U17561 (N_17561,N_15628,N_14835);
or U17562 (N_17562,N_14294,N_14596);
or U17563 (N_17563,N_14186,N_14683);
nand U17564 (N_17564,N_14965,N_15180);
and U17565 (N_17565,N_15444,N_14252);
and U17566 (N_17566,N_14096,N_15682);
nor U17567 (N_17567,N_14636,N_15557);
xnor U17568 (N_17568,N_15813,N_15775);
nor U17569 (N_17569,N_14730,N_15646);
or U17570 (N_17570,N_14491,N_14025);
and U17571 (N_17571,N_15127,N_15746);
and U17572 (N_17572,N_15195,N_15055);
xor U17573 (N_17573,N_14030,N_14996);
nor U17574 (N_17574,N_14705,N_15336);
nor U17575 (N_17575,N_14002,N_14450);
and U17576 (N_17576,N_14685,N_15004);
nor U17577 (N_17577,N_15981,N_15317);
nand U17578 (N_17578,N_14901,N_14859);
nand U17579 (N_17579,N_14993,N_15162);
and U17580 (N_17580,N_14900,N_14597);
nand U17581 (N_17581,N_15769,N_15290);
nor U17582 (N_17582,N_15774,N_15837);
xor U17583 (N_17583,N_15079,N_14793);
xor U17584 (N_17584,N_14814,N_15352);
xor U17585 (N_17585,N_15413,N_14256);
nand U17586 (N_17586,N_14680,N_15135);
xnor U17587 (N_17587,N_15670,N_14794);
nand U17588 (N_17588,N_15805,N_15311);
and U17589 (N_17589,N_14812,N_14238);
nand U17590 (N_17590,N_14661,N_15969);
and U17591 (N_17591,N_14715,N_15864);
and U17592 (N_17592,N_15216,N_15515);
nand U17593 (N_17593,N_15658,N_14910);
nand U17594 (N_17594,N_14120,N_14189);
and U17595 (N_17595,N_15578,N_14242);
xor U17596 (N_17596,N_15922,N_14827);
xor U17597 (N_17597,N_15272,N_14143);
nand U17598 (N_17598,N_15705,N_14861);
and U17599 (N_17599,N_14590,N_15827);
nand U17600 (N_17600,N_15493,N_14316);
xnor U17601 (N_17601,N_14122,N_15345);
xor U17602 (N_17602,N_15476,N_15423);
nand U17603 (N_17603,N_15039,N_14810);
nand U17604 (N_17604,N_15793,N_14812);
nand U17605 (N_17605,N_15429,N_14349);
and U17606 (N_17606,N_14487,N_14264);
nor U17607 (N_17607,N_14974,N_15034);
or U17608 (N_17608,N_15617,N_14053);
and U17609 (N_17609,N_14053,N_15306);
nand U17610 (N_17610,N_15899,N_14582);
xor U17611 (N_17611,N_14924,N_15946);
xnor U17612 (N_17612,N_15089,N_14302);
nor U17613 (N_17613,N_15483,N_14690);
nor U17614 (N_17614,N_14995,N_14834);
nand U17615 (N_17615,N_15451,N_15732);
xnor U17616 (N_17616,N_14606,N_15546);
nor U17617 (N_17617,N_14063,N_15844);
and U17618 (N_17618,N_15485,N_14800);
or U17619 (N_17619,N_15204,N_15446);
xor U17620 (N_17620,N_15985,N_15808);
nor U17621 (N_17621,N_15353,N_14699);
nor U17622 (N_17622,N_15813,N_14199);
xor U17623 (N_17623,N_14674,N_14084);
nand U17624 (N_17624,N_15696,N_14688);
and U17625 (N_17625,N_15557,N_14170);
nor U17626 (N_17626,N_15012,N_15733);
nor U17627 (N_17627,N_14757,N_15458);
nand U17628 (N_17628,N_15299,N_15208);
and U17629 (N_17629,N_15072,N_15736);
and U17630 (N_17630,N_15203,N_15929);
nor U17631 (N_17631,N_14503,N_15291);
nand U17632 (N_17632,N_15523,N_15500);
and U17633 (N_17633,N_14214,N_15782);
xnor U17634 (N_17634,N_15855,N_14582);
xnor U17635 (N_17635,N_14165,N_15711);
nand U17636 (N_17636,N_14754,N_14088);
nand U17637 (N_17637,N_15062,N_15247);
and U17638 (N_17638,N_14299,N_15924);
and U17639 (N_17639,N_15358,N_15490);
and U17640 (N_17640,N_14759,N_14807);
xnor U17641 (N_17641,N_14744,N_15718);
nand U17642 (N_17642,N_15048,N_15235);
nand U17643 (N_17643,N_15347,N_15965);
and U17644 (N_17644,N_15268,N_14992);
nand U17645 (N_17645,N_14956,N_14881);
and U17646 (N_17646,N_14437,N_15576);
and U17647 (N_17647,N_14308,N_15421);
and U17648 (N_17648,N_14811,N_15618);
or U17649 (N_17649,N_15231,N_14015);
nand U17650 (N_17650,N_15855,N_14458);
nor U17651 (N_17651,N_14039,N_14773);
nor U17652 (N_17652,N_14571,N_15847);
or U17653 (N_17653,N_14719,N_15080);
or U17654 (N_17654,N_15526,N_14324);
and U17655 (N_17655,N_15991,N_15345);
or U17656 (N_17656,N_14101,N_14719);
or U17657 (N_17657,N_14099,N_15247);
nor U17658 (N_17658,N_15798,N_14423);
nor U17659 (N_17659,N_14028,N_14255);
xnor U17660 (N_17660,N_14789,N_15131);
or U17661 (N_17661,N_14391,N_15419);
xor U17662 (N_17662,N_15497,N_14859);
or U17663 (N_17663,N_14536,N_15859);
xnor U17664 (N_17664,N_14746,N_14053);
xor U17665 (N_17665,N_15366,N_15511);
nand U17666 (N_17666,N_15618,N_15093);
nor U17667 (N_17667,N_15016,N_15450);
nand U17668 (N_17668,N_15963,N_15206);
nand U17669 (N_17669,N_15906,N_15867);
or U17670 (N_17670,N_15525,N_14781);
or U17671 (N_17671,N_14208,N_14867);
xnor U17672 (N_17672,N_15472,N_15045);
or U17673 (N_17673,N_15448,N_14121);
xor U17674 (N_17674,N_15635,N_14638);
nor U17675 (N_17675,N_14268,N_14301);
nor U17676 (N_17676,N_15240,N_14743);
nor U17677 (N_17677,N_14577,N_14220);
xnor U17678 (N_17678,N_15668,N_14287);
nand U17679 (N_17679,N_14513,N_14501);
xnor U17680 (N_17680,N_15548,N_15904);
nand U17681 (N_17681,N_15872,N_15023);
xor U17682 (N_17682,N_14976,N_15326);
nor U17683 (N_17683,N_15592,N_15091);
nand U17684 (N_17684,N_14210,N_14700);
nor U17685 (N_17685,N_14881,N_14952);
xor U17686 (N_17686,N_14959,N_15107);
or U17687 (N_17687,N_14614,N_14195);
xor U17688 (N_17688,N_14441,N_15920);
and U17689 (N_17689,N_14076,N_14340);
xor U17690 (N_17690,N_14467,N_15429);
nor U17691 (N_17691,N_14345,N_15597);
xnor U17692 (N_17692,N_15525,N_14898);
xnor U17693 (N_17693,N_15037,N_15686);
and U17694 (N_17694,N_15350,N_15875);
nand U17695 (N_17695,N_14691,N_14467);
and U17696 (N_17696,N_15309,N_15668);
nor U17697 (N_17697,N_14714,N_14013);
nand U17698 (N_17698,N_15733,N_15787);
or U17699 (N_17699,N_14374,N_14001);
or U17700 (N_17700,N_14879,N_15450);
xnor U17701 (N_17701,N_15951,N_15318);
and U17702 (N_17702,N_14755,N_15428);
nand U17703 (N_17703,N_14343,N_15387);
xor U17704 (N_17704,N_15482,N_15236);
nor U17705 (N_17705,N_14180,N_15023);
and U17706 (N_17706,N_14850,N_14880);
nand U17707 (N_17707,N_15243,N_15977);
or U17708 (N_17708,N_14734,N_14193);
or U17709 (N_17709,N_14424,N_14448);
nor U17710 (N_17710,N_15095,N_15377);
nand U17711 (N_17711,N_15314,N_15895);
xor U17712 (N_17712,N_15580,N_14031);
xnor U17713 (N_17713,N_14499,N_15850);
and U17714 (N_17714,N_15756,N_15548);
nand U17715 (N_17715,N_15971,N_14103);
xor U17716 (N_17716,N_15658,N_14745);
nor U17717 (N_17717,N_15287,N_15715);
and U17718 (N_17718,N_14576,N_14411);
nor U17719 (N_17719,N_15448,N_14599);
xor U17720 (N_17720,N_14296,N_14111);
or U17721 (N_17721,N_15466,N_15647);
nand U17722 (N_17722,N_14298,N_15709);
xor U17723 (N_17723,N_15684,N_15465);
nor U17724 (N_17724,N_14020,N_14763);
nand U17725 (N_17725,N_15751,N_14707);
nor U17726 (N_17726,N_15024,N_15958);
nor U17727 (N_17727,N_15619,N_15701);
nand U17728 (N_17728,N_14095,N_15109);
nand U17729 (N_17729,N_15749,N_15928);
xor U17730 (N_17730,N_14969,N_15824);
xnor U17731 (N_17731,N_15642,N_14692);
nand U17732 (N_17732,N_15076,N_14335);
and U17733 (N_17733,N_14520,N_15145);
xnor U17734 (N_17734,N_14555,N_15914);
xnor U17735 (N_17735,N_15582,N_15135);
nor U17736 (N_17736,N_14669,N_15598);
nand U17737 (N_17737,N_15450,N_15146);
or U17738 (N_17738,N_15753,N_15145);
nand U17739 (N_17739,N_14867,N_14224);
nor U17740 (N_17740,N_15846,N_15995);
nand U17741 (N_17741,N_14375,N_14002);
nand U17742 (N_17742,N_15592,N_15550);
and U17743 (N_17743,N_14260,N_15931);
nor U17744 (N_17744,N_14253,N_14245);
nor U17745 (N_17745,N_14255,N_15684);
and U17746 (N_17746,N_14626,N_15084);
and U17747 (N_17747,N_14890,N_14588);
nor U17748 (N_17748,N_15832,N_15393);
nor U17749 (N_17749,N_15452,N_14711);
and U17750 (N_17750,N_14434,N_15926);
xnor U17751 (N_17751,N_14709,N_14441);
and U17752 (N_17752,N_15694,N_14525);
or U17753 (N_17753,N_15128,N_15290);
xnor U17754 (N_17754,N_15819,N_15799);
nor U17755 (N_17755,N_14720,N_15818);
and U17756 (N_17756,N_14276,N_14239);
and U17757 (N_17757,N_14301,N_14514);
and U17758 (N_17758,N_14583,N_15308);
xor U17759 (N_17759,N_15625,N_15332);
and U17760 (N_17760,N_15173,N_14473);
nor U17761 (N_17761,N_14571,N_15937);
or U17762 (N_17762,N_15129,N_15577);
nand U17763 (N_17763,N_15359,N_15825);
or U17764 (N_17764,N_15373,N_14716);
or U17765 (N_17765,N_15457,N_15602);
xor U17766 (N_17766,N_14154,N_15281);
or U17767 (N_17767,N_14700,N_14640);
nor U17768 (N_17768,N_15896,N_15505);
nor U17769 (N_17769,N_15141,N_15014);
or U17770 (N_17770,N_15149,N_15998);
nand U17771 (N_17771,N_14569,N_15618);
nand U17772 (N_17772,N_15767,N_15681);
and U17773 (N_17773,N_15291,N_15616);
and U17774 (N_17774,N_15218,N_14831);
and U17775 (N_17775,N_15503,N_14791);
or U17776 (N_17776,N_14211,N_14579);
and U17777 (N_17777,N_15233,N_15004);
nand U17778 (N_17778,N_15618,N_14332);
nand U17779 (N_17779,N_14575,N_14566);
nor U17780 (N_17780,N_14467,N_14902);
and U17781 (N_17781,N_14887,N_15293);
xnor U17782 (N_17782,N_14329,N_14010);
nor U17783 (N_17783,N_15428,N_14374);
nand U17784 (N_17784,N_15361,N_15814);
nand U17785 (N_17785,N_15259,N_14188);
and U17786 (N_17786,N_14382,N_15055);
nor U17787 (N_17787,N_15515,N_15974);
or U17788 (N_17788,N_15449,N_15002);
or U17789 (N_17789,N_15093,N_15917);
and U17790 (N_17790,N_15802,N_15277);
xnor U17791 (N_17791,N_15275,N_14363);
nand U17792 (N_17792,N_14356,N_15583);
xnor U17793 (N_17793,N_14363,N_15521);
or U17794 (N_17794,N_14904,N_15776);
or U17795 (N_17795,N_15429,N_15126);
nor U17796 (N_17796,N_14544,N_15180);
nand U17797 (N_17797,N_15988,N_14028);
or U17798 (N_17798,N_15736,N_14926);
or U17799 (N_17799,N_15947,N_14900);
nand U17800 (N_17800,N_14106,N_15933);
xnor U17801 (N_17801,N_14229,N_15127);
or U17802 (N_17802,N_14437,N_14669);
and U17803 (N_17803,N_14006,N_15390);
or U17804 (N_17804,N_14674,N_14589);
and U17805 (N_17805,N_15765,N_15799);
or U17806 (N_17806,N_15138,N_15179);
and U17807 (N_17807,N_14939,N_14197);
nor U17808 (N_17808,N_15931,N_14778);
xnor U17809 (N_17809,N_15517,N_15059);
or U17810 (N_17810,N_14521,N_14276);
nor U17811 (N_17811,N_15968,N_14129);
or U17812 (N_17812,N_15275,N_14597);
nand U17813 (N_17813,N_15459,N_14069);
nor U17814 (N_17814,N_15448,N_14968);
and U17815 (N_17815,N_15117,N_14071);
nor U17816 (N_17816,N_15298,N_14735);
or U17817 (N_17817,N_14714,N_15377);
nor U17818 (N_17818,N_15114,N_14393);
nand U17819 (N_17819,N_15844,N_15006);
or U17820 (N_17820,N_15452,N_15843);
or U17821 (N_17821,N_15894,N_15744);
nand U17822 (N_17822,N_15886,N_15818);
and U17823 (N_17823,N_15340,N_14806);
and U17824 (N_17824,N_14651,N_15884);
nor U17825 (N_17825,N_14956,N_15385);
or U17826 (N_17826,N_15094,N_15116);
or U17827 (N_17827,N_15479,N_15892);
nand U17828 (N_17828,N_15580,N_14087);
or U17829 (N_17829,N_15757,N_14930);
or U17830 (N_17830,N_15917,N_14150);
nand U17831 (N_17831,N_15429,N_15227);
and U17832 (N_17832,N_15009,N_15541);
nor U17833 (N_17833,N_14230,N_14837);
xnor U17834 (N_17834,N_15560,N_14840);
or U17835 (N_17835,N_15153,N_14363);
nor U17836 (N_17836,N_15351,N_14575);
or U17837 (N_17837,N_14553,N_15103);
or U17838 (N_17838,N_14528,N_14077);
or U17839 (N_17839,N_15529,N_15722);
xnor U17840 (N_17840,N_14145,N_14092);
or U17841 (N_17841,N_14113,N_14661);
or U17842 (N_17842,N_14204,N_15485);
and U17843 (N_17843,N_14587,N_15470);
and U17844 (N_17844,N_14791,N_14614);
nand U17845 (N_17845,N_15671,N_14341);
and U17846 (N_17846,N_14876,N_15651);
xor U17847 (N_17847,N_15240,N_14742);
nor U17848 (N_17848,N_14162,N_15635);
nand U17849 (N_17849,N_14750,N_15580);
nand U17850 (N_17850,N_14676,N_14925);
xor U17851 (N_17851,N_14479,N_15047);
or U17852 (N_17852,N_14874,N_15271);
nor U17853 (N_17853,N_14427,N_14968);
or U17854 (N_17854,N_15487,N_14635);
xor U17855 (N_17855,N_14496,N_14748);
or U17856 (N_17856,N_14666,N_15405);
nor U17857 (N_17857,N_14096,N_14588);
nor U17858 (N_17858,N_14481,N_14868);
and U17859 (N_17859,N_14079,N_14470);
or U17860 (N_17860,N_14275,N_14469);
nand U17861 (N_17861,N_14663,N_15271);
nor U17862 (N_17862,N_14309,N_15134);
and U17863 (N_17863,N_14929,N_14821);
and U17864 (N_17864,N_14077,N_15050);
and U17865 (N_17865,N_15359,N_15832);
xnor U17866 (N_17866,N_15929,N_15286);
nand U17867 (N_17867,N_14186,N_14115);
nand U17868 (N_17868,N_15904,N_15931);
nand U17869 (N_17869,N_15988,N_14119);
and U17870 (N_17870,N_15741,N_15357);
nand U17871 (N_17871,N_14394,N_14051);
or U17872 (N_17872,N_15443,N_15905);
nand U17873 (N_17873,N_15235,N_15292);
nand U17874 (N_17874,N_14562,N_15321);
xor U17875 (N_17875,N_14514,N_14269);
nor U17876 (N_17876,N_15327,N_14712);
and U17877 (N_17877,N_14064,N_15492);
or U17878 (N_17878,N_14031,N_15814);
nor U17879 (N_17879,N_14293,N_15186);
nor U17880 (N_17880,N_14194,N_14714);
xnor U17881 (N_17881,N_14102,N_15420);
nand U17882 (N_17882,N_15249,N_15127);
xor U17883 (N_17883,N_15057,N_15151);
or U17884 (N_17884,N_14664,N_15156);
or U17885 (N_17885,N_14047,N_14119);
nand U17886 (N_17886,N_15502,N_15983);
and U17887 (N_17887,N_14843,N_15592);
xor U17888 (N_17888,N_14673,N_15747);
nor U17889 (N_17889,N_14052,N_15312);
nor U17890 (N_17890,N_14703,N_15644);
nand U17891 (N_17891,N_14116,N_15216);
nand U17892 (N_17892,N_14367,N_14066);
xnor U17893 (N_17893,N_14770,N_15834);
and U17894 (N_17894,N_15179,N_14554);
nor U17895 (N_17895,N_14286,N_15290);
nand U17896 (N_17896,N_14196,N_14526);
xor U17897 (N_17897,N_15544,N_14123);
xor U17898 (N_17898,N_15955,N_14025);
nand U17899 (N_17899,N_15043,N_15742);
or U17900 (N_17900,N_15129,N_14307);
xor U17901 (N_17901,N_14815,N_14821);
xnor U17902 (N_17902,N_15615,N_15239);
xor U17903 (N_17903,N_14249,N_15071);
xnor U17904 (N_17904,N_14238,N_14358);
or U17905 (N_17905,N_15569,N_15315);
xor U17906 (N_17906,N_14451,N_15447);
nor U17907 (N_17907,N_14058,N_14044);
nand U17908 (N_17908,N_14667,N_15673);
or U17909 (N_17909,N_15829,N_15542);
xor U17910 (N_17910,N_14294,N_15410);
and U17911 (N_17911,N_15341,N_15635);
nor U17912 (N_17912,N_14629,N_15573);
nand U17913 (N_17913,N_14489,N_14557);
nor U17914 (N_17914,N_14000,N_14861);
and U17915 (N_17915,N_14327,N_14452);
nor U17916 (N_17916,N_14221,N_15254);
and U17917 (N_17917,N_15565,N_15077);
or U17918 (N_17918,N_14606,N_14472);
or U17919 (N_17919,N_14644,N_15823);
nor U17920 (N_17920,N_14382,N_14642);
and U17921 (N_17921,N_15899,N_14385);
or U17922 (N_17922,N_15274,N_15606);
nor U17923 (N_17923,N_14340,N_14040);
or U17924 (N_17924,N_14182,N_14120);
nand U17925 (N_17925,N_14479,N_14590);
xor U17926 (N_17926,N_14458,N_15426);
and U17927 (N_17927,N_14311,N_15623);
xor U17928 (N_17928,N_15755,N_15420);
or U17929 (N_17929,N_14633,N_14549);
and U17930 (N_17930,N_15008,N_14395);
nor U17931 (N_17931,N_15600,N_15252);
nand U17932 (N_17932,N_15016,N_14373);
xor U17933 (N_17933,N_15844,N_14097);
and U17934 (N_17934,N_15397,N_15353);
and U17935 (N_17935,N_15888,N_14732);
or U17936 (N_17936,N_14556,N_14600);
or U17937 (N_17937,N_15204,N_14018);
nand U17938 (N_17938,N_15896,N_14907);
xor U17939 (N_17939,N_15044,N_15938);
nand U17940 (N_17940,N_14384,N_14143);
and U17941 (N_17941,N_14542,N_14560);
and U17942 (N_17942,N_15498,N_14542);
and U17943 (N_17943,N_14760,N_14665);
nand U17944 (N_17944,N_14948,N_15212);
nand U17945 (N_17945,N_14209,N_14563);
xnor U17946 (N_17946,N_14006,N_15903);
nand U17947 (N_17947,N_15445,N_14015);
nand U17948 (N_17948,N_14880,N_15142);
and U17949 (N_17949,N_14506,N_15815);
and U17950 (N_17950,N_15139,N_15507);
nand U17951 (N_17951,N_15260,N_14331);
or U17952 (N_17952,N_15678,N_15426);
xnor U17953 (N_17953,N_14160,N_14933);
nor U17954 (N_17954,N_14054,N_14255);
nor U17955 (N_17955,N_14757,N_15730);
xor U17956 (N_17956,N_15814,N_14048);
nand U17957 (N_17957,N_15154,N_14585);
and U17958 (N_17958,N_14069,N_14053);
or U17959 (N_17959,N_14996,N_15155);
and U17960 (N_17960,N_14401,N_14616);
xnor U17961 (N_17961,N_15463,N_14460);
nand U17962 (N_17962,N_14949,N_14839);
or U17963 (N_17963,N_14908,N_14345);
and U17964 (N_17964,N_15868,N_15650);
or U17965 (N_17965,N_15420,N_15535);
xnor U17966 (N_17966,N_14017,N_15226);
or U17967 (N_17967,N_15223,N_14066);
or U17968 (N_17968,N_15247,N_15404);
nor U17969 (N_17969,N_15352,N_15902);
xnor U17970 (N_17970,N_14897,N_15280);
and U17971 (N_17971,N_15677,N_15370);
xnor U17972 (N_17972,N_15964,N_15015);
xnor U17973 (N_17973,N_15711,N_14084);
or U17974 (N_17974,N_15837,N_15548);
xnor U17975 (N_17975,N_15082,N_15947);
nor U17976 (N_17976,N_14903,N_15134);
xnor U17977 (N_17977,N_15850,N_15480);
nand U17978 (N_17978,N_15211,N_14638);
or U17979 (N_17979,N_15229,N_15213);
or U17980 (N_17980,N_14454,N_14527);
or U17981 (N_17981,N_15520,N_14389);
xor U17982 (N_17982,N_15354,N_14933);
xor U17983 (N_17983,N_14785,N_14310);
or U17984 (N_17984,N_14880,N_15988);
xnor U17985 (N_17985,N_15846,N_15947);
xor U17986 (N_17986,N_15906,N_15771);
or U17987 (N_17987,N_15250,N_15807);
and U17988 (N_17988,N_14792,N_14948);
nor U17989 (N_17989,N_15852,N_14739);
xor U17990 (N_17990,N_15628,N_14599);
nor U17991 (N_17991,N_14214,N_15536);
nor U17992 (N_17992,N_14851,N_14721);
nor U17993 (N_17993,N_14355,N_14754);
nand U17994 (N_17994,N_14664,N_15394);
nand U17995 (N_17995,N_15117,N_15977);
nand U17996 (N_17996,N_15801,N_15842);
nand U17997 (N_17997,N_14512,N_14275);
and U17998 (N_17998,N_15724,N_15552);
xnor U17999 (N_17999,N_15760,N_15923);
nand U18000 (N_18000,N_16268,N_16229);
xnor U18001 (N_18001,N_17226,N_17662);
and U18002 (N_18002,N_17134,N_17568);
or U18003 (N_18003,N_16176,N_17592);
nand U18004 (N_18004,N_16575,N_17557);
xnor U18005 (N_18005,N_16494,N_17511);
or U18006 (N_18006,N_17092,N_16251);
and U18007 (N_18007,N_17259,N_17274);
nand U18008 (N_18008,N_17993,N_17110);
nand U18009 (N_18009,N_17117,N_17795);
nor U18010 (N_18010,N_17326,N_16996);
nor U18011 (N_18011,N_16782,N_16682);
nand U18012 (N_18012,N_16164,N_17058);
xor U18013 (N_18013,N_17497,N_16359);
nor U18014 (N_18014,N_16777,N_16814);
nand U18015 (N_18015,N_17124,N_17199);
nand U18016 (N_18016,N_17344,N_16526);
nor U18017 (N_18017,N_17096,N_17059);
nand U18018 (N_18018,N_16562,N_17031);
and U18019 (N_18019,N_17131,N_17216);
nor U18020 (N_18020,N_16568,N_16248);
and U18021 (N_18021,N_17069,N_16276);
nor U18022 (N_18022,N_17706,N_16025);
nand U18023 (N_18023,N_17841,N_16637);
or U18024 (N_18024,N_16375,N_17189);
xor U18025 (N_18025,N_17112,N_17487);
or U18026 (N_18026,N_17918,N_16872);
nor U18027 (N_18027,N_16324,N_16305);
nor U18028 (N_18028,N_17994,N_17252);
or U18029 (N_18029,N_16976,N_16593);
and U18030 (N_18030,N_17267,N_16982);
or U18031 (N_18031,N_17379,N_16937);
and U18032 (N_18032,N_16977,N_16502);
nor U18033 (N_18033,N_17996,N_17543);
nand U18034 (N_18034,N_17647,N_17775);
nor U18035 (N_18035,N_16288,N_16916);
or U18036 (N_18036,N_16220,N_16764);
nor U18037 (N_18037,N_16130,N_17399);
or U18038 (N_18038,N_16205,N_16731);
or U18039 (N_18039,N_16888,N_16363);
or U18040 (N_18040,N_17997,N_17292);
and U18041 (N_18041,N_17300,N_17439);
and U18042 (N_18042,N_16497,N_16675);
and U18043 (N_18043,N_17355,N_17605);
nor U18044 (N_18044,N_17505,N_17298);
nor U18045 (N_18045,N_16067,N_16341);
and U18046 (N_18046,N_17322,N_17545);
nand U18047 (N_18047,N_16501,N_17416);
and U18048 (N_18048,N_16558,N_16713);
nand U18049 (N_18049,N_16667,N_17974);
and U18050 (N_18050,N_16813,N_17411);
nor U18051 (N_18051,N_16401,N_17196);
and U18052 (N_18052,N_16153,N_16127);
nand U18053 (N_18053,N_16880,N_17296);
or U18054 (N_18054,N_16831,N_16170);
nand U18055 (N_18055,N_17752,N_17661);
nand U18056 (N_18056,N_17220,N_16296);
xnor U18057 (N_18057,N_16907,N_16047);
nor U18058 (N_18058,N_17025,N_16257);
nor U18059 (N_18059,N_17162,N_16676);
nand U18060 (N_18060,N_17395,N_17089);
or U18061 (N_18061,N_17366,N_17209);
or U18062 (N_18062,N_17085,N_17716);
nor U18063 (N_18063,N_16274,N_16587);
and U18064 (N_18064,N_16459,N_16409);
nand U18065 (N_18065,N_16998,N_17167);
or U18066 (N_18066,N_17781,N_16427);
nand U18067 (N_18067,N_17554,N_17075);
xnor U18068 (N_18068,N_17718,N_16661);
nand U18069 (N_18069,N_16510,N_16147);
or U18070 (N_18070,N_17707,N_17520);
and U18071 (N_18071,N_17897,N_17123);
nor U18072 (N_18072,N_17797,N_17137);
or U18073 (N_18073,N_16590,N_17359);
xor U18074 (N_18074,N_17287,N_16235);
nand U18075 (N_18075,N_16895,N_17597);
nand U18076 (N_18076,N_17817,N_17023);
xor U18077 (N_18077,N_17810,N_16543);
nor U18078 (N_18078,N_17796,N_17792);
xnor U18079 (N_18079,N_17933,N_17643);
nor U18080 (N_18080,N_17135,N_16602);
nand U18081 (N_18081,N_16043,N_16358);
and U18082 (N_18082,N_16546,N_16356);
or U18083 (N_18083,N_17780,N_17442);
nand U18084 (N_18084,N_17051,N_17422);
xnor U18085 (N_18085,N_17800,N_17742);
or U18086 (N_18086,N_16418,N_16760);
nand U18087 (N_18087,N_16853,N_17281);
and U18088 (N_18088,N_17712,N_16965);
xnor U18089 (N_18089,N_16385,N_16962);
nand U18090 (N_18090,N_17246,N_16095);
or U18091 (N_18091,N_17308,N_16351);
nand U18092 (N_18092,N_17822,N_17163);
nor U18093 (N_18093,N_17930,N_17338);
or U18094 (N_18094,N_16617,N_16722);
nor U18095 (N_18095,N_17481,N_17409);
and U18096 (N_18096,N_16697,N_16640);
and U18097 (N_18097,N_16978,N_16460);
nand U18098 (N_18098,N_16495,N_17140);
xnor U18099 (N_18099,N_17127,N_17490);
nand U18100 (N_18100,N_16215,N_16330);
nand U18101 (N_18101,N_16834,N_16589);
nand U18102 (N_18102,N_16733,N_16098);
or U18103 (N_18103,N_16243,N_17523);
xor U18104 (N_18104,N_17604,N_17036);
and U18105 (N_18105,N_16429,N_17510);
and U18106 (N_18106,N_16333,N_17938);
and U18107 (N_18107,N_17939,N_16538);
and U18108 (N_18108,N_16088,N_17719);
xor U18109 (N_18109,N_16044,N_17835);
nand U18110 (N_18110,N_17202,N_16979);
and U18111 (N_18111,N_16340,N_17552);
or U18112 (N_18112,N_16491,N_17669);
and U18113 (N_18113,N_17048,N_16129);
xnor U18114 (N_18114,N_17968,N_17887);
xor U18115 (N_18115,N_17736,N_17384);
nor U18116 (N_18116,N_17114,N_17213);
nand U18117 (N_18117,N_17369,N_17599);
nor U18118 (N_18118,N_16817,N_17690);
and U18119 (N_18119,N_17757,N_16860);
nand U18120 (N_18120,N_16124,N_16918);
nand U18121 (N_18121,N_17266,N_16975);
xor U18122 (N_18122,N_17747,N_17517);
and U18123 (N_18123,N_17172,N_17697);
or U18124 (N_18124,N_16809,N_16306);
xnor U18125 (N_18125,N_17845,N_16138);
nor U18126 (N_18126,N_16011,N_17854);
or U18127 (N_18127,N_16107,N_17181);
and U18128 (N_18128,N_16023,N_17040);
nand U18129 (N_18129,N_16457,N_17896);
or U18130 (N_18130,N_17519,N_17150);
xor U18131 (N_18131,N_17404,N_17726);
and U18132 (N_18132,N_17803,N_17417);
and U18133 (N_18133,N_16493,N_16755);
nor U18134 (N_18134,N_16055,N_17415);
or U18135 (N_18135,N_17190,N_16840);
nand U18136 (N_18136,N_17595,N_17231);
xor U18137 (N_18137,N_16065,N_17122);
xor U18138 (N_18138,N_16111,N_16580);
or U18139 (N_18139,N_16818,N_17437);
and U18140 (N_18140,N_17013,N_16717);
and U18141 (N_18141,N_17157,N_17488);
and U18142 (N_18142,N_16400,N_17495);
xnor U18143 (N_18143,N_16522,N_17971);
or U18144 (N_18144,N_16553,N_16901);
nand U18145 (N_18145,N_16197,N_17895);
nor U18146 (N_18146,N_17879,N_16606);
nand U18147 (N_18147,N_16613,N_17323);
nand U18148 (N_18148,N_16284,N_16527);
xnor U18149 (N_18149,N_16792,N_17876);
nor U18150 (N_18150,N_17492,N_16779);
and U18151 (N_18151,N_16654,N_17087);
or U18152 (N_18152,N_17650,N_16623);
and U18153 (N_18153,N_17911,N_16455);
nor U18154 (N_18154,N_16225,N_17363);
xnor U18155 (N_18155,N_16174,N_17353);
nand U18156 (N_18156,N_16287,N_17079);
xnor U18157 (N_18157,N_17826,N_16796);
nor U18158 (N_18158,N_17158,N_17965);
or U18159 (N_18159,N_17329,N_17567);
and U18160 (N_18160,N_16403,N_17857);
xnor U18161 (N_18161,N_17589,N_17341);
nand U18162 (N_18162,N_17708,N_16956);
or U18163 (N_18163,N_17192,N_17548);
nand U18164 (N_18164,N_17086,N_16433);
nor U18165 (N_18165,N_17531,N_16766);
or U18166 (N_18166,N_17864,N_16985);
xnor U18167 (N_18167,N_17247,N_17861);
or U18168 (N_18168,N_17152,N_17514);
or U18169 (N_18169,N_16845,N_16847);
xnor U18170 (N_18170,N_17999,N_16443);
and U18171 (N_18171,N_16159,N_17104);
nor U18172 (N_18172,N_17116,N_16173);
and U18173 (N_18173,N_17204,N_17614);
or U18174 (N_18174,N_17633,N_17739);
xor U18175 (N_18175,N_17253,N_17642);
nor U18176 (N_18176,N_17465,N_17277);
nor U18177 (N_18177,N_17952,N_17340);
nand U18178 (N_18178,N_17691,N_17333);
xor U18179 (N_18179,N_17766,N_16968);
xnor U18180 (N_18180,N_17834,N_17769);
xor U18181 (N_18181,N_16581,N_17536);
nand U18182 (N_18182,N_17912,N_16031);
or U18183 (N_18183,N_16304,N_16677);
nand U18184 (N_18184,N_16783,N_17419);
or U18185 (N_18185,N_17011,N_17449);
or U18186 (N_18186,N_16320,N_16277);
and U18187 (N_18187,N_17045,N_17676);
and U18188 (N_18188,N_16269,N_17774);
or U18189 (N_18189,N_16635,N_16994);
nand U18190 (N_18190,N_17414,N_17821);
nand U18191 (N_18191,N_17327,N_16134);
nand U18192 (N_18192,N_16877,N_16332);
xnor U18193 (N_18193,N_16083,N_16253);
or U18194 (N_18194,N_17244,N_17223);
and U18195 (N_18195,N_17161,N_17951);
and U18196 (N_18196,N_17348,N_16074);
nand U18197 (N_18197,N_17154,N_16687);
xnor U18198 (N_18198,N_16050,N_17831);
and U18199 (N_18199,N_17090,N_17892);
xnor U18200 (N_18200,N_16788,N_17148);
xnor U18201 (N_18201,N_16533,N_17015);
xor U18202 (N_18202,N_17584,N_16549);
and U18203 (N_18203,N_17856,N_16832);
nand U18204 (N_18204,N_16614,N_16308);
nand U18205 (N_18205,N_16850,N_16370);
and U18206 (N_18206,N_17107,N_17645);
nand U18207 (N_18207,N_16540,N_16481);
or U18208 (N_18208,N_16371,N_16941);
xnor U18209 (N_18209,N_16078,N_16206);
nand U18210 (N_18210,N_17397,N_17637);
nor U18211 (N_18211,N_17236,N_16283);
nor U18212 (N_18212,N_16193,N_17881);
or U18213 (N_18213,N_17789,N_17755);
or U18214 (N_18214,N_16041,N_16202);
xnor U18215 (N_18215,N_16136,N_17607);
nor U18216 (N_18216,N_16106,N_17073);
nor U18217 (N_18217,N_17016,N_17233);
xor U18218 (N_18218,N_16952,N_17351);
or U18219 (N_18219,N_17566,N_17037);
nand U18220 (N_18220,N_17787,N_16437);
xnor U18221 (N_18221,N_17908,N_16072);
xnor U18222 (N_18222,N_17171,N_16891);
nor U18223 (N_18223,N_16146,N_17130);
and U18224 (N_18224,N_16003,N_16987);
or U18225 (N_18225,N_16112,N_16149);
nor U18226 (N_18226,N_16607,N_17812);
and U18227 (N_18227,N_17020,N_17120);
nand U18228 (N_18228,N_16660,N_16275);
nand U18229 (N_18229,N_17648,N_17230);
nor U18230 (N_18230,N_17046,N_17318);
xor U18231 (N_18231,N_17940,N_16959);
xnor U18232 (N_18232,N_17931,N_17248);
xor U18233 (N_18233,N_16309,N_17883);
or U18234 (N_18234,N_16312,N_17047);
nor U18235 (N_18235,N_16123,N_16439);
or U18236 (N_18236,N_17555,N_16113);
or U18237 (N_18237,N_17227,N_17990);
nand U18238 (N_18238,N_17860,N_16335);
and U18239 (N_18239,N_16420,N_17392);
nor U18240 (N_18240,N_17724,N_16042);
and U18241 (N_18241,N_17334,N_16221);
xor U18242 (N_18242,N_17663,N_17866);
and U18243 (N_18243,N_16970,N_17467);
or U18244 (N_18244,N_17560,N_16051);
nand U18245 (N_18245,N_17989,N_17108);
nand U18246 (N_18246,N_17054,N_17504);
and U18247 (N_18247,N_17738,N_17958);
or U18248 (N_18248,N_16539,N_17242);
and U18249 (N_18249,N_16523,N_17986);
nor U18250 (N_18250,N_16644,N_16828);
xnor U18251 (N_18251,N_17722,N_16585);
and U18252 (N_18252,N_17286,N_17578);
nand U18253 (N_18253,N_16512,N_16757);
or U18254 (N_18254,N_16869,N_17547);
nor U18255 (N_18255,N_17237,N_16761);
xor U18256 (N_18256,N_16339,N_17283);
and U18257 (N_18257,N_16360,N_17955);
nand U18258 (N_18258,N_17677,N_17193);
or U18259 (N_18259,N_16210,N_16913);
or U18260 (N_18260,N_16505,N_16228);
and U18261 (N_18261,N_17966,N_16171);
nor U18262 (N_18262,N_16574,N_16695);
xor U18263 (N_18263,N_17256,N_17598);
nand U18264 (N_18264,N_16983,N_17390);
nand U18265 (N_18265,N_17763,N_17546);
xnor U18266 (N_18266,N_17961,N_16663);
nor U18267 (N_18267,N_16314,N_17301);
xnor U18268 (N_18268,N_16762,N_17003);
or U18269 (N_18269,N_16372,N_16318);
and U18270 (N_18270,N_17423,N_16326);
and U18271 (N_18271,N_16839,N_16488);
or U18272 (N_18272,N_16423,N_17463);
nand U18273 (N_18273,N_16485,N_17184);
xnor U18274 (N_18274,N_16621,N_16099);
nor U18275 (N_18275,N_16086,N_17109);
and U18276 (N_18276,N_16062,N_17418);
nor U18277 (N_18277,N_17033,N_17493);
nor U18278 (N_18278,N_16133,N_16870);
xor U18279 (N_18279,N_16925,N_17024);
xor U18280 (N_18280,N_17466,N_17197);
xor U18281 (N_18281,N_16852,N_16658);
nor U18282 (N_18282,N_17455,N_17391);
xor U18283 (N_18283,N_17410,N_16411);
xor U18284 (N_18284,N_17225,N_17634);
xnor U18285 (N_18285,N_16754,N_16462);
nand U18286 (N_18286,N_16195,N_17027);
xnor U18287 (N_18287,N_17980,N_17977);
xor U18288 (N_18288,N_17367,N_17014);
nand U18289 (N_18289,N_16059,N_17711);
nor U18290 (N_18290,N_16725,N_16236);
or U18291 (N_18291,N_17689,N_16529);
or U18292 (N_18292,N_17710,N_16417);
xor U18293 (N_18293,N_17907,N_17970);
and U18294 (N_18294,N_17867,N_17473);
nand U18295 (N_18295,N_16378,N_17177);
xnor U18296 (N_18296,N_17731,N_17535);
xnor U18297 (N_18297,N_17594,N_17332);
nand U18298 (N_18298,N_16851,N_16247);
and U18299 (N_18299,N_16807,N_17666);
xnor U18300 (N_18300,N_17464,N_17540);
or U18301 (N_18301,N_16947,N_17639);
and U18302 (N_18302,N_16576,N_17936);
or U18303 (N_18303,N_17573,N_16863);
xor U18304 (N_18304,N_16154,N_17901);
or U18305 (N_18305,N_17146,N_16520);
nand U18306 (N_18306,N_17099,N_17412);
nand U18307 (N_18307,N_16069,N_16477);
or U18308 (N_18308,N_17638,N_17849);
xnor U18309 (N_18309,N_17571,N_17026);
or U18310 (N_18310,N_16264,N_16957);
xor U18311 (N_18311,N_17581,N_16855);
xor U18312 (N_18312,N_17593,N_16728);
nand U18313 (N_18313,N_16185,N_16014);
or U18314 (N_18314,N_16995,N_17331);
and U18315 (N_18315,N_17434,N_17963);
nor U18316 (N_18316,N_17692,N_17919);
nand U18317 (N_18317,N_16953,N_17457);
nand U18318 (N_18318,N_17635,N_17139);
xor U18319 (N_18319,N_17920,N_16989);
nand U18320 (N_18320,N_16873,N_16303);
xor U18321 (N_18321,N_16945,N_16186);
xor U18322 (N_18322,N_16273,N_16026);
and U18323 (N_18323,N_16604,N_17756);
nand U18324 (N_18324,N_16161,N_17610);
nand U18325 (N_18325,N_16896,N_16190);
nor U18326 (N_18326,N_17444,N_17836);
nor U18327 (N_18327,N_17541,N_16861);
nor U18328 (N_18328,N_17922,N_16142);
nor U18329 (N_18329,N_16293,N_16883);
xnor U18330 (N_18330,N_17299,N_16507);
nor U18331 (N_18331,N_16745,N_17673);
nor U18332 (N_18332,N_17705,N_17767);
and U18333 (N_18333,N_16969,N_16037);
and U18334 (N_18334,N_16601,N_17556);
and U18335 (N_18335,N_16890,N_16163);
and U18336 (N_18336,N_17316,N_16569);
or U18337 (N_18337,N_16374,N_16742);
and U18338 (N_18338,N_16948,N_17325);
nand U18339 (N_18339,N_16775,N_17288);
or U18340 (N_18340,N_16710,N_16881);
and U18341 (N_18341,N_17622,N_16929);
nand U18342 (N_18342,N_17262,N_17585);
xor U18343 (N_18343,N_17270,N_16216);
or U18344 (N_18344,N_17979,N_16912);
or U18345 (N_18345,N_17273,N_16282);
nor U18346 (N_18346,N_17337,N_16906);
nand U18347 (N_18347,N_17884,N_17586);
xor U18348 (N_18348,N_17371,N_17704);
xnor U18349 (N_18349,N_16350,N_16213);
nand U18350 (N_18350,N_17271,N_16781);
nand U18351 (N_18351,N_16352,N_17018);
and U18352 (N_18352,N_17583,N_16398);
nand U18353 (N_18353,N_17491,N_17660);
nor U18354 (N_18354,N_16033,N_16651);
nor U18355 (N_18355,N_16992,N_17007);
or U18356 (N_18356,N_16625,N_17533);
or U18357 (N_18357,N_17043,N_17229);
xor U18358 (N_18358,N_16620,N_16795);
nor U18359 (N_18359,N_17790,N_16563);
xor U18360 (N_18360,N_17451,N_17132);
and U18361 (N_18361,N_16232,N_16366);
xor U18362 (N_18362,N_16917,N_17839);
nand U18363 (N_18363,N_17064,N_17732);
or U18364 (N_18364,N_16577,N_16121);
nand U18365 (N_18365,N_17649,N_17214);
xor U18366 (N_18366,N_17913,N_17681);
and U18367 (N_18367,N_16899,N_17203);
or U18368 (N_18368,N_16081,N_17400);
and U18369 (N_18369,N_17658,N_17032);
nor U18370 (N_18370,N_17667,N_17498);
or U18371 (N_18371,N_16431,N_17886);
nand U18372 (N_18372,N_17241,N_17057);
and U18373 (N_18373,N_16271,N_17373);
or U18374 (N_18374,N_17254,N_17474);
or U18375 (N_18375,N_16555,N_16810);
xnor U18376 (N_18376,N_16445,N_16097);
and U18377 (N_18377,N_17728,N_17848);
nand U18378 (N_18378,N_17055,N_16862);
xnor U18379 (N_18379,N_16468,N_16804);
xnor U18380 (N_18380,N_16703,N_17580);
or U18381 (N_18381,N_17311,N_17456);
nand U18382 (N_18382,N_17034,N_17264);
or U18383 (N_18383,N_17715,N_16610);
nor U18384 (N_18384,N_16674,N_17169);
nand U18385 (N_18385,N_17759,N_16940);
nand U18386 (N_18386,N_17078,N_17928);
and U18387 (N_18387,N_17530,N_16944);
or U18388 (N_18388,N_17102,N_16647);
xnor U18389 (N_18389,N_16004,N_16842);
xnor U18390 (N_18390,N_16950,N_17569);
and U18391 (N_18391,N_17394,N_16642);
xnor U18392 (N_18392,N_16826,N_17601);
nand U18393 (N_18393,N_16038,N_17820);
nand U18394 (N_18394,N_17342,N_17129);
nand U18395 (N_18395,N_16207,N_17364);
or U18396 (N_18396,N_16833,N_17080);
xor U18397 (N_18397,N_16552,N_17462);
or U18398 (N_18398,N_16560,N_16369);
xnor U18399 (N_18399,N_16278,N_17703);
xor U18400 (N_18400,N_17263,N_16249);
and U18401 (N_18401,N_17851,N_16368);
and U18402 (N_18402,N_17119,N_17582);
nand U18403 (N_18403,N_17729,N_17954);
and U18404 (N_18404,N_17050,N_17611);
or U18405 (N_18405,N_17022,N_16737);
or U18406 (N_18406,N_16573,N_16955);
and U18407 (N_18407,N_16325,N_16611);
nand U18408 (N_18408,N_17304,N_17091);
xnor U18409 (N_18409,N_16683,N_17179);
xor U18410 (N_18410,N_17923,N_17762);
nand U18411 (N_18411,N_17613,N_17501);
and U18412 (N_18412,N_16448,N_17577);
and U18413 (N_18413,N_16222,N_17380);
and U18414 (N_18414,N_17088,N_16645);
and U18415 (N_18415,N_17255,N_17430);
and U18416 (N_18416,N_17061,N_16518);
xor U18417 (N_18417,N_16165,N_16467);
and U18418 (N_18418,N_17679,N_16492);
and U18419 (N_18419,N_16414,N_17950);
or U18420 (N_18420,N_17828,N_17000);
nand U18421 (N_18421,N_17624,N_17383);
xor U18422 (N_18422,N_17093,N_17943);
xor U18423 (N_18423,N_17272,N_16157);
xnor U18424 (N_18424,N_16797,N_17865);
nand U18425 (N_18425,N_17753,N_17824);
and U18426 (N_18426,N_16662,N_16071);
or U18427 (N_18427,N_16046,N_17195);
nand U18428 (N_18428,N_16101,N_16691);
nand U18429 (N_18429,N_17903,N_17071);
and U18430 (N_18430,N_16730,N_17785);
nand U18431 (N_18431,N_16672,N_17238);
xor U18432 (N_18432,N_17778,N_16786);
or U18433 (N_18433,N_16724,N_16297);
nor U18434 (N_18434,N_16049,N_16572);
xnor U18435 (N_18435,N_17309,N_17698);
or U18436 (N_18436,N_17591,N_16187);
and U18437 (N_18437,N_16648,N_16075);
or U18438 (N_18438,N_16039,N_17160);
and U18439 (N_18439,N_17587,N_16551);
nor U18440 (N_18440,N_16933,N_17748);
or U18441 (N_18441,N_16889,N_16922);
nand U18442 (N_18442,N_17563,N_17471);
xor U18443 (N_18443,N_17542,N_16416);
xor U18444 (N_18444,N_17653,N_17798);
and U18445 (N_18445,N_17068,N_16438);
nand U18446 (N_18446,N_17837,N_16032);
and U18447 (N_18447,N_16451,N_16544);
or U18448 (N_18448,N_16487,N_17072);
nor U18449 (N_18449,N_17362,N_16397);
and U18450 (N_18450,N_16511,N_16270);
nor U18451 (N_18451,N_17562,N_16260);
and U18452 (N_18452,N_17111,N_16698);
and U18453 (N_18453,N_16652,N_17709);
nor U18454 (N_18454,N_17403,N_17927);
xor U18455 (N_18455,N_16857,N_17118);
or U18456 (N_18456,N_17935,N_16226);
xnor U18457 (N_18457,N_16189,N_17084);
or U18458 (N_18458,N_17891,N_16636);
nor U18459 (N_18459,N_16156,N_17217);
and U18460 (N_18460,N_16272,N_16615);
or U18461 (N_18461,N_16364,N_17807);
and U18462 (N_18462,N_16354,N_17670);
and U18463 (N_18463,N_17945,N_17066);
and U18464 (N_18464,N_17870,N_16772);
nand U18465 (N_18465,N_17811,N_16599);
and U18466 (N_18466,N_16456,N_16704);
nand U18467 (N_18467,N_16020,N_17953);
nor U18468 (N_18468,N_16391,N_17576);
or U18469 (N_18469,N_16096,N_16155);
xnor U18470 (N_18470,N_16432,N_16699);
nand U18471 (N_18471,N_16999,N_17387);
or U18472 (N_18472,N_17210,N_17324);
or U18473 (N_18473,N_16089,N_17564);
nand U18474 (N_18474,N_17446,N_16738);
and U18475 (N_18475,N_16013,N_17279);
xor U18476 (N_18476,N_16634,N_16478);
xor U18477 (N_18477,N_17001,N_16864);
xor U18478 (N_18478,N_16087,N_17310);
or U18479 (N_18479,N_17948,N_17675);
nor U18480 (N_18480,N_17644,N_16515);
and U18481 (N_18481,N_16915,N_17745);
nor U18482 (N_18482,N_16879,N_17374);
and U18483 (N_18483,N_16167,N_17532);
nor U18484 (N_18484,N_16148,N_16465);
and U18485 (N_18485,N_17855,N_16294);
or U18486 (N_18486,N_16082,N_16405);
nand U18487 (N_18487,N_16811,N_17981);
or U18488 (N_18488,N_16627,N_16981);
nand U18489 (N_18489,N_16390,N_17469);
or U18490 (N_18490,N_17646,N_17559);
xor U18491 (N_18491,N_16085,N_17074);
nand U18492 (N_18492,N_16219,N_16958);
or U18493 (N_18493,N_16489,N_17094);
nand U18494 (N_18494,N_16441,N_16412);
xor U18495 (N_18495,N_16291,N_17813);
and U18496 (N_18496,N_17029,N_17313);
or U18497 (N_18497,N_16504,N_17773);
nand U18498 (N_18498,N_17873,N_16212);
and U18499 (N_18499,N_16169,N_16218);
or U18500 (N_18500,N_16770,N_17499);
and U18501 (N_18501,N_16854,N_17992);
or U18502 (N_18502,N_16482,N_16723);
or U18503 (N_18503,N_16750,N_17044);
nor U18504 (N_18504,N_17809,N_17890);
xor U18505 (N_18505,N_17700,N_17529);
nand U18506 (N_18506,N_16310,N_17983);
or U18507 (N_18507,N_17882,N_16752);
xnor U18508 (N_18508,N_17378,N_16116);
nand U18509 (N_18509,N_16000,N_17844);
nor U18510 (N_18510,N_17436,N_17544);
and U18511 (N_18511,N_16240,N_17852);
or U18512 (N_18512,N_16559,N_17282);
or U18513 (N_18513,N_16259,N_17405);
and U18514 (N_18514,N_17121,N_17915);
nor U18515 (N_18515,N_16759,N_17278);
and U18516 (N_18516,N_17347,N_17625);
nor U18517 (N_18517,N_16125,N_16882);
nor U18518 (N_18518,N_16670,N_17232);
nand U18519 (N_18519,N_16858,N_17425);
xor U18520 (N_18520,N_17062,N_17136);
and U18521 (N_18521,N_17534,N_17804);
xnor U18522 (N_18522,N_16486,N_17850);
xnor U18523 (N_18523,N_17429,N_16805);
xnor U18524 (N_18524,N_17749,N_17388);
nand U18525 (N_18525,N_17426,N_17106);
xnor U18526 (N_18526,N_16110,N_17524);
or U18527 (N_18527,N_16784,N_17115);
nand U18528 (N_18528,N_16517,N_16141);
nand U18529 (N_18529,N_16910,N_17816);
or U18530 (N_18530,N_16380,N_17777);
xor U18531 (N_18531,N_17618,N_17240);
xnor U18532 (N_18532,N_16384,N_16619);
nand U18533 (N_18533,N_17275,N_16094);
xor U18534 (N_18534,N_16974,N_17261);
or U18535 (N_18535,N_16932,N_16452);
or U18536 (N_18536,N_17432,N_17623);
or U18537 (N_18537,N_17668,N_16612);
and U18538 (N_18538,N_17407,N_17761);
or U18539 (N_18539,N_17343,N_17486);
xnor U18540 (N_18540,N_16624,N_16566);
nand U18541 (N_18541,N_17537,N_16347);
xor U18542 (N_18542,N_17791,N_17636);
nand U18543 (N_18543,N_17260,N_17503);
nor U18544 (N_18544,N_16104,N_17889);
nand U18545 (N_18545,N_17454,N_16689);
xnor U18546 (N_18546,N_16630,N_16570);
and U18547 (N_18547,N_17829,N_16597);
nor U18548 (N_18548,N_17632,N_16245);
xor U18549 (N_18549,N_17833,N_16886);
nor U18550 (N_18550,N_17615,N_17725);
nand U18551 (N_18551,N_17733,N_16241);
or U18552 (N_18552,N_16990,N_17336);
nand U18553 (N_18553,N_16255,N_16824);
or U18554 (N_18554,N_16399,N_17946);
nor U18555 (N_18555,N_16541,N_16827);
xnor U18556 (N_18556,N_16177,N_16716);
nor U18557 (N_18557,N_16935,N_17863);
nor U18558 (N_18558,N_17627,N_16066);
and U18559 (N_18559,N_17458,N_17616);
nor U18560 (N_18560,N_17349,N_16694);
or U18561 (N_18561,N_16763,N_16030);
or U18562 (N_18562,N_17783,N_17460);
nor U18563 (N_18563,N_16388,N_16639);
nand U18564 (N_18564,N_17480,N_16466);
or U18565 (N_18565,N_16231,N_17421);
and U18566 (N_18566,N_16556,N_17941);
xnor U18567 (N_18567,N_16198,N_17406);
nor U18568 (N_18568,N_16239,N_17218);
nand U18569 (N_18569,N_17174,N_16659);
nor U18570 (N_18570,N_16105,N_17103);
and U18571 (N_18571,N_17788,N_16849);
and U18572 (N_18572,N_17030,N_16567);
nand U18573 (N_18573,N_16843,N_16093);
and U18574 (N_18574,N_17894,N_17985);
xor U18575 (N_18575,N_16564,N_17100);
and U18576 (N_18576,N_17714,N_17239);
xor U18577 (N_18577,N_17360,N_17452);
or U18578 (N_18578,N_17827,N_16476);
nand U18579 (N_18579,N_17328,N_17975);
and U18580 (N_18580,N_17606,N_17687);
nor U18581 (N_18581,N_16942,N_17314);
xnor U18582 (N_18582,N_17802,N_16426);
and U18583 (N_18583,N_16821,N_16265);
or U18584 (N_18584,N_16377,N_17838);
nand U18585 (N_18585,N_17973,N_16054);
or U18586 (N_18586,N_16790,N_16302);
and U18587 (N_18587,N_17060,N_16744);
and U18588 (N_18588,N_16252,N_16464);
or U18589 (N_18589,N_17178,N_17987);
and U18590 (N_18590,N_17441,N_17019);
and U18591 (N_18591,N_17877,N_17183);
xor U18592 (N_18592,N_16203,N_17579);
nand U18593 (N_18593,N_17801,N_16868);
xnor U18594 (N_18594,N_16406,N_17976);
or U18595 (N_18595,N_17438,N_16829);
and U18596 (N_18596,N_16470,N_16701);
and U18597 (N_18597,N_16596,N_17382);
nand U18598 (N_18598,N_16927,N_17306);
or U18599 (N_18599,N_17832,N_16997);
nor U18600 (N_18600,N_17868,N_16616);
or U18601 (N_18601,N_16139,N_17159);
nor U18602 (N_18602,N_17212,N_17268);
xnor U18603 (N_18603,N_16022,N_17793);
nor U18604 (N_18604,N_16812,N_17898);
or U18605 (N_18605,N_16668,N_16756);
xor U18606 (N_18606,N_16909,N_16160);
or U18607 (N_18607,N_16588,N_17631);
nand U18608 (N_18608,N_16289,N_17799);
nor U18609 (N_18609,N_16707,N_17558);
or U18610 (N_18610,N_17427,N_16665);
nand U18611 (N_18611,N_16319,N_16618);
or U18612 (N_18612,N_17695,N_17483);
xor U18613 (N_18613,N_16471,N_16237);
xnor U18614 (N_18614,N_16295,N_16018);
nand U18615 (N_18615,N_16867,N_17147);
or U18616 (N_18616,N_16657,N_17358);
or U18617 (N_18617,N_16966,N_16531);
nor U18618 (N_18618,N_17512,N_16328);
and U18619 (N_18619,N_17741,N_16181);
or U18620 (N_18620,N_17847,N_16928);
or U18621 (N_18621,N_16496,N_17251);
nand U18622 (N_18622,N_17056,N_16629);
or U18623 (N_18623,N_17862,N_16108);
and U18624 (N_18624,N_17723,N_16673);
nand U18625 (N_18625,N_16172,N_16815);
xnor U18626 (N_18626,N_16537,N_17957);
nand U18627 (N_18627,N_16017,N_16246);
and U18628 (N_18628,N_16806,N_16286);
nor U18629 (N_18629,N_16980,N_16600);
or U18630 (N_18630,N_16469,N_16622);
nor U18631 (N_18631,N_16964,N_16234);
or U18632 (N_18632,N_17307,N_16736);
nand U18633 (N_18633,N_16184,N_16064);
and U18634 (N_18634,N_16951,N_17959);
or U18635 (N_18635,N_17880,N_16162);
and U18636 (N_18636,N_17956,N_17285);
nor U18637 (N_18637,N_16939,N_16327);
nand U18638 (N_18638,N_17201,N_16337);
nand U18639 (N_18639,N_16988,N_17746);
and U18640 (N_18640,N_16734,N_16008);
xor U18641 (N_18641,N_17734,N_16479);
nor U18642 (N_18642,N_16475,N_16726);
or U18643 (N_18643,N_17693,N_17853);
xnor U18644 (N_18644,N_16946,N_17461);
or U18645 (N_18645,N_16052,N_16638);
xnor U18646 (N_18646,N_17095,N_16727);
xor U18647 (N_18647,N_17433,N_17871);
xor U18648 (N_18648,N_16217,N_17005);
nand U18649 (N_18649,N_17424,N_17859);
xnor U18650 (N_18650,N_16109,N_16799);
xnor U18651 (N_18651,N_16758,N_17926);
nor U18652 (N_18652,N_16938,N_17786);
nor U18653 (N_18653,N_17042,N_16450);
xnor U18654 (N_18654,N_16776,N_16056);
nor U18655 (N_18655,N_17699,N_17794);
and U18656 (N_18656,N_16179,N_16244);
xnor U18657 (N_18657,N_16285,N_16741);
xor U18658 (N_18658,N_17155,N_16706);
nor U18659 (N_18659,N_17297,N_16060);
nor U18660 (N_18660,N_16077,N_17081);
and U18661 (N_18661,N_16150,N_16063);
or U18662 (N_18662,N_16846,N_16199);
or U18663 (N_18663,N_16211,N_16453);
nor U18664 (N_18664,N_17303,N_17038);
nand U18665 (N_18665,N_16323,N_17942);
and U18666 (N_18666,N_17751,N_17905);
xor U18667 (N_18667,N_17224,N_16057);
and U18668 (N_18668,N_17041,N_17250);
nand U18669 (N_18669,N_16943,N_17315);
xnor U18670 (N_18670,N_16329,N_16898);
or U18671 (N_18671,N_17105,N_16407);
and U18672 (N_18672,N_17335,N_16128);
nor U18673 (N_18673,N_16048,N_16175);
xnor U18674 (N_18674,N_16434,N_16705);
and U18675 (N_18675,N_16135,N_16382);
and U18676 (N_18676,N_16586,N_16700);
or U18677 (N_18677,N_16914,N_16718);
nand U18678 (N_18678,N_17166,N_16373);
xnor U18679 (N_18679,N_16313,N_17164);
nand U18680 (N_18680,N_16183,N_17097);
and U18681 (N_18681,N_16449,N_17521);
nor U18682 (N_18682,N_16793,N_17489);
or U18683 (N_18683,N_16499,N_17222);
nor U18684 (N_18684,N_16131,N_16002);
or U18685 (N_18685,N_16029,N_16926);
xnor U18686 (N_18686,N_16751,N_17445);
and U18687 (N_18687,N_16015,N_16076);
or U18688 (N_18688,N_16609,N_17295);
xnor U18689 (N_18689,N_17921,N_17678);
nor U18690 (N_18690,N_16348,N_17640);
or U18691 (N_18691,N_16034,N_17875);
or U18692 (N_18692,N_16509,N_16920);
or U18693 (N_18693,N_16856,N_17590);
or U18694 (N_18694,N_17198,N_17513);
nor U18695 (N_18695,N_16765,N_17596);
or U18696 (N_18696,N_17538,N_17949);
nor U18697 (N_18697,N_16345,N_17750);
nand U18698 (N_18698,N_16747,N_17206);
xor U18699 (N_18699,N_16798,N_17470);
xnor U18700 (N_18700,N_16961,N_17289);
nor U18701 (N_18701,N_16746,N_16641);
and U18702 (N_18702,N_16349,N_16921);
and U18703 (N_18703,N_17720,N_16859);
xor U18704 (N_18704,N_16425,N_16904);
or U18705 (N_18705,N_16092,N_17083);
nand U18706 (N_18706,N_17808,N_17825);
or U18707 (N_18707,N_16911,N_17900);
and U18708 (N_18708,N_17173,N_16732);
nor U18709 (N_18709,N_16789,N_16579);
and U18710 (N_18710,N_16404,N_16103);
nor U18711 (N_18711,N_16986,N_17840);
nand U18712 (N_18712,N_17730,N_16415);
nand U18713 (N_18713,N_16073,N_17290);
or U18714 (N_18714,N_16005,N_16317);
nor U18715 (N_18715,N_16045,N_16338);
nor U18716 (N_18716,N_16357,N_16513);
nor U18717 (N_18717,N_16389,N_17929);
nor U18718 (N_18718,N_16336,N_16519);
or U18719 (N_18719,N_17772,N_16379);
xnor U18720 (N_18720,N_16311,N_16791);
and U18721 (N_18721,N_16440,N_16021);
and U18722 (N_18722,N_17652,N_17806);
nor U18723 (N_18723,N_17302,N_16794);
and U18724 (N_18724,N_17659,N_16280);
nand U18725 (N_18725,N_17435,N_17602);
and U18726 (N_18726,N_16960,N_17187);
xnor U18727 (N_18727,N_17574,N_16534);
xnor U18728 (N_18728,N_17006,N_17641);
and U18729 (N_18729,N_16743,N_17028);
xor U18730 (N_18730,N_16435,N_16152);
nand U18731 (N_18731,N_17478,N_16740);
nand U18732 (N_18732,N_16500,N_16735);
xor U18733 (N_18733,N_17447,N_16714);
nor U18734 (N_18734,N_16353,N_16679);
nand U18735 (N_18735,N_16822,N_17550);
and U18736 (N_18736,N_17684,N_17508);
and U18737 (N_18737,N_17070,N_17153);
xor U18738 (N_18738,N_17176,N_17656);
or U18739 (N_18739,N_17570,N_17156);
nor U18740 (N_18740,N_17215,N_16646);
xnor U18741 (N_18741,N_16422,N_16653);
and U18742 (N_18742,N_17010,N_17494);
nor U18743 (N_18743,N_17626,N_16688);
nor U18744 (N_18744,N_16693,N_17701);
and U18745 (N_18745,N_16362,N_17502);
nor U18746 (N_18746,N_16785,N_17522);
xor U18747 (N_18747,N_17191,N_17932);
and U18748 (N_18748,N_16267,N_16748);
or U18749 (N_18749,N_16068,N_17370);
nand U18750 (N_18750,N_16774,N_16053);
nand U18751 (N_18751,N_16548,N_17694);
nand U18752 (N_18752,N_17219,N_17651);
and U18753 (N_18753,N_16408,N_16685);
and U18754 (N_18754,N_17904,N_16396);
nand U18755 (N_18755,N_17969,N_16019);
and U18756 (N_18756,N_17549,N_16191);
nor U18757 (N_18757,N_17960,N_16012);
or U18758 (N_18758,N_17484,N_16608);
xnor U18759 (N_18759,N_16035,N_17620);
and U18760 (N_18760,N_16678,N_17052);
xor U18761 (N_18761,N_16582,N_17525);
nand U18762 (N_18762,N_17702,N_16830);
and U18763 (N_18763,N_17317,N_16196);
or U18764 (N_18764,N_16595,N_16201);
nand U18765 (N_18765,N_17228,N_17339);
and U18766 (N_18766,N_16238,N_17207);
xor U18767 (N_18767,N_17063,N_17575);
nand U18768 (N_18768,N_17375,N_16633);
or U18769 (N_18769,N_17770,N_16702);
nand U18770 (N_18770,N_16819,N_17600);
nand U18771 (N_18771,N_17686,N_16300);
or U18772 (N_18772,N_17572,N_17396);
xnor U18773 (N_18773,N_16993,N_17988);
nor U18774 (N_18774,N_17878,N_17138);
nand U18775 (N_18775,N_16753,N_16143);
or U18776 (N_18776,N_17784,N_16376);
or U18777 (N_18777,N_17995,N_17142);
and U18778 (N_18778,N_16841,N_17257);
nor U18779 (N_18779,N_17914,N_17321);
xor U18780 (N_18780,N_17962,N_17688);
nand U18781 (N_18781,N_16801,N_16498);
nor U18782 (N_18782,N_16919,N_16436);
nand U18783 (N_18783,N_17479,N_16395);
nand U18784 (N_18784,N_16258,N_16530);
or U18785 (N_18785,N_17180,N_17143);
xnor U18786 (N_18786,N_17144,N_17937);
or U18787 (N_18787,N_16410,N_16214);
xnor U18788 (N_18788,N_16490,N_16343);
nor U18789 (N_18789,N_16550,N_16844);
nor U18790 (N_18790,N_17113,N_16594);
xnor U18791 (N_18791,N_17453,N_16137);
xor U18792 (N_18792,N_17330,N_16773);
or U18793 (N_18793,N_16402,N_16816);
nor U18794 (N_18794,N_16036,N_16301);
nand U18795 (N_18795,N_17768,N_17211);
nand U18796 (N_18796,N_17500,N_16878);
nand U18797 (N_18797,N_17909,N_17133);
and U18798 (N_18798,N_17874,N_17482);
and U18799 (N_18799,N_17408,N_17629);
and U18800 (N_18800,N_16058,N_17431);
xnor U18801 (N_18801,N_16331,N_16684);
or U18802 (N_18802,N_17280,N_17967);
or U18803 (N_18803,N_16578,N_16070);
or U18804 (N_18804,N_17420,N_17293);
xnor U18805 (N_18805,N_16708,N_17760);
nor U18806 (N_18806,N_17125,N_16126);
or U18807 (N_18807,N_16091,N_16102);
nand U18808 (N_18808,N_17476,N_16692);
nand U18809 (N_18809,N_17245,N_16631);
or U18810 (N_18810,N_16242,N_16561);
and U18811 (N_18811,N_17386,N_17021);
xor U18812 (N_18812,N_16383,N_16991);
xnor U18813 (N_18813,N_17145,N_17674);
or U18814 (N_18814,N_16209,N_17978);
nor U18815 (N_18815,N_16823,N_16632);
xor U18816 (N_18816,N_17779,N_16836);
nor U18817 (N_18817,N_17507,N_17294);
nor U18818 (N_18818,N_17221,N_17049);
and U18819 (N_18819,N_16524,N_17128);
xor U18820 (N_18820,N_16972,N_16224);
or U18821 (N_18821,N_16316,N_16009);
nand U18822 (N_18822,N_16835,N_17389);
xnor U18823 (N_18823,N_16266,N_16140);
nand U18824 (N_18824,N_16545,N_17401);
or U18825 (N_18825,N_17815,N_16346);
nor U18826 (N_18826,N_16605,N_17518);
and U18827 (N_18827,N_16535,N_17528);
or U18828 (N_18828,N_17035,N_16963);
nor U18829 (N_18829,N_17098,N_17368);
or U18830 (N_18830,N_16118,N_16122);
or U18831 (N_18831,N_17682,N_17168);
nand U18832 (N_18832,N_17765,N_16825);
or U18833 (N_18833,N_16194,N_16542);
and U18834 (N_18834,N_17654,N_17740);
nand U18835 (N_18835,N_17249,N_17356);
nand U18836 (N_18836,N_17619,N_17776);
nor U18837 (N_18837,N_16516,N_17440);
xnor U18838 (N_18838,N_16603,N_16114);
xor U18839 (N_18839,N_16521,N_16591);
and U18840 (N_18840,N_16281,N_16650);
nand U18841 (N_18841,N_16837,N_17872);
xnor U18842 (N_18842,N_16583,N_16892);
xnor U18843 (N_18843,N_16007,N_17539);
or U18844 (N_18844,N_17782,N_17485);
nand U18845 (N_18845,N_16780,N_17077);
xnor U18846 (N_18846,N_16419,N_17185);
or U18847 (N_18847,N_17561,N_16874);
xor U18848 (N_18848,N_16290,N_17984);
nand U18849 (N_18849,N_17893,N_17553);
xnor U18850 (N_18850,N_16307,N_16808);
and U18851 (N_18851,N_17377,N_17291);
xor U18852 (N_18852,N_16536,N_17665);
xnor U18853 (N_18853,N_17393,N_17888);
nor U18854 (N_18854,N_17846,N_17621);
nor U18855 (N_18855,N_17376,N_17346);
or U18856 (N_18856,N_16256,N_16315);
or U18857 (N_18857,N_16696,N_16865);
nor U18858 (N_18858,N_17516,N_16528);
nand U18859 (N_18859,N_16838,N_16802);
xor U18860 (N_18860,N_16483,N_16887);
nand U18861 (N_18861,N_16848,N_16342);
nand U18862 (N_18862,N_17902,N_16503);
xor U18863 (N_18863,N_16061,N_17991);
nor U18864 (N_18864,N_16508,N_17964);
nand U18865 (N_18865,N_17243,N_17842);
nor U18866 (N_18866,N_16233,N_16686);
xnor U18867 (N_18867,N_17982,N_16263);
or U18868 (N_18868,N_16664,N_16024);
xnor U18869 (N_18869,N_16884,N_16971);
or U18870 (N_18870,N_17910,N_16712);
nor U18871 (N_18871,N_17200,N_17628);
nor U18872 (N_18872,N_16584,N_17814);
nand U18873 (N_18873,N_16715,N_16480);
nand U18874 (N_18874,N_17843,N_16984);
nor U18875 (N_18875,N_16681,N_17443);
nand U18876 (N_18876,N_17526,N_16204);
or U18877 (N_18877,N_17617,N_16875);
xnor U18878 (N_18878,N_17603,N_17165);
or U18879 (N_18879,N_17398,N_17527);
nor U18880 (N_18880,N_16361,N_16626);
or U18881 (N_18881,N_16080,N_16473);
nand U18882 (N_18882,N_16387,N_16192);
xor U18883 (N_18883,N_16392,N_17002);
xor U18884 (N_18884,N_16787,N_17771);
nand U18885 (N_18885,N_17906,N_16680);
xnor U18886 (N_18886,N_17671,N_16769);
nand U18887 (N_18887,N_16084,N_17372);
and U18888 (N_18888,N_16923,N_16525);
xor U18889 (N_18889,N_17657,N_17664);
and U18890 (N_18890,N_16200,N_16557);
nand U18891 (N_18891,N_17680,N_16158);
and U18892 (N_18892,N_16936,N_17823);
or U18893 (N_18893,N_16132,N_17805);
nor U18894 (N_18894,N_17234,N_16299);
xor U18895 (N_18895,N_16949,N_16394);
or U18896 (N_18896,N_17101,N_16151);
or U18897 (N_18897,N_17151,N_16261);
nand U18898 (N_18898,N_17170,N_17917);
nor U18899 (N_18899,N_16028,N_16442);
and U18900 (N_18900,N_17194,N_17265);
xnor U18901 (N_18901,N_16532,N_17305);
and U18902 (N_18902,N_17008,N_16381);
or U18903 (N_18903,N_17208,N_16145);
nor U18904 (N_18904,N_16768,N_16902);
nand U18905 (N_18905,N_16458,N_16908);
nor U18906 (N_18906,N_17869,N_16367);
nor U18907 (N_18907,N_16166,N_16115);
or U18908 (N_18908,N_17039,N_16592);
xnor U18909 (N_18909,N_16771,N_16446);
xnor U18910 (N_18910,N_16010,N_16671);
nand U18911 (N_18911,N_16223,N_16292);
xor U18912 (N_18912,N_17459,N_16393);
xor U18913 (N_18913,N_16893,N_17276);
nand U18914 (N_18914,N_16934,N_16711);
xnor U18915 (N_18915,N_17475,N_17506);
or U18916 (N_18916,N_17947,N_17858);
nor U18917 (N_18917,N_16334,N_17672);
nor U18918 (N_18918,N_16973,N_16719);
or U18919 (N_18919,N_17258,N_16006);
nand U18920 (N_18920,N_16454,N_17721);
nand U18921 (N_18921,N_17082,N_17685);
xnor U18922 (N_18922,N_17472,N_16120);
and U18923 (N_18923,N_17899,N_17696);
and U18924 (N_18924,N_17141,N_16250);
and U18925 (N_18925,N_17357,N_17235);
or U18926 (N_18926,N_16484,N_16227);
and U18927 (N_18927,N_17924,N_16413);
xor U18928 (N_18928,N_17944,N_16079);
nand U18929 (N_18929,N_17608,N_16778);
or U18930 (N_18930,N_16430,N_17012);
and U18931 (N_18931,N_16447,N_17188);
nand U18932 (N_18932,N_17361,N_16721);
nor U18933 (N_18933,N_17009,N_16180);
or U18934 (N_18934,N_16803,N_16897);
nor U18935 (N_18935,N_17365,N_17609);
and U18936 (N_18936,N_17017,N_16931);
nand U18937 (N_18937,N_16655,N_17743);
or U18938 (N_18938,N_16900,N_17385);
and U18939 (N_18939,N_17588,N_17345);
nand U18940 (N_18940,N_17655,N_16230);
and U18941 (N_18941,N_17819,N_17916);
nor U18942 (N_18942,N_17754,N_16930);
xnor U18943 (N_18943,N_16178,N_16365);
nand U18944 (N_18944,N_17350,N_17186);
xnor U18945 (N_18945,N_16090,N_16474);
or U18946 (N_18946,N_17717,N_17175);
and U18947 (N_18947,N_17413,N_16709);
or U18948 (N_18948,N_16871,N_17998);
xnor U18949 (N_18949,N_17509,N_16729);
nand U18950 (N_18950,N_16168,N_17972);
nor U18951 (N_18951,N_16720,N_17065);
nand U18952 (N_18952,N_17402,N_16666);
or U18953 (N_18953,N_16040,N_16428);
nand U18954 (N_18954,N_16598,N_16027);
and U18955 (N_18955,N_17727,N_16739);
nand U18956 (N_18956,N_16547,N_16182);
nor U18957 (N_18957,N_17352,N_17448);
or U18958 (N_18958,N_16554,N_17182);
or U18959 (N_18959,N_17737,N_17312);
nor U18960 (N_18960,N_16298,N_16322);
or U18961 (N_18961,N_16656,N_17818);
xor U18962 (N_18962,N_17925,N_17683);
nand U18963 (N_18963,N_16571,N_16444);
nor U18964 (N_18964,N_16967,N_16254);
or U18965 (N_18965,N_16144,N_16117);
or U18966 (N_18966,N_16866,N_16506);
xnor U18967 (N_18967,N_17744,N_16321);
xnor U18968 (N_18968,N_17126,N_16954);
nand U18969 (N_18969,N_16119,N_17551);
nor U18970 (N_18970,N_16767,N_16514);
and U18971 (N_18971,N_16344,N_16820);
nor U18972 (N_18972,N_17612,N_16262);
nand U18973 (N_18973,N_17468,N_17076);
nand U18974 (N_18974,N_17320,N_16565);
and U18975 (N_18975,N_17565,N_16208);
xnor U18976 (N_18976,N_16355,N_17354);
nor U18977 (N_18977,N_17067,N_17284);
and U18978 (N_18978,N_16424,N_16100);
or U18979 (N_18979,N_16800,N_16188);
xor U18980 (N_18980,N_17477,N_16001);
and U18981 (N_18981,N_16628,N_16279);
xnor U18982 (N_18982,N_17515,N_16649);
nand U18983 (N_18983,N_17428,N_17205);
or U18984 (N_18984,N_17934,N_16894);
and U18985 (N_18985,N_17630,N_16905);
nor U18986 (N_18986,N_17758,N_16690);
nand U18987 (N_18987,N_17885,N_16669);
xor U18988 (N_18988,N_16463,N_16924);
nor U18989 (N_18989,N_16876,N_17764);
xor U18990 (N_18990,N_16903,N_17053);
and U18991 (N_18991,N_17149,N_16421);
nor U18992 (N_18992,N_17830,N_16016);
nor U18993 (N_18993,N_16472,N_16386);
nor U18994 (N_18994,N_17269,N_17004);
nand U18995 (N_18995,N_16885,N_16643);
nor U18996 (N_18996,N_17735,N_17713);
or U18997 (N_18997,N_16461,N_17450);
and U18998 (N_18998,N_17496,N_17319);
xnor U18999 (N_18999,N_17381,N_16749);
xnor U19000 (N_19000,N_16284,N_17456);
nand U19001 (N_19001,N_17142,N_17679);
xnor U19002 (N_19002,N_16703,N_17385);
nor U19003 (N_19003,N_16706,N_16947);
xor U19004 (N_19004,N_16677,N_16823);
nand U19005 (N_19005,N_16757,N_16729);
or U19006 (N_19006,N_17215,N_17708);
xnor U19007 (N_19007,N_16001,N_16002);
nand U19008 (N_19008,N_17720,N_17464);
nor U19009 (N_19009,N_17000,N_16492);
and U19010 (N_19010,N_16242,N_17113);
and U19011 (N_19011,N_17048,N_16409);
nor U19012 (N_19012,N_17510,N_17773);
or U19013 (N_19013,N_17279,N_16721);
xnor U19014 (N_19014,N_17389,N_17684);
and U19015 (N_19015,N_17171,N_17445);
nor U19016 (N_19016,N_16576,N_17337);
or U19017 (N_19017,N_16493,N_17640);
or U19018 (N_19018,N_16364,N_16065);
nor U19019 (N_19019,N_17921,N_16893);
or U19020 (N_19020,N_17326,N_16514);
xor U19021 (N_19021,N_17375,N_17529);
xnor U19022 (N_19022,N_17728,N_16425);
nor U19023 (N_19023,N_16228,N_17180);
and U19024 (N_19024,N_17834,N_17149);
nor U19025 (N_19025,N_16535,N_16265);
and U19026 (N_19026,N_17569,N_17187);
xor U19027 (N_19027,N_17524,N_17695);
xor U19028 (N_19028,N_17301,N_17318);
xor U19029 (N_19029,N_17400,N_17419);
xnor U19030 (N_19030,N_17803,N_17754);
and U19031 (N_19031,N_16148,N_17737);
and U19032 (N_19032,N_16124,N_16934);
and U19033 (N_19033,N_16233,N_17577);
or U19034 (N_19034,N_17271,N_16543);
nor U19035 (N_19035,N_16454,N_17434);
or U19036 (N_19036,N_16161,N_17328);
xor U19037 (N_19037,N_16857,N_17136);
nand U19038 (N_19038,N_17722,N_16095);
or U19039 (N_19039,N_16140,N_16959);
or U19040 (N_19040,N_16538,N_17305);
or U19041 (N_19041,N_17301,N_16602);
nand U19042 (N_19042,N_17991,N_17678);
xor U19043 (N_19043,N_17645,N_16606);
or U19044 (N_19044,N_16549,N_16343);
nor U19045 (N_19045,N_16226,N_16332);
nand U19046 (N_19046,N_17799,N_16581);
nand U19047 (N_19047,N_16924,N_17181);
and U19048 (N_19048,N_17876,N_16775);
nand U19049 (N_19049,N_17553,N_16564);
nand U19050 (N_19050,N_17197,N_17907);
or U19051 (N_19051,N_17146,N_17768);
xor U19052 (N_19052,N_17887,N_17715);
nand U19053 (N_19053,N_16668,N_16759);
or U19054 (N_19054,N_16163,N_16314);
xnor U19055 (N_19055,N_17582,N_16041);
nand U19056 (N_19056,N_17615,N_16420);
and U19057 (N_19057,N_16936,N_16840);
nand U19058 (N_19058,N_16156,N_17501);
xor U19059 (N_19059,N_16493,N_17298);
and U19060 (N_19060,N_16083,N_16719);
xor U19061 (N_19061,N_16804,N_16784);
nor U19062 (N_19062,N_17935,N_16701);
nand U19063 (N_19063,N_16727,N_16211);
nor U19064 (N_19064,N_16382,N_16503);
nor U19065 (N_19065,N_17220,N_16720);
and U19066 (N_19066,N_17704,N_16865);
and U19067 (N_19067,N_16530,N_17354);
nor U19068 (N_19068,N_16192,N_17043);
nand U19069 (N_19069,N_16905,N_17717);
xor U19070 (N_19070,N_16035,N_16643);
and U19071 (N_19071,N_16595,N_16562);
or U19072 (N_19072,N_16962,N_17023);
nand U19073 (N_19073,N_17274,N_17489);
or U19074 (N_19074,N_16037,N_16386);
nand U19075 (N_19075,N_17897,N_17335);
nand U19076 (N_19076,N_16230,N_16991);
nand U19077 (N_19077,N_16787,N_17960);
and U19078 (N_19078,N_17164,N_16723);
nor U19079 (N_19079,N_16596,N_17075);
xor U19080 (N_19080,N_17929,N_16830);
nor U19081 (N_19081,N_17880,N_17418);
xnor U19082 (N_19082,N_17750,N_16524);
or U19083 (N_19083,N_16307,N_16611);
xor U19084 (N_19084,N_16019,N_17987);
or U19085 (N_19085,N_16454,N_16732);
nand U19086 (N_19086,N_17077,N_17729);
and U19087 (N_19087,N_16348,N_16918);
or U19088 (N_19088,N_16556,N_16924);
and U19089 (N_19089,N_17645,N_16987);
and U19090 (N_19090,N_16608,N_16118);
xnor U19091 (N_19091,N_17084,N_17444);
nand U19092 (N_19092,N_17268,N_17685);
nand U19093 (N_19093,N_17874,N_16425);
and U19094 (N_19094,N_17695,N_16230);
or U19095 (N_19095,N_16367,N_17485);
or U19096 (N_19096,N_16010,N_16012);
or U19097 (N_19097,N_17113,N_17762);
xor U19098 (N_19098,N_17044,N_16154);
and U19099 (N_19099,N_17743,N_16532);
xor U19100 (N_19100,N_16978,N_17721);
or U19101 (N_19101,N_16828,N_17042);
and U19102 (N_19102,N_17021,N_17269);
or U19103 (N_19103,N_16311,N_17705);
nor U19104 (N_19104,N_16856,N_16862);
xor U19105 (N_19105,N_17891,N_17057);
and U19106 (N_19106,N_16559,N_16841);
or U19107 (N_19107,N_16951,N_17786);
xnor U19108 (N_19108,N_16626,N_17517);
nor U19109 (N_19109,N_17396,N_16307);
nand U19110 (N_19110,N_17930,N_17079);
or U19111 (N_19111,N_17464,N_17994);
or U19112 (N_19112,N_16703,N_16694);
nor U19113 (N_19113,N_16127,N_17675);
nor U19114 (N_19114,N_16022,N_16756);
and U19115 (N_19115,N_17667,N_17806);
and U19116 (N_19116,N_16003,N_16310);
nor U19117 (N_19117,N_17478,N_16949);
nand U19118 (N_19118,N_17254,N_17109);
nor U19119 (N_19119,N_16781,N_17019);
or U19120 (N_19120,N_17055,N_16567);
nand U19121 (N_19121,N_17772,N_17962);
nor U19122 (N_19122,N_16861,N_17080);
xor U19123 (N_19123,N_17082,N_17513);
and U19124 (N_19124,N_16850,N_16961);
xnor U19125 (N_19125,N_16086,N_17459);
or U19126 (N_19126,N_17387,N_16342);
nand U19127 (N_19127,N_17429,N_17852);
or U19128 (N_19128,N_16766,N_16833);
and U19129 (N_19129,N_16126,N_16778);
and U19130 (N_19130,N_17633,N_16773);
or U19131 (N_19131,N_16232,N_17465);
nor U19132 (N_19132,N_16257,N_17967);
or U19133 (N_19133,N_16361,N_16025);
xor U19134 (N_19134,N_16961,N_16848);
or U19135 (N_19135,N_17930,N_17369);
or U19136 (N_19136,N_16439,N_17798);
nand U19137 (N_19137,N_16824,N_17222);
and U19138 (N_19138,N_16191,N_16406);
nor U19139 (N_19139,N_17194,N_17251);
nand U19140 (N_19140,N_16748,N_17497);
nand U19141 (N_19141,N_17564,N_16976);
nor U19142 (N_19142,N_17302,N_16993);
xnor U19143 (N_19143,N_16390,N_16638);
xnor U19144 (N_19144,N_16748,N_16393);
nand U19145 (N_19145,N_17399,N_17739);
xnor U19146 (N_19146,N_17472,N_17889);
xnor U19147 (N_19147,N_17712,N_17192);
or U19148 (N_19148,N_17403,N_16820);
and U19149 (N_19149,N_16679,N_17117);
or U19150 (N_19150,N_16516,N_17909);
and U19151 (N_19151,N_16136,N_17774);
or U19152 (N_19152,N_16031,N_17999);
and U19153 (N_19153,N_16515,N_17185);
or U19154 (N_19154,N_16947,N_16862);
nor U19155 (N_19155,N_16907,N_17272);
xnor U19156 (N_19156,N_17691,N_17817);
and U19157 (N_19157,N_17846,N_16357);
nor U19158 (N_19158,N_17130,N_16367);
nand U19159 (N_19159,N_16132,N_16283);
nor U19160 (N_19160,N_17991,N_16547);
nand U19161 (N_19161,N_16689,N_16171);
nand U19162 (N_19162,N_17702,N_17168);
and U19163 (N_19163,N_16864,N_17484);
nand U19164 (N_19164,N_17274,N_16368);
nor U19165 (N_19165,N_17137,N_16402);
xnor U19166 (N_19166,N_17900,N_17354);
nor U19167 (N_19167,N_17245,N_17234);
xor U19168 (N_19168,N_16339,N_17616);
nor U19169 (N_19169,N_17123,N_16762);
nand U19170 (N_19170,N_17752,N_16385);
and U19171 (N_19171,N_16264,N_17312);
nor U19172 (N_19172,N_16569,N_16302);
and U19173 (N_19173,N_17085,N_16722);
nor U19174 (N_19174,N_17612,N_17766);
or U19175 (N_19175,N_16488,N_16453);
and U19176 (N_19176,N_16003,N_16461);
nor U19177 (N_19177,N_16032,N_16925);
nand U19178 (N_19178,N_16703,N_17054);
nand U19179 (N_19179,N_16182,N_16795);
and U19180 (N_19180,N_16009,N_16193);
xor U19181 (N_19181,N_17514,N_16738);
and U19182 (N_19182,N_16083,N_17148);
xor U19183 (N_19183,N_17670,N_16718);
nor U19184 (N_19184,N_16724,N_17282);
or U19185 (N_19185,N_16975,N_17841);
nand U19186 (N_19186,N_17586,N_16776);
nand U19187 (N_19187,N_16125,N_16328);
and U19188 (N_19188,N_16406,N_16767);
nor U19189 (N_19189,N_16217,N_17414);
nand U19190 (N_19190,N_17263,N_17796);
xnor U19191 (N_19191,N_17473,N_16884);
nor U19192 (N_19192,N_17563,N_17056);
xnor U19193 (N_19193,N_17875,N_16983);
xor U19194 (N_19194,N_16182,N_16647);
nor U19195 (N_19195,N_16749,N_17166);
nor U19196 (N_19196,N_17625,N_17258);
and U19197 (N_19197,N_17468,N_16316);
nor U19198 (N_19198,N_17865,N_16560);
nor U19199 (N_19199,N_17822,N_16460);
nand U19200 (N_19200,N_16299,N_16735);
nand U19201 (N_19201,N_17860,N_16380);
and U19202 (N_19202,N_17291,N_17251);
and U19203 (N_19203,N_16724,N_17112);
xnor U19204 (N_19204,N_17792,N_16312);
nor U19205 (N_19205,N_17118,N_16589);
and U19206 (N_19206,N_16230,N_17613);
nand U19207 (N_19207,N_17374,N_17809);
nand U19208 (N_19208,N_17278,N_16188);
and U19209 (N_19209,N_16681,N_16656);
nor U19210 (N_19210,N_17868,N_17445);
or U19211 (N_19211,N_17991,N_16795);
nor U19212 (N_19212,N_17495,N_17995);
or U19213 (N_19213,N_17965,N_17968);
nand U19214 (N_19214,N_17211,N_17888);
nor U19215 (N_19215,N_17522,N_17961);
or U19216 (N_19216,N_17650,N_16775);
or U19217 (N_19217,N_16819,N_16606);
or U19218 (N_19218,N_17633,N_16703);
or U19219 (N_19219,N_16880,N_17526);
nand U19220 (N_19220,N_17584,N_16472);
nor U19221 (N_19221,N_16601,N_16782);
nor U19222 (N_19222,N_16892,N_16978);
nand U19223 (N_19223,N_16078,N_17569);
nor U19224 (N_19224,N_16187,N_16932);
nor U19225 (N_19225,N_17423,N_16346);
nor U19226 (N_19226,N_17896,N_17748);
nand U19227 (N_19227,N_17045,N_17917);
xnor U19228 (N_19228,N_17212,N_16431);
and U19229 (N_19229,N_16120,N_16978);
xor U19230 (N_19230,N_17161,N_16213);
xor U19231 (N_19231,N_17850,N_16848);
xor U19232 (N_19232,N_16229,N_16217);
xnor U19233 (N_19233,N_17903,N_16389);
and U19234 (N_19234,N_17825,N_16838);
xnor U19235 (N_19235,N_16083,N_17765);
and U19236 (N_19236,N_16660,N_16091);
xnor U19237 (N_19237,N_16524,N_17823);
or U19238 (N_19238,N_16163,N_17443);
or U19239 (N_19239,N_16033,N_16605);
xor U19240 (N_19240,N_17270,N_17442);
or U19241 (N_19241,N_17987,N_17157);
xor U19242 (N_19242,N_16494,N_16237);
or U19243 (N_19243,N_16746,N_17420);
xnor U19244 (N_19244,N_16028,N_16659);
nor U19245 (N_19245,N_16709,N_17555);
and U19246 (N_19246,N_16788,N_16923);
and U19247 (N_19247,N_17684,N_16498);
nand U19248 (N_19248,N_16737,N_16176);
or U19249 (N_19249,N_16508,N_16266);
xor U19250 (N_19250,N_16077,N_16881);
and U19251 (N_19251,N_16065,N_16769);
xor U19252 (N_19252,N_17230,N_16219);
and U19253 (N_19253,N_17196,N_17284);
and U19254 (N_19254,N_16824,N_17925);
nand U19255 (N_19255,N_16208,N_16534);
and U19256 (N_19256,N_17079,N_17772);
and U19257 (N_19257,N_17252,N_16195);
nor U19258 (N_19258,N_16310,N_17160);
and U19259 (N_19259,N_17044,N_17741);
nor U19260 (N_19260,N_17450,N_17403);
nor U19261 (N_19261,N_16623,N_17223);
or U19262 (N_19262,N_16415,N_17213);
or U19263 (N_19263,N_16105,N_16386);
nor U19264 (N_19264,N_16332,N_17638);
xnor U19265 (N_19265,N_16886,N_17606);
or U19266 (N_19266,N_17230,N_16066);
xor U19267 (N_19267,N_17881,N_17260);
nand U19268 (N_19268,N_17395,N_16253);
xor U19269 (N_19269,N_16192,N_17762);
nand U19270 (N_19270,N_17143,N_17598);
xor U19271 (N_19271,N_16784,N_16800);
nor U19272 (N_19272,N_16696,N_17318);
nor U19273 (N_19273,N_16513,N_17331);
and U19274 (N_19274,N_17994,N_16554);
xor U19275 (N_19275,N_17071,N_16115);
and U19276 (N_19276,N_16614,N_17885);
nand U19277 (N_19277,N_17588,N_17186);
nor U19278 (N_19278,N_17838,N_17185);
nor U19279 (N_19279,N_17605,N_16391);
nand U19280 (N_19280,N_16108,N_16231);
xor U19281 (N_19281,N_16116,N_17507);
or U19282 (N_19282,N_16250,N_16247);
or U19283 (N_19283,N_17210,N_17872);
and U19284 (N_19284,N_16636,N_16277);
and U19285 (N_19285,N_17928,N_16952);
nand U19286 (N_19286,N_16080,N_17792);
or U19287 (N_19287,N_17505,N_16437);
nor U19288 (N_19288,N_17387,N_16805);
or U19289 (N_19289,N_17278,N_16295);
and U19290 (N_19290,N_17193,N_16410);
xor U19291 (N_19291,N_16919,N_16851);
or U19292 (N_19292,N_17304,N_16098);
or U19293 (N_19293,N_17427,N_16235);
or U19294 (N_19294,N_16605,N_17833);
nand U19295 (N_19295,N_16547,N_17413);
nand U19296 (N_19296,N_16758,N_17919);
and U19297 (N_19297,N_17523,N_16363);
nor U19298 (N_19298,N_16703,N_17446);
and U19299 (N_19299,N_17438,N_16379);
nor U19300 (N_19300,N_17122,N_17158);
and U19301 (N_19301,N_16202,N_16275);
xor U19302 (N_19302,N_17521,N_16056);
xor U19303 (N_19303,N_16770,N_17522);
and U19304 (N_19304,N_17656,N_16649);
nand U19305 (N_19305,N_17776,N_17146);
nor U19306 (N_19306,N_17064,N_17412);
nor U19307 (N_19307,N_17464,N_16067);
and U19308 (N_19308,N_16198,N_16131);
nor U19309 (N_19309,N_17453,N_16420);
and U19310 (N_19310,N_17142,N_17070);
nor U19311 (N_19311,N_17506,N_16578);
or U19312 (N_19312,N_16809,N_17729);
nor U19313 (N_19313,N_16607,N_17894);
xor U19314 (N_19314,N_17077,N_17061);
or U19315 (N_19315,N_17633,N_16939);
xor U19316 (N_19316,N_16656,N_16766);
or U19317 (N_19317,N_17271,N_17316);
nor U19318 (N_19318,N_17165,N_16334);
nor U19319 (N_19319,N_17609,N_17079);
xnor U19320 (N_19320,N_17144,N_16464);
xor U19321 (N_19321,N_16973,N_17704);
or U19322 (N_19322,N_17264,N_16336);
xor U19323 (N_19323,N_16372,N_16472);
and U19324 (N_19324,N_16527,N_17872);
nor U19325 (N_19325,N_16337,N_17897);
or U19326 (N_19326,N_17519,N_17502);
and U19327 (N_19327,N_17705,N_17910);
nor U19328 (N_19328,N_16677,N_16885);
and U19329 (N_19329,N_16827,N_16658);
or U19330 (N_19330,N_16893,N_17849);
and U19331 (N_19331,N_17934,N_16456);
or U19332 (N_19332,N_17336,N_16511);
and U19333 (N_19333,N_16603,N_17686);
or U19334 (N_19334,N_17493,N_17075);
nand U19335 (N_19335,N_16664,N_17258);
nor U19336 (N_19336,N_16409,N_16103);
xor U19337 (N_19337,N_16737,N_16154);
xor U19338 (N_19338,N_16860,N_17185);
and U19339 (N_19339,N_17655,N_16380);
nand U19340 (N_19340,N_17998,N_16655);
nand U19341 (N_19341,N_16623,N_17946);
and U19342 (N_19342,N_16761,N_16388);
and U19343 (N_19343,N_16310,N_16090);
nand U19344 (N_19344,N_17617,N_16642);
and U19345 (N_19345,N_17499,N_17467);
xor U19346 (N_19346,N_16965,N_16359);
or U19347 (N_19347,N_16771,N_17035);
xnor U19348 (N_19348,N_16297,N_17514);
or U19349 (N_19349,N_16270,N_17199);
and U19350 (N_19350,N_16425,N_16114);
nand U19351 (N_19351,N_16430,N_16332);
xnor U19352 (N_19352,N_16492,N_17184);
nor U19353 (N_19353,N_17246,N_17126);
nand U19354 (N_19354,N_16745,N_17047);
and U19355 (N_19355,N_16204,N_16606);
and U19356 (N_19356,N_16756,N_17958);
and U19357 (N_19357,N_16194,N_17455);
xor U19358 (N_19358,N_16859,N_16913);
and U19359 (N_19359,N_17598,N_16720);
nand U19360 (N_19360,N_17331,N_16227);
nand U19361 (N_19361,N_17167,N_17704);
xor U19362 (N_19362,N_17113,N_16304);
nand U19363 (N_19363,N_16927,N_16110);
nand U19364 (N_19364,N_16732,N_17984);
nor U19365 (N_19365,N_16962,N_17387);
or U19366 (N_19366,N_16448,N_17664);
or U19367 (N_19367,N_17777,N_17449);
nand U19368 (N_19368,N_17669,N_16027);
nand U19369 (N_19369,N_16150,N_16974);
xor U19370 (N_19370,N_17406,N_17436);
xor U19371 (N_19371,N_17475,N_16277);
nand U19372 (N_19372,N_17509,N_16490);
xnor U19373 (N_19373,N_17309,N_17552);
or U19374 (N_19374,N_17351,N_17949);
and U19375 (N_19375,N_16325,N_16798);
xor U19376 (N_19376,N_16553,N_16600);
nand U19377 (N_19377,N_17215,N_17176);
nor U19378 (N_19378,N_16728,N_17336);
nand U19379 (N_19379,N_17461,N_16817);
or U19380 (N_19380,N_16409,N_16138);
and U19381 (N_19381,N_16484,N_17914);
and U19382 (N_19382,N_16990,N_16957);
xor U19383 (N_19383,N_17057,N_16278);
and U19384 (N_19384,N_16126,N_16322);
nand U19385 (N_19385,N_16899,N_17961);
xor U19386 (N_19386,N_16845,N_16343);
nand U19387 (N_19387,N_16905,N_17293);
or U19388 (N_19388,N_16714,N_17240);
and U19389 (N_19389,N_17093,N_16430);
nor U19390 (N_19390,N_16274,N_17211);
nand U19391 (N_19391,N_17946,N_16397);
nand U19392 (N_19392,N_17376,N_16659);
xnor U19393 (N_19393,N_16285,N_17688);
nor U19394 (N_19394,N_17685,N_16298);
or U19395 (N_19395,N_17051,N_17992);
xor U19396 (N_19396,N_16221,N_17870);
nand U19397 (N_19397,N_17738,N_16412);
or U19398 (N_19398,N_17682,N_16683);
and U19399 (N_19399,N_17332,N_16650);
or U19400 (N_19400,N_16473,N_17248);
nand U19401 (N_19401,N_17471,N_16086);
or U19402 (N_19402,N_16292,N_17235);
and U19403 (N_19403,N_16836,N_17736);
xor U19404 (N_19404,N_16305,N_17225);
nand U19405 (N_19405,N_17088,N_16969);
or U19406 (N_19406,N_17572,N_17000);
or U19407 (N_19407,N_17787,N_16895);
nor U19408 (N_19408,N_16482,N_16452);
xnor U19409 (N_19409,N_16343,N_16726);
or U19410 (N_19410,N_16189,N_17422);
xnor U19411 (N_19411,N_16736,N_17256);
nand U19412 (N_19412,N_16528,N_16539);
nor U19413 (N_19413,N_16435,N_16127);
nand U19414 (N_19414,N_17460,N_17826);
xnor U19415 (N_19415,N_16141,N_16742);
nor U19416 (N_19416,N_17713,N_16931);
nand U19417 (N_19417,N_16194,N_16188);
nor U19418 (N_19418,N_16519,N_16095);
and U19419 (N_19419,N_17185,N_17693);
xnor U19420 (N_19420,N_16075,N_16155);
and U19421 (N_19421,N_16463,N_16865);
nor U19422 (N_19422,N_17097,N_16394);
xor U19423 (N_19423,N_16818,N_17906);
or U19424 (N_19424,N_16250,N_17058);
and U19425 (N_19425,N_17729,N_16766);
or U19426 (N_19426,N_17096,N_17546);
nor U19427 (N_19427,N_16701,N_16069);
and U19428 (N_19428,N_17836,N_17432);
nor U19429 (N_19429,N_16105,N_16754);
nand U19430 (N_19430,N_16362,N_17189);
and U19431 (N_19431,N_16658,N_17164);
nand U19432 (N_19432,N_17609,N_17236);
and U19433 (N_19433,N_16739,N_17811);
nand U19434 (N_19434,N_17266,N_17953);
nand U19435 (N_19435,N_17900,N_16424);
nor U19436 (N_19436,N_16670,N_17646);
nor U19437 (N_19437,N_16536,N_16394);
or U19438 (N_19438,N_16573,N_16241);
xor U19439 (N_19439,N_17190,N_16122);
nand U19440 (N_19440,N_17902,N_16773);
xor U19441 (N_19441,N_17574,N_16958);
nor U19442 (N_19442,N_17445,N_16123);
or U19443 (N_19443,N_17892,N_17911);
or U19444 (N_19444,N_16265,N_16469);
xnor U19445 (N_19445,N_17374,N_16373);
nor U19446 (N_19446,N_16624,N_16425);
and U19447 (N_19447,N_16150,N_17499);
nor U19448 (N_19448,N_17836,N_16149);
nand U19449 (N_19449,N_16854,N_17847);
xor U19450 (N_19450,N_17784,N_17052);
nor U19451 (N_19451,N_16306,N_16450);
and U19452 (N_19452,N_16492,N_16266);
nor U19453 (N_19453,N_17754,N_16032);
nor U19454 (N_19454,N_17877,N_16134);
nor U19455 (N_19455,N_17056,N_16162);
and U19456 (N_19456,N_16488,N_17340);
nor U19457 (N_19457,N_17596,N_16307);
nor U19458 (N_19458,N_17016,N_17608);
xnor U19459 (N_19459,N_17473,N_16451);
or U19460 (N_19460,N_17238,N_16142);
and U19461 (N_19461,N_16218,N_16083);
and U19462 (N_19462,N_16973,N_17405);
or U19463 (N_19463,N_16592,N_16426);
nand U19464 (N_19464,N_17922,N_17113);
xnor U19465 (N_19465,N_17056,N_17697);
or U19466 (N_19466,N_17608,N_17764);
nand U19467 (N_19467,N_16960,N_16184);
and U19468 (N_19468,N_16661,N_17155);
or U19469 (N_19469,N_17700,N_16664);
xor U19470 (N_19470,N_16715,N_17631);
or U19471 (N_19471,N_17108,N_16647);
nor U19472 (N_19472,N_17542,N_16742);
nand U19473 (N_19473,N_17318,N_16478);
or U19474 (N_19474,N_17833,N_17295);
nor U19475 (N_19475,N_17862,N_16215);
nand U19476 (N_19476,N_16333,N_16633);
nor U19477 (N_19477,N_16621,N_16061);
nor U19478 (N_19478,N_16537,N_17271);
nor U19479 (N_19479,N_16087,N_16002);
nand U19480 (N_19480,N_17459,N_17042);
nand U19481 (N_19481,N_17008,N_16460);
or U19482 (N_19482,N_17618,N_17651);
xnor U19483 (N_19483,N_16223,N_17259);
nor U19484 (N_19484,N_17971,N_17497);
xnor U19485 (N_19485,N_17333,N_17618);
or U19486 (N_19486,N_17639,N_16724);
nand U19487 (N_19487,N_17074,N_17897);
and U19488 (N_19488,N_17492,N_17095);
xor U19489 (N_19489,N_16191,N_16167);
nand U19490 (N_19490,N_16790,N_16705);
nand U19491 (N_19491,N_16973,N_16052);
or U19492 (N_19492,N_16821,N_17881);
xnor U19493 (N_19493,N_17552,N_17627);
or U19494 (N_19494,N_16370,N_16865);
xnor U19495 (N_19495,N_16086,N_17963);
nor U19496 (N_19496,N_17852,N_17180);
and U19497 (N_19497,N_17882,N_17272);
xnor U19498 (N_19498,N_17607,N_16773);
and U19499 (N_19499,N_17032,N_17610);
nor U19500 (N_19500,N_17306,N_17168);
xor U19501 (N_19501,N_16728,N_16425);
and U19502 (N_19502,N_16145,N_17919);
and U19503 (N_19503,N_16220,N_16400);
or U19504 (N_19504,N_17674,N_16775);
nor U19505 (N_19505,N_17029,N_16722);
nor U19506 (N_19506,N_16686,N_16610);
xor U19507 (N_19507,N_16107,N_17192);
nor U19508 (N_19508,N_17368,N_16263);
xor U19509 (N_19509,N_17493,N_17688);
or U19510 (N_19510,N_17376,N_17952);
nor U19511 (N_19511,N_17557,N_16441);
xor U19512 (N_19512,N_16566,N_16794);
nor U19513 (N_19513,N_16245,N_17081);
and U19514 (N_19514,N_17002,N_16737);
nor U19515 (N_19515,N_17059,N_17691);
nor U19516 (N_19516,N_17443,N_17295);
xor U19517 (N_19517,N_17530,N_17323);
nor U19518 (N_19518,N_17082,N_17331);
nor U19519 (N_19519,N_17661,N_16745);
or U19520 (N_19520,N_17622,N_17746);
nor U19521 (N_19521,N_17861,N_17265);
and U19522 (N_19522,N_17043,N_17013);
xor U19523 (N_19523,N_17418,N_17601);
nand U19524 (N_19524,N_17606,N_16839);
nor U19525 (N_19525,N_16986,N_17081);
and U19526 (N_19526,N_16508,N_17659);
and U19527 (N_19527,N_17281,N_17006);
or U19528 (N_19528,N_16632,N_17470);
or U19529 (N_19529,N_16403,N_17618);
and U19530 (N_19530,N_17469,N_17438);
nand U19531 (N_19531,N_16585,N_17691);
and U19532 (N_19532,N_16350,N_17851);
nand U19533 (N_19533,N_16483,N_16999);
and U19534 (N_19534,N_17497,N_16394);
or U19535 (N_19535,N_17480,N_16161);
and U19536 (N_19536,N_16447,N_17463);
xor U19537 (N_19537,N_17106,N_16804);
and U19538 (N_19538,N_16516,N_17010);
nor U19539 (N_19539,N_16525,N_17393);
or U19540 (N_19540,N_16871,N_16706);
and U19541 (N_19541,N_17655,N_17939);
and U19542 (N_19542,N_17450,N_17702);
nor U19543 (N_19543,N_17321,N_16095);
nand U19544 (N_19544,N_17744,N_17128);
xnor U19545 (N_19545,N_17993,N_16559);
nor U19546 (N_19546,N_16213,N_17475);
and U19547 (N_19547,N_17733,N_17662);
nor U19548 (N_19548,N_16673,N_17640);
nor U19549 (N_19549,N_17878,N_16368);
and U19550 (N_19550,N_16765,N_16955);
nand U19551 (N_19551,N_16602,N_16183);
and U19552 (N_19552,N_16214,N_16357);
nor U19553 (N_19553,N_17146,N_17916);
xor U19554 (N_19554,N_16578,N_16708);
or U19555 (N_19555,N_17502,N_16843);
and U19556 (N_19556,N_17916,N_17991);
or U19557 (N_19557,N_16736,N_17669);
nand U19558 (N_19558,N_16698,N_17477);
or U19559 (N_19559,N_17402,N_16948);
and U19560 (N_19560,N_16074,N_16814);
nand U19561 (N_19561,N_17377,N_17068);
or U19562 (N_19562,N_17657,N_16944);
nand U19563 (N_19563,N_17068,N_16387);
xor U19564 (N_19564,N_17357,N_17262);
and U19565 (N_19565,N_16639,N_17680);
xnor U19566 (N_19566,N_17090,N_17403);
and U19567 (N_19567,N_16533,N_17663);
xnor U19568 (N_19568,N_17298,N_17653);
xor U19569 (N_19569,N_16508,N_16099);
and U19570 (N_19570,N_17006,N_16528);
or U19571 (N_19571,N_17472,N_16821);
nor U19572 (N_19572,N_16185,N_17132);
nor U19573 (N_19573,N_16478,N_16953);
or U19574 (N_19574,N_16980,N_17431);
xor U19575 (N_19575,N_17164,N_16326);
and U19576 (N_19576,N_17416,N_16050);
or U19577 (N_19577,N_16528,N_17708);
or U19578 (N_19578,N_17174,N_17826);
xnor U19579 (N_19579,N_16611,N_17694);
and U19580 (N_19580,N_17693,N_17245);
and U19581 (N_19581,N_17674,N_17305);
nor U19582 (N_19582,N_16463,N_16108);
nand U19583 (N_19583,N_16360,N_17831);
xor U19584 (N_19584,N_17818,N_16092);
or U19585 (N_19585,N_16682,N_16777);
or U19586 (N_19586,N_16202,N_16120);
and U19587 (N_19587,N_17197,N_17917);
and U19588 (N_19588,N_16181,N_16715);
xnor U19589 (N_19589,N_17555,N_17421);
xnor U19590 (N_19590,N_16749,N_17748);
xor U19591 (N_19591,N_17821,N_16601);
nor U19592 (N_19592,N_17437,N_16762);
and U19593 (N_19593,N_17386,N_17545);
xor U19594 (N_19594,N_16606,N_17282);
xor U19595 (N_19595,N_16324,N_17426);
nand U19596 (N_19596,N_17781,N_16893);
or U19597 (N_19597,N_17724,N_17060);
xor U19598 (N_19598,N_17694,N_17510);
nor U19599 (N_19599,N_17529,N_16819);
nand U19600 (N_19600,N_16257,N_16759);
xnor U19601 (N_19601,N_17022,N_17690);
nand U19602 (N_19602,N_16223,N_16837);
or U19603 (N_19603,N_17038,N_17010);
nand U19604 (N_19604,N_17625,N_16336);
nand U19605 (N_19605,N_17105,N_16087);
or U19606 (N_19606,N_17624,N_16548);
or U19607 (N_19607,N_16952,N_17037);
xor U19608 (N_19608,N_17274,N_16366);
nor U19609 (N_19609,N_17677,N_17900);
nand U19610 (N_19610,N_16931,N_16090);
nand U19611 (N_19611,N_17422,N_16446);
or U19612 (N_19612,N_16879,N_16355);
nor U19613 (N_19613,N_17061,N_17133);
and U19614 (N_19614,N_17037,N_17848);
and U19615 (N_19615,N_16662,N_16585);
and U19616 (N_19616,N_17992,N_16533);
nand U19617 (N_19617,N_17637,N_16570);
xnor U19618 (N_19618,N_17950,N_16751);
and U19619 (N_19619,N_16867,N_17632);
and U19620 (N_19620,N_17522,N_17703);
xnor U19621 (N_19621,N_17323,N_17324);
xor U19622 (N_19622,N_16696,N_16841);
nand U19623 (N_19623,N_17803,N_17700);
and U19624 (N_19624,N_16935,N_17799);
nand U19625 (N_19625,N_17649,N_16912);
xnor U19626 (N_19626,N_16912,N_17861);
xor U19627 (N_19627,N_16976,N_17768);
xnor U19628 (N_19628,N_16826,N_16053);
xnor U19629 (N_19629,N_17004,N_17436);
or U19630 (N_19630,N_16924,N_17632);
or U19631 (N_19631,N_16293,N_17484);
nand U19632 (N_19632,N_16022,N_16475);
and U19633 (N_19633,N_16551,N_16510);
nand U19634 (N_19634,N_17542,N_16143);
or U19635 (N_19635,N_16790,N_16418);
nand U19636 (N_19636,N_17291,N_17264);
nor U19637 (N_19637,N_16311,N_16850);
nand U19638 (N_19638,N_17019,N_16178);
and U19639 (N_19639,N_17114,N_16318);
nor U19640 (N_19640,N_16514,N_17140);
xnor U19641 (N_19641,N_16661,N_17981);
and U19642 (N_19642,N_16825,N_16129);
and U19643 (N_19643,N_16182,N_16822);
or U19644 (N_19644,N_16067,N_16500);
or U19645 (N_19645,N_16768,N_16457);
nand U19646 (N_19646,N_17568,N_16067);
xor U19647 (N_19647,N_16549,N_17941);
and U19648 (N_19648,N_16242,N_16110);
or U19649 (N_19649,N_17441,N_17459);
or U19650 (N_19650,N_16785,N_16833);
nand U19651 (N_19651,N_16819,N_16761);
and U19652 (N_19652,N_16832,N_16985);
nand U19653 (N_19653,N_17685,N_16335);
nand U19654 (N_19654,N_17331,N_17629);
nand U19655 (N_19655,N_17658,N_17705);
or U19656 (N_19656,N_17105,N_16940);
nor U19657 (N_19657,N_17861,N_17934);
or U19658 (N_19658,N_17869,N_16008);
or U19659 (N_19659,N_16385,N_17289);
or U19660 (N_19660,N_16723,N_17458);
nand U19661 (N_19661,N_16921,N_16576);
or U19662 (N_19662,N_16602,N_16430);
or U19663 (N_19663,N_16549,N_16453);
xnor U19664 (N_19664,N_16302,N_17817);
and U19665 (N_19665,N_17456,N_17777);
or U19666 (N_19666,N_16900,N_16160);
nand U19667 (N_19667,N_16825,N_17304);
xor U19668 (N_19668,N_16000,N_17575);
nor U19669 (N_19669,N_16288,N_16286);
xor U19670 (N_19670,N_17780,N_16761);
nor U19671 (N_19671,N_17130,N_17966);
nor U19672 (N_19672,N_16489,N_17297);
nor U19673 (N_19673,N_16308,N_16491);
xor U19674 (N_19674,N_16604,N_17158);
nor U19675 (N_19675,N_16170,N_16425);
xor U19676 (N_19676,N_16541,N_16657);
or U19677 (N_19677,N_16654,N_16275);
and U19678 (N_19678,N_16347,N_16410);
xnor U19679 (N_19679,N_16870,N_17539);
nand U19680 (N_19680,N_16919,N_16150);
or U19681 (N_19681,N_17166,N_17953);
xnor U19682 (N_19682,N_16175,N_17520);
nor U19683 (N_19683,N_16424,N_17204);
xor U19684 (N_19684,N_17729,N_17909);
or U19685 (N_19685,N_17049,N_16044);
nand U19686 (N_19686,N_16539,N_17737);
and U19687 (N_19687,N_16961,N_16835);
nand U19688 (N_19688,N_17945,N_16703);
or U19689 (N_19689,N_16512,N_16992);
nand U19690 (N_19690,N_17850,N_16046);
nand U19691 (N_19691,N_17840,N_16045);
nor U19692 (N_19692,N_17811,N_17723);
nor U19693 (N_19693,N_16234,N_16385);
nor U19694 (N_19694,N_17942,N_16647);
xor U19695 (N_19695,N_16981,N_17230);
nor U19696 (N_19696,N_17765,N_17995);
nand U19697 (N_19697,N_16858,N_16116);
xnor U19698 (N_19698,N_17281,N_16880);
and U19699 (N_19699,N_17050,N_16049);
or U19700 (N_19700,N_16417,N_16460);
xnor U19701 (N_19701,N_16676,N_17336);
nand U19702 (N_19702,N_17674,N_17052);
xor U19703 (N_19703,N_17130,N_17404);
nor U19704 (N_19704,N_16242,N_16459);
nor U19705 (N_19705,N_17894,N_17907);
or U19706 (N_19706,N_16744,N_17536);
nor U19707 (N_19707,N_16259,N_17205);
nand U19708 (N_19708,N_16526,N_16177);
nand U19709 (N_19709,N_17671,N_17733);
nand U19710 (N_19710,N_17552,N_17088);
or U19711 (N_19711,N_17183,N_16600);
xnor U19712 (N_19712,N_17596,N_17263);
xor U19713 (N_19713,N_16932,N_16553);
and U19714 (N_19714,N_16222,N_16243);
and U19715 (N_19715,N_17478,N_16561);
nor U19716 (N_19716,N_17510,N_16847);
xor U19717 (N_19717,N_17782,N_16527);
nor U19718 (N_19718,N_16066,N_16153);
and U19719 (N_19719,N_16969,N_17354);
nand U19720 (N_19720,N_17718,N_17018);
nor U19721 (N_19721,N_16599,N_16978);
nand U19722 (N_19722,N_17579,N_16235);
nand U19723 (N_19723,N_16088,N_16743);
xnor U19724 (N_19724,N_17670,N_17921);
xnor U19725 (N_19725,N_17939,N_16416);
nand U19726 (N_19726,N_17369,N_17453);
xor U19727 (N_19727,N_17867,N_16877);
nand U19728 (N_19728,N_16605,N_17031);
nor U19729 (N_19729,N_16466,N_16807);
nand U19730 (N_19730,N_17704,N_17196);
or U19731 (N_19731,N_17973,N_16466);
nand U19732 (N_19732,N_16008,N_17856);
nor U19733 (N_19733,N_17497,N_16535);
or U19734 (N_19734,N_16967,N_17705);
nand U19735 (N_19735,N_16477,N_17106);
nand U19736 (N_19736,N_17149,N_17880);
xor U19737 (N_19737,N_17364,N_16041);
and U19738 (N_19738,N_17616,N_17457);
xor U19739 (N_19739,N_17081,N_17326);
or U19740 (N_19740,N_16964,N_17983);
and U19741 (N_19741,N_17588,N_17221);
xnor U19742 (N_19742,N_17679,N_17673);
and U19743 (N_19743,N_16423,N_17012);
nand U19744 (N_19744,N_16163,N_17592);
nand U19745 (N_19745,N_17502,N_17731);
or U19746 (N_19746,N_16543,N_17101);
or U19747 (N_19747,N_17002,N_17350);
nand U19748 (N_19748,N_16377,N_17480);
nand U19749 (N_19749,N_16297,N_17725);
xor U19750 (N_19750,N_17764,N_17706);
and U19751 (N_19751,N_17055,N_16307);
and U19752 (N_19752,N_16511,N_17912);
xnor U19753 (N_19753,N_17278,N_17386);
xnor U19754 (N_19754,N_16177,N_17752);
and U19755 (N_19755,N_16105,N_17881);
nand U19756 (N_19756,N_17049,N_16265);
nor U19757 (N_19757,N_17073,N_16089);
nand U19758 (N_19758,N_16139,N_16503);
nand U19759 (N_19759,N_17818,N_17786);
or U19760 (N_19760,N_17700,N_16565);
xor U19761 (N_19761,N_17839,N_17323);
and U19762 (N_19762,N_16381,N_17915);
xnor U19763 (N_19763,N_17963,N_16597);
or U19764 (N_19764,N_17549,N_17732);
nor U19765 (N_19765,N_16644,N_17271);
nor U19766 (N_19766,N_16348,N_16111);
nor U19767 (N_19767,N_16472,N_16206);
or U19768 (N_19768,N_17804,N_16576);
nor U19769 (N_19769,N_17275,N_16558);
xnor U19770 (N_19770,N_17925,N_16507);
nor U19771 (N_19771,N_16397,N_17291);
and U19772 (N_19772,N_17435,N_17564);
xnor U19773 (N_19773,N_16615,N_16423);
nor U19774 (N_19774,N_16109,N_17824);
or U19775 (N_19775,N_16474,N_16348);
and U19776 (N_19776,N_17197,N_16906);
or U19777 (N_19777,N_16677,N_16128);
and U19778 (N_19778,N_17945,N_16021);
or U19779 (N_19779,N_16977,N_16571);
nand U19780 (N_19780,N_16135,N_16523);
nand U19781 (N_19781,N_16414,N_16667);
or U19782 (N_19782,N_17414,N_17895);
xor U19783 (N_19783,N_16545,N_17555);
or U19784 (N_19784,N_16356,N_16548);
and U19785 (N_19785,N_16457,N_16607);
and U19786 (N_19786,N_17265,N_16822);
xor U19787 (N_19787,N_17421,N_17047);
xnor U19788 (N_19788,N_16213,N_16079);
xor U19789 (N_19789,N_16561,N_16732);
and U19790 (N_19790,N_16815,N_16640);
nor U19791 (N_19791,N_17640,N_17516);
nor U19792 (N_19792,N_16704,N_17077);
and U19793 (N_19793,N_17364,N_16381);
or U19794 (N_19794,N_17338,N_17592);
or U19795 (N_19795,N_17171,N_16191);
nand U19796 (N_19796,N_17446,N_17193);
xnor U19797 (N_19797,N_16704,N_17053);
nand U19798 (N_19798,N_16229,N_17763);
xor U19799 (N_19799,N_17075,N_16039);
and U19800 (N_19800,N_17126,N_16169);
nand U19801 (N_19801,N_16704,N_16718);
xor U19802 (N_19802,N_17858,N_16357);
or U19803 (N_19803,N_16380,N_16131);
and U19804 (N_19804,N_16828,N_17450);
and U19805 (N_19805,N_17118,N_17700);
nor U19806 (N_19806,N_17710,N_17423);
xnor U19807 (N_19807,N_17524,N_16828);
xnor U19808 (N_19808,N_17581,N_16831);
xor U19809 (N_19809,N_17541,N_16829);
and U19810 (N_19810,N_17439,N_16897);
and U19811 (N_19811,N_16932,N_17841);
xor U19812 (N_19812,N_17377,N_17190);
and U19813 (N_19813,N_17238,N_16873);
nand U19814 (N_19814,N_16939,N_16398);
nand U19815 (N_19815,N_16614,N_17869);
nand U19816 (N_19816,N_16076,N_17622);
and U19817 (N_19817,N_17790,N_17175);
xnor U19818 (N_19818,N_16994,N_17497);
and U19819 (N_19819,N_17484,N_17949);
nand U19820 (N_19820,N_17657,N_16730);
nor U19821 (N_19821,N_17543,N_16428);
and U19822 (N_19822,N_16639,N_17774);
and U19823 (N_19823,N_16377,N_17588);
and U19824 (N_19824,N_17115,N_17207);
and U19825 (N_19825,N_17720,N_16302);
xor U19826 (N_19826,N_17322,N_16904);
or U19827 (N_19827,N_17859,N_17643);
and U19828 (N_19828,N_16272,N_17700);
nor U19829 (N_19829,N_16729,N_17157);
or U19830 (N_19830,N_17552,N_16883);
nor U19831 (N_19831,N_16289,N_17714);
xnor U19832 (N_19832,N_16439,N_16271);
nor U19833 (N_19833,N_17243,N_17129);
xnor U19834 (N_19834,N_17943,N_17904);
nor U19835 (N_19835,N_17002,N_17150);
and U19836 (N_19836,N_16087,N_17312);
and U19837 (N_19837,N_17355,N_16534);
or U19838 (N_19838,N_17901,N_17673);
and U19839 (N_19839,N_16584,N_16442);
nor U19840 (N_19840,N_17883,N_17713);
and U19841 (N_19841,N_16367,N_16094);
xor U19842 (N_19842,N_16106,N_17925);
and U19843 (N_19843,N_17592,N_17222);
nor U19844 (N_19844,N_16498,N_16394);
nor U19845 (N_19845,N_16737,N_17283);
nand U19846 (N_19846,N_17002,N_16874);
and U19847 (N_19847,N_17090,N_17852);
or U19848 (N_19848,N_16754,N_16714);
or U19849 (N_19849,N_17463,N_16378);
or U19850 (N_19850,N_17819,N_16882);
nor U19851 (N_19851,N_16447,N_17285);
or U19852 (N_19852,N_17540,N_17557);
xnor U19853 (N_19853,N_17751,N_16762);
xor U19854 (N_19854,N_17441,N_16277);
and U19855 (N_19855,N_17215,N_16365);
nand U19856 (N_19856,N_16497,N_17344);
or U19857 (N_19857,N_16515,N_17437);
or U19858 (N_19858,N_17800,N_16191);
nor U19859 (N_19859,N_16814,N_17636);
xor U19860 (N_19860,N_17961,N_17446);
nand U19861 (N_19861,N_16842,N_17098);
nor U19862 (N_19862,N_17417,N_16133);
nor U19863 (N_19863,N_17745,N_16437);
or U19864 (N_19864,N_16024,N_16521);
nor U19865 (N_19865,N_16094,N_17467);
or U19866 (N_19866,N_17438,N_17670);
nor U19867 (N_19867,N_17439,N_16571);
or U19868 (N_19868,N_16700,N_17518);
or U19869 (N_19869,N_17015,N_17692);
nor U19870 (N_19870,N_16204,N_16884);
xor U19871 (N_19871,N_17933,N_16499);
nand U19872 (N_19872,N_16544,N_17213);
nor U19873 (N_19873,N_17497,N_17929);
or U19874 (N_19874,N_17606,N_17455);
or U19875 (N_19875,N_16655,N_16966);
nand U19876 (N_19876,N_17099,N_16696);
or U19877 (N_19877,N_17209,N_16759);
xor U19878 (N_19878,N_17518,N_17351);
and U19879 (N_19879,N_17521,N_17289);
and U19880 (N_19880,N_16709,N_16668);
and U19881 (N_19881,N_16130,N_16037);
and U19882 (N_19882,N_16207,N_17465);
or U19883 (N_19883,N_16097,N_16928);
xnor U19884 (N_19884,N_17019,N_16895);
nor U19885 (N_19885,N_17348,N_17857);
nor U19886 (N_19886,N_17063,N_16824);
nor U19887 (N_19887,N_16822,N_16781);
and U19888 (N_19888,N_17766,N_17136);
nor U19889 (N_19889,N_17988,N_17337);
or U19890 (N_19890,N_17947,N_17938);
xor U19891 (N_19891,N_16510,N_17290);
or U19892 (N_19892,N_16782,N_17210);
xor U19893 (N_19893,N_17349,N_16255);
and U19894 (N_19894,N_17579,N_16318);
or U19895 (N_19895,N_17579,N_16154);
nand U19896 (N_19896,N_16487,N_16109);
and U19897 (N_19897,N_16520,N_17297);
nand U19898 (N_19898,N_16023,N_16062);
xnor U19899 (N_19899,N_17626,N_17930);
or U19900 (N_19900,N_16660,N_16692);
and U19901 (N_19901,N_16414,N_17991);
nor U19902 (N_19902,N_16518,N_17492);
and U19903 (N_19903,N_17400,N_17282);
or U19904 (N_19904,N_17652,N_16503);
or U19905 (N_19905,N_16402,N_16182);
and U19906 (N_19906,N_17464,N_16605);
xor U19907 (N_19907,N_16227,N_16524);
or U19908 (N_19908,N_17288,N_17684);
or U19909 (N_19909,N_17089,N_16371);
nand U19910 (N_19910,N_17080,N_17668);
and U19911 (N_19911,N_16010,N_16776);
or U19912 (N_19912,N_16444,N_17016);
or U19913 (N_19913,N_17642,N_17488);
nand U19914 (N_19914,N_17568,N_16931);
xor U19915 (N_19915,N_16272,N_17064);
nor U19916 (N_19916,N_16795,N_17999);
xor U19917 (N_19917,N_16852,N_16475);
and U19918 (N_19918,N_17619,N_17598);
nand U19919 (N_19919,N_17942,N_17902);
nand U19920 (N_19920,N_16302,N_17154);
nor U19921 (N_19921,N_16614,N_17087);
nor U19922 (N_19922,N_17090,N_16131);
nor U19923 (N_19923,N_17621,N_16474);
nand U19924 (N_19924,N_16642,N_16552);
or U19925 (N_19925,N_16521,N_17000);
xor U19926 (N_19926,N_17829,N_16989);
and U19927 (N_19927,N_17749,N_16600);
nor U19928 (N_19928,N_16054,N_16337);
and U19929 (N_19929,N_16003,N_17093);
and U19930 (N_19930,N_17735,N_17442);
nand U19931 (N_19931,N_16243,N_17248);
nor U19932 (N_19932,N_16601,N_16881);
xor U19933 (N_19933,N_17077,N_17051);
nand U19934 (N_19934,N_17538,N_17516);
and U19935 (N_19935,N_17103,N_16836);
or U19936 (N_19936,N_16660,N_16011);
and U19937 (N_19937,N_17960,N_16369);
nor U19938 (N_19938,N_17198,N_17954);
xor U19939 (N_19939,N_17488,N_16394);
nor U19940 (N_19940,N_17859,N_16179);
or U19941 (N_19941,N_17003,N_16088);
and U19942 (N_19942,N_17506,N_17835);
or U19943 (N_19943,N_17018,N_17404);
nand U19944 (N_19944,N_16135,N_16889);
xor U19945 (N_19945,N_16528,N_16194);
xnor U19946 (N_19946,N_16176,N_16105);
nand U19947 (N_19947,N_17346,N_17715);
xnor U19948 (N_19948,N_17390,N_17130);
nor U19949 (N_19949,N_16454,N_17465);
nand U19950 (N_19950,N_16814,N_17095);
or U19951 (N_19951,N_17784,N_16468);
and U19952 (N_19952,N_17645,N_17943);
nand U19953 (N_19953,N_17534,N_17171);
nor U19954 (N_19954,N_16376,N_16975);
nor U19955 (N_19955,N_16247,N_16463);
nand U19956 (N_19956,N_17596,N_17133);
nand U19957 (N_19957,N_16984,N_16038);
or U19958 (N_19958,N_17055,N_16433);
and U19959 (N_19959,N_17518,N_17627);
nand U19960 (N_19960,N_16577,N_16175);
and U19961 (N_19961,N_16799,N_16089);
xor U19962 (N_19962,N_17446,N_17962);
or U19963 (N_19963,N_17539,N_17736);
nand U19964 (N_19964,N_17906,N_16676);
or U19965 (N_19965,N_17217,N_16785);
nor U19966 (N_19966,N_16576,N_17552);
xnor U19967 (N_19967,N_17111,N_17001);
and U19968 (N_19968,N_16544,N_17055);
or U19969 (N_19969,N_17163,N_17549);
or U19970 (N_19970,N_17060,N_17912);
nand U19971 (N_19971,N_17742,N_17151);
nor U19972 (N_19972,N_17236,N_17630);
xor U19973 (N_19973,N_17745,N_17249);
and U19974 (N_19974,N_16546,N_16207);
and U19975 (N_19975,N_17454,N_17876);
and U19976 (N_19976,N_17789,N_16692);
nand U19977 (N_19977,N_17801,N_16047);
and U19978 (N_19978,N_17227,N_16884);
and U19979 (N_19979,N_17282,N_16368);
and U19980 (N_19980,N_16941,N_16251);
nor U19981 (N_19981,N_17855,N_17476);
xnor U19982 (N_19982,N_16231,N_16053);
xor U19983 (N_19983,N_17986,N_17783);
xnor U19984 (N_19984,N_16045,N_16593);
xnor U19985 (N_19985,N_16681,N_16245);
xor U19986 (N_19986,N_16179,N_17889);
xnor U19987 (N_19987,N_17568,N_16510);
and U19988 (N_19988,N_17826,N_16076);
nor U19989 (N_19989,N_17160,N_16606);
nand U19990 (N_19990,N_16709,N_17613);
or U19991 (N_19991,N_17396,N_16303);
nand U19992 (N_19992,N_16703,N_16182);
or U19993 (N_19993,N_17461,N_16391);
nand U19994 (N_19994,N_16233,N_16611);
or U19995 (N_19995,N_17737,N_17979);
and U19996 (N_19996,N_17247,N_16191);
and U19997 (N_19997,N_16049,N_16636);
or U19998 (N_19998,N_16925,N_17763);
xnor U19999 (N_19999,N_17554,N_17766);
and UO_0 (O_0,N_18551,N_18176);
nor UO_1 (O_1,N_18914,N_19734);
xnor UO_2 (O_2,N_18869,N_18406);
and UO_3 (O_3,N_18634,N_19532);
and UO_4 (O_4,N_18941,N_18938);
xor UO_5 (O_5,N_19741,N_18433);
and UO_6 (O_6,N_19529,N_19425);
nor UO_7 (O_7,N_19203,N_18726);
xnor UO_8 (O_8,N_18244,N_19449);
and UO_9 (O_9,N_18959,N_19353);
nand UO_10 (O_10,N_19910,N_19962);
nand UO_11 (O_11,N_18876,N_19816);
nor UO_12 (O_12,N_19326,N_18628);
nor UO_13 (O_13,N_18654,N_18723);
and UO_14 (O_14,N_19728,N_19123);
nor UO_15 (O_15,N_18684,N_18187);
nor UO_16 (O_16,N_18161,N_18750);
nand UO_17 (O_17,N_19506,N_19496);
and UO_18 (O_18,N_18758,N_18565);
and UO_19 (O_19,N_19813,N_19551);
nand UO_20 (O_20,N_18698,N_18686);
nor UO_21 (O_21,N_18219,N_18868);
or UO_22 (O_22,N_18909,N_18663);
xor UO_23 (O_23,N_19825,N_18745);
nor UO_24 (O_24,N_18969,N_18353);
nor UO_25 (O_25,N_19137,N_18798);
xor UO_26 (O_26,N_19034,N_18140);
and UO_27 (O_27,N_18057,N_18871);
or UO_28 (O_28,N_18437,N_18232);
or UO_29 (O_29,N_19987,N_19254);
nand UO_30 (O_30,N_18248,N_18329);
and UO_31 (O_31,N_19947,N_18385);
and UO_32 (O_32,N_18811,N_18442);
nor UO_33 (O_33,N_18369,N_19598);
nor UO_34 (O_34,N_19671,N_19427);
nand UO_35 (O_35,N_19836,N_18711);
and UO_36 (O_36,N_19380,N_19284);
and UO_37 (O_37,N_18229,N_19858);
or UO_38 (O_38,N_19490,N_19870);
nor UO_39 (O_39,N_19038,N_18878);
nor UO_40 (O_40,N_19046,N_18364);
xor UO_41 (O_41,N_18728,N_19324);
nor UO_42 (O_42,N_18131,N_19125);
nor UO_43 (O_43,N_19132,N_18933);
and UO_44 (O_44,N_19941,N_18597);
nand UO_45 (O_45,N_18481,N_18655);
xnor UO_46 (O_46,N_19288,N_18886);
nand UO_47 (O_47,N_18340,N_18271);
nand UO_48 (O_48,N_18472,N_18827);
and UO_49 (O_49,N_19452,N_18840);
or UO_50 (O_50,N_18790,N_18136);
and UO_51 (O_51,N_19537,N_18756);
nor UO_52 (O_52,N_19637,N_19155);
xor UO_53 (O_53,N_18260,N_18712);
or UO_54 (O_54,N_19863,N_19851);
xnor UO_55 (O_55,N_18036,N_19662);
or UO_56 (O_56,N_19442,N_18135);
and UO_57 (O_57,N_18138,N_19811);
nand UO_58 (O_58,N_19277,N_18178);
nor UO_59 (O_59,N_19651,N_18095);
or UO_60 (O_60,N_19607,N_19860);
or UO_61 (O_61,N_18861,N_18570);
nand UO_62 (O_62,N_18793,N_19828);
xnor UO_63 (O_63,N_18245,N_18425);
xor UO_64 (O_64,N_19902,N_19823);
nor UO_65 (O_65,N_19698,N_19697);
nand UO_66 (O_66,N_18530,N_19877);
xor UO_67 (O_67,N_18328,N_19437);
nor UO_68 (O_68,N_19867,N_18865);
or UO_69 (O_69,N_19041,N_19348);
nor UO_70 (O_70,N_19781,N_19623);
and UO_71 (O_71,N_19318,N_18851);
or UO_72 (O_72,N_18124,N_18262);
and UO_73 (O_73,N_19293,N_18848);
or UO_74 (O_74,N_18916,N_19417);
nand UO_75 (O_75,N_18638,N_18584);
nor UO_76 (O_76,N_19934,N_18403);
or UO_77 (O_77,N_18130,N_18942);
nor UO_78 (O_78,N_18574,N_18267);
or UO_79 (O_79,N_19766,N_19684);
or UO_80 (O_80,N_18335,N_18354);
nor UO_81 (O_81,N_18247,N_18699);
nand UO_82 (O_82,N_19821,N_19120);
nor UO_83 (O_83,N_18533,N_18467);
and UO_84 (O_84,N_19289,N_18429);
and UO_85 (O_85,N_18853,N_19161);
or UO_86 (O_86,N_19482,N_19719);
and UO_87 (O_87,N_18413,N_19475);
xor UO_88 (O_88,N_19259,N_18208);
nand UO_89 (O_89,N_18078,N_18133);
nor UO_90 (O_90,N_18559,N_18754);
nand UO_91 (O_91,N_18116,N_18822);
and UO_92 (O_92,N_19384,N_19977);
xor UO_93 (O_93,N_19635,N_18650);
xnor UO_94 (O_94,N_18908,N_18348);
and UO_95 (O_95,N_19398,N_18360);
or UO_96 (O_96,N_19503,N_19233);
nor UO_97 (O_97,N_19704,N_19007);
nand UO_98 (O_98,N_19378,N_19024);
and UO_99 (O_99,N_18681,N_19830);
nor UO_100 (O_100,N_18872,N_18150);
nand UO_101 (O_101,N_18257,N_19750);
xnor UO_102 (O_102,N_18334,N_19481);
nor UO_103 (O_103,N_19622,N_19979);
and UO_104 (O_104,N_19385,N_19356);
nand UO_105 (O_105,N_18749,N_18004);
xor UO_106 (O_106,N_19916,N_18186);
nor UO_107 (O_107,N_18311,N_18603);
and UO_108 (O_108,N_19394,N_18833);
or UO_109 (O_109,N_19911,N_19748);
or UO_110 (O_110,N_18153,N_18605);
nor UO_111 (O_111,N_19957,N_18881);
xor UO_112 (O_112,N_18981,N_19265);
and UO_113 (O_113,N_18240,N_19773);
or UO_114 (O_114,N_18202,N_18185);
nor UO_115 (O_115,N_19932,N_18904);
and UO_116 (O_116,N_18792,N_18852);
nor UO_117 (O_117,N_18322,N_18234);
nor UO_118 (O_118,N_18616,N_18256);
nand UO_119 (O_119,N_18787,N_18645);
xnor UO_120 (O_120,N_18893,N_19817);
and UO_121 (O_121,N_19371,N_18714);
nor UO_122 (O_122,N_18776,N_19925);
xor UO_123 (O_123,N_18387,N_19804);
or UO_124 (O_124,N_18007,N_18103);
and UO_125 (O_125,N_19843,N_18330);
nor UO_126 (O_126,N_18374,N_19098);
nor UO_127 (O_127,N_18884,N_19679);
nand UO_128 (O_128,N_18527,N_19168);
nand UO_129 (O_129,N_18390,N_19295);
and UO_130 (O_130,N_19292,N_19924);
and UO_131 (O_131,N_18098,N_18225);
nand UO_132 (O_132,N_19997,N_18464);
and UO_133 (O_133,N_19862,N_18094);
nand UO_134 (O_134,N_18180,N_19221);
nand UO_135 (O_135,N_18174,N_19114);
nor UO_136 (O_136,N_18294,N_19527);
nor UO_137 (O_137,N_18082,N_18598);
nand UO_138 (O_138,N_18773,N_19919);
nand UO_139 (O_139,N_19775,N_19239);
and UO_140 (O_140,N_18236,N_18190);
and UO_141 (O_141,N_18469,N_19770);
xnor UO_142 (O_142,N_18394,N_18155);
or UO_143 (O_143,N_19524,N_18503);
nand UO_144 (O_144,N_19177,N_19632);
and UO_145 (O_145,N_19247,N_19146);
nand UO_146 (O_146,N_19140,N_19727);
and UO_147 (O_147,N_18775,N_18146);
nor UO_148 (O_148,N_19810,N_19470);
nor UO_149 (O_149,N_18285,N_19197);
nand UO_150 (O_150,N_19900,N_19584);
and UO_151 (O_151,N_19269,N_19065);
and UO_152 (O_152,N_19777,N_19627);
or UO_153 (O_153,N_18371,N_19274);
and UO_154 (O_154,N_18310,N_18492);
nor UO_155 (O_155,N_18372,N_19762);
nor UO_156 (O_156,N_18218,N_19225);
xnor UO_157 (O_157,N_19476,N_18621);
xnor UO_158 (O_158,N_18170,N_19213);
and UO_159 (O_159,N_19631,N_19642);
nand UO_160 (O_160,N_18383,N_18120);
and UO_161 (O_161,N_19141,N_19946);
nor UO_162 (O_162,N_19788,N_19959);
and UO_163 (O_163,N_18960,N_18418);
and UO_164 (O_164,N_19515,N_18434);
and UO_165 (O_165,N_18898,N_18831);
and UO_166 (O_166,N_19691,N_18156);
nand UO_167 (O_167,N_18906,N_18541);
and UO_168 (O_168,N_19783,N_19854);
nand UO_169 (O_169,N_18587,N_18777);
nor UO_170 (O_170,N_19174,N_18314);
nor UO_171 (O_171,N_18580,N_18629);
nor UO_172 (O_172,N_18599,N_18099);
nor UO_173 (O_173,N_18378,N_18733);
and UO_174 (O_174,N_19388,N_19036);
nand UO_175 (O_175,N_18556,N_18992);
nor UO_176 (O_176,N_18063,N_18062);
or UO_177 (O_177,N_19207,N_19159);
or UO_178 (O_178,N_18452,N_18891);
or UO_179 (O_179,N_19364,N_18582);
nand UO_180 (O_180,N_18676,N_19311);
nor UO_181 (O_181,N_19409,N_18615);
or UO_182 (O_182,N_18357,N_18991);
nor UO_183 (O_183,N_19771,N_18243);
xnor UO_184 (O_184,N_19117,N_19373);
nand UO_185 (O_185,N_19226,N_19696);
nand UO_186 (O_186,N_19250,N_18934);
nand UO_187 (O_187,N_19834,N_18944);
xnor UO_188 (O_188,N_19855,N_19536);
nand UO_189 (O_189,N_18496,N_19614);
nand UO_190 (O_190,N_19395,N_19915);
xnor UO_191 (O_191,N_19595,N_19359);
xnor UO_192 (O_192,N_18043,N_18930);
nand UO_193 (O_193,N_18892,N_18367);
xnor UO_194 (O_194,N_19908,N_18212);
nand UO_195 (O_195,N_19624,N_19907);
nand UO_196 (O_196,N_19521,N_19342);
xor UO_197 (O_197,N_18689,N_19228);
and UO_198 (O_198,N_19070,N_18671);
xor UO_199 (O_199,N_19838,N_19018);
or UO_200 (O_200,N_19878,N_19063);
and UO_201 (O_201,N_19302,N_19673);
nor UO_202 (O_202,N_18744,N_18823);
nor UO_203 (O_203,N_18123,N_19795);
xnor UO_204 (O_204,N_18552,N_18015);
and UO_205 (O_205,N_18896,N_19211);
or UO_206 (O_206,N_19413,N_18854);
xor UO_207 (O_207,N_18951,N_19666);
nor UO_208 (O_208,N_18788,N_18962);
nor UO_209 (O_209,N_19438,N_19291);
xor UO_210 (O_210,N_19803,N_19998);
nor UO_211 (O_211,N_18973,N_18618);
xor UO_212 (O_212,N_18297,N_19973);
xor UO_213 (O_213,N_18384,N_18067);
or UO_214 (O_214,N_18569,N_18303);
nand UO_215 (O_215,N_19661,N_18313);
or UO_216 (O_216,N_18048,N_18058);
and UO_217 (O_217,N_19343,N_19154);
nand UO_218 (O_218,N_19191,N_19706);
or UO_219 (O_219,N_18477,N_19261);
nor UO_220 (O_220,N_19577,N_18769);
xnor UO_221 (O_221,N_19656,N_19848);
or UO_222 (O_222,N_19352,N_19334);
xor UO_223 (O_223,N_19866,N_18958);
nand UO_224 (O_224,N_18915,N_18149);
and UO_225 (O_225,N_19149,N_19921);
or UO_226 (O_226,N_18729,N_19365);
and UO_227 (O_227,N_18619,N_19004);
nor UO_228 (O_228,N_18517,N_18889);
nor UO_229 (O_229,N_19682,N_18538);
and UO_230 (O_230,N_18268,N_19057);
xor UO_231 (O_231,N_18590,N_18986);
nor UO_232 (O_232,N_19178,N_19309);
xor UO_233 (O_233,N_18596,N_19319);
and UO_234 (O_234,N_18639,N_18836);
xnor UO_235 (O_235,N_18691,N_18101);
nand UO_236 (O_236,N_18209,N_19489);
xnor UO_237 (O_237,N_19504,N_18781);
and UO_238 (O_238,N_19290,N_18441);
and UO_239 (O_239,N_18030,N_18059);
and UO_240 (O_240,N_19280,N_19712);
nor UO_241 (O_241,N_19093,N_19849);
nand UO_242 (O_242,N_19346,N_19760);
nor UO_243 (O_243,N_18122,N_19165);
nor UO_244 (O_244,N_18046,N_19659);
nor UO_245 (O_245,N_19549,N_18325);
nor UO_246 (O_246,N_19794,N_18679);
and UO_247 (O_247,N_19738,N_18727);
xnor UO_248 (O_248,N_19067,N_18796);
and UO_249 (O_249,N_19031,N_18768);
nand UO_250 (O_250,N_19565,N_18341);
and UO_251 (O_251,N_18839,N_18657);
nand UO_252 (O_252,N_18502,N_18771);
nand UO_253 (O_253,N_19264,N_19091);
nand UO_254 (O_254,N_18537,N_19074);
nand UO_255 (O_255,N_19006,N_19769);
or UO_256 (O_256,N_19135,N_19485);
or UO_257 (O_257,N_18976,N_19235);
and UO_258 (O_258,N_19298,N_18778);
nor UO_259 (O_259,N_18395,N_19391);
nor UO_260 (O_260,N_19757,N_18897);
or UO_261 (O_261,N_18662,N_19049);
and UO_262 (O_262,N_19538,N_19231);
and UO_263 (O_263,N_18952,N_19325);
nand UO_264 (O_264,N_18824,N_19208);
or UO_265 (O_265,N_19895,N_19668);
or UO_266 (O_266,N_18143,N_18794);
xor UO_267 (O_267,N_19732,N_18774);
nor UO_268 (O_268,N_18068,N_18820);
nand UO_269 (O_269,N_19652,N_18215);
xor UO_270 (O_270,N_18801,N_19369);
nor UO_271 (O_271,N_19639,N_19791);
xnor UO_272 (O_272,N_19405,N_19820);
and UO_273 (O_273,N_19890,N_19965);
nor UO_274 (O_274,N_19188,N_19865);
nand UO_275 (O_275,N_19003,N_18242);
or UO_276 (O_276,N_19301,N_18443);
and UO_277 (O_277,N_19955,N_19570);
nand UO_278 (O_278,N_19847,N_18031);
nand UO_279 (O_279,N_18214,N_18119);
nand UO_280 (O_280,N_19575,N_18841);
nand UO_281 (O_281,N_19990,N_19107);
nor UO_282 (O_282,N_19985,N_19456);
nand UO_283 (O_283,N_19993,N_18431);
or UO_284 (O_284,N_18375,N_18762);
nor UO_285 (O_285,N_19060,N_18859);
nand UO_286 (O_286,N_19724,N_18857);
xnor UO_287 (O_287,N_19156,N_19960);
nor UO_288 (O_288,N_19009,N_18018);
xor UO_289 (O_289,N_19025,N_18049);
nor UO_290 (O_290,N_18830,N_18928);
nor UO_291 (O_291,N_19045,N_18069);
or UO_292 (O_292,N_18002,N_18542);
xnor UO_293 (O_293,N_18770,N_18377);
or UO_294 (O_294,N_19106,N_19884);
nand UO_295 (O_295,N_19448,N_19224);
and UO_296 (O_296,N_18578,N_19234);
nor UO_297 (O_297,N_18498,N_19660);
nor UO_298 (O_298,N_19210,N_19829);
xor UO_299 (O_299,N_19628,N_19227);
or UO_300 (O_300,N_19143,N_19818);
and UO_301 (O_301,N_18401,N_19643);
nand UO_302 (O_302,N_19667,N_18845);
or UO_303 (O_303,N_18937,N_19824);
xor UO_304 (O_304,N_19723,N_18804);
or UO_305 (O_305,N_19392,N_19455);
nor UO_306 (O_306,N_19048,N_18494);
nor UO_307 (O_307,N_19037,N_18905);
nand UO_308 (O_308,N_18090,N_19753);
xor UO_309 (O_309,N_18412,N_18465);
and UO_310 (O_310,N_19459,N_18998);
or UO_311 (O_311,N_18550,N_19505);
or UO_312 (O_312,N_19896,N_18461);
nor UO_313 (O_313,N_19541,N_19731);
xnor UO_314 (O_314,N_18995,N_18152);
xnor UO_315 (O_315,N_18291,N_19053);
xor UO_316 (O_316,N_19021,N_19307);
nor UO_317 (O_317,N_19814,N_18344);
and UO_318 (O_318,N_18713,N_18764);
and UO_319 (O_319,N_18665,N_18748);
nand UO_320 (O_320,N_18368,N_18490);
nor UO_321 (O_321,N_19026,N_18978);
xnor UO_322 (O_322,N_18519,N_19717);
or UO_323 (O_323,N_19263,N_19194);
and UO_324 (O_324,N_18718,N_19815);
nor UO_325 (O_325,N_18040,N_18253);
and UO_326 (O_326,N_19948,N_19591);
nand UO_327 (O_327,N_19699,N_18339);
xnor UO_328 (O_328,N_19216,N_18731);
and UO_329 (O_329,N_19601,N_19118);
xor UO_330 (O_330,N_18188,N_19271);
nand UO_331 (O_331,N_18264,N_19871);
xnor UO_332 (O_332,N_19418,N_19440);
xnor UO_333 (O_333,N_19454,N_19267);
nor UO_334 (O_334,N_18561,N_19430);
xnor UO_335 (O_335,N_18485,N_19972);
xnor UO_336 (O_336,N_18860,N_18070);
xor UO_337 (O_337,N_19488,N_19412);
or UO_338 (O_338,N_18927,N_19509);
and UO_339 (O_339,N_18436,N_19519);
xnor UO_340 (O_340,N_19126,N_18290);
nor UO_341 (O_341,N_19381,N_19872);
nor UO_342 (O_342,N_19322,N_19163);
xor UO_343 (O_343,N_19054,N_18419);
nand UO_344 (O_344,N_19525,N_18555);
and UO_345 (O_345,N_19205,N_18834);
and UO_346 (O_346,N_18534,N_19615);
or UO_347 (O_347,N_18623,N_19655);
or UO_348 (O_348,N_18486,N_19966);
and UO_349 (O_349,N_18947,N_19103);
nor UO_350 (O_350,N_18125,N_18147);
or UO_351 (O_351,N_19500,N_19879);
nand UO_352 (O_352,N_18200,N_18614);
or UO_353 (O_353,N_18308,N_18641);
xnor UO_354 (O_354,N_18193,N_18276);
nand UO_355 (O_355,N_19995,N_18342);
nand UO_356 (O_356,N_18987,N_18967);
xnor UO_357 (O_357,N_19569,N_18604);
nor UO_358 (O_358,N_19217,N_19222);
nand UO_359 (O_359,N_18332,N_19257);
and UO_360 (O_360,N_19784,N_19200);
nand UO_361 (O_361,N_18279,N_18021);
or UO_362 (O_362,N_18025,N_18595);
or UO_363 (O_363,N_19789,N_18482);
nand UO_364 (O_364,N_19526,N_19469);
nor UO_365 (O_365,N_18894,N_19169);
nand UO_366 (O_366,N_19733,N_18805);
xor UO_367 (O_367,N_18782,N_18213);
nor UO_368 (O_368,N_19432,N_18447);
nand UO_369 (O_369,N_19183,N_18563);
nand UO_370 (O_370,N_19081,N_18270);
xnor UO_371 (O_371,N_18880,N_19323);
or UO_372 (O_372,N_19885,N_19453);
and UO_373 (O_373,N_19061,N_18050);
nand UO_374 (O_374,N_19328,N_18703);
and UO_375 (O_375,N_19142,N_19550);
xnor UO_376 (O_376,N_19131,N_19279);
or UO_377 (O_377,N_19912,N_18807);
nor UO_378 (O_378,N_18522,N_18115);
or UO_379 (O_379,N_18284,N_19287);
nor UO_380 (O_380,N_18283,N_19138);
and UO_381 (O_381,N_18439,N_18331);
xor UO_382 (O_382,N_18814,N_19320);
and UO_383 (O_383,N_18012,N_18266);
nor UO_384 (O_384,N_19032,N_18539);
or UO_385 (O_385,N_18510,N_19097);
nand UO_386 (O_386,N_19076,N_19458);
nand UO_387 (O_387,N_19968,N_19883);
or UO_388 (O_388,N_19914,N_19576);
and UO_389 (O_389,N_18014,N_19176);
and UO_390 (O_390,N_19088,N_19075);
or UO_391 (O_391,N_18725,N_19001);
nor UO_392 (O_392,N_18620,N_18631);
nor UO_393 (O_393,N_18760,N_19180);
and UO_394 (O_394,N_19787,N_19875);
nor UO_395 (O_395,N_19446,N_19195);
nand UO_396 (O_396,N_18409,N_18356);
nand UO_397 (O_397,N_19214,N_19134);
nor UO_398 (O_398,N_18196,N_19558);
nor UO_399 (O_399,N_18935,N_19079);
and UO_400 (O_400,N_19510,N_18414);
and UO_401 (O_401,N_19242,N_18763);
nand UO_402 (O_402,N_18277,N_19206);
nor UO_403 (O_403,N_19282,N_19013);
nand UO_404 (O_404,N_18104,N_19219);
nor UO_405 (O_405,N_18626,N_18081);
and UO_406 (O_406,N_18060,N_19597);
xor UO_407 (O_407,N_19636,N_19864);
nor UO_408 (O_408,N_19403,N_19028);
xnor UO_409 (O_409,N_18767,N_18653);
nor UO_410 (O_410,N_18269,N_19850);
xor UO_411 (O_411,N_18226,N_18887);
or UO_412 (O_412,N_19019,N_18061);
or UO_413 (O_413,N_18903,N_18716);
nor UO_414 (O_414,N_18661,N_19801);
nor UO_415 (O_415,N_19893,N_19377);
nand UO_416 (O_416,N_19023,N_18709);
nand UO_417 (O_417,N_19545,N_19670);
nand UO_418 (O_418,N_18168,N_18444);
nor UO_419 (O_419,N_18066,N_19602);
nand UO_420 (O_420,N_18006,N_19743);
xnor UO_421 (O_421,N_18761,N_18052);
nor UO_422 (O_422,N_19136,N_18558);
nor UO_423 (O_423,N_18993,N_19119);
and UO_424 (O_424,N_19585,N_19522);
or UO_425 (O_425,N_19646,N_19594);
or UO_426 (O_426,N_19423,N_19175);
xnor UO_427 (O_427,N_18493,N_19167);
and UO_428 (O_428,N_19735,N_18129);
nand UO_429 (O_429,N_18459,N_18504);
nor UO_430 (O_430,N_19415,N_18165);
or UO_431 (O_431,N_19826,N_18238);
nor UO_432 (O_432,N_18740,N_19337);
xnor UO_433 (O_433,N_18890,N_19940);
nand UO_434 (O_434,N_18112,N_19742);
nand UO_435 (O_435,N_18013,N_19244);
nand UO_436 (O_436,N_19853,N_19000);
nand UO_437 (O_437,N_19832,N_18877);
or UO_438 (O_438,N_19300,N_18399);
nand UO_439 (O_439,N_18719,N_19095);
nor UO_440 (O_440,N_18843,N_19445);
nor UO_441 (O_441,N_18289,N_18318);
nor UO_442 (O_442,N_19421,N_18426);
nor UO_443 (O_443,N_19980,N_19182);
nor UO_444 (O_444,N_19797,N_19121);
nor UO_445 (O_445,N_18786,N_18688);
nand UO_446 (O_446,N_19589,N_18382);
and UO_447 (O_447,N_18454,N_18637);
nor UO_448 (O_448,N_19790,N_19043);
or UO_449 (O_449,N_18977,N_18659);
nor UO_450 (O_450,N_19202,N_18028);
nand UO_451 (O_451,N_18151,N_18093);
or UO_452 (O_452,N_18241,N_19082);
nand UO_453 (O_453,N_18592,N_19297);
xnor UO_454 (O_454,N_18779,N_18446);
and UO_455 (O_455,N_19349,N_18042);
nand UO_456 (O_456,N_18535,N_19332);
xor UO_457 (O_457,N_18056,N_18026);
nor UO_458 (O_458,N_18842,N_18064);
nand UO_459 (O_459,N_18296,N_19184);
or UO_460 (O_460,N_18221,N_18815);
nor UO_461 (O_461,N_19331,N_18707);
nand UO_462 (O_462,N_18586,N_19590);
or UO_463 (O_463,N_18957,N_18305);
or UO_464 (O_464,N_18432,N_18988);
nand UO_465 (O_465,N_19073,N_18516);
or UO_466 (O_466,N_18440,N_18692);
nand UO_467 (O_467,N_19466,N_19996);
and UO_468 (O_468,N_19675,N_18694);
nand UO_469 (O_469,N_18320,N_19516);
or UO_470 (O_470,N_19083,N_19901);
xnor UO_471 (O_471,N_19444,N_19531);
xnor UO_472 (O_472,N_19923,N_19110);
or UO_473 (O_473,N_19354,N_18720);
nor UO_474 (O_474,N_19982,N_19544);
or UO_475 (O_475,N_18483,N_18005);
or UO_476 (O_476,N_19802,N_18797);
xor UO_477 (O_477,N_18074,N_18696);
nand UO_478 (O_478,N_18102,N_18220);
and UO_479 (O_479,N_18451,N_18254);
nor UO_480 (O_480,N_19016,N_19172);
nor UO_481 (O_481,N_18380,N_19358);
or UO_482 (O_482,N_19881,N_18500);
nor UO_483 (O_483,N_18177,N_19650);
nor UO_484 (O_484,N_18721,N_19367);
xor UO_485 (O_485,N_19620,N_18870);
nand UO_486 (O_486,N_18083,N_18420);
nor UO_487 (O_487,N_18813,N_18345);
nand UO_488 (O_488,N_18803,N_19321);
nor UO_489 (O_489,N_19108,N_18453);
or UO_490 (O_490,N_19010,N_19179);
and UO_491 (O_491,N_18879,N_18108);
or UO_492 (O_492,N_18191,N_19127);
xnor UO_493 (O_493,N_18054,N_19389);
nand UO_494 (O_494,N_18075,N_19313);
nor UO_495 (O_495,N_18984,N_18100);
and UO_496 (O_496,N_19721,N_19756);
or UO_497 (O_497,N_18497,N_18480);
xnor UO_498 (O_498,N_19839,N_18251);
nand UO_499 (O_499,N_18003,N_19546);
or UO_500 (O_500,N_19681,N_18210);
and UO_501 (O_501,N_18347,N_19022);
and UO_502 (O_502,N_18982,N_18071);
or UO_503 (O_503,N_19572,N_18397);
or UO_504 (O_504,N_19874,N_19514);
or UO_505 (O_505,N_19726,N_19451);
and UO_506 (O_506,N_19593,N_19938);
xnor UO_507 (O_507,N_18685,N_18617);
nor UO_508 (O_508,N_19111,N_18478);
or UO_509 (O_509,N_19897,N_19669);
nor UO_510 (O_510,N_18110,N_18359);
nor UO_511 (O_511,N_19062,N_19693);
xor UO_512 (O_512,N_19528,N_19833);
or UO_513 (O_513,N_19314,N_19238);
or UO_514 (O_514,N_19491,N_18381);
or UO_515 (O_515,N_19580,N_19841);
and UO_516 (O_516,N_18261,N_19612);
nor UO_517 (O_517,N_18513,N_19153);
and UO_518 (O_518,N_19248,N_18065);
or UO_519 (O_519,N_19692,N_18233);
nand UO_520 (O_520,N_18222,N_19251);
and UO_521 (O_521,N_19272,N_18199);
nand UO_522 (O_522,N_18032,N_19310);
nor UO_523 (O_523,N_18281,N_18034);
and UO_524 (O_524,N_19144,N_18415);
xnor UO_525 (O_525,N_19819,N_18487);
nor UO_526 (O_526,N_18818,N_18990);
and UO_527 (O_527,N_18471,N_19695);
nor UO_528 (O_528,N_18817,N_19276);
or UO_529 (O_529,N_19513,N_19689);
nand UO_530 (O_530,N_18020,N_18239);
nor UO_531 (O_531,N_18263,N_18427);
nor UO_532 (O_532,N_18673,N_18337);
nand UO_533 (O_533,N_18073,N_19868);
and UO_534 (O_534,N_18484,N_19033);
and UO_535 (O_535,N_18087,N_18273);
nor UO_536 (O_536,N_18816,N_18518);
nand UO_537 (O_537,N_19749,N_18515);
xnor UO_538 (O_538,N_19701,N_18821);
nand UO_539 (O_539,N_19329,N_18211);
nor UO_540 (O_540,N_19610,N_18362);
nor UO_541 (O_541,N_18918,N_18983);
nand UO_542 (O_542,N_19441,N_18450);
and UO_543 (O_543,N_19419,N_19209);
or UO_544 (O_544,N_19059,N_19767);
and UO_545 (O_545,N_18573,N_19909);
nor UO_546 (O_546,N_19193,N_19683);
and UO_547 (O_547,N_18708,N_19150);
and UO_548 (O_548,N_19435,N_19051);
and UO_549 (O_549,N_19249,N_18470);
and UO_550 (O_550,N_18752,N_18295);
xnor UO_551 (O_551,N_19360,N_18033);
or UO_552 (O_552,N_19688,N_18683);
or UO_553 (O_553,N_18445,N_18172);
and UO_554 (O_554,N_19559,N_18545);
nor UO_555 (O_555,N_19479,N_19520);
nand UO_556 (O_556,N_18001,N_18602);
and UO_557 (O_557,N_18755,N_18117);
nor UO_558 (O_558,N_19856,N_18902);
or UO_559 (O_559,N_19619,N_19961);
nor UO_560 (O_560,N_18953,N_19722);
xor UO_561 (O_561,N_19986,N_18554);
and UO_562 (O_562,N_18571,N_18008);
xor UO_563 (O_563,N_19017,N_19991);
xor UO_564 (O_564,N_18784,N_19936);
nor UO_565 (O_565,N_19462,N_19714);
xnor UO_566 (O_566,N_18300,N_18508);
xor UO_567 (O_567,N_18966,N_19012);
nor UO_568 (O_568,N_19375,N_19583);
and UO_569 (O_569,N_19196,N_18252);
xnor UO_570 (O_570,N_19641,N_19303);
or UO_571 (O_571,N_18919,N_19092);
nor UO_572 (O_572,N_19613,N_18301);
or UO_573 (O_573,N_18734,N_19090);
nand UO_574 (O_574,N_18473,N_19014);
or UO_575 (O_575,N_19086,N_18351);
nor UO_576 (O_576,N_18873,N_19935);
xnor UO_577 (O_577,N_19069,N_18948);
nor UO_578 (O_578,N_18521,N_19633);
nand UO_579 (O_579,N_18376,N_19999);
and UO_580 (O_580,N_19887,N_18495);
nand UO_581 (O_581,N_19511,N_19744);
nand UO_582 (O_582,N_18921,N_19578);
xor UO_583 (O_583,N_18017,N_18636);
xnor UO_584 (O_584,N_19629,N_19799);
or UO_585 (O_585,N_19926,N_19401);
nor UO_586 (O_586,N_18456,N_19710);
xor UO_587 (O_587,N_18509,N_19039);
nor UO_588 (O_588,N_18389,N_19976);
nand UO_589 (O_589,N_19533,N_18096);
nor UO_590 (O_590,N_19534,N_18024);
nor UO_591 (O_591,N_19929,N_19133);
nor UO_592 (O_592,N_19852,N_18785);
nor UO_593 (O_593,N_19084,N_19588);
nor UO_594 (O_594,N_18016,N_18695);
nand UO_595 (O_595,N_18475,N_18408);
nand UO_596 (O_596,N_19157,N_19917);
nor UO_597 (O_597,N_18668,N_18581);
xor UO_598 (O_598,N_18651,N_18730);
and UO_599 (O_599,N_18609,N_19189);
xnor UO_600 (O_600,N_18591,N_19535);
and UO_601 (O_601,N_18386,N_19411);
and UO_602 (O_602,N_19339,N_18677);
nand UO_603 (O_603,N_19782,N_19487);
xnor UO_604 (O_604,N_19596,N_18808);
nor UO_605 (O_605,N_18206,N_19621);
nor UO_606 (O_606,N_18265,N_19716);
or UO_607 (O_607,N_18920,N_18835);
nand UO_608 (O_608,N_18832,N_19680);
xor UO_609 (O_609,N_19547,N_19434);
xor UO_610 (O_610,N_19964,N_19431);
and UO_611 (O_611,N_19989,N_19467);
nand UO_612 (O_612,N_19981,N_18549);
xor UO_613 (O_613,N_19027,N_19793);
or UO_614 (O_614,N_19357,N_19765);
and UO_615 (O_615,N_19665,N_18349);
nor UO_616 (O_616,N_18885,N_19861);
or UO_617 (O_617,N_19145,N_18867);
or UO_618 (O_618,N_18693,N_19956);
and UO_619 (O_619,N_19173,N_19657);
and UO_620 (O_620,N_19939,N_19005);
or UO_621 (O_621,N_18583,N_19988);
nor UO_622 (O_622,N_19739,N_18577);
and UO_623 (O_623,N_19220,N_18652);
and UO_624 (O_624,N_18505,N_19471);
nor UO_625 (O_625,N_18438,N_19812);
nor UO_626 (O_626,N_19382,N_19345);
xor UO_627 (O_627,N_18405,N_18622);
and UO_628 (O_628,N_18589,N_19586);
nand UO_629 (O_629,N_18491,N_18682);
and UO_630 (O_630,N_18299,N_19243);
xor UO_631 (O_631,N_18901,N_18204);
nand UO_632 (O_632,N_19560,N_19809);
xnor UO_633 (O_633,N_19306,N_19778);
nand UO_634 (O_634,N_19256,N_18166);
xnor UO_635 (O_635,N_19842,N_18955);
nor UO_636 (O_636,N_18627,N_19164);
and UO_637 (O_637,N_18819,N_19835);
xnor UO_638 (O_638,N_19402,N_18907);
nor UO_639 (O_639,N_18037,N_18258);
xor UO_640 (O_640,N_19374,N_19502);
or UO_641 (O_641,N_18506,N_19747);
nor UO_642 (O_642,N_18917,N_18407);
and UO_643 (O_643,N_19338,N_19258);
nor UO_644 (O_644,N_18144,N_18079);
nor UO_645 (O_645,N_19429,N_19420);
nand UO_646 (O_646,N_19556,N_19857);
xor UO_647 (O_647,N_19611,N_18825);
xor UO_648 (O_648,N_18687,N_18421);
and UO_649 (O_649,N_19554,N_18945);
xor UO_650 (O_650,N_19779,N_19327);
or UO_651 (O_651,N_18874,N_18838);
nor UO_652 (O_652,N_18392,N_18511);
nand UO_653 (O_653,N_18751,N_18388);
and UO_654 (O_654,N_18970,N_18985);
nand UO_655 (O_655,N_18009,N_19312);
nand UO_656 (O_656,N_19754,N_18216);
and UO_657 (O_657,N_18996,N_18361);
nor UO_658 (O_658,N_19796,N_19952);
xor UO_659 (O_659,N_18722,N_18086);
nor UO_660 (O_660,N_19071,N_18312);
or UO_661 (O_661,N_18259,N_18940);
nand UO_662 (O_662,N_19050,N_19889);
nand UO_663 (O_663,N_18572,N_19880);
nand UO_664 (O_664,N_19994,N_18961);
and UO_665 (O_665,N_19056,N_18772);
and UO_666 (O_666,N_19844,N_18142);
nand UO_667 (O_667,N_19647,N_18741);
nand UO_668 (O_668,N_19776,N_18975);
xnor UO_669 (O_669,N_19786,N_18235);
nand UO_670 (O_670,N_18275,N_18167);
or UO_671 (O_671,N_19151,N_18946);
or UO_672 (O_672,N_18293,N_19201);
and UO_673 (O_673,N_19068,N_19386);
xor UO_674 (O_674,N_18528,N_18106);
xor UO_675 (O_675,N_18979,N_18548);
nor UO_676 (O_676,N_18593,N_18738);
nand UO_677 (O_677,N_18806,N_19971);
or UO_678 (O_678,N_19105,N_18743);
or UO_679 (O_679,N_18184,N_19755);
or UO_680 (O_680,N_18849,N_18700);
nand UO_681 (O_681,N_19626,N_19355);
and UO_682 (O_682,N_18567,N_19187);
nand UO_683 (O_683,N_18217,N_19700);
xnor UO_684 (O_684,N_18203,N_19336);
nor UO_685 (O_685,N_19192,N_19493);
xor UO_686 (O_686,N_19685,N_18600);
and UO_687 (O_687,N_18194,N_19553);
xnor UO_688 (O_688,N_19840,N_19152);
nand UO_689 (O_689,N_19461,N_18154);
nor UO_690 (O_690,N_19974,N_19617);
and UO_691 (O_691,N_18971,N_18704);
xnor UO_692 (O_692,N_18667,N_19798);
and UO_693 (O_693,N_18732,N_19255);
xnor UO_694 (O_694,N_19992,N_18702);
xnor UO_695 (O_695,N_19846,N_19190);
and UO_696 (O_696,N_18366,N_18363);
nand UO_697 (O_697,N_19362,N_19882);
nand UO_698 (O_698,N_18624,N_19304);
nand UO_699 (O_699,N_18766,N_18643);
xnor UO_700 (O_700,N_18460,N_18192);
nor UO_701 (O_701,N_19943,N_18039);
and UO_702 (O_702,N_18162,N_18608);
and UO_703 (O_703,N_18642,N_18324);
or UO_704 (O_704,N_19147,N_19379);
and UO_705 (O_705,N_18697,N_19030);
xnor UO_706 (O_706,N_19281,N_19296);
and UO_707 (O_707,N_18023,N_19087);
or UO_708 (O_708,N_19245,N_18566);
or UO_709 (O_709,N_19618,N_19888);
or UO_710 (O_710,N_19603,N_18649);
and UO_711 (O_711,N_18989,N_18802);
nand UO_712 (O_712,N_19305,N_19869);
nand UO_713 (O_713,N_18791,N_18198);
nand UO_714 (O_714,N_19218,N_19780);
xor UO_715 (O_715,N_18055,N_19937);
nand UO_716 (O_716,N_18109,N_18435);
or UO_717 (O_717,N_18810,N_19492);
nor UO_718 (O_718,N_19891,N_18863);
nand UO_719 (O_719,N_18462,N_19484);
or UO_720 (O_720,N_18132,N_18925);
xnor UO_721 (O_721,N_19315,N_19718);
xor UO_722 (O_722,N_18759,N_19625);
nand UO_723 (O_723,N_18089,N_18664);
and UO_724 (O_724,N_18428,N_19237);
or UO_725 (O_725,N_18323,N_18183);
nand UO_726 (O_726,N_18846,N_18404);
nand UO_727 (O_727,N_19566,N_19407);
nor UO_728 (O_728,N_18974,N_19927);
nand UO_729 (O_729,N_18304,N_18633);
or UO_730 (O_730,N_18949,N_19085);
nor UO_731 (O_731,N_18051,N_19945);
and UO_732 (O_732,N_19229,N_19599);
and UO_733 (O_733,N_19845,N_19042);
and UO_734 (O_734,N_19275,N_19730);
nand UO_735 (O_735,N_19568,N_19260);
and UO_736 (O_736,N_19751,N_18646);
nand UO_737 (O_737,N_19397,N_18742);
xor UO_738 (O_738,N_19709,N_19763);
nor UO_739 (O_739,N_18111,N_19581);
nor UO_740 (O_740,N_18647,N_19286);
xnor UO_741 (O_741,N_19557,N_19299);
nand UO_742 (O_742,N_19501,N_18455);
and UO_743 (O_743,N_19984,N_18568);
nor UO_744 (O_744,N_19408,N_18632);
nor UO_745 (O_745,N_18690,N_18343);
and UO_746 (O_746,N_18019,N_18338);
or UO_747 (O_747,N_18780,N_18575);
nor UO_748 (O_748,N_19406,N_19066);
or UO_749 (O_749,N_19387,N_19115);
xnor UO_750 (O_750,N_18994,N_18171);
xor UO_751 (O_751,N_18899,N_19122);
nand UO_752 (O_752,N_19166,N_18246);
nor UO_753 (O_753,N_19262,N_19089);
nand UO_754 (O_754,N_18980,N_19630);
nand UO_755 (O_755,N_19913,N_19368);
nor UO_756 (O_756,N_19859,N_18278);
xor UO_757 (O_757,N_19443,N_18333);
and UO_758 (O_758,N_19772,N_18292);
xnor UO_759 (O_759,N_18118,N_19563);
or UO_760 (O_760,N_19101,N_18520);
or UO_761 (O_761,N_19294,N_18856);
xnor UO_762 (O_762,N_18173,N_18175);
xnor UO_763 (O_763,N_19029,N_19953);
or UO_764 (O_764,N_19283,N_19344);
nor UO_765 (O_765,N_19285,N_19605);
nand UO_766 (O_766,N_18080,N_18855);
nand UO_767 (O_767,N_19740,N_18809);
and UO_768 (O_768,N_18670,N_19677);
and UO_769 (O_769,N_19737,N_18352);
xor UO_770 (O_770,N_19905,N_18547);
nand UO_771 (O_771,N_19414,N_19609);
xor UO_772 (O_772,N_18795,N_18799);
nand UO_773 (O_773,N_18022,N_19465);
or UO_774 (O_774,N_19705,N_18739);
nand UO_775 (O_775,N_19604,N_18858);
nand UO_776 (O_776,N_18678,N_18936);
nand UO_777 (O_777,N_19707,N_18141);
nand UO_778 (O_778,N_18084,N_19002);
nand UO_779 (O_779,N_18402,N_18044);
xor UO_780 (O_780,N_18302,N_18114);
or UO_781 (O_781,N_18644,N_18181);
or UO_782 (O_782,N_18092,N_18474);
nor UO_783 (O_783,N_19058,N_19450);
or UO_784 (O_784,N_19078,N_19703);
nand UO_785 (O_785,N_19499,N_18326);
and UO_786 (O_786,N_18943,N_18724);
xor UO_787 (O_787,N_18424,N_18157);
nand UO_788 (O_788,N_19400,N_19094);
or UO_789 (O_789,N_19273,N_19564);
and UO_790 (O_790,N_19827,N_18926);
and UO_791 (O_791,N_19160,N_19436);
nand UO_792 (O_792,N_19186,N_18091);
nor UO_793 (O_793,N_19463,N_18306);
or UO_794 (O_794,N_18765,N_19831);
nor UO_795 (O_795,N_18449,N_19792);
and UO_796 (O_796,N_19052,N_19170);
nor UO_797 (O_797,N_18585,N_18205);
xor UO_798 (O_798,N_19561,N_18231);
nor UO_799 (O_799,N_18468,N_18564);
nand UO_800 (O_800,N_19426,N_19512);
nand UO_801 (O_801,N_18540,N_19530);
nor UO_802 (O_802,N_19672,N_18317);
or UO_803 (O_803,N_19634,N_18410);
or UO_804 (O_804,N_19240,N_19800);
nand UO_805 (O_805,N_19950,N_19969);
and UO_806 (O_806,N_19433,N_19904);
or UO_807 (O_807,N_19649,N_19096);
or UO_808 (O_808,N_18365,N_18422);
or UO_809 (O_809,N_19567,N_18601);
and UO_810 (O_810,N_18029,N_19736);
and UO_811 (O_811,N_18850,N_18145);
and UO_812 (O_812,N_19539,N_18336);
nor UO_813 (O_813,N_19543,N_19370);
and UO_814 (O_814,N_19678,N_19020);
xnor UO_815 (O_815,N_19104,N_18189);
or UO_816 (O_816,N_19548,N_18396);
nand UO_817 (O_817,N_18648,N_19015);
nand UO_818 (O_818,N_19808,N_19158);
xnor UO_819 (O_819,N_19694,N_19495);
or UO_820 (O_820,N_19477,N_19930);
or UO_821 (O_821,N_18588,N_18812);
and UO_822 (O_822,N_19702,N_19162);
nor UO_823 (O_823,N_19746,N_19933);
nor UO_824 (O_824,N_18612,N_19774);
nor UO_825 (O_825,N_19518,N_18321);
and UO_826 (O_826,N_19729,N_19129);
and UO_827 (O_827,N_19922,N_19100);
nand UO_828 (O_828,N_18753,N_18327);
or UO_829 (O_829,N_19340,N_18476);
nor UO_830 (O_830,N_19640,N_19745);
xor UO_831 (O_831,N_18546,N_18532);
nor UO_832 (O_832,N_18997,N_19759);
and UO_833 (O_833,N_18309,N_18900);
and UO_834 (O_834,N_19764,N_18250);
nor UO_835 (O_835,N_19215,N_19212);
or UO_836 (O_836,N_18159,N_18526);
and UO_837 (O_837,N_19894,N_19308);
xnor UO_838 (O_838,N_19241,N_19944);
or UO_839 (O_839,N_19920,N_18282);
and UO_840 (O_840,N_18400,N_19478);
xnor UO_841 (O_841,N_19072,N_18126);
xnor UO_842 (O_842,N_18701,N_19761);
nor UO_843 (O_843,N_19983,N_19899);
or UO_844 (O_844,N_19422,N_18737);
or UO_845 (O_845,N_19113,N_18611);
nand UO_846 (O_846,N_19011,N_18525);
and UO_847 (O_847,N_18128,N_19540);
nand UO_848 (O_848,N_19725,N_18888);
nand UO_849 (O_849,N_19758,N_19676);
nand UO_850 (O_850,N_18411,N_19341);
and UO_851 (O_851,N_18134,N_19486);
nand UO_852 (O_852,N_18557,N_19562);
and UO_853 (O_853,N_18393,N_19474);
or UO_854 (O_854,N_18148,N_18736);
xnor UO_855 (O_855,N_18370,N_18228);
xor UO_856 (O_856,N_18544,N_19376);
and UO_857 (O_857,N_18307,N_19686);
or UO_858 (O_858,N_19204,N_19139);
nor UO_859 (O_859,N_19587,N_19822);
nand UO_860 (O_860,N_19645,N_19008);
xor UO_861 (O_861,N_19892,N_19390);
or UO_862 (O_862,N_18828,N_18430);
nand UO_863 (O_863,N_19473,N_19077);
xor UO_864 (O_864,N_19963,N_19080);
or UO_865 (O_865,N_19047,N_19644);
nor UO_866 (O_866,N_18223,N_19439);
xnor UO_867 (O_867,N_19571,N_19363);
nor UO_868 (O_868,N_18227,N_18560);
nand UO_869 (O_869,N_19064,N_18466);
and UO_870 (O_870,N_18011,N_19600);
nand UO_871 (O_871,N_19109,N_19715);
and UO_872 (O_872,N_18669,N_18862);
nand UO_873 (O_873,N_19573,N_18287);
or UO_874 (O_874,N_19873,N_19055);
xor UO_875 (O_875,N_19886,N_19713);
or UO_876 (O_876,N_19638,N_19606);
nor UO_877 (O_877,N_18717,N_19148);
or UO_878 (O_878,N_18085,N_18735);
and UO_879 (O_879,N_18837,N_18035);
nor UO_880 (O_880,N_18910,N_18932);
xnor UO_881 (O_881,N_18182,N_18105);
xor UO_882 (O_882,N_18398,N_19472);
xor UO_883 (O_883,N_18391,N_18706);
xor UO_884 (O_884,N_19361,N_18635);
and UO_885 (O_885,N_18666,N_18747);
or UO_886 (O_886,N_18463,N_19954);
and UO_887 (O_887,N_19333,N_18864);
xnor UO_888 (O_888,N_18923,N_18965);
nor UO_889 (O_889,N_19464,N_19230);
or UO_890 (O_890,N_19876,N_18507);
or UO_891 (O_891,N_18053,N_18576);
and UO_892 (O_892,N_18956,N_19949);
nand UO_893 (O_893,N_18579,N_18319);
or UO_894 (O_894,N_18423,N_18829);
nor UO_895 (O_895,N_19653,N_18963);
or UO_896 (O_896,N_18715,N_19232);
nor UO_897 (O_897,N_19542,N_18640);
nor UO_898 (O_898,N_19687,N_19664);
xnor UO_899 (O_899,N_19942,N_18674);
xor UO_900 (O_900,N_19898,N_19978);
nand UO_901 (O_901,N_18705,N_18844);
nand UO_902 (O_902,N_19711,N_18315);
nor UO_903 (O_903,N_18656,N_19918);
or UO_904 (O_904,N_18607,N_19404);
nand UO_905 (O_905,N_19270,N_19330);
or UO_906 (O_906,N_18489,N_18911);
or UO_907 (O_907,N_19785,N_19690);
xnor UO_908 (O_908,N_18160,N_18660);
xnor UO_909 (O_909,N_18594,N_19975);
xnor UO_910 (O_910,N_18895,N_19497);
nand UO_911 (O_911,N_18479,N_19424);
or UO_912 (O_912,N_19460,N_19102);
xnor UO_913 (O_913,N_19447,N_19366);
nand UO_914 (O_914,N_18195,N_18625);
xnor UO_915 (O_915,N_18107,N_19428);
and UO_916 (O_916,N_18286,N_18847);
or UO_917 (O_917,N_19498,N_19035);
nor UO_918 (O_918,N_18524,N_19494);
or UO_919 (O_919,N_19720,N_19608);
nand UO_920 (O_920,N_19223,N_18680);
or UO_921 (O_921,N_19552,N_18350);
and UO_922 (O_922,N_19399,N_19967);
or UO_923 (O_923,N_18929,N_18499);
xnor UO_924 (O_924,N_18038,N_18088);
xnor UO_925 (O_925,N_19507,N_19246);
nor UO_926 (O_926,N_19648,N_18163);
and UO_927 (O_927,N_18882,N_18358);
xor UO_928 (O_928,N_19268,N_18630);
xnor UO_929 (O_929,N_18924,N_18010);
and UO_930 (O_930,N_18230,N_19266);
and UO_931 (O_931,N_18562,N_19171);
nand UO_932 (O_932,N_18346,N_19185);
nand UO_933 (O_933,N_18045,N_18047);
or UO_934 (O_934,N_19582,N_18553);
xnor UO_935 (O_935,N_19393,N_19372);
and UO_936 (O_936,N_18237,N_18488);
nor UO_937 (O_937,N_19805,N_18041);
xnor UO_938 (O_938,N_18127,N_19347);
and UO_939 (O_939,N_19480,N_19253);
or UO_940 (O_940,N_18121,N_19396);
and UO_941 (O_941,N_18197,N_18514);
or UO_942 (O_942,N_19416,N_18972);
and UO_943 (O_943,N_18746,N_19903);
or UO_944 (O_944,N_18448,N_18458);
nor UO_945 (O_945,N_18710,N_18255);
nand UO_946 (O_946,N_19807,N_18789);
and UO_947 (O_947,N_18272,N_18280);
nor UO_948 (O_948,N_18501,N_19350);
nand UO_949 (O_949,N_19124,N_18875);
or UO_950 (O_950,N_19317,N_19457);
nor UO_951 (O_951,N_18417,N_19278);
or UO_952 (O_952,N_18912,N_19410);
and UO_953 (O_953,N_18139,N_19468);
or UO_954 (O_954,N_18164,N_18201);
and UO_955 (O_955,N_19708,N_19658);
xnor UO_956 (O_956,N_19383,N_18783);
nand UO_957 (O_957,N_19351,N_18373);
and UO_958 (O_958,N_19335,N_18999);
xnor UO_959 (O_959,N_18207,N_18800);
xor UO_960 (O_960,N_18613,N_19181);
xor UO_961 (O_961,N_19970,N_18866);
nor UO_962 (O_962,N_19252,N_18964);
nor UO_963 (O_963,N_19592,N_19616);
nand UO_964 (O_964,N_19236,N_18316);
or UO_965 (O_965,N_19044,N_18158);
nor UO_966 (O_966,N_18658,N_18950);
xnor UO_967 (O_967,N_18416,N_18512);
nand UO_968 (O_968,N_18606,N_18249);
and UO_969 (O_969,N_19483,N_19654);
nand UO_970 (O_970,N_18883,N_18355);
xnor UO_971 (O_971,N_18027,N_18531);
nor UO_972 (O_972,N_18523,N_19928);
and UO_973 (O_973,N_18000,N_18913);
xnor UO_974 (O_974,N_19768,N_19517);
or UO_975 (O_975,N_18610,N_18922);
nor UO_976 (O_976,N_18169,N_18954);
nand UO_977 (O_977,N_18097,N_18288);
nand UO_978 (O_978,N_18939,N_18529);
or UO_979 (O_979,N_18179,N_19931);
and UO_980 (O_980,N_18224,N_19508);
nand UO_981 (O_981,N_19579,N_19574);
and UO_982 (O_982,N_19752,N_18543);
nor UO_983 (O_983,N_18968,N_18298);
or UO_984 (O_984,N_19099,N_19116);
nor UO_985 (O_985,N_19523,N_18675);
and UO_986 (O_986,N_18536,N_18072);
or UO_987 (O_987,N_18076,N_18931);
nor UO_988 (O_988,N_18379,N_19951);
or UO_989 (O_989,N_19199,N_19663);
or UO_990 (O_990,N_19906,N_19128);
nand UO_991 (O_991,N_18672,N_19130);
and UO_992 (O_992,N_19806,N_19040);
nor UO_993 (O_993,N_18077,N_19198);
nor UO_994 (O_994,N_19674,N_19555);
nor UO_995 (O_995,N_19316,N_18113);
nand UO_996 (O_996,N_18137,N_18274);
xor UO_997 (O_997,N_19112,N_18826);
and UO_998 (O_998,N_19958,N_18757);
xnor UO_999 (O_999,N_19837,N_18457);
xnor UO_1000 (O_1000,N_19533,N_18250);
nor UO_1001 (O_1001,N_18703,N_18627);
xor UO_1002 (O_1002,N_19727,N_19200);
nand UO_1003 (O_1003,N_18193,N_18337);
or UO_1004 (O_1004,N_18088,N_18459);
nor UO_1005 (O_1005,N_18061,N_18127);
and UO_1006 (O_1006,N_19353,N_18634);
nand UO_1007 (O_1007,N_18345,N_18022);
xor UO_1008 (O_1008,N_18570,N_18427);
xor UO_1009 (O_1009,N_18421,N_19801);
nand UO_1010 (O_1010,N_19738,N_18598);
nand UO_1011 (O_1011,N_18976,N_18526);
xor UO_1012 (O_1012,N_18110,N_19335);
and UO_1013 (O_1013,N_18200,N_19179);
nand UO_1014 (O_1014,N_19827,N_18271);
nor UO_1015 (O_1015,N_18905,N_19965);
or UO_1016 (O_1016,N_18263,N_19413);
nor UO_1017 (O_1017,N_18938,N_19569);
or UO_1018 (O_1018,N_19509,N_19180);
or UO_1019 (O_1019,N_19451,N_18581);
xnor UO_1020 (O_1020,N_19780,N_19685);
nor UO_1021 (O_1021,N_18336,N_18022);
and UO_1022 (O_1022,N_18329,N_18832);
nor UO_1023 (O_1023,N_18171,N_18677);
and UO_1024 (O_1024,N_19001,N_18021);
nor UO_1025 (O_1025,N_18512,N_18314);
or UO_1026 (O_1026,N_18274,N_18319);
and UO_1027 (O_1027,N_19057,N_19361);
nand UO_1028 (O_1028,N_18527,N_19074);
xor UO_1029 (O_1029,N_18136,N_19216);
nand UO_1030 (O_1030,N_19795,N_19829);
and UO_1031 (O_1031,N_18454,N_19871);
and UO_1032 (O_1032,N_18101,N_19925);
nand UO_1033 (O_1033,N_19629,N_19257);
nor UO_1034 (O_1034,N_19016,N_18349);
nand UO_1035 (O_1035,N_18609,N_18688);
nand UO_1036 (O_1036,N_19143,N_18497);
nand UO_1037 (O_1037,N_18193,N_19108);
xor UO_1038 (O_1038,N_18011,N_18214);
nor UO_1039 (O_1039,N_18793,N_18910);
or UO_1040 (O_1040,N_19903,N_18712);
nand UO_1041 (O_1041,N_18782,N_19560);
xor UO_1042 (O_1042,N_19751,N_19421);
xnor UO_1043 (O_1043,N_19016,N_19085);
nand UO_1044 (O_1044,N_19604,N_19269);
nand UO_1045 (O_1045,N_18579,N_19614);
or UO_1046 (O_1046,N_19228,N_19245);
nand UO_1047 (O_1047,N_19678,N_19078);
nand UO_1048 (O_1048,N_19811,N_19598);
and UO_1049 (O_1049,N_19635,N_18586);
nand UO_1050 (O_1050,N_19247,N_19290);
nand UO_1051 (O_1051,N_19289,N_18273);
and UO_1052 (O_1052,N_18452,N_18693);
or UO_1053 (O_1053,N_18514,N_18327);
or UO_1054 (O_1054,N_19464,N_18500);
or UO_1055 (O_1055,N_18426,N_18256);
or UO_1056 (O_1056,N_19289,N_18577);
and UO_1057 (O_1057,N_19666,N_18600);
nand UO_1058 (O_1058,N_18355,N_19603);
nor UO_1059 (O_1059,N_19170,N_19221);
nor UO_1060 (O_1060,N_19665,N_19515);
nor UO_1061 (O_1061,N_19842,N_19337);
or UO_1062 (O_1062,N_18647,N_19044);
xor UO_1063 (O_1063,N_19271,N_18964);
xor UO_1064 (O_1064,N_18746,N_18289);
and UO_1065 (O_1065,N_19425,N_18256);
xnor UO_1066 (O_1066,N_19629,N_19747);
nand UO_1067 (O_1067,N_18903,N_18517);
nor UO_1068 (O_1068,N_19835,N_18287);
or UO_1069 (O_1069,N_18905,N_18298);
nand UO_1070 (O_1070,N_19266,N_19703);
nor UO_1071 (O_1071,N_18674,N_18097);
nand UO_1072 (O_1072,N_18955,N_19645);
and UO_1073 (O_1073,N_19043,N_18084);
and UO_1074 (O_1074,N_18363,N_18457);
nand UO_1075 (O_1075,N_18836,N_18098);
xnor UO_1076 (O_1076,N_18793,N_18242);
and UO_1077 (O_1077,N_18503,N_18242);
nor UO_1078 (O_1078,N_19608,N_18410);
nand UO_1079 (O_1079,N_18886,N_18663);
or UO_1080 (O_1080,N_19632,N_19503);
or UO_1081 (O_1081,N_18013,N_18822);
nand UO_1082 (O_1082,N_19542,N_19086);
and UO_1083 (O_1083,N_19889,N_19748);
or UO_1084 (O_1084,N_18315,N_18047);
and UO_1085 (O_1085,N_18354,N_18437);
xnor UO_1086 (O_1086,N_19685,N_19591);
nor UO_1087 (O_1087,N_19274,N_18347);
nand UO_1088 (O_1088,N_19862,N_19204);
or UO_1089 (O_1089,N_19324,N_19922);
nand UO_1090 (O_1090,N_19990,N_18543);
and UO_1091 (O_1091,N_19273,N_19656);
or UO_1092 (O_1092,N_19401,N_18401);
and UO_1093 (O_1093,N_18230,N_18616);
nor UO_1094 (O_1094,N_19882,N_19249);
nor UO_1095 (O_1095,N_18669,N_18487);
nand UO_1096 (O_1096,N_18261,N_18014);
or UO_1097 (O_1097,N_19962,N_19470);
and UO_1098 (O_1098,N_19297,N_18186);
or UO_1099 (O_1099,N_19267,N_19636);
xnor UO_1100 (O_1100,N_19063,N_18126);
xnor UO_1101 (O_1101,N_19455,N_19626);
or UO_1102 (O_1102,N_18520,N_19509);
nand UO_1103 (O_1103,N_18223,N_18592);
nor UO_1104 (O_1104,N_18813,N_19182);
xor UO_1105 (O_1105,N_19417,N_19831);
xor UO_1106 (O_1106,N_18676,N_19093);
nor UO_1107 (O_1107,N_19079,N_18620);
nor UO_1108 (O_1108,N_18783,N_18904);
nor UO_1109 (O_1109,N_18510,N_18185);
and UO_1110 (O_1110,N_18091,N_19780);
xnor UO_1111 (O_1111,N_18788,N_18978);
nand UO_1112 (O_1112,N_19051,N_19944);
or UO_1113 (O_1113,N_18440,N_19054);
and UO_1114 (O_1114,N_18142,N_18054);
and UO_1115 (O_1115,N_19303,N_18310);
or UO_1116 (O_1116,N_19215,N_18686);
or UO_1117 (O_1117,N_18801,N_19525);
nand UO_1118 (O_1118,N_18783,N_19469);
nor UO_1119 (O_1119,N_18384,N_19217);
nor UO_1120 (O_1120,N_18331,N_19925);
or UO_1121 (O_1121,N_19067,N_19519);
xnor UO_1122 (O_1122,N_19344,N_18015);
and UO_1123 (O_1123,N_19932,N_19597);
xor UO_1124 (O_1124,N_19186,N_18677);
nand UO_1125 (O_1125,N_19553,N_18702);
nor UO_1126 (O_1126,N_19371,N_18005);
or UO_1127 (O_1127,N_18049,N_19372);
xor UO_1128 (O_1128,N_18773,N_18844);
xor UO_1129 (O_1129,N_18076,N_19805);
or UO_1130 (O_1130,N_18971,N_19666);
or UO_1131 (O_1131,N_18030,N_18328);
nand UO_1132 (O_1132,N_18260,N_18570);
nand UO_1133 (O_1133,N_18178,N_18247);
and UO_1134 (O_1134,N_18522,N_18883);
nor UO_1135 (O_1135,N_19234,N_19242);
nor UO_1136 (O_1136,N_18304,N_19647);
nand UO_1137 (O_1137,N_19209,N_19889);
and UO_1138 (O_1138,N_18987,N_19233);
nand UO_1139 (O_1139,N_19775,N_18947);
nor UO_1140 (O_1140,N_18455,N_19659);
nand UO_1141 (O_1141,N_18295,N_18233);
nand UO_1142 (O_1142,N_18746,N_19461);
xnor UO_1143 (O_1143,N_19312,N_19665);
or UO_1144 (O_1144,N_19533,N_19680);
nand UO_1145 (O_1145,N_19642,N_19483);
xor UO_1146 (O_1146,N_19937,N_18977);
nor UO_1147 (O_1147,N_19352,N_19474);
or UO_1148 (O_1148,N_19831,N_19255);
nand UO_1149 (O_1149,N_18717,N_19162);
xnor UO_1150 (O_1150,N_18771,N_19457);
or UO_1151 (O_1151,N_18160,N_18054);
xor UO_1152 (O_1152,N_18752,N_18297);
or UO_1153 (O_1153,N_19470,N_19899);
xnor UO_1154 (O_1154,N_19327,N_18673);
nor UO_1155 (O_1155,N_18312,N_19798);
xnor UO_1156 (O_1156,N_19483,N_19918);
and UO_1157 (O_1157,N_19835,N_19849);
and UO_1158 (O_1158,N_19189,N_18659);
nor UO_1159 (O_1159,N_19776,N_19668);
and UO_1160 (O_1160,N_18847,N_18443);
xnor UO_1161 (O_1161,N_19495,N_19884);
xor UO_1162 (O_1162,N_19557,N_19988);
or UO_1163 (O_1163,N_19070,N_18714);
nor UO_1164 (O_1164,N_19894,N_19873);
or UO_1165 (O_1165,N_19714,N_19381);
or UO_1166 (O_1166,N_18750,N_18679);
nor UO_1167 (O_1167,N_18968,N_19460);
xor UO_1168 (O_1168,N_18024,N_19555);
and UO_1169 (O_1169,N_18983,N_18462);
or UO_1170 (O_1170,N_18764,N_18155);
nand UO_1171 (O_1171,N_19879,N_18754);
or UO_1172 (O_1172,N_19722,N_18800);
nor UO_1173 (O_1173,N_19533,N_18588);
xnor UO_1174 (O_1174,N_19656,N_19407);
nor UO_1175 (O_1175,N_19690,N_18906);
xnor UO_1176 (O_1176,N_19454,N_19888);
or UO_1177 (O_1177,N_19052,N_19133);
or UO_1178 (O_1178,N_18352,N_18665);
and UO_1179 (O_1179,N_19694,N_19575);
nor UO_1180 (O_1180,N_19632,N_18582);
xnor UO_1181 (O_1181,N_18243,N_19926);
or UO_1182 (O_1182,N_19646,N_19494);
nor UO_1183 (O_1183,N_18330,N_18194);
or UO_1184 (O_1184,N_18245,N_18931);
or UO_1185 (O_1185,N_18785,N_19215);
nand UO_1186 (O_1186,N_18267,N_18715);
and UO_1187 (O_1187,N_19719,N_19397);
nor UO_1188 (O_1188,N_19282,N_18559);
nand UO_1189 (O_1189,N_19041,N_18000);
nand UO_1190 (O_1190,N_18282,N_19666);
xnor UO_1191 (O_1191,N_19700,N_18203);
xnor UO_1192 (O_1192,N_19202,N_19981);
or UO_1193 (O_1193,N_18017,N_18153);
or UO_1194 (O_1194,N_19699,N_18069);
and UO_1195 (O_1195,N_19096,N_19994);
or UO_1196 (O_1196,N_18439,N_18598);
and UO_1197 (O_1197,N_19300,N_19799);
or UO_1198 (O_1198,N_18949,N_19554);
and UO_1199 (O_1199,N_19557,N_18171);
xnor UO_1200 (O_1200,N_18256,N_18958);
nand UO_1201 (O_1201,N_18290,N_18471);
and UO_1202 (O_1202,N_18513,N_18779);
nor UO_1203 (O_1203,N_19996,N_19684);
or UO_1204 (O_1204,N_18831,N_19429);
and UO_1205 (O_1205,N_19982,N_18496);
nor UO_1206 (O_1206,N_19234,N_18572);
and UO_1207 (O_1207,N_19075,N_18678);
and UO_1208 (O_1208,N_18200,N_19799);
or UO_1209 (O_1209,N_19670,N_18705);
nand UO_1210 (O_1210,N_18292,N_19666);
or UO_1211 (O_1211,N_19905,N_19661);
and UO_1212 (O_1212,N_19964,N_18529);
xnor UO_1213 (O_1213,N_18168,N_19964);
nor UO_1214 (O_1214,N_18752,N_19361);
xor UO_1215 (O_1215,N_19684,N_19208);
and UO_1216 (O_1216,N_19687,N_18817);
nor UO_1217 (O_1217,N_19482,N_19565);
nor UO_1218 (O_1218,N_19271,N_18073);
or UO_1219 (O_1219,N_18116,N_18199);
nor UO_1220 (O_1220,N_18344,N_19273);
and UO_1221 (O_1221,N_18969,N_19591);
xor UO_1222 (O_1222,N_19478,N_19929);
and UO_1223 (O_1223,N_18502,N_19271);
nand UO_1224 (O_1224,N_19844,N_19391);
xnor UO_1225 (O_1225,N_18104,N_18819);
and UO_1226 (O_1226,N_18779,N_18223);
or UO_1227 (O_1227,N_18223,N_18827);
xor UO_1228 (O_1228,N_19941,N_19837);
and UO_1229 (O_1229,N_19152,N_19276);
nand UO_1230 (O_1230,N_19117,N_18612);
and UO_1231 (O_1231,N_19413,N_19529);
nand UO_1232 (O_1232,N_18060,N_19194);
nand UO_1233 (O_1233,N_19190,N_19377);
xnor UO_1234 (O_1234,N_18029,N_18255);
xnor UO_1235 (O_1235,N_18921,N_19943);
nand UO_1236 (O_1236,N_19393,N_18888);
xnor UO_1237 (O_1237,N_19178,N_19182);
or UO_1238 (O_1238,N_18224,N_18697);
nand UO_1239 (O_1239,N_18069,N_18857);
nand UO_1240 (O_1240,N_18751,N_18089);
nand UO_1241 (O_1241,N_18280,N_19548);
nor UO_1242 (O_1242,N_19473,N_18962);
xor UO_1243 (O_1243,N_18551,N_18723);
nand UO_1244 (O_1244,N_19383,N_18750);
xnor UO_1245 (O_1245,N_19171,N_19023);
xor UO_1246 (O_1246,N_18427,N_19827);
nor UO_1247 (O_1247,N_19601,N_19538);
and UO_1248 (O_1248,N_19444,N_19138);
nor UO_1249 (O_1249,N_18497,N_18879);
or UO_1250 (O_1250,N_19503,N_19104);
nand UO_1251 (O_1251,N_19630,N_18774);
nor UO_1252 (O_1252,N_18216,N_19782);
nand UO_1253 (O_1253,N_18502,N_18913);
or UO_1254 (O_1254,N_18546,N_18678);
and UO_1255 (O_1255,N_18520,N_19479);
nor UO_1256 (O_1256,N_18342,N_18748);
nand UO_1257 (O_1257,N_18698,N_19650);
xor UO_1258 (O_1258,N_18940,N_19540);
and UO_1259 (O_1259,N_19029,N_18167);
nand UO_1260 (O_1260,N_18369,N_18255);
xor UO_1261 (O_1261,N_19006,N_19851);
nor UO_1262 (O_1262,N_18880,N_18324);
nand UO_1263 (O_1263,N_19588,N_18290);
nand UO_1264 (O_1264,N_19330,N_18193);
nand UO_1265 (O_1265,N_19218,N_18751);
nor UO_1266 (O_1266,N_18914,N_18695);
nor UO_1267 (O_1267,N_18167,N_19458);
or UO_1268 (O_1268,N_18176,N_19252);
xor UO_1269 (O_1269,N_19533,N_18554);
nor UO_1270 (O_1270,N_19314,N_18514);
nor UO_1271 (O_1271,N_18041,N_19089);
xor UO_1272 (O_1272,N_18809,N_18365);
xor UO_1273 (O_1273,N_18576,N_18771);
nand UO_1274 (O_1274,N_18171,N_19966);
and UO_1275 (O_1275,N_18468,N_19476);
or UO_1276 (O_1276,N_19730,N_19292);
or UO_1277 (O_1277,N_19116,N_19000);
nand UO_1278 (O_1278,N_18907,N_19075);
or UO_1279 (O_1279,N_18602,N_19674);
or UO_1280 (O_1280,N_18638,N_19702);
and UO_1281 (O_1281,N_18283,N_18084);
nand UO_1282 (O_1282,N_19825,N_19884);
or UO_1283 (O_1283,N_18308,N_19417);
nand UO_1284 (O_1284,N_18569,N_18671);
or UO_1285 (O_1285,N_18699,N_19297);
nand UO_1286 (O_1286,N_19020,N_18742);
or UO_1287 (O_1287,N_18028,N_18267);
xnor UO_1288 (O_1288,N_19206,N_19800);
xnor UO_1289 (O_1289,N_18668,N_18944);
nand UO_1290 (O_1290,N_18461,N_18968);
or UO_1291 (O_1291,N_19609,N_19651);
nand UO_1292 (O_1292,N_19656,N_19332);
or UO_1293 (O_1293,N_19132,N_19026);
nor UO_1294 (O_1294,N_19116,N_19139);
or UO_1295 (O_1295,N_19555,N_19829);
nor UO_1296 (O_1296,N_19359,N_19796);
xnor UO_1297 (O_1297,N_19456,N_18713);
xnor UO_1298 (O_1298,N_18580,N_19538);
nor UO_1299 (O_1299,N_19009,N_19072);
nor UO_1300 (O_1300,N_18625,N_18384);
or UO_1301 (O_1301,N_18369,N_18902);
nand UO_1302 (O_1302,N_19114,N_18883);
or UO_1303 (O_1303,N_19220,N_19209);
or UO_1304 (O_1304,N_18656,N_19919);
and UO_1305 (O_1305,N_18586,N_19736);
nand UO_1306 (O_1306,N_19390,N_19837);
nor UO_1307 (O_1307,N_19405,N_19835);
nand UO_1308 (O_1308,N_19580,N_19724);
nor UO_1309 (O_1309,N_19614,N_18438);
or UO_1310 (O_1310,N_19845,N_19392);
nor UO_1311 (O_1311,N_18537,N_18899);
nand UO_1312 (O_1312,N_18129,N_18982);
nor UO_1313 (O_1313,N_18108,N_19211);
xor UO_1314 (O_1314,N_18120,N_19377);
xor UO_1315 (O_1315,N_18030,N_19145);
xor UO_1316 (O_1316,N_18131,N_18555);
or UO_1317 (O_1317,N_18108,N_19749);
or UO_1318 (O_1318,N_19232,N_18741);
xnor UO_1319 (O_1319,N_19789,N_18668);
xor UO_1320 (O_1320,N_19765,N_18042);
xnor UO_1321 (O_1321,N_19150,N_18996);
xor UO_1322 (O_1322,N_18032,N_18899);
and UO_1323 (O_1323,N_19172,N_19293);
xnor UO_1324 (O_1324,N_18374,N_18471);
xor UO_1325 (O_1325,N_19345,N_19295);
and UO_1326 (O_1326,N_19710,N_18975);
nand UO_1327 (O_1327,N_19162,N_19546);
and UO_1328 (O_1328,N_19790,N_18520);
or UO_1329 (O_1329,N_18422,N_18971);
xor UO_1330 (O_1330,N_19840,N_19711);
nor UO_1331 (O_1331,N_18587,N_18193);
xor UO_1332 (O_1332,N_19172,N_18860);
nor UO_1333 (O_1333,N_18679,N_18178);
and UO_1334 (O_1334,N_18972,N_19022);
and UO_1335 (O_1335,N_18949,N_18197);
nand UO_1336 (O_1336,N_18608,N_19952);
and UO_1337 (O_1337,N_18438,N_18921);
nand UO_1338 (O_1338,N_18506,N_19891);
xnor UO_1339 (O_1339,N_19958,N_18247);
nor UO_1340 (O_1340,N_18805,N_19868);
xor UO_1341 (O_1341,N_19961,N_19001);
xnor UO_1342 (O_1342,N_18183,N_19249);
and UO_1343 (O_1343,N_18159,N_18044);
nand UO_1344 (O_1344,N_19099,N_18208);
and UO_1345 (O_1345,N_19721,N_18192);
xor UO_1346 (O_1346,N_19471,N_19712);
xor UO_1347 (O_1347,N_19606,N_19085);
nor UO_1348 (O_1348,N_19487,N_19069);
and UO_1349 (O_1349,N_18461,N_18288);
or UO_1350 (O_1350,N_19844,N_19093);
and UO_1351 (O_1351,N_18127,N_19674);
xor UO_1352 (O_1352,N_19363,N_18071);
and UO_1353 (O_1353,N_18972,N_19597);
nor UO_1354 (O_1354,N_19675,N_18336);
nor UO_1355 (O_1355,N_19434,N_19058);
xor UO_1356 (O_1356,N_19936,N_18583);
xnor UO_1357 (O_1357,N_18630,N_18629);
and UO_1358 (O_1358,N_19792,N_18401);
nor UO_1359 (O_1359,N_18610,N_19310);
xor UO_1360 (O_1360,N_18571,N_19076);
and UO_1361 (O_1361,N_19541,N_19249);
and UO_1362 (O_1362,N_19144,N_19050);
or UO_1363 (O_1363,N_19825,N_18841);
nand UO_1364 (O_1364,N_19978,N_18188);
and UO_1365 (O_1365,N_19113,N_18833);
nor UO_1366 (O_1366,N_19329,N_18203);
and UO_1367 (O_1367,N_18935,N_19995);
xnor UO_1368 (O_1368,N_18440,N_18613);
or UO_1369 (O_1369,N_19160,N_18762);
nor UO_1370 (O_1370,N_19289,N_18158);
nor UO_1371 (O_1371,N_18389,N_19076);
and UO_1372 (O_1372,N_18818,N_18640);
and UO_1373 (O_1373,N_18667,N_19047);
nand UO_1374 (O_1374,N_19279,N_18335);
xor UO_1375 (O_1375,N_18835,N_19999);
nand UO_1376 (O_1376,N_18827,N_18377);
xnor UO_1377 (O_1377,N_18150,N_18785);
xor UO_1378 (O_1378,N_18226,N_18026);
or UO_1379 (O_1379,N_19678,N_19692);
nand UO_1380 (O_1380,N_19781,N_18915);
nand UO_1381 (O_1381,N_19930,N_19111);
nor UO_1382 (O_1382,N_19976,N_18672);
or UO_1383 (O_1383,N_18091,N_19388);
xnor UO_1384 (O_1384,N_19997,N_18318);
nor UO_1385 (O_1385,N_18882,N_19990);
nand UO_1386 (O_1386,N_19728,N_18042);
xnor UO_1387 (O_1387,N_19307,N_19886);
and UO_1388 (O_1388,N_18397,N_18600);
or UO_1389 (O_1389,N_18264,N_18480);
nand UO_1390 (O_1390,N_18921,N_19069);
nand UO_1391 (O_1391,N_18774,N_18767);
and UO_1392 (O_1392,N_18770,N_19872);
nor UO_1393 (O_1393,N_18196,N_19505);
or UO_1394 (O_1394,N_19265,N_19191);
or UO_1395 (O_1395,N_19841,N_18867);
nor UO_1396 (O_1396,N_19940,N_18920);
nand UO_1397 (O_1397,N_18042,N_18139);
nor UO_1398 (O_1398,N_18815,N_19925);
and UO_1399 (O_1399,N_19638,N_19940);
nor UO_1400 (O_1400,N_19076,N_18436);
and UO_1401 (O_1401,N_19504,N_18552);
and UO_1402 (O_1402,N_19319,N_18693);
and UO_1403 (O_1403,N_18339,N_19758);
xor UO_1404 (O_1404,N_19437,N_18281);
nor UO_1405 (O_1405,N_18606,N_18109);
xor UO_1406 (O_1406,N_18128,N_18310);
or UO_1407 (O_1407,N_19013,N_18382);
and UO_1408 (O_1408,N_19308,N_19311);
or UO_1409 (O_1409,N_19116,N_19373);
or UO_1410 (O_1410,N_18743,N_18030);
or UO_1411 (O_1411,N_19146,N_18771);
nor UO_1412 (O_1412,N_18819,N_19410);
xor UO_1413 (O_1413,N_19912,N_18835);
nand UO_1414 (O_1414,N_18593,N_18591);
nand UO_1415 (O_1415,N_19166,N_18352);
and UO_1416 (O_1416,N_19591,N_19150);
nor UO_1417 (O_1417,N_18632,N_19876);
or UO_1418 (O_1418,N_18281,N_18465);
xnor UO_1419 (O_1419,N_19542,N_19340);
or UO_1420 (O_1420,N_18721,N_18223);
or UO_1421 (O_1421,N_18545,N_19439);
or UO_1422 (O_1422,N_18438,N_18181);
and UO_1423 (O_1423,N_19225,N_19413);
or UO_1424 (O_1424,N_19360,N_18696);
and UO_1425 (O_1425,N_18408,N_19068);
nor UO_1426 (O_1426,N_18609,N_19285);
xor UO_1427 (O_1427,N_18078,N_18770);
and UO_1428 (O_1428,N_18481,N_18767);
nor UO_1429 (O_1429,N_19024,N_18016);
and UO_1430 (O_1430,N_19435,N_19012);
and UO_1431 (O_1431,N_18596,N_19694);
nor UO_1432 (O_1432,N_18817,N_19787);
and UO_1433 (O_1433,N_19925,N_18873);
and UO_1434 (O_1434,N_19343,N_18270);
or UO_1435 (O_1435,N_19442,N_18334);
and UO_1436 (O_1436,N_19858,N_18893);
and UO_1437 (O_1437,N_19759,N_19323);
xor UO_1438 (O_1438,N_19957,N_18310);
nor UO_1439 (O_1439,N_19593,N_18710);
xnor UO_1440 (O_1440,N_18666,N_19803);
or UO_1441 (O_1441,N_18484,N_18471);
nand UO_1442 (O_1442,N_18783,N_18002);
and UO_1443 (O_1443,N_18262,N_18256);
nor UO_1444 (O_1444,N_19961,N_19805);
nor UO_1445 (O_1445,N_19180,N_18193);
nor UO_1446 (O_1446,N_19468,N_18798);
or UO_1447 (O_1447,N_18798,N_18899);
and UO_1448 (O_1448,N_18497,N_19565);
nor UO_1449 (O_1449,N_19576,N_18607);
or UO_1450 (O_1450,N_19166,N_18441);
or UO_1451 (O_1451,N_19881,N_18742);
xnor UO_1452 (O_1452,N_18917,N_19891);
and UO_1453 (O_1453,N_18672,N_18390);
nor UO_1454 (O_1454,N_18364,N_18177);
nand UO_1455 (O_1455,N_19287,N_19112);
nor UO_1456 (O_1456,N_19841,N_19218);
or UO_1457 (O_1457,N_18703,N_18749);
or UO_1458 (O_1458,N_19309,N_19375);
or UO_1459 (O_1459,N_18357,N_18450);
nor UO_1460 (O_1460,N_19035,N_19642);
xnor UO_1461 (O_1461,N_18840,N_19457);
nor UO_1462 (O_1462,N_19740,N_18783);
nand UO_1463 (O_1463,N_18010,N_19281);
xor UO_1464 (O_1464,N_18255,N_19964);
nor UO_1465 (O_1465,N_19475,N_19166);
nand UO_1466 (O_1466,N_19125,N_19483);
xnor UO_1467 (O_1467,N_18943,N_19991);
xor UO_1468 (O_1468,N_18665,N_19991);
nor UO_1469 (O_1469,N_19577,N_19984);
and UO_1470 (O_1470,N_19707,N_18211);
and UO_1471 (O_1471,N_18034,N_18155);
and UO_1472 (O_1472,N_18435,N_18650);
nand UO_1473 (O_1473,N_18193,N_18163);
or UO_1474 (O_1474,N_18827,N_19156);
nor UO_1475 (O_1475,N_19278,N_19171);
xnor UO_1476 (O_1476,N_19294,N_19457);
and UO_1477 (O_1477,N_19244,N_19400);
nor UO_1478 (O_1478,N_19039,N_18335);
nand UO_1479 (O_1479,N_18018,N_19352);
nor UO_1480 (O_1480,N_18992,N_19710);
nor UO_1481 (O_1481,N_18270,N_19939);
nor UO_1482 (O_1482,N_18223,N_18039);
or UO_1483 (O_1483,N_19535,N_18299);
and UO_1484 (O_1484,N_18717,N_19424);
nor UO_1485 (O_1485,N_19992,N_18457);
xnor UO_1486 (O_1486,N_19775,N_19554);
nor UO_1487 (O_1487,N_19999,N_18327);
xor UO_1488 (O_1488,N_19632,N_19522);
or UO_1489 (O_1489,N_18517,N_18879);
and UO_1490 (O_1490,N_18636,N_18226);
xnor UO_1491 (O_1491,N_19845,N_18713);
xnor UO_1492 (O_1492,N_19069,N_18455);
nor UO_1493 (O_1493,N_18838,N_18192);
xnor UO_1494 (O_1494,N_18042,N_18829);
and UO_1495 (O_1495,N_18498,N_19671);
or UO_1496 (O_1496,N_18572,N_18230);
nor UO_1497 (O_1497,N_19177,N_19418);
xor UO_1498 (O_1498,N_19099,N_18731);
nor UO_1499 (O_1499,N_18393,N_19000);
xor UO_1500 (O_1500,N_19570,N_18292);
and UO_1501 (O_1501,N_18073,N_18341);
nor UO_1502 (O_1502,N_19518,N_18466);
or UO_1503 (O_1503,N_18805,N_18574);
nor UO_1504 (O_1504,N_18582,N_19699);
nor UO_1505 (O_1505,N_18024,N_19448);
nor UO_1506 (O_1506,N_18992,N_18397);
xnor UO_1507 (O_1507,N_19178,N_19984);
and UO_1508 (O_1508,N_19398,N_19283);
nand UO_1509 (O_1509,N_19519,N_18622);
nor UO_1510 (O_1510,N_19126,N_18465);
nor UO_1511 (O_1511,N_19466,N_18177);
xnor UO_1512 (O_1512,N_18554,N_18502);
or UO_1513 (O_1513,N_18042,N_19742);
xnor UO_1514 (O_1514,N_19785,N_18896);
or UO_1515 (O_1515,N_18073,N_18041);
nor UO_1516 (O_1516,N_18225,N_19361);
or UO_1517 (O_1517,N_19087,N_19710);
and UO_1518 (O_1518,N_19829,N_18058);
or UO_1519 (O_1519,N_19095,N_18843);
xnor UO_1520 (O_1520,N_19187,N_19463);
nand UO_1521 (O_1521,N_19968,N_19989);
nor UO_1522 (O_1522,N_19282,N_19724);
xor UO_1523 (O_1523,N_19007,N_18732);
nor UO_1524 (O_1524,N_19211,N_18307);
xnor UO_1525 (O_1525,N_18072,N_19976);
and UO_1526 (O_1526,N_18567,N_18694);
and UO_1527 (O_1527,N_18682,N_19507);
and UO_1528 (O_1528,N_19215,N_19417);
nand UO_1529 (O_1529,N_19982,N_18681);
and UO_1530 (O_1530,N_19076,N_19027);
xor UO_1531 (O_1531,N_19033,N_18297);
xnor UO_1532 (O_1532,N_19763,N_18590);
or UO_1533 (O_1533,N_18808,N_18156);
xor UO_1534 (O_1534,N_18680,N_19239);
and UO_1535 (O_1535,N_19972,N_18938);
or UO_1536 (O_1536,N_19792,N_19819);
and UO_1537 (O_1537,N_18628,N_19084);
and UO_1538 (O_1538,N_19823,N_18949);
nand UO_1539 (O_1539,N_18230,N_19527);
or UO_1540 (O_1540,N_18861,N_19910);
and UO_1541 (O_1541,N_19388,N_19665);
and UO_1542 (O_1542,N_18734,N_19502);
nor UO_1543 (O_1543,N_18728,N_19093);
and UO_1544 (O_1544,N_18652,N_19040);
xnor UO_1545 (O_1545,N_19696,N_18262);
nor UO_1546 (O_1546,N_18666,N_19064);
and UO_1547 (O_1547,N_18675,N_18322);
nor UO_1548 (O_1548,N_19863,N_18398);
nand UO_1549 (O_1549,N_19642,N_19797);
and UO_1550 (O_1550,N_18991,N_19525);
or UO_1551 (O_1551,N_18624,N_19395);
nand UO_1552 (O_1552,N_18408,N_19081);
and UO_1553 (O_1553,N_19316,N_18683);
and UO_1554 (O_1554,N_19563,N_19120);
and UO_1555 (O_1555,N_18426,N_19316);
nor UO_1556 (O_1556,N_19023,N_19483);
or UO_1557 (O_1557,N_19491,N_18525);
and UO_1558 (O_1558,N_19498,N_18891);
or UO_1559 (O_1559,N_19534,N_18603);
xor UO_1560 (O_1560,N_19232,N_19196);
nor UO_1561 (O_1561,N_18074,N_18336);
or UO_1562 (O_1562,N_19923,N_18990);
or UO_1563 (O_1563,N_18740,N_19206);
and UO_1564 (O_1564,N_19428,N_19613);
nand UO_1565 (O_1565,N_18875,N_19505);
xnor UO_1566 (O_1566,N_19480,N_19125);
nor UO_1567 (O_1567,N_19381,N_18074);
nor UO_1568 (O_1568,N_18334,N_18802);
nor UO_1569 (O_1569,N_18142,N_19365);
xnor UO_1570 (O_1570,N_18055,N_18291);
nor UO_1571 (O_1571,N_19778,N_19404);
nand UO_1572 (O_1572,N_18466,N_19532);
nand UO_1573 (O_1573,N_18639,N_19499);
and UO_1574 (O_1574,N_18339,N_18492);
or UO_1575 (O_1575,N_19698,N_18976);
and UO_1576 (O_1576,N_18238,N_18340);
nor UO_1577 (O_1577,N_18111,N_19268);
or UO_1578 (O_1578,N_18548,N_18616);
nand UO_1579 (O_1579,N_19600,N_18285);
nand UO_1580 (O_1580,N_19211,N_19207);
or UO_1581 (O_1581,N_18832,N_19804);
and UO_1582 (O_1582,N_18158,N_18558);
nand UO_1583 (O_1583,N_19455,N_18944);
nand UO_1584 (O_1584,N_19745,N_19090);
and UO_1585 (O_1585,N_19436,N_18968);
nor UO_1586 (O_1586,N_19446,N_19899);
nand UO_1587 (O_1587,N_19650,N_18321);
xnor UO_1588 (O_1588,N_18214,N_19168);
or UO_1589 (O_1589,N_18037,N_19381);
or UO_1590 (O_1590,N_19338,N_18933);
or UO_1591 (O_1591,N_19695,N_18104);
and UO_1592 (O_1592,N_18344,N_18547);
and UO_1593 (O_1593,N_18480,N_18953);
xnor UO_1594 (O_1594,N_18753,N_18608);
nor UO_1595 (O_1595,N_18590,N_19822);
and UO_1596 (O_1596,N_18086,N_19207);
and UO_1597 (O_1597,N_19666,N_19735);
nor UO_1598 (O_1598,N_18681,N_19449);
nor UO_1599 (O_1599,N_18500,N_19859);
nor UO_1600 (O_1600,N_18600,N_18260);
or UO_1601 (O_1601,N_18862,N_19711);
and UO_1602 (O_1602,N_18180,N_19009);
nand UO_1603 (O_1603,N_18743,N_18696);
or UO_1604 (O_1604,N_18731,N_18523);
xnor UO_1605 (O_1605,N_19047,N_18406);
and UO_1606 (O_1606,N_18957,N_19248);
nor UO_1607 (O_1607,N_18063,N_19286);
and UO_1608 (O_1608,N_18751,N_18006);
or UO_1609 (O_1609,N_18633,N_18083);
nor UO_1610 (O_1610,N_18178,N_18493);
or UO_1611 (O_1611,N_19660,N_18510);
nor UO_1612 (O_1612,N_18851,N_19626);
or UO_1613 (O_1613,N_19847,N_18996);
nor UO_1614 (O_1614,N_18362,N_19123);
and UO_1615 (O_1615,N_18637,N_18779);
nor UO_1616 (O_1616,N_18949,N_18005);
xnor UO_1617 (O_1617,N_19846,N_18889);
nand UO_1618 (O_1618,N_19315,N_19895);
and UO_1619 (O_1619,N_18992,N_19383);
nand UO_1620 (O_1620,N_19335,N_19198);
nand UO_1621 (O_1621,N_18952,N_18581);
xnor UO_1622 (O_1622,N_19931,N_18848);
or UO_1623 (O_1623,N_18145,N_19154);
and UO_1624 (O_1624,N_19084,N_18940);
and UO_1625 (O_1625,N_19237,N_18118);
and UO_1626 (O_1626,N_18261,N_18353);
xor UO_1627 (O_1627,N_19487,N_18445);
nand UO_1628 (O_1628,N_19523,N_18359);
xor UO_1629 (O_1629,N_19489,N_19726);
or UO_1630 (O_1630,N_19869,N_19209);
and UO_1631 (O_1631,N_19074,N_18129);
or UO_1632 (O_1632,N_18191,N_19879);
nand UO_1633 (O_1633,N_19804,N_18210);
and UO_1634 (O_1634,N_18423,N_19155);
or UO_1635 (O_1635,N_18427,N_19659);
or UO_1636 (O_1636,N_19044,N_18402);
xnor UO_1637 (O_1637,N_19540,N_19992);
nand UO_1638 (O_1638,N_19832,N_18893);
xnor UO_1639 (O_1639,N_18653,N_18487);
or UO_1640 (O_1640,N_19560,N_18253);
xnor UO_1641 (O_1641,N_19603,N_18216);
nor UO_1642 (O_1642,N_19153,N_19128);
xor UO_1643 (O_1643,N_19876,N_18587);
and UO_1644 (O_1644,N_19880,N_19208);
nor UO_1645 (O_1645,N_18080,N_19001);
xnor UO_1646 (O_1646,N_19793,N_19468);
nand UO_1647 (O_1647,N_18967,N_19700);
nor UO_1648 (O_1648,N_18659,N_19389);
and UO_1649 (O_1649,N_19908,N_18411);
nand UO_1650 (O_1650,N_18535,N_19589);
nor UO_1651 (O_1651,N_19385,N_18774);
nor UO_1652 (O_1652,N_18317,N_18841);
xnor UO_1653 (O_1653,N_19409,N_19474);
and UO_1654 (O_1654,N_19539,N_18760);
or UO_1655 (O_1655,N_18469,N_19841);
or UO_1656 (O_1656,N_19434,N_19009);
and UO_1657 (O_1657,N_19886,N_19155);
nor UO_1658 (O_1658,N_18658,N_19542);
and UO_1659 (O_1659,N_19960,N_18906);
nor UO_1660 (O_1660,N_18350,N_18213);
or UO_1661 (O_1661,N_19600,N_18818);
nor UO_1662 (O_1662,N_19248,N_18857);
nand UO_1663 (O_1663,N_19313,N_19551);
or UO_1664 (O_1664,N_18863,N_18979);
nor UO_1665 (O_1665,N_18673,N_18148);
nor UO_1666 (O_1666,N_18632,N_18410);
nor UO_1667 (O_1667,N_19443,N_19026);
nor UO_1668 (O_1668,N_18521,N_18311);
and UO_1669 (O_1669,N_18747,N_19553);
xor UO_1670 (O_1670,N_18889,N_18961);
xor UO_1671 (O_1671,N_19049,N_19913);
nand UO_1672 (O_1672,N_19760,N_19349);
nor UO_1673 (O_1673,N_19799,N_19699);
nor UO_1674 (O_1674,N_18228,N_19820);
xor UO_1675 (O_1675,N_19863,N_18525);
nand UO_1676 (O_1676,N_19216,N_19127);
nor UO_1677 (O_1677,N_18157,N_18380);
xnor UO_1678 (O_1678,N_19409,N_19415);
and UO_1679 (O_1679,N_18599,N_19991);
nand UO_1680 (O_1680,N_19602,N_18631);
or UO_1681 (O_1681,N_18899,N_19069);
and UO_1682 (O_1682,N_18435,N_19531);
and UO_1683 (O_1683,N_18136,N_19494);
xor UO_1684 (O_1684,N_18070,N_18498);
nand UO_1685 (O_1685,N_18006,N_18944);
xor UO_1686 (O_1686,N_19257,N_18441);
nand UO_1687 (O_1687,N_19324,N_19407);
nand UO_1688 (O_1688,N_19393,N_18344);
xnor UO_1689 (O_1689,N_18686,N_19123);
and UO_1690 (O_1690,N_19471,N_18813);
or UO_1691 (O_1691,N_18028,N_19785);
and UO_1692 (O_1692,N_19897,N_18042);
and UO_1693 (O_1693,N_18193,N_18706);
xor UO_1694 (O_1694,N_18761,N_18714);
and UO_1695 (O_1695,N_19059,N_19867);
xnor UO_1696 (O_1696,N_18096,N_19366);
nor UO_1697 (O_1697,N_19955,N_18891);
xnor UO_1698 (O_1698,N_19636,N_18687);
and UO_1699 (O_1699,N_19688,N_19468);
nand UO_1700 (O_1700,N_19187,N_18943);
nand UO_1701 (O_1701,N_19513,N_19687);
nand UO_1702 (O_1702,N_19708,N_19979);
xnor UO_1703 (O_1703,N_18187,N_19982);
xor UO_1704 (O_1704,N_18195,N_18005);
or UO_1705 (O_1705,N_19902,N_18756);
nand UO_1706 (O_1706,N_18075,N_18909);
and UO_1707 (O_1707,N_19613,N_19442);
and UO_1708 (O_1708,N_18523,N_19716);
xnor UO_1709 (O_1709,N_19725,N_18715);
or UO_1710 (O_1710,N_19323,N_18201);
xor UO_1711 (O_1711,N_19999,N_18231);
and UO_1712 (O_1712,N_19894,N_18710);
or UO_1713 (O_1713,N_19467,N_19300);
or UO_1714 (O_1714,N_19869,N_19366);
or UO_1715 (O_1715,N_19078,N_19509);
or UO_1716 (O_1716,N_18852,N_18411);
nor UO_1717 (O_1717,N_19682,N_18104);
or UO_1718 (O_1718,N_18759,N_18829);
nand UO_1719 (O_1719,N_18994,N_19142);
or UO_1720 (O_1720,N_19741,N_18777);
and UO_1721 (O_1721,N_19636,N_19817);
and UO_1722 (O_1722,N_18648,N_19411);
nor UO_1723 (O_1723,N_18023,N_18661);
and UO_1724 (O_1724,N_18566,N_18530);
nor UO_1725 (O_1725,N_18387,N_18401);
xor UO_1726 (O_1726,N_18386,N_18121);
or UO_1727 (O_1727,N_19520,N_19788);
xor UO_1728 (O_1728,N_19380,N_18166);
xnor UO_1729 (O_1729,N_18932,N_19416);
and UO_1730 (O_1730,N_19813,N_18398);
and UO_1731 (O_1731,N_19410,N_18942);
and UO_1732 (O_1732,N_18051,N_19047);
nand UO_1733 (O_1733,N_18365,N_19117);
and UO_1734 (O_1734,N_18333,N_18900);
xor UO_1735 (O_1735,N_19765,N_18208);
nand UO_1736 (O_1736,N_19304,N_19399);
nor UO_1737 (O_1737,N_18561,N_19883);
or UO_1738 (O_1738,N_18636,N_19718);
xor UO_1739 (O_1739,N_19950,N_19061);
nand UO_1740 (O_1740,N_19877,N_19082);
nand UO_1741 (O_1741,N_19815,N_18202);
or UO_1742 (O_1742,N_18137,N_18831);
nor UO_1743 (O_1743,N_19415,N_19898);
nor UO_1744 (O_1744,N_18611,N_18733);
and UO_1745 (O_1745,N_18115,N_19015);
xnor UO_1746 (O_1746,N_19680,N_19314);
nor UO_1747 (O_1747,N_18846,N_18844);
nand UO_1748 (O_1748,N_19738,N_19044);
or UO_1749 (O_1749,N_19238,N_18498);
xnor UO_1750 (O_1750,N_19883,N_18280);
nor UO_1751 (O_1751,N_18434,N_18375);
and UO_1752 (O_1752,N_19020,N_18990);
and UO_1753 (O_1753,N_18310,N_19201);
or UO_1754 (O_1754,N_19935,N_19407);
nand UO_1755 (O_1755,N_19352,N_19146);
nand UO_1756 (O_1756,N_19107,N_18093);
nand UO_1757 (O_1757,N_18985,N_19612);
or UO_1758 (O_1758,N_18262,N_19407);
and UO_1759 (O_1759,N_19586,N_19801);
nor UO_1760 (O_1760,N_18574,N_18186);
xnor UO_1761 (O_1761,N_18010,N_19083);
nor UO_1762 (O_1762,N_18112,N_18412);
xor UO_1763 (O_1763,N_19528,N_19511);
nand UO_1764 (O_1764,N_19869,N_19999);
or UO_1765 (O_1765,N_18502,N_19378);
nor UO_1766 (O_1766,N_18933,N_18664);
nor UO_1767 (O_1767,N_18522,N_19335);
xor UO_1768 (O_1768,N_19250,N_19461);
or UO_1769 (O_1769,N_19750,N_18426);
or UO_1770 (O_1770,N_19625,N_19924);
xor UO_1771 (O_1771,N_19201,N_18729);
xnor UO_1772 (O_1772,N_18989,N_19058);
or UO_1773 (O_1773,N_18396,N_19760);
nand UO_1774 (O_1774,N_19914,N_18496);
nor UO_1775 (O_1775,N_19971,N_18087);
and UO_1776 (O_1776,N_18920,N_19568);
nand UO_1777 (O_1777,N_18124,N_18084);
nand UO_1778 (O_1778,N_19824,N_18319);
xor UO_1779 (O_1779,N_18357,N_19340);
nand UO_1780 (O_1780,N_18214,N_18740);
and UO_1781 (O_1781,N_18944,N_19325);
nor UO_1782 (O_1782,N_18621,N_18316);
nand UO_1783 (O_1783,N_19360,N_19454);
and UO_1784 (O_1784,N_18121,N_19268);
xor UO_1785 (O_1785,N_18713,N_18863);
xnor UO_1786 (O_1786,N_19522,N_19071);
nand UO_1787 (O_1787,N_19851,N_18675);
nand UO_1788 (O_1788,N_18046,N_19662);
xor UO_1789 (O_1789,N_18880,N_18681);
or UO_1790 (O_1790,N_19411,N_18833);
nor UO_1791 (O_1791,N_18336,N_18733);
xor UO_1792 (O_1792,N_19347,N_18798);
or UO_1793 (O_1793,N_19354,N_19594);
nand UO_1794 (O_1794,N_18220,N_19047);
xor UO_1795 (O_1795,N_19447,N_18483);
or UO_1796 (O_1796,N_18175,N_19574);
nand UO_1797 (O_1797,N_18056,N_19201);
xnor UO_1798 (O_1798,N_19580,N_18630);
nand UO_1799 (O_1799,N_18284,N_19391);
or UO_1800 (O_1800,N_19615,N_18996);
xor UO_1801 (O_1801,N_19533,N_19090);
nand UO_1802 (O_1802,N_18746,N_19106);
xor UO_1803 (O_1803,N_18320,N_18852);
or UO_1804 (O_1804,N_19275,N_19364);
and UO_1805 (O_1805,N_19024,N_18688);
and UO_1806 (O_1806,N_18063,N_19678);
or UO_1807 (O_1807,N_19600,N_18463);
or UO_1808 (O_1808,N_18795,N_19153);
and UO_1809 (O_1809,N_18745,N_18927);
nand UO_1810 (O_1810,N_18978,N_18404);
and UO_1811 (O_1811,N_18009,N_19057);
nor UO_1812 (O_1812,N_18823,N_18440);
xnor UO_1813 (O_1813,N_19631,N_18185);
nand UO_1814 (O_1814,N_19065,N_19327);
nor UO_1815 (O_1815,N_18370,N_18890);
nand UO_1816 (O_1816,N_19291,N_19140);
xnor UO_1817 (O_1817,N_19234,N_18748);
and UO_1818 (O_1818,N_19910,N_19270);
or UO_1819 (O_1819,N_18747,N_19452);
nor UO_1820 (O_1820,N_19102,N_18293);
nor UO_1821 (O_1821,N_18552,N_19451);
nor UO_1822 (O_1822,N_19921,N_18348);
nand UO_1823 (O_1823,N_18972,N_19654);
or UO_1824 (O_1824,N_18210,N_19749);
nor UO_1825 (O_1825,N_19604,N_19067);
nor UO_1826 (O_1826,N_19147,N_18733);
nand UO_1827 (O_1827,N_18307,N_18106);
and UO_1828 (O_1828,N_19984,N_19307);
nor UO_1829 (O_1829,N_19755,N_18011);
nand UO_1830 (O_1830,N_19973,N_19999);
and UO_1831 (O_1831,N_18733,N_19394);
xor UO_1832 (O_1832,N_18284,N_19199);
xnor UO_1833 (O_1833,N_19524,N_18533);
or UO_1834 (O_1834,N_19128,N_18184);
or UO_1835 (O_1835,N_19836,N_19095);
and UO_1836 (O_1836,N_18810,N_18212);
nor UO_1837 (O_1837,N_18095,N_19933);
or UO_1838 (O_1838,N_18289,N_19417);
nor UO_1839 (O_1839,N_18104,N_18612);
nor UO_1840 (O_1840,N_18346,N_19082);
xnor UO_1841 (O_1841,N_18580,N_19514);
nand UO_1842 (O_1842,N_19923,N_19509);
xor UO_1843 (O_1843,N_18264,N_19388);
nor UO_1844 (O_1844,N_19703,N_18853);
and UO_1845 (O_1845,N_19360,N_19101);
and UO_1846 (O_1846,N_18018,N_18163);
and UO_1847 (O_1847,N_18875,N_19612);
nor UO_1848 (O_1848,N_19275,N_19552);
and UO_1849 (O_1849,N_19620,N_18939);
nand UO_1850 (O_1850,N_18471,N_19716);
nor UO_1851 (O_1851,N_19613,N_19423);
nand UO_1852 (O_1852,N_18538,N_19776);
or UO_1853 (O_1853,N_18935,N_18046);
xnor UO_1854 (O_1854,N_19082,N_19935);
and UO_1855 (O_1855,N_19725,N_18747);
nand UO_1856 (O_1856,N_19915,N_19751);
nand UO_1857 (O_1857,N_19116,N_18810);
or UO_1858 (O_1858,N_18428,N_18041);
or UO_1859 (O_1859,N_19996,N_19130);
nand UO_1860 (O_1860,N_18502,N_19723);
or UO_1861 (O_1861,N_18656,N_18029);
or UO_1862 (O_1862,N_19955,N_18005);
or UO_1863 (O_1863,N_18697,N_18968);
and UO_1864 (O_1864,N_18343,N_19509);
nor UO_1865 (O_1865,N_18797,N_18357);
or UO_1866 (O_1866,N_18694,N_19178);
nand UO_1867 (O_1867,N_19744,N_19395);
xor UO_1868 (O_1868,N_19670,N_18869);
xor UO_1869 (O_1869,N_19620,N_19392);
xnor UO_1870 (O_1870,N_19569,N_19615);
nor UO_1871 (O_1871,N_18389,N_19509);
xnor UO_1872 (O_1872,N_18173,N_18927);
nand UO_1873 (O_1873,N_19322,N_19079);
nor UO_1874 (O_1874,N_19935,N_19693);
nor UO_1875 (O_1875,N_19078,N_18551);
nand UO_1876 (O_1876,N_19250,N_19414);
xnor UO_1877 (O_1877,N_19222,N_19484);
xor UO_1878 (O_1878,N_19105,N_19853);
nor UO_1879 (O_1879,N_19415,N_19712);
nand UO_1880 (O_1880,N_19993,N_18347);
and UO_1881 (O_1881,N_18315,N_19306);
nor UO_1882 (O_1882,N_19740,N_19802);
or UO_1883 (O_1883,N_18751,N_19717);
nand UO_1884 (O_1884,N_19734,N_19888);
nand UO_1885 (O_1885,N_19395,N_19637);
and UO_1886 (O_1886,N_18465,N_18325);
and UO_1887 (O_1887,N_18729,N_19174);
nor UO_1888 (O_1888,N_19044,N_19158);
nand UO_1889 (O_1889,N_18865,N_18593);
or UO_1890 (O_1890,N_18184,N_19488);
or UO_1891 (O_1891,N_18649,N_18876);
nor UO_1892 (O_1892,N_18628,N_19773);
nor UO_1893 (O_1893,N_19200,N_18190);
or UO_1894 (O_1894,N_19844,N_18753);
nand UO_1895 (O_1895,N_18613,N_19635);
nor UO_1896 (O_1896,N_18115,N_19400);
and UO_1897 (O_1897,N_19345,N_19863);
or UO_1898 (O_1898,N_18724,N_18576);
nand UO_1899 (O_1899,N_19666,N_18042);
or UO_1900 (O_1900,N_18191,N_19172);
nor UO_1901 (O_1901,N_19021,N_19399);
nand UO_1902 (O_1902,N_18273,N_18791);
nand UO_1903 (O_1903,N_18185,N_18976);
nand UO_1904 (O_1904,N_18713,N_19710);
and UO_1905 (O_1905,N_18846,N_19933);
and UO_1906 (O_1906,N_18798,N_19456);
or UO_1907 (O_1907,N_19582,N_19837);
xor UO_1908 (O_1908,N_18710,N_18123);
nor UO_1909 (O_1909,N_18337,N_18832);
nand UO_1910 (O_1910,N_19785,N_19404);
and UO_1911 (O_1911,N_19031,N_18330);
xor UO_1912 (O_1912,N_18429,N_18996);
xnor UO_1913 (O_1913,N_19238,N_18549);
and UO_1914 (O_1914,N_18569,N_19649);
and UO_1915 (O_1915,N_19246,N_18139);
nor UO_1916 (O_1916,N_19447,N_19257);
xor UO_1917 (O_1917,N_18794,N_19082);
or UO_1918 (O_1918,N_18079,N_19048);
nand UO_1919 (O_1919,N_19716,N_18300);
nand UO_1920 (O_1920,N_19402,N_18404);
xor UO_1921 (O_1921,N_19536,N_19069);
nor UO_1922 (O_1922,N_18578,N_18841);
nor UO_1923 (O_1923,N_19969,N_18071);
nor UO_1924 (O_1924,N_19748,N_19591);
nand UO_1925 (O_1925,N_18443,N_18315);
nand UO_1926 (O_1926,N_19885,N_19299);
and UO_1927 (O_1927,N_19123,N_19896);
or UO_1928 (O_1928,N_18169,N_19253);
xor UO_1929 (O_1929,N_19736,N_19636);
or UO_1930 (O_1930,N_19544,N_19803);
xor UO_1931 (O_1931,N_19599,N_19751);
and UO_1932 (O_1932,N_18542,N_19876);
or UO_1933 (O_1933,N_18965,N_18121);
xnor UO_1934 (O_1934,N_19982,N_18133);
nor UO_1935 (O_1935,N_19550,N_18879);
nand UO_1936 (O_1936,N_18205,N_18042);
and UO_1937 (O_1937,N_19958,N_18846);
and UO_1938 (O_1938,N_18647,N_19669);
xnor UO_1939 (O_1939,N_18121,N_19313);
or UO_1940 (O_1940,N_18301,N_19085);
xor UO_1941 (O_1941,N_18167,N_19407);
and UO_1942 (O_1942,N_18932,N_18702);
or UO_1943 (O_1943,N_19253,N_19746);
and UO_1944 (O_1944,N_18815,N_19060);
nand UO_1945 (O_1945,N_19167,N_18940);
and UO_1946 (O_1946,N_19625,N_18667);
or UO_1947 (O_1947,N_19525,N_18700);
nand UO_1948 (O_1948,N_18767,N_19807);
or UO_1949 (O_1949,N_18919,N_18668);
nand UO_1950 (O_1950,N_19722,N_19721);
or UO_1951 (O_1951,N_18659,N_18132);
nor UO_1952 (O_1952,N_18506,N_19426);
or UO_1953 (O_1953,N_18213,N_19984);
xor UO_1954 (O_1954,N_19862,N_18418);
and UO_1955 (O_1955,N_19254,N_19442);
xor UO_1956 (O_1956,N_19297,N_18841);
or UO_1957 (O_1957,N_19337,N_18549);
and UO_1958 (O_1958,N_18992,N_18174);
xnor UO_1959 (O_1959,N_18797,N_19279);
and UO_1960 (O_1960,N_18520,N_18217);
nor UO_1961 (O_1961,N_18548,N_18686);
and UO_1962 (O_1962,N_19550,N_19233);
nand UO_1963 (O_1963,N_19794,N_19427);
or UO_1964 (O_1964,N_18266,N_18691);
or UO_1965 (O_1965,N_18136,N_19566);
or UO_1966 (O_1966,N_19256,N_18067);
nand UO_1967 (O_1967,N_19605,N_19858);
xnor UO_1968 (O_1968,N_19161,N_19312);
xor UO_1969 (O_1969,N_18195,N_18072);
xor UO_1970 (O_1970,N_19477,N_18029);
nand UO_1971 (O_1971,N_18439,N_19057);
or UO_1972 (O_1972,N_18976,N_18849);
nand UO_1973 (O_1973,N_18647,N_19027);
and UO_1974 (O_1974,N_19620,N_19450);
or UO_1975 (O_1975,N_19615,N_19299);
or UO_1976 (O_1976,N_18317,N_18742);
nand UO_1977 (O_1977,N_18259,N_19515);
and UO_1978 (O_1978,N_18554,N_18691);
nand UO_1979 (O_1979,N_19384,N_19986);
nor UO_1980 (O_1980,N_19968,N_18522);
nor UO_1981 (O_1981,N_18078,N_19273);
xor UO_1982 (O_1982,N_19866,N_18322);
nand UO_1983 (O_1983,N_18844,N_18067);
and UO_1984 (O_1984,N_19740,N_19931);
xnor UO_1985 (O_1985,N_18259,N_18836);
and UO_1986 (O_1986,N_18984,N_18982);
nand UO_1987 (O_1987,N_19534,N_19456);
nor UO_1988 (O_1988,N_18056,N_18016);
and UO_1989 (O_1989,N_18561,N_18197);
nor UO_1990 (O_1990,N_19485,N_19979);
xnor UO_1991 (O_1991,N_19284,N_18774);
xor UO_1992 (O_1992,N_19786,N_19716);
nor UO_1993 (O_1993,N_18101,N_18402);
nand UO_1994 (O_1994,N_19546,N_19406);
xor UO_1995 (O_1995,N_18027,N_18757);
or UO_1996 (O_1996,N_19276,N_19475);
xor UO_1997 (O_1997,N_18346,N_19102);
nor UO_1998 (O_1998,N_19073,N_18626);
or UO_1999 (O_1999,N_19354,N_19269);
and UO_2000 (O_2000,N_19832,N_18544);
nor UO_2001 (O_2001,N_19458,N_19135);
xor UO_2002 (O_2002,N_18845,N_19143);
or UO_2003 (O_2003,N_19965,N_19960);
xnor UO_2004 (O_2004,N_18934,N_18840);
nand UO_2005 (O_2005,N_18114,N_19847);
nand UO_2006 (O_2006,N_18610,N_18488);
nor UO_2007 (O_2007,N_18752,N_19900);
nor UO_2008 (O_2008,N_18456,N_19321);
xor UO_2009 (O_2009,N_19265,N_19897);
nand UO_2010 (O_2010,N_18942,N_18460);
nand UO_2011 (O_2011,N_18957,N_19510);
nor UO_2012 (O_2012,N_19021,N_18072);
or UO_2013 (O_2013,N_19699,N_19106);
or UO_2014 (O_2014,N_18196,N_19527);
and UO_2015 (O_2015,N_18147,N_18675);
and UO_2016 (O_2016,N_19344,N_18088);
or UO_2017 (O_2017,N_19425,N_18038);
or UO_2018 (O_2018,N_18564,N_19502);
nor UO_2019 (O_2019,N_18852,N_18948);
or UO_2020 (O_2020,N_19869,N_19259);
and UO_2021 (O_2021,N_18471,N_18584);
or UO_2022 (O_2022,N_18276,N_18054);
nand UO_2023 (O_2023,N_19918,N_18475);
and UO_2024 (O_2024,N_18832,N_18601);
nor UO_2025 (O_2025,N_18581,N_19006);
or UO_2026 (O_2026,N_19278,N_18459);
nor UO_2027 (O_2027,N_18907,N_18941);
or UO_2028 (O_2028,N_19827,N_18426);
nand UO_2029 (O_2029,N_18802,N_18057);
nand UO_2030 (O_2030,N_18974,N_18638);
nand UO_2031 (O_2031,N_19033,N_18712);
nor UO_2032 (O_2032,N_18169,N_19462);
xnor UO_2033 (O_2033,N_18557,N_19553);
nand UO_2034 (O_2034,N_18090,N_19579);
xnor UO_2035 (O_2035,N_18976,N_18479);
nand UO_2036 (O_2036,N_19584,N_19912);
nand UO_2037 (O_2037,N_19131,N_19493);
and UO_2038 (O_2038,N_18264,N_19440);
nand UO_2039 (O_2039,N_18873,N_19003);
nand UO_2040 (O_2040,N_19736,N_18778);
nand UO_2041 (O_2041,N_18472,N_18618);
nand UO_2042 (O_2042,N_18102,N_19192);
nor UO_2043 (O_2043,N_19361,N_18247);
or UO_2044 (O_2044,N_19793,N_19210);
nand UO_2045 (O_2045,N_18862,N_19198);
nor UO_2046 (O_2046,N_18183,N_18787);
nor UO_2047 (O_2047,N_19115,N_19265);
nand UO_2048 (O_2048,N_18005,N_18484);
nand UO_2049 (O_2049,N_18567,N_18033);
and UO_2050 (O_2050,N_18185,N_18689);
nor UO_2051 (O_2051,N_19843,N_18935);
nand UO_2052 (O_2052,N_18513,N_19366);
nor UO_2053 (O_2053,N_19439,N_18505);
nand UO_2054 (O_2054,N_19014,N_19159);
xnor UO_2055 (O_2055,N_18031,N_19434);
or UO_2056 (O_2056,N_19425,N_18935);
and UO_2057 (O_2057,N_18879,N_19057);
xnor UO_2058 (O_2058,N_18114,N_19208);
xnor UO_2059 (O_2059,N_18854,N_18617);
or UO_2060 (O_2060,N_19361,N_18021);
nand UO_2061 (O_2061,N_18218,N_18398);
or UO_2062 (O_2062,N_18088,N_19297);
nor UO_2063 (O_2063,N_18648,N_18229);
nand UO_2064 (O_2064,N_18023,N_18339);
nor UO_2065 (O_2065,N_18973,N_18232);
and UO_2066 (O_2066,N_18233,N_19114);
or UO_2067 (O_2067,N_18081,N_18966);
xnor UO_2068 (O_2068,N_19460,N_18169);
xnor UO_2069 (O_2069,N_18558,N_19812);
nand UO_2070 (O_2070,N_18527,N_19918);
or UO_2071 (O_2071,N_18903,N_19645);
xor UO_2072 (O_2072,N_18749,N_19622);
or UO_2073 (O_2073,N_19169,N_19870);
nand UO_2074 (O_2074,N_19127,N_19902);
nor UO_2075 (O_2075,N_19402,N_18142);
and UO_2076 (O_2076,N_18352,N_19252);
xor UO_2077 (O_2077,N_19200,N_19748);
xnor UO_2078 (O_2078,N_18650,N_19843);
nand UO_2079 (O_2079,N_18195,N_18052);
and UO_2080 (O_2080,N_19918,N_19139);
nor UO_2081 (O_2081,N_19763,N_18880);
nor UO_2082 (O_2082,N_18767,N_19474);
nand UO_2083 (O_2083,N_19542,N_19775);
xnor UO_2084 (O_2084,N_18816,N_18390);
and UO_2085 (O_2085,N_19289,N_18446);
nor UO_2086 (O_2086,N_19578,N_19697);
nand UO_2087 (O_2087,N_18693,N_19145);
nor UO_2088 (O_2088,N_19741,N_19320);
or UO_2089 (O_2089,N_18824,N_19918);
and UO_2090 (O_2090,N_18725,N_18542);
xnor UO_2091 (O_2091,N_18079,N_19300);
nor UO_2092 (O_2092,N_19021,N_18209);
or UO_2093 (O_2093,N_18960,N_18452);
nand UO_2094 (O_2094,N_19464,N_18555);
nand UO_2095 (O_2095,N_18531,N_19803);
nand UO_2096 (O_2096,N_19675,N_19131);
xor UO_2097 (O_2097,N_19902,N_19099);
nor UO_2098 (O_2098,N_19187,N_19306);
xor UO_2099 (O_2099,N_19780,N_19783);
nand UO_2100 (O_2100,N_18892,N_18186);
and UO_2101 (O_2101,N_18686,N_18635);
xnor UO_2102 (O_2102,N_18547,N_19035);
nand UO_2103 (O_2103,N_18809,N_19633);
nand UO_2104 (O_2104,N_18137,N_19568);
xnor UO_2105 (O_2105,N_18280,N_19636);
or UO_2106 (O_2106,N_18626,N_18080);
xor UO_2107 (O_2107,N_19943,N_19179);
xor UO_2108 (O_2108,N_19008,N_18700);
nand UO_2109 (O_2109,N_18899,N_19486);
and UO_2110 (O_2110,N_19177,N_19000);
nand UO_2111 (O_2111,N_19888,N_19553);
nand UO_2112 (O_2112,N_19508,N_19644);
nor UO_2113 (O_2113,N_19848,N_18141);
and UO_2114 (O_2114,N_19478,N_19580);
xor UO_2115 (O_2115,N_19288,N_18053);
or UO_2116 (O_2116,N_19097,N_19079);
and UO_2117 (O_2117,N_19957,N_18941);
nand UO_2118 (O_2118,N_18640,N_19049);
xor UO_2119 (O_2119,N_18038,N_19479);
or UO_2120 (O_2120,N_19174,N_19983);
nor UO_2121 (O_2121,N_18840,N_18740);
or UO_2122 (O_2122,N_19889,N_18202);
xnor UO_2123 (O_2123,N_18117,N_19194);
and UO_2124 (O_2124,N_19108,N_18041);
xnor UO_2125 (O_2125,N_18535,N_18024);
nand UO_2126 (O_2126,N_19599,N_19898);
or UO_2127 (O_2127,N_19780,N_19059);
or UO_2128 (O_2128,N_18524,N_18715);
and UO_2129 (O_2129,N_19054,N_18420);
nand UO_2130 (O_2130,N_19028,N_19445);
or UO_2131 (O_2131,N_19460,N_18683);
nand UO_2132 (O_2132,N_18961,N_18094);
or UO_2133 (O_2133,N_19962,N_18056);
xnor UO_2134 (O_2134,N_19749,N_19431);
or UO_2135 (O_2135,N_19093,N_18040);
and UO_2136 (O_2136,N_19590,N_19088);
and UO_2137 (O_2137,N_19894,N_18099);
and UO_2138 (O_2138,N_18750,N_19128);
or UO_2139 (O_2139,N_19397,N_18550);
nor UO_2140 (O_2140,N_19028,N_19355);
and UO_2141 (O_2141,N_19057,N_19150);
or UO_2142 (O_2142,N_18558,N_19552);
nor UO_2143 (O_2143,N_19582,N_18600);
nor UO_2144 (O_2144,N_18907,N_19437);
xor UO_2145 (O_2145,N_18196,N_18954);
nand UO_2146 (O_2146,N_19441,N_19729);
and UO_2147 (O_2147,N_19137,N_19414);
or UO_2148 (O_2148,N_18323,N_19128);
nand UO_2149 (O_2149,N_18093,N_19795);
nand UO_2150 (O_2150,N_18782,N_18706);
and UO_2151 (O_2151,N_18434,N_18685);
nor UO_2152 (O_2152,N_19990,N_18686);
nor UO_2153 (O_2153,N_18350,N_18033);
nor UO_2154 (O_2154,N_19912,N_18694);
and UO_2155 (O_2155,N_19277,N_19204);
or UO_2156 (O_2156,N_18821,N_19908);
or UO_2157 (O_2157,N_19899,N_18962);
or UO_2158 (O_2158,N_19382,N_18196);
xor UO_2159 (O_2159,N_19174,N_18462);
nor UO_2160 (O_2160,N_18152,N_18001);
or UO_2161 (O_2161,N_18597,N_19957);
xor UO_2162 (O_2162,N_19555,N_18418);
xnor UO_2163 (O_2163,N_18580,N_19786);
and UO_2164 (O_2164,N_19171,N_19123);
xor UO_2165 (O_2165,N_19260,N_18424);
and UO_2166 (O_2166,N_19318,N_19900);
and UO_2167 (O_2167,N_19497,N_19239);
or UO_2168 (O_2168,N_18435,N_19243);
nor UO_2169 (O_2169,N_19956,N_18065);
or UO_2170 (O_2170,N_19925,N_19842);
nor UO_2171 (O_2171,N_18991,N_18941);
nand UO_2172 (O_2172,N_18323,N_18168);
and UO_2173 (O_2173,N_19957,N_18434);
or UO_2174 (O_2174,N_19865,N_19361);
xnor UO_2175 (O_2175,N_19164,N_18115);
nand UO_2176 (O_2176,N_19342,N_19647);
and UO_2177 (O_2177,N_18150,N_18546);
nor UO_2178 (O_2178,N_19413,N_19952);
and UO_2179 (O_2179,N_18267,N_18684);
nor UO_2180 (O_2180,N_19707,N_19272);
nand UO_2181 (O_2181,N_19166,N_18366);
xor UO_2182 (O_2182,N_19567,N_19934);
nor UO_2183 (O_2183,N_18872,N_18897);
nand UO_2184 (O_2184,N_18832,N_18854);
nor UO_2185 (O_2185,N_18760,N_19194);
nor UO_2186 (O_2186,N_18494,N_19724);
nor UO_2187 (O_2187,N_18713,N_18004);
and UO_2188 (O_2188,N_18559,N_18642);
xnor UO_2189 (O_2189,N_18701,N_18725);
nor UO_2190 (O_2190,N_19414,N_18540);
or UO_2191 (O_2191,N_19456,N_18549);
and UO_2192 (O_2192,N_19488,N_19316);
xor UO_2193 (O_2193,N_18809,N_18632);
or UO_2194 (O_2194,N_18192,N_19833);
xor UO_2195 (O_2195,N_19743,N_18901);
nand UO_2196 (O_2196,N_18337,N_19574);
nor UO_2197 (O_2197,N_18995,N_19839);
xnor UO_2198 (O_2198,N_19497,N_18431);
xnor UO_2199 (O_2199,N_19863,N_19585);
and UO_2200 (O_2200,N_18160,N_19220);
nor UO_2201 (O_2201,N_18220,N_18702);
xor UO_2202 (O_2202,N_19803,N_19811);
or UO_2203 (O_2203,N_18458,N_19867);
and UO_2204 (O_2204,N_19501,N_19244);
xor UO_2205 (O_2205,N_18182,N_18332);
and UO_2206 (O_2206,N_19230,N_19056);
nand UO_2207 (O_2207,N_18586,N_19950);
nand UO_2208 (O_2208,N_19326,N_18421);
and UO_2209 (O_2209,N_18871,N_18076);
and UO_2210 (O_2210,N_19701,N_19935);
nand UO_2211 (O_2211,N_19949,N_18251);
nor UO_2212 (O_2212,N_19556,N_19892);
or UO_2213 (O_2213,N_19733,N_19371);
nand UO_2214 (O_2214,N_18643,N_18144);
and UO_2215 (O_2215,N_18506,N_18341);
and UO_2216 (O_2216,N_19713,N_19159);
nand UO_2217 (O_2217,N_19823,N_18602);
nor UO_2218 (O_2218,N_18482,N_19236);
or UO_2219 (O_2219,N_19232,N_18772);
nand UO_2220 (O_2220,N_18171,N_18865);
nand UO_2221 (O_2221,N_19091,N_19919);
nand UO_2222 (O_2222,N_19389,N_19260);
nor UO_2223 (O_2223,N_18261,N_19636);
or UO_2224 (O_2224,N_18707,N_19231);
and UO_2225 (O_2225,N_18923,N_18076);
or UO_2226 (O_2226,N_19570,N_19968);
nand UO_2227 (O_2227,N_19724,N_19120);
nand UO_2228 (O_2228,N_18899,N_19839);
nor UO_2229 (O_2229,N_19875,N_18386);
and UO_2230 (O_2230,N_18361,N_18287);
xor UO_2231 (O_2231,N_18019,N_18313);
nand UO_2232 (O_2232,N_19220,N_19885);
xor UO_2233 (O_2233,N_19245,N_19412);
xnor UO_2234 (O_2234,N_19139,N_18413);
nand UO_2235 (O_2235,N_19492,N_18781);
xnor UO_2236 (O_2236,N_18816,N_18720);
or UO_2237 (O_2237,N_18869,N_18852);
and UO_2238 (O_2238,N_18767,N_18661);
nor UO_2239 (O_2239,N_18716,N_19539);
xnor UO_2240 (O_2240,N_18798,N_19731);
xnor UO_2241 (O_2241,N_18836,N_18034);
or UO_2242 (O_2242,N_18576,N_19427);
nand UO_2243 (O_2243,N_19462,N_19749);
nor UO_2244 (O_2244,N_18201,N_19937);
nor UO_2245 (O_2245,N_19126,N_18352);
and UO_2246 (O_2246,N_18238,N_18286);
or UO_2247 (O_2247,N_19024,N_19685);
xnor UO_2248 (O_2248,N_19429,N_19534);
xnor UO_2249 (O_2249,N_18065,N_19906);
xnor UO_2250 (O_2250,N_18902,N_19908);
nor UO_2251 (O_2251,N_18401,N_19556);
xnor UO_2252 (O_2252,N_18083,N_18884);
xnor UO_2253 (O_2253,N_19468,N_18339);
nor UO_2254 (O_2254,N_18651,N_19505);
nor UO_2255 (O_2255,N_19383,N_19779);
nor UO_2256 (O_2256,N_19268,N_19225);
nand UO_2257 (O_2257,N_18818,N_19441);
and UO_2258 (O_2258,N_19568,N_19776);
xor UO_2259 (O_2259,N_18843,N_18964);
xor UO_2260 (O_2260,N_19495,N_18700);
nand UO_2261 (O_2261,N_19024,N_19990);
nand UO_2262 (O_2262,N_18424,N_19610);
xor UO_2263 (O_2263,N_18650,N_18566);
nand UO_2264 (O_2264,N_18523,N_18522);
or UO_2265 (O_2265,N_18898,N_18192);
or UO_2266 (O_2266,N_18664,N_18135);
and UO_2267 (O_2267,N_18033,N_19634);
and UO_2268 (O_2268,N_18992,N_18104);
xor UO_2269 (O_2269,N_19018,N_18928);
or UO_2270 (O_2270,N_18621,N_18231);
or UO_2271 (O_2271,N_18952,N_18072);
and UO_2272 (O_2272,N_19731,N_19960);
or UO_2273 (O_2273,N_18173,N_18596);
nor UO_2274 (O_2274,N_19937,N_19986);
or UO_2275 (O_2275,N_18308,N_19303);
nand UO_2276 (O_2276,N_19482,N_18647);
or UO_2277 (O_2277,N_18751,N_18081);
xor UO_2278 (O_2278,N_18566,N_19078);
nor UO_2279 (O_2279,N_19404,N_18972);
or UO_2280 (O_2280,N_19994,N_18797);
nor UO_2281 (O_2281,N_19244,N_18110);
nor UO_2282 (O_2282,N_18835,N_18771);
nor UO_2283 (O_2283,N_19296,N_19759);
nand UO_2284 (O_2284,N_19507,N_19691);
nor UO_2285 (O_2285,N_19438,N_19668);
nor UO_2286 (O_2286,N_18094,N_18416);
and UO_2287 (O_2287,N_18862,N_18080);
nor UO_2288 (O_2288,N_18094,N_18156);
nor UO_2289 (O_2289,N_19681,N_18659);
or UO_2290 (O_2290,N_19914,N_18769);
or UO_2291 (O_2291,N_18357,N_19645);
xor UO_2292 (O_2292,N_18382,N_19476);
nor UO_2293 (O_2293,N_18564,N_19988);
and UO_2294 (O_2294,N_18079,N_19988);
or UO_2295 (O_2295,N_19383,N_19767);
xnor UO_2296 (O_2296,N_19389,N_18141);
nor UO_2297 (O_2297,N_18262,N_18828);
xor UO_2298 (O_2298,N_19909,N_19391);
xor UO_2299 (O_2299,N_18665,N_19636);
nand UO_2300 (O_2300,N_19033,N_19456);
xnor UO_2301 (O_2301,N_18483,N_18428);
and UO_2302 (O_2302,N_19548,N_18536);
nor UO_2303 (O_2303,N_18709,N_19437);
and UO_2304 (O_2304,N_18263,N_18821);
xnor UO_2305 (O_2305,N_18328,N_18963);
nand UO_2306 (O_2306,N_18086,N_19181);
nand UO_2307 (O_2307,N_19111,N_18868);
and UO_2308 (O_2308,N_19286,N_19257);
nand UO_2309 (O_2309,N_18646,N_19992);
or UO_2310 (O_2310,N_18778,N_18648);
xnor UO_2311 (O_2311,N_18169,N_18613);
nand UO_2312 (O_2312,N_18996,N_19584);
xnor UO_2313 (O_2313,N_19599,N_19735);
nor UO_2314 (O_2314,N_18272,N_18662);
nor UO_2315 (O_2315,N_19621,N_19110);
nor UO_2316 (O_2316,N_18487,N_19192);
nor UO_2317 (O_2317,N_19421,N_18590);
xnor UO_2318 (O_2318,N_18468,N_18666);
nand UO_2319 (O_2319,N_18095,N_18958);
or UO_2320 (O_2320,N_19911,N_19437);
and UO_2321 (O_2321,N_18110,N_18788);
nand UO_2322 (O_2322,N_19702,N_19193);
nor UO_2323 (O_2323,N_19030,N_18788);
nand UO_2324 (O_2324,N_18406,N_18655);
nand UO_2325 (O_2325,N_18512,N_19262);
xor UO_2326 (O_2326,N_18831,N_19849);
and UO_2327 (O_2327,N_18162,N_19457);
and UO_2328 (O_2328,N_18913,N_18983);
or UO_2329 (O_2329,N_18233,N_19243);
or UO_2330 (O_2330,N_19136,N_19170);
or UO_2331 (O_2331,N_19243,N_18978);
or UO_2332 (O_2332,N_18681,N_19008);
or UO_2333 (O_2333,N_19425,N_19050);
or UO_2334 (O_2334,N_19196,N_18368);
xor UO_2335 (O_2335,N_18165,N_19324);
xnor UO_2336 (O_2336,N_19636,N_19734);
nand UO_2337 (O_2337,N_18678,N_19382);
or UO_2338 (O_2338,N_19478,N_18114);
nand UO_2339 (O_2339,N_18106,N_19432);
nand UO_2340 (O_2340,N_18205,N_19844);
or UO_2341 (O_2341,N_19472,N_19117);
or UO_2342 (O_2342,N_18247,N_19843);
nand UO_2343 (O_2343,N_18739,N_19714);
and UO_2344 (O_2344,N_18577,N_18032);
nand UO_2345 (O_2345,N_18999,N_19407);
or UO_2346 (O_2346,N_19097,N_19061);
nor UO_2347 (O_2347,N_19929,N_19375);
xor UO_2348 (O_2348,N_18055,N_18865);
or UO_2349 (O_2349,N_18262,N_19643);
xnor UO_2350 (O_2350,N_18175,N_18846);
xnor UO_2351 (O_2351,N_19065,N_19993);
and UO_2352 (O_2352,N_18459,N_18769);
or UO_2353 (O_2353,N_19469,N_19041);
or UO_2354 (O_2354,N_19877,N_18320);
nor UO_2355 (O_2355,N_18678,N_19344);
or UO_2356 (O_2356,N_18528,N_18823);
and UO_2357 (O_2357,N_19242,N_18775);
and UO_2358 (O_2358,N_18440,N_19519);
nand UO_2359 (O_2359,N_18231,N_18348);
nand UO_2360 (O_2360,N_18411,N_18419);
nand UO_2361 (O_2361,N_18868,N_19360);
nor UO_2362 (O_2362,N_19482,N_18726);
and UO_2363 (O_2363,N_18173,N_19880);
and UO_2364 (O_2364,N_18978,N_18792);
and UO_2365 (O_2365,N_19378,N_19903);
nand UO_2366 (O_2366,N_19679,N_19272);
or UO_2367 (O_2367,N_19571,N_18582);
or UO_2368 (O_2368,N_19079,N_19151);
nand UO_2369 (O_2369,N_19895,N_18176);
or UO_2370 (O_2370,N_19796,N_19553);
nor UO_2371 (O_2371,N_18668,N_19050);
xor UO_2372 (O_2372,N_19107,N_19784);
and UO_2373 (O_2373,N_18876,N_18760);
nand UO_2374 (O_2374,N_19734,N_19309);
nor UO_2375 (O_2375,N_19004,N_19245);
or UO_2376 (O_2376,N_18606,N_18527);
and UO_2377 (O_2377,N_18775,N_18440);
or UO_2378 (O_2378,N_18473,N_18958);
and UO_2379 (O_2379,N_19982,N_18727);
nand UO_2380 (O_2380,N_19633,N_19107);
nor UO_2381 (O_2381,N_19938,N_19381);
and UO_2382 (O_2382,N_19506,N_18900);
and UO_2383 (O_2383,N_19967,N_18241);
nand UO_2384 (O_2384,N_18627,N_19844);
xnor UO_2385 (O_2385,N_19557,N_19960);
or UO_2386 (O_2386,N_19680,N_18257);
nand UO_2387 (O_2387,N_19543,N_19206);
nand UO_2388 (O_2388,N_19638,N_18592);
or UO_2389 (O_2389,N_19445,N_18962);
and UO_2390 (O_2390,N_18172,N_18625);
nor UO_2391 (O_2391,N_18551,N_19116);
xor UO_2392 (O_2392,N_19377,N_18746);
and UO_2393 (O_2393,N_19336,N_18325);
nor UO_2394 (O_2394,N_19808,N_19906);
nor UO_2395 (O_2395,N_19075,N_19658);
and UO_2396 (O_2396,N_19394,N_18089);
or UO_2397 (O_2397,N_19932,N_18500);
or UO_2398 (O_2398,N_18187,N_18117);
or UO_2399 (O_2399,N_19400,N_18983);
or UO_2400 (O_2400,N_19031,N_18114);
xnor UO_2401 (O_2401,N_18451,N_18770);
or UO_2402 (O_2402,N_18120,N_18394);
xor UO_2403 (O_2403,N_19413,N_18999);
nor UO_2404 (O_2404,N_18410,N_18514);
xnor UO_2405 (O_2405,N_19178,N_18220);
or UO_2406 (O_2406,N_18395,N_19583);
xor UO_2407 (O_2407,N_18263,N_18855);
nor UO_2408 (O_2408,N_19145,N_19947);
nand UO_2409 (O_2409,N_19470,N_19512);
nor UO_2410 (O_2410,N_19347,N_19752);
and UO_2411 (O_2411,N_19903,N_18876);
xnor UO_2412 (O_2412,N_19075,N_18133);
xnor UO_2413 (O_2413,N_19868,N_18445);
and UO_2414 (O_2414,N_19359,N_18278);
nor UO_2415 (O_2415,N_18485,N_18649);
or UO_2416 (O_2416,N_18204,N_19036);
nor UO_2417 (O_2417,N_18712,N_18418);
or UO_2418 (O_2418,N_18380,N_19240);
xor UO_2419 (O_2419,N_19332,N_19391);
and UO_2420 (O_2420,N_18710,N_18907);
and UO_2421 (O_2421,N_19607,N_18855);
or UO_2422 (O_2422,N_19593,N_19705);
nor UO_2423 (O_2423,N_18623,N_18730);
nand UO_2424 (O_2424,N_18678,N_18349);
xnor UO_2425 (O_2425,N_18497,N_18638);
or UO_2426 (O_2426,N_18013,N_18737);
nor UO_2427 (O_2427,N_19390,N_19377);
nand UO_2428 (O_2428,N_18939,N_18432);
and UO_2429 (O_2429,N_18774,N_18373);
and UO_2430 (O_2430,N_18364,N_19403);
nand UO_2431 (O_2431,N_18130,N_19736);
nor UO_2432 (O_2432,N_18641,N_19718);
nand UO_2433 (O_2433,N_19510,N_19048);
nor UO_2434 (O_2434,N_18351,N_18467);
and UO_2435 (O_2435,N_19612,N_19336);
xor UO_2436 (O_2436,N_18909,N_19919);
nand UO_2437 (O_2437,N_18117,N_18453);
or UO_2438 (O_2438,N_18500,N_18451);
nor UO_2439 (O_2439,N_19516,N_18534);
and UO_2440 (O_2440,N_18988,N_18650);
nand UO_2441 (O_2441,N_19692,N_18361);
nand UO_2442 (O_2442,N_18921,N_19063);
and UO_2443 (O_2443,N_18866,N_18676);
or UO_2444 (O_2444,N_18187,N_19891);
and UO_2445 (O_2445,N_19441,N_18010);
and UO_2446 (O_2446,N_18132,N_19683);
nand UO_2447 (O_2447,N_19420,N_19082);
xor UO_2448 (O_2448,N_19345,N_18934);
nor UO_2449 (O_2449,N_18729,N_19631);
nand UO_2450 (O_2450,N_18594,N_18954);
nor UO_2451 (O_2451,N_18536,N_18163);
xor UO_2452 (O_2452,N_18544,N_18236);
xnor UO_2453 (O_2453,N_18463,N_19291);
and UO_2454 (O_2454,N_18222,N_18999);
nand UO_2455 (O_2455,N_18073,N_18924);
nor UO_2456 (O_2456,N_18408,N_19406);
nand UO_2457 (O_2457,N_18862,N_19750);
nor UO_2458 (O_2458,N_19544,N_18359);
xor UO_2459 (O_2459,N_18290,N_18148);
nand UO_2460 (O_2460,N_19530,N_18053);
nand UO_2461 (O_2461,N_18009,N_19725);
or UO_2462 (O_2462,N_18409,N_19776);
xnor UO_2463 (O_2463,N_19719,N_18716);
nor UO_2464 (O_2464,N_18147,N_18097);
nand UO_2465 (O_2465,N_19078,N_19039);
and UO_2466 (O_2466,N_18046,N_18466);
or UO_2467 (O_2467,N_18464,N_19437);
xor UO_2468 (O_2468,N_18310,N_18268);
and UO_2469 (O_2469,N_18167,N_19965);
nor UO_2470 (O_2470,N_18985,N_19906);
or UO_2471 (O_2471,N_19601,N_19701);
and UO_2472 (O_2472,N_18365,N_19951);
xnor UO_2473 (O_2473,N_19865,N_18083);
nor UO_2474 (O_2474,N_19538,N_19611);
or UO_2475 (O_2475,N_19955,N_19672);
and UO_2476 (O_2476,N_18507,N_19874);
nor UO_2477 (O_2477,N_18923,N_19991);
and UO_2478 (O_2478,N_18371,N_18564);
and UO_2479 (O_2479,N_19361,N_19440);
xnor UO_2480 (O_2480,N_18439,N_19420);
and UO_2481 (O_2481,N_19824,N_19602);
nand UO_2482 (O_2482,N_18760,N_19749);
xor UO_2483 (O_2483,N_19301,N_18592);
or UO_2484 (O_2484,N_18923,N_18458);
nor UO_2485 (O_2485,N_19320,N_18723);
or UO_2486 (O_2486,N_19278,N_18270);
and UO_2487 (O_2487,N_18894,N_19932);
and UO_2488 (O_2488,N_19293,N_19779);
xor UO_2489 (O_2489,N_18455,N_18667);
nand UO_2490 (O_2490,N_18471,N_19872);
xor UO_2491 (O_2491,N_18127,N_18281);
nand UO_2492 (O_2492,N_18730,N_19293);
and UO_2493 (O_2493,N_19061,N_18653);
nor UO_2494 (O_2494,N_19033,N_18225);
xor UO_2495 (O_2495,N_19994,N_18269);
nor UO_2496 (O_2496,N_19842,N_19834);
and UO_2497 (O_2497,N_19468,N_18012);
nand UO_2498 (O_2498,N_18381,N_19268);
nand UO_2499 (O_2499,N_18619,N_18559);
endmodule