module basic_3000_30000_3500_30_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xnor U0 (N_0,In_2720,In_2879);
xnor U1 (N_1,In_2774,In_1597);
nor U2 (N_2,In_2678,In_1401);
nor U3 (N_3,In_21,In_1820);
or U4 (N_4,In_1625,In_668);
nor U5 (N_5,In_1069,In_1480);
or U6 (N_6,In_1816,In_1445);
nand U7 (N_7,In_2583,In_906);
and U8 (N_8,In_1240,In_1925);
or U9 (N_9,In_2865,In_1224);
and U10 (N_10,In_956,In_128);
nor U11 (N_11,In_1471,In_1253);
nand U12 (N_12,In_2902,In_1587);
xnor U13 (N_13,In_309,In_508);
nor U14 (N_14,In_2735,In_1773);
nand U15 (N_15,In_151,In_2743);
nor U16 (N_16,In_45,In_327);
nand U17 (N_17,In_2688,In_85);
nand U18 (N_18,In_1135,In_422);
and U19 (N_19,In_2385,In_758);
or U20 (N_20,In_2518,In_1398);
nand U21 (N_21,In_199,In_1723);
nand U22 (N_22,In_1121,In_2940);
or U23 (N_23,In_2207,In_1032);
or U24 (N_24,In_1279,In_2021);
nor U25 (N_25,In_655,In_1477);
and U26 (N_26,In_790,In_548);
or U27 (N_27,In_22,In_576);
nand U28 (N_28,In_2777,In_1428);
or U29 (N_29,In_2004,In_2556);
nand U30 (N_30,In_1713,In_2151);
nor U31 (N_31,In_2223,In_1647);
nand U32 (N_32,In_1159,In_2499);
xnor U33 (N_33,In_100,In_775);
nor U34 (N_34,In_2833,In_2367);
or U35 (N_35,In_1975,In_1999);
nand U36 (N_36,In_2477,In_250);
xnor U37 (N_37,In_2226,In_2256);
nand U38 (N_38,In_397,In_392);
and U39 (N_39,In_1856,In_101);
nand U40 (N_40,In_1803,In_1619);
nand U41 (N_41,In_705,In_163);
or U42 (N_42,In_2449,In_2211);
xor U43 (N_43,In_1793,In_1276);
or U44 (N_44,In_2103,In_2338);
nor U45 (N_45,In_2962,In_1048);
and U46 (N_46,In_657,In_2277);
nor U47 (N_47,In_2278,In_653);
nor U48 (N_48,In_504,In_835);
nor U49 (N_49,In_1940,In_446);
or U50 (N_50,In_1890,In_2347);
and U51 (N_51,In_2623,In_2576);
nand U52 (N_52,In_1570,In_2780);
xnor U53 (N_53,In_2936,In_982);
xor U54 (N_54,In_2569,In_649);
nor U55 (N_55,In_1060,In_278);
or U56 (N_56,In_67,In_1823);
and U57 (N_57,In_2817,In_2716);
xor U58 (N_58,In_2221,In_2630);
or U59 (N_59,In_164,In_2174);
nand U60 (N_60,In_641,In_453);
nand U61 (N_61,In_1854,In_300);
and U62 (N_62,In_2984,In_2);
and U63 (N_63,In_511,In_1110);
nor U64 (N_64,In_2648,In_1039);
and U65 (N_65,In_2590,In_1315);
and U66 (N_66,In_1661,In_771);
or U67 (N_67,In_2549,In_2788);
and U68 (N_68,In_2572,In_419);
or U69 (N_69,In_2608,In_2228);
and U70 (N_70,In_1553,In_1677);
nor U71 (N_71,In_1111,In_2983);
or U72 (N_72,In_1754,In_1789);
nor U73 (N_73,In_1105,In_2649);
nand U74 (N_74,In_166,In_2547);
nand U75 (N_75,In_1298,In_2712);
or U76 (N_76,In_2677,In_1444);
nand U77 (N_77,In_939,In_2670);
or U78 (N_78,In_1629,In_320);
nand U79 (N_79,In_2265,In_934);
xnor U80 (N_80,In_2076,In_132);
nor U81 (N_81,In_2302,In_630);
nor U82 (N_82,In_1431,In_1651);
and U83 (N_83,In_1148,In_2708);
nor U84 (N_84,In_1044,In_1182);
or U85 (N_85,In_2316,In_957);
nand U86 (N_86,In_1139,In_1404);
and U87 (N_87,In_615,In_2158);
or U88 (N_88,In_492,In_2083);
nor U89 (N_89,In_2908,In_274);
xor U90 (N_90,In_2880,In_1372);
nand U91 (N_91,In_1842,In_2717);
or U92 (N_92,In_1680,In_2749);
xnor U93 (N_93,In_2822,In_2399);
and U94 (N_94,In_2327,In_1607);
and U95 (N_95,In_1905,In_2467);
or U96 (N_96,In_2516,In_1157);
xnor U97 (N_97,In_496,In_334);
nand U98 (N_98,In_1106,In_776);
and U99 (N_99,In_747,In_1806);
xnor U100 (N_100,In_2182,In_1951);
and U101 (N_101,In_525,In_581);
and U102 (N_102,In_2172,In_811);
xnor U103 (N_103,In_1528,In_1154);
xnor U104 (N_104,In_1388,In_2424);
or U105 (N_105,In_283,In_733);
and U106 (N_106,In_2905,In_2136);
xor U107 (N_107,In_1019,In_2317);
nor U108 (N_108,In_1799,In_524);
xor U109 (N_109,In_933,In_2289);
nand U110 (N_110,In_1129,In_1420);
and U111 (N_111,In_204,In_2740);
and U112 (N_112,In_1235,In_987);
and U113 (N_113,In_1515,In_56);
and U114 (N_114,In_537,In_610);
or U115 (N_115,In_1558,In_2819);
nand U116 (N_116,In_779,In_2168);
and U117 (N_117,In_1338,In_769);
xor U118 (N_118,In_2884,In_1817);
and U119 (N_119,In_1426,In_777);
xor U120 (N_120,In_1700,In_382);
or U121 (N_121,In_952,In_2640);
and U122 (N_122,In_2563,In_1517);
xor U123 (N_123,In_42,In_2292);
nor U124 (N_124,In_901,In_1221);
nand U125 (N_125,In_2016,In_2000);
xnor U126 (N_126,In_1473,In_1920);
nand U127 (N_127,In_2821,In_116);
nor U128 (N_128,In_1813,In_583);
or U129 (N_129,In_2929,In_1170);
xnor U130 (N_130,In_1311,In_1965);
or U131 (N_131,In_839,In_2089);
nor U132 (N_132,In_1772,In_1829);
nor U133 (N_133,In_1871,In_214);
nor U134 (N_134,In_1861,In_2836);
or U135 (N_135,In_348,In_2489);
xor U136 (N_136,In_2233,In_2726);
nor U137 (N_137,In_2546,In_12);
and U138 (N_138,In_1695,In_596);
xnor U139 (N_139,In_1676,In_1821);
xnor U140 (N_140,In_595,In_1917);
xor U141 (N_141,In_1491,In_891);
and U142 (N_142,In_1826,In_1881);
or U143 (N_143,In_2269,In_1012);
or U144 (N_144,In_2533,In_2795);
or U145 (N_145,In_903,In_2188);
or U146 (N_146,In_39,In_817);
or U147 (N_147,In_49,In_1664);
nand U148 (N_148,In_1561,In_2508);
or U149 (N_149,In_2617,In_1163);
and U150 (N_150,In_2112,In_2970);
nand U151 (N_151,In_2117,In_171);
nand U152 (N_152,In_1008,In_828);
nor U153 (N_153,In_236,In_735);
nand U154 (N_154,In_2279,In_804);
nor U155 (N_155,In_408,In_846);
and U156 (N_156,In_2017,In_2229);
nor U157 (N_157,In_1175,In_1027);
nand U158 (N_158,In_119,In_2619);
xnor U159 (N_159,In_764,In_1482);
or U160 (N_160,In_1234,In_1396);
nor U161 (N_161,In_470,In_883);
nor U162 (N_162,In_456,In_824);
xor U163 (N_163,In_2032,In_1208);
xor U164 (N_164,In_1874,In_1758);
or U165 (N_165,In_99,In_2213);
xnor U166 (N_166,In_2283,In_2039);
or U167 (N_167,In_326,In_2133);
nor U168 (N_168,In_1931,In_1631);
xor U169 (N_169,In_1215,In_1063);
nor U170 (N_170,In_1853,In_393);
nor U171 (N_171,In_2540,In_2679);
and U172 (N_172,In_2268,In_213);
xnor U173 (N_173,In_2320,In_2014);
and U174 (N_174,In_245,In_2602);
nor U175 (N_175,In_1565,In_910);
and U176 (N_176,In_2309,In_748);
or U177 (N_177,In_2513,In_1801);
and U178 (N_178,In_2830,In_1857);
or U179 (N_179,In_399,In_1082);
nor U180 (N_180,In_2995,In_1675);
nand U181 (N_181,In_688,In_1369);
and U182 (N_182,In_1072,In_1912);
nor U183 (N_183,In_1589,In_2628);
or U184 (N_184,In_2621,In_1132);
nor U185 (N_185,In_922,In_1074);
nand U186 (N_186,In_1366,In_2593);
nand U187 (N_187,In_279,In_1996);
xnor U188 (N_188,In_2090,In_979);
or U189 (N_189,In_9,In_1930);
xnor U190 (N_190,In_2991,In_2994);
nor U191 (N_191,In_2762,In_2371);
or U192 (N_192,In_1704,In_2646);
and U193 (N_193,In_1374,In_1417);
nor U194 (N_194,In_2642,In_1083);
xor U195 (N_195,In_1638,In_2956);
or U196 (N_196,In_1418,In_1569);
nand U197 (N_197,In_1606,In_2791);
and U198 (N_198,In_795,In_385);
or U199 (N_199,In_2531,In_520);
nor U200 (N_200,In_2056,In_505);
and U201 (N_201,In_2336,In_4);
and U202 (N_202,In_2482,In_485);
or U203 (N_203,In_1540,In_555);
xor U204 (N_204,In_486,In_2715);
nor U205 (N_205,In_2887,In_458);
and U206 (N_206,In_2051,In_369);
nor U207 (N_207,In_2658,In_292);
and U208 (N_208,In_1024,In_338);
xnor U209 (N_209,In_2775,In_570);
nand U210 (N_210,In_1467,In_1299);
xor U211 (N_211,In_1893,In_1249);
nor U212 (N_212,In_2093,In_2118);
nand U213 (N_213,In_566,In_1909);
nand U214 (N_214,In_2250,In_1499);
or U215 (N_215,In_1204,In_700);
or U216 (N_216,In_2573,In_2859);
or U217 (N_217,In_1641,In_2344);
and U218 (N_218,In_175,In_2684);
and U219 (N_219,In_1453,In_315);
and U220 (N_220,In_416,In_988);
nor U221 (N_221,In_1440,In_2178);
or U222 (N_222,In_1013,In_980);
and U223 (N_223,In_440,In_442);
and U224 (N_224,In_156,In_2258);
xnor U225 (N_225,In_2035,In_1167);
nor U226 (N_226,In_746,In_1708);
or U227 (N_227,In_322,In_2522);
or U228 (N_228,In_83,In_1058);
xnor U229 (N_229,In_2007,In_1261);
nand U230 (N_230,In_469,In_1584);
nor U231 (N_231,In_2696,In_1284);
nand U232 (N_232,In_1971,In_117);
nand U233 (N_233,In_905,In_1673);
or U234 (N_234,In_693,In_2730);
nor U235 (N_235,In_2537,In_1860);
xor U236 (N_236,In_1352,In_154);
and U237 (N_237,In_765,In_1452);
or U238 (N_238,In_2129,In_1578);
xnor U239 (N_239,In_1686,In_1034);
and U240 (N_240,In_951,In_639);
xor U241 (N_241,In_1066,In_174);
or U242 (N_242,In_1679,In_2374);
nor U243 (N_243,In_2186,In_1603);
nand U244 (N_244,In_142,In_2615);
or U245 (N_245,In_2350,In_1510);
and U246 (N_246,In_281,In_1811);
nand U247 (N_247,In_493,In_1674);
nand U248 (N_248,In_2806,In_2885);
or U249 (N_249,In_227,In_2781);
nor U250 (N_250,In_2393,In_604);
or U251 (N_251,In_620,In_450);
and U252 (N_252,In_256,In_311);
nand U253 (N_253,In_1877,In_1290);
xor U254 (N_254,In_698,In_473);
nor U255 (N_255,In_2511,In_1796);
or U256 (N_256,In_2818,In_1539);
nand U257 (N_257,In_345,In_2377);
nor U258 (N_258,In_2725,In_478);
nand U259 (N_259,In_517,In_2542);
xnor U260 (N_260,In_896,In_1825);
nand U261 (N_261,In_884,In_1898);
xnor U262 (N_262,In_1283,In_2834);
nor U263 (N_263,In_31,In_378);
and U264 (N_264,In_1405,In_2661);
nor U265 (N_265,In_146,In_2579);
nand U266 (N_266,In_2381,In_1333);
xor U267 (N_267,In_2194,In_2690);
and U268 (N_268,In_1255,In_471);
xor U269 (N_269,In_2974,In_2175);
nand U270 (N_270,In_2939,In_1943);
nor U271 (N_271,In_1351,In_659);
nand U272 (N_272,In_360,In_179);
or U273 (N_273,In_387,In_529);
nand U274 (N_274,In_2029,In_1936);
xor U275 (N_275,In_2699,In_1688);
or U276 (N_276,In_2237,In_1757);
xor U277 (N_277,In_2030,In_1133);
and U278 (N_278,In_1002,In_2967);
and U279 (N_279,In_660,In_2564);
and U280 (N_280,In_945,In_876);
xor U281 (N_281,In_1814,In_1748);
nand U282 (N_282,In_2999,In_983);
xnor U283 (N_283,In_1775,In_193);
and U284 (N_284,In_304,In_401);
or U285 (N_285,In_102,In_2724);
and U286 (N_286,In_2741,In_2733);
xor U287 (N_287,In_2812,In_1150);
or U288 (N_288,In_2494,In_1070);
nand U289 (N_289,In_2747,In_1838);
nor U290 (N_290,In_2084,In_1870);
nor U291 (N_291,In_1531,In_1228);
xnor U292 (N_292,In_2744,In_1541);
nor U293 (N_293,In_2758,In_538);
nor U294 (N_294,In_2916,In_96);
nand U295 (N_295,In_133,In_1736);
xnor U296 (N_296,In_940,In_1800);
and U297 (N_297,In_1161,In_807);
nand U298 (N_298,In_995,In_1939);
nand U299 (N_299,In_1545,In_1859);
nor U300 (N_300,In_72,In_1468);
nor U301 (N_301,In_1265,In_1892);
xnor U302 (N_302,In_1644,In_192);
or U303 (N_303,In_1325,In_1997);
xnor U304 (N_304,In_1572,In_230);
and U305 (N_305,In_452,In_895);
nand U306 (N_306,In_2404,In_833);
xor U307 (N_307,In_2378,In_1178);
or U308 (N_308,In_302,In_1031);
xor U309 (N_309,In_1025,In_2846);
and U310 (N_310,In_2322,In_2917);
xnor U311 (N_311,In_1119,In_1096);
nor U312 (N_312,In_1463,In_2691);
xor U313 (N_313,In_388,In_1579);
nor U314 (N_314,In_1502,In_977);
nor U315 (N_315,In_1866,In_135);
xor U316 (N_316,In_1145,In_1582);
xor U317 (N_317,In_861,In_1714);
and U318 (N_318,In_2306,In_1273);
or U319 (N_319,In_637,In_561);
and U320 (N_320,In_1551,In_2180);
nand U321 (N_321,In_865,In_293);
or U322 (N_322,In_1899,In_830);
xnor U323 (N_323,In_2011,In_165);
nor U324 (N_324,In_1537,In_1383);
or U325 (N_325,In_715,In_2711);
xnor U326 (N_326,In_209,In_2308);
nand U327 (N_327,In_986,In_2847);
and U328 (N_328,In_1164,In_2526);
and U329 (N_329,In_2413,In_2061);
nand U330 (N_330,In_2465,In_887);
xor U331 (N_331,In_2584,In_1250);
and U332 (N_332,In_2675,In_722);
and U333 (N_333,In_2636,In_1845);
nand U334 (N_334,In_202,In_1506);
and U335 (N_335,In_51,In_1962);
xor U336 (N_336,In_244,In_1252);
and U337 (N_337,In_1655,In_201);
and U338 (N_338,In_1743,In_2271);
or U339 (N_339,In_2510,In_1851);
and U340 (N_340,In_1568,In_2550);
and U341 (N_341,In_1323,In_946);
and U342 (N_342,In_2270,In_1321);
nor U343 (N_343,In_2527,In_2881);
and U344 (N_344,In_2848,In_2509);
xnor U345 (N_345,In_1872,In_349);
and U346 (N_346,In_1518,In_20);
and U347 (N_347,In_1294,In_1219);
nand U348 (N_348,In_624,In_2938);
nand U349 (N_349,In_1200,In_183);
nor U350 (N_350,In_1436,In_2096);
xor U351 (N_351,In_2582,In_2605);
nor U352 (N_352,In_61,In_1470);
and U353 (N_353,In_1529,In_2387);
or U354 (N_354,In_1465,In_554);
nor U355 (N_355,In_2689,In_459);
xnor U356 (N_356,In_2548,In_2931);
or U357 (N_357,In_1009,In_2596);
or U358 (N_358,In_2832,In_673);
nor U359 (N_359,In_1264,In_918);
and U360 (N_360,In_1068,In_2495);
and U361 (N_361,In_358,In_2372);
nand U362 (N_362,In_73,In_2941);
xnor U363 (N_363,In_2086,In_2355);
nor U364 (N_364,In_2107,In_2475);
nor U365 (N_365,In_2654,In_2875);
nor U366 (N_366,In_1292,In_70);
nor U367 (N_367,In_1310,In_275);
or U368 (N_368,In_2959,In_2366);
nand U369 (N_369,In_516,In_1441);
or U370 (N_370,In_1165,In_1071);
or U371 (N_371,In_2454,In_1991);
nor U372 (N_372,In_229,In_1409);
xnor U373 (N_373,In_2328,In_1730);
or U374 (N_374,In_1256,In_778);
nor U375 (N_375,In_707,In_531);
xnor U376 (N_376,In_1370,In_1867);
and U377 (N_377,In_1018,In_1633);
xor U378 (N_378,In_1717,In_2814);
xnor U379 (N_379,In_1573,In_435);
or U380 (N_380,In_2438,In_2502);
xnor U381 (N_381,In_1160,In_1636);
and U382 (N_382,In_1144,In_1056);
and U383 (N_383,In_1014,In_860);
xor U384 (N_384,In_1424,In_1771);
nand U385 (N_385,In_1972,In_1776);
nand U386 (N_386,In_938,In_2215);
or U387 (N_387,In_1974,In_853);
nor U388 (N_388,In_28,In_2653);
and U389 (N_389,In_1976,In_181);
xor U390 (N_390,In_683,In_2342);
xor U391 (N_391,In_2199,In_75);
or U392 (N_392,In_370,In_2315);
nand U393 (N_393,In_186,In_476);
or U394 (N_394,In_2957,In_2784);
nand U395 (N_395,In_2468,In_1314);
nor U396 (N_396,In_1319,In_2723);
or U397 (N_397,In_943,In_10);
xnor U398 (N_398,In_605,In_2388);
or U399 (N_399,In_2041,In_1488);
nor U400 (N_400,In_336,In_2667);
xor U401 (N_401,In_1266,In_766);
and U402 (N_402,In_791,In_1672);
and U403 (N_403,In_1852,In_2910);
nand U404 (N_404,In_120,In_2249);
and U405 (N_405,In_1855,In_1028);
nor U406 (N_406,In_305,In_2329);
and U407 (N_407,In_1001,In_2487);
nor U408 (N_408,In_1836,In_2068);
nand U409 (N_409,In_1320,In_2113);
xnor U410 (N_410,In_1822,In_2709);
nor U411 (N_411,In_1828,In_2925);
or U412 (N_412,In_1837,In_1623);
xor U413 (N_413,In_27,In_2165);
nor U414 (N_414,In_2290,In_850);
and U415 (N_415,In_2559,In_503);
or U416 (N_416,In_68,In_749);
nor U417 (N_417,In_2052,In_1611);
nand U418 (N_418,In_932,In_645);
or U419 (N_419,In_2230,In_547);
nor U420 (N_420,In_1514,In_1097);
nand U421 (N_421,In_2868,In_961);
or U422 (N_422,In_2447,In_110);
or U423 (N_423,In_955,In_2862);
and U424 (N_424,In_2973,In_793);
and U425 (N_425,In_1654,In_1935);
nand U426 (N_426,In_2247,In_1302);
nand U427 (N_427,In_2166,In_719);
or U428 (N_428,In_420,In_1538);
or U429 (N_429,In_2826,In_1146);
nand U430 (N_430,In_2722,In_2924);
nor U431 (N_431,In_2567,In_118);
and U432 (N_432,In_325,In_1262);
xor U433 (N_433,In_1438,In_168);
nor U434 (N_434,In_984,In_1696);
or U435 (N_435,In_2988,In_2321);
xnor U436 (N_436,In_391,In_1594);
nor U437 (N_437,In_1613,In_2202);
nor U438 (N_438,In_2861,In_1040);
or U439 (N_439,In_2571,In_224);
nor U440 (N_440,In_2702,In_314);
or U441 (N_441,In_2038,In_522);
and U442 (N_442,In_366,In_2672);
nor U443 (N_443,In_80,In_1508);
and U444 (N_444,In_740,In_1968);
nand U445 (N_445,In_1251,In_991);
nand U446 (N_446,In_2053,In_2243);
or U447 (N_447,In_2443,In_1990);
nand U448 (N_448,In_2288,In_541);
xor U449 (N_449,In_2356,In_2624);
xnor U450 (N_450,In_1894,In_1626);
nand U451 (N_451,In_188,In_2431);
and U452 (N_452,In_2142,In_1429);
or U453 (N_453,In_507,In_2330);
nand U454 (N_454,In_2534,In_290);
nor U455 (N_455,In_243,In_1332);
or U456 (N_456,In_1630,In_1022);
xnor U457 (N_457,In_2274,In_1762);
xnor U458 (N_458,In_103,In_1765);
or U459 (N_459,In_2358,In_569);
nor U460 (N_460,In_2219,In_2512);
and U461 (N_461,In_1094,In_1459);
nor U462 (N_462,In_2073,In_838);
and U463 (N_463,In_1658,In_720);
or U464 (N_464,In_2947,In_2200);
and U465 (N_465,In_246,In_2173);
and U466 (N_466,In_1493,In_2234);
and U467 (N_467,In_1478,In_1634);
or U468 (N_468,In_2609,In_2622);
nor U469 (N_469,In_1802,In_2102);
nand U470 (N_470,In_1992,In_1648);
xnor U471 (N_471,In_413,In_1557);
nor U472 (N_472,In_1928,In_947);
nor U473 (N_473,In_871,In_1196);
nand U474 (N_474,In_1339,In_1079);
nor U475 (N_475,In_1687,In_837);
nand U476 (N_476,In_223,In_1891);
and U477 (N_477,In_1199,In_1073);
nand U478 (N_478,In_1516,In_2769);
nor U479 (N_479,In_1412,In_2799);
or U480 (N_480,In_260,In_307);
or U481 (N_481,In_55,In_126);
nor U482 (N_482,In_2162,In_2335);
or U483 (N_483,In_584,In_1458);
xor U484 (N_484,In_129,In_2303);
and U485 (N_485,In_78,In_1632);
and U486 (N_486,In_536,In_1795);
nand U487 (N_487,In_597,In_613);
and U488 (N_488,In_226,In_1141);
and U489 (N_489,In_759,In_2209);
or U490 (N_490,In_1649,In_781);
xor U491 (N_491,In_234,In_1317);
xnor U492 (N_492,In_985,In_1878);
and U493 (N_493,In_593,In_1140);
nand U494 (N_494,In_2115,In_2909);
and U495 (N_495,In_498,In_2024);
xor U496 (N_496,In_929,In_2078);
xor U497 (N_497,In_2240,In_879);
and U498 (N_498,In_2488,In_1722);
nand U499 (N_499,In_754,In_2960);
or U500 (N_500,In_2177,In_2490);
nor U501 (N_501,In_1354,In_94);
and U502 (N_502,In_2034,In_2169);
or U503 (N_503,In_2792,In_974);
nand U504 (N_504,In_1527,In_2864);
or U505 (N_505,In_2284,In_261);
nand U506 (N_506,In_1300,In_914);
or U507 (N_507,In_724,In_629);
and U508 (N_508,In_621,In_1747);
nand U509 (N_509,In_159,In_788);
nand U510 (N_510,In_1371,In_418);
and U511 (N_511,In_559,In_8);
nand U512 (N_512,In_1639,In_2314);
or U513 (N_513,In_2515,In_730);
nand U514 (N_514,In_454,In_2850);
and U515 (N_515,In_232,In_1535);
nor U516 (N_516,In_975,In_2866);
nor U517 (N_517,In_1995,In_1202);
nand U518 (N_518,In_867,In_331);
and U519 (N_519,In_316,In_97);
or U520 (N_520,In_701,In_1421);
or U521 (N_521,In_1733,In_332);
nor U522 (N_522,In_1504,In_1662);
nor U523 (N_523,In_2532,In_869);
or U524 (N_524,In_2707,In_2587);
xnor U525 (N_525,In_303,In_2281);
nand U526 (N_526,In_512,In_2236);
nor U527 (N_527,In_1189,In_1970);
nor U528 (N_528,In_149,In_2578);
nand U529 (N_529,In_1174,In_1850);
xor U530 (N_530,In_821,In_877);
and U531 (N_531,In_2524,In_1343);
and U532 (N_532,In_2616,In_2803);
nand U533 (N_533,In_1117,In_1843);
and U534 (N_534,In_2020,In_2380);
nand U535 (N_535,In_1267,In_87);
nand U536 (N_536,In_2926,In_1918);
and U537 (N_537,In_1604,In_2445);
and U538 (N_538,In_1635,In_1394);
nor U539 (N_539,In_592,In_1941);
and U540 (N_540,In_1443,In_455);
and U541 (N_541,In_1566,In_2625);
or U542 (N_542,In_2131,In_367);
nor U543 (N_543,In_2555,In_251);
and U544 (N_544,In_2354,In_1884);
nor U545 (N_545,In_115,In_2008);
or U546 (N_546,In_1749,In_2565);
xor U547 (N_547,In_1500,In_681);
nor U548 (N_548,In_794,In_286);
xnor U549 (N_549,In_1581,In_2701);
xnor U550 (N_550,In_2643,In_2514);
xor U551 (N_551,In_2987,In_675);
and U552 (N_552,In_2227,In_997);
xor U553 (N_553,In_79,In_130);
nor U554 (N_554,In_2976,In_430);
nand U555 (N_555,In_1684,In_1978);
xnor U556 (N_556,In_2085,In_718);
or U557 (N_557,In_2192,In_534);
and U558 (N_558,In_373,In_184);
and U559 (N_559,In_1798,In_1787);
nor U560 (N_560,In_1065,In_2633);
and U561 (N_561,In_589,In_2224);
and U562 (N_562,In_356,In_2721);
or U563 (N_563,In_1462,In_2300);
or U564 (N_564,In_488,In_1542);
and U565 (N_565,In_1501,In_176);
nand U566 (N_566,In_598,In_1128);
nand U567 (N_567,In_2789,In_958);
xor U568 (N_568,In_1143,In_1481);
and U569 (N_569,In_1184,In_1947);
nand U570 (N_570,In_66,In_90);
nor U571 (N_571,In_2440,In_2553);
or U572 (N_572,In_157,In_448);
xor U573 (N_573,In_990,In_964);
nor U574 (N_574,In_2075,In_1454);
nand U575 (N_575,In_390,In_2964);
xnor U576 (N_576,In_677,In_996);
xnor U577 (N_577,In_1301,In_1967);
or U578 (N_578,In_2614,In_1910);
nor U579 (N_579,In_15,In_1608);
and U580 (N_580,In_1287,In_2139);
and U581 (N_581,In_1247,In_301);
or U582 (N_582,In_1407,In_1191);
and U583 (N_583,In_2889,In_1122);
or U584 (N_584,In_2787,In_1092);
xnor U585 (N_585,In_1327,In_1588);
nor U586 (N_586,In_1331,In_2466);
nand U587 (N_587,In_1791,In_479);
or U588 (N_588,In_622,In_2242);
xor U589 (N_589,In_844,In_206);
nand U590 (N_590,In_734,In_976);
or U591 (N_591,In_2694,In_484);
nor U592 (N_592,In_900,In_2921);
or U593 (N_593,In_405,In_2433);
or U594 (N_594,In_1567,In_2410);
and U595 (N_595,In_2206,In_864);
nor U596 (N_596,In_682,In_2928);
and U597 (N_597,In_616,In_1815);
or U598 (N_598,In_2755,In_1835);
nor U599 (N_599,In_2181,In_1591);
or U600 (N_600,In_1739,In_2164);
and U601 (N_601,In_1702,In_1770);
and U602 (N_602,In_1595,In_2503);
or U603 (N_603,In_1263,In_402);
nand U604 (N_604,In_575,In_2363);
or U605 (N_605,In_2122,In_2225);
or U606 (N_606,In_1393,In_2049);
xor U607 (N_607,In_1245,In_2001);
and U608 (N_608,In_556,In_2856);
or U609 (N_609,In_2459,In_704);
or U610 (N_610,In_1296,In_723);
xor U611 (N_611,In_783,In_2852);
and U612 (N_612,In_2800,In_2023);
nand U613 (N_613,In_1742,In_571);
nand U614 (N_614,In_2379,In_2807);
nor U615 (N_615,In_1562,In_2927);
nor U616 (N_616,In_1667,In_729);
nand U617 (N_617,In_1668,In_2551);
and U618 (N_618,In_2116,In_2692);
or U619 (N_619,In_1994,In_1681);
and U620 (N_620,In_1238,In_1042);
and U621 (N_621,In_123,In_1177);
or U622 (N_622,In_880,In_1084);
nor U623 (N_623,In_672,In_1342);
and U624 (N_624,In_363,In_60);
and U625 (N_625,In_1479,In_515);
and U626 (N_626,In_2886,In_1960);
or U627 (N_627,In_1373,In_1977);
nor U628 (N_628,In_1316,In_196);
nand U629 (N_629,In_810,In_530);
and U630 (N_630,In_1180,In_582);
and U631 (N_631,In_2680,In_2953);
xnor U632 (N_632,In_2906,In_2287);
nor U633 (N_633,In_1896,In_1906);
and U634 (N_634,In_711,In_1669);
and U635 (N_635,In_2801,In_1600);
xor U636 (N_636,In_1764,In_679);
xnor U637 (N_637,In_1780,In_761);
and U638 (N_638,In_1166,In_1218);
xor U639 (N_639,In_50,In_215);
nand U640 (N_640,In_1173,In_2072);
or U641 (N_641,In_2275,In_1364);
and U642 (N_642,In_1334,In_1380);
and U643 (N_643,In_1387,In_407);
nor U644 (N_644,In_365,In_1660);
nor U645 (N_645,In_1403,In_1819);
xor U646 (N_646,In_1483,In_941);
nand U647 (N_647,In_2607,In_403);
or U648 (N_648,In_1929,In_41);
xor U649 (N_649,In_1193,In_1304);
and U650 (N_650,In_2087,In_2837);
and U651 (N_651,In_927,In_2652);
and U652 (N_652,In_550,In_2401);
xnor U653 (N_653,In_2239,In_1737);
and U654 (N_654,In_1761,In_2476);
or U655 (N_655,In_1000,In_443);
nand U656 (N_656,In_1485,In_1385);
xnor U657 (N_657,In_1492,In_1659);
nand U658 (N_658,In_1203,In_2718);
nand U659 (N_659,In_44,In_1958);
and U660 (N_660,In_1503,In_2185);
and U661 (N_661,In_148,In_2048);
nor U662 (N_662,In_2998,In_856);
nor U663 (N_663,In_2634,In_328);
xor U664 (N_664,In_1185,In_2773);
and U665 (N_665,In_1423,In_1439);
or U666 (N_666,In_1670,In_1155);
xor U667 (N_667,In_1904,In_490);
or U668 (N_668,In_1862,In_889);
nand U669 (N_669,In_2797,In_1046);
or U670 (N_670,In_1427,In_185);
nand U671 (N_671,In_1476,In_1559);
xnor U672 (N_672,In_1169,In_809);
or U673 (N_673,In_2155,In_1390);
nand U674 (N_674,In_1270,In_1987);
and U675 (N_675,In_1945,In_427);
and U676 (N_676,In_1699,In_2552);
or U677 (N_677,In_1665,In_36);
nand U678 (N_678,In_2899,In_542);
or U679 (N_679,In_2340,In_676);
nand U680 (N_680,In_728,In_2154);
or U681 (N_681,In_1788,In_2160);
nor U682 (N_682,In_848,In_173);
and U683 (N_683,In_2232,In_1098);
nor U684 (N_684,In_2216,In_2492);
xor U685 (N_685,In_796,In_2975);
xor U686 (N_686,In_2019,In_34);
and U687 (N_687,In_750,In_409);
and U688 (N_688,In_1419,In_2260);
nand U689 (N_689,In_380,In_2062);
and U690 (N_690,In_2635,In_1449);
and U691 (N_691,In_2697,In_2519);
nand U692 (N_692,In_2420,In_732);
or U693 (N_693,In_421,In_1602);
xnor U694 (N_694,In_2853,In_24);
or U695 (N_695,In_270,In_1624);
nand U696 (N_696,In_921,In_1363);
nor U697 (N_697,In_1963,In_651);
nor U698 (N_698,In_1446,In_1399);
xnor U699 (N_699,In_2759,In_528);
and U700 (N_700,In_98,In_1759);
and U701 (N_701,In_2132,In_1848);
and U702 (N_702,In_863,In_2415);
nor U703 (N_703,In_600,In_1671);
nand U704 (N_704,In_1889,In_1340);
nor U705 (N_705,In_228,In_1411);
nor U706 (N_706,In_211,In_1888);
or U707 (N_707,In_182,In_962);
and U708 (N_708,In_568,In_65);
and U709 (N_709,In_178,In_2040);
xnor U710 (N_710,In_467,In_1937);
nand U711 (N_711,In_1902,In_2337);
nand U712 (N_712,In_2891,In_1985);
or U713 (N_713,In_1690,In_242);
and U714 (N_714,In_189,In_1295);
xnor U715 (N_715,In_2325,In_2458);
or U716 (N_716,In_1536,In_752);
or U717 (N_717,In_2191,In_1601);
nand U718 (N_718,In_1349,In_875);
nand U719 (N_719,In_266,In_1786);
xnor U720 (N_720,In_1280,In_1763);
xnor U721 (N_721,In_2351,In_1003);
xor U722 (N_722,In_2505,In_2212);
and U723 (N_723,In_1067,In_787);
and U724 (N_724,In_855,In_295);
nand U725 (N_725,In_636,In_2161);
and U726 (N_726,In_2560,In_350);
or U727 (N_727,In_2841,In_2823);
or U728 (N_728,In_2262,In_2754);
xor U729 (N_729,In_2738,In_917);
xor U730 (N_730,In_2047,In_2804);
xnor U731 (N_731,In_913,In_1162);
xor U732 (N_732,In_2601,In_2626);
nor U733 (N_733,In_1422,In_1222);
nand U734 (N_734,In_2119,In_457);
xnor U735 (N_735,In_1348,In_2408);
or U736 (N_736,In_2942,In_2293);
and U737 (N_737,In_2554,In_1693);
or U738 (N_738,In_1766,In_1402);
nor U739 (N_739,In_1580,In_1395);
nand U740 (N_740,In_2913,In_1627);
nor U741 (N_741,In_935,In_2033);
or U742 (N_742,In_2373,In_2581);
or U743 (N_743,In_2171,In_2659);
xnor U744 (N_744,In_2423,In_510);
xnor U745 (N_745,In_2353,In_1408);
nand U746 (N_746,In_805,In_1313);
and U747 (N_747,In_2966,In_882);
nor U748 (N_748,In_1505,In_925);
xnor U749 (N_749,In_2650,In_240);
and U750 (N_750,In_2389,In_2778);
and U751 (N_751,In_2183,In_1875);
nor U752 (N_752,In_2365,In_558);
and U753 (N_753,In_1377,In_942);
or U754 (N_754,In_216,In_1358);
and U755 (N_755,In_527,In_2911);
nand U756 (N_756,In_259,In_881);
xnor U757 (N_757,In_695,In_2339);
nor U758 (N_758,In_618,In_2915);
and U759 (N_759,In_1979,In_2706);
and U760 (N_760,In_1715,In_2827);
xor U761 (N_761,In_680,In_2108);
nand U762 (N_762,In_2944,In_239);
xnor U763 (N_763,In_2100,In_62);
xnor U764 (N_764,In_551,In_1437);
nand U765 (N_765,In_7,In_1596);
nor U766 (N_766,In_2179,In_2657);
or U767 (N_767,In_736,In_2319);
and U768 (N_768,In_2345,In_2860);
and U769 (N_769,In_1466,In_2058);
nor U770 (N_770,In_2055,In_114);
and U771 (N_771,In_1701,In_2441);
nor U772 (N_772,In_960,In_2469);
xor U773 (N_773,In_1093,In_1158);
nand U774 (N_774,In_2156,In_2442);
nor U775 (N_775,In_2828,In_2525);
xor U776 (N_776,In_1831,In_1942);
nor U777 (N_777,In_1544,In_741);
nand U778 (N_778,In_899,In_562);
and U779 (N_779,In_774,In_1986);
nand U780 (N_780,In_2810,In_2176);
nor U781 (N_781,In_1109,In_198);
nor U782 (N_782,In_737,In_1207);
nand U783 (N_783,In_1895,In_916);
nand U784 (N_784,In_2323,In_2645);
nand U785 (N_785,In_2411,In_2703);
and U786 (N_786,In_1489,In_2187);
or U787 (N_787,In_1151,In_738);
xnor U788 (N_788,In_43,In_2144);
xnor U789 (N_789,In_1621,In_586);
and U790 (N_790,In_2010,In_784);
nand U791 (N_791,In_773,In_1646);
nand U792 (N_792,In_1546,In_888);
and U793 (N_793,In_1102,In_1460);
nand U794 (N_794,In_1242,In_1220);
nor U795 (N_795,In_2046,In_1745);
nand U796 (N_796,In_1085,In_658);
and U797 (N_797,In_611,In_890);
nor U798 (N_798,In_1725,In_2464);
or U799 (N_799,In_2005,In_937);
nand U800 (N_800,In_1171,In_2098);
nand U801 (N_801,In_1513,In_967);
and U802 (N_802,In_667,In_1118);
nor U803 (N_803,In_885,In_1833);
nand U804 (N_804,In_2662,In_923);
nor U805 (N_805,In_546,In_254);
or U806 (N_806,In_1005,In_480);
or U807 (N_807,In_866,In_1685);
xor U808 (N_808,In_272,In_669);
nand U809 (N_809,In_1181,In_1447);
or U810 (N_810,In_1127,In_670);
xnor U811 (N_811,In_2517,In_2597);
nor U812 (N_812,In_106,In_276);
xor U813 (N_813,In_2686,In_125);
nand U814 (N_814,In_2599,In_2483);
xor U815 (N_815,In_1147,In_2346);
xnor U816 (N_816,In_1824,In_180);
or U817 (N_817,In_249,In_2235);
nand U818 (N_818,In_1125,In_1434);
nand U819 (N_819,In_585,In_2474);
nand U820 (N_820,In_1706,In_1054);
nor U821 (N_821,In_2746,In_2395);
nor U822 (N_822,In_121,In_1076);
nor U823 (N_823,In_2935,In_105);
nor U824 (N_824,In_330,In_428);
or U825 (N_825,In_11,In_1487);
xnor U826 (N_826,In_601,In_59);
xnor U827 (N_827,In_1368,In_565);
nor U828 (N_828,In_1575,In_2403);
xnor U829 (N_829,In_2752,In_1225);
nand U830 (N_830,In_280,In_973);
xnor U831 (N_831,In_560,In_23);
or U832 (N_832,In_2655,In_1322);
nor U833 (N_833,In_1993,In_398);
nand U834 (N_834,In_48,In_235);
nor U835 (N_835,In_2446,In_1081);
nor U836 (N_836,In_2753,In_1642);
nor U837 (N_837,In_207,In_2394);
nor U838 (N_838,In_1100,In_364);
nor U839 (N_839,In_2150,In_1879);
or U840 (N_840,In_2252,In_357);
nand U841 (N_841,In_2101,In_2170);
nand U842 (N_842,In_2729,In_2082);
and U843 (N_843,In_2892,In_449);
or U844 (N_844,In_2349,In_1229);
and U845 (N_845,In_1550,In_2748);
and U846 (N_846,In_1260,In_2111);
nand U847 (N_847,In_111,In_1318);
nor U848 (N_848,In_2460,In_2945);
and U849 (N_849,In_1033,In_92);
nand U850 (N_850,In_2561,In_543);
or U851 (N_851,In_1574,In_2159);
nand U852 (N_852,In_803,In_706);
xnor U853 (N_853,In_1378,In_1710);
or U854 (N_854,In_1435,In_2362);
and U855 (N_855,In_1709,In_2570);
xnor U856 (N_856,In_1045,In_2205);
or U857 (N_857,In_82,In_2529);
nand U858 (N_858,In_2390,In_396);
or U859 (N_859,In_298,In_2871);
nand U860 (N_860,In_1099,In_1104);
nor U861 (N_861,In_104,In_2854);
nor U862 (N_862,In_799,In_928);
xnor U863 (N_863,In_2121,In_1682);
nand U864 (N_864,In_2064,In_2106);
xnor U865 (N_865,In_2025,In_268);
nor U866 (N_866,In_2015,In_1038);
and U867 (N_867,In_1523,In_288);
xnor U868 (N_868,In_1598,In_2455);
and U869 (N_869,In_2214,In_2368);
and U870 (N_870,In_2756,In_1326);
and U871 (N_871,In_640,In_2088);
or U872 (N_872,In_1955,In_1617);
xor U873 (N_873,In_1430,In_2562);
nor U874 (N_874,In_2419,In_2585);
xor U875 (N_875,In_2855,In_2409);
nor U876 (N_876,In_30,In_1188);
nor U877 (N_877,In_717,In_2104);
xor U878 (N_878,In_2669,In_18);
xor U879 (N_879,In_646,In_1077);
xnor U880 (N_880,In_845,In_2427);
nor U881 (N_881,In_2948,In_2783);
xnor U882 (N_882,In_2665,In_981);
and U883 (N_883,In_347,In_2036);
xnor U884 (N_884,In_664,In_145);
nor U885 (N_885,In_1948,In_1486);
and U886 (N_886,In_205,In_1305);
or U887 (N_887,In_1425,In_1645);
nor U888 (N_888,In_2963,In_1753);
xor U889 (N_889,In_2146,In_2137);
nand U890 (N_890,In_1908,In_1194);
nand U891 (N_891,In_2453,In_2507);
nor U892 (N_892,In_432,In_221);
or U893 (N_893,In_2618,In_1330);
nand U894 (N_894,In_1498,In_394);
xnor U895 (N_895,In_2324,In_17);
nor U896 (N_896,In_2375,In_1921);
xor U897 (N_897,In_1886,In_187);
xnor U898 (N_898,In_1563,In_633);
and U899 (N_899,In_753,In_353);
or U900 (N_900,In_2248,In_721);
nand U901 (N_901,In_2473,In_355);
nand U902 (N_902,In_1053,In_1414);
or U903 (N_903,In_1392,In_172);
or U904 (N_904,In_1885,In_1980);
nand U905 (N_905,In_992,In_930);
and U906 (N_906,In_1142,In_138);
or U907 (N_907,In_878,In_2835);
or U908 (N_908,In_337,In_1376);
or U909 (N_909,In_836,In_2264);
or U910 (N_910,In_346,In_1030);
xor U911 (N_911,In_2498,In_2950);
and U912 (N_912,In_81,In_47);
xor U913 (N_913,In_1769,In_265);
xnor U914 (N_914,In_1195,In_2091);
xor U915 (N_915,In_2932,In_1156);
xnor U916 (N_916,In_1051,In_2127);
nor U917 (N_917,In_2434,In_628);
or U918 (N_918,In_950,In_1457);
or U919 (N_919,In_1809,In_1719);
nor U920 (N_920,In_549,In_2629);
or U921 (N_921,In_868,In_2580);
xor U922 (N_922,In_2751,In_1810);
nand U923 (N_923,In_2920,In_1876);
nand U924 (N_924,In_2745,In_218);
nand U925 (N_925,In_1214,In_2045);
nor U926 (N_926,In_2606,In_2666);
and U927 (N_927,In_1356,In_1827);
nor U928 (N_928,In_1172,In_1035);
and U929 (N_929,In_35,In_2876);
nand U930 (N_930,In_361,In_1610);
nor U931 (N_931,In_1112,In_1620);
nand U932 (N_932,In_909,In_2543);
xnor U933 (N_933,In_1201,In_296);
nand U934 (N_934,In_1882,In_1210);
or U935 (N_935,In_77,In_590);
or U936 (N_936,In_2110,In_2398);
and U937 (N_937,In_2996,In_1293);
or U938 (N_938,In_840,In_2245);
nand U939 (N_939,In_1004,In_2786);
nand U940 (N_940,In_2124,In_1560);
xnor U941 (N_941,In_2463,In_499);
and U942 (N_942,In_2683,In_2641);
nand U943 (N_943,In_1346,In_843);
nor U944 (N_944,In_757,In_1006);
xor U945 (N_945,In_2491,In_1286);
or U946 (N_946,In_1731,In_627);
and U947 (N_947,In_1919,In_379);
and U948 (N_948,In_1416,In_2604);
nor U949 (N_949,In_822,In_208);
xnor U950 (N_950,In_841,In_2776);
or U951 (N_951,In_2802,In_1017);
nor U952 (N_952,In_2520,In_907);
and U953 (N_953,In_612,In_2044);
xnor U954 (N_954,In_359,In_297);
nand U955 (N_955,In_1168,In_468);
nand U956 (N_956,In_2528,In_1521);
or U957 (N_957,In_389,In_2825);
or U958 (N_958,In_434,In_2425);
and U959 (N_959,In_140,In_789);
and U960 (N_960,In_2710,In_255);
nor U961 (N_961,In_500,In_1197);
and U962 (N_962,In_2903,In_2060);
xnor U963 (N_963,In_212,In_441);
nor U964 (N_964,In_241,In_710);
nand U965 (N_965,In_2437,In_1807);
xnor U966 (N_966,In_1911,In_1490);
xor U967 (N_967,In_603,In_1913);
and U968 (N_968,In_2627,In_2930);
or U969 (N_969,In_2147,In_343);
nor U970 (N_970,In_2577,In_858);
or U971 (N_971,In_2276,In_310);
nor U972 (N_972,In_1271,In_993);
xor U973 (N_973,In_2244,In_1778);
nor U974 (N_974,In_424,In_1101);
and U975 (N_975,In_842,In_1415);
and U976 (N_976,In_1989,In_2094);
and U977 (N_977,In_40,In_1808);
or U978 (N_978,In_832,In_1131);
xnor U979 (N_979,In_532,In_2280);
nand U980 (N_980,In_1849,In_2768);
and U981 (N_981,In_772,In_631);
and U982 (N_982,In_1205,In_2071);
and U983 (N_983,In_1149,In_1933);
or U984 (N_984,In_1057,In_1868);
and U985 (N_985,In_743,In_1484);
xor U986 (N_986,In_2796,In_1397);
xnor U987 (N_987,In_2907,In_978);
nor U988 (N_988,In_1656,In_1618);
and U989 (N_989,In_540,In_2197);
nand U990 (N_990,In_2671,In_2461);
xor U991 (N_991,In_665,In_2360);
and U992 (N_992,In_2301,In_2779);
and U993 (N_993,In_2311,In_1832);
and U994 (N_994,In_1413,In_2934);
xnor U995 (N_995,In_2863,In_2500);
nand U996 (N_996,In_1781,In_2977);
nor U997 (N_997,In_1049,In_1577);
nand U998 (N_998,In_926,In_1124);
and U999 (N_999,In_2451,In_920);
or U1000 (N_1000,N_682,In_2031);
nand U1001 (N_1001,N_564,In_1973);
nor U1002 (N_1002,N_405,In_642);
xor U1003 (N_1003,N_415,In_1774);
nand U1004 (N_1004,N_59,In_2506);
nor U1005 (N_1005,N_219,In_1552);
nor U1006 (N_1006,N_105,In_1134);
xnor U1007 (N_1007,In_411,N_749);
xnor U1008 (N_1008,N_681,In_2429);
nand U1009 (N_1009,In_1887,N_584);
or U1010 (N_1010,In_545,In_1406);
nor U1011 (N_1011,In_1512,In_2598);
xor U1012 (N_1012,In_436,In_643);
or U1013 (N_1013,N_407,In_2480);
xnor U1014 (N_1014,In_1209,N_756);
xor U1015 (N_1015,In_834,In_557);
or U1016 (N_1016,In_1724,N_347);
and U1017 (N_1017,N_947,N_959);
or U1018 (N_1018,In_282,N_953);
or U1019 (N_1019,In_1901,N_905);
or U1020 (N_1020,N_689,In_139);
nor U1021 (N_1021,N_15,N_208);
or U1022 (N_1022,In_902,N_739);
nor U1023 (N_1023,N_424,N_194);
xor U1024 (N_1024,N_439,N_534);
xor U1025 (N_1025,In_2997,N_671);
and U1026 (N_1026,In_1291,In_2979);
or U1027 (N_1027,In_949,In_2808);
nand U1028 (N_1028,In_257,N_805);
xor U1029 (N_1029,In_2217,N_256);
nor U1030 (N_1030,In_2766,In_2050);
nor U1031 (N_1031,In_786,In_0);
nand U1032 (N_1032,N_381,In_2254);
and U1033 (N_1033,In_2734,N_449);
nand U1034 (N_1034,In_1328,In_137);
nor U1035 (N_1035,N_538,In_948);
nand U1036 (N_1036,N_241,N_275);
xor U1037 (N_1037,N_984,In_2586);
and U1038 (N_1038,In_2422,N_127);
nor U1039 (N_1039,In_1236,N_317);
nor U1040 (N_1040,In_2949,N_448);
xor U1041 (N_1041,In_972,N_459);
nand U1042 (N_1042,In_483,N_206);
and U1043 (N_1043,N_40,In_1176);
and U1044 (N_1044,In_966,In_2444);
nor U1045 (N_1045,N_986,In_564);
or U1046 (N_1046,N_606,N_556);
and U1047 (N_1047,In_1522,N_997);
nand U1048 (N_1048,N_649,N_164);
xor U1049 (N_1049,In_2135,In_1259);
or U1050 (N_1050,N_622,N_142);
nor U1051 (N_1051,N_304,N_234);
nor U1052 (N_1052,N_670,In_1953);
nor U1053 (N_1053,In_1442,In_291);
and U1054 (N_1054,In_2484,N_875);
nand U1055 (N_1055,N_550,In_2273);
and U1056 (N_1056,In_1650,N_460);
or U1057 (N_1057,In_2043,In_1367);
xor U1058 (N_1058,In_2396,In_167);
nand U1059 (N_1059,In_1834,N_532);
or U1060 (N_1060,In_523,In_632);
nand U1061 (N_1061,N_829,N_627);
xnor U1062 (N_1062,N_176,N_854);
and U1063 (N_1063,In_1223,In_384);
xor U1064 (N_1064,In_2295,In_1237);
and U1065 (N_1065,In_802,N_477);
or U1066 (N_1066,N_966,N_189);
nand U1067 (N_1067,In_2263,N_510);
xor U1068 (N_1068,In_893,In_1464);
and U1069 (N_1069,N_714,In_1880);
nand U1070 (N_1070,N_620,N_363);
nand U1071 (N_1071,In_2872,N_675);
nor U1072 (N_1072,N_560,N_161);
nand U1073 (N_1073,In_1830,In_1389);
nor U1074 (N_1074,N_549,In_2978);
xor U1075 (N_1075,N_131,N_95);
xor U1076 (N_1076,In_1020,N_143);
nor U1077 (N_1077,In_607,In_1075);
and U1078 (N_1078,In_2439,N_170);
or U1079 (N_1079,N_83,N_154);
nor U1080 (N_1080,In_535,N_987);
and U1081 (N_1081,N_96,In_1496);
or U1082 (N_1082,In_2432,In_1729);
and U1083 (N_1083,N_245,N_404);
nand U1084 (N_1084,In_1691,N_438);
or U1085 (N_1085,In_825,N_691);
nor U1086 (N_1086,In_238,In_617);
and U1087 (N_1087,N_557,In_1047);
nand U1088 (N_1088,N_937,N_529);
nand U1089 (N_1089,In_2114,In_447);
nand U1090 (N_1090,In_2128,In_1272);
nor U1091 (N_1091,N_158,N_904);
nor U1092 (N_1092,In_661,N_846);
and U1093 (N_1093,N_686,In_1924);
or U1094 (N_1094,N_802,In_678);
nor U1095 (N_1095,In_1768,In_1938);
nor U1096 (N_1096,In_963,N_777);
nand U1097 (N_1097,In_2238,N_299);
nand U1098 (N_1098,In_594,N_737);
nand U1099 (N_1099,N_362,In_313);
nor U1100 (N_1100,N_361,N_284);
and U1101 (N_1101,N_64,In_1329);
and U1102 (N_1102,In_1115,N_352);
xnor U1103 (N_1103,In_1308,In_1037);
xnor U1104 (N_1104,In_767,N_168);
nand U1105 (N_1105,N_43,In_699);
or U1106 (N_1106,N_778,In_2603);
nor U1107 (N_1107,In_1694,In_1055);
nand U1108 (N_1108,In_1949,N_588);
nor U1109 (N_1109,In_1309,N_48);
or U1110 (N_1110,N_166,In_1797);
or U1111 (N_1111,N_853,N_456);
nor U1112 (N_1112,In_2092,In_2304);
nor U1113 (N_1113,In_2912,N_630);
or U1114 (N_1114,In_904,In_136);
or U1115 (N_1115,In_2820,In_2839);
and U1116 (N_1116,N_963,In_1728);
xor U1117 (N_1117,N_874,In_284);
or U1118 (N_1118,In_2933,In_2149);
or U1119 (N_1119,In_2386,N_491);
nand U1120 (N_1120,N_396,In_1932);
or U1121 (N_1121,In_798,N_278);
xor U1122 (N_1122,N_791,N_25);
or U1123 (N_1123,In_2333,In_2858);
and U1124 (N_1124,N_619,In_404);
nor U1125 (N_1125,In_1007,In_691);
nand U1126 (N_1126,In_273,N_835);
and U1127 (N_1127,N_625,In_1183);
nor U1128 (N_1128,In_2059,In_2557);
xor U1129 (N_1129,N_787,N_740);
nor U1130 (N_1130,N_962,N_933);
nand U1131 (N_1131,In_954,In_1015);
xnor U1132 (N_1132,N_608,N_667);
xor U1133 (N_1133,In_2727,In_588);
nand U1134 (N_1134,In_2656,N_437);
xnor U1135 (N_1135,In_2594,In_2285);
and U1136 (N_1136,N_581,N_523);
nor U1137 (N_1137,In_755,In_190);
xnor U1138 (N_1138,N_928,N_772);
or U1139 (N_1139,N_900,In_1381);
nand U1140 (N_1140,N_697,N_162);
or U1141 (N_1141,In_1213,In_437);
and U1142 (N_1142,N_497,In_2037);
nor U1143 (N_1143,N_748,In_1023);
and U1144 (N_1144,In_1206,In_1091);
xnor U1145 (N_1145,N_809,In_2095);
nand U1146 (N_1146,N_935,In_2210);
or U1147 (N_1147,In_33,N_475);
nor U1148 (N_1148,N_653,In_1751);
nor U1149 (N_1149,N_988,N_723);
nand U1150 (N_1150,In_2893,In_2620);
or U1151 (N_1151,N_521,In_2764);
or U1152 (N_1152,In_2719,N_688);
nor U1153 (N_1153,In_1755,In_2361);
xnor U1154 (N_1154,In_1016,In_1086);
or U1155 (N_1155,In_1556,N_42);
and U1156 (N_1156,N_86,N_145);
nor U1157 (N_1157,N_328,N_231);
nand U1158 (N_1158,N_906,N_629);
nand U1159 (N_1159,N_146,N_470);
nor U1160 (N_1160,In_127,In_1410);
xor U1161 (N_1161,In_2591,In_851);
nand U1162 (N_1162,N_609,In_1988);
nand U1163 (N_1163,N_747,In_2989);
and U1164 (N_1164,In_1883,In_2664);
nand U1165 (N_1165,In_2851,N_893);
and U1166 (N_1166,N_401,N_598);
and U1167 (N_1167,N_762,N_792);
and U1168 (N_1168,In_475,N_885);
nand U1169 (N_1169,N_499,N_775);
or U1170 (N_1170,N_3,In_1059);
or U1171 (N_1171,In_2757,N_199);
nor U1172 (N_1172,In_2685,In_687);
or U1173 (N_1173,In_1520,N_218);
xor U1174 (N_1174,N_482,In_14);
nor U1175 (N_1175,N_165,In_210);
nor U1176 (N_1176,N_98,In_2343);
nand U1177 (N_1177,N_29,N_215);
xor U1178 (N_1178,N_57,N_376);
nor U1179 (N_1179,N_298,N_952);
or U1180 (N_1180,In_739,N_23);
xor U1181 (N_1181,In_1812,In_1805);
or U1182 (N_1182,N_728,In_1244);
nor U1183 (N_1183,In_340,In_1268);
and U1184 (N_1184,In_2558,N_335);
or U1185 (N_1185,N_472,In_2013);
nor U1186 (N_1186,In_644,In_1966);
nand U1187 (N_1187,N_274,In_1740);
nand U1188 (N_1188,N_996,In_1456);
nand U1189 (N_1189,N_827,In_2359);
or U1190 (N_1190,In_1957,In_2272);
or U1191 (N_1191,In_2310,In_1915);
nor U1192 (N_1192,In_2595,N_80);
nand U1193 (N_1193,In_2993,In_2816);
and U1194 (N_1194,N_876,N_295);
and U1195 (N_1195,In_2123,N_110);
or U1196 (N_1196,N_204,In_2771);
nand U1197 (N_1197,N_440,N_950);
nor U1198 (N_1198,In_970,N_195);
nor U1199 (N_1199,In_1846,N_55);
xnor U1200 (N_1200,N_706,N_500);
nor U1201 (N_1201,In_1592,N_799);
xor U1202 (N_1202,N_724,In_1961);
nand U1203 (N_1203,N_857,In_577);
xor U1204 (N_1204,N_708,N_350);
xor U1205 (N_1205,In_1357,N_569);
or U1206 (N_1206,In_312,N_4);
and U1207 (N_1207,N_559,In_625);
xor U1208 (N_1208,N_153,In_2897);
and U1209 (N_1209,In_1289,N_602);
and U1210 (N_1210,N_30,In_381);
nor U1211 (N_1211,N_610,N_578);
and U1212 (N_1212,N_931,N_710);
or U1213 (N_1213,N_377,In_2831);
xnor U1214 (N_1214,N_21,In_1784);
or U1215 (N_1215,In_2637,N_591);
nor U1216 (N_1216,N_938,N_993);
nor U1217 (N_1217,In_2731,In_666);
or U1218 (N_1218,N_561,In_1064);
or U1219 (N_1219,N_54,N_616);
or U1220 (N_1220,In_122,In_2857);
and U1221 (N_1221,N_895,N_862);
nand U1222 (N_1222,In_762,N_109);
xnor U1223 (N_1223,In_1432,In_518);
nor U1224 (N_1224,N_695,In_2003);
xnor U1225 (N_1225,N_280,In_2231);
nand U1226 (N_1226,N_640,In_319);
nor U1227 (N_1227,In_2452,In_429);
nor U1228 (N_1228,In_474,In_1087);
nand U1229 (N_1229,In_2873,In_2297);
xnor U1230 (N_1230,In_919,N_253);
and U1231 (N_1231,In_3,N_157);
xor U1232 (N_1232,In_383,In_1227);
and U1233 (N_1233,N_468,In_377);
and U1234 (N_1234,N_97,In_410);
or U1235 (N_1235,N_908,In_521);
xnor U1236 (N_1236,In_1571,N_650);
or U1237 (N_1237,N_832,In_1777);
or U1238 (N_1238,In_2767,In_445);
or U1239 (N_1239,In_2070,In_333);
xnor U1240 (N_1240,N_180,In_2985);
xnor U1241 (N_1241,In_2448,N_845);
nor U1242 (N_1242,N_287,In_1288);
xor U1243 (N_1243,In_91,N_979);
or U1244 (N_1244,N_150,N_509);
or U1245 (N_1245,In_2312,In_2456);
and U1246 (N_1246,In_2687,N_301);
nor U1247 (N_1247,In_2982,In_1964);
xnor U1248 (N_1248,N_956,In_417);
xor U1249 (N_1249,N_882,N_364);
and U1250 (N_1250,In_143,N_782);
and U1251 (N_1251,In_994,In_2574);
nand U1252 (N_1252,N_525,N_156);
xnor U1253 (N_1253,In_2251,N_998);
nor U1254 (N_1254,In_912,In_2589);
nor U1255 (N_1255,In_1455,In_574);
or U1256 (N_1256,In_219,N_93);
and U1257 (N_1257,N_319,In_2027);
xor U1258 (N_1258,In_2972,N_541);
xor U1259 (N_1259,N_0,In_2334);
xnor U1260 (N_1260,N_50,In_1248);
nand U1261 (N_1261,In_1998,N_112);
and U1262 (N_1262,N_248,In_2681);
or U1263 (N_1263,N_639,N_453);
nand U1264 (N_1264,In_423,In_544);
or U1265 (N_1265,In_2152,In_414);
nor U1266 (N_1266,N_634,In_2673);
nand U1267 (N_1267,In_1226,In_152);
nor U1268 (N_1268,In_460,N_160);
xnor U1269 (N_1269,In_477,N_949);
and U1270 (N_1270,In_872,N_213);
xnor U1271 (N_1271,N_467,In_2042);
or U1272 (N_1272,N_228,In_1353);
nand U1273 (N_1273,In_936,In_1337);
or U1274 (N_1274,N_191,In_2600);
nand U1275 (N_1275,N_327,In_623);
nand U1276 (N_1276,In_1564,N_599);
nand U1277 (N_1277,In_481,In_2798);
xnor U1278 (N_1278,In_487,N_912);
or U1279 (N_1279,N_251,N_261);
and U1280 (N_1280,In_2732,N_542);
or U1281 (N_1281,N_957,N_555);
nand U1282 (N_1282,N_436,N_849);
and U1283 (N_1283,N_891,In_2805);
nor U1284 (N_1284,N_519,N_801);
nand U1285 (N_1285,N_265,N_767);
nor U1286 (N_1286,N_431,N_694);
nor U1287 (N_1287,N_575,In_217);
xnor U1288 (N_1288,N_693,N_51);
xor U1289 (N_1289,In_58,N_202);
or U1290 (N_1290,N_973,In_2782);
nand U1291 (N_1291,In_770,N_883);
nand U1292 (N_1292,N_547,In_609);
or U1293 (N_1293,In_1934,N_994);
nor U1294 (N_1294,N_626,In_2693);
xnor U1295 (N_1295,N_461,In_847);
or U1296 (N_1296,N_886,N_445);
and U1297 (N_1297,N_267,In_1379);
and U1298 (N_1298,In_2402,N_426);
or U1299 (N_1299,In_2631,In_626);
or U1300 (N_1300,N_669,In_686);
or U1301 (N_1301,N_184,N_577);
xor U1302 (N_1302,In_2705,In_253);
or U1303 (N_1303,In_170,N_340);
nor U1304 (N_1304,In_220,N_786);
nor U1305 (N_1305,N_585,N_508);
or U1306 (N_1306,N_249,In_1341);
xor U1307 (N_1307,N_824,In_806);
nand U1308 (N_1308,In_153,In_426);
xor U1309 (N_1309,In_150,N_66);
xnor U1310 (N_1310,In_539,N_655);
xnor U1311 (N_1311,In_1391,N_137);
nor U1312 (N_1312,N_2,In_1900);
nand U1313 (N_1313,N_360,N_932);
nand U1314 (N_1314,N_858,N_394);
and U1315 (N_1315,In_2486,N_727);
nor U1316 (N_1316,N_818,N_188);
nor U1317 (N_1317,In_2079,N_53);
or U1318 (N_1318,N_969,N_924);
nand U1319 (N_1319,N_387,N_659);
or U1320 (N_1320,In_2736,N_763);
and U1321 (N_1321,In_2566,N_712);
nand U1322 (N_1322,In_1495,In_567);
nand U1323 (N_1323,In_203,N_624);
nand U1324 (N_1324,In_2120,N_114);
nand U1325 (N_1325,N_526,N_911);
and U1326 (N_1326,N_128,In_25);
nor U1327 (N_1327,N_38,N_964);
nor U1328 (N_1328,N_582,In_813);
and U1329 (N_1329,N_558,N_781);
nor U1330 (N_1330,In_482,In_2493);
nand U1331 (N_1331,N_915,In_785);
or U1332 (N_1332,N_735,N_149);
and U1333 (N_1333,In_1469,In_1705);
xnor U1334 (N_1334,In_1451,N_32);
nand U1335 (N_1335,In_2417,In_1840);
and U1336 (N_1336,N_31,In_1524);
nor U1337 (N_1337,In_2838,In_374);
nor U1338 (N_1338,N_85,N_971);
xor U1339 (N_1339,N_631,In_1107);
xnor U1340 (N_1340,N_117,N_917);
and U1341 (N_1341,In_64,In_563);
nand U1342 (N_1342,N_663,In_1347);
nand U1343 (N_1343,N_921,In_2700);
nand U1344 (N_1344,In_634,N_201);
xnor U1345 (N_1345,In_731,N_785);
xnor U1346 (N_1346,In_1946,N_118);
xnor U1347 (N_1347,In_2539,N_894);
xnor U1348 (N_1348,In_1782,N_13);
or U1349 (N_1349,N_305,N_730);
or U1350 (N_1350,N_243,In_2714);
or U1351 (N_1351,In_2840,In_2126);
nor U1352 (N_1352,In_2521,In_2888);
nand U1353 (N_1353,N_435,N_540);
xor U1354 (N_1354,In_1543,In_2611);
xor U1355 (N_1355,N_719,In_2937);
nor U1356 (N_1356,In_526,N_613);
and U1357 (N_1357,N_263,In_1614);
and U1358 (N_1358,N_567,In_2299);
xor U1359 (N_1359,N_193,In_2054);
and U1360 (N_1360,N_684,N_545);
and U1361 (N_1361,In_1903,N_746);
and U1362 (N_1362,In_329,N_339);
or U1363 (N_1363,N_185,N_122);
nor U1364 (N_1364,In_1461,N_873);
xnor U1365 (N_1365,In_553,In_2130);
nand U1366 (N_1366,N_152,N_77);
or U1367 (N_1367,N_553,N_830);
nor U1368 (N_1368,In_2298,N_410);
xnor U1369 (N_1369,N_722,N_484);
nor U1370 (N_1370,In_1400,In_351);
nand U1371 (N_1371,N_637,In_13);
or U1372 (N_1372,In_1137,N_18);
and U1373 (N_1373,N_985,In_1586);
and U1374 (N_1374,N_779,N_863);
nand U1375 (N_1375,N_812,N_67);
or U1376 (N_1376,N_896,In_1036);
and U1377 (N_1377,N_738,N_187);
and U1378 (N_1378,In_6,In_299);
and U1379 (N_1379,In_2575,In_169);
xor U1380 (N_1380,In_1718,N_690);
nor U1381 (N_1381,In_177,N_923);
nor U1382 (N_1382,N_447,N_539);
nor U1383 (N_1383,N_133,N_443);
nand U1384 (N_1384,In_1361,In_439);
nor U1385 (N_1385,In_1954,N_621);
or U1386 (N_1386,N_378,In_1360);
and U1387 (N_1387,N_74,In_2009);
nand U1388 (N_1388,N_565,In_335);
xnor U1389 (N_1389,In_267,In_826);
and U1390 (N_1390,N_797,In_2845);
xnor U1391 (N_1391,In_2296,N_715);
nor U1392 (N_1392,N_399,In_1375);
or U1393 (N_1393,In_1278,In_2874);
or U1394 (N_1394,In_262,In_2647);
nand U1395 (N_1395,N_236,N_246);
nand U1396 (N_1396,In_2305,In_2952);
xor U1397 (N_1397,N_179,In_2898);
and U1398 (N_1398,In_1982,In_608);
and U1399 (N_1399,N_342,In_671);
or U1400 (N_1400,In_197,N_125);
or U1401 (N_1401,In_2824,In_1359);
nand U1402 (N_1402,In_2961,In_602);
nand U1403 (N_1403,In_1983,N_418);
nor U1404 (N_1404,In_2544,N_496);
nand U1405 (N_1405,In_2074,In_2485);
or U1406 (N_1406,In_1657,In_2870);
and U1407 (N_1407,In_2391,In_674);
xor U1408 (N_1408,N_977,N_847);
nor U1409 (N_1409,N_600,N_276);
and U1410 (N_1410,N_934,N_713);
nand U1411 (N_1411,N_106,In_849);
or U1412 (N_1412,In_1783,N_61);
nand U1413 (N_1413,In_2097,In_2737);
nor U1414 (N_1414,In_1897,In_2923);
and U1415 (N_1415,N_868,N_103);
or U1416 (N_1416,In_709,In_808);
nor U1417 (N_1417,In_1345,N_186);
nand U1418 (N_1418,In_287,N_702);
nand U1419 (N_1419,N_850,N_413);
or U1420 (N_1420,N_692,In_1269);
nand U1421 (N_1421,N_828,N_825);
nor U1422 (N_1422,In_306,In_2057);
and U1423 (N_1423,In_2145,In_191);
nor U1424 (N_1424,N_623,N_768);
nor U1425 (N_1425,In_2668,N_795);
nand U1426 (N_1426,N_235,In_2369);
or U1427 (N_1427,N_593,N_306);
nand U1428 (N_1428,In_2918,In_1187);
xor U1429 (N_1429,N_752,N_607);
or U1430 (N_1430,In_1697,In_2674);
and U1431 (N_1431,N_991,N_878);
nand U1432 (N_1432,N_940,In_2006);
nand U1433 (N_1433,In_2971,N_411);
and U1434 (N_1434,N_658,N_877);
or U1435 (N_1435,In_2208,In_354);
nor U1436 (N_1436,N_469,N_196);
or U1437 (N_1437,N_326,N_704);
nand U1438 (N_1438,In_1689,N_220);
xnor U1439 (N_1439,N_331,N_790);
xnor U1440 (N_1440,N_212,N_592);
or U1441 (N_1441,N_349,N_200);
and U1442 (N_1442,In_2198,N_207);
nor U1443 (N_1443,In_2138,N_674);
and U1444 (N_1444,N_916,N_918);
nor U1445 (N_1445,N_776,N_155);
nand U1446 (N_1446,N_535,In_1285);
nand U1447 (N_1447,N_489,In_2760);
xor U1448 (N_1448,N_100,In_638);
or U1449 (N_1449,N_283,N_769);
xor U1450 (N_1450,In_19,In_2291);
or U1451 (N_1451,N_833,In_1152);
and U1452 (N_1452,In_52,N_119);
and U1453 (N_1453,In_969,N_88);
and U1454 (N_1454,N_974,In_908);
and U1455 (N_1455,N_107,In_2613);
and U1456 (N_1456,In_2022,In_444);
nor U1457 (N_1457,In_2919,In_1738);
nor U1458 (N_1458,In_2326,N_34);
and U1459 (N_1459,N_87,N_652);
nor U1460 (N_1460,In_2844,In_1095);
or U1461 (N_1461,In_406,N_594);
or U1462 (N_1462,In_1241,N_169);
or U1463 (N_1463,In_431,In_2663);
and U1464 (N_1464,In_823,In_1735);
nor U1465 (N_1465,In_1062,N_506);
nand U1466 (N_1466,N_182,N_473);
nand U1467 (N_1467,In_1984,N_409);
nand U1468 (N_1468,In_1547,N_380);
nand U1469 (N_1469,In_2307,In_689);
and U1470 (N_1470,N_576,N_851);
or U1471 (N_1471,N_580,N_548);
or U1472 (N_1472,N_60,In_965);
nor U1473 (N_1473,N_358,In_71);
xor U1474 (N_1474,N_343,N_595);
nor U1475 (N_1475,In_1041,In_32);
nor U1476 (N_1476,In_2698,In_294);
nor U1477 (N_1477,In_800,N_99);
and U1478 (N_1478,In_1233,In_400);
nand U1479 (N_1479,In_1090,In_2523);
nor U1480 (N_1480,N_803,N_229);
nor U1481 (N_1481,In_819,N_840);
xnor U1482 (N_1482,N_211,N_764);
and U1483 (N_1483,N_10,N_628);
nand U1484 (N_1484,N_941,In_1969);
and U1485 (N_1485,In_578,In_2765);
nor U1486 (N_1486,N_226,In_725);
nand U1487 (N_1487,In_1450,N_981);
nor U1488 (N_1488,N_741,N_351);
nor U1489 (N_1489,N_843,In_2109);
or U1490 (N_1490,N_820,N_699);
or U1491 (N_1491,In_1138,N_716);
or U1492 (N_1492,N_315,In_1727);
xnor U1493 (N_1493,N_841,In_1186);
and U1494 (N_1494,N_661,N_209);
nor U1495 (N_1495,N_672,In_2077);
nor U1496 (N_1496,In_690,In_2644);
nor U1497 (N_1497,In_1844,N_901);
nor U1498 (N_1498,N_960,In_2943);
and U1499 (N_1499,N_385,In_1756);
or U1500 (N_1500,N_141,N_861);
nand U1501 (N_1501,In_2352,N_992);
or U1502 (N_1502,In_1108,In_466);
and U1503 (N_1503,N_56,In_2536);
nor U1504 (N_1504,In_1956,N_210);
nand U1505 (N_1505,In_362,In_1585);
nor U1506 (N_1506,N_416,In_1116);
nand U1507 (N_1507,In_1507,N_33);
and U1508 (N_1508,N_839,N_913);
nor U1509 (N_1509,N_134,In_2530);
nand U1510 (N_1510,N_471,In_1533);
nor U1511 (N_1511,N_552,N_668);
and U1512 (N_1512,N_414,In_124);
and U1513 (N_1513,In_289,N_264);
or U1514 (N_1514,In_112,In_491);
xnor U1515 (N_1515,In_2481,N_909);
or U1516 (N_1516,In_635,N_403);
nand U1517 (N_1517,N_78,N_148);
nand U1518 (N_1518,In_2167,In_107);
or U1519 (N_1519,N_887,N_574);
and U1520 (N_1520,In_599,N_102);
and U1521 (N_1521,N_721,In_2157);
and U1522 (N_1522,N_700,In_1497);
xnor U1523 (N_1523,N_902,In_1746);
and U1524 (N_1524,N_94,N_603);
nand U1525 (N_1525,N_743,In_591);
and U1526 (N_1526,N_879,In_692);
nor U1527 (N_1527,In_2968,In_2141);
xor U1528 (N_1528,In_2125,N_124);
xor U1529 (N_1529,In_2462,N_174);
xor U1530 (N_1530,N_810,N_601);
and U1531 (N_1531,N_239,In_727);
nand U1532 (N_1532,N_753,N_572);
xor U1533 (N_1533,In_324,N_203);
xor U1534 (N_1534,N_89,In_712);
or U1535 (N_1535,N_451,In_862);
nand U1536 (N_1536,In_1212,In_1907);
xnor U1537 (N_1537,In_1120,In_1258);
or U1538 (N_1538,In_2267,N_462);
or U1539 (N_1539,In_1050,N_314);
or U1540 (N_1540,N_586,N_345);
nand U1541 (N_1541,N_808,N_866);
or U1542 (N_1542,N_222,N_217);
and U1543 (N_1543,In_318,N_823);
nand U1544 (N_1544,In_2286,In_2376);
nand U1545 (N_1545,In_2954,N_494);
or U1546 (N_1546,In_2545,In_2065);
or U1547 (N_1547,In_1864,In_1509);
nand U1548 (N_1548,In_1643,N_698);
nor U1549 (N_1549,In_2501,In_386);
xnor U1550 (N_1550,N_546,N_47);
nand U1551 (N_1551,N_371,In_572);
or U1552 (N_1552,N_726,N_837);
and U1553 (N_1553,N_943,In_1525);
nor U1554 (N_1554,N_766,In_375);
or U1555 (N_1555,N_951,N_22);
nand U1556 (N_1556,In_924,N_198);
and U1557 (N_1557,In_1472,N_238);
or U1558 (N_1558,In_780,In_1089);
nand U1559 (N_1559,In_147,In_894);
and U1560 (N_1560,N_814,In_1336);
nor U1561 (N_1561,N_501,N_811);
xor U1562 (N_1562,In_1678,In_1703);
nor U1563 (N_1563,In_2829,In_2471);
xnor U1564 (N_1564,N_230,N_505);
and U1565 (N_1565,In_1637,In_1230);
or U1566 (N_1566,In_1355,In_873);
nand U1567 (N_1567,In_2541,N_566);
nand U1568 (N_1568,In_579,N_914);
or U1569 (N_1569,In_827,In_26);
xor U1570 (N_1570,In_953,In_726);
and U1571 (N_1571,In_2220,N_975);
xnor U1572 (N_1572,N_58,In_237);
nand U1573 (N_1573,N_257,N_664);
nor U1574 (N_1574,In_352,In_161);
or U1575 (N_1575,In_2849,N_750);
nor U1576 (N_1576,N_259,In_1663);
xnor U1577 (N_1577,In_1198,In_1365);
and U1578 (N_1578,N_270,N_742);
nand U1579 (N_1579,N_375,In_2241);
or U1580 (N_1580,N_368,In_339);
nand U1581 (N_1581,In_1043,In_134);
or U1582 (N_1582,In_857,N_454);
xnor U1583 (N_1583,In_2713,In_2218);
nor U1584 (N_1584,N_880,N_536);
or U1585 (N_1585,In_2986,In_2407);
xor U1586 (N_1586,N_341,In_2080);
and U1587 (N_1587,In_1804,N_167);
nand U1588 (N_1588,N_826,N_804);
xor U1589 (N_1589,N_425,In_1103);
xnor U1590 (N_1590,N_379,In_514);
nand U1591 (N_1591,In_2196,N_478);
and U1592 (N_1592,N_14,N_771);
xnor U1593 (N_1593,N_590,N_242);
xnor U1594 (N_1594,N_897,N_926);
nand U1595 (N_1595,In_368,In_2163);
nand U1596 (N_1596,N_711,N_7);
and U1597 (N_1597,N_269,In_2255);
and U1598 (N_1598,In_1324,N_731);
xnor U1599 (N_1599,In_815,In_2331);
nand U1600 (N_1600,In_341,N_113);
and U1601 (N_1601,In_2400,N_617);
and U1602 (N_1602,In_2134,In_2436);
or U1603 (N_1603,In_1760,In_2535);
nor U1604 (N_1604,In_2785,In_1914);
nand U1605 (N_1605,In_1944,In_84);
or U1606 (N_1606,In_2895,In_1576);
or U1607 (N_1607,N_190,In_662);
and U1608 (N_1608,N_982,In_2002);
and U1609 (N_1609,N_312,N_192);
xnor U1610 (N_1610,N_507,N_6);
nor U1611 (N_1611,N_487,In_2877);
or U1612 (N_1612,N_642,In_2470);
nor U1613 (N_1613,N_334,N_406);
or U1614 (N_1614,In_2842,In_744);
nand U1615 (N_1615,In_5,In_2969);
xor U1616 (N_1616,N_511,In_2063);
nand U1617 (N_1617,N_612,N_427);
and U1618 (N_1618,In_2794,In_663);
nand U1619 (N_1619,In_1548,In_1952);
nor U1620 (N_1620,N_486,In_1475);
nand U1621 (N_1621,In_708,N_1);
and U1622 (N_1622,In_1384,In_1274);
or U1623 (N_1623,N_970,N_570);
or U1624 (N_1624,N_954,In_395);
nor U1625 (N_1625,In_1386,In_2382);
xor U1626 (N_1626,In_703,In_2992);
and U1627 (N_1627,In_2497,N_968);
or U1628 (N_1628,N_729,N_369);
and U1629 (N_1629,In_464,N_216);
nor U1630 (N_1630,N_68,In_438);
or U1631 (N_1631,In_2012,N_120);
nor U1632 (N_1632,In_1858,N_899);
and U1633 (N_1633,In_1599,N_537);
nor U1634 (N_1634,N_225,In_2896);
xor U1635 (N_1635,In_2222,N_17);
nand U1636 (N_1636,N_816,In_1254);
nand U1637 (N_1637,In_760,N_844);
xnor U1638 (N_1638,In_2364,N_479);
and U1639 (N_1639,N_852,In_2946);
nor U1640 (N_1640,N_927,N_277);
nor U1641 (N_1641,N_869,N_322);
nor U1642 (N_1642,N_392,In_233);
nand U1643 (N_1643,N_614,In_1217);
xnor U1644 (N_1644,In_1981,In_742);
nor U1645 (N_1645,N_420,N_297);
and U1646 (N_1646,In_1615,In_2676);
and U1647 (N_1647,N_325,N_285);
nor U1648 (N_1648,In_1959,In_54);
or U1649 (N_1649,N_101,N_571);
nor U1650 (N_1650,N_648,N_817);
xor U1651 (N_1651,In_86,N_754);
and U1652 (N_1652,In_801,In_131);
and U1653 (N_1653,In_654,N_796);
and U1654 (N_1654,N_770,In_509);
and U1655 (N_1655,In_57,N_75);
and U1656 (N_1656,In_2588,N_644);
and U1657 (N_1657,In_113,In_2357);
or U1658 (N_1658,N_635,In_1609);
and U1659 (N_1659,In_1767,In_989);
nand U1660 (N_1660,N_318,N_367);
or U1661 (N_1661,In_1192,N_310);
or U1662 (N_1662,N_898,In_321);
and U1663 (N_1663,N_302,In_2900);
or U1664 (N_1664,In_911,N_573);
nor U1665 (N_1665,N_942,In_1474);
nor U1666 (N_1666,N_870,In_144);
nand U1667 (N_1667,N_881,N_976);
nand U1668 (N_1668,N_831,N_504);
nand U1669 (N_1669,In_502,N_49);
xor U1670 (N_1670,N_463,In_415);
or U1671 (N_1671,In_1692,In_1532);
or U1672 (N_1672,In_1029,N_255);
nor U1673 (N_1673,In_2405,N_815);
or U1674 (N_1674,In_814,In_782);
and U1675 (N_1675,In_74,In_2478);
and U1676 (N_1676,In_870,N_517);
nor U1677 (N_1677,N_389,N_121);
or U1678 (N_1678,In_2890,N_967);
xor U1679 (N_1679,N_955,In_999);
and U1680 (N_1680,N_958,N_641);
or U1681 (N_1681,N_524,N_919);
nor U1682 (N_1682,In_854,In_2266);
nand U1683 (N_1683,In_716,In_1126);
nand U1684 (N_1684,N_408,N_513);
nor U1685 (N_1685,In_797,In_37);
nor U1686 (N_1686,N_402,In_2099);
nor U1687 (N_1687,In_886,In_2318);
or U1688 (N_1688,N_980,N_422);
nor U1689 (N_1689,N_458,N_82);
nand U1690 (N_1690,In_1741,N_205);
or U1691 (N_1691,N_647,In_1927);
and U1692 (N_1692,In_2201,In_2190);
xnor U1693 (N_1693,N_244,N_794);
nor U1694 (N_1694,N_8,In_2414);
or U1695 (N_1695,N_417,N_466);
and U1696 (N_1696,N_308,In_818);
or U1697 (N_1697,N_587,In_812);
xnor U1698 (N_1698,N_44,In_1010);
xnor U1699 (N_1699,In_497,In_2282);
or U1700 (N_1700,In_1698,N_39);
xor U1701 (N_1701,In_323,N_488);
nand U1702 (N_1702,In_2660,N_268);
nand U1703 (N_1703,In_376,N_247);
nand U1704 (N_1704,In_1011,In_1683);
nand U1705 (N_1705,In_433,N_136);
and U1706 (N_1706,In_852,N_293);
nor U1707 (N_1707,In_2069,N_656);
xor U1708 (N_1708,N_965,In_1246);
nor U1709 (N_1709,In_1752,N_323);
nor U1710 (N_1710,In_1616,N_551);
nor U1711 (N_1711,In_2728,N_999);
and U1712 (N_1712,N_26,N_806);
or U1713 (N_1713,In_768,N_633);
or U1714 (N_1714,N_272,In_1744);
nand U1715 (N_1715,N_382,N_291);
nor U1716 (N_1716,In_38,N_332);
nand U1717 (N_1717,N_355,N_733);
xor U1718 (N_1718,In_2914,In_2397);
nor U1719 (N_1719,N_884,N_432);
and U1720 (N_1720,In_1088,In_1);
nand U1721 (N_1721,N_944,N_563);
or U1722 (N_1722,N_765,N_384);
and U1723 (N_1723,In_1923,N_597);
and U1724 (N_1724,N_159,N_720);
nor U1725 (N_1725,N_348,N_262);
xnor U1726 (N_1726,In_489,In_1593);
or U1727 (N_1727,In_108,N_848);
xor U1728 (N_1728,In_619,In_1494);
xnor U1729 (N_1729,N_429,In_494);
and U1730 (N_1730,In_792,In_1026);
nand U1731 (N_1731,In_1312,In_2883);
nand U1732 (N_1732,In_158,In_1790);
nand U1733 (N_1733,N_543,N_615);
xor U1734 (N_1734,In_2632,In_1216);
or U1735 (N_1735,N_939,In_1666);
or U1736 (N_1736,N_636,In_2682);
nand U1737 (N_1737,In_2739,N_171);
or U1738 (N_1738,In_2203,In_751);
nor U1739 (N_1739,In_2809,N_254);
or U1740 (N_1740,In_874,In_2348);
xnor U1741 (N_1741,In_614,N_140);
and U1742 (N_1742,N_660,N_734);
xor U1743 (N_1743,N_28,In_2472);
nor U1744 (N_1744,In_2750,N_391);
nand U1745 (N_1745,In_344,N_197);
and U1746 (N_1746,N_502,In_1153);
or U1747 (N_1747,In_2341,In_222);
or U1748 (N_1748,In_2894,N_455);
nand U1749 (N_1749,In_998,In_200);
and U1750 (N_1750,N_221,N_583);
or U1751 (N_1751,In_2990,In_1865);
nor U1752 (N_1752,In_820,N_19);
or U1753 (N_1753,N_52,In_1721);
or U1754 (N_1754,N_929,N_393);
and U1755 (N_1755,In_2479,N_930);
nor U1756 (N_1756,In_2901,N_45);
xor U1757 (N_1757,In_88,In_1344);
nor U1758 (N_1758,N_69,N_495);
nand U1759 (N_1759,N_223,In_1847);
or U1760 (N_1760,N_266,In_1922);
or U1761 (N_1761,In_2965,In_1612);
nor U1762 (N_1762,N_450,N_685);
and U1763 (N_1763,N_925,N_527);
or U1764 (N_1764,N_5,In_1720);
nor U1765 (N_1765,N_441,N_683);
or U1766 (N_1766,N_233,In_160);
xor U1767 (N_1767,In_2504,In_2538);
nand U1768 (N_1768,In_1583,N_855);
nand U1769 (N_1769,N_457,In_1113);
xor U1770 (N_1770,In_269,N_834);
nor U1771 (N_1771,N_135,In_263);
and U1772 (N_1772,N_822,N_485);
xor U1773 (N_1773,In_1712,In_1726);
xor U1774 (N_1774,In_2204,N_330);
xnor U1775 (N_1775,In_2435,In_1307);
and U1776 (N_1776,N_707,N_643);
nand U1777 (N_1777,In_231,In_1530);
or U1778 (N_1778,N_662,N_678);
or U1779 (N_1779,N_329,N_618);
and U1780 (N_1780,In_1707,N_516);
nand U1781 (N_1781,In_944,N_773);
or U1782 (N_1782,In_2922,In_277);
nand U1783 (N_1783,N_271,In_308);
or U1784 (N_1784,In_2140,In_1916);
nand U1785 (N_1785,In_2951,N_36);
and U1786 (N_1786,In_2811,In_2610);
nor U1787 (N_1787,N_789,In_2018);
or U1788 (N_1788,N_838,N_91);
nor U1789 (N_1789,N_518,In_1061);
xor U1790 (N_1790,N_800,N_111);
and U1791 (N_1791,N_357,In_533);
xor U1792 (N_1792,In_2638,In_2105);
nand U1793 (N_1793,In_2763,In_519);
xnor U1794 (N_1794,In_2384,In_2568);
nor U1795 (N_1795,N_474,N_821);
nor U1796 (N_1796,N_41,N_476);
or U1797 (N_1797,N_139,N_147);
and U1798 (N_1798,In_1873,In_285);
or U1799 (N_1799,In_425,In_685);
nand U1800 (N_1800,In_2026,In_2259);
nor U1801 (N_1801,N_503,In_2980);
nand U1802 (N_1802,In_2313,In_2412);
nor U1803 (N_1803,N_442,N_227);
and U1804 (N_1804,N_864,In_412);
or U1805 (N_1805,In_1190,N_760);
xnor U1806 (N_1806,N_725,In_258);
nor U1807 (N_1807,N_842,N_240);
nor U1808 (N_1808,N_983,N_309);
xor U1809 (N_1809,N_687,In_1653);
xnor U1810 (N_1810,N_151,N_337);
nand U1811 (N_1811,N_755,N_288);
xnor U1812 (N_1812,N_71,In_2450);
nor U1813 (N_1813,N_948,In_702);
or U1814 (N_1814,N_132,N_481);
nand U1815 (N_1815,N_676,In_1231);
and U1816 (N_1816,In_2790,N_757);
nand U1817 (N_1817,In_2651,N_303);
xor U1818 (N_1818,N_316,In_29);
or U1819 (N_1819,N_514,In_2639);
nand U1820 (N_1820,N_313,In_745);
nand U1821 (N_1821,In_1303,N_859);
xor U1822 (N_1822,In_714,N_492);
nor U1823 (N_1823,In_1511,In_859);
nand U1824 (N_1824,N_286,N_181);
xor U1825 (N_1825,N_515,N_430);
nor U1826 (N_1826,N_373,In_2418);
nand U1827 (N_1827,N_709,N_751);
and U1828 (N_1828,In_109,In_1243);
nor U1829 (N_1829,N_289,N_27);
and U1830 (N_1830,In_1232,In_2496);
and U1831 (N_1831,N_605,In_897);
nand U1832 (N_1832,N_282,In_1519);
nand U1833 (N_1833,In_1590,In_959);
or U1834 (N_1834,N_871,N_172);
xor U1835 (N_1835,N_353,In_506);
nor U1836 (N_1836,N_354,In_513);
nor U1837 (N_1837,N_972,N_703);
nor U1838 (N_1838,N_632,N_638);
or U1839 (N_1839,In_2195,In_247);
and U1840 (N_1840,N_978,N_130);
or U1841 (N_1841,In_697,N_745);
and U1842 (N_1842,N_493,In_2813);
or U1843 (N_1843,N_232,N_294);
nor U1844 (N_1844,N_890,In_1628);
xor U1845 (N_1845,In_2261,In_892);
or U1846 (N_1846,N_657,N_990);
xor U1847 (N_1847,In_1211,In_1734);
and U1848 (N_1848,In_342,In_1136);
and U1849 (N_1849,In_2421,In_2193);
xor U1850 (N_1850,In_652,In_141);
or U1851 (N_1851,In_195,In_2793);
or U1852 (N_1852,N_784,In_2392);
nor U1853 (N_1853,N_252,N_798);
xnor U1854 (N_1854,N_372,In_1549);
nand U1855 (N_1855,N_673,N_324);
and U1856 (N_1856,In_1818,N_646);
nand U1857 (N_1857,N_175,N_273);
or U1858 (N_1858,In_2869,N_533);
or U1859 (N_1859,N_279,N_237);
xnor U1860 (N_1860,In_580,In_2770);
or U1861 (N_1861,In_1021,N_76);
nor U1862 (N_1862,N_718,In_1277);
or U1863 (N_1863,In_1555,N_37);
nand U1864 (N_1864,In_271,In_76);
and U1865 (N_1865,In_684,N_126);
or U1866 (N_1866,In_2878,N_311);
and U1867 (N_1867,N_70,In_2612);
or U1868 (N_1868,In_46,N_84);
nor U1869 (N_1869,In_162,N_651);
xnor U1870 (N_1870,N_696,N_79);
nor U1871 (N_1871,N_554,N_679);
nor U1872 (N_1872,N_705,N_434);
or U1873 (N_1873,In_1448,In_573);
nor U1874 (N_1874,N_464,N_889);
or U1875 (N_1875,N_946,N_611);
or U1876 (N_1876,N_104,In_252);
nor U1877 (N_1877,In_2815,N_444);
and U1878 (N_1878,In_915,In_756);
nand U1879 (N_1879,N_356,N_321);
nand U1880 (N_1880,N_744,In_2184);
nor U1881 (N_1881,In_2695,N_480);
and U1882 (N_1882,In_1130,N_398);
xor U1883 (N_1883,In_465,In_2067);
xnor U1884 (N_1884,N_62,N_108);
nand U1885 (N_1885,N_446,In_1335);
or U1886 (N_1886,N_214,N_645);
and U1887 (N_1887,N_452,In_1297);
and U1888 (N_1888,N_793,N_412);
xor U1889 (N_1889,In_2416,In_696);
and U1890 (N_1890,N_989,N_995);
xnor U1891 (N_1891,In_1779,N_522);
nor U1892 (N_1892,N_654,N_892);
xor U1893 (N_1893,In_1306,N_604);
nand U1894 (N_1894,In_16,N_856);
and U1895 (N_1895,In_1362,N_115);
nor U1896 (N_1896,N_945,N_65);
nor U1897 (N_1897,In_1732,In_2958);
nor U1898 (N_1898,N_907,N_397);
or U1899 (N_1899,N_92,N_224);
and U1900 (N_1900,N_365,In_1554);
nor U1901 (N_1901,N_498,N_680);
nand U1902 (N_1902,N_250,In_2457);
nand U1903 (N_1903,N_320,N_867);
and U1904 (N_1904,N_129,N_483);
and U1905 (N_1905,In_463,In_713);
nor U1906 (N_1906,N_260,N_11);
nand U1907 (N_1907,In_501,In_1281);
and U1908 (N_1908,In_2955,N_16);
nand U1909 (N_1909,In_931,In_194);
nor U1910 (N_1910,In_372,N_281);
nor U1911 (N_1911,In_1839,N_73);
nand U1912 (N_1912,In_2246,In_2294);
nor U1913 (N_1913,N_423,N_903);
nor U1914 (N_1914,N_421,In_1841);
nand U1915 (N_1915,In_1926,In_2148);
and U1916 (N_1916,In_1640,In_1534);
nand U1917 (N_1917,In_647,N_292);
nor U1918 (N_1918,In_552,In_248);
xnor U1919 (N_1919,N_579,N_774);
or U1920 (N_1920,N_388,In_2426);
and U1921 (N_1921,N_428,N_116);
and U1922 (N_1922,N_758,In_2383);
and U1923 (N_1923,N_910,N_90);
nor U1924 (N_1924,In_2370,In_69);
xnor U1925 (N_1925,N_258,N_512);
xnor U1926 (N_1926,In_694,In_93);
nor U1927 (N_1927,In_2332,In_155);
nor U1928 (N_1928,In_2406,N_666);
nor U1929 (N_1929,In_95,N_520);
nand U1930 (N_1930,N_400,N_807);
nor U1931 (N_1931,N_872,In_1605);
and U1932 (N_1932,In_2843,In_648);
or U1933 (N_1933,N_296,N_390);
nor U1934 (N_1934,In_1282,N_860);
xor U1935 (N_1935,In_2153,N_562);
and U1936 (N_1936,In_971,In_2428);
or U1937 (N_1937,N_788,In_1123);
nand U1938 (N_1938,In_606,N_46);
nor U1939 (N_1939,In_371,In_587);
xnor U1940 (N_1940,N_177,N_732);
xor U1941 (N_1941,In_1622,In_831);
nor U1942 (N_1942,N_163,In_1114);
nand U1943 (N_1943,N_419,N_761);
xnor U1944 (N_1944,N_531,N_24);
and U1945 (N_1945,In_1711,In_1275);
nand U1946 (N_1946,N_865,N_544);
and U1947 (N_1947,In_462,N_123);
and U1948 (N_1948,In_2189,In_2981);
and U1949 (N_1949,N_35,N_568);
nand U1950 (N_1950,In_1716,In_1794);
nor U1951 (N_1951,N_374,In_1080);
xor U1952 (N_1952,N_366,In_2772);
or U1953 (N_1953,N_813,N_528);
nor U1954 (N_1954,N_433,In_1750);
nand U1955 (N_1955,In_451,In_2430);
nand U1956 (N_1956,In_2761,N_183);
nand U1957 (N_1957,In_2904,N_336);
xor U1958 (N_1958,In_1863,N_9);
or U1959 (N_1959,In_1526,In_1785);
nor U1960 (N_1960,In_2742,N_370);
nor U1961 (N_1961,N_383,N_490);
or U1962 (N_1962,N_395,N_589);
and U1963 (N_1963,N_836,In_2704);
nor U1964 (N_1964,In_1239,N_780);
and U1965 (N_1965,N_920,N_596);
and U1966 (N_1966,N_12,N_819);
nand U1967 (N_1967,N_736,In_1052);
nor U1968 (N_1968,In_763,N_178);
and U1969 (N_1969,N_346,In_317);
nand U1970 (N_1970,In_1350,N_333);
or U1971 (N_1971,N_717,N_81);
xnor U1972 (N_1972,In_2882,N_530);
nand U1973 (N_1973,N_465,In_829);
or U1974 (N_1974,N_922,In_63);
nor U1975 (N_1975,N_386,In_89);
xor U1976 (N_1976,In_2066,In_898);
and U1977 (N_1977,In_2253,N_344);
nor U1978 (N_1978,N_783,N_338);
xor U1979 (N_1979,N_300,In_495);
nor U1980 (N_1980,In_968,In_1433);
nor U1981 (N_1981,In_461,In_1382);
and U1982 (N_1982,N_936,N_72);
xor U1983 (N_1983,N_290,In_2028);
xnor U1984 (N_1984,In_53,In_1869);
nor U1985 (N_1985,In_225,In_650);
or U1986 (N_1986,In_2257,N_63);
nand U1987 (N_1987,N_701,In_2081);
nand U1988 (N_1988,In_1179,In_1950);
or U1989 (N_1989,In_264,N_173);
or U1990 (N_1990,In_816,In_2143);
nand U1991 (N_1991,N_677,In_472);
or U1992 (N_1992,N_759,In_1078);
and U1993 (N_1993,In_1257,N_144);
or U1994 (N_1994,N_665,N_307);
or U1995 (N_1995,In_1792,In_2867);
and U1996 (N_1996,N_138,N_20);
nand U1997 (N_1997,N_888,In_1652);
nand U1998 (N_1998,In_656,N_961);
nand U1999 (N_1999,N_359,In_2592);
or U2000 (N_2000,N_1646,N_1797);
nor U2001 (N_2001,N_1953,N_1166);
nor U2002 (N_2002,N_1380,N_1134);
xor U2003 (N_2003,N_1067,N_1463);
nand U2004 (N_2004,N_1679,N_1939);
xnor U2005 (N_2005,N_1061,N_1268);
and U2006 (N_2006,N_1219,N_1818);
xor U2007 (N_2007,N_1577,N_1556);
or U2008 (N_2008,N_1882,N_1719);
xor U2009 (N_2009,N_1014,N_1831);
nor U2010 (N_2010,N_1040,N_1596);
or U2011 (N_2011,N_1736,N_1641);
nor U2012 (N_2012,N_1922,N_1343);
or U2013 (N_2013,N_1782,N_1001);
or U2014 (N_2014,N_1251,N_1649);
nor U2015 (N_2015,N_1206,N_1483);
or U2016 (N_2016,N_1100,N_1430);
and U2017 (N_2017,N_1481,N_1650);
nand U2018 (N_2018,N_1868,N_1064);
nand U2019 (N_2019,N_1033,N_1357);
nand U2020 (N_2020,N_1562,N_1169);
and U2021 (N_2021,N_1408,N_1377);
or U2022 (N_2022,N_1290,N_1202);
and U2023 (N_2023,N_1824,N_1150);
or U2024 (N_2024,N_1954,N_1437);
nand U2025 (N_2025,N_1688,N_1045);
and U2026 (N_2026,N_1926,N_1386);
nor U2027 (N_2027,N_1029,N_1837);
xnor U2028 (N_2028,N_1574,N_1945);
or U2029 (N_2029,N_1088,N_1956);
nand U2030 (N_2030,N_1648,N_1960);
nor U2031 (N_2031,N_1404,N_1355);
nor U2032 (N_2032,N_1994,N_1976);
and U2033 (N_2033,N_1398,N_1457);
xnor U2034 (N_2034,N_1581,N_1199);
nand U2035 (N_2035,N_1286,N_1222);
nand U2036 (N_2036,N_1758,N_1419);
nand U2037 (N_2037,N_1167,N_1966);
and U2038 (N_2038,N_1018,N_1030);
nor U2039 (N_2039,N_1579,N_1242);
nand U2040 (N_2040,N_1750,N_1850);
xnor U2041 (N_2041,N_1348,N_1936);
nor U2042 (N_2042,N_1247,N_1342);
nor U2043 (N_2043,N_1157,N_1684);
xor U2044 (N_2044,N_1791,N_1937);
xnor U2045 (N_2045,N_1560,N_1883);
and U2046 (N_2046,N_1591,N_1110);
nand U2047 (N_2047,N_1112,N_1142);
nand U2048 (N_2048,N_1527,N_1474);
nor U2049 (N_2049,N_1393,N_1547);
and U2050 (N_2050,N_1390,N_1164);
xnor U2051 (N_2051,N_1839,N_1707);
and U2052 (N_2052,N_1830,N_1848);
or U2053 (N_2053,N_1148,N_1967);
or U2054 (N_2054,N_1987,N_1710);
or U2055 (N_2055,N_1432,N_1345);
nand U2056 (N_2056,N_1344,N_1520);
and U2057 (N_2057,N_1042,N_1827);
and U2058 (N_2058,N_1754,N_1210);
nand U2059 (N_2059,N_1168,N_1723);
xnor U2060 (N_2060,N_1454,N_1031);
and U2061 (N_2061,N_1270,N_1125);
and U2062 (N_2062,N_1655,N_1821);
and U2063 (N_2063,N_1993,N_1312);
or U2064 (N_2064,N_1834,N_1863);
and U2065 (N_2065,N_1808,N_1948);
or U2066 (N_2066,N_1693,N_1915);
and U2067 (N_2067,N_1517,N_1084);
xnor U2068 (N_2068,N_1026,N_1442);
nand U2069 (N_2069,N_1443,N_1949);
and U2070 (N_2070,N_1196,N_1198);
xnor U2071 (N_2071,N_1768,N_1041);
or U2072 (N_2072,N_1846,N_1606);
xnor U2073 (N_2073,N_1983,N_1347);
and U2074 (N_2074,N_1047,N_1385);
and U2075 (N_2075,N_1958,N_1910);
nor U2076 (N_2076,N_1739,N_1070);
xnor U2077 (N_2077,N_1594,N_1424);
xor U2078 (N_2078,N_1970,N_1476);
and U2079 (N_2079,N_1217,N_1304);
nand U2080 (N_2080,N_1654,N_1094);
nand U2081 (N_2081,N_1322,N_1158);
nor U2082 (N_2082,N_1721,N_1779);
nand U2083 (N_2083,N_1711,N_1301);
or U2084 (N_2084,N_1121,N_1551);
nor U2085 (N_2085,N_1644,N_1115);
nor U2086 (N_2086,N_1749,N_1531);
and U2087 (N_2087,N_1906,N_1192);
nand U2088 (N_2088,N_1942,N_1440);
or U2089 (N_2089,N_1610,N_1506);
and U2090 (N_2090,N_1459,N_1996);
or U2091 (N_2091,N_1384,N_1809);
xnor U2092 (N_2092,N_1287,N_1081);
and U2093 (N_2093,N_1914,N_1456);
xnor U2094 (N_2094,N_1555,N_1232);
or U2095 (N_2095,N_1665,N_1066);
xor U2096 (N_2096,N_1248,N_1093);
nand U2097 (N_2097,N_1672,N_1132);
and U2098 (N_2098,N_1427,N_1608);
and U2099 (N_2099,N_1775,N_1753);
and U2100 (N_2100,N_1661,N_1737);
and U2101 (N_2101,N_1174,N_1571);
and U2102 (N_2102,N_1896,N_1969);
nor U2103 (N_2103,N_1681,N_1674);
or U2104 (N_2104,N_1544,N_1752);
nand U2105 (N_2105,N_1341,N_1726);
nor U2106 (N_2106,N_1801,N_1616);
nand U2107 (N_2107,N_1120,N_1193);
nor U2108 (N_2108,N_1776,N_1911);
xor U2109 (N_2109,N_1812,N_1642);
nor U2110 (N_2110,N_1010,N_1173);
or U2111 (N_2111,N_1558,N_1549);
nor U2112 (N_2112,N_1756,N_1659);
and U2113 (N_2113,N_1091,N_1647);
and U2114 (N_2114,N_1059,N_1441);
xor U2115 (N_2115,N_1292,N_1773);
or U2116 (N_2116,N_1853,N_1034);
and U2117 (N_2117,N_1515,N_1260);
and U2118 (N_2118,N_1358,N_1645);
xor U2119 (N_2119,N_1930,N_1493);
xor U2120 (N_2120,N_1327,N_1306);
and U2121 (N_2121,N_1036,N_1777);
nor U2122 (N_2122,N_1485,N_1625);
and U2123 (N_2123,N_1262,N_1369);
and U2124 (N_2124,N_1058,N_1622);
and U2125 (N_2125,N_1620,N_1643);
nand U2126 (N_2126,N_1467,N_1184);
xor U2127 (N_2127,N_1267,N_1657);
nand U2128 (N_2128,N_1634,N_1855);
and U2129 (N_2129,N_1353,N_1871);
nor U2130 (N_2130,N_1767,N_1607);
nand U2131 (N_2131,N_1052,N_1630);
xnor U2132 (N_2132,N_1139,N_1367);
or U2133 (N_2133,N_1941,N_1195);
xnor U2134 (N_2134,N_1313,N_1946);
and U2135 (N_2135,N_1772,N_1144);
nand U2136 (N_2136,N_1155,N_1235);
or U2137 (N_2137,N_1806,N_1351);
nor U2138 (N_2138,N_1107,N_1748);
and U2139 (N_2139,N_1455,N_1567);
or U2140 (N_2140,N_1046,N_1228);
nor U2141 (N_2141,N_1538,N_1734);
and U2142 (N_2142,N_1704,N_1225);
nor U2143 (N_2143,N_1407,N_1133);
and U2144 (N_2144,N_1460,N_1552);
or U2145 (N_2145,N_1305,N_1986);
nor U2146 (N_2146,N_1981,N_1920);
nor U2147 (N_2147,N_1618,N_1955);
or U2148 (N_2148,N_1103,N_1480);
nand U2149 (N_2149,N_1931,N_1141);
nand U2150 (N_2150,N_1448,N_1951);
nand U2151 (N_2151,N_1479,N_1609);
and U2152 (N_2152,N_1213,N_1578);
nor U2153 (N_2153,N_1019,N_1470);
nor U2154 (N_2154,N_1800,N_1436);
nor U2155 (N_2155,N_1504,N_1502);
xnor U2156 (N_2156,N_1867,N_1671);
nand U2157 (N_2157,N_1988,N_1000);
nor U2158 (N_2158,N_1200,N_1147);
xor U2159 (N_2159,N_1374,N_1289);
nor U2160 (N_2160,N_1513,N_1016);
or U2161 (N_2161,N_1114,N_1127);
nor U2162 (N_2162,N_1316,N_1098);
nand U2163 (N_2163,N_1396,N_1604);
xnor U2164 (N_2164,N_1537,N_1395);
or U2165 (N_2165,N_1523,N_1256);
nand U2166 (N_2166,N_1843,N_1412);
and U2167 (N_2167,N_1445,N_1275);
and U2168 (N_2168,N_1415,N_1866);
nand U2169 (N_2169,N_1165,N_1239);
and U2170 (N_2170,N_1838,N_1337);
xor U2171 (N_2171,N_1478,N_1011);
xnor U2172 (N_2172,N_1947,N_1022);
and U2173 (N_2173,N_1592,N_1580);
nor U2174 (N_2174,N_1680,N_1979);
xnor U2175 (N_2175,N_1980,N_1216);
or U2176 (N_2176,N_1439,N_1220);
xnor U2177 (N_2177,N_1279,N_1743);
and U2178 (N_2178,N_1472,N_1897);
or U2179 (N_2179,N_1600,N_1813);
xor U2180 (N_2180,N_1745,N_1170);
nor U2181 (N_2181,N_1308,N_1261);
nor U2182 (N_2182,N_1140,N_1546);
nand U2183 (N_2183,N_1392,N_1338);
nand U2184 (N_2184,N_1762,N_1633);
nor U2185 (N_2185,N_1152,N_1177);
xor U2186 (N_2186,N_1835,N_1788);
nor U2187 (N_2187,N_1231,N_1944);
nand U2188 (N_2188,N_1530,N_1488);
and U2189 (N_2189,N_1899,N_1324);
or U2190 (N_2190,N_1397,N_1105);
nand U2191 (N_2191,N_1695,N_1639);
nor U2192 (N_2192,N_1664,N_1588);
nor U2193 (N_2193,N_1807,N_1602);
nand U2194 (N_2194,N_1413,N_1400);
nor U2195 (N_2195,N_1746,N_1590);
nor U2196 (N_2196,N_1917,N_1083);
nand U2197 (N_2197,N_1720,N_1733);
nand U2198 (N_2198,N_1027,N_1792);
nor U2199 (N_2199,N_1656,N_1466);
or U2200 (N_2200,N_1833,N_1038);
xor U2201 (N_2201,N_1852,N_1712);
nand U2202 (N_2202,N_1653,N_1469);
xor U2203 (N_2203,N_1875,N_1893);
and U2204 (N_2204,N_1522,N_1934);
and U2205 (N_2205,N_1929,N_1113);
xor U2206 (N_2206,N_1569,N_1051);
and U2207 (N_2207,N_1526,N_1740);
or U2208 (N_2208,N_1399,N_1820);
xnor U2209 (N_2209,N_1370,N_1375);
and U2210 (N_2210,N_1770,N_1182);
nand U2211 (N_2211,N_1468,N_1130);
nand U2212 (N_2212,N_1814,N_1971);
xnor U2213 (N_2213,N_1111,N_1742);
and U2214 (N_2214,N_1236,N_1933);
xor U2215 (N_2215,N_1887,N_1787);
and U2216 (N_2216,N_1728,N_1190);
or U2217 (N_2217,N_1007,N_1371);
nor U2218 (N_2218,N_1116,N_1593);
xnor U2219 (N_2219,N_1346,N_1096);
and U2220 (N_2220,N_1984,N_1889);
nor U2221 (N_2221,N_1487,N_1361);
or U2222 (N_2222,N_1092,N_1543);
and U2223 (N_2223,N_1884,N_1730);
and U2224 (N_2224,N_1296,N_1539);
and U2225 (N_2225,N_1662,N_1802);
xor U2226 (N_2226,N_1964,N_1696);
xnor U2227 (N_2227,N_1450,N_1410);
xnor U2228 (N_2228,N_1008,N_1329);
and U2229 (N_2229,N_1626,N_1461);
nand U2230 (N_2230,N_1209,N_1145);
nor U2231 (N_2231,N_1160,N_1918);
and U2232 (N_2232,N_1420,N_1619);
and U2233 (N_2233,N_1597,N_1589);
nor U2234 (N_2234,N_1708,N_1912);
or U2235 (N_2235,N_1854,N_1281);
nor U2236 (N_2236,N_1585,N_1938);
nand U2237 (N_2237,N_1595,N_1499);
xor U2238 (N_2238,N_1055,N_1423);
nand U2239 (N_2239,N_1885,N_1426);
and U2240 (N_2240,N_1069,N_1940);
nor U2241 (N_2241,N_1117,N_1627);
xnor U2242 (N_2242,N_1796,N_1378);
or U2243 (N_2243,N_1605,N_1126);
or U2244 (N_2244,N_1446,N_1999);
and U2245 (N_2245,N_1240,N_1844);
xnor U2246 (N_2246,N_1965,N_1482);
or U2247 (N_2247,N_1161,N_1372);
and U2248 (N_2248,N_1628,N_1054);
xor U2249 (N_2249,N_1265,N_1335);
nor U2250 (N_2250,N_1901,N_1729);
or U2251 (N_2251,N_1181,N_1360);
or U2252 (N_2252,N_1858,N_1873);
and U2253 (N_2253,N_1722,N_1637);
nor U2254 (N_2254,N_1223,N_1277);
nor U2255 (N_2255,N_1611,N_1149);
nor U2256 (N_2256,N_1387,N_1391);
or U2257 (N_2257,N_1414,N_1266);
xor U2258 (N_2258,N_1354,N_1204);
xor U2259 (N_2259,N_1293,N_1409);
or U2260 (N_2260,N_1851,N_1795);
and U2261 (N_2261,N_1118,N_1179);
nor U2262 (N_2262,N_1285,N_1128);
nand U2263 (N_2263,N_1559,N_1421);
nand U2264 (N_2264,N_1194,N_1841);
nand U2265 (N_2265,N_1307,N_1550);
nand U2266 (N_2266,N_1352,N_1484);
nand U2267 (N_2267,N_1326,N_1362);
nand U2268 (N_2268,N_1238,N_1904);
nor U2269 (N_2269,N_1651,N_1254);
nor U2270 (N_2270,N_1715,N_1632);
nand U2271 (N_2271,N_1186,N_1143);
nand U2272 (N_2272,N_1032,N_1491);
nand U2273 (N_2273,N_1163,N_1511);
nor U2274 (N_2274,N_1603,N_1845);
xor U2275 (N_2275,N_1631,N_1124);
xnor U2276 (N_2276,N_1294,N_1935);
nand U2277 (N_2277,N_1815,N_1138);
xor U2278 (N_2278,N_1280,N_1025);
xor U2279 (N_2279,N_1438,N_1245);
xnor U2280 (N_2280,N_1548,N_1519);
or U2281 (N_2281,N_1810,N_1009);
nor U2282 (N_2282,N_1895,N_1135);
nor U2283 (N_2283,N_1747,N_1013);
and U2284 (N_2284,N_1699,N_1477);
or U2285 (N_2285,N_1525,N_1176);
xnor U2286 (N_2286,N_1146,N_1529);
or U2287 (N_2287,N_1892,N_1330);
or U2288 (N_2288,N_1044,N_1295);
xor U2289 (N_2289,N_1876,N_1489);
nand U2290 (N_2290,N_1565,N_1601);
and U2291 (N_2291,N_1826,N_1274);
nand U2292 (N_2292,N_1237,N_1908);
and U2293 (N_2293,N_1003,N_1458);
nand U2294 (N_2294,N_1402,N_1617);
or U2295 (N_2295,N_1624,N_1921);
nor U2296 (N_2296,N_1973,N_1255);
nand U2297 (N_2297,N_1874,N_1498);
nor U2298 (N_2298,N_1823,N_1898);
nor U2299 (N_2299,N_1670,N_1886);
or U2300 (N_2300,N_1043,N_1687);
and U2301 (N_2301,N_1211,N_1180);
and U2302 (N_2302,N_1162,N_1663);
nor U2303 (N_2303,N_1784,N_1203);
nand U2304 (N_2304,N_1183,N_1284);
nand U2305 (N_2305,N_1989,N_1060);
or U2306 (N_2306,N_1677,N_1794);
xnor U2307 (N_2307,N_1218,N_1510);
nor U2308 (N_2308,N_1789,N_1303);
xnor U2309 (N_2309,N_1761,N_1024);
or U2310 (N_2310,N_1447,N_1686);
or U2311 (N_2311,N_1576,N_1471);
nor U2312 (N_2312,N_1288,N_1257);
nor U2313 (N_2313,N_1464,N_1119);
and U2314 (N_2314,N_1388,N_1435);
xor U2315 (N_2315,N_1366,N_1961);
nand U2316 (N_2316,N_1405,N_1071);
nor U2317 (N_2317,N_1943,N_1249);
or U2318 (N_2318,N_1963,N_1101);
xnor U2319 (N_2319,N_1089,N_1350);
xor U2320 (N_2320,N_1518,N_1108);
nor U2321 (N_2321,N_1978,N_1535);
nor U2322 (N_2322,N_1990,N_1977);
nor U2323 (N_2323,N_1263,N_1512);
nor U2324 (N_2324,N_1842,N_1997);
xnor U2325 (N_2325,N_1859,N_1205);
nand U2326 (N_2326,N_1568,N_1339);
nor U2327 (N_2327,N_1077,N_1252);
xnor U2328 (N_2328,N_1185,N_1349);
xor U2329 (N_2329,N_1129,N_1959);
xor U2330 (N_2330,N_1233,N_1403);
or U2331 (N_2331,N_1545,N_1658);
or U2332 (N_2332,N_1613,N_1497);
xnor U2333 (N_2333,N_1612,N_1271);
nand U2334 (N_2334,N_1283,N_1928);
or U2335 (N_2335,N_1226,N_1159);
nor U2336 (N_2336,N_1713,N_1297);
or U2337 (N_2337,N_1678,N_1706);
xor U2338 (N_2338,N_1475,N_1724);
or U2339 (N_2339,N_1401,N_1153);
or U2340 (N_2340,N_1137,N_1102);
and U2341 (N_2341,N_1431,N_1072);
nand U2342 (N_2342,N_1425,N_1765);
and U2343 (N_2343,N_1718,N_1541);
nand U2344 (N_2344,N_1907,N_1865);
nand U2345 (N_2345,N_1381,N_1697);
xnor U2346 (N_2346,N_1763,N_1599);
and U2347 (N_2347,N_1328,N_1073);
nand U2348 (N_2348,N_1923,N_1816);
nor U2349 (N_2349,N_1334,N_1406);
nor U2350 (N_2350,N_1501,N_1175);
nor U2351 (N_2351,N_1080,N_1382);
nor U2352 (N_2352,N_1079,N_1278);
and U2353 (N_2353,N_1785,N_1258);
nor U2354 (N_2354,N_1516,N_1566);
xnor U2355 (N_2355,N_1311,N_1264);
and U2356 (N_2356,N_1982,N_1669);
nand U2357 (N_2357,N_1197,N_1187);
nand U2358 (N_2358,N_1916,N_1751);
or U2359 (N_2359,N_1774,N_1760);
and U2360 (N_2360,N_1972,N_1836);
and U2361 (N_2361,N_1171,N_1974);
nor U2362 (N_2362,N_1764,N_1573);
nor U2363 (N_2363,N_1952,N_1891);
and U2364 (N_2364,N_1790,N_1056);
nor U2365 (N_2365,N_1319,N_1241);
nand U2366 (N_2366,N_1793,N_1786);
or U2367 (N_2367,N_1356,N_1919);
and U2368 (N_2368,N_1564,N_1074);
nand U2369 (N_2369,N_1856,N_1048);
nor U2370 (N_2370,N_1321,N_1065);
nand U2371 (N_2371,N_1717,N_1021);
nand U2372 (N_2372,N_1227,N_1698);
and U2373 (N_2373,N_1212,N_1700);
or U2374 (N_2374,N_1514,N_1207);
and U2375 (N_2375,N_1099,N_1985);
nor U2376 (N_2376,N_1189,N_1068);
and U2377 (N_2377,N_1359,N_1243);
xnor U2378 (N_2378,N_1444,N_1417);
or U2379 (N_2379,N_1085,N_1178);
xor U2380 (N_2380,N_1039,N_1496);
or U2381 (N_2381,N_1214,N_1318);
and U2382 (N_2382,N_1509,N_1861);
and U2383 (N_2383,N_1095,N_1554);
nand U2384 (N_2384,N_1500,N_1870);
nor U2385 (N_2385,N_1379,N_1716);
xor U2386 (N_2386,N_1667,N_1104);
or U2387 (N_2387,N_1635,N_1462);
xnor U2388 (N_2388,N_1368,N_1583);
nand U2389 (N_2389,N_1582,N_1172);
nand U2390 (N_2390,N_1273,N_1224);
and U2391 (N_2391,N_1890,N_1683);
or U2392 (N_2392,N_1614,N_1453);
and U2393 (N_2393,N_1309,N_1629);
nand U2394 (N_2394,N_1057,N_1002);
and U2395 (N_2395,N_1738,N_1727);
nand U2396 (N_2396,N_1615,N_1598);
xnor U2397 (N_2397,N_1798,N_1894);
nand U2398 (N_2398,N_1492,N_1825);
and U2399 (N_2399,N_1817,N_1584);
xnor U2400 (N_2400,N_1062,N_1741);
xor U2401 (N_2401,N_1735,N_1004);
xnor U2402 (N_2402,N_1422,N_1528);
and U2403 (N_2403,N_1314,N_1636);
or U2404 (N_2404,N_1320,N_1905);
xnor U2405 (N_2405,N_1106,N_1803);
nand U2406 (N_2406,N_1878,N_1832);
or U2407 (N_2407,N_1006,N_1725);
nand U2408 (N_2408,N_1151,N_1269);
and U2409 (N_2409,N_1924,N_1012);
nand U2410 (N_2410,N_1900,N_1299);
and U2411 (N_2411,N_1536,N_1097);
and U2412 (N_2412,N_1995,N_1418);
nor U2413 (N_2413,N_1714,N_1557);
and U2414 (N_2414,N_1811,N_1563);
nor U2415 (N_2415,N_1962,N_1847);
nor U2416 (N_2416,N_1364,N_1154);
nor U2417 (N_2417,N_1005,N_1780);
and U2418 (N_2418,N_1215,N_1822);
and U2419 (N_2419,N_1575,N_1122);
and U2420 (N_2420,N_1053,N_1587);
nor U2421 (N_2421,N_1201,N_1524);
xor U2422 (N_2422,N_1690,N_1666);
and U2423 (N_2423,N_1676,N_1769);
nand U2424 (N_2424,N_1298,N_1668);
or U2425 (N_2425,N_1340,N_1333);
or U2426 (N_2426,N_1136,N_1692);
xnor U2427 (N_2427,N_1473,N_1682);
nand U2428 (N_2428,N_1416,N_1234);
and U2429 (N_2429,N_1428,N_1660);
nor U2430 (N_2430,N_1759,N_1703);
and U2431 (N_2431,N_1376,N_1086);
xnor U2432 (N_2432,N_1829,N_1521);
and U2433 (N_2433,N_1037,N_1494);
nor U2434 (N_2434,N_1805,N_1804);
nor U2435 (N_2435,N_1394,N_1230);
nand U2436 (N_2436,N_1879,N_1015);
and U2437 (N_2437,N_1975,N_1433);
nand U2438 (N_2438,N_1250,N_1927);
xnor U2439 (N_2439,N_1389,N_1035);
or U2440 (N_2440,N_1302,N_1495);
xor U2441 (N_2441,N_1877,N_1049);
nor U2442 (N_2442,N_1486,N_1490);
nand U2443 (N_2443,N_1272,N_1766);
nor U2444 (N_2444,N_1325,N_1429);
nand U2445 (N_2445,N_1363,N_1623);
and U2446 (N_2446,N_1849,N_1840);
or U2447 (N_2447,N_1701,N_1869);
xnor U2448 (N_2448,N_1050,N_1323);
and U2449 (N_2449,N_1731,N_1451);
and U2450 (N_2450,N_1276,N_1411);
xnor U2451 (N_2451,N_1465,N_1702);
nor U2452 (N_2452,N_1259,N_1336);
xnor U2453 (N_2453,N_1572,N_1503);
nand U2454 (N_2454,N_1075,N_1783);
nor U2455 (N_2455,N_1913,N_1188);
and U2456 (N_2456,N_1123,N_1208);
nor U2457 (N_2457,N_1638,N_1534);
or U2458 (N_2458,N_1689,N_1023);
and U2459 (N_2459,N_1621,N_1076);
nor U2460 (N_2460,N_1998,N_1449);
or U2461 (N_2461,N_1909,N_1586);
xnor U2462 (N_2462,N_1991,N_1156);
xnor U2463 (N_2463,N_1640,N_1332);
xnor U2464 (N_2464,N_1968,N_1755);
nor U2465 (N_2465,N_1872,N_1992);
and U2466 (N_2466,N_1819,N_1191);
nor U2467 (N_2467,N_1561,N_1315);
and U2468 (N_2468,N_1020,N_1881);
nand U2469 (N_2469,N_1957,N_1902);
and U2470 (N_2470,N_1950,N_1282);
xnor U2471 (N_2471,N_1652,N_1570);
nand U2472 (N_2472,N_1063,N_1507);
nand U2473 (N_2473,N_1880,N_1828);
and U2474 (N_2474,N_1310,N_1781);
nor U2475 (N_2475,N_1778,N_1860);
nor U2476 (N_2476,N_1028,N_1540);
xor U2477 (N_2477,N_1244,N_1542);
or U2478 (N_2478,N_1373,N_1331);
nor U2479 (N_2479,N_1673,N_1757);
nand U2480 (N_2480,N_1434,N_1862);
nand U2481 (N_2481,N_1675,N_1685);
and U2482 (N_2482,N_1082,N_1300);
nand U2483 (N_2483,N_1799,N_1109);
nand U2484 (N_2484,N_1365,N_1888);
or U2485 (N_2485,N_1291,N_1864);
nor U2486 (N_2486,N_1508,N_1090);
and U2487 (N_2487,N_1903,N_1744);
or U2488 (N_2488,N_1532,N_1246);
nor U2489 (N_2489,N_1131,N_1694);
or U2490 (N_2490,N_1553,N_1533);
nor U2491 (N_2491,N_1709,N_1317);
nor U2492 (N_2492,N_1017,N_1925);
and U2493 (N_2493,N_1078,N_1229);
or U2494 (N_2494,N_1771,N_1705);
xor U2495 (N_2495,N_1857,N_1383);
nor U2496 (N_2496,N_1221,N_1253);
xnor U2497 (N_2497,N_1732,N_1505);
nor U2498 (N_2498,N_1452,N_1932);
xnor U2499 (N_2499,N_1691,N_1087);
and U2500 (N_2500,N_1625,N_1552);
or U2501 (N_2501,N_1861,N_1002);
nand U2502 (N_2502,N_1485,N_1240);
nor U2503 (N_2503,N_1534,N_1165);
or U2504 (N_2504,N_1409,N_1673);
nand U2505 (N_2505,N_1631,N_1333);
nor U2506 (N_2506,N_1310,N_1101);
nor U2507 (N_2507,N_1386,N_1896);
xnor U2508 (N_2508,N_1704,N_1057);
or U2509 (N_2509,N_1468,N_1548);
or U2510 (N_2510,N_1019,N_1910);
nor U2511 (N_2511,N_1500,N_1545);
or U2512 (N_2512,N_1829,N_1197);
xnor U2513 (N_2513,N_1354,N_1922);
xnor U2514 (N_2514,N_1197,N_1711);
or U2515 (N_2515,N_1862,N_1601);
xor U2516 (N_2516,N_1163,N_1013);
nand U2517 (N_2517,N_1155,N_1003);
and U2518 (N_2518,N_1226,N_1476);
or U2519 (N_2519,N_1869,N_1226);
and U2520 (N_2520,N_1260,N_1952);
nand U2521 (N_2521,N_1721,N_1812);
or U2522 (N_2522,N_1370,N_1593);
nand U2523 (N_2523,N_1811,N_1355);
nand U2524 (N_2524,N_1639,N_1119);
nand U2525 (N_2525,N_1830,N_1127);
and U2526 (N_2526,N_1397,N_1328);
xor U2527 (N_2527,N_1508,N_1990);
or U2528 (N_2528,N_1219,N_1075);
xnor U2529 (N_2529,N_1022,N_1253);
or U2530 (N_2530,N_1620,N_1793);
nand U2531 (N_2531,N_1124,N_1608);
or U2532 (N_2532,N_1020,N_1981);
nor U2533 (N_2533,N_1258,N_1791);
and U2534 (N_2534,N_1282,N_1450);
or U2535 (N_2535,N_1570,N_1811);
or U2536 (N_2536,N_1251,N_1499);
nor U2537 (N_2537,N_1438,N_1689);
or U2538 (N_2538,N_1142,N_1428);
nand U2539 (N_2539,N_1659,N_1118);
and U2540 (N_2540,N_1275,N_1929);
or U2541 (N_2541,N_1706,N_1814);
nand U2542 (N_2542,N_1931,N_1875);
or U2543 (N_2543,N_1458,N_1587);
nand U2544 (N_2544,N_1154,N_1623);
and U2545 (N_2545,N_1624,N_1745);
xnor U2546 (N_2546,N_1581,N_1457);
xnor U2547 (N_2547,N_1316,N_1874);
and U2548 (N_2548,N_1510,N_1662);
or U2549 (N_2549,N_1423,N_1062);
and U2550 (N_2550,N_1457,N_1887);
and U2551 (N_2551,N_1935,N_1636);
and U2552 (N_2552,N_1810,N_1611);
xnor U2553 (N_2553,N_1429,N_1129);
nand U2554 (N_2554,N_1699,N_1221);
or U2555 (N_2555,N_1396,N_1150);
nand U2556 (N_2556,N_1229,N_1606);
nor U2557 (N_2557,N_1346,N_1133);
nor U2558 (N_2558,N_1329,N_1555);
nor U2559 (N_2559,N_1018,N_1986);
and U2560 (N_2560,N_1141,N_1797);
or U2561 (N_2561,N_1646,N_1864);
xor U2562 (N_2562,N_1680,N_1632);
nor U2563 (N_2563,N_1120,N_1924);
xor U2564 (N_2564,N_1733,N_1381);
nor U2565 (N_2565,N_1551,N_1126);
xor U2566 (N_2566,N_1186,N_1051);
nor U2567 (N_2567,N_1168,N_1245);
nand U2568 (N_2568,N_1561,N_1593);
nand U2569 (N_2569,N_1425,N_1867);
or U2570 (N_2570,N_1259,N_1828);
xnor U2571 (N_2571,N_1189,N_1492);
or U2572 (N_2572,N_1288,N_1208);
nor U2573 (N_2573,N_1746,N_1655);
xor U2574 (N_2574,N_1590,N_1233);
nand U2575 (N_2575,N_1313,N_1914);
nor U2576 (N_2576,N_1135,N_1700);
or U2577 (N_2577,N_1651,N_1695);
and U2578 (N_2578,N_1941,N_1853);
nand U2579 (N_2579,N_1082,N_1208);
nand U2580 (N_2580,N_1138,N_1299);
or U2581 (N_2581,N_1469,N_1490);
xor U2582 (N_2582,N_1399,N_1283);
xnor U2583 (N_2583,N_1340,N_1846);
or U2584 (N_2584,N_1181,N_1576);
and U2585 (N_2585,N_1212,N_1935);
and U2586 (N_2586,N_1294,N_1162);
nand U2587 (N_2587,N_1294,N_1654);
or U2588 (N_2588,N_1805,N_1627);
xnor U2589 (N_2589,N_1598,N_1377);
and U2590 (N_2590,N_1271,N_1190);
nand U2591 (N_2591,N_1784,N_1958);
or U2592 (N_2592,N_1024,N_1728);
xor U2593 (N_2593,N_1162,N_1419);
nor U2594 (N_2594,N_1986,N_1926);
xnor U2595 (N_2595,N_1861,N_1314);
nor U2596 (N_2596,N_1157,N_1369);
xor U2597 (N_2597,N_1513,N_1818);
nand U2598 (N_2598,N_1899,N_1491);
and U2599 (N_2599,N_1183,N_1706);
xor U2600 (N_2600,N_1715,N_1166);
nor U2601 (N_2601,N_1482,N_1880);
or U2602 (N_2602,N_1965,N_1549);
xor U2603 (N_2603,N_1714,N_1420);
or U2604 (N_2604,N_1117,N_1178);
xor U2605 (N_2605,N_1616,N_1749);
nor U2606 (N_2606,N_1004,N_1161);
and U2607 (N_2607,N_1746,N_1663);
or U2608 (N_2608,N_1609,N_1177);
nor U2609 (N_2609,N_1111,N_1114);
or U2610 (N_2610,N_1044,N_1173);
nor U2611 (N_2611,N_1786,N_1855);
nand U2612 (N_2612,N_1421,N_1473);
and U2613 (N_2613,N_1418,N_1797);
nand U2614 (N_2614,N_1846,N_1560);
xor U2615 (N_2615,N_1003,N_1372);
nand U2616 (N_2616,N_1591,N_1543);
or U2617 (N_2617,N_1602,N_1315);
nor U2618 (N_2618,N_1734,N_1645);
and U2619 (N_2619,N_1597,N_1476);
nor U2620 (N_2620,N_1434,N_1566);
nor U2621 (N_2621,N_1900,N_1625);
nor U2622 (N_2622,N_1139,N_1483);
nor U2623 (N_2623,N_1068,N_1792);
nand U2624 (N_2624,N_1500,N_1941);
and U2625 (N_2625,N_1782,N_1407);
nor U2626 (N_2626,N_1125,N_1557);
and U2627 (N_2627,N_1778,N_1429);
and U2628 (N_2628,N_1676,N_1277);
nand U2629 (N_2629,N_1487,N_1024);
nor U2630 (N_2630,N_1036,N_1941);
nand U2631 (N_2631,N_1525,N_1597);
and U2632 (N_2632,N_1252,N_1525);
nand U2633 (N_2633,N_1009,N_1065);
xor U2634 (N_2634,N_1046,N_1239);
and U2635 (N_2635,N_1495,N_1991);
nor U2636 (N_2636,N_1552,N_1453);
or U2637 (N_2637,N_1825,N_1462);
nor U2638 (N_2638,N_1177,N_1817);
nor U2639 (N_2639,N_1843,N_1031);
or U2640 (N_2640,N_1461,N_1391);
xnor U2641 (N_2641,N_1533,N_1380);
or U2642 (N_2642,N_1014,N_1753);
nor U2643 (N_2643,N_1559,N_1534);
xor U2644 (N_2644,N_1793,N_1385);
xor U2645 (N_2645,N_1318,N_1930);
or U2646 (N_2646,N_1489,N_1412);
nand U2647 (N_2647,N_1647,N_1496);
and U2648 (N_2648,N_1888,N_1046);
nand U2649 (N_2649,N_1948,N_1819);
xnor U2650 (N_2650,N_1665,N_1814);
nand U2651 (N_2651,N_1574,N_1308);
or U2652 (N_2652,N_1074,N_1283);
nand U2653 (N_2653,N_1397,N_1901);
or U2654 (N_2654,N_1925,N_1313);
or U2655 (N_2655,N_1505,N_1758);
and U2656 (N_2656,N_1988,N_1474);
xor U2657 (N_2657,N_1087,N_1970);
nand U2658 (N_2658,N_1724,N_1263);
and U2659 (N_2659,N_1096,N_1608);
xor U2660 (N_2660,N_1150,N_1400);
nand U2661 (N_2661,N_1935,N_1359);
nand U2662 (N_2662,N_1811,N_1476);
nor U2663 (N_2663,N_1469,N_1399);
and U2664 (N_2664,N_1814,N_1653);
xor U2665 (N_2665,N_1101,N_1341);
nor U2666 (N_2666,N_1756,N_1644);
or U2667 (N_2667,N_1783,N_1789);
and U2668 (N_2668,N_1378,N_1747);
or U2669 (N_2669,N_1882,N_1262);
xnor U2670 (N_2670,N_1052,N_1274);
nor U2671 (N_2671,N_1156,N_1708);
nor U2672 (N_2672,N_1560,N_1212);
or U2673 (N_2673,N_1613,N_1263);
nor U2674 (N_2674,N_1640,N_1743);
nand U2675 (N_2675,N_1045,N_1973);
xor U2676 (N_2676,N_1374,N_1251);
and U2677 (N_2677,N_1906,N_1344);
or U2678 (N_2678,N_1439,N_1035);
nor U2679 (N_2679,N_1519,N_1847);
or U2680 (N_2680,N_1119,N_1185);
or U2681 (N_2681,N_1327,N_1325);
nor U2682 (N_2682,N_1931,N_1582);
or U2683 (N_2683,N_1800,N_1983);
or U2684 (N_2684,N_1182,N_1518);
and U2685 (N_2685,N_1650,N_1396);
xor U2686 (N_2686,N_1290,N_1580);
and U2687 (N_2687,N_1176,N_1479);
xnor U2688 (N_2688,N_1182,N_1425);
or U2689 (N_2689,N_1495,N_1227);
xor U2690 (N_2690,N_1386,N_1133);
nand U2691 (N_2691,N_1656,N_1237);
or U2692 (N_2692,N_1090,N_1997);
xor U2693 (N_2693,N_1661,N_1994);
or U2694 (N_2694,N_1559,N_1217);
xor U2695 (N_2695,N_1523,N_1817);
nor U2696 (N_2696,N_1311,N_1562);
xor U2697 (N_2697,N_1369,N_1068);
nand U2698 (N_2698,N_1981,N_1299);
nand U2699 (N_2699,N_1421,N_1357);
nand U2700 (N_2700,N_1336,N_1328);
or U2701 (N_2701,N_1670,N_1198);
xnor U2702 (N_2702,N_1504,N_1594);
and U2703 (N_2703,N_1669,N_1367);
nand U2704 (N_2704,N_1997,N_1178);
nand U2705 (N_2705,N_1794,N_1342);
nand U2706 (N_2706,N_1862,N_1365);
xor U2707 (N_2707,N_1027,N_1240);
and U2708 (N_2708,N_1037,N_1263);
and U2709 (N_2709,N_1286,N_1968);
nand U2710 (N_2710,N_1328,N_1079);
nor U2711 (N_2711,N_1976,N_1231);
nor U2712 (N_2712,N_1368,N_1934);
or U2713 (N_2713,N_1465,N_1920);
nand U2714 (N_2714,N_1392,N_1293);
or U2715 (N_2715,N_1906,N_1846);
and U2716 (N_2716,N_1056,N_1709);
xnor U2717 (N_2717,N_1604,N_1940);
xnor U2718 (N_2718,N_1286,N_1719);
xor U2719 (N_2719,N_1221,N_1362);
nor U2720 (N_2720,N_1002,N_1015);
xnor U2721 (N_2721,N_1133,N_1382);
nor U2722 (N_2722,N_1897,N_1602);
nand U2723 (N_2723,N_1419,N_1158);
or U2724 (N_2724,N_1607,N_1460);
nor U2725 (N_2725,N_1246,N_1738);
nor U2726 (N_2726,N_1202,N_1122);
xnor U2727 (N_2727,N_1196,N_1164);
xor U2728 (N_2728,N_1003,N_1506);
nand U2729 (N_2729,N_1769,N_1235);
or U2730 (N_2730,N_1603,N_1944);
nand U2731 (N_2731,N_1102,N_1380);
or U2732 (N_2732,N_1314,N_1480);
nand U2733 (N_2733,N_1002,N_1698);
xnor U2734 (N_2734,N_1930,N_1938);
or U2735 (N_2735,N_1656,N_1086);
xor U2736 (N_2736,N_1562,N_1656);
nand U2737 (N_2737,N_1257,N_1088);
xnor U2738 (N_2738,N_1786,N_1842);
nor U2739 (N_2739,N_1037,N_1314);
or U2740 (N_2740,N_1609,N_1406);
and U2741 (N_2741,N_1174,N_1737);
and U2742 (N_2742,N_1370,N_1136);
nand U2743 (N_2743,N_1253,N_1166);
nand U2744 (N_2744,N_1688,N_1825);
nor U2745 (N_2745,N_1233,N_1944);
nor U2746 (N_2746,N_1535,N_1322);
or U2747 (N_2747,N_1210,N_1341);
and U2748 (N_2748,N_1975,N_1072);
nor U2749 (N_2749,N_1884,N_1630);
nand U2750 (N_2750,N_1915,N_1559);
or U2751 (N_2751,N_1001,N_1701);
nor U2752 (N_2752,N_1622,N_1347);
nand U2753 (N_2753,N_1228,N_1150);
and U2754 (N_2754,N_1449,N_1802);
xnor U2755 (N_2755,N_1066,N_1183);
nand U2756 (N_2756,N_1117,N_1294);
or U2757 (N_2757,N_1276,N_1371);
nor U2758 (N_2758,N_1291,N_1703);
nand U2759 (N_2759,N_1202,N_1707);
or U2760 (N_2760,N_1781,N_1801);
nor U2761 (N_2761,N_1833,N_1672);
nand U2762 (N_2762,N_1836,N_1469);
nand U2763 (N_2763,N_1601,N_1557);
or U2764 (N_2764,N_1361,N_1023);
nand U2765 (N_2765,N_1154,N_1547);
and U2766 (N_2766,N_1528,N_1082);
or U2767 (N_2767,N_1560,N_1042);
xnor U2768 (N_2768,N_1782,N_1812);
nor U2769 (N_2769,N_1897,N_1550);
nand U2770 (N_2770,N_1292,N_1215);
xor U2771 (N_2771,N_1855,N_1850);
xor U2772 (N_2772,N_1636,N_1416);
and U2773 (N_2773,N_1016,N_1394);
nand U2774 (N_2774,N_1583,N_1967);
or U2775 (N_2775,N_1608,N_1492);
nor U2776 (N_2776,N_1930,N_1492);
xor U2777 (N_2777,N_1714,N_1906);
nor U2778 (N_2778,N_1476,N_1900);
xor U2779 (N_2779,N_1591,N_1776);
nor U2780 (N_2780,N_1807,N_1585);
or U2781 (N_2781,N_1586,N_1741);
nand U2782 (N_2782,N_1248,N_1592);
nand U2783 (N_2783,N_1757,N_1690);
nand U2784 (N_2784,N_1001,N_1462);
xnor U2785 (N_2785,N_1409,N_1950);
or U2786 (N_2786,N_1084,N_1357);
and U2787 (N_2787,N_1965,N_1270);
nor U2788 (N_2788,N_1083,N_1878);
or U2789 (N_2789,N_1328,N_1706);
and U2790 (N_2790,N_1113,N_1766);
nor U2791 (N_2791,N_1284,N_1929);
and U2792 (N_2792,N_1322,N_1285);
xnor U2793 (N_2793,N_1983,N_1909);
nor U2794 (N_2794,N_1346,N_1220);
or U2795 (N_2795,N_1694,N_1079);
nand U2796 (N_2796,N_1083,N_1615);
xnor U2797 (N_2797,N_1203,N_1806);
or U2798 (N_2798,N_1618,N_1380);
or U2799 (N_2799,N_1459,N_1082);
nand U2800 (N_2800,N_1022,N_1625);
and U2801 (N_2801,N_1874,N_1674);
and U2802 (N_2802,N_1921,N_1329);
or U2803 (N_2803,N_1409,N_1424);
and U2804 (N_2804,N_1395,N_1965);
nor U2805 (N_2805,N_1081,N_1368);
or U2806 (N_2806,N_1773,N_1783);
nor U2807 (N_2807,N_1887,N_1753);
or U2808 (N_2808,N_1889,N_1756);
nor U2809 (N_2809,N_1759,N_1230);
xor U2810 (N_2810,N_1571,N_1878);
nand U2811 (N_2811,N_1230,N_1073);
or U2812 (N_2812,N_1730,N_1370);
and U2813 (N_2813,N_1284,N_1674);
or U2814 (N_2814,N_1007,N_1820);
and U2815 (N_2815,N_1477,N_1051);
nor U2816 (N_2816,N_1893,N_1319);
or U2817 (N_2817,N_1430,N_1282);
nor U2818 (N_2818,N_1582,N_1081);
and U2819 (N_2819,N_1600,N_1566);
or U2820 (N_2820,N_1519,N_1887);
nand U2821 (N_2821,N_1980,N_1559);
or U2822 (N_2822,N_1907,N_1331);
or U2823 (N_2823,N_1649,N_1695);
and U2824 (N_2824,N_1200,N_1654);
xnor U2825 (N_2825,N_1962,N_1971);
or U2826 (N_2826,N_1274,N_1201);
nor U2827 (N_2827,N_1944,N_1882);
nor U2828 (N_2828,N_1304,N_1547);
and U2829 (N_2829,N_1344,N_1915);
and U2830 (N_2830,N_1592,N_1112);
nand U2831 (N_2831,N_1925,N_1139);
nand U2832 (N_2832,N_1813,N_1072);
or U2833 (N_2833,N_1849,N_1664);
nor U2834 (N_2834,N_1802,N_1683);
nand U2835 (N_2835,N_1689,N_1887);
or U2836 (N_2836,N_1523,N_1127);
nand U2837 (N_2837,N_1270,N_1960);
nor U2838 (N_2838,N_1887,N_1972);
nor U2839 (N_2839,N_1441,N_1585);
xor U2840 (N_2840,N_1298,N_1506);
and U2841 (N_2841,N_1553,N_1869);
and U2842 (N_2842,N_1331,N_1887);
nand U2843 (N_2843,N_1022,N_1603);
xnor U2844 (N_2844,N_1011,N_1475);
xnor U2845 (N_2845,N_1543,N_1526);
and U2846 (N_2846,N_1235,N_1821);
and U2847 (N_2847,N_1922,N_1624);
or U2848 (N_2848,N_1327,N_1534);
nand U2849 (N_2849,N_1626,N_1112);
nand U2850 (N_2850,N_1756,N_1634);
nand U2851 (N_2851,N_1594,N_1588);
or U2852 (N_2852,N_1282,N_1523);
xnor U2853 (N_2853,N_1195,N_1101);
nor U2854 (N_2854,N_1079,N_1413);
or U2855 (N_2855,N_1016,N_1635);
nand U2856 (N_2856,N_1417,N_1850);
nor U2857 (N_2857,N_1978,N_1014);
nand U2858 (N_2858,N_1094,N_1081);
nand U2859 (N_2859,N_1506,N_1402);
or U2860 (N_2860,N_1569,N_1477);
or U2861 (N_2861,N_1283,N_1467);
and U2862 (N_2862,N_1989,N_1541);
and U2863 (N_2863,N_1848,N_1750);
or U2864 (N_2864,N_1067,N_1005);
nand U2865 (N_2865,N_1992,N_1423);
or U2866 (N_2866,N_1801,N_1937);
nand U2867 (N_2867,N_1510,N_1142);
and U2868 (N_2868,N_1224,N_1876);
nand U2869 (N_2869,N_1739,N_1006);
or U2870 (N_2870,N_1946,N_1580);
or U2871 (N_2871,N_1450,N_1499);
or U2872 (N_2872,N_1869,N_1033);
and U2873 (N_2873,N_1045,N_1214);
and U2874 (N_2874,N_1208,N_1230);
nand U2875 (N_2875,N_1469,N_1956);
or U2876 (N_2876,N_1511,N_1117);
and U2877 (N_2877,N_1402,N_1828);
nand U2878 (N_2878,N_1077,N_1056);
xnor U2879 (N_2879,N_1961,N_1438);
xnor U2880 (N_2880,N_1005,N_1482);
xor U2881 (N_2881,N_1351,N_1501);
and U2882 (N_2882,N_1766,N_1561);
xor U2883 (N_2883,N_1879,N_1489);
and U2884 (N_2884,N_1214,N_1546);
nor U2885 (N_2885,N_1010,N_1480);
xnor U2886 (N_2886,N_1953,N_1548);
or U2887 (N_2887,N_1018,N_1553);
or U2888 (N_2888,N_1788,N_1084);
nor U2889 (N_2889,N_1307,N_1390);
xor U2890 (N_2890,N_1429,N_1229);
or U2891 (N_2891,N_1331,N_1308);
nor U2892 (N_2892,N_1782,N_1940);
nor U2893 (N_2893,N_1019,N_1100);
nand U2894 (N_2894,N_1722,N_1365);
nor U2895 (N_2895,N_1601,N_1284);
nand U2896 (N_2896,N_1836,N_1732);
nand U2897 (N_2897,N_1146,N_1125);
nand U2898 (N_2898,N_1758,N_1088);
nand U2899 (N_2899,N_1686,N_1790);
or U2900 (N_2900,N_1706,N_1398);
and U2901 (N_2901,N_1221,N_1516);
and U2902 (N_2902,N_1622,N_1559);
nand U2903 (N_2903,N_1321,N_1402);
nand U2904 (N_2904,N_1679,N_1764);
or U2905 (N_2905,N_1649,N_1283);
nand U2906 (N_2906,N_1780,N_1412);
and U2907 (N_2907,N_1393,N_1900);
or U2908 (N_2908,N_1998,N_1432);
nor U2909 (N_2909,N_1301,N_1417);
or U2910 (N_2910,N_1890,N_1481);
and U2911 (N_2911,N_1549,N_1399);
or U2912 (N_2912,N_1125,N_1407);
nor U2913 (N_2913,N_1591,N_1743);
or U2914 (N_2914,N_1877,N_1153);
nand U2915 (N_2915,N_1794,N_1335);
and U2916 (N_2916,N_1688,N_1387);
and U2917 (N_2917,N_1515,N_1961);
xnor U2918 (N_2918,N_1259,N_1983);
or U2919 (N_2919,N_1085,N_1720);
and U2920 (N_2920,N_1139,N_1653);
nand U2921 (N_2921,N_1547,N_1301);
nand U2922 (N_2922,N_1425,N_1490);
nand U2923 (N_2923,N_1249,N_1138);
xor U2924 (N_2924,N_1569,N_1260);
or U2925 (N_2925,N_1498,N_1935);
and U2926 (N_2926,N_1502,N_1445);
nor U2927 (N_2927,N_1004,N_1736);
nor U2928 (N_2928,N_1552,N_1452);
xor U2929 (N_2929,N_1273,N_1413);
xor U2930 (N_2930,N_1359,N_1020);
nor U2931 (N_2931,N_1934,N_1806);
and U2932 (N_2932,N_1333,N_1858);
nor U2933 (N_2933,N_1877,N_1657);
xor U2934 (N_2934,N_1885,N_1477);
xnor U2935 (N_2935,N_1743,N_1956);
xor U2936 (N_2936,N_1976,N_1549);
or U2937 (N_2937,N_1094,N_1949);
xnor U2938 (N_2938,N_1007,N_1589);
nor U2939 (N_2939,N_1057,N_1578);
and U2940 (N_2940,N_1070,N_1010);
and U2941 (N_2941,N_1889,N_1498);
nand U2942 (N_2942,N_1105,N_1884);
and U2943 (N_2943,N_1176,N_1335);
nand U2944 (N_2944,N_1556,N_1569);
xnor U2945 (N_2945,N_1574,N_1102);
xor U2946 (N_2946,N_1926,N_1916);
or U2947 (N_2947,N_1702,N_1028);
or U2948 (N_2948,N_1314,N_1540);
and U2949 (N_2949,N_1166,N_1945);
and U2950 (N_2950,N_1933,N_1137);
or U2951 (N_2951,N_1747,N_1472);
nor U2952 (N_2952,N_1931,N_1773);
and U2953 (N_2953,N_1978,N_1517);
xor U2954 (N_2954,N_1027,N_1552);
or U2955 (N_2955,N_1691,N_1417);
or U2956 (N_2956,N_1844,N_1575);
nor U2957 (N_2957,N_1087,N_1295);
nand U2958 (N_2958,N_1109,N_1023);
nor U2959 (N_2959,N_1441,N_1606);
and U2960 (N_2960,N_1015,N_1818);
nor U2961 (N_2961,N_1241,N_1801);
xor U2962 (N_2962,N_1520,N_1632);
and U2963 (N_2963,N_1523,N_1552);
and U2964 (N_2964,N_1985,N_1861);
or U2965 (N_2965,N_1301,N_1717);
or U2966 (N_2966,N_1028,N_1363);
and U2967 (N_2967,N_1960,N_1507);
or U2968 (N_2968,N_1575,N_1916);
and U2969 (N_2969,N_1978,N_1338);
nand U2970 (N_2970,N_1655,N_1443);
nand U2971 (N_2971,N_1841,N_1226);
or U2972 (N_2972,N_1397,N_1622);
and U2973 (N_2973,N_1620,N_1476);
or U2974 (N_2974,N_1373,N_1196);
xor U2975 (N_2975,N_1945,N_1416);
or U2976 (N_2976,N_1654,N_1481);
nand U2977 (N_2977,N_1557,N_1242);
or U2978 (N_2978,N_1874,N_1863);
xnor U2979 (N_2979,N_1384,N_1737);
nand U2980 (N_2980,N_1618,N_1978);
nor U2981 (N_2981,N_1505,N_1801);
nor U2982 (N_2982,N_1938,N_1362);
nand U2983 (N_2983,N_1463,N_1886);
and U2984 (N_2984,N_1792,N_1519);
nand U2985 (N_2985,N_1619,N_1587);
and U2986 (N_2986,N_1702,N_1314);
or U2987 (N_2987,N_1375,N_1900);
nand U2988 (N_2988,N_1023,N_1954);
xnor U2989 (N_2989,N_1938,N_1947);
and U2990 (N_2990,N_1594,N_1547);
nor U2991 (N_2991,N_1247,N_1023);
or U2992 (N_2992,N_1929,N_1736);
or U2993 (N_2993,N_1392,N_1543);
nor U2994 (N_2994,N_1346,N_1867);
xor U2995 (N_2995,N_1791,N_1732);
or U2996 (N_2996,N_1036,N_1603);
nor U2997 (N_2997,N_1986,N_1971);
nand U2998 (N_2998,N_1418,N_1153);
and U2999 (N_2999,N_1995,N_1177);
nor U3000 (N_3000,N_2500,N_2557);
or U3001 (N_3001,N_2106,N_2674);
xor U3002 (N_3002,N_2747,N_2108);
and U3003 (N_3003,N_2635,N_2559);
nor U3004 (N_3004,N_2488,N_2280);
nand U3005 (N_3005,N_2840,N_2105);
nor U3006 (N_3006,N_2489,N_2494);
or U3007 (N_3007,N_2117,N_2383);
and U3008 (N_3008,N_2192,N_2510);
nor U3009 (N_3009,N_2846,N_2671);
nor U3010 (N_3010,N_2087,N_2495);
nand U3011 (N_3011,N_2947,N_2235);
and U3012 (N_3012,N_2449,N_2194);
xor U3013 (N_3013,N_2516,N_2853);
or U3014 (N_3014,N_2109,N_2216);
nor U3015 (N_3015,N_2252,N_2163);
xor U3016 (N_3016,N_2518,N_2411);
nor U3017 (N_3017,N_2612,N_2342);
or U3018 (N_3018,N_2689,N_2148);
or U3019 (N_3019,N_2377,N_2440);
xnor U3020 (N_3020,N_2995,N_2521);
or U3021 (N_3021,N_2776,N_2804);
xnor U3022 (N_3022,N_2960,N_2887);
or U3023 (N_3023,N_2309,N_2834);
nand U3024 (N_3024,N_2811,N_2872);
or U3025 (N_3025,N_2768,N_2295);
and U3026 (N_3026,N_2427,N_2463);
nand U3027 (N_3027,N_2785,N_2751);
and U3028 (N_3028,N_2882,N_2487);
nand U3029 (N_3029,N_2934,N_2800);
nor U3030 (N_3030,N_2076,N_2878);
and U3031 (N_3031,N_2993,N_2199);
and U3032 (N_3032,N_2291,N_2017);
xnor U3033 (N_3033,N_2909,N_2704);
xnor U3034 (N_3034,N_2088,N_2599);
xnor U3035 (N_3035,N_2444,N_2234);
xnor U3036 (N_3036,N_2118,N_2517);
nand U3037 (N_3037,N_2658,N_2842);
nand U3038 (N_3038,N_2877,N_2945);
and U3039 (N_3039,N_2164,N_2292);
xor U3040 (N_3040,N_2641,N_2374);
nor U3041 (N_3041,N_2240,N_2573);
xnor U3042 (N_3042,N_2176,N_2784);
or U3043 (N_3043,N_2997,N_2208);
xor U3044 (N_3044,N_2661,N_2034);
nand U3045 (N_3045,N_2367,N_2155);
and U3046 (N_3046,N_2926,N_2056);
nor U3047 (N_3047,N_2525,N_2803);
or U3048 (N_3048,N_2224,N_2839);
nor U3049 (N_3049,N_2459,N_2986);
xor U3050 (N_3050,N_2347,N_2262);
or U3051 (N_3051,N_2639,N_2448);
or U3052 (N_3052,N_2278,N_2649);
nand U3053 (N_3053,N_2685,N_2301);
or U3054 (N_3054,N_2959,N_2548);
and U3055 (N_3055,N_2503,N_2043);
or U3056 (N_3056,N_2426,N_2369);
or U3057 (N_3057,N_2093,N_2596);
nand U3058 (N_3058,N_2771,N_2675);
and U3059 (N_3059,N_2754,N_2037);
or U3060 (N_3060,N_2364,N_2820);
nand U3061 (N_3061,N_2471,N_2786);
nor U3062 (N_3062,N_2697,N_2227);
nor U3063 (N_3063,N_2334,N_2482);
xnor U3064 (N_3064,N_2919,N_2901);
xor U3065 (N_3065,N_2568,N_2466);
or U3066 (N_3066,N_2578,N_2066);
and U3067 (N_3067,N_2756,N_2617);
or U3068 (N_3068,N_2157,N_2423);
nor U3069 (N_3069,N_2244,N_2654);
xnor U3070 (N_3070,N_2018,N_2543);
or U3071 (N_3071,N_2373,N_2779);
or U3072 (N_3072,N_2223,N_2167);
or U3073 (N_3073,N_2418,N_2188);
and U3074 (N_3074,N_2329,N_2506);
xnor U3075 (N_3075,N_2847,N_2467);
and U3076 (N_3076,N_2614,N_2065);
nor U3077 (N_3077,N_2363,N_2089);
nand U3078 (N_3078,N_2207,N_2529);
and U3079 (N_3079,N_2538,N_2469);
nor U3080 (N_3080,N_2132,N_2563);
nand U3081 (N_3081,N_2542,N_2719);
xor U3082 (N_3082,N_2791,N_2468);
xnor U3083 (N_3083,N_2987,N_2415);
and U3084 (N_3084,N_2399,N_2832);
and U3085 (N_3085,N_2273,N_2409);
nand U3086 (N_3086,N_2583,N_2958);
xor U3087 (N_3087,N_2916,N_2628);
and U3088 (N_3088,N_2237,N_2371);
and U3089 (N_3089,N_2856,N_2990);
and U3090 (N_3090,N_2370,N_2978);
xor U3091 (N_3091,N_2836,N_2582);
nand U3092 (N_3092,N_2620,N_2414);
nand U3093 (N_3093,N_2205,N_2151);
and U3094 (N_3094,N_2597,N_2186);
nor U3095 (N_3095,N_2730,N_2047);
nand U3096 (N_3096,N_2522,N_2724);
or U3097 (N_3097,N_2007,N_2509);
and U3098 (N_3098,N_2677,N_2837);
nor U3099 (N_3099,N_2158,N_2187);
or U3100 (N_3100,N_2816,N_2338);
nor U3101 (N_3101,N_2673,N_2220);
or U3102 (N_3102,N_2330,N_2360);
or U3103 (N_3103,N_2044,N_2410);
and U3104 (N_3104,N_2052,N_2261);
and U3105 (N_3105,N_2739,N_2899);
nand U3106 (N_3106,N_2711,N_2356);
nand U3107 (N_3107,N_2792,N_2149);
xor U3108 (N_3108,N_2404,N_2527);
xnor U3109 (N_3109,N_2615,N_2598);
nor U3110 (N_3110,N_2134,N_2567);
nand U3111 (N_3111,N_2021,N_2217);
or U3112 (N_3112,N_2777,N_2143);
and U3113 (N_3113,N_2336,N_2060);
and U3114 (N_3114,N_2144,N_2300);
and U3115 (N_3115,N_2113,N_2375);
nand U3116 (N_3116,N_2452,N_2643);
and U3117 (N_3117,N_2888,N_2812);
xnor U3118 (N_3118,N_2257,N_2595);
nand U3119 (N_3119,N_2593,N_2202);
nand U3120 (N_3120,N_2064,N_2095);
xnor U3121 (N_3121,N_2605,N_2028);
nor U3122 (N_3122,N_2512,N_2880);
xnor U3123 (N_3123,N_2722,N_2868);
nor U3124 (N_3124,N_2124,N_2378);
or U3125 (N_3125,N_2077,N_2337);
nor U3126 (N_3126,N_2646,N_2446);
nor U3127 (N_3127,N_2014,N_2627);
nor U3128 (N_3128,N_2528,N_2138);
or U3129 (N_3129,N_2465,N_2491);
or U3130 (N_3130,N_2607,N_2102);
or U3131 (N_3131,N_2546,N_2700);
nor U3132 (N_3132,N_2530,N_2429);
and U3133 (N_3133,N_2384,N_2835);
nor U3134 (N_3134,N_2752,N_2706);
nor U3135 (N_3135,N_2902,N_2998);
xor U3136 (N_3136,N_2749,N_2308);
nor U3137 (N_3137,N_2903,N_2507);
xor U3138 (N_3138,N_2195,N_2474);
and U3139 (N_3139,N_2968,N_2636);
nand U3140 (N_3140,N_2744,N_2335);
xnor U3141 (N_3141,N_2428,N_2304);
and U3142 (N_3142,N_2456,N_2023);
and U3143 (N_3143,N_2279,N_2083);
nor U3144 (N_3144,N_2558,N_2497);
and U3145 (N_3145,N_2953,N_2588);
xor U3146 (N_3146,N_2432,N_2633);
xor U3147 (N_3147,N_2358,N_2473);
xnor U3148 (N_3148,N_2566,N_2112);
nor U3149 (N_3149,N_2353,N_2226);
nor U3150 (N_3150,N_2855,N_2579);
xor U3151 (N_3151,N_2398,N_2002);
nor U3152 (N_3152,N_2943,N_2807);
or U3153 (N_3153,N_2642,N_2590);
nor U3154 (N_3154,N_2139,N_2119);
xor U3155 (N_3155,N_2198,N_2669);
xor U3156 (N_3156,N_2259,N_2110);
and U3157 (N_3157,N_2003,N_2447);
and U3158 (N_3158,N_2179,N_2104);
nor U3159 (N_3159,N_2349,N_2190);
nor U3160 (N_3160,N_2561,N_2225);
or U3161 (N_3161,N_2039,N_2656);
nor U3162 (N_3162,N_2948,N_2221);
or U3163 (N_3163,N_2933,N_2787);
xor U3164 (N_3164,N_2325,N_2284);
or U3165 (N_3165,N_2725,N_2867);
and U3166 (N_3166,N_2838,N_2696);
xor U3167 (N_3167,N_2897,N_2041);
or U3168 (N_3168,N_2601,N_2746);
xnor U3169 (N_3169,N_2866,N_2232);
xnor U3170 (N_3170,N_2655,N_2092);
nor U3171 (N_3171,N_2541,N_2608);
nand U3172 (N_3172,N_2735,N_2254);
or U3173 (N_3173,N_2708,N_2434);
nand U3174 (N_3174,N_2798,N_2876);
nor U3175 (N_3175,N_2750,N_2022);
nand U3176 (N_3176,N_2204,N_2504);
and U3177 (N_3177,N_2939,N_2475);
nand U3178 (N_3178,N_2822,N_2793);
and U3179 (N_3179,N_2769,N_2736);
xor U3180 (N_3180,N_2574,N_2894);
xor U3181 (N_3181,N_2801,N_2029);
nor U3182 (N_3182,N_2775,N_2778);
nor U3183 (N_3183,N_2180,N_2293);
and U3184 (N_3184,N_2984,N_2222);
nor U3185 (N_3185,N_2681,N_2055);
or U3186 (N_3186,N_2946,N_2417);
nor U3187 (N_3187,N_2854,N_2441);
or U3188 (N_3188,N_2971,N_2025);
and U3189 (N_3189,N_2587,N_2533);
and U3190 (N_3190,N_2584,N_2571);
nor U3191 (N_3191,N_2780,N_2860);
xnor U3192 (N_3192,N_2956,N_2540);
or U3193 (N_3193,N_2988,N_2405);
nand U3194 (N_3194,N_2328,N_2738);
nor U3195 (N_3195,N_2652,N_2238);
or U3196 (N_3196,N_2630,N_2274);
and U3197 (N_3197,N_2191,N_2665);
and U3198 (N_3198,N_2992,N_2267);
xnor U3199 (N_3199,N_2720,N_2264);
and U3200 (N_3200,N_2382,N_2453);
nand U3201 (N_3201,N_2631,N_2515);
nor U3202 (N_3202,N_2702,N_2004);
and U3203 (N_3203,N_2603,N_2142);
nor U3204 (N_3204,N_2162,N_2016);
nand U3205 (N_3205,N_2146,N_2890);
nor U3206 (N_3206,N_2121,N_2551);
or U3207 (N_3207,N_2153,N_2058);
nand U3208 (N_3208,N_2431,N_2898);
nand U3209 (N_3209,N_2015,N_2318);
nand U3210 (N_3210,N_2251,N_2263);
xor U3211 (N_3211,N_2006,N_2457);
xnor U3212 (N_3212,N_2687,N_2670);
nor U3213 (N_3213,N_2594,N_2536);
nor U3214 (N_3214,N_2905,N_2009);
nor U3215 (N_3215,N_2306,N_2098);
and U3216 (N_3216,N_2442,N_2718);
or U3217 (N_3217,N_2214,N_2844);
nand U3218 (N_3218,N_2758,N_2366);
xnor U3219 (N_3219,N_2618,N_2827);
nand U3220 (N_3220,N_2281,N_2075);
nor U3221 (N_3221,N_2012,N_2591);
or U3222 (N_3222,N_2114,N_2450);
and U3223 (N_3223,N_2362,N_2403);
or U3224 (N_3224,N_2874,N_2393);
nand U3225 (N_3225,N_2526,N_2623);
nor U3226 (N_3226,N_2532,N_2795);
xor U3227 (N_3227,N_2478,N_2137);
xor U3228 (N_3228,N_2760,N_2392);
nand U3229 (N_3229,N_2765,N_2556);
nand U3230 (N_3230,N_2236,N_2717);
or U3231 (N_3231,N_2954,N_2397);
and U3232 (N_3232,N_2537,N_2813);
nand U3233 (N_3233,N_2554,N_2458);
nor U3234 (N_3234,N_2451,N_2935);
nand U3235 (N_3235,N_2365,N_2312);
nor U3236 (N_3236,N_2733,N_2774);
xnor U3237 (N_3237,N_2904,N_2298);
nand U3238 (N_3238,N_2388,N_2351);
nand U3239 (N_3239,N_2664,N_2975);
nor U3240 (N_3240,N_2057,N_2299);
or U3241 (N_3241,N_2435,N_2394);
nand U3242 (N_3242,N_2511,N_2078);
xnor U3243 (N_3243,N_2930,N_2177);
or U3244 (N_3244,N_2972,N_2637);
xnor U3245 (N_3245,N_2983,N_2454);
nor U3246 (N_3246,N_2297,N_2707);
and U3247 (N_3247,N_2498,N_2182);
nand U3248 (N_3248,N_2070,N_2455);
and U3249 (N_3249,N_2924,N_2638);
or U3250 (N_3250,N_2680,N_2061);
nor U3251 (N_3251,N_2991,N_2402);
nor U3252 (N_3252,N_2662,N_2348);
xor U3253 (N_3253,N_2891,N_2289);
nor U3254 (N_3254,N_2831,N_2433);
or U3255 (N_3255,N_2307,N_2354);
nand U3256 (N_3256,N_2485,N_2107);
xor U3257 (N_3257,N_2327,N_2809);
nor U3258 (N_3258,N_2350,N_2256);
nand U3259 (N_3259,N_2914,N_2520);
or U3260 (N_3260,N_2477,N_2539);
and U3261 (N_3261,N_2985,N_2799);
and U3262 (N_3262,N_2085,N_2100);
or U3263 (N_3263,N_2091,N_2479);
nand U3264 (N_3264,N_2843,N_2046);
nor U3265 (N_3265,N_2586,N_2303);
nor U3266 (N_3266,N_2248,N_2053);
nand U3267 (N_3267,N_2071,N_2211);
xnor U3268 (N_3268,N_2322,N_2966);
xor U3269 (N_3269,N_2782,N_2097);
xnor U3270 (N_3270,N_2357,N_2229);
xor U3271 (N_3271,N_2131,N_2931);
xor U3272 (N_3272,N_2712,N_2818);
nand U3273 (N_3273,N_2174,N_2950);
nand U3274 (N_3274,N_2239,N_2406);
xnor U3275 (N_3275,N_2438,N_2920);
or U3276 (N_3276,N_2320,N_2123);
nand U3277 (N_3277,N_2727,N_2833);
nor U3278 (N_3278,N_2713,N_2806);
or U3279 (N_3279,N_2686,N_2437);
nor U3280 (N_3280,N_2302,N_2197);
xnor U3281 (N_3281,N_2421,N_2622);
or U3282 (N_3282,N_2808,N_2464);
or U3283 (N_3283,N_2624,N_2443);
and U3284 (N_3284,N_2535,N_2710);
nor U3285 (N_3285,N_2376,N_2401);
nand U3286 (N_3286,N_2970,N_2828);
or U3287 (N_3287,N_2326,N_2709);
xor U3288 (N_3288,N_2419,N_2111);
nand U3289 (N_3289,N_2266,N_2734);
nor U3290 (N_3290,N_2941,N_2159);
nand U3291 (N_3291,N_2857,N_2609);
nor U3292 (N_3292,N_2230,N_2977);
and U3293 (N_3293,N_2928,N_2082);
xor U3294 (N_3294,N_2648,N_2989);
and U3295 (N_3295,N_2116,N_2841);
or U3296 (N_3296,N_2923,N_2570);
xor U3297 (N_3297,N_2027,N_2797);
nand U3298 (N_3298,N_2343,N_2183);
or U3299 (N_3299,N_2486,N_2575);
or U3300 (N_3300,N_2886,N_2439);
xor U3301 (N_3301,N_2171,N_2729);
nand U3302 (N_3302,N_2932,N_2560);
xnor U3303 (N_3303,N_2255,N_2690);
nand U3304 (N_3304,N_2980,N_2210);
nor U3305 (N_3305,N_2921,N_2156);
nand U3306 (N_3306,N_2967,N_2900);
and U3307 (N_3307,N_2147,N_2829);
xor U3308 (N_3308,N_2391,N_2387);
and U3309 (N_3309,N_2810,N_2850);
and U3310 (N_3310,N_2368,N_2974);
and U3311 (N_3311,N_2889,N_2416);
and U3312 (N_3312,N_2359,N_2745);
nor U3313 (N_3313,N_2436,N_2869);
xor U3314 (N_3314,N_2253,N_2981);
or U3315 (N_3315,N_2870,N_2695);
or U3316 (N_3316,N_2271,N_2871);
nor U3317 (N_3317,N_2250,N_2008);
xnor U3318 (N_3318,N_2385,N_2764);
xnor U3319 (N_3319,N_2625,N_2699);
xnor U3320 (N_3320,N_2576,N_2128);
nand U3321 (N_3321,N_2361,N_2678);
and U3322 (N_3322,N_2740,N_2592);
xor U3323 (N_3323,N_2346,N_2896);
xnor U3324 (N_3324,N_2413,N_2400);
xor U3325 (N_3325,N_2125,N_2490);
xnor U3326 (N_3326,N_2269,N_2691);
or U3327 (N_3327,N_2963,N_2026);
xnor U3328 (N_3328,N_2305,N_2040);
xor U3329 (N_3329,N_2203,N_2781);
nand U3330 (N_3330,N_2245,N_2682);
xor U3331 (N_3331,N_2613,N_2938);
xor U3332 (N_3332,N_2277,N_2863);
nand U3333 (N_3333,N_2296,N_2676);
xnor U3334 (N_3334,N_2688,N_2175);
nor U3335 (N_3335,N_2859,N_2629);
nor U3336 (N_3336,N_2258,N_2714);
xnor U3337 (N_3337,N_2493,N_2247);
and U3338 (N_3338,N_2381,N_2731);
and U3339 (N_3339,N_2483,N_2496);
xnor U3340 (N_3340,N_2219,N_2524);
or U3341 (N_3341,N_2552,N_2600);
and U3342 (N_3342,N_2311,N_2602);
nand U3343 (N_3343,N_2010,N_2054);
and U3344 (N_3344,N_2042,N_2462);
xor U3345 (N_3345,N_2915,N_2858);
nand U3346 (N_3346,N_2032,N_2160);
nand U3347 (N_3347,N_2130,N_2036);
nand U3348 (N_3348,N_2165,N_2942);
nand U3349 (N_3349,N_2141,N_2033);
xor U3350 (N_3350,N_2895,N_2090);
and U3351 (N_3351,N_2789,N_2819);
nand U3352 (N_3352,N_2755,N_2790);
or U3353 (N_3353,N_2201,N_2339);
or U3354 (N_3354,N_2861,N_2951);
or U3355 (N_3355,N_2616,N_2825);
nand U3356 (N_3356,N_2660,N_2513);
and U3357 (N_3357,N_2461,N_2233);
and U3358 (N_3358,N_2703,N_2723);
xor U3359 (N_3359,N_2310,N_2879);
or U3360 (N_3360,N_2213,N_2737);
xnor U3361 (N_3361,N_2341,N_2683);
or U3362 (N_3362,N_2422,N_2480);
xnor U3363 (N_3363,N_2964,N_2120);
xor U3364 (N_3364,N_2632,N_2352);
nor U3365 (N_3365,N_2184,N_2865);
and U3366 (N_3366,N_2881,N_2189);
or U3367 (N_3367,N_2285,N_2742);
or U3368 (N_3368,N_2514,N_2973);
nand U3369 (N_3369,N_2161,N_2672);
or U3370 (N_3370,N_2577,N_2231);
nand U3371 (N_3371,N_2830,N_2355);
xor U3372 (N_3372,N_2802,N_2955);
nand U3373 (N_3373,N_2906,N_2484);
nand U3374 (N_3374,N_2024,N_2767);
nand U3375 (N_3375,N_2168,N_2936);
xnor U3376 (N_3376,N_2408,N_2531);
nor U3377 (N_3377,N_2817,N_2129);
and U3378 (N_3378,N_2845,N_2716);
xor U3379 (N_3379,N_2606,N_2965);
xor U3380 (N_3380,N_2196,N_2640);
nand U3381 (N_3381,N_2395,N_2585);
nor U3382 (N_3382,N_2260,N_2659);
or U3383 (N_3383,N_2380,N_2604);
nor U3384 (N_3384,N_2796,N_2086);
and U3385 (N_3385,N_2994,N_2663);
xnor U3386 (N_3386,N_2794,N_2961);
and U3387 (N_3387,N_2173,N_2753);
xor U3388 (N_3388,N_2815,N_2912);
nand U3389 (N_3389,N_2067,N_2396);
or U3390 (N_3390,N_2059,N_2332);
and U3391 (N_3391,N_2610,N_2884);
nor U3392 (N_3392,N_2270,N_2547);
nand U3393 (N_3393,N_2505,N_2290);
nor U3394 (N_3394,N_2424,N_2748);
or U3395 (N_3395,N_2826,N_2372);
or U3396 (N_3396,N_2081,N_2757);
and U3397 (N_3397,N_2979,N_2181);
nand U3398 (N_3398,N_2481,N_2323);
nand U3399 (N_3399,N_2243,N_2386);
or U3400 (N_3400,N_2650,N_2063);
xnor U3401 (N_3401,N_2313,N_2073);
and U3402 (N_3402,N_2331,N_2805);
xnor U3403 (N_3403,N_2875,N_2611);
nor U3404 (N_3404,N_2265,N_2910);
xor U3405 (N_3405,N_2565,N_2344);
or U3406 (N_3406,N_2645,N_2314);
or U3407 (N_3407,N_2684,N_2929);
or U3408 (N_3408,N_2922,N_2030);
or U3409 (N_3409,N_2883,N_2101);
or U3410 (N_3410,N_2653,N_2761);
xnor U3411 (N_3411,N_2553,N_2925);
or U3412 (N_3412,N_2549,N_2048);
or U3413 (N_3413,N_2940,N_2701);
and U3414 (N_3414,N_2694,N_2545);
nor U3415 (N_3415,N_2045,N_2492);
and U3416 (N_3416,N_2476,N_2268);
nor U3417 (N_3417,N_2907,N_2705);
or U3418 (N_3418,N_2550,N_2084);
or U3419 (N_3419,N_2679,N_2407);
xor U3420 (N_3420,N_2893,N_2619);
nand U3421 (N_3421,N_2848,N_2501);
xnor U3422 (N_3422,N_2976,N_2913);
nor U3423 (N_3423,N_2644,N_2741);
xnor U3424 (N_3424,N_2319,N_2873);
xnor U3425 (N_3425,N_2294,N_2049);
xor U3426 (N_3426,N_2242,N_2762);
and U3427 (N_3427,N_2732,N_2031);
xnor U3428 (N_3428,N_2657,N_2996);
and U3429 (N_3429,N_2178,N_2944);
nor U3430 (N_3430,N_2287,N_2715);
xor U3431 (N_3431,N_2094,N_2050);
nand U3432 (N_3432,N_2564,N_2759);
and U3433 (N_3433,N_2145,N_2763);
nand U3434 (N_3434,N_2911,N_2079);
nand U3435 (N_3435,N_2519,N_2862);
or U3436 (N_3436,N_2952,N_2555);
nand U3437 (N_3437,N_2103,N_2918);
or U3438 (N_3438,N_2206,N_2283);
nand U3439 (N_3439,N_2115,N_2122);
and U3440 (N_3440,N_2698,N_2788);
nand U3441 (N_3441,N_2389,N_2212);
nand U3442 (N_3442,N_2246,N_2726);
xor U3443 (N_3443,N_2340,N_2589);
nand U3444 (N_3444,N_2770,N_2420);
nand U3445 (N_3445,N_2150,N_2200);
and U3446 (N_3446,N_2908,N_2508);
or U3447 (N_3447,N_2080,N_2321);
and U3448 (N_3448,N_2412,N_2460);
or U3449 (N_3449,N_2999,N_2154);
xnor U3450 (N_3450,N_2135,N_2020);
and U3451 (N_3451,N_2544,N_2692);
xor U3452 (N_3452,N_2166,N_2470);
nor U3453 (N_3453,N_2062,N_2249);
nor U3454 (N_3454,N_2651,N_2892);
nand U3455 (N_3455,N_2773,N_2286);
nand U3456 (N_3456,N_2472,N_2185);
and U3457 (N_3457,N_2068,N_2051);
nand U3458 (N_3458,N_2127,N_2430);
or U3459 (N_3459,N_2634,N_2885);
nor U3460 (N_3460,N_2814,N_2136);
and U3461 (N_3461,N_2851,N_2969);
nor U3462 (N_3462,N_2569,N_2626);
nor U3463 (N_3463,N_2390,N_2001);
or U3464 (N_3464,N_2276,N_2152);
xor U3465 (N_3465,N_2743,N_2000);
or U3466 (N_3466,N_2035,N_2957);
and U3467 (N_3467,N_2917,N_2011);
and U3468 (N_3468,N_2324,N_2534);
or U3469 (N_3469,N_2272,N_2038);
nand U3470 (N_3470,N_2766,N_2647);
xnor U3471 (N_3471,N_2288,N_2962);
and U3472 (N_3472,N_2140,N_2721);
nor U3473 (N_3473,N_2621,N_2864);
or U3474 (N_3474,N_2228,N_2333);
or U3475 (N_3475,N_2581,N_2668);
or U3476 (N_3476,N_2949,N_2425);
xnor U3477 (N_3477,N_2379,N_2580);
nand U3478 (N_3478,N_2772,N_2172);
or U3479 (N_3479,N_2523,N_2666);
or U3480 (N_3480,N_2852,N_2937);
nand U3481 (N_3481,N_2693,N_2317);
and U3482 (N_3482,N_2069,N_2275);
nand U3483 (N_3483,N_2133,N_2074);
xor U3484 (N_3484,N_2193,N_2282);
and U3485 (N_3485,N_2445,N_2005);
nand U3486 (N_3486,N_2572,N_2499);
xnor U3487 (N_3487,N_2209,N_2099);
nand U3488 (N_3488,N_2562,N_2096);
nand U3489 (N_3489,N_2824,N_2728);
and U3490 (N_3490,N_2345,N_2502);
or U3491 (N_3491,N_2982,N_2849);
nor U3492 (N_3492,N_2126,N_2241);
xor U3493 (N_3493,N_2316,N_2013);
nand U3494 (N_3494,N_2072,N_2927);
or U3495 (N_3495,N_2667,N_2315);
nand U3496 (N_3496,N_2218,N_2170);
nor U3497 (N_3497,N_2783,N_2215);
nor U3498 (N_3498,N_2169,N_2821);
nand U3499 (N_3499,N_2823,N_2019);
nand U3500 (N_3500,N_2327,N_2538);
nand U3501 (N_3501,N_2405,N_2526);
or U3502 (N_3502,N_2621,N_2070);
or U3503 (N_3503,N_2932,N_2276);
nand U3504 (N_3504,N_2286,N_2837);
nand U3505 (N_3505,N_2895,N_2008);
or U3506 (N_3506,N_2252,N_2999);
xnor U3507 (N_3507,N_2648,N_2449);
and U3508 (N_3508,N_2788,N_2185);
and U3509 (N_3509,N_2586,N_2849);
nor U3510 (N_3510,N_2963,N_2443);
or U3511 (N_3511,N_2435,N_2931);
nand U3512 (N_3512,N_2879,N_2724);
nand U3513 (N_3513,N_2041,N_2987);
nand U3514 (N_3514,N_2582,N_2050);
and U3515 (N_3515,N_2747,N_2826);
or U3516 (N_3516,N_2377,N_2203);
nand U3517 (N_3517,N_2544,N_2816);
nor U3518 (N_3518,N_2405,N_2050);
or U3519 (N_3519,N_2702,N_2608);
or U3520 (N_3520,N_2102,N_2824);
nor U3521 (N_3521,N_2858,N_2454);
nor U3522 (N_3522,N_2232,N_2390);
xnor U3523 (N_3523,N_2627,N_2780);
or U3524 (N_3524,N_2258,N_2444);
xor U3525 (N_3525,N_2692,N_2777);
nand U3526 (N_3526,N_2871,N_2130);
xnor U3527 (N_3527,N_2364,N_2418);
nand U3528 (N_3528,N_2045,N_2938);
and U3529 (N_3529,N_2239,N_2031);
or U3530 (N_3530,N_2964,N_2079);
and U3531 (N_3531,N_2889,N_2804);
or U3532 (N_3532,N_2289,N_2995);
nor U3533 (N_3533,N_2378,N_2003);
and U3534 (N_3534,N_2578,N_2704);
or U3535 (N_3535,N_2011,N_2710);
and U3536 (N_3536,N_2285,N_2856);
or U3537 (N_3537,N_2586,N_2883);
nor U3538 (N_3538,N_2825,N_2372);
xnor U3539 (N_3539,N_2027,N_2097);
nor U3540 (N_3540,N_2425,N_2627);
or U3541 (N_3541,N_2119,N_2284);
or U3542 (N_3542,N_2756,N_2818);
and U3543 (N_3543,N_2368,N_2544);
and U3544 (N_3544,N_2000,N_2415);
or U3545 (N_3545,N_2773,N_2941);
nand U3546 (N_3546,N_2482,N_2065);
nor U3547 (N_3547,N_2684,N_2348);
nand U3548 (N_3548,N_2323,N_2038);
nand U3549 (N_3549,N_2006,N_2553);
xnor U3550 (N_3550,N_2100,N_2343);
nor U3551 (N_3551,N_2691,N_2750);
xor U3552 (N_3552,N_2358,N_2407);
nor U3553 (N_3553,N_2482,N_2780);
nor U3554 (N_3554,N_2222,N_2669);
or U3555 (N_3555,N_2496,N_2942);
or U3556 (N_3556,N_2609,N_2913);
and U3557 (N_3557,N_2623,N_2696);
nand U3558 (N_3558,N_2873,N_2403);
and U3559 (N_3559,N_2278,N_2475);
xor U3560 (N_3560,N_2434,N_2429);
and U3561 (N_3561,N_2618,N_2123);
xor U3562 (N_3562,N_2378,N_2556);
nand U3563 (N_3563,N_2246,N_2881);
and U3564 (N_3564,N_2958,N_2869);
and U3565 (N_3565,N_2163,N_2511);
and U3566 (N_3566,N_2644,N_2064);
and U3567 (N_3567,N_2486,N_2259);
nor U3568 (N_3568,N_2316,N_2082);
xnor U3569 (N_3569,N_2946,N_2912);
nor U3570 (N_3570,N_2998,N_2023);
nor U3571 (N_3571,N_2836,N_2762);
and U3572 (N_3572,N_2821,N_2863);
nand U3573 (N_3573,N_2033,N_2699);
nand U3574 (N_3574,N_2871,N_2521);
and U3575 (N_3575,N_2498,N_2527);
nand U3576 (N_3576,N_2658,N_2593);
xnor U3577 (N_3577,N_2178,N_2531);
xnor U3578 (N_3578,N_2510,N_2680);
nand U3579 (N_3579,N_2588,N_2430);
or U3580 (N_3580,N_2485,N_2162);
and U3581 (N_3581,N_2398,N_2287);
nand U3582 (N_3582,N_2962,N_2489);
xnor U3583 (N_3583,N_2845,N_2748);
and U3584 (N_3584,N_2783,N_2260);
xnor U3585 (N_3585,N_2244,N_2700);
nand U3586 (N_3586,N_2772,N_2118);
or U3587 (N_3587,N_2222,N_2657);
and U3588 (N_3588,N_2550,N_2377);
or U3589 (N_3589,N_2918,N_2976);
nand U3590 (N_3590,N_2272,N_2509);
xnor U3591 (N_3591,N_2339,N_2174);
or U3592 (N_3592,N_2241,N_2218);
nand U3593 (N_3593,N_2103,N_2130);
xnor U3594 (N_3594,N_2709,N_2470);
nor U3595 (N_3595,N_2753,N_2877);
xor U3596 (N_3596,N_2225,N_2243);
and U3597 (N_3597,N_2133,N_2702);
xor U3598 (N_3598,N_2339,N_2553);
nor U3599 (N_3599,N_2695,N_2964);
xnor U3600 (N_3600,N_2547,N_2848);
or U3601 (N_3601,N_2188,N_2905);
nand U3602 (N_3602,N_2788,N_2879);
nand U3603 (N_3603,N_2508,N_2536);
xor U3604 (N_3604,N_2217,N_2048);
or U3605 (N_3605,N_2954,N_2218);
xnor U3606 (N_3606,N_2718,N_2794);
xor U3607 (N_3607,N_2770,N_2935);
and U3608 (N_3608,N_2898,N_2360);
and U3609 (N_3609,N_2011,N_2783);
nand U3610 (N_3610,N_2317,N_2555);
xnor U3611 (N_3611,N_2295,N_2595);
xnor U3612 (N_3612,N_2213,N_2864);
nor U3613 (N_3613,N_2253,N_2989);
or U3614 (N_3614,N_2163,N_2302);
and U3615 (N_3615,N_2691,N_2229);
nor U3616 (N_3616,N_2096,N_2413);
or U3617 (N_3617,N_2470,N_2392);
and U3618 (N_3618,N_2287,N_2631);
xnor U3619 (N_3619,N_2865,N_2774);
nand U3620 (N_3620,N_2323,N_2419);
nand U3621 (N_3621,N_2516,N_2101);
or U3622 (N_3622,N_2971,N_2970);
or U3623 (N_3623,N_2874,N_2770);
nor U3624 (N_3624,N_2026,N_2662);
nor U3625 (N_3625,N_2546,N_2115);
xnor U3626 (N_3626,N_2235,N_2372);
and U3627 (N_3627,N_2714,N_2489);
and U3628 (N_3628,N_2940,N_2018);
xnor U3629 (N_3629,N_2264,N_2238);
nand U3630 (N_3630,N_2030,N_2404);
nand U3631 (N_3631,N_2928,N_2508);
nor U3632 (N_3632,N_2940,N_2596);
or U3633 (N_3633,N_2416,N_2014);
nor U3634 (N_3634,N_2660,N_2029);
xor U3635 (N_3635,N_2207,N_2139);
or U3636 (N_3636,N_2104,N_2364);
nor U3637 (N_3637,N_2126,N_2277);
or U3638 (N_3638,N_2265,N_2628);
xnor U3639 (N_3639,N_2439,N_2097);
nand U3640 (N_3640,N_2720,N_2422);
nand U3641 (N_3641,N_2014,N_2175);
nor U3642 (N_3642,N_2120,N_2247);
nand U3643 (N_3643,N_2800,N_2591);
and U3644 (N_3644,N_2462,N_2411);
and U3645 (N_3645,N_2973,N_2468);
nor U3646 (N_3646,N_2195,N_2918);
nand U3647 (N_3647,N_2723,N_2432);
xnor U3648 (N_3648,N_2286,N_2367);
and U3649 (N_3649,N_2669,N_2941);
or U3650 (N_3650,N_2658,N_2763);
xor U3651 (N_3651,N_2317,N_2129);
nand U3652 (N_3652,N_2065,N_2727);
nand U3653 (N_3653,N_2027,N_2004);
nand U3654 (N_3654,N_2617,N_2171);
xor U3655 (N_3655,N_2272,N_2985);
or U3656 (N_3656,N_2740,N_2310);
or U3657 (N_3657,N_2888,N_2404);
or U3658 (N_3658,N_2082,N_2693);
and U3659 (N_3659,N_2125,N_2135);
and U3660 (N_3660,N_2504,N_2664);
and U3661 (N_3661,N_2067,N_2650);
nand U3662 (N_3662,N_2710,N_2002);
xor U3663 (N_3663,N_2704,N_2679);
nor U3664 (N_3664,N_2829,N_2151);
and U3665 (N_3665,N_2745,N_2833);
or U3666 (N_3666,N_2777,N_2903);
nand U3667 (N_3667,N_2975,N_2860);
nor U3668 (N_3668,N_2731,N_2533);
nor U3669 (N_3669,N_2706,N_2141);
nand U3670 (N_3670,N_2482,N_2434);
xnor U3671 (N_3671,N_2086,N_2573);
and U3672 (N_3672,N_2273,N_2762);
nand U3673 (N_3673,N_2575,N_2827);
and U3674 (N_3674,N_2687,N_2795);
nor U3675 (N_3675,N_2963,N_2893);
xnor U3676 (N_3676,N_2975,N_2513);
and U3677 (N_3677,N_2355,N_2548);
nand U3678 (N_3678,N_2561,N_2537);
or U3679 (N_3679,N_2163,N_2077);
or U3680 (N_3680,N_2625,N_2772);
nand U3681 (N_3681,N_2307,N_2018);
nand U3682 (N_3682,N_2777,N_2370);
or U3683 (N_3683,N_2750,N_2163);
and U3684 (N_3684,N_2189,N_2796);
nand U3685 (N_3685,N_2341,N_2031);
nand U3686 (N_3686,N_2919,N_2308);
and U3687 (N_3687,N_2662,N_2913);
or U3688 (N_3688,N_2421,N_2616);
xor U3689 (N_3689,N_2883,N_2993);
nor U3690 (N_3690,N_2020,N_2331);
nor U3691 (N_3691,N_2760,N_2879);
and U3692 (N_3692,N_2037,N_2809);
xor U3693 (N_3693,N_2712,N_2477);
nand U3694 (N_3694,N_2228,N_2840);
and U3695 (N_3695,N_2690,N_2682);
or U3696 (N_3696,N_2659,N_2091);
nor U3697 (N_3697,N_2022,N_2646);
nor U3698 (N_3698,N_2259,N_2481);
and U3699 (N_3699,N_2214,N_2814);
xnor U3700 (N_3700,N_2669,N_2232);
nor U3701 (N_3701,N_2088,N_2436);
or U3702 (N_3702,N_2557,N_2978);
or U3703 (N_3703,N_2609,N_2651);
or U3704 (N_3704,N_2027,N_2268);
or U3705 (N_3705,N_2646,N_2070);
or U3706 (N_3706,N_2010,N_2407);
or U3707 (N_3707,N_2735,N_2194);
and U3708 (N_3708,N_2771,N_2726);
or U3709 (N_3709,N_2570,N_2648);
xor U3710 (N_3710,N_2641,N_2351);
nand U3711 (N_3711,N_2894,N_2528);
nand U3712 (N_3712,N_2108,N_2448);
xor U3713 (N_3713,N_2807,N_2838);
nand U3714 (N_3714,N_2209,N_2111);
nand U3715 (N_3715,N_2875,N_2219);
nand U3716 (N_3716,N_2809,N_2591);
or U3717 (N_3717,N_2611,N_2046);
or U3718 (N_3718,N_2843,N_2153);
nand U3719 (N_3719,N_2676,N_2305);
or U3720 (N_3720,N_2038,N_2201);
or U3721 (N_3721,N_2851,N_2230);
xnor U3722 (N_3722,N_2118,N_2420);
nor U3723 (N_3723,N_2325,N_2800);
nand U3724 (N_3724,N_2840,N_2171);
nor U3725 (N_3725,N_2747,N_2335);
nand U3726 (N_3726,N_2152,N_2287);
nand U3727 (N_3727,N_2835,N_2948);
and U3728 (N_3728,N_2023,N_2333);
xnor U3729 (N_3729,N_2474,N_2080);
or U3730 (N_3730,N_2350,N_2129);
nor U3731 (N_3731,N_2765,N_2425);
xor U3732 (N_3732,N_2514,N_2957);
or U3733 (N_3733,N_2556,N_2742);
or U3734 (N_3734,N_2921,N_2227);
xnor U3735 (N_3735,N_2151,N_2302);
nor U3736 (N_3736,N_2802,N_2874);
and U3737 (N_3737,N_2380,N_2736);
xnor U3738 (N_3738,N_2009,N_2685);
nand U3739 (N_3739,N_2221,N_2675);
xor U3740 (N_3740,N_2085,N_2616);
and U3741 (N_3741,N_2318,N_2595);
xnor U3742 (N_3742,N_2665,N_2932);
and U3743 (N_3743,N_2151,N_2452);
or U3744 (N_3744,N_2634,N_2238);
and U3745 (N_3745,N_2873,N_2789);
nand U3746 (N_3746,N_2899,N_2489);
xnor U3747 (N_3747,N_2409,N_2436);
xor U3748 (N_3748,N_2680,N_2056);
and U3749 (N_3749,N_2329,N_2445);
xor U3750 (N_3750,N_2949,N_2294);
nor U3751 (N_3751,N_2053,N_2227);
or U3752 (N_3752,N_2113,N_2623);
and U3753 (N_3753,N_2155,N_2162);
nor U3754 (N_3754,N_2407,N_2576);
nand U3755 (N_3755,N_2454,N_2379);
nor U3756 (N_3756,N_2381,N_2221);
nand U3757 (N_3757,N_2821,N_2259);
nand U3758 (N_3758,N_2561,N_2654);
xor U3759 (N_3759,N_2998,N_2306);
nand U3760 (N_3760,N_2505,N_2561);
or U3761 (N_3761,N_2756,N_2974);
xnor U3762 (N_3762,N_2632,N_2158);
nor U3763 (N_3763,N_2694,N_2888);
or U3764 (N_3764,N_2464,N_2577);
xnor U3765 (N_3765,N_2978,N_2729);
nand U3766 (N_3766,N_2087,N_2300);
and U3767 (N_3767,N_2573,N_2053);
or U3768 (N_3768,N_2636,N_2652);
xnor U3769 (N_3769,N_2722,N_2794);
nand U3770 (N_3770,N_2869,N_2769);
or U3771 (N_3771,N_2343,N_2537);
nand U3772 (N_3772,N_2529,N_2201);
xnor U3773 (N_3773,N_2087,N_2534);
and U3774 (N_3774,N_2803,N_2030);
and U3775 (N_3775,N_2739,N_2094);
and U3776 (N_3776,N_2856,N_2846);
xnor U3777 (N_3777,N_2484,N_2244);
xor U3778 (N_3778,N_2073,N_2008);
nor U3779 (N_3779,N_2329,N_2437);
xor U3780 (N_3780,N_2174,N_2723);
xor U3781 (N_3781,N_2626,N_2822);
and U3782 (N_3782,N_2544,N_2117);
or U3783 (N_3783,N_2931,N_2718);
nand U3784 (N_3784,N_2651,N_2509);
or U3785 (N_3785,N_2562,N_2942);
xnor U3786 (N_3786,N_2665,N_2860);
nand U3787 (N_3787,N_2452,N_2861);
nand U3788 (N_3788,N_2840,N_2860);
or U3789 (N_3789,N_2367,N_2479);
and U3790 (N_3790,N_2184,N_2693);
xor U3791 (N_3791,N_2804,N_2411);
nand U3792 (N_3792,N_2137,N_2250);
nand U3793 (N_3793,N_2182,N_2465);
or U3794 (N_3794,N_2111,N_2674);
and U3795 (N_3795,N_2815,N_2108);
nor U3796 (N_3796,N_2527,N_2208);
nor U3797 (N_3797,N_2050,N_2888);
and U3798 (N_3798,N_2699,N_2539);
or U3799 (N_3799,N_2321,N_2306);
or U3800 (N_3800,N_2289,N_2788);
and U3801 (N_3801,N_2847,N_2871);
or U3802 (N_3802,N_2390,N_2199);
and U3803 (N_3803,N_2338,N_2442);
nand U3804 (N_3804,N_2507,N_2189);
nor U3805 (N_3805,N_2590,N_2734);
nor U3806 (N_3806,N_2269,N_2805);
xnor U3807 (N_3807,N_2889,N_2701);
nand U3808 (N_3808,N_2951,N_2926);
and U3809 (N_3809,N_2422,N_2608);
xor U3810 (N_3810,N_2433,N_2364);
xnor U3811 (N_3811,N_2914,N_2660);
xnor U3812 (N_3812,N_2472,N_2314);
xnor U3813 (N_3813,N_2181,N_2995);
nand U3814 (N_3814,N_2626,N_2767);
xnor U3815 (N_3815,N_2706,N_2653);
or U3816 (N_3816,N_2425,N_2319);
nor U3817 (N_3817,N_2178,N_2719);
or U3818 (N_3818,N_2839,N_2160);
xnor U3819 (N_3819,N_2698,N_2337);
nand U3820 (N_3820,N_2426,N_2924);
xnor U3821 (N_3821,N_2527,N_2622);
xnor U3822 (N_3822,N_2311,N_2569);
xor U3823 (N_3823,N_2067,N_2232);
and U3824 (N_3824,N_2614,N_2646);
and U3825 (N_3825,N_2891,N_2388);
or U3826 (N_3826,N_2114,N_2001);
nand U3827 (N_3827,N_2224,N_2809);
nor U3828 (N_3828,N_2557,N_2219);
nor U3829 (N_3829,N_2267,N_2023);
nor U3830 (N_3830,N_2234,N_2639);
nand U3831 (N_3831,N_2414,N_2337);
or U3832 (N_3832,N_2396,N_2163);
xnor U3833 (N_3833,N_2891,N_2344);
nand U3834 (N_3834,N_2256,N_2145);
nand U3835 (N_3835,N_2728,N_2645);
or U3836 (N_3836,N_2920,N_2004);
and U3837 (N_3837,N_2172,N_2618);
and U3838 (N_3838,N_2646,N_2164);
nand U3839 (N_3839,N_2199,N_2702);
and U3840 (N_3840,N_2691,N_2621);
or U3841 (N_3841,N_2756,N_2509);
nand U3842 (N_3842,N_2326,N_2501);
nor U3843 (N_3843,N_2120,N_2085);
nor U3844 (N_3844,N_2158,N_2760);
nor U3845 (N_3845,N_2603,N_2295);
nor U3846 (N_3846,N_2925,N_2164);
nand U3847 (N_3847,N_2688,N_2263);
and U3848 (N_3848,N_2557,N_2569);
xnor U3849 (N_3849,N_2195,N_2850);
nor U3850 (N_3850,N_2580,N_2658);
xnor U3851 (N_3851,N_2331,N_2244);
or U3852 (N_3852,N_2587,N_2489);
nand U3853 (N_3853,N_2168,N_2058);
xor U3854 (N_3854,N_2371,N_2155);
or U3855 (N_3855,N_2485,N_2224);
or U3856 (N_3856,N_2561,N_2596);
or U3857 (N_3857,N_2227,N_2763);
and U3858 (N_3858,N_2908,N_2856);
or U3859 (N_3859,N_2673,N_2119);
or U3860 (N_3860,N_2931,N_2103);
nand U3861 (N_3861,N_2675,N_2359);
or U3862 (N_3862,N_2157,N_2641);
and U3863 (N_3863,N_2344,N_2366);
nor U3864 (N_3864,N_2295,N_2519);
or U3865 (N_3865,N_2020,N_2930);
or U3866 (N_3866,N_2735,N_2464);
nand U3867 (N_3867,N_2419,N_2079);
and U3868 (N_3868,N_2263,N_2248);
and U3869 (N_3869,N_2832,N_2785);
and U3870 (N_3870,N_2906,N_2734);
or U3871 (N_3871,N_2757,N_2867);
nor U3872 (N_3872,N_2486,N_2621);
nand U3873 (N_3873,N_2953,N_2560);
nor U3874 (N_3874,N_2375,N_2114);
xnor U3875 (N_3875,N_2496,N_2482);
xor U3876 (N_3876,N_2453,N_2432);
nand U3877 (N_3877,N_2551,N_2785);
nor U3878 (N_3878,N_2515,N_2221);
nand U3879 (N_3879,N_2066,N_2247);
nor U3880 (N_3880,N_2523,N_2767);
nor U3881 (N_3881,N_2005,N_2340);
and U3882 (N_3882,N_2153,N_2367);
or U3883 (N_3883,N_2759,N_2362);
nand U3884 (N_3884,N_2318,N_2701);
nand U3885 (N_3885,N_2576,N_2585);
or U3886 (N_3886,N_2208,N_2496);
or U3887 (N_3887,N_2811,N_2144);
and U3888 (N_3888,N_2378,N_2145);
nor U3889 (N_3889,N_2006,N_2859);
nand U3890 (N_3890,N_2645,N_2126);
nor U3891 (N_3891,N_2454,N_2692);
nand U3892 (N_3892,N_2464,N_2209);
nor U3893 (N_3893,N_2576,N_2378);
nand U3894 (N_3894,N_2440,N_2746);
nor U3895 (N_3895,N_2110,N_2671);
or U3896 (N_3896,N_2600,N_2931);
and U3897 (N_3897,N_2396,N_2381);
and U3898 (N_3898,N_2053,N_2417);
and U3899 (N_3899,N_2927,N_2012);
nand U3900 (N_3900,N_2716,N_2415);
xor U3901 (N_3901,N_2234,N_2073);
nor U3902 (N_3902,N_2902,N_2257);
and U3903 (N_3903,N_2015,N_2206);
nor U3904 (N_3904,N_2541,N_2872);
xor U3905 (N_3905,N_2447,N_2102);
or U3906 (N_3906,N_2155,N_2721);
nand U3907 (N_3907,N_2239,N_2774);
xor U3908 (N_3908,N_2344,N_2442);
nor U3909 (N_3909,N_2480,N_2018);
nor U3910 (N_3910,N_2857,N_2303);
xor U3911 (N_3911,N_2950,N_2213);
xnor U3912 (N_3912,N_2045,N_2440);
nor U3913 (N_3913,N_2077,N_2027);
nand U3914 (N_3914,N_2661,N_2949);
or U3915 (N_3915,N_2467,N_2869);
nand U3916 (N_3916,N_2751,N_2309);
or U3917 (N_3917,N_2810,N_2673);
or U3918 (N_3918,N_2960,N_2901);
nor U3919 (N_3919,N_2084,N_2896);
and U3920 (N_3920,N_2493,N_2629);
nand U3921 (N_3921,N_2646,N_2315);
nand U3922 (N_3922,N_2477,N_2065);
and U3923 (N_3923,N_2850,N_2984);
nand U3924 (N_3924,N_2423,N_2390);
and U3925 (N_3925,N_2819,N_2902);
nand U3926 (N_3926,N_2921,N_2443);
and U3927 (N_3927,N_2203,N_2284);
nand U3928 (N_3928,N_2481,N_2336);
nor U3929 (N_3929,N_2596,N_2487);
nor U3930 (N_3930,N_2329,N_2642);
or U3931 (N_3931,N_2350,N_2121);
nor U3932 (N_3932,N_2527,N_2469);
nand U3933 (N_3933,N_2016,N_2445);
nand U3934 (N_3934,N_2033,N_2168);
nor U3935 (N_3935,N_2140,N_2592);
xnor U3936 (N_3936,N_2307,N_2165);
nand U3937 (N_3937,N_2143,N_2174);
nor U3938 (N_3938,N_2152,N_2841);
and U3939 (N_3939,N_2697,N_2440);
nor U3940 (N_3940,N_2254,N_2407);
and U3941 (N_3941,N_2832,N_2038);
nand U3942 (N_3942,N_2075,N_2489);
and U3943 (N_3943,N_2353,N_2270);
and U3944 (N_3944,N_2324,N_2656);
nor U3945 (N_3945,N_2658,N_2565);
nand U3946 (N_3946,N_2811,N_2636);
or U3947 (N_3947,N_2825,N_2490);
and U3948 (N_3948,N_2948,N_2193);
and U3949 (N_3949,N_2606,N_2298);
nand U3950 (N_3950,N_2942,N_2567);
xnor U3951 (N_3951,N_2261,N_2900);
nor U3952 (N_3952,N_2790,N_2745);
and U3953 (N_3953,N_2516,N_2671);
or U3954 (N_3954,N_2429,N_2636);
nand U3955 (N_3955,N_2123,N_2182);
xor U3956 (N_3956,N_2978,N_2841);
nand U3957 (N_3957,N_2526,N_2972);
nand U3958 (N_3958,N_2240,N_2819);
nand U3959 (N_3959,N_2428,N_2541);
and U3960 (N_3960,N_2512,N_2754);
xnor U3961 (N_3961,N_2969,N_2976);
nor U3962 (N_3962,N_2205,N_2464);
nor U3963 (N_3963,N_2794,N_2189);
and U3964 (N_3964,N_2683,N_2936);
nand U3965 (N_3965,N_2555,N_2156);
and U3966 (N_3966,N_2220,N_2981);
xor U3967 (N_3967,N_2680,N_2506);
or U3968 (N_3968,N_2966,N_2904);
and U3969 (N_3969,N_2780,N_2643);
or U3970 (N_3970,N_2096,N_2546);
xor U3971 (N_3971,N_2674,N_2123);
or U3972 (N_3972,N_2452,N_2697);
or U3973 (N_3973,N_2203,N_2892);
nor U3974 (N_3974,N_2195,N_2987);
and U3975 (N_3975,N_2039,N_2910);
or U3976 (N_3976,N_2869,N_2658);
and U3977 (N_3977,N_2920,N_2052);
nand U3978 (N_3978,N_2137,N_2734);
xor U3979 (N_3979,N_2289,N_2931);
nand U3980 (N_3980,N_2026,N_2268);
xnor U3981 (N_3981,N_2383,N_2355);
nand U3982 (N_3982,N_2594,N_2990);
or U3983 (N_3983,N_2580,N_2626);
or U3984 (N_3984,N_2530,N_2554);
nor U3985 (N_3985,N_2927,N_2641);
nand U3986 (N_3986,N_2332,N_2545);
or U3987 (N_3987,N_2533,N_2604);
nand U3988 (N_3988,N_2777,N_2994);
nor U3989 (N_3989,N_2633,N_2635);
or U3990 (N_3990,N_2711,N_2354);
nand U3991 (N_3991,N_2083,N_2504);
xor U3992 (N_3992,N_2633,N_2764);
nor U3993 (N_3993,N_2161,N_2879);
or U3994 (N_3994,N_2314,N_2993);
and U3995 (N_3995,N_2663,N_2630);
or U3996 (N_3996,N_2645,N_2928);
and U3997 (N_3997,N_2707,N_2626);
or U3998 (N_3998,N_2222,N_2085);
nor U3999 (N_3999,N_2086,N_2239);
and U4000 (N_4000,N_3905,N_3166);
xor U4001 (N_4001,N_3473,N_3726);
nor U4002 (N_4002,N_3915,N_3836);
nand U4003 (N_4003,N_3320,N_3614);
and U4004 (N_4004,N_3510,N_3758);
nand U4005 (N_4005,N_3385,N_3045);
xor U4006 (N_4006,N_3828,N_3759);
or U4007 (N_4007,N_3893,N_3435);
or U4008 (N_4008,N_3953,N_3808);
nor U4009 (N_4009,N_3192,N_3978);
and U4010 (N_4010,N_3232,N_3704);
nor U4011 (N_4011,N_3351,N_3838);
and U4012 (N_4012,N_3445,N_3273);
and U4013 (N_4013,N_3989,N_3881);
nand U4014 (N_4014,N_3007,N_3408);
nand U4015 (N_4015,N_3278,N_3847);
nor U4016 (N_4016,N_3244,N_3465);
xnor U4017 (N_4017,N_3238,N_3246);
nand U4018 (N_4018,N_3610,N_3991);
xnor U4019 (N_4019,N_3210,N_3720);
xor U4020 (N_4020,N_3426,N_3670);
xor U4021 (N_4021,N_3032,N_3139);
and U4022 (N_4022,N_3441,N_3622);
or U4023 (N_4023,N_3528,N_3060);
nand U4024 (N_4024,N_3804,N_3392);
and U4025 (N_4025,N_3458,N_3715);
xnor U4026 (N_4026,N_3163,N_3005);
nor U4027 (N_4027,N_3697,N_3906);
and U4028 (N_4028,N_3405,N_3855);
nand U4029 (N_4029,N_3868,N_3523);
nor U4030 (N_4030,N_3197,N_3586);
xnor U4031 (N_4031,N_3652,N_3269);
nand U4032 (N_4032,N_3006,N_3186);
xnor U4033 (N_4033,N_3409,N_3829);
and U4034 (N_4034,N_3695,N_3690);
and U4035 (N_4035,N_3677,N_3290);
xnor U4036 (N_4036,N_3171,N_3025);
and U4037 (N_4037,N_3329,N_3038);
or U4038 (N_4038,N_3455,N_3875);
or U4039 (N_4039,N_3575,N_3433);
nand U4040 (N_4040,N_3599,N_3755);
nand U4041 (N_4041,N_3135,N_3041);
and U4042 (N_4042,N_3822,N_3176);
nand U4043 (N_4043,N_3093,N_3365);
xor U4044 (N_4044,N_3656,N_3647);
or U4045 (N_4045,N_3084,N_3352);
and U4046 (N_4046,N_3078,N_3902);
nand U4047 (N_4047,N_3292,N_3702);
and U4048 (N_4048,N_3860,N_3361);
xor U4049 (N_4049,N_3844,N_3810);
or U4050 (N_4050,N_3371,N_3977);
and U4051 (N_4051,N_3559,N_3850);
and U4052 (N_4052,N_3423,N_3250);
nor U4053 (N_4053,N_3223,N_3574);
xor U4054 (N_4054,N_3536,N_3279);
xnor U4055 (N_4055,N_3616,N_3681);
nor U4056 (N_4056,N_3260,N_3551);
nand U4057 (N_4057,N_3098,N_3722);
xor U4058 (N_4058,N_3561,N_3733);
or U4059 (N_4059,N_3555,N_3706);
and U4060 (N_4060,N_3598,N_3628);
nand U4061 (N_4061,N_3427,N_3799);
and U4062 (N_4062,N_3519,N_3757);
nor U4063 (N_4063,N_3132,N_3456);
nand U4064 (N_4064,N_3499,N_3079);
xnor U4065 (N_4065,N_3887,N_3737);
xor U4066 (N_4066,N_3992,N_3149);
xnor U4067 (N_4067,N_3676,N_3595);
and U4068 (N_4068,N_3699,N_3222);
nand U4069 (N_4069,N_3162,N_3212);
and U4070 (N_4070,N_3861,N_3487);
xnor U4071 (N_4071,N_3907,N_3087);
nor U4072 (N_4072,N_3151,N_3106);
nor U4073 (N_4073,N_3332,N_3736);
nand U4074 (N_4074,N_3515,N_3783);
nand U4075 (N_4075,N_3619,N_3140);
and U4076 (N_4076,N_3023,N_3390);
and U4077 (N_4077,N_3539,N_3230);
xnor U4078 (N_4078,N_3065,N_3888);
nand U4079 (N_4079,N_3129,N_3201);
xnor U4080 (N_4080,N_3634,N_3734);
xnor U4081 (N_4081,N_3476,N_3741);
nor U4082 (N_4082,N_3196,N_3679);
or U4083 (N_4083,N_3374,N_3285);
xor U4084 (N_4084,N_3781,N_3090);
nand U4085 (N_4085,N_3957,N_3096);
xnor U4086 (N_4086,N_3545,N_3483);
xnor U4087 (N_4087,N_3767,N_3771);
and U4088 (N_4088,N_3571,N_3011);
xnor U4089 (N_4089,N_3412,N_3434);
nor U4090 (N_4090,N_3621,N_3219);
and U4091 (N_4091,N_3117,N_3908);
xor U4092 (N_4092,N_3788,N_3251);
or U4093 (N_4093,N_3396,N_3931);
nand U4094 (N_4094,N_3694,N_3589);
nand U4095 (N_4095,N_3958,N_3389);
nand U4096 (N_4096,N_3698,N_3101);
nor U4097 (N_4097,N_3313,N_3198);
nor U4098 (N_4098,N_3266,N_3233);
nor U4099 (N_4099,N_3779,N_3322);
or U4100 (N_4100,N_3760,N_3933);
nor U4101 (N_4101,N_3301,N_3059);
or U4102 (N_4102,N_3752,N_3504);
xnor U4103 (N_4103,N_3972,N_3985);
nand U4104 (N_4104,N_3790,N_3089);
and U4105 (N_4105,N_3270,N_3814);
or U4106 (N_4106,N_3912,N_3770);
and U4107 (N_4107,N_3310,N_3832);
nor U4108 (N_4108,N_3379,N_3378);
nand U4109 (N_4109,N_3410,N_3961);
xnor U4110 (N_4110,N_3144,N_3597);
nor U4111 (N_4111,N_3497,N_3833);
or U4112 (N_4112,N_3926,N_3678);
and U4113 (N_4113,N_3029,N_3347);
xnor U4114 (N_4114,N_3827,N_3801);
and U4115 (N_4115,N_3248,N_3463);
xor U4116 (N_4116,N_3319,N_3493);
nor U4117 (N_4117,N_3054,N_3094);
or U4118 (N_4118,N_3451,N_3877);
or U4119 (N_4119,N_3685,N_3959);
or U4120 (N_4120,N_3184,N_3466);
nand U4121 (N_4121,N_3395,N_3500);
or U4122 (N_4122,N_3126,N_3540);
or U4123 (N_4123,N_3928,N_3590);
xor U4124 (N_4124,N_3274,N_3026);
and U4125 (N_4125,N_3208,N_3398);
nor U4126 (N_4126,N_3729,N_3717);
or U4127 (N_4127,N_3055,N_3406);
and U4128 (N_4128,N_3228,N_3929);
and U4129 (N_4129,N_3563,N_3343);
xnor U4130 (N_4130,N_3603,N_3857);
nor U4131 (N_4131,N_3107,N_3088);
nand U4132 (N_4132,N_3271,N_3159);
xor U4133 (N_4133,N_3534,N_3582);
nand U4134 (N_4134,N_3448,N_3360);
nor U4135 (N_4135,N_3998,N_3321);
nand U4136 (N_4136,N_3588,N_3158);
nor U4137 (N_4137,N_3895,N_3138);
or U4138 (N_4138,N_3180,N_3155);
nand U4139 (N_4139,N_3524,N_3795);
nor U4140 (N_4140,N_3963,N_3482);
nor U4141 (N_4141,N_3876,N_3130);
or U4142 (N_4142,N_3899,N_3359);
or U4143 (N_4143,N_3843,N_3592);
and U4144 (N_4144,N_3606,N_3852);
and U4145 (N_4145,N_3886,N_3520);
nand U4146 (N_4146,N_3743,N_3607);
nand U4147 (N_4147,N_3775,N_3999);
nand U4148 (N_4148,N_3214,N_3203);
or U4149 (N_4149,N_3567,N_3542);
or U4150 (N_4150,N_3348,N_3611);
and U4151 (N_4151,N_3327,N_3917);
or U4152 (N_4152,N_3921,N_3234);
and U4153 (N_4153,N_3751,N_3630);
and U4154 (N_4154,N_3550,N_3108);
nand U4155 (N_4155,N_3115,N_3541);
nor U4156 (N_4156,N_3514,N_3627);
and U4157 (N_4157,N_3768,N_3629);
or U4158 (N_4158,N_3284,N_3331);
and U4159 (N_4159,N_3420,N_3552);
and U4160 (N_4160,N_3370,N_3046);
and U4161 (N_4161,N_3037,N_3485);
nor U4162 (N_4162,N_3909,N_3478);
or U4163 (N_4163,N_3438,N_3930);
or U4164 (N_4164,N_3713,N_3355);
xor U4165 (N_4165,N_3245,N_3511);
nor U4166 (N_4166,N_3402,N_3587);
or U4167 (N_4167,N_3030,N_3071);
nand U4168 (N_4168,N_3095,N_3732);
nor U4169 (N_4169,N_3145,N_3063);
nor U4170 (N_4170,N_3318,N_3707);
or U4171 (N_4171,N_3010,N_3818);
xor U4172 (N_4172,N_3177,N_3739);
xor U4173 (N_4173,N_3692,N_3718);
xnor U4174 (N_4174,N_3668,N_3995);
nor U4175 (N_4175,N_3572,N_3501);
nor U4176 (N_4176,N_3287,N_3787);
xnor U4177 (N_4177,N_3874,N_3394);
or U4178 (N_4178,N_3036,N_3489);
xnor U4179 (N_4179,N_3048,N_3944);
nor U4180 (N_4180,N_3967,N_3856);
or U4181 (N_4181,N_3017,N_3137);
or U4182 (N_4182,N_3807,N_3068);
and U4183 (N_4183,N_3311,N_3666);
and U4184 (N_4184,N_3724,N_3892);
or U4185 (N_4185,N_3020,N_3502);
or U4186 (N_4186,N_3073,N_3765);
and U4187 (N_4187,N_3806,N_3104);
or U4188 (N_4188,N_3649,N_3798);
or U4189 (N_4189,N_3064,N_3546);
xor U4190 (N_4190,N_3811,N_3272);
or U4191 (N_4191,N_3018,N_3033);
nor U4192 (N_4192,N_3253,N_3125);
nand U4193 (N_4193,N_3820,N_3609);
or U4194 (N_4194,N_3070,N_3053);
or U4195 (N_4195,N_3143,N_3112);
and U4196 (N_4196,N_3263,N_3825);
nand U4197 (N_4197,N_3935,N_3920);
and U4198 (N_4198,N_3276,N_3031);
nor U4199 (N_4199,N_3333,N_3134);
and U4200 (N_4200,N_3951,N_3740);
nand U4201 (N_4201,N_3674,N_3305);
or U4202 (N_4202,N_3687,N_3527);
nand U4203 (N_4203,N_3646,N_3291);
or U4204 (N_4204,N_3346,N_3488);
or U4205 (N_4205,N_3858,N_3748);
or U4206 (N_4206,N_3211,N_3579);
and U4207 (N_4207,N_3675,N_3264);
xnor U4208 (N_4208,N_3657,N_3444);
xor U4209 (N_4209,N_3436,N_3239);
nand U4210 (N_4210,N_3190,N_3517);
nand U4211 (N_4211,N_3911,N_3826);
nor U4212 (N_4212,N_3954,N_3086);
xor U4213 (N_4213,N_3034,N_3625);
xor U4214 (N_4214,N_3518,N_3167);
nand U4215 (N_4215,N_3979,N_3131);
nand U4216 (N_4216,N_3334,N_3654);
nand U4217 (N_4217,N_3160,N_3056);
nand U4218 (N_4218,N_3941,N_3593);
xor U4219 (N_4219,N_3753,N_3633);
nand U4220 (N_4220,N_3261,N_3372);
and U4221 (N_4221,N_3735,N_3462);
and U4222 (N_4222,N_3164,N_3342);
nor U4223 (N_4223,N_3047,N_3431);
or U4224 (N_4224,N_3994,N_3267);
or U4225 (N_4225,N_3114,N_3213);
and U4226 (N_4226,N_3452,N_3797);
and U4227 (N_4227,N_3050,N_3354);
nor U4228 (N_4228,N_3884,N_3437);
or U4229 (N_4229,N_3612,N_3848);
nand U4230 (N_4230,N_3618,N_3682);
nor U4231 (N_4231,N_3224,N_3146);
xor U4232 (N_4232,N_3865,N_3309);
xnor U4233 (N_4233,N_3472,N_3731);
or U4234 (N_4234,N_3866,N_3387);
or U4235 (N_4235,N_3430,N_3522);
and U4236 (N_4236,N_3468,N_3871);
nor U4237 (N_4237,N_3328,N_3965);
nor U4238 (N_4238,N_3058,N_3791);
and U4239 (N_4239,N_3357,N_3154);
nor U4240 (N_4240,N_3632,N_3624);
xor U4241 (N_4241,N_3970,N_3557);
nand U4242 (N_4242,N_3716,N_3766);
nor U4243 (N_4243,N_3450,N_3968);
nor U4244 (N_4244,N_3072,N_3035);
xnor U4245 (N_4245,N_3262,N_3415);
nor U4246 (N_4246,N_3532,N_3446);
or U4247 (N_4247,N_3174,N_3764);
xnor U4248 (N_4248,N_3317,N_3794);
or U4249 (N_4249,N_3604,N_3216);
nand U4250 (N_4250,N_3742,N_3853);
nand U4251 (N_4251,N_3120,N_3560);
and U4252 (N_4252,N_3596,N_3282);
nand U4253 (N_4253,N_3424,N_3823);
nor U4254 (N_4254,N_3118,N_3157);
nand U4255 (N_4255,N_3353,N_3001);
or U4256 (N_4256,N_3756,N_3252);
nand U4257 (N_4257,N_3181,N_3401);
nand U4258 (N_4258,N_3513,N_3529);
nor U4259 (N_4259,N_3123,N_3039);
or U4260 (N_4260,N_3049,N_3383);
nand U4261 (N_4261,N_3531,N_3012);
or U4262 (N_4262,N_3636,N_3496);
nand U4263 (N_4263,N_3439,N_3846);
or U4264 (N_4264,N_3635,N_3242);
nand U4265 (N_4265,N_3200,N_3339);
or U4266 (N_4266,N_3639,N_3879);
nor U4267 (N_4267,N_3870,N_3377);
nand U4268 (N_4268,N_3367,N_3659);
and U4269 (N_4269,N_3882,N_3962);
xnor U4270 (N_4270,N_3363,N_3470);
and U4271 (N_4271,N_3845,N_3165);
nor U4272 (N_4272,N_3976,N_3044);
xor U4273 (N_4273,N_3939,N_3916);
xor U4274 (N_4274,N_3074,N_3591);
or U4275 (N_4275,N_3016,N_3404);
nor U4276 (N_4276,N_3169,N_3308);
nor U4277 (N_4277,N_3386,N_3314);
or U4278 (N_4278,N_3113,N_3092);
xnor U4279 (N_4279,N_3672,N_3507);
or U4280 (N_4280,N_3231,N_3744);
and U4281 (N_4281,N_3240,N_3340);
xor U4282 (N_4282,N_3133,N_3793);
nor U4283 (N_4283,N_3658,N_3417);
nor U4284 (N_4284,N_3076,N_3295);
xnor U4285 (N_4285,N_3680,N_3964);
nor U4286 (N_4286,N_3600,N_3701);
and U4287 (N_4287,N_3110,N_3102);
nand U4288 (N_4288,N_3014,N_3040);
nor U4289 (N_4289,N_3924,N_3443);
and U4290 (N_4290,N_3300,N_3696);
or U4291 (N_4291,N_3819,N_3194);
and U4292 (N_4292,N_3221,N_3003);
nand U4293 (N_4293,N_3712,N_3277);
nor U4294 (N_4294,N_3471,N_3283);
or U4295 (N_4295,N_3000,N_3583);
xor U4296 (N_4296,N_3459,N_3626);
or U4297 (N_4297,N_3193,N_3185);
xor U4298 (N_4298,N_3199,N_3710);
and U4299 (N_4299,N_3693,N_3449);
and U4300 (N_4300,N_3225,N_3650);
and U4301 (N_4301,N_3854,N_3631);
nand U4302 (N_4302,N_3684,N_3189);
nor U4303 (N_4303,N_3898,N_3565);
nor U4304 (N_4304,N_3350,N_3432);
nand U4305 (N_4305,N_3268,N_3306);
or U4306 (N_4306,N_3457,N_3467);
nand U4307 (N_4307,N_3413,N_3477);
or U4308 (N_4308,N_3368,N_3688);
xor U4309 (N_4309,N_3303,N_3175);
nor U4310 (N_4310,N_3913,N_3091);
nand U4311 (N_4311,N_3027,N_3265);
or U4312 (N_4312,N_3789,N_3229);
and U4313 (N_4313,N_3289,N_3883);
nand U4314 (N_4314,N_3453,N_3393);
xnor U4315 (N_4315,N_3066,N_3548);
and U4316 (N_4316,N_3356,N_3111);
xor U4317 (N_4317,N_3705,N_3925);
and U4318 (N_4318,N_3547,N_3864);
nand U4319 (N_4319,N_3975,N_3516);
xnor U4320 (N_4320,N_3460,N_3100);
nor U4321 (N_4321,N_3172,N_3996);
or U4322 (N_4322,N_3257,N_3577);
or U4323 (N_4323,N_3168,N_3227);
nor U4324 (N_4324,N_3824,N_3894);
nor U4325 (N_4325,N_3554,N_3640);
nand U4326 (N_4326,N_3950,N_3971);
nor U4327 (N_4327,N_3099,N_3642);
nand U4328 (N_4328,N_3486,N_3097);
nand U4329 (N_4329,N_3982,N_3254);
and U4330 (N_4330,N_3558,N_3419);
and U4331 (N_4331,N_3136,N_3400);
and U4332 (N_4332,N_3296,N_3988);
and U4333 (N_4333,N_3904,N_3878);
xor U4334 (N_4334,N_3147,N_3745);
nand U4335 (N_4335,N_3608,N_3660);
or U4336 (N_4336,N_3324,N_3969);
nand U4337 (N_4337,N_3960,N_3564);
nor U4338 (N_4338,N_3298,N_3307);
xnor U4339 (N_4339,N_3543,N_3637);
xor U4340 (N_4340,N_3206,N_3304);
nor U4341 (N_4341,N_3188,N_3947);
nor U4342 (N_4342,N_3416,N_3837);
nand U4343 (N_4343,N_3121,N_3683);
nor U4344 (N_4344,N_3815,N_3537);
nor U4345 (N_4345,N_3966,N_3021);
nand U4346 (N_4346,N_3220,N_3255);
nand U4347 (N_4347,N_3335,N_3336);
xor U4348 (N_4348,N_3051,N_3341);
nor U4349 (N_4349,N_3152,N_3484);
and U4350 (N_4350,N_3873,N_3601);
nand U4351 (N_4351,N_3803,N_3015);
and U4352 (N_4352,N_3568,N_3330);
xor U4353 (N_4353,N_3421,N_3491);
nand U4354 (N_4354,N_3796,N_3566);
nand U4355 (N_4355,N_3780,N_3105);
or U4356 (N_4356,N_3890,N_3075);
nand U4357 (N_4357,N_3358,N_3019);
or U4358 (N_4358,N_3669,N_3187);
nor U4359 (N_4359,N_3830,N_3281);
nor U4360 (N_4360,N_3872,N_3956);
or U4361 (N_4361,N_3721,N_3122);
or U4362 (N_4362,N_3509,N_3384);
or U4363 (N_4363,N_3952,N_3506);
or U4364 (N_4364,N_3573,N_3288);
or U4365 (N_4365,N_3127,N_3119);
and U4366 (N_4366,N_3161,N_3946);
nor U4367 (N_4367,N_3576,N_3889);
and U4368 (N_4368,N_3299,N_3142);
and U4369 (N_4369,N_3425,N_3345);
nand U4370 (N_4370,N_3776,N_3259);
nor U4371 (N_4371,N_3762,N_3816);
nor U4372 (N_4372,N_3839,N_3024);
nor U4373 (N_4373,N_3191,N_3851);
and U4374 (N_4374,N_3863,N_3247);
or U4375 (N_4375,N_3938,N_3241);
nand U4376 (N_4376,N_3217,N_3062);
and U4377 (N_4377,N_3205,N_3662);
and U4378 (N_4378,N_3813,N_3556);
nor U4379 (N_4379,N_3580,N_3043);
nor U4380 (N_4380,N_3570,N_3936);
xor U4381 (N_4381,N_3834,N_3900);
and U4382 (N_4382,N_3215,N_3664);
and U4383 (N_4383,N_3562,N_3178);
and U4384 (N_4384,N_3842,N_3042);
nand U4385 (N_4385,N_3896,N_3381);
and U4386 (N_4386,N_3613,N_3934);
and U4387 (N_4387,N_3725,N_3464);
or U4388 (N_4388,N_3312,N_3256);
xor U4389 (N_4389,N_3337,N_3204);
xnor U4390 (N_4390,N_3326,N_3578);
nand U4391 (N_4391,N_3376,N_3763);
and U4392 (N_4392,N_3237,N_3508);
nand U4393 (N_4393,N_3981,N_3013);
or U4394 (N_4394,N_3785,N_3773);
nor U4395 (N_4395,N_3746,N_3083);
xor U4396 (N_4396,N_3569,N_3218);
and U4397 (N_4397,N_3057,N_3605);
and U4398 (N_4398,N_3835,N_3533);
or U4399 (N_4399,N_3081,N_3403);
nor U4400 (N_4400,N_3480,N_3802);
or U4401 (N_4401,N_3997,N_3974);
nand U4402 (N_4402,N_3280,N_3648);
xnor U4403 (N_4403,N_3148,N_3711);
xor U4404 (N_4404,N_3859,N_3004);
and U4405 (N_4405,N_3407,N_3769);
and U4406 (N_4406,N_3067,N_3170);
xnor U4407 (N_4407,N_3525,N_3549);
xnor U4408 (N_4408,N_3922,N_3109);
or U4409 (N_4409,N_3236,N_3077);
nor U4410 (N_4410,N_3620,N_3869);
nor U4411 (N_4411,N_3812,N_3945);
and U4412 (N_4412,N_3082,N_3469);
nand U4413 (N_4413,N_3862,N_3990);
xnor U4414 (N_4414,N_3885,N_3479);
nand U4415 (N_4415,N_3923,N_3919);
and U4416 (N_4416,N_3901,N_3349);
xor U4417 (N_4417,N_3738,N_3209);
xnor U4418 (N_4418,N_3411,N_3891);
nor U4419 (N_4419,N_3987,N_3986);
nand U4420 (N_4420,N_3344,N_3821);
xor U4421 (N_4421,N_3526,N_3382);
nand U4422 (N_4422,N_3817,N_3623);
nand U4423 (N_4423,N_3831,N_3243);
or U4424 (N_4424,N_3297,N_3362);
nand U4425 (N_4425,N_3927,N_3418);
or U4426 (N_4426,N_3645,N_3428);
and U4427 (N_4427,N_3505,N_3202);
or U4428 (N_4428,N_3153,N_3602);
nor U4429 (N_4429,N_3943,N_3156);
or U4430 (N_4430,N_3942,N_3615);
xnor U4431 (N_4431,N_3521,N_3375);
nor U4432 (N_4432,N_3440,N_3897);
and U4433 (N_4433,N_3708,N_3293);
nand U4434 (N_4434,N_3369,N_3691);
nand U4435 (N_4435,N_3128,N_3399);
xor U4436 (N_4436,N_3124,N_3069);
and U4437 (N_4437,N_3494,N_3723);
nand U4438 (N_4438,N_3786,N_3849);
nor U4439 (N_4439,N_3008,N_3700);
and U4440 (N_4440,N_3388,N_3338);
xor U4441 (N_4441,N_3584,N_3495);
xor U4442 (N_4442,N_3009,N_3761);
and U4443 (N_4443,N_3910,N_3714);
xor U4444 (N_4444,N_3538,N_3782);
nand U4445 (N_4445,N_3414,N_3784);
nor U4446 (N_4446,N_3183,N_3323);
and U4447 (N_4447,N_3754,N_3052);
xnor U4448 (N_4448,N_3366,N_3841);
xor U4449 (N_4449,N_3553,N_3903);
and U4450 (N_4450,N_3195,N_3727);
or U4451 (N_4451,N_3594,N_3644);
xor U4452 (N_4452,N_3778,N_3749);
xnor U4453 (N_4453,N_3286,N_3535);
and U4454 (N_4454,N_3249,N_3948);
nand U4455 (N_4455,N_3937,N_3973);
nand U4456 (N_4456,N_3772,N_3373);
xnor U4457 (N_4457,N_3641,N_3429);
nand U4458 (N_4458,N_3673,N_3686);
nand U4459 (N_4459,N_3481,N_3617);
nor U4460 (N_4460,N_3103,N_3391);
nor U4461 (N_4461,N_3651,N_3294);
or U4462 (N_4462,N_3980,N_3179);
xor U4463 (N_4463,N_3914,N_3235);
or U4464 (N_4464,N_3316,N_3800);
or U4465 (N_4465,N_3728,N_3442);
xnor U4466 (N_4466,N_3581,N_3173);
nor U4467 (N_4467,N_3774,N_3325);
nor U4468 (N_4468,N_3275,N_3150);
nor U4469 (N_4469,N_3747,N_3474);
and U4470 (N_4470,N_3984,N_3719);
and U4471 (N_4471,N_3490,N_3585);
nand U4472 (N_4472,N_3544,N_3805);
nor U4473 (N_4473,N_3867,N_3840);
and U4474 (N_4474,N_3949,N_3638);
xor U4475 (N_4475,N_3258,N_3703);
and U4476 (N_4476,N_3475,N_3498);
nand U4477 (N_4477,N_3461,N_3880);
or U4478 (N_4478,N_3022,N_3116);
or U4479 (N_4479,N_3364,N_3653);
xnor U4480 (N_4480,N_3028,N_3932);
nand U4481 (N_4481,N_3315,N_3809);
and U4482 (N_4482,N_3643,N_3302);
or U4483 (N_4483,N_3492,N_3380);
nor U4484 (N_4484,N_3397,N_3422);
xor U4485 (N_4485,N_3940,N_3447);
nor U4486 (N_4486,N_3512,N_3709);
and U4487 (N_4487,N_3689,N_3002);
and U4488 (N_4488,N_3983,N_3993);
nand U4489 (N_4489,N_3730,N_3061);
or U4490 (N_4490,N_3503,N_3655);
nand U4491 (N_4491,N_3226,N_3665);
nor U4492 (N_4492,N_3750,N_3792);
nor U4493 (N_4493,N_3667,N_3080);
nor U4494 (N_4494,N_3661,N_3671);
or U4495 (N_4495,N_3454,N_3207);
nand U4496 (N_4496,N_3530,N_3182);
and U4497 (N_4497,N_3918,N_3777);
xnor U4498 (N_4498,N_3141,N_3955);
or U4499 (N_4499,N_3663,N_3085);
and U4500 (N_4500,N_3093,N_3879);
or U4501 (N_4501,N_3976,N_3004);
nand U4502 (N_4502,N_3962,N_3499);
nor U4503 (N_4503,N_3006,N_3845);
or U4504 (N_4504,N_3390,N_3538);
xnor U4505 (N_4505,N_3569,N_3401);
nor U4506 (N_4506,N_3217,N_3931);
nor U4507 (N_4507,N_3176,N_3268);
and U4508 (N_4508,N_3573,N_3358);
nor U4509 (N_4509,N_3057,N_3895);
nand U4510 (N_4510,N_3328,N_3511);
or U4511 (N_4511,N_3285,N_3348);
xnor U4512 (N_4512,N_3331,N_3013);
xnor U4513 (N_4513,N_3509,N_3747);
xor U4514 (N_4514,N_3289,N_3863);
xor U4515 (N_4515,N_3013,N_3804);
or U4516 (N_4516,N_3687,N_3912);
nor U4517 (N_4517,N_3126,N_3631);
nor U4518 (N_4518,N_3559,N_3498);
xnor U4519 (N_4519,N_3889,N_3191);
xnor U4520 (N_4520,N_3001,N_3452);
and U4521 (N_4521,N_3641,N_3655);
xor U4522 (N_4522,N_3151,N_3759);
xor U4523 (N_4523,N_3585,N_3765);
and U4524 (N_4524,N_3328,N_3446);
nand U4525 (N_4525,N_3672,N_3580);
nand U4526 (N_4526,N_3884,N_3017);
or U4527 (N_4527,N_3994,N_3680);
nor U4528 (N_4528,N_3891,N_3840);
and U4529 (N_4529,N_3733,N_3244);
nand U4530 (N_4530,N_3741,N_3514);
xnor U4531 (N_4531,N_3443,N_3688);
xnor U4532 (N_4532,N_3857,N_3521);
and U4533 (N_4533,N_3277,N_3179);
nor U4534 (N_4534,N_3767,N_3208);
or U4535 (N_4535,N_3234,N_3602);
nor U4536 (N_4536,N_3780,N_3644);
xnor U4537 (N_4537,N_3244,N_3712);
and U4538 (N_4538,N_3662,N_3875);
or U4539 (N_4539,N_3033,N_3513);
xor U4540 (N_4540,N_3656,N_3711);
xnor U4541 (N_4541,N_3523,N_3746);
nor U4542 (N_4542,N_3493,N_3182);
xnor U4543 (N_4543,N_3906,N_3511);
nor U4544 (N_4544,N_3772,N_3698);
nand U4545 (N_4545,N_3521,N_3258);
or U4546 (N_4546,N_3389,N_3135);
or U4547 (N_4547,N_3423,N_3188);
nor U4548 (N_4548,N_3009,N_3624);
nor U4549 (N_4549,N_3983,N_3547);
and U4550 (N_4550,N_3693,N_3194);
xor U4551 (N_4551,N_3543,N_3035);
and U4552 (N_4552,N_3111,N_3025);
or U4553 (N_4553,N_3408,N_3724);
nand U4554 (N_4554,N_3745,N_3079);
nand U4555 (N_4555,N_3441,N_3084);
nand U4556 (N_4556,N_3833,N_3144);
nand U4557 (N_4557,N_3620,N_3039);
and U4558 (N_4558,N_3209,N_3983);
and U4559 (N_4559,N_3684,N_3573);
nand U4560 (N_4560,N_3304,N_3521);
nand U4561 (N_4561,N_3998,N_3792);
nand U4562 (N_4562,N_3221,N_3669);
or U4563 (N_4563,N_3598,N_3774);
xor U4564 (N_4564,N_3594,N_3398);
nand U4565 (N_4565,N_3604,N_3758);
or U4566 (N_4566,N_3808,N_3196);
and U4567 (N_4567,N_3322,N_3876);
or U4568 (N_4568,N_3253,N_3988);
or U4569 (N_4569,N_3661,N_3989);
xnor U4570 (N_4570,N_3680,N_3671);
or U4571 (N_4571,N_3527,N_3186);
or U4572 (N_4572,N_3649,N_3342);
or U4573 (N_4573,N_3782,N_3366);
xnor U4574 (N_4574,N_3480,N_3006);
or U4575 (N_4575,N_3237,N_3964);
nand U4576 (N_4576,N_3083,N_3981);
xor U4577 (N_4577,N_3228,N_3404);
xnor U4578 (N_4578,N_3531,N_3082);
nand U4579 (N_4579,N_3170,N_3366);
and U4580 (N_4580,N_3160,N_3461);
nand U4581 (N_4581,N_3542,N_3810);
and U4582 (N_4582,N_3089,N_3201);
or U4583 (N_4583,N_3622,N_3442);
nor U4584 (N_4584,N_3231,N_3872);
xor U4585 (N_4585,N_3999,N_3656);
and U4586 (N_4586,N_3572,N_3417);
xnor U4587 (N_4587,N_3211,N_3502);
and U4588 (N_4588,N_3638,N_3690);
xnor U4589 (N_4589,N_3541,N_3714);
xnor U4590 (N_4590,N_3128,N_3724);
xnor U4591 (N_4591,N_3689,N_3923);
and U4592 (N_4592,N_3606,N_3902);
nand U4593 (N_4593,N_3736,N_3902);
or U4594 (N_4594,N_3648,N_3149);
xnor U4595 (N_4595,N_3608,N_3953);
xor U4596 (N_4596,N_3688,N_3913);
xor U4597 (N_4597,N_3873,N_3262);
or U4598 (N_4598,N_3163,N_3879);
xor U4599 (N_4599,N_3115,N_3196);
and U4600 (N_4600,N_3514,N_3341);
and U4601 (N_4601,N_3032,N_3875);
nor U4602 (N_4602,N_3670,N_3971);
and U4603 (N_4603,N_3174,N_3195);
and U4604 (N_4604,N_3101,N_3723);
and U4605 (N_4605,N_3021,N_3600);
or U4606 (N_4606,N_3899,N_3024);
nor U4607 (N_4607,N_3554,N_3996);
nand U4608 (N_4608,N_3359,N_3048);
or U4609 (N_4609,N_3182,N_3729);
nor U4610 (N_4610,N_3544,N_3360);
or U4611 (N_4611,N_3313,N_3111);
nor U4612 (N_4612,N_3210,N_3025);
nor U4613 (N_4613,N_3620,N_3022);
nand U4614 (N_4614,N_3123,N_3047);
nand U4615 (N_4615,N_3543,N_3211);
nand U4616 (N_4616,N_3391,N_3957);
or U4617 (N_4617,N_3342,N_3544);
and U4618 (N_4618,N_3382,N_3876);
or U4619 (N_4619,N_3418,N_3662);
and U4620 (N_4620,N_3148,N_3276);
nor U4621 (N_4621,N_3128,N_3102);
nor U4622 (N_4622,N_3263,N_3853);
nand U4623 (N_4623,N_3046,N_3229);
and U4624 (N_4624,N_3985,N_3628);
or U4625 (N_4625,N_3163,N_3669);
and U4626 (N_4626,N_3362,N_3106);
and U4627 (N_4627,N_3588,N_3689);
xor U4628 (N_4628,N_3017,N_3853);
nand U4629 (N_4629,N_3017,N_3033);
xor U4630 (N_4630,N_3901,N_3636);
xnor U4631 (N_4631,N_3752,N_3254);
nand U4632 (N_4632,N_3860,N_3913);
or U4633 (N_4633,N_3514,N_3455);
or U4634 (N_4634,N_3360,N_3827);
xnor U4635 (N_4635,N_3845,N_3039);
nor U4636 (N_4636,N_3807,N_3794);
or U4637 (N_4637,N_3394,N_3830);
nor U4638 (N_4638,N_3052,N_3912);
or U4639 (N_4639,N_3669,N_3953);
or U4640 (N_4640,N_3727,N_3938);
and U4641 (N_4641,N_3707,N_3890);
and U4642 (N_4642,N_3760,N_3159);
xnor U4643 (N_4643,N_3197,N_3387);
nor U4644 (N_4644,N_3129,N_3289);
nor U4645 (N_4645,N_3320,N_3101);
nand U4646 (N_4646,N_3992,N_3668);
nor U4647 (N_4647,N_3144,N_3272);
xor U4648 (N_4648,N_3723,N_3027);
nand U4649 (N_4649,N_3397,N_3030);
xor U4650 (N_4650,N_3210,N_3330);
and U4651 (N_4651,N_3172,N_3779);
nand U4652 (N_4652,N_3843,N_3341);
nand U4653 (N_4653,N_3423,N_3826);
or U4654 (N_4654,N_3266,N_3952);
nand U4655 (N_4655,N_3517,N_3100);
nand U4656 (N_4656,N_3231,N_3458);
and U4657 (N_4657,N_3935,N_3047);
nand U4658 (N_4658,N_3975,N_3986);
nor U4659 (N_4659,N_3410,N_3770);
nand U4660 (N_4660,N_3133,N_3382);
or U4661 (N_4661,N_3805,N_3317);
nor U4662 (N_4662,N_3688,N_3222);
and U4663 (N_4663,N_3969,N_3428);
xnor U4664 (N_4664,N_3199,N_3143);
and U4665 (N_4665,N_3362,N_3726);
nand U4666 (N_4666,N_3141,N_3864);
xor U4667 (N_4667,N_3974,N_3432);
nor U4668 (N_4668,N_3156,N_3454);
and U4669 (N_4669,N_3035,N_3447);
or U4670 (N_4670,N_3905,N_3153);
or U4671 (N_4671,N_3146,N_3314);
or U4672 (N_4672,N_3725,N_3812);
or U4673 (N_4673,N_3006,N_3625);
or U4674 (N_4674,N_3703,N_3284);
or U4675 (N_4675,N_3021,N_3618);
nand U4676 (N_4676,N_3482,N_3796);
nor U4677 (N_4677,N_3538,N_3213);
nand U4678 (N_4678,N_3086,N_3451);
nor U4679 (N_4679,N_3387,N_3900);
and U4680 (N_4680,N_3001,N_3262);
nand U4681 (N_4681,N_3950,N_3553);
and U4682 (N_4682,N_3893,N_3135);
or U4683 (N_4683,N_3536,N_3563);
and U4684 (N_4684,N_3513,N_3269);
and U4685 (N_4685,N_3679,N_3267);
or U4686 (N_4686,N_3317,N_3848);
and U4687 (N_4687,N_3894,N_3779);
or U4688 (N_4688,N_3322,N_3644);
nand U4689 (N_4689,N_3130,N_3356);
xnor U4690 (N_4690,N_3507,N_3657);
xnor U4691 (N_4691,N_3595,N_3652);
nand U4692 (N_4692,N_3285,N_3471);
nor U4693 (N_4693,N_3301,N_3691);
nor U4694 (N_4694,N_3780,N_3649);
xor U4695 (N_4695,N_3151,N_3640);
and U4696 (N_4696,N_3326,N_3769);
xnor U4697 (N_4697,N_3087,N_3540);
and U4698 (N_4698,N_3370,N_3604);
xnor U4699 (N_4699,N_3193,N_3761);
or U4700 (N_4700,N_3070,N_3329);
xnor U4701 (N_4701,N_3394,N_3931);
nor U4702 (N_4702,N_3632,N_3659);
or U4703 (N_4703,N_3494,N_3842);
or U4704 (N_4704,N_3639,N_3010);
xnor U4705 (N_4705,N_3910,N_3595);
nand U4706 (N_4706,N_3507,N_3449);
and U4707 (N_4707,N_3230,N_3449);
xnor U4708 (N_4708,N_3119,N_3631);
nand U4709 (N_4709,N_3958,N_3629);
and U4710 (N_4710,N_3036,N_3430);
or U4711 (N_4711,N_3392,N_3329);
or U4712 (N_4712,N_3397,N_3448);
and U4713 (N_4713,N_3334,N_3045);
xor U4714 (N_4714,N_3147,N_3585);
nor U4715 (N_4715,N_3037,N_3755);
nor U4716 (N_4716,N_3370,N_3207);
nand U4717 (N_4717,N_3639,N_3634);
xnor U4718 (N_4718,N_3417,N_3253);
xor U4719 (N_4719,N_3894,N_3935);
xor U4720 (N_4720,N_3051,N_3513);
xor U4721 (N_4721,N_3413,N_3245);
or U4722 (N_4722,N_3632,N_3821);
and U4723 (N_4723,N_3100,N_3924);
nand U4724 (N_4724,N_3595,N_3752);
and U4725 (N_4725,N_3853,N_3083);
nand U4726 (N_4726,N_3910,N_3354);
xnor U4727 (N_4727,N_3343,N_3368);
xor U4728 (N_4728,N_3358,N_3825);
xnor U4729 (N_4729,N_3534,N_3959);
or U4730 (N_4730,N_3438,N_3172);
nor U4731 (N_4731,N_3268,N_3278);
or U4732 (N_4732,N_3026,N_3356);
xnor U4733 (N_4733,N_3495,N_3151);
xor U4734 (N_4734,N_3987,N_3317);
nand U4735 (N_4735,N_3253,N_3736);
xnor U4736 (N_4736,N_3653,N_3880);
nand U4737 (N_4737,N_3018,N_3710);
nor U4738 (N_4738,N_3724,N_3469);
or U4739 (N_4739,N_3910,N_3639);
nor U4740 (N_4740,N_3877,N_3568);
and U4741 (N_4741,N_3874,N_3805);
and U4742 (N_4742,N_3672,N_3186);
and U4743 (N_4743,N_3025,N_3262);
nand U4744 (N_4744,N_3701,N_3425);
or U4745 (N_4745,N_3471,N_3927);
and U4746 (N_4746,N_3926,N_3129);
or U4747 (N_4747,N_3931,N_3174);
xnor U4748 (N_4748,N_3340,N_3562);
or U4749 (N_4749,N_3106,N_3285);
xor U4750 (N_4750,N_3039,N_3881);
or U4751 (N_4751,N_3876,N_3375);
or U4752 (N_4752,N_3501,N_3645);
nand U4753 (N_4753,N_3949,N_3916);
xor U4754 (N_4754,N_3177,N_3603);
xor U4755 (N_4755,N_3331,N_3189);
and U4756 (N_4756,N_3076,N_3084);
xor U4757 (N_4757,N_3797,N_3092);
nand U4758 (N_4758,N_3001,N_3623);
and U4759 (N_4759,N_3872,N_3736);
or U4760 (N_4760,N_3826,N_3521);
nor U4761 (N_4761,N_3158,N_3972);
and U4762 (N_4762,N_3474,N_3092);
and U4763 (N_4763,N_3561,N_3719);
or U4764 (N_4764,N_3665,N_3394);
and U4765 (N_4765,N_3152,N_3738);
xnor U4766 (N_4766,N_3685,N_3182);
nor U4767 (N_4767,N_3777,N_3835);
and U4768 (N_4768,N_3605,N_3434);
xnor U4769 (N_4769,N_3795,N_3635);
nor U4770 (N_4770,N_3594,N_3956);
nor U4771 (N_4771,N_3511,N_3135);
or U4772 (N_4772,N_3879,N_3177);
and U4773 (N_4773,N_3274,N_3596);
nor U4774 (N_4774,N_3647,N_3127);
xnor U4775 (N_4775,N_3563,N_3358);
xnor U4776 (N_4776,N_3400,N_3959);
xor U4777 (N_4777,N_3078,N_3485);
xnor U4778 (N_4778,N_3761,N_3961);
nand U4779 (N_4779,N_3899,N_3948);
nand U4780 (N_4780,N_3952,N_3104);
nor U4781 (N_4781,N_3457,N_3315);
nor U4782 (N_4782,N_3324,N_3786);
nand U4783 (N_4783,N_3067,N_3781);
xnor U4784 (N_4784,N_3160,N_3412);
xnor U4785 (N_4785,N_3876,N_3098);
xor U4786 (N_4786,N_3777,N_3644);
nand U4787 (N_4787,N_3327,N_3756);
xor U4788 (N_4788,N_3366,N_3837);
nand U4789 (N_4789,N_3844,N_3074);
xnor U4790 (N_4790,N_3571,N_3869);
and U4791 (N_4791,N_3289,N_3758);
or U4792 (N_4792,N_3747,N_3052);
nand U4793 (N_4793,N_3626,N_3943);
and U4794 (N_4794,N_3249,N_3593);
nand U4795 (N_4795,N_3374,N_3545);
or U4796 (N_4796,N_3171,N_3282);
xnor U4797 (N_4797,N_3478,N_3473);
nor U4798 (N_4798,N_3628,N_3854);
nand U4799 (N_4799,N_3624,N_3836);
nand U4800 (N_4800,N_3170,N_3823);
and U4801 (N_4801,N_3837,N_3526);
or U4802 (N_4802,N_3107,N_3357);
and U4803 (N_4803,N_3694,N_3354);
and U4804 (N_4804,N_3216,N_3471);
xnor U4805 (N_4805,N_3756,N_3295);
nor U4806 (N_4806,N_3046,N_3235);
nor U4807 (N_4807,N_3798,N_3715);
nor U4808 (N_4808,N_3299,N_3108);
and U4809 (N_4809,N_3477,N_3100);
xnor U4810 (N_4810,N_3104,N_3655);
or U4811 (N_4811,N_3418,N_3305);
nand U4812 (N_4812,N_3407,N_3397);
and U4813 (N_4813,N_3921,N_3654);
or U4814 (N_4814,N_3082,N_3563);
nor U4815 (N_4815,N_3378,N_3659);
xnor U4816 (N_4816,N_3128,N_3470);
and U4817 (N_4817,N_3623,N_3657);
and U4818 (N_4818,N_3587,N_3264);
nor U4819 (N_4819,N_3784,N_3940);
or U4820 (N_4820,N_3607,N_3615);
or U4821 (N_4821,N_3628,N_3601);
and U4822 (N_4822,N_3676,N_3721);
nor U4823 (N_4823,N_3531,N_3968);
nand U4824 (N_4824,N_3911,N_3293);
xor U4825 (N_4825,N_3818,N_3786);
nand U4826 (N_4826,N_3142,N_3939);
nor U4827 (N_4827,N_3783,N_3891);
nor U4828 (N_4828,N_3302,N_3594);
and U4829 (N_4829,N_3753,N_3088);
xnor U4830 (N_4830,N_3192,N_3911);
nor U4831 (N_4831,N_3477,N_3545);
or U4832 (N_4832,N_3249,N_3175);
or U4833 (N_4833,N_3833,N_3717);
and U4834 (N_4834,N_3867,N_3008);
and U4835 (N_4835,N_3361,N_3823);
nand U4836 (N_4836,N_3657,N_3784);
nor U4837 (N_4837,N_3602,N_3654);
nand U4838 (N_4838,N_3291,N_3677);
nor U4839 (N_4839,N_3892,N_3268);
nor U4840 (N_4840,N_3042,N_3153);
or U4841 (N_4841,N_3275,N_3349);
xor U4842 (N_4842,N_3984,N_3581);
xor U4843 (N_4843,N_3316,N_3255);
xor U4844 (N_4844,N_3896,N_3779);
xor U4845 (N_4845,N_3612,N_3795);
nor U4846 (N_4846,N_3443,N_3418);
and U4847 (N_4847,N_3582,N_3050);
xnor U4848 (N_4848,N_3070,N_3782);
or U4849 (N_4849,N_3551,N_3165);
nand U4850 (N_4850,N_3321,N_3022);
nand U4851 (N_4851,N_3287,N_3068);
and U4852 (N_4852,N_3809,N_3721);
nor U4853 (N_4853,N_3750,N_3335);
or U4854 (N_4854,N_3360,N_3343);
nor U4855 (N_4855,N_3147,N_3636);
and U4856 (N_4856,N_3991,N_3366);
nor U4857 (N_4857,N_3537,N_3180);
and U4858 (N_4858,N_3164,N_3948);
or U4859 (N_4859,N_3435,N_3993);
nor U4860 (N_4860,N_3274,N_3976);
nand U4861 (N_4861,N_3976,N_3455);
nor U4862 (N_4862,N_3148,N_3633);
nor U4863 (N_4863,N_3735,N_3986);
or U4864 (N_4864,N_3267,N_3047);
nor U4865 (N_4865,N_3131,N_3362);
nand U4866 (N_4866,N_3747,N_3126);
or U4867 (N_4867,N_3375,N_3315);
or U4868 (N_4868,N_3004,N_3297);
xor U4869 (N_4869,N_3490,N_3745);
and U4870 (N_4870,N_3169,N_3740);
nand U4871 (N_4871,N_3118,N_3980);
nor U4872 (N_4872,N_3581,N_3987);
xnor U4873 (N_4873,N_3786,N_3889);
xor U4874 (N_4874,N_3761,N_3401);
nor U4875 (N_4875,N_3349,N_3558);
and U4876 (N_4876,N_3854,N_3698);
nand U4877 (N_4877,N_3294,N_3395);
or U4878 (N_4878,N_3899,N_3961);
or U4879 (N_4879,N_3421,N_3781);
nor U4880 (N_4880,N_3579,N_3285);
or U4881 (N_4881,N_3116,N_3893);
xor U4882 (N_4882,N_3507,N_3684);
or U4883 (N_4883,N_3192,N_3279);
xor U4884 (N_4884,N_3190,N_3964);
nand U4885 (N_4885,N_3601,N_3541);
or U4886 (N_4886,N_3161,N_3785);
nand U4887 (N_4887,N_3877,N_3510);
or U4888 (N_4888,N_3373,N_3811);
xor U4889 (N_4889,N_3287,N_3396);
or U4890 (N_4890,N_3530,N_3107);
or U4891 (N_4891,N_3096,N_3622);
nor U4892 (N_4892,N_3462,N_3082);
and U4893 (N_4893,N_3717,N_3620);
and U4894 (N_4894,N_3978,N_3337);
nand U4895 (N_4895,N_3763,N_3266);
or U4896 (N_4896,N_3772,N_3661);
or U4897 (N_4897,N_3042,N_3457);
nand U4898 (N_4898,N_3328,N_3774);
and U4899 (N_4899,N_3198,N_3694);
or U4900 (N_4900,N_3212,N_3898);
nor U4901 (N_4901,N_3170,N_3948);
nor U4902 (N_4902,N_3107,N_3490);
nor U4903 (N_4903,N_3926,N_3621);
and U4904 (N_4904,N_3033,N_3368);
nand U4905 (N_4905,N_3542,N_3694);
and U4906 (N_4906,N_3684,N_3026);
nand U4907 (N_4907,N_3864,N_3067);
and U4908 (N_4908,N_3146,N_3379);
nor U4909 (N_4909,N_3316,N_3390);
or U4910 (N_4910,N_3861,N_3891);
nand U4911 (N_4911,N_3199,N_3694);
xor U4912 (N_4912,N_3357,N_3205);
and U4913 (N_4913,N_3928,N_3408);
and U4914 (N_4914,N_3229,N_3584);
xor U4915 (N_4915,N_3466,N_3545);
nor U4916 (N_4916,N_3680,N_3546);
xor U4917 (N_4917,N_3025,N_3993);
or U4918 (N_4918,N_3395,N_3662);
and U4919 (N_4919,N_3929,N_3544);
xor U4920 (N_4920,N_3687,N_3017);
and U4921 (N_4921,N_3654,N_3186);
xnor U4922 (N_4922,N_3837,N_3905);
and U4923 (N_4923,N_3949,N_3287);
or U4924 (N_4924,N_3739,N_3094);
nor U4925 (N_4925,N_3425,N_3179);
nand U4926 (N_4926,N_3804,N_3521);
xor U4927 (N_4927,N_3797,N_3789);
xnor U4928 (N_4928,N_3084,N_3712);
and U4929 (N_4929,N_3589,N_3070);
xnor U4930 (N_4930,N_3396,N_3719);
nor U4931 (N_4931,N_3468,N_3097);
nor U4932 (N_4932,N_3723,N_3100);
and U4933 (N_4933,N_3649,N_3077);
xnor U4934 (N_4934,N_3851,N_3516);
nor U4935 (N_4935,N_3866,N_3672);
nand U4936 (N_4936,N_3015,N_3747);
and U4937 (N_4937,N_3720,N_3980);
nor U4938 (N_4938,N_3645,N_3142);
nor U4939 (N_4939,N_3488,N_3375);
or U4940 (N_4940,N_3933,N_3988);
nor U4941 (N_4941,N_3202,N_3341);
nor U4942 (N_4942,N_3011,N_3338);
xnor U4943 (N_4943,N_3036,N_3707);
and U4944 (N_4944,N_3556,N_3589);
nor U4945 (N_4945,N_3394,N_3579);
or U4946 (N_4946,N_3356,N_3005);
nor U4947 (N_4947,N_3011,N_3695);
nor U4948 (N_4948,N_3213,N_3253);
xor U4949 (N_4949,N_3690,N_3518);
nand U4950 (N_4950,N_3409,N_3060);
and U4951 (N_4951,N_3300,N_3485);
nor U4952 (N_4952,N_3206,N_3602);
xor U4953 (N_4953,N_3356,N_3717);
or U4954 (N_4954,N_3247,N_3983);
or U4955 (N_4955,N_3581,N_3073);
xnor U4956 (N_4956,N_3109,N_3431);
nand U4957 (N_4957,N_3372,N_3035);
or U4958 (N_4958,N_3035,N_3647);
nor U4959 (N_4959,N_3656,N_3148);
xor U4960 (N_4960,N_3356,N_3669);
nor U4961 (N_4961,N_3489,N_3348);
nand U4962 (N_4962,N_3796,N_3071);
or U4963 (N_4963,N_3594,N_3722);
or U4964 (N_4964,N_3002,N_3886);
or U4965 (N_4965,N_3311,N_3719);
nor U4966 (N_4966,N_3190,N_3655);
nand U4967 (N_4967,N_3576,N_3687);
nor U4968 (N_4968,N_3338,N_3534);
nor U4969 (N_4969,N_3570,N_3016);
nor U4970 (N_4970,N_3092,N_3352);
or U4971 (N_4971,N_3343,N_3191);
xor U4972 (N_4972,N_3967,N_3666);
nand U4973 (N_4973,N_3922,N_3946);
nand U4974 (N_4974,N_3612,N_3265);
nand U4975 (N_4975,N_3426,N_3393);
or U4976 (N_4976,N_3080,N_3388);
or U4977 (N_4977,N_3383,N_3505);
and U4978 (N_4978,N_3010,N_3376);
and U4979 (N_4979,N_3774,N_3687);
xor U4980 (N_4980,N_3852,N_3749);
xnor U4981 (N_4981,N_3711,N_3125);
nor U4982 (N_4982,N_3147,N_3285);
or U4983 (N_4983,N_3289,N_3566);
nor U4984 (N_4984,N_3346,N_3126);
or U4985 (N_4985,N_3114,N_3838);
xnor U4986 (N_4986,N_3528,N_3179);
nand U4987 (N_4987,N_3661,N_3397);
xnor U4988 (N_4988,N_3606,N_3358);
nor U4989 (N_4989,N_3288,N_3595);
nand U4990 (N_4990,N_3002,N_3519);
xnor U4991 (N_4991,N_3934,N_3390);
nand U4992 (N_4992,N_3947,N_3704);
and U4993 (N_4993,N_3704,N_3625);
nand U4994 (N_4994,N_3482,N_3437);
and U4995 (N_4995,N_3296,N_3288);
and U4996 (N_4996,N_3336,N_3080);
xor U4997 (N_4997,N_3281,N_3790);
or U4998 (N_4998,N_3717,N_3681);
xnor U4999 (N_4999,N_3501,N_3199);
or U5000 (N_5000,N_4219,N_4624);
nor U5001 (N_5001,N_4930,N_4365);
xor U5002 (N_5002,N_4266,N_4943);
nand U5003 (N_5003,N_4837,N_4575);
nor U5004 (N_5004,N_4671,N_4673);
and U5005 (N_5005,N_4042,N_4648);
nor U5006 (N_5006,N_4689,N_4633);
xnor U5007 (N_5007,N_4013,N_4323);
xor U5008 (N_5008,N_4600,N_4109);
nor U5009 (N_5009,N_4532,N_4435);
nand U5010 (N_5010,N_4080,N_4324);
nor U5011 (N_5011,N_4628,N_4970);
or U5012 (N_5012,N_4393,N_4209);
or U5013 (N_5013,N_4657,N_4142);
xor U5014 (N_5014,N_4057,N_4150);
nand U5015 (N_5015,N_4264,N_4986);
or U5016 (N_5016,N_4619,N_4678);
nor U5017 (N_5017,N_4661,N_4862);
nand U5018 (N_5018,N_4108,N_4818);
nand U5019 (N_5019,N_4426,N_4474);
nor U5020 (N_5020,N_4516,N_4065);
and U5021 (N_5021,N_4071,N_4213);
nand U5022 (N_5022,N_4895,N_4867);
xnor U5023 (N_5023,N_4552,N_4766);
nor U5024 (N_5024,N_4345,N_4546);
or U5025 (N_5025,N_4521,N_4461);
nor U5026 (N_5026,N_4642,N_4423);
xor U5027 (N_5027,N_4060,N_4896);
or U5028 (N_5028,N_4023,N_4127);
xnor U5029 (N_5029,N_4699,N_4351);
xnor U5030 (N_5030,N_4291,N_4471);
xor U5031 (N_5031,N_4972,N_4541);
and U5032 (N_5032,N_4355,N_4932);
nor U5033 (N_5033,N_4710,N_4669);
and U5034 (N_5034,N_4145,N_4372);
nor U5035 (N_5035,N_4430,N_4200);
xnor U5036 (N_5036,N_4156,N_4558);
or U5037 (N_5037,N_4909,N_4014);
or U5038 (N_5038,N_4233,N_4173);
xnor U5039 (N_5039,N_4043,N_4976);
xor U5040 (N_5040,N_4413,N_4242);
or U5041 (N_5041,N_4252,N_4543);
nand U5042 (N_5042,N_4592,N_4416);
and U5043 (N_5043,N_4696,N_4090);
and U5044 (N_5044,N_4447,N_4135);
and U5045 (N_5045,N_4215,N_4906);
nor U5046 (N_5046,N_4692,N_4808);
nor U5047 (N_5047,N_4882,N_4410);
nor U5048 (N_5048,N_4202,N_4183);
xnor U5049 (N_5049,N_4525,N_4615);
nor U5050 (N_5050,N_4500,N_4185);
xnor U5051 (N_5051,N_4220,N_4973);
nor U5052 (N_5052,N_4695,N_4064);
nor U5053 (N_5053,N_4576,N_4686);
nor U5054 (N_5054,N_4153,N_4462);
nand U5055 (N_5055,N_4371,N_4807);
and U5056 (N_5056,N_4451,N_4594);
or U5057 (N_5057,N_4983,N_4006);
nor U5058 (N_5058,N_4907,N_4046);
and U5059 (N_5059,N_4805,N_4399);
nor U5060 (N_5060,N_4578,N_4879);
xor U5061 (N_5061,N_4282,N_4095);
or U5062 (N_5062,N_4781,N_4102);
xnor U5063 (N_5063,N_4596,N_4729);
nor U5064 (N_5064,N_4515,N_4453);
nor U5065 (N_5065,N_4000,N_4314);
nand U5066 (N_5066,N_4420,N_4921);
xor U5067 (N_5067,N_4431,N_4201);
and U5068 (N_5068,N_4313,N_4418);
or U5069 (N_5069,N_4049,N_4853);
nor U5070 (N_5070,N_4364,N_4203);
xnor U5071 (N_5071,N_4773,N_4969);
nand U5072 (N_5072,N_4368,N_4101);
and U5073 (N_5073,N_4865,N_4590);
and U5074 (N_5074,N_4362,N_4743);
or U5075 (N_5075,N_4849,N_4616);
and U5076 (N_5076,N_4405,N_4744);
or U5077 (N_5077,N_4772,N_4106);
xnor U5078 (N_5078,N_4555,N_4164);
xnor U5079 (N_5079,N_4407,N_4995);
nor U5080 (N_5080,N_4840,N_4711);
and U5081 (N_5081,N_4666,N_4414);
nor U5082 (N_5082,N_4093,N_4366);
and U5083 (N_5083,N_4980,N_4519);
or U5084 (N_5084,N_4148,N_4409);
xnor U5085 (N_5085,N_4572,N_4786);
xnor U5086 (N_5086,N_4884,N_4449);
and U5087 (N_5087,N_4293,N_4512);
or U5088 (N_5088,N_4297,N_4813);
xor U5089 (N_5089,N_4990,N_4800);
xor U5090 (N_5090,N_4175,N_4994);
and U5091 (N_5091,N_4222,N_4883);
xnor U5092 (N_5092,N_4854,N_4070);
xor U5093 (N_5093,N_4121,N_4470);
or U5094 (N_5094,N_4803,N_4299);
and U5095 (N_5095,N_4408,N_4583);
nand U5096 (N_5096,N_4656,N_4212);
and U5097 (N_5097,N_4147,N_4269);
nor U5098 (N_5098,N_4776,N_4801);
or U5099 (N_5099,N_4246,N_4499);
or U5100 (N_5100,N_4775,N_4460);
and U5101 (N_5101,N_4636,N_4629);
xor U5102 (N_5102,N_4580,N_4835);
and U5103 (N_5103,N_4099,N_4702);
xor U5104 (N_5104,N_4251,N_4625);
and U5105 (N_5105,N_4253,N_4912);
nand U5106 (N_5106,N_4663,N_4454);
and U5107 (N_5107,N_4132,N_4476);
nor U5108 (N_5108,N_4588,N_4640);
nor U5109 (N_5109,N_4411,N_4363);
xor U5110 (N_5110,N_4717,N_4306);
and U5111 (N_5111,N_4257,N_4350);
or U5112 (N_5112,N_4340,N_4472);
and U5113 (N_5113,N_4505,N_4634);
xnor U5114 (N_5114,N_4789,N_4312);
nor U5115 (N_5115,N_4141,N_4063);
nor U5116 (N_5116,N_4052,N_4216);
nand U5117 (N_5117,N_4679,N_4281);
and U5118 (N_5118,N_4439,N_4359);
nor U5119 (N_5119,N_4685,N_4910);
xnor U5120 (N_5120,N_4484,N_4154);
or U5121 (N_5121,N_4001,N_4780);
nand U5122 (N_5122,N_4166,N_4022);
and U5123 (N_5123,N_4582,N_4181);
xnor U5124 (N_5124,N_4114,N_4611);
nand U5125 (N_5125,N_4701,N_4440);
nor U5126 (N_5126,N_4931,N_4660);
or U5127 (N_5127,N_4169,N_4851);
and U5128 (N_5128,N_4329,N_4612);
xor U5129 (N_5129,N_4131,N_4914);
nor U5130 (N_5130,N_4097,N_4311);
nand U5131 (N_5131,N_4991,N_4877);
xor U5132 (N_5132,N_4817,N_4079);
xor U5133 (N_5133,N_4709,N_4279);
and U5134 (N_5134,N_4791,N_4922);
xnor U5135 (N_5135,N_4855,N_4341);
and U5136 (N_5136,N_4740,N_4742);
nor U5137 (N_5137,N_4116,N_4165);
and U5138 (N_5138,N_4122,N_4802);
or U5139 (N_5139,N_4028,N_4275);
nand U5140 (N_5140,N_4231,N_4417);
xnor U5141 (N_5141,N_4876,N_4868);
nor U5142 (N_5142,N_4002,N_4824);
nand U5143 (N_5143,N_4003,N_4218);
nand U5144 (N_5144,N_4814,N_4077);
and U5145 (N_5145,N_4190,N_4607);
or U5146 (N_5146,N_4186,N_4204);
nand U5147 (N_5147,N_4459,N_4872);
nor U5148 (N_5148,N_4008,N_4873);
and U5149 (N_5149,N_4658,N_4852);
nor U5150 (N_5150,N_4794,N_4874);
or U5151 (N_5151,N_4292,N_4045);
nor U5152 (N_5152,N_4133,N_4513);
nand U5153 (N_5153,N_4386,N_4745);
nand U5154 (N_5154,N_4750,N_4728);
nand U5155 (N_5155,N_4507,N_4488);
nor U5156 (N_5156,N_4009,N_4026);
xnor U5157 (N_5157,N_4285,N_4730);
and U5158 (N_5158,N_4480,N_4086);
xor U5159 (N_5159,N_4665,N_4827);
nor U5160 (N_5160,N_4346,N_4396);
xor U5161 (N_5161,N_4024,N_4354);
nor U5162 (N_5162,N_4848,N_4347);
and U5163 (N_5163,N_4920,N_4146);
nor U5164 (N_5164,N_4739,N_4162);
and U5165 (N_5165,N_4105,N_4455);
xnor U5166 (N_5166,N_4258,N_4975);
and U5167 (N_5167,N_4191,N_4627);
and U5168 (N_5168,N_4170,N_4782);
or U5169 (N_5169,N_4958,N_4468);
xor U5170 (N_5170,N_4406,N_4645);
xnor U5171 (N_5171,N_4337,N_4621);
xor U5172 (N_5172,N_4381,N_4494);
or U5173 (N_5173,N_4760,N_4763);
nor U5174 (N_5174,N_4305,N_4288);
xor U5175 (N_5175,N_4569,N_4514);
xor U5176 (N_5176,N_4167,N_4704);
xor U5177 (N_5177,N_4981,N_4893);
xor U5178 (N_5178,N_4298,N_4676);
or U5179 (N_5179,N_4603,N_4984);
and U5180 (N_5180,N_4614,N_4107);
xor U5181 (N_5181,N_4935,N_4599);
nand U5182 (N_5182,N_4924,N_4965);
and U5183 (N_5183,N_4059,N_4038);
or U5184 (N_5184,N_4755,N_4604);
or U5185 (N_5185,N_4448,N_4927);
or U5186 (N_5186,N_4098,N_4517);
xnor U5187 (N_5187,N_4208,N_4498);
nor U5188 (N_5188,N_4529,N_4887);
nand U5189 (N_5189,N_4027,N_4320);
xnor U5190 (N_5190,N_4839,N_4947);
nor U5191 (N_5191,N_4829,N_4240);
and U5192 (N_5192,N_4248,N_4892);
or U5193 (N_5193,N_4978,N_4798);
nand U5194 (N_5194,N_4348,N_4094);
nand U5195 (N_5195,N_4904,N_4749);
or U5196 (N_5196,N_4992,N_4318);
or U5197 (N_5197,N_4081,N_4733);
xnor U5198 (N_5198,N_4178,N_4536);
or U5199 (N_5199,N_4662,N_4387);
xor U5200 (N_5200,N_4369,N_4769);
nor U5201 (N_5201,N_4759,N_4207);
nand U5202 (N_5202,N_4712,N_4724);
or U5203 (N_5203,N_4327,N_4950);
xor U5204 (N_5204,N_4068,N_4029);
and U5205 (N_5205,N_4570,N_4194);
nor U5206 (N_5206,N_4937,N_4300);
and U5207 (N_5207,N_4056,N_4916);
nand U5208 (N_5208,N_4971,N_4585);
and U5209 (N_5209,N_4509,N_4356);
and U5210 (N_5210,N_4360,N_4989);
xnor U5211 (N_5211,N_4573,N_4092);
or U5212 (N_5212,N_4339,N_4804);
xnor U5213 (N_5213,N_4442,N_4457);
xnor U5214 (N_5214,N_4124,N_4280);
or U5215 (N_5215,N_4402,N_4948);
nor U5216 (N_5216,N_4568,N_4718);
nand U5217 (N_5217,N_4650,N_4998);
nand U5218 (N_5218,N_4310,N_4574);
nand U5219 (N_5219,N_4774,N_4177);
or U5220 (N_5220,N_4062,N_4979);
nor U5221 (N_5221,N_4796,N_4731);
xor U5222 (N_5222,N_4319,N_4041);
xor U5223 (N_5223,N_4174,N_4664);
and U5224 (N_5224,N_4938,N_4700);
or U5225 (N_5225,N_4822,N_4171);
or U5226 (N_5226,N_4021,N_4490);
or U5227 (N_5227,N_4908,N_4234);
nor U5228 (N_5228,N_4672,N_4273);
or U5229 (N_5229,N_4858,N_4450);
or U5230 (N_5230,N_4284,N_4394);
or U5231 (N_5231,N_4495,N_4259);
or U5232 (N_5232,N_4296,N_4256);
or U5233 (N_5233,N_4261,N_4790);
xor U5234 (N_5234,N_4968,N_4559);
and U5235 (N_5235,N_4843,N_4952);
nor U5236 (N_5236,N_4271,N_4881);
nand U5237 (N_5237,N_4556,N_4757);
nand U5238 (N_5238,N_4765,N_4206);
xnor U5239 (N_5239,N_4746,N_4143);
nand U5240 (N_5240,N_4577,N_4267);
or U5241 (N_5241,N_4693,N_4084);
nand U5242 (N_5242,N_4539,N_4254);
xnor U5243 (N_5243,N_4214,N_4016);
xnor U5244 (N_5244,N_4630,N_4358);
and U5245 (N_5245,N_4917,N_4834);
and U5246 (N_5246,N_4388,N_4900);
nor U5247 (N_5247,N_4694,N_4492);
nor U5248 (N_5248,N_4561,N_4025);
and U5249 (N_5249,N_4184,N_4437);
nand U5250 (N_5250,N_4378,N_4089);
nor U5251 (N_5251,N_4199,N_4033);
nand U5252 (N_5252,N_4597,N_4939);
xor U5253 (N_5253,N_4223,N_4620);
nand U5254 (N_5254,N_4503,N_4523);
xnor U5255 (N_5255,N_4788,N_4385);
nor U5256 (N_5256,N_4117,N_4333);
xnor U5257 (N_5257,N_4287,N_4936);
xnor U5258 (N_5258,N_4168,N_4828);
xnor U5259 (N_5259,N_4289,N_4129);
and U5260 (N_5260,N_4428,N_4703);
or U5261 (N_5261,N_4493,N_4155);
or U5262 (N_5262,N_4825,N_4510);
nand U5263 (N_5263,N_4641,N_4545);
or U5264 (N_5264,N_4205,N_4705);
xnor U5265 (N_5265,N_4265,N_4250);
and U5266 (N_5266,N_4652,N_4623);
xor U5267 (N_5267,N_4608,N_4244);
or U5268 (N_5268,N_4771,N_4885);
or U5269 (N_5269,N_4085,N_4770);
nor U5270 (N_5270,N_4617,N_4110);
nor U5271 (N_5271,N_4096,N_4235);
xnor U5272 (N_5272,N_4964,N_4192);
nor U5273 (N_5273,N_4751,N_4263);
nor U5274 (N_5274,N_4847,N_4557);
or U5275 (N_5275,N_4030,N_4508);
nor U5276 (N_5276,N_4675,N_4959);
xor U5277 (N_5277,N_4072,N_4415);
xnor U5278 (N_5278,N_4015,N_4502);
xnor U5279 (N_5279,N_4714,N_4036);
nor U5280 (N_5280,N_4421,N_4832);
nor U5281 (N_5281,N_4799,N_4436);
nand U5282 (N_5282,N_4842,N_4878);
xnor U5283 (N_5283,N_4304,N_4584);
and U5284 (N_5284,N_4732,N_4768);
or U5285 (N_5285,N_4547,N_4446);
or U5286 (N_5286,N_4844,N_4520);
xnor U5287 (N_5287,N_4422,N_4397);
nand U5288 (N_5288,N_4687,N_4725);
or U5289 (N_5289,N_4441,N_4463);
xnor U5290 (N_5290,N_4152,N_4815);
nor U5291 (N_5291,N_4158,N_4126);
and U5292 (N_5292,N_4334,N_4587);
xnor U5293 (N_5293,N_4087,N_4445);
and U5294 (N_5294,N_4831,N_4290);
or U5295 (N_5295,N_4535,N_4074);
nand U5296 (N_5296,N_4227,N_4073);
or U5297 (N_5297,N_4295,N_4553);
or U5298 (N_5298,N_4343,N_4485);
nor U5299 (N_5299,N_4123,N_4708);
nor U5300 (N_5300,N_4741,N_4735);
nand U5301 (N_5301,N_4857,N_4944);
nand U5302 (N_5302,N_4897,N_4151);
xnor U5303 (N_5303,N_4886,N_4838);
and U5304 (N_5304,N_4217,N_4255);
or U5305 (N_5305,N_4277,N_4891);
and U5306 (N_5306,N_4315,N_4820);
or U5307 (N_5307,N_4047,N_4654);
or U5308 (N_5308,N_4860,N_4752);
and U5309 (N_5309,N_4856,N_4586);
xor U5310 (N_5310,N_4112,N_4458);
or U5311 (N_5311,N_4115,N_4134);
xor U5312 (N_5312,N_4875,N_4589);
or U5313 (N_5313,N_4179,N_4962);
nor U5314 (N_5314,N_4727,N_4826);
and U5315 (N_5315,N_4659,N_4342);
nand U5316 (N_5316,N_4270,N_4734);
nor U5317 (N_5317,N_4511,N_4674);
xor U5318 (N_5318,N_4144,N_4579);
nor U5319 (N_5319,N_4390,N_4988);
xnor U5320 (N_5320,N_4125,N_4863);
and U5321 (N_5321,N_4866,N_4894);
nor U5322 (N_5322,N_4538,N_4303);
xnor U5323 (N_5323,N_4668,N_4901);
and U5324 (N_5324,N_4682,N_4182);
or U5325 (N_5325,N_4933,N_4088);
and U5326 (N_5326,N_4486,N_4698);
nor U5327 (N_5327,N_4823,N_4707);
nor U5328 (N_5328,N_4139,N_4119);
or U5329 (N_5329,N_4374,N_4889);
xor U5330 (N_5330,N_4398,N_4841);
xor U5331 (N_5331,N_4903,N_4618);
and U5332 (N_5332,N_4335,N_4806);
nor U5333 (N_5333,N_4898,N_4104);
xnor U5334 (N_5334,N_4032,N_4483);
nor U5335 (N_5335,N_4985,N_4644);
xnor U5336 (N_5336,N_4083,N_4082);
nand U5337 (N_5337,N_4136,N_4330);
or U5338 (N_5338,N_4491,N_4534);
nor U5339 (N_5339,N_4317,N_4719);
nand U5340 (N_5340,N_4328,N_4530);
and U5341 (N_5341,N_4403,N_4560);
and U5342 (N_5342,N_4522,N_4325);
or U5343 (N_5343,N_4846,N_4138);
or U5344 (N_5344,N_4905,N_4433);
xor U5345 (N_5345,N_4562,N_4504);
and U5346 (N_5346,N_4163,N_4762);
or U5347 (N_5347,N_4966,N_4720);
or U5348 (N_5348,N_4011,N_4425);
nor U5349 (N_5349,N_4005,N_4792);
nand U5350 (N_5350,N_4925,N_4055);
or U5351 (N_5351,N_4716,N_4684);
and U5352 (N_5352,N_4400,N_4361);
nand U5353 (N_5353,N_4812,N_4391);
nor U5354 (N_5354,N_4412,N_4945);
nor U5355 (N_5355,N_4301,N_4819);
and U5356 (N_5356,N_4429,N_4999);
nor U5357 (N_5357,N_4637,N_4977);
or U5358 (N_5358,N_4591,N_4795);
and U5359 (N_5359,N_4527,N_4861);
nand U5360 (N_5360,N_4949,N_4836);
xnor U5361 (N_5361,N_4427,N_4308);
and U5362 (N_5362,N_4195,N_4850);
or U5363 (N_5363,N_4210,N_4050);
and U5364 (N_5364,N_4816,N_4232);
xor U5365 (N_5365,N_4272,N_4249);
nand U5366 (N_5366,N_4481,N_4928);
and U5367 (N_5367,N_4810,N_4646);
nand U5368 (N_5368,N_4069,N_4238);
and U5369 (N_5369,N_4276,N_4918);
xnor U5370 (N_5370,N_4078,N_4111);
nor U5371 (N_5371,N_4321,N_4956);
xnor U5372 (N_5372,N_4475,N_4019);
and U5373 (N_5373,N_4404,N_4353);
nand U5374 (N_5374,N_4037,N_4100);
and U5375 (N_5375,N_4149,N_4993);
nor U5376 (N_5376,N_4054,N_4683);
and U5377 (N_5377,N_4934,N_4655);
xor U5378 (N_5378,N_4061,N_4548);
or U5379 (N_5379,N_4649,N_4438);
nor U5380 (N_5380,N_4302,N_4767);
and U5381 (N_5381,N_4635,N_4224);
nand U5382 (N_5382,N_4344,N_4137);
nand U5383 (N_5383,N_4103,N_4286);
or U5384 (N_5384,N_4777,N_4778);
xnor U5385 (N_5385,N_4880,N_4542);
or U5386 (N_5386,N_4262,N_4567);
nand U5387 (N_5387,N_4197,N_4566);
nand U5388 (N_5388,N_4715,N_4007);
xor U5389 (N_5389,N_4738,N_4048);
nand U5390 (N_5390,N_4237,N_4338);
and U5391 (N_5391,N_4531,N_4899);
nor U5392 (N_5392,N_4389,N_4609);
nand U5393 (N_5393,N_4869,N_4370);
and U5394 (N_5394,N_4982,N_4518);
nor U5395 (N_5395,N_4466,N_4706);
xor U5396 (N_5396,N_4747,N_4225);
nor U5397 (N_5397,N_4554,N_4797);
nand U5398 (N_5398,N_4477,N_4395);
nor U5399 (N_5399,N_4758,N_4419);
and U5400 (N_5400,N_4053,N_4479);
nand U5401 (N_5401,N_4380,N_4761);
xor U5402 (N_5402,N_4469,N_4452);
or U5403 (N_5403,N_4954,N_4229);
or U5404 (N_5404,N_4383,N_4239);
xnor U5405 (N_5405,N_4432,N_4278);
or U5406 (N_5406,N_4871,N_4779);
nor U5407 (N_5407,N_4113,N_4357);
xor U5408 (N_5408,N_4748,N_4809);
and U5409 (N_5409,N_4322,N_4713);
or U5410 (N_5410,N_4540,N_4681);
and U5411 (N_5411,N_4524,N_4294);
xor U5412 (N_5412,N_4643,N_4316);
xnor U5413 (N_5413,N_4967,N_4890);
nor U5414 (N_5414,N_4140,N_4632);
xnor U5415 (N_5415,N_4639,N_4274);
nor U5416 (N_5416,N_4187,N_4919);
nor U5417 (N_5417,N_4957,N_4157);
xor U5418 (N_5418,N_4564,N_4497);
xor U5419 (N_5419,N_4785,N_4193);
xnor U5420 (N_5420,N_4888,N_4375);
and U5421 (N_5421,N_4221,N_4845);
or U5422 (N_5422,N_4018,N_4961);
or U5423 (N_5423,N_4601,N_4309);
nand U5424 (N_5424,N_4487,N_4189);
and U5425 (N_5425,N_4075,N_4951);
nor U5426 (N_5426,N_4496,N_4473);
nand U5427 (N_5427,N_4533,N_4811);
or U5428 (N_5428,N_4544,N_4902);
or U5429 (N_5429,N_4034,N_4245);
xnor U5430 (N_5430,N_4631,N_4960);
nand U5431 (N_5431,N_4196,N_4384);
xor U5432 (N_5432,N_4756,N_4044);
or U5433 (N_5433,N_4549,N_4581);
xnor U5434 (N_5434,N_4118,N_4373);
nand U5435 (N_5435,N_4434,N_4035);
and U5436 (N_5436,N_4613,N_4911);
xor U5437 (N_5437,N_4653,N_4367);
xor U5438 (N_5438,N_4004,N_4677);
xnor U5439 (N_5439,N_4550,N_4376);
xor U5440 (N_5440,N_4723,N_4058);
or U5441 (N_5441,N_4161,N_4467);
nor U5442 (N_5442,N_4352,N_4923);
nor U5443 (N_5443,N_4764,N_4870);
or U5444 (N_5444,N_4331,N_4651);
and U5445 (N_5445,N_4464,N_4670);
xor U5446 (N_5446,N_4180,N_4926);
nand U5447 (N_5447,N_4076,N_4942);
nand U5448 (N_5448,N_4721,N_4680);
or U5449 (N_5449,N_4754,N_4595);
nor U5450 (N_5450,N_4626,N_4020);
and U5451 (N_5451,N_4307,N_4172);
nor U5452 (N_5452,N_4444,N_4753);
and U5453 (N_5453,N_4066,N_4571);
xor U5454 (N_5454,N_4598,N_4211);
nand U5455 (N_5455,N_4783,N_4688);
or U5456 (N_5456,N_4040,N_4593);
and U5457 (N_5457,N_4130,N_4160);
nor U5458 (N_5458,N_4230,N_4226);
and U5459 (N_5459,N_4722,N_4198);
nand U5460 (N_5460,N_4915,N_4236);
or U5461 (N_5461,N_4946,N_4031);
nand U5462 (N_5462,N_4864,N_4610);
nand U5463 (N_5463,N_4913,N_4787);
xor U5464 (N_5464,N_4940,N_4176);
or U5465 (N_5465,N_4606,N_4736);
or U5466 (N_5466,N_4283,N_4501);
and U5467 (N_5467,N_4638,N_4228);
nand U5468 (N_5468,N_4010,N_4833);
and U5469 (N_5469,N_4478,N_4551);
nand U5470 (N_5470,N_4039,N_4268);
nor U5471 (N_5471,N_4784,N_4424);
nand U5472 (N_5472,N_4091,N_4565);
nor U5473 (N_5473,N_4605,N_4622);
nand U5474 (N_5474,N_4793,N_4691);
nor U5475 (N_5475,N_4349,N_4489);
or U5476 (N_5476,N_4379,N_4974);
nor U5477 (N_5477,N_4243,N_4859);
nand U5478 (N_5478,N_4821,N_4443);
nor U5479 (N_5479,N_4051,N_4456);
and U5480 (N_5480,N_4987,N_4997);
nand U5481 (N_5481,N_4012,N_4667);
xnor U5482 (N_5482,N_4326,N_4382);
xnor U5483 (N_5483,N_4953,N_4830);
or U5484 (N_5484,N_4482,N_4726);
or U5485 (N_5485,N_4737,N_4526);
or U5486 (N_5486,N_4392,N_4067);
nand U5487 (N_5487,N_4506,N_4017);
nor U5488 (N_5488,N_4159,N_4602);
nor U5489 (N_5489,N_4563,N_4247);
nand U5490 (N_5490,N_4929,N_4128);
nor U5491 (N_5491,N_4647,N_4260);
and U5492 (N_5492,N_4241,N_4537);
and U5493 (N_5493,N_4996,N_4332);
nand U5494 (N_5494,N_4336,N_4465);
nor U5495 (N_5495,N_4941,N_4697);
and U5496 (N_5496,N_4120,N_4377);
nor U5497 (N_5497,N_4963,N_4528);
xnor U5498 (N_5498,N_4690,N_4955);
nor U5499 (N_5499,N_4401,N_4188);
xor U5500 (N_5500,N_4360,N_4126);
xnor U5501 (N_5501,N_4454,N_4928);
and U5502 (N_5502,N_4203,N_4318);
or U5503 (N_5503,N_4350,N_4518);
nor U5504 (N_5504,N_4079,N_4071);
and U5505 (N_5505,N_4066,N_4301);
and U5506 (N_5506,N_4392,N_4334);
nand U5507 (N_5507,N_4993,N_4401);
nand U5508 (N_5508,N_4270,N_4945);
nor U5509 (N_5509,N_4143,N_4663);
nand U5510 (N_5510,N_4604,N_4832);
or U5511 (N_5511,N_4782,N_4595);
xor U5512 (N_5512,N_4548,N_4739);
or U5513 (N_5513,N_4393,N_4842);
or U5514 (N_5514,N_4576,N_4391);
and U5515 (N_5515,N_4327,N_4035);
or U5516 (N_5516,N_4662,N_4309);
xor U5517 (N_5517,N_4139,N_4529);
xnor U5518 (N_5518,N_4406,N_4622);
or U5519 (N_5519,N_4777,N_4290);
and U5520 (N_5520,N_4702,N_4461);
or U5521 (N_5521,N_4469,N_4532);
nand U5522 (N_5522,N_4594,N_4820);
and U5523 (N_5523,N_4837,N_4119);
nand U5524 (N_5524,N_4440,N_4796);
nor U5525 (N_5525,N_4572,N_4658);
xor U5526 (N_5526,N_4940,N_4184);
nand U5527 (N_5527,N_4652,N_4098);
and U5528 (N_5528,N_4116,N_4579);
xor U5529 (N_5529,N_4822,N_4402);
and U5530 (N_5530,N_4566,N_4845);
and U5531 (N_5531,N_4427,N_4524);
xnor U5532 (N_5532,N_4656,N_4937);
and U5533 (N_5533,N_4965,N_4651);
nor U5534 (N_5534,N_4113,N_4915);
nor U5535 (N_5535,N_4892,N_4111);
and U5536 (N_5536,N_4303,N_4181);
or U5537 (N_5537,N_4139,N_4327);
xnor U5538 (N_5538,N_4661,N_4657);
xnor U5539 (N_5539,N_4794,N_4328);
nor U5540 (N_5540,N_4381,N_4457);
nor U5541 (N_5541,N_4315,N_4155);
nor U5542 (N_5542,N_4837,N_4143);
xor U5543 (N_5543,N_4568,N_4519);
or U5544 (N_5544,N_4005,N_4850);
nor U5545 (N_5545,N_4377,N_4321);
xor U5546 (N_5546,N_4918,N_4858);
nor U5547 (N_5547,N_4642,N_4527);
nor U5548 (N_5548,N_4962,N_4207);
nor U5549 (N_5549,N_4228,N_4322);
or U5550 (N_5550,N_4291,N_4571);
or U5551 (N_5551,N_4444,N_4490);
or U5552 (N_5552,N_4273,N_4037);
or U5553 (N_5553,N_4048,N_4097);
nor U5554 (N_5554,N_4585,N_4731);
or U5555 (N_5555,N_4391,N_4185);
nor U5556 (N_5556,N_4301,N_4460);
xnor U5557 (N_5557,N_4887,N_4393);
nor U5558 (N_5558,N_4849,N_4688);
nor U5559 (N_5559,N_4299,N_4534);
or U5560 (N_5560,N_4123,N_4387);
or U5561 (N_5561,N_4340,N_4947);
nor U5562 (N_5562,N_4182,N_4708);
nand U5563 (N_5563,N_4635,N_4706);
xor U5564 (N_5564,N_4262,N_4835);
nand U5565 (N_5565,N_4280,N_4064);
nor U5566 (N_5566,N_4555,N_4265);
nor U5567 (N_5567,N_4305,N_4702);
xnor U5568 (N_5568,N_4394,N_4859);
and U5569 (N_5569,N_4752,N_4156);
and U5570 (N_5570,N_4216,N_4901);
and U5571 (N_5571,N_4409,N_4335);
nand U5572 (N_5572,N_4471,N_4648);
xor U5573 (N_5573,N_4545,N_4124);
or U5574 (N_5574,N_4557,N_4166);
nand U5575 (N_5575,N_4012,N_4684);
nand U5576 (N_5576,N_4270,N_4698);
or U5577 (N_5577,N_4660,N_4910);
xnor U5578 (N_5578,N_4138,N_4010);
nand U5579 (N_5579,N_4691,N_4642);
and U5580 (N_5580,N_4522,N_4315);
xor U5581 (N_5581,N_4161,N_4167);
nor U5582 (N_5582,N_4776,N_4509);
or U5583 (N_5583,N_4327,N_4678);
and U5584 (N_5584,N_4876,N_4073);
xnor U5585 (N_5585,N_4124,N_4505);
nand U5586 (N_5586,N_4031,N_4026);
xor U5587 (N_5587,N_4936,N_4860);
and U5588 (N_5588,N_4460,N_4503);
and U5589 (N_5589,N_4276,N_4962);
xnor U5590 (N_5590,N_4698,N_4191);
nor U5591 (N_5591,N_4537,N_4396);
nand U5592 (N_5592,N_4850,N_4764);
and U5593 (N_5593,N_4823,N_4329);
xnor U5594 (N_5594,N_4533,N_4987);
nand U5595 (N_5595,N_4504,N_4177);
xor U5596 (N_5596,N_4152,N_4283);
nand U5597 (N_5597,N_4209,N_4385);
nand U5598 (N_5598,N_4137,N_4090);
nor U5599 (N_5599,N_4557,N_4763);
nor U5600 (N_5600,N_4083,N_4877);
nor U5601 (N_5601,N_4814,N_4063);
or U5602 (N_5602,N_4780,N_4790);
and U5603 (N_5603,N_4040,N_4993);
xor U5604 (N_5604,N_4636,N_4642);
or U5605 (N_5605,N_4318,N_4536);
or U5606 (N_5606,N_4983,N_4339);
xor U5607 (N_5607,N_4458,N_4421);
nand U5608 (N_5608,N_4760,N_4224);
and U5609 (N_5609,N_4038,N_4395);
xor U5610 (N_5610,N_4308,N_4252);
xor U5611 (N_5611,N_4020,N_4091);
nor U5612 (N_5612,N_4077,N_4481);
nor U5613 (N_5613,N_4697,N_4659);
nand U5614 (N_5614,N_4138,N_4364);
or U5615 (N_5615,N_4211,N_4890);
and U5616 (N_5616,N_4184,N_4983);
xor U5617 (N_5617,N_4258,N_4412);
xor U5618 (N_5618,N_4651,N_4006);
nand U5619 (N_5619,N_4066,N_4659);
nor U5620 (N_5620,N_4943,N_4403);
and U5621 (N_5621,N_4008,N_4698);
and U5622 (N_5622,N_4100,N_4669);
nor U5623 (N_5623,N_4888,N_4148);
nor U5624 (N_5624,N_4569,N_4863);
nand U5625 (N_5625,N_4091,N_4702);
or U5626 (N_5626,N_4345,N_4451);
xnor U5627 (N_5627,N_4924,N_4440);
nand U5628 (N_5628,N_4589,N_4575);
nor U5629 (N_5629,N_4576,N_4655);
nand U5630 (N_5630,N_4174,N_4862);
nand U5631 (N_5631,N_4689,N_4774);
nor U5632 (N_5632,N_4747,N_4228);
or U5633 (N_5633,N_4570,N_4940);
nand U5634 (N_5634,N_4273,N_4269);
or U5635 (N_5635,N_4579,N_4698);
nor U5636 (N_5636,N_4722,N_4564);
xor U5637 (N_5637,N_4071,N_4617);
and U5638 (N_5638,N_4384,N_4868);
and U5639 (N_5639,N_4661,N_4823);
and U5640 (N_5640,N_4164,N_4710);
or U5641 (N_5641,N_4460,N_4432);
and U5642 (N_5642,N_4876,N_4940);
or U5643 (N_5643,N_4100,N_4636);
nand U5644 (N_5644,N_4097,N_4313);
or U5645 (N_5645,N_4939,N_4937);
xnor U5646 (N_5646,N_4084,N_4885);
and U5647 (N_5647,N_4314,N_4278);
and U5648 (N_5648,N_4336,N_4894);
and U5649 (N_5649,N_4076,N_4166);
nand U5650 (N_5650,N_4630,N_4219);
and U5651 (N_5651,N_4169,N_4325);
xnor U5652 (N_5652,N_4955,N_4277);
nand U5653 (N_5653,N_4888,N_4566);
nand U5654 (N_5654,N_4467,N_4898);
xor U5655 (N_5655,N_4124,N_4311);
xor U5656 (N_5656,N_4786,N_4038);
nand U5657 (N_5657,N_4430,N_4242);
or U5658 (N_5658,N_4983,N_4958);
nor U5659 (N_5659,N_4335,N_4420);
xnor U5660 (N_5660,N_4520,N_4861);
or U5661 (N_5661,N_4211,N_4641);
or U5662 (N_5662,N_4920,N_4386);
xor U5663 (N_5663,N_4670,N_4980);
xor U5664 (N_5664,N_4679,N_4247);
nor U5665 (N_5665,N_4058,N_4998);
and U5666 (N_5666,N_4689,N_4095);
xnor U5667 (N_5667,N_4296,N_4985);
nor U5668 (N_5668,N_4607,N_4965);
nand U5669 (N_5669,N_4727,N_4384);
nor U5670 (N_5670,N_4850,N_4979);
nor U5671 (N_5671,N_4592,N_4847);
nand U5672 (N_5672,N_4881,N_4644);
xor U5673 (N_5673,N_4929,N_4689);
and U5674 (N_5674,N_4273,N_4899);
nor U5675 (N_5675,N_4540,N_4942);
and U5676 (N_5676,N_4900,N_4812);
and U5677 (N_5677,N_4269,N_4845);
and U5678 (N_5678,N_4142,N_4766);
nand U5679 (N_5679,N_4054,N_4009);
xnor U5680 (N_5680,N_4826,N_4720);
or U5681 (N_5681,N_4365,N_4884);
or U5682 (N_5682,N_4310,N_4262);
nand U5683 (N_5683,N_4975,N_4683);
and U5684 (N_5684,N_4820,N_4000);
nor U5685 (N_5685,N_4383,N_4981);
and U5686 (N_5686,N_4651,N_4709);
nor U5687 (N_5687,N_4814,N_4016);
and U5688 (N_5688,N_4226,N_4481);
or U5689 (N_5689,N_4869,N_4953);
or U5690 (N_5690,N_4545,N_4501);
xor U5691 (N_5691,N_4718,N_4736);
nand U5692 (N_5692,N_4403,N_4459);
and U5693 (N_5693,N_4843,N_4336);
or U5694 (N_5694,N_4461,N_4515);
and U5695 (N_5695,N_4704,N_4370);
or U5696 (N_5696,N_4954,N_4245);
and U5697 (N_5697,N_4313,N_4586);
and U5698 (N_5698,N_4690,N_4958);
xnor U5699 (N_5699,N_4312,N_4244);
nor U5700 (N_5700,N_4113,N_4240);
nor U5701 (N_5701,N_4046,N_4706);
xor U5702 (N_5702,N_4211,N_4657);
and U5703 (N_5703,N_4142,N_4294);
or U5704 (N_5704,N_4425,N_4994);
nand U5705 (N_5705,N_4004,N_4237);
xnor U5706 (N_5706,N_4541,N_4265);
nor U5707 (N_5707,N_4433,N_4244);
nor U5708 (N_5708,N_4961,N_4999);
nand U5709 (N_5709,N_4958,N_4052);
nor U5710 (N_5710,N_4625,N_4787);
nand U5711 (N_5711,N_4255,N_4164);
xnor U5712 (N_5712,N_4827,N_4196);
xnor U5713 (N_5713,N_4420,N_4959);
nand U5714 (N_5714,N_4283,N_4601);
nor U5715 (N_5715,N_4005,N_4214);
or U5716 (N_5716,N_4194,N_4167);
or U5717 (N_5717,N_4532,N_4240);
nand U5718 (N_5718,N_4078,N_4691);
nand U5719 (N_5719,N_4464,N_4515);
xnor U5720 (N_5720,N_4777,N_4242);
xnor U5721 (N_5721,N_4117,N_4005);
nand U5722 (N_5722,N_4467,N_4384);
or U5723 (N_5723,N_4488,N_4655);
or U5724 (N_5724,N_4342,N_4593);
xor U5725 (N_5725,N_4891,N_4133);
nand U5726 (N_5726,N_4730,N_4310);
nand U5727 (N_5727,N_4572,N_4600);
nor U5728 (N_5728,N_4652,N_4121);
nand U5729 (N_5729,N_4117,N_4622);
nand U5730 (N_5730,N_4493,N_4519);
xor U5731 (N_5731,N_4187,N_4179);
nand U5732 (N_5732,N_4833,N_4074);
nor U5733 (N_5733,N_4626,N_4388);
nor U5734 (N_5734,N_4659,N_4011);
xor U5735 (N_5735,N_4793,N_4620);
nand U5736 (N_5736,N_4001,N_4944);
and U5737 (N_5737,N_4122,N_4368);
and U5738 (N_5738,N_4354,N_4553);
xnor U5739 (N_5739,N_4726,N_4537);
nand U5740 (N_5740,N_4495,N_4257);
nand U5741 (N_5741,N_4553,N_4261);
and U5742 (N_5742,N_4822,N_4770);
and U5743 (N_5743,N_4338,N_4642);
nand U5744 (N_5744,N_4727,N_4218);
and U5745 (N_5745,N_4803,N_4759);
xor U5746 (N_5746,N_4659,N_4681);
nand U5747 (N_5747,N_4103,N_4792);
or U5748 (N_5748,N_4216,N_4835);
xor U5749 (N_5749,N_4631,N_4803);
nor U5750 (N_5750,N_4735,N_4311);
or U5751 (N_5751,N_4835,N_4489);
or U5752 (N_5752,N_4563,N_4576);
or U5753 (N_5753,N_4972,N_4024);
or U5754 (N_5754,N_4829,N_4947);
xnor U5755 (N_5755,N_4826,N_4660);
xnor U5756 (N_5756,N_4491,N_4423);
or U5757 (N_5757,N_4127,N_4979);
or U5758 (N_5758,N_4668,N_4272);
xnor U5759 (N_5759,N_4398,N_4434);
or U5760 (N_5760,N_4015,N_4411);
nand U5761 (N_5761,N_4671,N_4150);
and U5762 (N_5762,N_4739,N_4273);
and U5763 (N_5763,N_4863,N_4109);
or U5764 (N_5764,N_4552,N_4883);
and U5765 (N_5765,N_4172,N_4885);
or U5766 (N_5766,N_4462,N_4476);
nand U5767 (N_5767,N_4425,N_4566);
and U5768 (N_5768,N_4910,N_4065);
or U5769 (N_5769,N_4817,N_4723);
nor U5770 (N_5770,N_4903,N_4332);
or U5771 (N_5771,N_4130,N_4364);
nand U5772 (N_5772,N_4693,N_4475);
nor U5773 (N_5773,N_4979,N_4117);
xnor U5774 (N_5774,N_4415,N_4035);
xnor U5775 (N_5775,N_4575,N_4548);
or U5776 (N_5776,N_4618,N_4175);
nor U5777 (N_5777,N_4788,N_4564);
nor U5778 (N_5778,N_4498,N_4780);
nand U5779 (N_5779,N_4488,N_4125);
nor U5780 (N_5780,N_4395,N_4734);
and U5781 (N_5781,N_4047,N_4899);
or U5782 (N_5782,N_4220,N_4818);
nor U5783 (N_5783,N_4807,N_4767);
nor U5784 (N_5784,N_4295,N_4991);
and U5785 (N_5785,N_4044,N_4204);
or U5786 (N_5786,N_4311,N_4250);
and U5787 (N_5787,N_4343,N_4978);
and U5788 (N_5788,N_4471,N_4570);
nor U5789 (N_5789,N_4294,N_4089);
nand U5790 (N_5790,N_4125,N_4609);
nor U5791 (N_5791,N_4313,N_4707);
nor U5792 (N_5792,N_4103,N_4276);
nor U5793 (N_5793,N_4858,N_4813);
and U5794 (N_5794,N_4363,N_4835);
and U5795 (N_5795,N_4491,N_4510);
nor U5796 (N_5796,N_4237,N_4617);
nor U5797 (N_5797,N_4410,N_4971);
and U5798 (N_5798,N_4018,N_4590);
xnor U5799 (N_5799,N_4749,N_4667);
nand U5800 (N_5800,N_4452,N_4356);
nor U5801 (N_5801,N_4608,N_4249);
nand U5802 (N_5802,N_4637,N_4033);
nor U5803 (N_5803,N_4753,N_4746);
and U5804 (N_5804,N_4923,N_4347);
nand U5805 (N_5805,N_4593,N_4388);
xnor U5806 (N_5806,N_4651,N_4335);
nor U5807 (N_5807,N_4709,N_4139);
nor U5808 (N_5808,N_4017,N_4755);
or U5809 (N_5809,N_4477,N_4244);
nand U5810 (N_5810,N_4474,N_4852);
xnor U5811 (N_5811,N_4779,N_4395);
xnor U5812 (N_5812,N_4725,N_4976);
nor U5813 (N_5813,N_4495,N_4608);
xnor U5814 (N_5814,N_4923,N_4117);
nor U5815 (N_5815,N_4442,N_4336);
or U5816 (N_5816,N_4475,N_4334);
or U5817 (N_5817,N_4289,N_4256);
and U5818 (N_5818,N_4366,N_4941);
or U5819 (N_5819,N_4748,N_4862);
nand U5820 (N_5820,N_4330,N_4420);
xnor U5821 (N_5821,N_4081,N_4854);
nand U5822 (N_5822,N_4589,N_4615);
nor U5823 (N_5823,N_4219,N_4982);
xor U5824 (N_5824,N_4834,N_4588);
or U5825 (N_5825,N_4728,N_4049);
nand U5826 (N_5826,N_4146,N_4571);
nor U5827 (N_5827,N_4428,N_4778);
xnor U5828 (N_5828,N_4929,N_4114);
nor U5829 (N_5829,N_4445,N_4831);
nor U5830 (N_5830,N_4264,N_4018);
nand U5831 (N_5831,N_4191,N_4106);
or U5832 (N_5832,N_4384,N_4466);
or U5833 (N_5833,N_4395,N_4155);
xor U5834 (N_5834,N_4386,N_4471);
or U5835 (N_5835,N_4403,N_4297);
or U5836 (N_5836,N_4799,N_4638);
xor U5837 (N_5837,N_4289,N_4318);
xnor U5838 (N_5838,N_4904,N_4836);
or U5839 (N_5839,N_4553,N_4032);
xor U5840 (N_5840,N_4004,N_4683);
nor U5841 (N_5841,N_4761,N_4514);
nand U5842 (N_5842,N_4226,N_4539);
and U5843 (N_5843,N_4945,N_4239);
or U5844 (N_5844,N_4393,N_4295);
and U5845 (N_5845,N_4150,N_4457);
nand U5846 (N_5846,N_4219,N_4791);
and U5847 (N_5847,N_4394,N_4905);
nor U5848 (N_5848,N_4893,N_4120);
and U5849 (N_5849,N_4338,N_4718);
and U5850 (N_5850,N_4058,N_4030);
nand U5851 (N_5851,N_4272,N_4038);
nor U5852 (N_5852,N_4640,N_4842);
and U5853 (N_5853,N_4337,N_4797);
xnor U5854 (N_5854,N_4839,N_4079);
or U5855 (N_5855,N_4414,N_4124);
or U5856 (N_5856,N_4655,N_4672);
or U5857 (N_5857,N_4724,N_4526);
nor U5858 (N_5858,N_4886,N_4427);
nand U5859 (N_5859,N_4934,N_4888);
or U5860 (N_5860,N_4191,N_4866);
nor U5861 (N_5861,N_4760,N_4349);
nor U5862 (N_5862,N_4254,N_4324);
xnor U5863 (N_5863,N_4481,N_4112);
xor U5864 (N_5864,N_4668,N_4144);
or U5865 (N_5865,N_4922,N_4545);
nor U5866 (N_5866,N_4431,N_4437);
nor U5867 (N_5867,N_4272,N_4721);
xor U5868 (N_5868,N_4197,N_4556);
xor U5869 (N_5869,N_4556,N_4484);
nor U5870 (N_5870,N_4077,N_4723);
or U5871 (N_5871,N_4502,N_4205);
xor U5872 (N_5872,N_4047,N_4637);
nand U5873 (N_5873,N_4601,N_4468);
nand U5874 (N_5874,N_4915,N_4135);
xor U5875 (N_5875,N_4335,N_4011);
nand U5876 (N_5876,N_4114,N_4354);
nand U5877 (N_5877,N_4780,N_4201);
nand U5878 (N_5878,N_4001,N_4681);
nand U5879 (N_5879,N_4164,N_4735);
xnor U5880 (N_5880,N_4647,N_4604);
and U5881 (N_5881,N_4832,N_4670);
xor U5882 (N_5882,N_4986,N_4960);
xnor U5883 (N_5883,N_4583,N_4085);
and U5884 (N_5884,N_4171,N_4391);
nand U5885 (N_5885,N_4930,N_4706);
xnor U5886 (N_5886,N_4117,N_4672);
nor U5887 (N_5887,N_4516,N_4926);
nand U5888 (N_5888,N_4233,N_4079);
and U5889 (N_5889,N_4752,N_4791);
and U5890 (N_5890,N_4698,N_4825);
xnor U5891 (N_5891,N_4061,N_4971);
and U5892 (N_5892,N_4164,N_4850);
xor U5893 (N_5893,N_4666,N_4304);
or U5894 (N_5894,N_4086,N_4862);
and U5895 (N_5895,N_4863,N_4138);
nor U5896 (N_5896,N_4013,N_4819);
or U5897 (N_5897,N_4090,N_4629);
and U5898 (N_5898,N_4818,N_4535);
nand U5899 (N_5899,N_4883,N_4367);
nand U5900 (N_5900,N_4058,N_4421);
nor U5901 (N_5901,N_4547,N_4241);
or U5902 (N_5902,N_4634,N_4881);
and U5903 (N_5903,N_4983,N_4265);
nor U5904 (N_5904,N_4861,N_4087);
nor U5905 (N_5905,N_4910,N_4337);
and U5906 (N_5906,N_4098,N_4741);
nor U5907 (N_5907,N_4093,N_4875);
xor U5908 (N_5908,N_4855,N_4631);
and U5909 (N_5909,N_4512,N_4341);
xor U5910 (N_5910,N_4804,N_4643);
and U5911 (N_5911,N_4376,N_4542);
nand U5912 (N_5912,N_4504,N_4604);
nand U5913 (N_5913,N_4952,N_4788);
xor U5914 (N_5914,N_4625,N_4529);
nand U5915 (N_5915,N_4250,N_4526);
nor U5916 (N_5916,N_4512,N_4288);
xor U5917 (N_5917,N_4025,N_4437);
and U5918 (N_5918,N_4626,N_4586);
nand U5919 (N_5919,N_4115,N_4677);
or U5920 (N_5920,N_4520,N_4812);
and U5921 (N_5921,N_4056,N_4799);
nor U5922 (N_5922,N_4949,N_4972);
or U5923 (N_5923,N_4152,N_4831);
nand U5924 (N_5924,N_4682,N_4373);
and U5925 (N_5925,N_4366,N_4026);
and U5926 (N_5926,N_4979,N_4788);
nor U5927 (N_5927,N_4764,N_4121);
and U5928 (N_5928,N_4655,N_4463);
and U5929 (N_5929,N_4222,N_4610);
nor U5930 (N_5930,N_4498,N_4764);
xor U5931 (N_5931,N_4248,N_4352);
nor U5932 (N_5932,N_4949,N_4230);
nand U5933 (N_5933,N_4462,N_4294);
and U5934 (N_5934,N_4592,N_4697);
nand U5935 (N_5935,N_4959,N_4025);
and U5936 (N_5936,N_4871,N_4795);
and U5937 (N_5937,N_4557,N_4569);
nand U5938 (N_5938,N_4100,N_4552);
nor U5939 (N_5939,N_4202,N_4311);
or U5940 (N_5940,N_4013,N_4903);
and U5941 (N_5941,N_4555,N_4728);
nand U5942 (N_5942,N_4713,N_4211);
and U5943 (N_5943,N_4052,N_4514);
nor U5944 (N_5944,N_4836,N_4244);
or U5945 (N_5945,N_4563,N_4490);
or U5946 (N_5946,N_4330,N_4739);
nor U5947 (N_5947,N_4408,N_4745);
nand U5948 (N_5948,N_4705,N_4475);
nand U5949 (N_5949,N_4532,N_4238);
xor U5950 (N_5950,N_4045,N_4617);
nand U5951 (N_5951,N_4842,N_4107);
or U5952 (N_5952,N_4846,N_4938);
or U5953 (N_5953,N_4067,N_4780);
or U5954 (N_5954,N_4790,N_4593);
nand U5955 (N_5955,N_4633,N_4519);
and U5956 (N_5956,N_4772,N_4694);
nor U5957 (N_5957,N_4746,N_4274);
nor U5958 (N_5958,N_4935,N_4967);
nor U5959 (N_5959,N_4932,N_4836);
xor U5960 (N_5960,N_4292,N_4587);
xor U5961 (N_5961,N_4654,N_4806);
nand U5962 (N_5962,N_4795,N_4998);
nor U5963 (N_5963,N_4981,N_4765);
or U5964 (N_5964,N_4445,N_4478);
xor U5965 (N_5965,N_4237,N_4449);
nor U5966 (N_5966,N_4231,N_4195);
or U5967 (N_5967,N_4220,N_4294);
or U5968 (N_5968,N_4527,N_4982);
xnor U5969 (N_5969,N_4432,N_4170);
or U5970 (N_5970,N_4361,N_4545);
nor U5971 (N_5971,N_4408,N_4664);
xor U5972 (N_5972,N_4054,N_4411);
or U5973 (N_5973,N_4066,N_4101);
or U5974 (N_5974,N_4027,N_4039);
xor U5975 (N_5975,N_4902,N_4960);
nand U5976 (N_5976,N_4782,N_4747);
and U5977 (N_5977,N_4466,N_4498);
nand U5978 (N_5978,N_4789,N_4210);
xor U5979 (N_5979,N_4712,N_4608);
and U5980 (N_5980,N_4957,N_4687);
nor U5981 (N_5981,N_4358,N_4301);
nand U5982 (N_5982,N_4170,N_4799);
and U5983 (N_5983,N_4106,N_4233);
xnor U5984 (N_5984,N_4450,N_4724);
nand U5985 (N_5985,N_4042,N_4110);
xor U5986 (N_5986,N_4764,N_4186);
xnor U5987 (N_5987,N_4769,N_4963);
nor U5988 (N_5988,N_4303,N_4096);
or U5989 (N_5989,N_4884,N_4732);
nand U5990 (N_5990,N_4657,N_4087);
nand U5991 (N_5991,N_4679,N_4129);
or U5992 (N_5992,N_4012,N_4579);
nand U5993 (N_5993,N_4354,N_4483);
nor U5994 (N_5994,N_4282,N_4767);
and U5995 (N_5995,N_4947,N_4911);
and U5996 (N_5996,N_4179,N_4827);
or U5997 (N_5997,N_4111,N_4720);
nand U5998 (N_5998,N_4425,N_4661);
and U5999 (N_5999,N_4498,N_4932);
or U6000 (N_6000,N_5987,N_5099);
and U6001 (N_6001,N_5983,N_5362);
nor U6002 (N_6002,N_5677,N_5676);
xnor U6003 (N_6003,N_5960,N_5997);
and U6004 (N_6004,N_5013,N_5111);
and U6005 (N_6005,N_5233,N_5882);
and U6006 (N_6006,N_5338,N_5282);
nand U6007 (N_6007,N_5656,N_5605);
xnor U6008 (N_6008,N_5312,N_5352);
nor U6009 (N_6009,N_5105,N_5924);
or U6010 (N_6010,N_5119,N_5116);
nor U6011 (N_6011,N_5059,N_5660);
and U6012 (N_6012,N_5829,N_5556);
xnor U6013 (N_6013,N_5745,N_5032);
and U6014 (N_6014,N_5106,N_5768);
or U6015 (N_6015,N_5216,N_5847);
nand U6016 (N_6016,N_5658,N_5690);
or U6017 (N_6017,N_5365,N_5182);
xnor U6018 (N_6018,N_5292,N_5540);
and U6019 (N_6019,N_5158,N_5699);
nand U6020 (N_6020,N_5388,N_5856);
or U6021 (N_6021,N_5323,N_5469);
or U6022 (N_6022,N_5998,N_5104);
and U6023 (N_6023,N_5194,N_5543);
and U6024 (N_6024,N_5439,N_5327);
nand U6025 (N_6025,N_5669,N_5070);
xor U6026 (N_6026,N_5319,N_5253);
nor U6027 (N_6027,N_5207,N_5057);
xor U6028 (N_6028,N_5552,N_5991);
nand U6029 (N_6029,N_5386,N_5189);
or U6030 (N_6030,N_5947,N_5376);
and U6031 (N_6031,N_5822,N_5892);
and U6032 (N_6032,N_5243,N_5524);
nor U6033 (N_6033,N_5979,N_5037);
nor U6034 (N_6034,N_5113,N_5795);
nand U6035 (N_6035,N_5023,N_5334);
or U6036 (N_6036,N_5891,N_5497);
nand U6037 (N_6037,N_5166,N_5068);
nor U6038 (N_6038,N_5496,N_5721);
nor U6039 (N_6039,N_5484,N_5051);
or U6040 (N_6040,N_5739,N_5094);
or U6041 (N_6041,N_5844,N_5849);
xor U6042 (N_6042,N_5575,N_5980);
xnor U6043 (N_6043,N_5049,N_5830);
xor U6044 (N_6044,N_5781,N_5747);
and U6045 (N_6045,N_5761,N_5949);
nor U6046 (N_6046,N_5221,N_5817);
and U6047 (N_6047,N_5904,N_5261);
and U6048 (N_6048,N_5090,N_5010);
nor U6049 (N_6049,N_5145,N_5294);
nand U6050 (N_6050,N_5283,N_5564);
nand U6051 (N_6051,N_5277,N_5918);
xnor U6052 (N_6052,N_5887,N_5246);
nor U6053 (N_6053,N_5250,N_5984);
nor U6054 (N_6054,N_5193,N_5837);
nand U6055 (N_6055,N_5160,N_5164);
or U6056 (N_6056,N_5877,N_5616);
xor U6057 (N_6057,N_5908,N_5176);
and U6058 (N_6058,N_5625,N_5003);
nand U6059 (N_6059,N_5255,N_5736);
and U6060 (N_6060,N_5228,N_5153);
and U6061 (N_6061,N_5371,N_5492);
nand U6062 (N_6062,N_5775,N_5760);
nor U6063 (N_6063,N_5071,N_5159);
nor U6064 (N_6064,N_5195,N_5171);
or U6065 (N_6065,N_5652,N_5405);
xnor U6066 (N_6066,N_5594,N_5401);
nor U6067 (N_6067,N_5619,N_5092);
xor U6068 (N_6068,N_5035,N_5417);
or U6069 (N_6069,N_5936,N_5640);
xor U6070 (N_6070,N_5396,N_5664);
or U6071 (N_6071,N_5331,N_5724);
xnor U6072 (N_6072,N_5535,N_5890);
and U6073 (N_6073,N_5462,N_5144);
or U6074 (N_6074,N_5500,N_5336);
nor U6075 (N_6075,N_5265,N_5266);
nor U6076 (N_6076,N_5612,N_5898);
and U6077 (N_6077,N_5999,N_5911);
and U6078 (N_6078,N_5796,N_5852);
nand U6079 (N_6079,N_5038,N_5722);
or U6080 (N_6080,N_5648,N_5379);
xor U6081 (N_6081,N_5063,N_5082);
nand U6082 (N_6082,N_5900,N_5709);
and U6083 (N_6083,N_5028,N_5916);
or U6084 (N_6084,N_5345,N_5222);
nand U6085 (N_6085,N_5298,N_5181);
or U6086 (N_6086,N_5783,N_5123);
xor U6087 (N_6087,N_5322,N_5878);
nor U6088 (N_6088,N_5374,N_5416);
nor U6089 (N_6089,N_5521,N_5742);
and U6090 (N_6090,N_5458,N_5730);
and U6091 (N_6091,N_5083,N_5039);
xnor U6092 (N_6092,N_5093,N_5131);
and U6093 (N_6093,N_5758,N_5438);
xor U6094 (N_6094,N_5787,N_5637);
nor U6095 (N_6095,N_5433,N_5180);
xor U6096 (N_6096,N_5102,N_5529);
nor U6097 (N_6097,N_5383,N_5456);
and U6098 (N_6098,N_5513,N_5988);
nor U6099 (N_6099,N_5128,N_5996);
nand U6100 (N_6100,N_5303,N_5451);
nand U6101 (N_6101,N_5251,N_5689);
or U6102 (N_6102,N_5151,N_5806);
nor U6103 (N_6103,N_5259,N_5910);
or U6104 (N_6104,N_5271,N_5315);
nor U6105 (N_6105,N_5413,N_5499);
or U6106 (N_6106,N_5792,N_5431);
nor U6107 (N_6107,N_5707,N_5974);
nor U6108 (N_6108,N_5268,N_5241);
or U6109 (N_6109,N_5297,N_5651);
nand U6110 (N_6110,N_5753,N_5380);
and U6111 (N_6111,N_5737,N_5710);
xnor U6112 (N_6112,N_5369,N_5686);
nor U6113 (N_6113,N_5186,N_5884);
xor U6114 (N_6114,N_5069,N_5992);
and U6115 (N_6115,N_5349,N_5870);
and U6116 (N_6116,N_5247,N_5940);
or U6117 (N_6117,N_5718,N_5248);
nor U6118 (N_6118,N_5986,N_5426);
xor U6119 (N_6119,N_5672,N_5667);
nor U6120 (N_6120,N_5725,N_5871);
nand U6121 (N_6121,N_5596,N_5206);
xnor U6122 (N_6122,N_5731,N_5236);
and U6123 (N_6123,N_5223,N_5569);
nor U6124 (N_6124,N_5634,N_5771);
nand U6125 (N_6125,N_5354,N_5138);
nand U6126 (N_6126,N_5534,N_5022);
nand U6127 (N_6127,N_5278,N_5378);
or U6128 (N_6128,N_5593,N_5002);
xor U6129 (N_6129,N_5237,N_5928);
nand U6130 (N_6130,N_5344,N_5025);
or U6131 (N_6131,N_5729,N_5628);
or U6132 (N_6132,N_5889,N_5422);
xor U6133 (N_6133,N_5165,N_5385);
nor U6134 (N_6134,N_5033,N_5894);
nand U6135 (N_6135,N_5136,N_5178);
nor U6136 (N_6136,N_5544,N_5864);
or U6137 (N_6137,N_5445,N_5395);
xnor U6138 (N_6138,N_5518,N_5860);
nor U6139 (N_6139,N_5079,N_5842);
or U6140 (N_6140,N_5018,N_5200);
or U6141 (N_6141,N_5767,N_5258);
nand U6142 (N_6142,N_5262,N_5715);
nor U6143 (N_6143,N_5876,N_5012);
or U6144 (N_6144,N_5693,N_5666);
nor U6145 (N_6145,N_5784,N_5957);
nor U6146 (N_6146,N_5735,N_5506);
nand U6147 (N_6147,N_5091,N_5542);
or U6148 (N_6148,N_5218,N_5252);
and U6149 (N_6149,N_5343,N_5565);
and U6150 (N_6150,N_5804,N_5415);
nand U6151 (N_6151,N_5559,N_5351);
nand U6152 (N_6152,N_5821,N_5608);
or U6153 (N_6153,N_5211,N_5580);
nand U6154 (N_6154,N_5779,N_5454);
xor U6155 (N_6155,N_5342,N_5016);
xnor U6156 (N_6156,N_5636,N_5762);
xor U6157 (N_6157,N_5641,N_5448);
nand U6158 (N_6158,N_5948,N_5697);
xor U6159 (N_6159,N_5647,N_5224);
and U6160 (N_6160,N_5723,N_5600);
xor U6161 (N_6161,N_5525,N_5526);
or U6162 (N_6162,N_5883,N_5240);
and U6163 (N_6163,N_5538,N_5360);
and U6164 (N_6164,N_5897,N_5520);
nor U6165 (N_6165,N_5087,N_5219);
or U6166 (N_6166,N_5464,N_5649);
nand U6167 (N_6167,N_5851,N_5537);
nand U6168 (N_6168,N_5711,N_5845);
nor U6169 (N_6169,N_5933,N_5481);
or U6170 (N_6170,N_5156,N_5147);
xor U6171 (N_6171,N_5930,N_5843);
or U6172 (N_6172,N_5316,N_5814);
or U6173 (N_6173,N_5973,N_5389);
xnor U6174 (N_6174,N_5313,N_5067);
nor U6175 (N_6175,N_5981,N_5811);
nor U6176 (N_6176,N_5777,N_5375);
or U6177 (N_6177,N_5807,N_5027);
nand U6178 (N_6178,N_5623,N_5727);
or U6179 (N_6179,N_5956,N_5053);
and U6180 (N_6180,N_5961,N_5286);
nor U6181 (N_6181,N_5474,N_5923);
xor U6182 (N_6182,N_5635,N_5531);
and U6183 (N_6183,N_5793,N_5185);
or U6184 (N_6184,N_5065,N_5561);
and U6185 (N_6185,N_5553,N_5129);
nand U6186 (N_6186,N_5587,N_5472);
xor U6187 (N_6187,N_5225,N_5942);
nor U6188 (N_6188,N_5260,N_5337);
or U6189 (N_6189,N_5455,N_5467);
nand U6190 (N_6190,N_5072,N_5560);
or U6191 (N_6191,N_5075,N_5485);
xor U6192 (N_6192,N_5643,N_5205);
xnor U6193 (N_6193,N_5137,N_5734);
and U6194 (N_6194,N_5938,N_5061);
xor U6195 (N_6195,N_5886,N_5846);
or U6196 (N_6196,N_5631,N_5790);
nor U6197 (N_6197,N_5550,N_5966);
nand U6198 (N_6198,N_5749,N_5130);
xor U6199 (N_6199,N_5488,N_5346);
or U6200 (N_6200,N_5632,N_5601);
nor U6201 (N_6201,N_5468,N_5935);
xnor U6202 (N_6202,N_5473,N_5859);
or U6203 (N_6203,N_5517,N_5486);
and U6204 (N_6204,N_5763,N_5339);
or U6205 (N_6205,N_5659,N_5058);
nor U6206 (N_6206,N_5572,N_5769);
xor U6207 (N_6207,N_5915,N_5579);
nor U6208 (N_6208,N_5650,N_5630);
xor U6209 (N_6209,N_5397,N_5217);
or U6210 (N_6210,N_5008,N_5245);
xnor U6211 (N_6211,N_5080,N_5620);
xor U6212 (N_6212,N_5357,N_5394);
or U6213 (N_6213,N_5967,N_5364);
xor U6214 (N_6214,N_5163,N_5203);
xor U6215 (N_6215,N_5755,N_5198);
nor U6216 (N_6216,N_5183,N_5744);
nor U6217 (N_6217,N_5424,N_5511);
xor U6218 (N_6218,N_5532,N_5429);
nand U6219 (N_6219,N_5654,N_5952);
nor U6220 (N_6220,N_5305,N_5503);
and U6221 (N_6221,N_5421,N_5411);
and U6222 (N_6222,N_5828,N_5528);
and U6223 (N_6223,N_5665,N_5645);
nand U6224 (N_6224,N_5668,N_5021);
nor U6225 (N_6225,N_5042,N_5671);
nor U6226 (N_6226,N_5126,N_5698);
nand U6227 (N_6227,N_5150,N_5704);
xor U6228 (N_6228,N_5085,N_5172);
nor U6229 (N_6229,N_5533,N_5382);
xor U6230 (N_6230,N_5614,N_5340);
and U6231 (N_6231,N_5404,N_5662);
or U6232 (N_6232,N_5865,N_5447);
nand U6233 (N_6233,N_5452,N_5308);
or U6234 (N_6234,N_5302,N_5490);
nor U6235 (N_6235,N_5853,N_5854);
and U6236 (N_6236,N_5306,N_5293);
nor U6237 (N_6237,N_5043,N_5873);
or U6238 (N_6238,N_5155,N_5201);
nand U6239 (N_6239,N_5937,N_5475);
nor U6240 (N_6240,N_5504,N_5419);
xor U6241 (N_6241,N_5695,N_5459);
xor U6242 (N_6242,N_5964,N_5366);
nand U6243 (N_6243,N_5902,N_5242);
xor U6244 (N_6244,N_5231,N_5780);
nand U6245 (N_6245,N_5489,N_5899);
nor U6246 (N_6246,N_5188,N_5570);
nor U6247 (N_6247,N_5196,N_5922);
xor U6248 (N_6248,N_5311,N_5152);
or U6249 (N_6249,N_5096,N_5017);
nand U6250 (N_6250,N_5990,N_5670);
nor U6251 (N_6251,N_5446,N_5962);
or U6252 (N_6252,N_5861,N_5140);
xnor U6253 (N_6253,N_5406,N_5696);
nor U6254 (N_6254,N_5493,N_5191);
and U6255 (N_6255,N_5402,N_5434);
nand U6256 (N_6256,N_5480,N_5300);
and U6257 (N_6257,N_5751,N_5318);
nor U6258 (N_6258,N_5358,N_5809);
nor U6259 (N_6259,N_5329,N_5232);
or U6260 (N_6260,N_5494,N_5442);
nor U6261 (N_6261,N_5591,N_5951);
and U6262 (N_6262,N_5309,N_5428);
or U6263 (N_6263,N_5945,N_5972);
and U6264 (N_6264,N_5210,N_5187);
xor U6265 (N_6265,N_5505,N_5786);
or U6266 (N_6266,N_5436,N_5443);
nor U6267 (N_6267,N_5244,N_5179);
xnor U6268 (N_6268,N_5420,N_5098);
or U6269 (N_6269,N_5192,N_5571);
and U6270 (N_6270,N_5355,N_5133);
nor U6271 (N_6271,N_5026,N_5862);
nor U6272 (N_6272,N_5269,N_5024);
or U6273 (N_6273,N_5976,N_5954);
nor U6274 (N_6274,N_5674,N_5052);
xnor U6275 (N_6275,N_5994,N_5284);
or U6276 (N_6276,N_5348,N_5603);
nor U6277 (N_6277,N_5705,N_5040);
or U6278 (N_6278,N_5530,N_5523);
nand U6279 (N_6279,N_5885,N_5879);
or U6280 (N_6280,N_5373,N_5800);
xnor U6281 (N_6281,N_5978,N_5062);
nor U6282 (N_6282,N_5273,N_5554);
nor U6283 (N_6283,N_5341,N_5363);
or U6284 (N_6284,N_5400,N_5606);
nor U6285 (N_6285,N_5076,N_5479);
nand U6286 (N_6286,N_5384,N_5437);
and U6287 (N_6287,N_5077,N_5955);
xnor U6288 (N_6288,N_5617,N_5418);
and U6289 (N_6289,N_5307,N_5127);
xor U6290 (N_6290,N_5169,N_5675);
xor U6291 (N_6291,N_5778,N_5757);
and U6292 (N_6292,N_5719,N_5613);
nand U6293 (N_6293,N_5799,N_5791);
or U6294 (N_6294,N_5320,N_5820);
nor U6295 (N_6295,N_5254,N_5919);
xor U6296 (N_6296,N_5581,N_5177);
and U6297 (N_6297,N_5726,N_5673);
and U6298 (N_6298,N_5272,N_5546);
nor U6299 (N_6299,N_5754,N_5512);
nor U6300 (N_6300,N_5819,N_5574);
nor U6301 (N_6301,N_5107,N_5141);
and U6302 (N_6302,N_5408,N_5638);
and U6303 (N_6303,N_5970,N_5208);
and U6304 (N_6304,N_5713,N_5963);
or U6305 (N_6305,N_5202,N_5772);
nand U6306 (N_6306,N_5005,N_5679);
or U6307 (N_6307,N_5212,N_5470);
nand U6308 (N_6308,N_5190,N_5112);
or U6309 (N_6309,N_5314,N_5483);
xnor U6310 (N_6310,N_5607,N_5234);
nand U6311 (N_6311,N_5858,N_5646);
xnor U6312 (N_6312,N_5678,N_5036);
nand U6313 (N_6313,N_5162,N_5326);
and U6314 (N_6314,N_5088,N_5353);
nor U6315 (N_6315,N_5597,N_5808);
xnor U6316 (N_6316,N_5466,N_5683);
or U6317 (N_6317,N_5827,N_5450);
nand U6318 (N_6318,N_5797,N_5491);
nand U6319 (N_6319,N_5618,N_5423);
xnor U6320 (N_6320,N_5281,N_5465);
nor U6321 (N_6321,N_5680,N_5595);
nor U6322 (N_6322,N_5831,N_5114);
xnor U6323 (N_6323,N_5598,N_5100);
nor U6324 (N_6324,N_5142,N_5330);
nand U6325 (N_6325,N_5582,N_5931);
xor U6326 (N_6326,N_5044,N_5425);
nand U6327 (N_6327,N_5545,N_5084);
nand U6328 (N_6328,N_5161,N_5139);
nand U6329 (N_6329,N_5004,N_5290);
xnor U6330 (N_6330,N_5551,N_5220);
nand U6331 (N_6331,N_5122,N_5276);
or U6332 (N_6332,N_5001,N_5839);
and U6333 (N_6333,N_5154,N_5317);
nor U6334 (N_6334,N_5782,N_5081);
nand U6335 (N_6335,N_5982,N_5056);
xor U6336 (N_6336,N_5971,N_5167);
or U6337 (N_6337,N_5946,N_5498);
xor U6338 (N_6338,N_5132,N_5818);
nand U6339 (N_6339,N_5019,N_5295);
or U6340 (N_6340,N_5324,N_5953);
nand U6341 (N_6341,N_5086,N_5014);
or U6342 (N_6342,N_5841,N_5350);
nand U6343 (N_6343,N_5875,N_5639);
xnor U6344 (N_6344,N_5562,N_5548);
nand U6345 (N_6345,N_5449,N_5684);
and U6346 (N_6346,N_5287,N_5288);
and U6347 (N_6347,N_5975,N_5732);
nor U6348 (N_6348,N_5381,N_5785);
xor U6349 (N_6349,N_5304,N_5661);
nor U6350 (N_6350,N_5020,N_5440);
or U6351 (N_6351,N_5586,N_5888);
and U6352 (N_6352,N_5078,N_5321);
or U6353 (N_6353,N_5299,N_5706);
nor U6354 (N_6354,N_5399,N_5692);
nor U6355 (N_6355,N_5563,N_5622);
nand U6356 (N_6356,N_5653,N_5274);
nand U6357 (N_6357,N_5146,N_5691);
or U6358 (N_6358,N_5229,N_5627);
or U6359 (N_6359,N_5700,N_5694);
xnor U6360 (N_6360,N_5507,N_5110);
or U6361 (N_6361,N_5633,N_5912);
nor U6362 (N_6362,N_5174,N_5584);
nor U6363 (N_6363,N_5759,N_5514);
and U6364 (N_6364,N_5738,N_5515);
nor U6365 (N_6365,N_5913,N_5066);
nand U6366 (N_6366,N_5270,N_5642);
xnor U6367 (N_6367,N_5685,N_5235);
or U6368 (N_6368,N_5810,N_5264);
nand U6369 (N_6369,N_5588,N_5377);
xor U6370 (N_6370,N_5748,N_5741);
nor U6371 (N_6371,N_5046,N_5011);
nand U6372 (N_6372,N_5624,N_5301);
and U6373 (N_6373,N_5566,N_5604);
xor U6374 (N_6374,N_5527,N_5041);
nand U6375 (N_6375,N_5427,N_5412);
xnor U6376 (N_6376,N_5495,N_5239);
and U6377 (N_6377,N_5789,N_5770);
and U6378 (N_6378,N_5134,N_5432);
xor U6379 (N_6379,N_5108,N_5589);
nand U6380 (N_6380,N_5609,N_5501);
xnor U6381 (N_6381,N_5850,N_5204);
nor U6382 (N_6382,N_5249,N_5280);
and U6383 (N_6383,N_5097,N_5279);
or U6384 (N_6384,N_5907,N_5708);
nor U6385 (N_6385,N_5143,N_5215);
nand U6386 (N_6386,N_5905,N_5199);
or U6387 (N_6387,N_5578,N_5536);
nand U6388 (N_6388,N_5929,N_5788);
nand U6389 (N_6389,N_5407,N_5644);
nand U6390 (N_6390,N_5168,N_5743);
or U6391 (N_6391,N_5773,N_5109);
nand U6392 (N_6392,N_5958,N_5539);
nand U6393 (N_6393,N_5989,N_5558);
xor U6394 (N_6394,N_5914,N_5444);
nor U6395 (N_6395,N_5510,N_5868);
xnor U6396 (N_6396,N_5663,N_5629);
xor U6397 (N_6397,N_5335,N_5920);
xor U6398 (N_6398,N_5977,N_5476);
xnor U6399 (N_6399,N_5173,N_5801);
or U6400 (N_6400,N_5615,N_5157);
or U6401 (N_6401,N_5688,N_5824);
nand U6402 (N_6402,N_5602,N_5256);
xor U6403 (N_6403,N_5117,N_5909);
and U6404 (N_6404,N_5263,N_5519);
nor U6405 (N_6405,N_5881,N_5508);
xor U6406 (N_6406,N_5895,N_5869);
nand U6407 (N_6407,N_5590,N_5047);
and U6408 (N_6408,N_5740,N_5720);
or U6409 (N_6409,N_5657,N_5866);
or U6410 (N_6410,N_5390,N_5227);
nor U6411 (N_6411,N_5985,N_5863);
nor U6412 (N_6412,N_5387,N_5009);
nor U6413 (N_6413,N_5457,N_5880);
and U6414 (N_6414,N_5682,N_5815);
and U6415 (N_6415,N_5502,N_5555);
xor U6416 (N_6416,N_5776,N_5702);
xor U6417 (N_6417,N_5124,N_5175);
nor U6418 (N_6418,N_5393,N_5074);
nor U6419 (N_6419,N_5823,N_5714);
or U6420 (N_6420,N_5712,N_5054);
or U6421 (N_6421,N_5872,N_5611);
and U6422 (N_6422,N_5006,N_5917);
nand U6423 (N_6423,N_5592,N_5968);
or U6424 (N_6424,N_5214,N_5029);
nor U6425 (N_6425,N_5701,N_5209);
xor U6426 (N_6426,N_5257,N_5549);
and U6427 (N_6427,N_5230,N_5944);
and U6428 (N_6428,N_5120,N_5655);
and U6429 (N_6429,N_5766,N_5728);
nand U6430 (N_6430,N_5803,N_5626);
and U6431 (N_6431,N_5568,N_5703);
nand U6432 (N_6432,N_5328,N_5487);
or U6433 (N_6433,N_5332,N_5893);
xnor U6434 (N_6434,N_5943,N_5838);
nor U6435 (N_6435,N_5347,N_5681);
and U6436 (N_6436,N_5926,N_5836);
or U6437 (N_6437,N_5356,N_5541);
nor U6438 (N_6438,N_5361,N_5927);
xor U6439 (N_6439,N_5995,N_5950);
xnor U6440 (N_6440,N_5045,N_5857);
nor U6441 (N_6441,N_5576,N_5925);
xor U6442 (N_6442,N_5765,N_5599);
and U6443 (N_6443,N_5547,N_5463);
nor U6444 (N_6444,N_5372,N_5939);
or U6445 (N_6445,N_5573,N_5932);
nor U6446 (N_6446,N_5840,N_5125);
nand U6447 (N_6447,N_5752,N_5055);
and U6448 (N_6448,N_5073,N_5170);
xnor U6449 (N_6449,N_5410,N_5118);
or U6450 (N_6450,N_5965,N_5833);
or U6451 (N_6451,N_5941,N_5367);
and U6452 (N_6452,N_5813,N_5184);
nand U6453 (N_6453,N_5048,N_5805);
xnor U6454 (N_6454,N_5750,N_5414);
and U6455 (N_6455,N_5398,N_5289);
and U6456 (N_6456,N_5060,N_5848);
and U6457 (N_6457,N_5430,N_5103);
nand U6458 (N_6458,N_5934,N_5148);
xor U6459 (N_6459,N_5370,N_5435);
xor U6460 (N_6460,N_5064,N_5213);
or U6461 (N_6461,N_5007,N_5409);
nor U6462 (N_6462,N_5567,N_5050);
and U6463 (N_6463,N_5522,N_5906);
nor U6464 (N_6464,N_5557,N_5717);
nor U6465 (N_6465,N_5764,N_5798);
or U6466 (N_6466,N_5969,N_5135);
and U6467 (N_6467,N_5296,N_5610);
nand U6468 (N_6468,N_5482,N_5756);
nand U6469 (N_6469,N_5746,N_5325);
and U6470 (N_6470,N_5441,N_5460);
nor U6471 (N_6471,N_5903,N_5477);
and U6472 (N_6472,N_5275,N_5359);
nand U6473 (N_6473,N_5115,N_5816);
nand U6474 (N_6474,N_5867,N_5015);
and U6475 (N_6475,N_5333,N_5392);
or U6476 (N_6476,N_5687,N_5095);
nand U6477 (N_6477,N_5101,N_5461);
xnor U6478 (N_6478,N_5403,N_5000);
and U6479 (N_6479,N_5621,N_5832);
or U6480 (N_6480,N_5197,N_5921);
xnor U6481 (N_6481,N_5774,N_5577);
nand U6482 (N_6482,N_5855,N_5226);
xor U6483 (N_6483,N_5034,N_5516);
nand U6484 (N_6484,N_5391,N_5149);
nor U6485 (N_6485,N_5291,N_5802);
or U6486 (N_6486,N_5267,N_5874);
nor U6487 (N_6487,N_5794,N_5959);
and U6488 (N_6488,N_5585,N_5368);
xor U6489 (N_6489,N_5716,N_5901);
xnor U6490 (N_6490,N_5993,N_5238);
and U6491 (N_6491,N_5834,N_5825);
or U6492 (N_6492,N_5896,N_5285);
nand U6493 (N_6493,N_5509,N_5812);
nor U6494 (N_6494,N_5835,N_5310);
or U6495 (N_6495,N_5826,N_5583);
xor U6496 (N_6496,N_5453,N_5478);
nor U6497 (N_6497,N_5089,N_5031);
xnor U6498 (N_6498,N_5733,N_5471);
nor U6499 (N_6499,N_5030,N_5121);
nand U6500 (N_6500,N_5269,N_5897);
xor U6501 (N_6501,N_5456,N_5156);
and U6502 (N_6502,N_5222,N_5375);
and U6503 (N_6503,N_5786,N_5351);
or U6504 (N_6504,N_5287,N_5710);
and U6505 (N_6505,N_5792,N_5610);
xnor U6506 (N_6506,N_5448,N_5944);
and U6507 (N_6507,N_5136,N_5593);
xnor U6508 (N_6508,N_5563,N_5139);
or U6509 (N_6509,N_5187,N_5706);
xnor U6510 (N_6510,N_5032,N_5536);
or U6511 (N_6511,N_5952,N_5567);
and U6512 (N_6512,N_5906,N_5033);
xor U6513 (N_6513,N_5819,N_5006);
nor U6514 (N_6514,N_5149,N_5833);
and U6515 (N_6515,N_5622,N_5242);
or U6516 (N_6516,N_5148,N_5551);
or U6517 (N_6517,N_5108,N_5049);
and U6518 (N_6518,N_5245,N_5917);
or U6519 (N_6519,N_5039,N_5483);
nand U6520 (N_6520,N_5854,N_5665);
or U6521 (N_6521,N_5166,N_5984);
xnor U6522 (N_6522,N_5286,N_5887);
xor U6523 (N_6523,N_5510,N_5439);
or U6524 (N_6524,N_5245,N_5296);
nand U6525 (N_6525,N_5683,N_5282);
xor U6526 (N_6526,N_5084,N_5017);
xnor U6527 (N_6527,N_5437,N_5594);
and U6528 (N_6528,N_5394,N_5140);
nand U6529 (N_6529,N_5932,N_5454);
or U6530 (N_6530,N_5200,N_5229);
nand U6531 (N_6531,N_5281,N_5048);
nand U6532 (N_6532,N_5324,N_5746);
xor U6533 (N_6533,N_5355,N_5326);
or U6534 (N_6534,N_5149,N_5573);
nor U6535 (N_6535,N_5263,N_5777);
and U6536 (N_6536,N_5848,N_5503);
nand U6537 (N_6537,N_5077,N_5474);
or U6538 (N_6538,N_5065,N_5573);
nor U6539 (N_6539,N_5628,N_5339);
xnor U6540 (N_6540,N_5251,N_5838);
xnor U6541 (N_6541,N_5084,N_5580);
nor U6542 (N_6542,N_5244,N_5677);
or U6543 (N_6543,N_5346,N_5878);
and U6544 (N_6544,N_5258,N_5365);
xnor U6545 (N_6545,N_5665,N_5096);
nand U6546 (N_6546,N_5796,N_5660);
and U6547 (N_6547,N_5904,N_5488);
xnor U6548 (N_6548,N_5243,N_5052);
and U6549 (N_6549,N_5863,N_5338);
or U6550 (N_6550,N_5086,N_5443);
and U6551 (N_6551,N_5290,N_5843);
nor U6552 (N_6552,N_5343,N_5606);
nand U6553 (N_6553,N_5966,N_5399);
nor U6554 (N_6554,N_5054,N_5725);
xor U6555 (N_6555,N_5247,N_5534);
or U6556 (N_6556,N_5467,N_5995);
and U6557 (N_6557,N_5654,N_5424);
xnor U6558 (N_6558,N_5937,N_5747);
and U6559 (N_6559,N_5358,N_5688);
nor U6560 (N_6560,N_5602,N_5641);
and U6561 (N_6561,N_5020,N_5225);
or U6562 (N_6562,N_5560,N_5614);
nor U6563 (N_6563,N_5427,N_5313);
nor U6564 (N_6564,N_5779,N_5010);
nand U6565 (N_6565,N_5273,N_5497);
nand U6566 (N_6566,N_5135,N_5001);
xnor U6567 (N_6567,N_5912,N_5128);
or U6568 (N_6568,N_5568,N_5887);
or U6569 (N_6569,N_5750,N_5029);
nor U6570 (N_6570,N_5788,N_5831);
nor U6571 (N_6571,N_5466,N_5740);
or U6572 (N_6572,N_5693,N_5107);
or U6573 (N_6573,N_5207,N_5538);
or U6574 (N_6574,N_5627,N_5995);
or U6575 (N_6575,N_5497,N_5155);
xor U6576 (N_6576,N_5965,N_5210);
nor U6577 (N_6577,N_5672,N_5374);
nor U6578 (N_6578,N_5286,N_5336);
nor U6579 (N_6579,N_5600,N_5049);
nand U6580 (N_6580,N_5684,N_5010);
and U6581 (N_6581,N_5045,N_5569);
or U6582 (N_6582,N_5957,N_5713);
and U6583 (N_6583,N_5987,N_5118);
xnor U6584 (N_6584,N_5500,N_5219);
xor U6585 (N_6585,N_5225,N_5509);
nand U6586 (N_6586,N_5279,N_5368);
nand U6587 (N_6587,N_5214,N_5500);
and U6588 (N_6588,N_5516,N_5743);
xnor U6589 (N_6589,N_5701,N_5872);
nand U6590 (N_6590,N_5470,N_5992);
or U6591 (N_6591,N_5466,N_5478);
and U6592 (N_6592,N_5766,N_5363);
and U6593 (N_6593,N_5471,N_5632);
or U6594 (N_6594,N_5433,N_5490);
nor U6595 (N_6595,N_5675,N_5701);
and U6596 (N_6596,N_5640,N_5794);
or U6597 (N_6597,N_5967,N_5814);
nand U6598 (N_6598,N_5357,N_5009);
nor U6599 (N_6599,N_5240,N_5624);
or U6600 (N_6600,N_5183,N_5642);
and U6601 (N_6601,N_5765,N_5156);
or U6602 (N_6602,N_5004,N_5181);
or U6603 (N_6603,N_5933,N_5009);
nor U6604 (N_6604,N_5541,N_5676);
or U6605 (N_6605,N_5230,N_5888);
nor U6606 (N_6606,N_5296,N_5096);
and U6607 (N_6607,N_5162,N_5437);
nand U6608 (N_6608,N_5193,N_5902);
nand U6609 (N_6609,N_5251,N_5053);
and U6610 (N_6610,N_5663,N_5284);
nor U6611 (N_6611,N_5823,N_5273);
nand U6612 (N_6612,N_5487,N_5392);
or U6613 (N_6613,N_5949,N_5680);
nor U6614 (N_6614,N_5362,N_5984);
and U6615 (N_6615,N_5462,N_5515);
and U6616 (N_6616,N_5896,N_5231);
nor U6617 (N_6617,N_5105,N_5542);
nor U6618 (N_6618,N_5207,N_5820);
nor U6619 (N_6619,N_5029,N_5364);
xor U6620 (N_6620,N_5891,N_5853);
and U6621 (N_6621,N_5557,N_5168);
or U6622 (N_6622,N_5383,N_5638);
nand U6623 (N_6623,N_5420,N_5515);
nand U6624 (N_6624,N_5975,N_5958);
nor U6625 (N_6625,N_5415,N_5044);
and U6626 (N_6626,N_5070,N_5645);
nor U6627 (N_6627,N_5339,N_5850);
nor U6628 (N_6628,N_5529,N_5560);
xor U6629 (N_6629,N_5511,N_5455);
nor U6630 (N_6630,N_5473,N_5708);
nand U6631 (N_6631,N_5569,N_5519);
xnor U6632 (N_6632,N_5690,N_5270);
xnor U6633 (N_6633,N_5696,N_5105);
and U6634 (N_6634,N_5785,N_5793);
and U6635 (N_6635,N_5951,N_5398);
and U6636 (N_6636,N_5612,N_5752);
nor U6637 (N_6637,N_5428,N_5765);
nor U6638 (N_6638,N_5969,N_5466);
nor U6639 (N_6639,N_5395,N_5167);
or U6640 (N_6640,N_5964,N_5806);
and U6641 (N_6641,N_5914,N_5358);
or U6642 (N_6642,N_5341,N_5980);
xor U6643 (N_6643,N_5735,N_5707);
and U6644 (N_6644,N_5745,N_5713);
nor U6645 (N_6645,N_5574,N_5078);
nand U6646 (N_6646,N_5031,N_5192);
nand U6647 (N_6647,N_5580,N_5674);
nor U6648 (N_6648,N_5438,N_5728);
xnor U6649 (N_6649,N_5775,N_5124);
or U6650 (N_6650,N_5511,N_5082);
xor U6651 (N_6651,N_5838,N_5458);
and U6652 (N_6652,N_5969,N_5945);
xor U6653 (N_6653,N_5951,N_5280);
or U6654 (N_6654,N_5513,N_5790);
or U6655 (N_6655,N_5067,N_5139);
and U6656 (N_6656,N_5837,N_5131);
xnor U6657 (N_6657,N_5150,N_5742);
xor U6658 (N_6658,N_5329,N_5942);
xor U6659 (N_6659,N_5228,N_5333);
xor U6660 (N_6660,N_5326,N_5538);
and U6661 (N_6661,N_5533,N_5832);
and U6662 (N_6662,N_5710,N_5908);
xor U6663 (N_6663,N_5497,N_5003);
nand U6664 (N_6664,N_5775,N_5720);
or U6665 (N_6665,N_5528,N_5638);
xnor U6666 (N_6666,N_5273,N_5210);
nor U6667 (N_6667,N_5847,N_5073);
nand U6668 (N_6668,N_5080,N_5981);
nor U6669 (N_6669,N_5471,N_5741);
and U6670 (N_6670,N_5355,N_5035);
and U6671 (N_6671,N_5788,N_5765);
nand U6672 (N_6672,N_5911,N_5954);
or U6673 (N_6673,N_5980,N_5563);
nand U6674 (N_6674,N_5089,N_5100);
xnor U6675 (N_6675,N_5620,N_5114);
nand U6676 (N_6676,N_5619,N_5723);
or U6677 (N_6677,N_5563,N_5820);
xor U6678 (N_6678,N_5886,N_5508);
xor U6679 (N_6679,N_5020,N_5082);
xnor U6680 (N_6680,N_5801,N_5860);
xor U6681 (N_6681,N_5136,N_5831);
xnor U6682 (N_6682,N_5973,N_5021);
or U6683 (N_6683,N_5037,N_5428);
nor U6684 (N_6684,N_5071,N_5149);
nand U6685 (N_6685,N_5338,N_5721);
and U6686 (N_6686,N_5940,N_5331);
and U6687 (N_6687,N_5813,N_5176);
nand U6688 (N_6688,N_5924,N_5494);
and U6689 (N_6689,N_5760,N_5442);
nand U6690 (N_6690,N_5414,N_5618);
and U6691 (N_6691,N_5626,N_5686);
or U6692 (N_6692,N_5531,N_5434);
or U6693 (N_6693,N_5624,N_5167);
or U6694 (N_6694,N_5324,N_5873);
nor U6695 (N_6695,N_5182,N_5892);
nand U6696 (N_6696,N_5368,N_5312);
nor U6697 (N_6697,N_5120,N_5631);
xor U6698 (N_6698,N_5234,N_5159);
nor U6699 (N_6699,N_5720,N_5482);
nand U6700 (N_6700,N_5012,N_5682);
or U6701 (N_6701,N_5848,N_5498);
nor U6702 (N_6702,N_5686,N_5954);
or U6703 (N_6703,N_5820,N_5293);
and U6704 (N_6704,N_5412,N_5735);
nand U6705 (N_6705,N_5593,N_5999);
xor U6706 (N_6706,N_5198,N_5694);
xnor U6707 (N_6707,N_5887,N_5888);
nand U6708 (N_6708,N_5891,N_5049);
nor U6709 (N_6709,N_5871,N_5282);
nor U6710 (N_6710,N_5404,N_5171);
and U6711 (N_6711,N_5181,N_5943);
nor U6712 (N_6712,N_5281,N_5830);
xor U6713 (N_6713,N_5107,N_5365);
nor U6714 (N_6714,N_5774,N_5827);
xor U6715 (N_6715,N_5481,N_5903);
xnor U6716 (N_6716,N_5486,N_5935);
nand U6717 (N_6717,N_5051,N_5066);
or U6718 (N_6718,N_5849,N_5436);
or U6719 (N_6719,N_5990,N_5969);
xnor U6720 (N_6720,N_5750,N_5325);
nand U6721 (N_6721,N_5597,N_5128);
nand U6722 (N_6722,N_5871,N_5037);
xor U6723 (N_6723,N_5897,N_5642);
nand U6724 (N_6724,N_5704,N_5521);
and U6725 (N_6725,N_5921,N_5574);
nand U6726 (N_6726,N_5604,N_5424);
or U6727 (N_6727,N_5490,N_5422);
nand U6728 (N_6728,N_5124,N_5848);
nor U6729 (N_6729,N_5339,N_5275);
xor U6730 (N_6730,N_5347,N_5468);
nor U6731 (N_6731,N_5398,N_5902);
or U6732 (N_6732,N_5392,N_5061);
xor U6733 (N_6733,N_5749,N_5839);
nand U6734 (N_6734,N_5814,N_5248);
and U6735 (N_6735,N_5937,N_5232);
or U6736 (N_6736,N_5781,N_5816);
or U6737 (N_6737,N_5880,N_5677);
and U6738 (N_6738,N_5970,N_5237);
nor U6739 (N_6739,N_5662,N_5210);
nor U6740 (N_6740,N_5194,N_5451);
xnor U6741 (N_6741,N_5876,N_5304);
xnor U6742 (N_6742,N_5874,N_5430);
nand U6743 (N_6743,N_5415,N_5634);
nand U6744 (N_6744,N_5151,N_5378);
and U6745 (N_6745,N_5947,N_5137);
nor U6746 (N_6746,N_5381,N_5710);
nand U6747 (N_6747,N_5245,N_5932);
nor U6748 (N_6748,N_5971,N_5289);
and U6749 (N_6749,N_5304,N_5842);
xnor U6750 (N_6750,N_5124,N_5023);
or U6751 (N_6751,N_5236,N_5851);
and U6752 (N_6752,N_5154,N_5065);
and U6753 (N_6753,N_5908,N_5361);
nand U6754 (N_6754,N_5211,N_5892);
xor U6755 (N_6755,N_5122,N_5509);
or U6756 (N_6756,N_5290,N_5875);
nand U6757 (N_6757,N_5124,N_5336);
nor U6758 (N_6758,N_5065,N_5179);
xnor U6759 (N_6759,N_5319,N_5576);
xor U6760 (N_6760,N_5611,N_5339);
nor U6761 (N_6761,N_5197,N_5594);
nor U6762 (N_6762,N_5552,N_5367);
nand U6763 (N_6763,N_5583,N_5995);
nand U6764 (N_6764,N_5533,N_5204);
nand U6765 (N_6765,N_5166,N_5821);
xnor U6766 (N_6766,N_5990,N_5111);
xor U6767 (N_6767,N_5356,N_5423);
and U6768 (N_6768,N_5606,N_5485);
and U6769 (N_6769,N_5478,N_5462);
or U6770 (N_6770,N_5238,N_5715);
or U6771 (N_6771,N_5888,N_5079);
or U6772 (N_6772,N_5330,N_5579);
xor U6773 (N_6773,N_5982,N_5131);
and U6774 (N_6774,N_5040,N_5937);
or U6775 (N_6775,N_5159,N_5209);
and U6776 (N_6776,N_5304,N_5024);
xnor U6777 (N_6777,N_5186,N_5046);
and U6778 (N_6778,N_5474,N_5245);
or U6779 (N_6779,N_5097,N_5183);
nand U6780 (N_6780,N_5055,N_5990);
and U6781 (N_6781,N_5081,N_5113);
and U6782 (N_6782,N_5273,N_5372);
or U6783 (N_6783,N_5444,N_5296);
nor U6784 (N_6784,N_5630,N_5059);
xnor U6785 (N_6785,N_5899,N_5908);
nand U6786 (N_6786,N_5842,N_5388);
nand U6787 (N_6787,N_5884,N_5923);
or U6788 (N_6788,N_5620,N_5434);
and U6789 (N_6789,N_5969,N_5763);
nand U6790 (N_6790,N_5323,N_5098);
and U6791 (N_6791,N_5424,N_5997);
and U6792 (N_6792,N_5132,N_5235);
and U6793 (N_6793,N_5155,N_5823);
or U6794 (N_6794,N_5727,N_5587);
xnor U6795 (N_6795,N_5962,N_5503);
xnor U6796 (N_6796,N_5431,N_5268);
or U6797 (N_6797,N_5063,N_5670);
or U6798 (N_6798,N_5078,N_5745);
or U6799 (N_6799,N_5134,N_5511);
and U6800 (N_6800,N_5290,N_5627);
nand U6801 (N_6801,N_5536,N_5642);
nor U6802 (N_6802,N_5655,N_5788);
and U6803 (N_6803,N_5080,N_5081);
nor U6804 (N_6804,N_5327,N_5731);
xor U6805 (N_6805,N_5121,N_5672);
nor U6806 (N_6806,N_5261,N_5834);
or U6807 (N_6807,N_5143,N_5083);
nand U6808 (N_6808,N_5655,N_5985);
xor U6809 (N_6809,N_5629,N_5583);
xor U6810 (N_6810,N_5417,N_5283);
nand U6811 (N_6811,N_5011,N_5563);
or U6812 (N_6812,N_5748,N_5252);
xnor U6813 (N_6813,N_5311,N_5478);
nor U6814 (N_6814,N_5281,N_5160);
nor U6815 (N_6815,N_5520,N_5415);
nor U6816 (N_6816,N_5034,N_5159);
nand U6817 (N_6817,N_5540,N_5162);
xor U6818 (N_6818,N_5640,N_5281);
xor U6819 (N_6819,N_5330,N_5187);
xor U6820 (N_6820,N_5406,N_5226);
nand U6821 (N_6821,N_5631,N_5877);
or U6822 (N_6822,N_5941,N_5576);
nand U6823 (N_6823,N_5725,N_5168);
and U6824 (N_6824,N_5515,N_5285);
and U6825 (N_6825,N_5599,N_5629);
xnor U6826 (N_6826,N_5282,N_5329);
and U6827 (N_6827,N_5907,N_5840);
nor U6828 (N_6828,N_5714,N_5103);
and U6829 (N_6829,N_5363,N_5447);
or U6830 (N_6830,N_5937,N_5622);
and U6831 (N_6831,N_5447,N_5589);
or U6832 (N_6832,N_5137,N_5748);
or U6833 (N_6833,N_5841,N_5383);
nand U6834 (N_6834,N_5078,N_5006);
nand U6835 (N_6835,N_5852,N_5913);
or U6836 (N_6836,N_5867,N_5557);
nor U6837 (N_6837,N_5604,N_5498);
nand U6838 (N_6838,N_5320,N_5488);
nor U6839 (N_6839,N_5173,N_5702);
or U6840 (N_6840,N_5926,N_5816);
or U6841 (N_6841,N_5572,N_5640);
and U6842 (N_6842,N_5211,N_5552);
nor U6843 (N_6843,N_5324,N_5243);
and U6844 (N_6844,N_5596,N_5144);
and U6845 (N_6845,N_5088,N_5264);
or U6846 (N_6846,N_5586,N_5136);
and U6847 (N_6847,N_5842,N_5245);
or U6848 (N_6848,N_5021,N_5675);
or U6849 (N_6849,N_5640,N_5553);
xor U6850 (N_6850,N_5115,N_5090);
or U6851 (N_6851,N_5644,N_5296);
and U6852 (N_6852,N_5238,N_5720);
nor U6853 (N_6853,N_5525,N_5476);
or U6854 (N_6854,N_5860,N_5915);
nor U6855 (N_6855,N_5889,N_5620);
or U6856 (N_6856,N_5571,N_5379);
or U6857 (N_6857,N_5644,N_5195);
and U6858 (N_6858,N_5259,N_5273);
xnor U6859 (N_6859,N_5072,N_5961);
nand U6860 (N_6860,N_5961,N_5049);
xor U6861 (N_6861,N_5593,N_5261);
xnor U6862 (N_6862,N_5552,N_5817);
nand U6863 (N_6863,N_5654,N_5454);
nor U6864 (N_6864,N_5871,N_5809);
or U6865 (N_6865,N_5437,N_5343);
xor U6866 (N_6866,N_5442,N_5036);
or U6867 (N_6867,N_5935,N_5951);
or U6868 (N_6868,N_5232,N_5379);
nor U6869 (N_6869,N_5904,N_5916);
xnor U6870 (N_6870,N_5395,N_5496);
and U6871 (N_6871,N_5251,N_5353);
nor U6872 (N_6872,N_5455,N_5707);
nand U6873 (N_6873,N_5628,N_5614);
nor U6874 (N_6874,N_5950,N_5058);
xnor U6875 (N_6875,N_5107,N_5463);
nand U6876 (N_6876,N_5519,N_5232);
and U6877 (N_6877,N_5465,N_5073);
nor U6878 (N_6878,N_5892,N_5475);
nand U6879 (N_6879,N_5668,N_5057);
xnor U6880 (N_6880,N_5805,N_5132);
nor U6881 (N_6881,N_5627,N_5024);
and U6882 (N_6882,N_5994,N_5402);
xnor U6883 (N_6883,N_5069,N_5744);
nand U6884 (N_6884,N_5814,N_5177);
nor U6885 (N_6885,N_5549,N_5851);
or U6886 (N_6886,N_5683,N_5624);
xnor U6887 (N_6887,N_5798,N_5835);
or U6888 (N_6888,N_5145,N_5784);
nand U6889 (N_6889,N_5951,N_5729);
or U6890 (N_6890,N_5236,N_5655);
or U6891 (N_6891,N_5980,N_5778);
nor U6892 (N_6892,N_5553,N_5393);
and U6893 (N_6893,N_5261,N_5384);
and U6894 (N_6894,N_5907,N_5568);
xor U6895 (N_6895,N_5079,N_5748);
xnor U6896 (N_6896,N_5695,N_5261);
xnor U6897 (N_6897,N_5259,N_5003);
nand U6898 (N_6898,N_5970,N_5073);
xor U6899 (N_6899,N_5414,N_5542);
xnor U6900 (N_6900,N_5295,N_5207);
xnor U6901 (N_6901,N_5448,N_5234);
xor U6902 (N_6902,N_5566,N_5192);
or U6903 (N_6903,N_5618,N_5446);
or U6904 (N_6904,N_5469,N_5949);
nor U6905 (N_6905,N_5716,N_5718);
nand U6906 (N_6906,N_5859,N_5462);
nor U6907 (N_6907,N_5570,N_5915);
nor U6908 (N_6908,N_5564,N_5440);
or U6909 (N_6909,N_5131,N_5681);
and U6910 (N_6910,N_5984,N_5763);
xnor U6911 (N_6911,N_5253,N_5107);
nor U6912 (N_6912,N_5114,N_5338);
or U6913 (N_6913,N_5631,N_5984);
or U6914 (N_6914,N_5925,N_5781);
xnor U6915 (N_6915,N_5756,N_5936);
nand U6916 (N_6916,N_5270,N_5515);
and U6917 (N_6917,N_5812,N_5791);
xnor U6918 (N_6918,N_5215,N_5654);
and U6919 (N_6919,N_5679,N_5825);
xnor U6920 (N_6920,N_5723,N_5203);
or U6921 (N_6921,N_5147,N_5432);
and U6922 (N_6922,N_5021,N_5057);
nand U6923 (N_6923,N_5966,N_5036);
or U6924 (N_6924,N_5906,N_5804);
xor U6925 (N_6925,N_5920,N_5047);
nor U6926 (N_6926,N_5834,N_5643);
or U6927 (N_6927,N_5919,N_5894);
nor U6928 (N_6928,N_5080,N_5431);
nor U6929 (N_6929,N_5909,N_5459);
or U6930 (N_6930,N_5524,N_5994);
xnor U6931 (N_6931,N_5987,N_5157);
nor U6932 (N_6932,N_5238,N_5065);
nor U6933 (N_6933,N_5458,N_5038);
xor U6934 (N_6934,N_5090,N_5112);
and U6935 (N_6935,N_5948,N_5929);
or U6936 (N_6936,N_5601,N_5619);
nand U6937 (N_6937,N_5499,N_5736);
nand U6938 (N_6938,N_5237,N_5473);
nand U6939 (N_6939,N_5234,N_5054);
and U6940 (N_6940,N_5012,N_5627);
xor U6941 (N_6941,N_5928,N_5773);
nor U6942 (N_6942,N_5197,N_5699);
or U6943 (N_6943,N_5823,N_5254);
xor U6944 (N_6944,N_5299,N_5066);
nor U6945 (N_6945,N_5864,N_5937);
or U6946 (N_6946,N_5092,N_5670);
or U6947 (N_6947,N_5145,N_5743);
and U6948 (N_6948,N_5675,N_5742);
nand U6949 (N_6949,N_5224,N_5921);
nor U6950 (N_6950,N_5914,N_5675);
nor U6951 (N_6951,N_5030,N_5517);
nand U6952 (N_6952,N_5699,N_5270);
and U6953 (N_6953,N_5566,N_5721);
and U6954 (N_6954,N_5693,N_5002);
nor U6955 (N_6955,N_5108,N_5608);
and U6956 (N_6956,N_5562,N_5146);
xor U6957 (N_6957,N_5167,N_5318);
nor U6958 (N_6958,N_5574,N_5387);
nor U6959 (N_6959,N_5239,N_5339);
or U6960 (N_6960,N_5442,N_5210);
nand U6961 (N_6961,N_5847,N_5097);
nand U6962 (N_6962,N_5132,N_5385);
nand U6963 (N_6963,N_5953,N_5297);
xor U6964 (N_6964,N_5689,N_5623);
and U6965 (N_6965,N_5688,N_5999);
nand U6966 (N_6966,N_5594,N_5669);
xor U6967 (N_6967,N_5361,N_5983);
xnor U6968 (N_6968,N_5823,N_5227);
nand U6969 (N_6969,N_5720,N_5756);
xnor U6970 (N_6970,N_5507,N_5044);
nor U6971 (N_6971,N_5815,N_5470);
xor U6972 (N_6972,N_5154,N_5092);
and U6973 (N_6973,N_5440,N_5134);
nor U6974 (N_6974,N_5423,N_5225);
nor U6975 (N_6975,N_5475,N_5675);
nor U6976 (N_6976,N_5368,N_5965);
xor U6977 (N_6977,N_5495,N_5164);
nand U6978 (N_6978,N_5355,N_5230);
nor U6979 (N_6979,N_5782,N_5834);
nand U6980 (N_6980,N_5626,N_5322);
nand U6981 (N_6981,N_5518,N_5613);
and U6982 (N_6982,N_5912,N_5908);
nand U6983 (N_6983,N_5526,N_5022);
nand U6984 (N_6984,N_5665,N_5101);
nor U6985 (N_6985,N_5978,N_5183);
nand U6986 (N_6986,N_5141,N_5371);
and U6987 (N_6987,N_5170,N_5703);
xor U6988 (N_6988,N_5300,N_5902);
nand U6989 (N_6989,N_5203,N_5225);
nor U6990 (N_6990,N_5704,N_5788);
nor U6991 (N_6991,N_5985,N_5030);
nand U6992 (N_6992,N_5774,N_5099);
xnor U6993 (N_6993,N_5674,N_5687);
or U6994 (N_6994,N_5731,N_5735);
nand U6995 (N_6995,N_5191,N_5327);
or U6996 (N_6996,N_5229,N_5774);
xor U6997 (N_6997,N_5080,N_5833);
or U6998 (N_6998,N_5484,N_5830);
xor U6999 (N_6999,N_5858,N_5880);
nand U7000 (N_7000,N_6482,N_6696);
nand U7001 (N_7001,N_6456,N_6236);
or U7002 (N_7002,N_6868,N_6202);
and U7003 (N_7003,N_6005,N_6145);
and U7004 (N_7004,N_6462,N_6280);
or U7005 (N_7005,N_6554,N_6724);
nor U7006 (N_7006,N_6582,N_6031);
and U7007 (N_7007,N_6337,N_6458);
or U7008 (N_7008,N_6644,N_6684);
and U7009 (N_7009,N_6555,N_6949);
nor U7010 (N_7010,N_6593,N_6537);
nor U7011 (N_7011,N_6241,N_6412);
or U7012 (N_7012,N_6743,N_6927);
or U7013 (N_7013,N_6415,N_6818);
nor U7014 (N_7014,N_6703,N_6519);
and U7015 (N_7015,N_6713,N_6316);
and U7016 (N_7016,N_6066,N_6497);
or U7017 (N_7017,N_6796,N_6972);
nor U7018 (N_7018,N_6451,N_6536);
and U7019 (N_7019,N_6650,N_6774);
xor U7020 (N_7020,N_6237,N_6506);
nand U7021 (N_7021,N_6504,N_6626);
nand U7022 (N_7022,N_6449,N_6278);
nor U7023 (N_7023,N_6034,N_6538);
and U7024 (N_7024,N_6550,N_6999);
or U7025 (N_7025,N_6087,N_6384);
xnor U7026 (N_7026,N_6362,N_6764);
nand U7027 (N_7027,N_6956,N_6775);
xnor U7028 (N_7028,N_6753,N_6809);
nor U7029 (N_7029,N_6046,N_6836);
or U7030 (N_7030,N_6778,N_6030);
nand U7031 (N_7031,N_6491,N_6891);
and U7032 (N_7032,N_6111,N_6985);
or U7033 (N_7033,N_6799,N_6396);
or U7034 (N_7034,N_6833,N_6893);
and U7035 (N_7035,N_6043,N_6940);
nand U7036 (N_7036,N_6473,N_6688);
nand U7037 (N_7037,N_6975,N_6459);
or U7038 (N_7038,N_6069,N_6589);
or U7039 (N_7039,N_6392,N_6134);
and U7040 (N_7040,N_6223,N_6751);
nor U7041 (N_7041,N_6428,N_6557);
nand U7042 (N_7042,N_6932,N_6591);
xor U7043 (N_7043,N_6023,N_6705);
nor U7044 (N_7044,N_6405,N_6305);
and U7045 (N_7045,N_6991,N_6944);
xnor U7046 (N_7046,N_6240,N_6431);
and U7047 (N_7047,N_6802,N_6853);
nand U7048 (N_7048,N_6152,N_6787);
xor U7049 (N_7049,N_6026,N_6281);
and U7050 (N_7050,N_6843,N_6502);
or U7051 (N_7051,N_6277,N_6096);
xor U7052 (N_7052,N_6676,N_6664);
nor U7053 (N_7053,N_6338,N_6074);
and U7054 (N_7054,N_6749,N_6494);
nor U7055 (N_7055,N_6822,N_6807);
nor U7056 (N_7056,N_6156,N_6130);
nor U7057 (N_7057,N_6358,N_6624);
or U7058 (N_7058,N_6048,N_6974);
or U7059 (N_7059,N_6516,N_6808);
and U7060 (N_7060,N_6575,N_6307);
xnor U7061 (N_7061,N_6518,N_6413);
nor U7062 (N_7062,N_6224,N_6024);
or U7063 (N_7063,N_6765,N_6183);
or U7064 (N_7064,N_6505,N_6526);
and U7065 (N_7065,N_6158,N_6948);
xor U7066 (N_7066,N_6939,N_6056);
nand U7067 (N_7067,N_6033,N_6247);
or U7068 (N_7068,N_6792,N_6826);
and U7069 (N_7069,N_6600,N_6806);
xor U7070 (N_7070,N_6206,N_6186);
nand U7071 (N_7071,N_6585,N_6854);
nor U7072 (N_7072,N_6571,N_6106);
nor U7073 (N_7073,N_6895,N_6515);
or U7074 (N_7074,N_6539,N_6229);
or U7075 (N_7075,N_6867,N_6613);
and U7076 (N_7076,N_6093,N_6894);
or U7077 (N_7077,N_6243,N_6552);
nand U7078 (N_7078,N_6172,N_6349);
or U7079 (N_7079,N_6231,N_6119);
nor U7080 (N_7080,N_6366,N_6308);
and U7081 (N_7081,N_6101,N_6001);
nand U7082 (N_7082,N_6434,N_6865);
nand U7083 (N_7083,N_6641,N_6430);
or U7084 (N_7084,N_6579,N_6263);
xnor U7085 (N_7085,N_6837,N_6697);
nor U7086 (N_7086,N_6723,N_6282);
nor U7087 (N_7087,N_6495,N_6699);
nand U7088 (N_7088,N_6065,N_6789);
nand U7089 (N_7089,N_6059,N_6370);
xnor U7090 (N_7090,N_6100,N_6633);
nor U7091 (N_7091,N_6076,N_6672);
or U7092 (N_7092,N_6272,N_6782);
nand U7093 (N_7093,N_6943,N_6219);
xor U7094 (N_7094,N_6409,N_6619);
xor U7095 (N_7095,N_6376,N_6834);
xnor U7096 (N_7096,N_6880,N_6286);
nand U7097 (N_7097,N_6062,N_6153);
nand U7098 (N_7098,N_6524,N_6565);
and U7099 (N_7099,N_6094,N_6653);
and U7100 (N_7100,N_6900,N_6973);
nor U7101 (N_7101,N_6637,N_6324);
nand U7102 (N_7102,N_6746,N_6133);
or U7103 (N_7103,N_6884,N_6909);
or U7104 (N_7104,N_6721,N_6745);
nand U7105 (N_7105,N_6475,N_6309);
or U7106 (N_7106,N_6418,N_6549);
xor U7107 (N_7107,N_6658,N_6173);
nor U7108 (N_7108,N_6089,N_6105);
or U7109 (N_7109,N_6887,N_6192);
and U7110 (N_7110,N_6689,N_6288);
xnor U7111 (N_7111,N_6194,N_6327);
or U7112 (N_7112,N_6000,N_6960);
or U7113 (N_7113,N_6284,N_6058);
and U7114 (N_7114,N_6813,N_6769);
and U7115 (N_7115,N_6463,N_6612);
or U7116 (N_7116,N_6271,N_6332);
nor U7117 (N_7117,N_6047,N_6639);
xnor U7118 (N_7118,N_6385,N_6189);
nor U7119 (N_7119,N_6244,N_6568);
nand U7120 (N_7120,N_6828,N_6700);
or U7121 (N_7121,N_6627,N_6323);
xnor U7122 (N_7122,N_6545,N_6845);
or U7123 (N_7123,N_6166,N_6830);
and U7124 (N_7124,N_6514,N_6291);
and U7125 (N_7125,N_6762,N_6139);
or U7126 (N_7126,N_6803,N_6424);
and U7127 (N_7127,N_6197,N_6661);
nor U7128 (N_7128,N_6042,N_6322);
xnor U7129 (N_7129,N_6603,N_6343);
nand U7130 (N_7130,N_6503,N_6861);
and U7131 (N_7131,N_6544,N_6679);
and U7132 (N_7132,N_6636,N_6951);
nand U7133 (N_7133,N_6912,N_6098);
or U7134 (N_7134,N_6992,N_6786);
nand U7135 (N_7135,N_6730,N_6419);
and U7136 (N_7136,N_6262,N_6732);
xnor U7137 (N_7137,N_6234,N_6246);
xnor U7138 (N_7138,N_6325,N_6196);
and U7139 (N_7139,N_6875,N_6354);
nand U7140 (N_7140,N_6294,N_6242);
or U7141 (N_7141,N_6317,N_6261);
and U7142 (N_7142,N_6312,N_6760);
or U7143 (N_7143,N_6982,N_6274);
and U7144 (N_7144,N_6488,N_6099);
nor U7145 (N_7145,N_6566,N_6489);
or U7146 (N_7146,N_6580,N_6154);
nor U7147 (N_7147,N_6116,N_6443);
xnor U7148 (N_7148,N_6390,N_6542);
xor U7149 (N_7149,N_6090,N_6551);
or U7150 (N_7150,N_6766,N_6285);
or U7151 (N_7151,N_6731,N_6903);
nor U7152 (N_7152,N_6752,N_6962);
or U7153 (N_7153,N_6964,N_6102);
xnor U7154 (N_7154,N_6501,N_6480);
nand U7155 (N_7155,N_6330,N_6199);
or U7156 (N_7156,N_6931,N_6364);
nand U7157 (N_7157,N_6883,N_6213);
and U7158 (N_7158,N_6656,N_6870);
and U7159 (N_7159,N_6694,N_6402);
and U7160 (N_7160,N_6979,N_6435);
nand U7161 (N_7161,N_6256,N_6329);
nand U7162 (N_7162,N_6622,N_6977);
nand U7163 (N_7163,N_6588,N_6935);
xor U7164 (N_7164,N_6378,N_6556);
nand U7165 (N_7165,N_6227,N_6856);
nand U7166 (N_7166,N_6035,N_6109);
nor U7167 (N_7167,N_6107,N_6386);
xor U7168 (N_7168,N_6389,N_6669);
and U7169 (N_7169,N_6407,N_6235);
nor U7170 (N_7170,N_6598,N_6356);
xor U7171 (N_7171,N_6981,N_6850);
xnor U7172 (N_7172,N_6297,N_6476);
nand U7173 (N_7173,N_6293,N_6665);
xor U7174 (N_7174,N_6507,N_6953);
and U7175 (N_7175,N_6345,N_6768);
and U7176 (N_7176,N_6300,N_6771);
xor U7177 (N_7177,N_6645,N_6744);
nand U7178 (N_7178,N_6132,N_6060);
xnor U7179 (N_7179,N_6226,N_6313);
nor U7180 (N_7180,N_6326,N_6120);
nor U7181 (N_7181,N_6547,N_6611);
xnor U7182 (N_7182,N_6823,N_6170);
nor U7183 (N_7183,N_6399,N_6104);
or U7184 (N_7184,N_6251,N_6899);
nor U7185 (N_7185,N_6128,N_6606);
nand U7186 (N_7186,N_6904,N_6310);
and U7187 (N_7187,N_6208,N_6368);
nor U7188 (N_7188,N_6216,N_6728);
and U7189 (N_7189,N_6725,N_6414);
or U7190 (N_7190,N_6264,N_6022);
or U7191 (N_7191,N_6086,N_6441);
xnor U7192 (N_7192,N_6780,N_6188);
nor U7193 (N_7193,N_6230,N_6342);
nand U7194 (N_7194,N_6408,N_6290);
nor U7195 (N_7195,N_6773,N_6238);
nand U7196 (N_7196,N_6010,N_6432);
or U7197 (N_7197,N_6508,N_6204);
or U7198 (N_7198,N_6182,N_6155);
nand U7199 (N_7199,N_6693,N_6862);
nand U7200 (N_7200,N_6015,N_6623);
or U7201 (N_7201,N_6529,N_6602);
and U7202 (N_7202,N_6253,N_6527);
nor U7203 (N_7203,N_6346,N_6080);
nand U7204 (N_7204,N_6360,N_6011);
nor U7205 (N_7205,N_6279,N_6220);
or U7206 (N_7206,N_6680,N_6470);
and U7207 (N_7207,N_6070,N_6648);
nand U7208 (N_7208,N_6934,N_6677);
xor U7209 (N_7209,N_6314,N_6083);
xnor U7210 (N_7210,N_6455,N_6161);
nand U7211 (N_7211,N_6168,N_6250);
nor U7212 (N_7212,N_6761,N_6686);
and U7213 (N_7213,N_6930,N_6339);
or U7214 (N_7214,N_6675,N_6634);
and U7215 (N_7215,N_6481,N_6915);
nand U7216 (N_7216,N_6667,N_6484);
or U7217 (N_7217,N_6737,N_6838);
nor U7218 (N_7218,N_6925,N_6871);
and U7219 (N_7219,N_6164,N_6791);
or U7220 (N_7220,N_6423,N_6417);
and U7221 (N_7221,N_6232,N_6984);
and U7222 (N_7222,N_6049,N_6570);
nor U7223 (N_7223,N_6876,N_6827);
xor U7224 (N_7224,N_6268,N_6275);
nand U7225 (N_7225,N_6009,N_6578);
nand U7226 (N_7226,N_6006,N_6072);
xor U7227 (N_7227,N_6530,N_6304);
nor U7228 (N_7228,N_6882,N_6355);
nand U7229 (N_7229,N_6162,N_6259);
or U7230 (N_7230,N_6525,N_6397);
nand U7231 (N_7231,N_6149,N_6541);
nand U7232 (N_7232,N_6976,N_6365);
or U7233 (N_7233,N_6474,N_6276);
and U7234 (N_7234,N_6668,N_6388);
and U7235 (N_7235,N_6657,N_6453);
nand U7236 (N_7236,N_6118,N_6841);
nand U7237 (N_7237,N_6855,N_6963);
nand U7238 (N_7238,N_6905,N_6198);
nor U7239 (N_7239,N_6750,N_6215);
nor U7240 (N_7240,N_6735,N_6002);
nor U7241 (N_7241,N_6758,N_6879);
or U7242 (N_7242,N_6959,N_6564);
xor U7243 (N_7243,N_6788,N_6890);
or U7244 (N_7244,N_6692,N_6671);
or U7245 (N_7245,N_6707,N_6742);
xnor U7246 (N_7246,N_6734,N_6248);
or U7247 (N_7247,N_6496,N_6922);
xor U7248 (N_7248,N_6928,N_6805);
and U7249 (N_7249,N_6652,N_6863);
nor U7250 (N_7250,N_6517,N_6174);
and U7251 (N_7251,N_6690,N_6559);
nand U7252 (N_7252,N_6007,N_6319);
nand U7253 (N_7253,N_6763,N_6727);
xnor U7254 (N_7254,N_6531,N_6112);
nor U7255 (N_7255,N_6654,N_6151);
nor U7256 (N_7256,N_6095,N_6596);
nand U7257 (N_7257,N_6628,N_6824);
nand U7258 (N_7258,N_6126,N_6510);
or U7259 (N_7259,N_6967,N_6306);
nor U7260 (N_7260,N_6136,N_6410);
and U7261 (N_7261,N_6379,N_6500);
nor U7262 (N_7262,N_6594,N_6492);
nand U7263 (N_7263,N_6543,N_6367);
nor U7264 (N_7264,N_6228,N_6068);
nand U7265 (N_7265,N_6478,N_6157);
xnor U7266 (N_7266,N_6708,N_6181);
xnor U7267 (N_7267,N_6874,N_6950);
nand U7268 (N_7268,N_6754,N_6759);
or U7269 (N_7269,N_6642,N_6287);
or U7270 (N_7270,N_6553,N_6344);
xor U7271 (N_7271,N_6203,N_6315);
xnor U7272 (N_7272,N_6036,N_6159);
or U7273 (N_7273,N_6361,N_6144);
nor U7274 (N_7274,N_6615,N_6437);
nor U7275 (N_7275,N_6110,N_6607);
nor U7276 (N_7276,N_6886,N_6587);
and U7277 (N_7277,N_6719,N_6857);
nor U7278 (N_7278,N_6632,N_6483);
xnor U7279 (N_7279,N_6840,N_6296);
nand U7280 (N_7280,N_6438,N_6740);
nor U7281 (N_7281,N_6466,N_6937);
and U7282 (N_7282,N_6958,N_6872);
or U7283 (N_7283,N_6169,N_6866);
nand U7284 (N_7284,N_6520,N_6618);
nand U7285 (N_7285,N_6695,N_6714);
xnor U7286 (N_7286,N_6479,N_6334);
nand U7287 (N_7287,N_6584,N_6528);
and U7288 (N_7288,N_6576,N_6218);
and U7289 (N_7289,N_6121,N_6382);
nand U7290 (N_7290,N_6180,N_6425);
nor U7291 (N_7291,N_6395,N_6785);
xnor U7292 (N_7292,N_6123,N_6722);
xnor U7293 (N_7293,N_6638,N_6881);
and U7294 (N_7294,N_6336,N_6233);
and U7295 (N_7295,N_6609,N_6590);
or U7296 (N_7296,N_6113,N_6446);
and U7297 (N_7297,N_6888,N_6490);
nand U7298 (N_7298,N_6914,N_6946);
nand U7299 (N_7299,N_6640,N_6212);
or U7300 (N_7300,N_6037,N_6055);
xnor U7301 (N_7301,N_6563,N_6381);
xnor U7302 (N_7302,N_6993,N_6472);
xor U7303 (N_7303,N_6465,N_6924);
nor U7304 (N_7304,N_6698,N_6498);
and U7305 (N_7305,N_6616,N_6635);
and U7306 (N_7306,N_6968,N_6560);
xor U7307 (N_7307,N_6258,N_6117);
nor U7308 (N_7308,N_6340,N_6767);
and U7309 (N_7309,N_6835,N_6040);
nand U7310 (N_7310,N_6075,N_6393);
and U7311 (N_7311,N_6348,N_6605);
nand U7312 (N_7312,N_6630,N_6878);
xor U7313 (N_7313,N_6401,N_6165);
or U7314 (N_7314,N_6190,N_6601);
nor U7315 (N_7315,N_6885,N_6998);
nor U7316 (N_7316,N_6829,N_6269);
or U7317 (N_7317,N_6333,N_6318);
xor U7318 (N_7318,N_6921,N_6947);
nand U7319 (N_7319,N_6014,N_6077);
or U7320 (N_7320,N_6178,N_6561);
nand U7321 (N_7321,N_6273,N_6468);
or U7322 (N_7322,N_6436,N_6864);
and U7323 (N_7323,N_6716,N_6631);
nor U7324 (N_7324,N_6374,N_6179);
nand U7325 (N_7325,N_6608,N_6908);
nor U7326 (N_7326,N_6377,N_6177);
or U7327 (N_7327,N_6783,N_6629);
xor U7328 (N_7328,N_6819,N_6770);
xor U7329 (N_7329,N_6320,N_6936);
and U7330 (N_7330,N_6994,N_6917);
nor U7331 (N_7331,N_6471,N_6877);
nor U7332 (N_7332,N_6569,N_6499);
nor U7333 (N_7333,N_6896,N_6583);
nand U7334 (N_7334,N_6729,N_6018);
and U7335 (N_7335,N_6387,N_6574);
nand U7336 (N_7336,N_6039,N_6053);
and U7337 (N_7337,N_6717,N_6595);
and U7338 (N_7338,N_6997,N_6978);
or U7339 (N_7339,N_6200,N_6045);
nor U7340 (N_7340,N_6321,N_6025);
nor U7341 (N_7341,N_6439,N_6701);
nand U7342 (N_7342,N_6655,N_6239);
or U7343 (N_7343,N_6851,N_6422);
or U7344 (N_7344,N_6114,N_6777);
nor U7345 (N_7345,N_6493,N_6918);
nor U7346 (N_7346,N_6148,N_6255);
or U7347 (N_7347,N_6748,N_6711);
xnor U7348 (N_7348,N_6739,N_6146);
and U7349 (N_7349,N_6012,N_6662);
xor U7350 (N_7350,N_6184,N_6535);
nand U7351 (N_7351,N_6429,N_6050);
or U7352 (N_7352,N_6041,N_6811);
nor U7353 (N_7353,N_6311,N_6142);
or U7354 (N_7354,N_6920,N_6797);
or U7355 (N_7355,N_6678,N_6573);
nand U7356 (N_7356,N_6052,N_6398);
xor U7357 (N_7357,N_6923,N_6383);
nand U7358 (N_7358,N_6801,N_6108);
or U7359 (N_7359,N_6427,N_6741);
or U7360 (N_7360,N_6509,N_6403);
xnor U7361 (N_7361,N_6747,N_6254);
and U7362 (N_7362,N_6467,N_6683);
and U7363 (N_7363,N_6400,N_6647);
nand U7364 (N_7364,N_6426,N_6193);
or U7365 (N_7365,N_6673,N_6245);
or U7366 (N_7366,N_6084,N_6019);
xor U7367 (N_7367,N_6965,N_6757);
nand U7368 (N_7368,N_6546,N_6558);
or U7369 (N_7369,N_6511,N_6810);
and U7370 (N_7370,N_6008,N_6260);
and U7371 (N_7371,N_6457,N_6341);
xnor U7372 (N_7372,N_6902,N_6143);
xor U7373 (N_7373,N_6163,N_6670);
and U7374 (N_7374,N_6357,N_6860);
nand U7375 (N_7375,N_6176,N_6125);
nor U7376 (N_7376,N_6798,N_6625);
or U7377 (N_7377,N_6846,N_6825);
nor U7378 (N_7378,N_6996,N_6800);
xnor U7379 (N_7379,N_6267,N_6682);
nor U7380 (N_7380,N_6225,N_6444);
xnor U7381 (N_7381,N_6957,N_6421);
nand U7382 (N_7382,N_6485,N_6452);
and U7383 (N_7383,N_6597,N_6733);
and U7384 (N_7384,N_6970,N_6532);
nand U7385 (N_7385,N_6445,N_6610);
nand U7386 (N_7386,N_6523,N_6450);
or U7387 (N_7387,N_6815,N_6303);
nor U7388 (N_7388,N_6990,N_6614);
and U7389 (N_7389,N_6726,N_6859);
or U7390 (N_7390,N_6794,N_6980);
and U7391 (N_7391,N_6852,N_6351);
nand U7392 (N_7392,N_6205,N_6391);
and U7393 (N_7393,N_6933,N_6265);
nor U7394 (N_7394,N_6191,N_6869);
or U7395 (N_7395,N_6027,N_6945);
or U7396 (N_7396,N_6211,N_6844);
and U7397 (N_7397,N_6461,N_6420);
nor U7398 (N_7398,N_6522,N_6781);
xnor U7399 (N_7399,N_6987,N_6548);
and U7400 (N_7400,N_6091,N_6715);
xnor U7401 (N_7401,N_6486,N_6185);
and U7402 (N_7402,N_6270,N_6756);
nand U7403 (N_7403,N_6897,N_6704);
or U7404 (N_7404,N_6175,N_6839);
nor U7405 (N_7405,N_6129,N_6755);
and U7406 (N_7406,N_6266,N_6847);
nand U7407 (N_7407,N_6738,N_6141);
nand U7408 (N_7408,N_6460,N_6513);
xor U7409 (N_7409,N_6581,N_6988);
or U7410 (N_7410,N_6057,N_6989);
and U7411 (N_7411,N_6051,N_6941);
nor U7412 (N_7412,N_6375,N_6620);
nand U7413 (N_7413,N_6061,N_6209);
or U7414 (N_7414,N_6712,N_6350);
nor U7415 (N_7415,N_6299,N_6533);
and U7416 (N_7416,N_6586,N_6359);
and U7417 (N_7417,N_6201,N_6122);
or U7418 (N_7418,N_6849,N_6371);
xnor U7419 (N_7419,N_6659,N_6906);
xor U7420 (N_7420,N_6966,N_6831);
or U7421 (N_7421,N_6649,N_6487);
nor U7422 (N_7422,N_6454,N_6440);
nand U7423 (N_7423,N_6702,N_6044);
and U7424 (N_7424,N_6892,N_6433);
nor U7425 (N_7425,N_6814,N_6032);
nand U7426 (N_7426,N_6302,N_6352);
or U7427 (N_7427,N_6038,N_6085);
nor U7428 (N_7428,N_6131,N_6842);
and U7429 (N_7429,N_6167,N_6135);
and U7430 (N_7430,N_6150,N_6081);
xnor U7431 (N_7431,N_6898,N_6016);
and U7432 (N_7432,N_6063,N_6411);
or U7433 (N_7433,N_6889,N_6938);
or U7434 (N_7434,N_6779,N_6289);
xor U7435 (N_7435,N_6687,N_6790);
or U7436 (N_7436,N_6983,N_6369);
nand U7437 (N_7437,N_6955,N_6477);
nand U7438 (N_7438,N_6464,N_6160);
nand U7439 (N_7439,N_6078,N_6643);
or U7440 (N_7440,N_6394,N_6221);
xor U7441 (N_7441,N_6140,N_6592);
xnor U7442 (N_7442,N_6147,N_6115);
nand U7443 (N_7443,N_6404,N_6138);
nand U7444 (N_7444,N_6651,N_6907);
nand U7445 (N_7445,N_6347,N_6187);
and U7446 (N_7446,N_6406,N_6328);
and U7447 (N_7447,N_6512,N_6013);
nor U7448 (N_7448,N_6736,N_6858);
and U7449 (N_7449,N_6092,N_6812);
nand U7450 (N_7450,N_6685,N_6916);
or U7451 (N_7451,N_6848,N_6249);
nor U7452 (N_7452,N_6772,N_6222);
xnor U7453 (N_7453,N_6901,N_6252);
xnor U7454 (N_7454,N_6709,N_6660);
nand U7455 (N_7455,N_6097,N_6363);
xor U7456 (N_7456,N_6817,N_6540);
nor U7457 (N_7457,N_6416,N_6691);
nand U7458 (N_7458,N_6969,N_6919);
xor U7459 (N_7459,N_6599,N_6301);
xnor U7460 (N_7460,N_6913,N_6380);
and U7461 (N_7461,N_6674,N_6681);
and U7462 (N_7462,N_6873,N_6567);
and U7463 (N_7463,N_6710,N_6617);
nor U7464 (N_7464,N_6995,N_6028);
or U7465 (N_7465,N_6952,N_6217);
nand U7466 (N_7466,N_6521,N_6986);
xor U7467 (N_7467,N_6666,N_6562);
or U7468 (N_7468,N_6929,N_6171);
nand U7469 (N_7469,N_6832,N_6793);
nand U7470 (N_7470,N_6137,N_6706);
and U7471 (N_7471,N_6821,N_6073);
or U7472 (N_7472,N_6353,N_6292);
xor U7473 (N_7473,N_6017,N_6718);
and U7474 (N_7474,N_6816,N_6298);
nand U7475 (N_7475,N_6534,N_6804);
and U7476 (N_7476,N_6283,N_6971);
and U7477 (N_7477,N_6942,N_6447);
or U7478 (N_7478,N_6961,N_6054);
nand U7479 (N_7479,N_6373,N_6372);
xnor U7480 (N_7480,N_6448,N_6604);
or U7481 (N_7481,N_6442,N_6214);
xor U7482 (N_7482,N_6020,N_6577);
xor U7483 (N_7483,N_6021,N_6295);
and U7484 (N_7484,N_6088,N_6004);
nand U7485 (N_7485,N_6820,N_6207);
and U7486 (N_7486,N_6646,N_6911);
xor U7487 (N_7487,N_6071,N_6926);
and U7488 (N_7488,N_6067,N_6029);
nand U7489 (N_7489,N_6910,N_6335);
nor U7490 (N_7490,N_6663,N_6469);
nand U7491 (N_7491,N_6331,N_6124);
nor U7492 (N_7492,N_6064,N_6103);
xnor U7493 (N_7493,N_6082,N_6003);
or U7494 (N_7494,N_6127,N_6195);
nor U7495 (N_7495,N_6784,N_6572);
or U7496 (N_7496,N_6954,N_6795);
and U7497 (N_7497,N_6720,N_6079);
nand U7498 (N_7498,N_6776,N_6210);
nor U7499 (N_7499,N_6621,N_6257);
and U7500 (N_7500,N_6698,N_6095);
or U7501 (N_7501,N_6699,N_6007);
nor U7502 (N_7502,N_6631,N_6950);
nand U7503 (N_7503,N_6660,N_6241);
nor U7504 (N_7504,N_6049,N_6729);
or U7505 (N_7505,N_6039,N_6389);
nand U7506 (N_7506,N_6702,N_6154);
or U7507 (N_7507,N_6674,N_6179);
xor U7508 (N_7508,N_6312,N_6759);
nor U7509 (N_7509,N_6533,N_6089);
nand U7510 (N_7510,N_6521,N_6957);
xnor U7511 (N_7511,N_6976,N_6138);
xor U7512 (N_7512,N_6325,N_6776);
and U7513 (N_7513,N_6484,N_6717);
xnor U7514 (N_7514,N_6897,N_6320);
and U7515 (N_7515,N_6192,N_6261);
or U7516 (N_7516,N_6027,N_6819);
nor U7517 (N_7517,N_6781,N_6854);
or U7518 (N_7518,N_6053,N_6693);
xnor U7519 (N_7519,N_6848,N_6917);
xnor U7520 (N_7520,N_6884,N_6387);
and U7521 (N_7521,N_6419,N_6103);
or U7522 (N_7522,N_6133,N_6604);
or U7523 (N_7523,N_6123,N_6350);
or U7524 (N_7524,N_6244,N_6503);
and U7525 (N_7525,N_6454,N_6735);
and U7526 (N_7526,N_6350,N_6938);
nand U7527 (N_7527,N_6914,N_6325);
nand U7528 (N_7528,N_6419,N_6381);
or U7529 (N_7529,N_6854,N_6359);
nor U7530 (N_7530,N_6644,N_6045);
or U7531 (N_7531,N_6135,N_6108);
and U7532 (N_7532,N_6776,N_6499);
or U7533 (N_7533,N_6206,N_6687);
and U7534 (N_7534,N_6602,N_6498);
nand U7535 (N_7535,N_6179,N_6354);
nand U7536 (N_7536,N_6944,N_6093);
or U7537 (N_7537,N_6041,N_6522);
and U7538 (N_7538,N_6384,N_6907);
xnor U7539 (N_7539,N_6080,N_6443);
and U7540 (N_7540,N_6052,N_6988);
or U7541 (N_7541,N_6017,N_6211);
or U7542 (N_7542,N_6706,N_6500);
and U7543 (N_7543,N_6544,N_6080);
or U7544 (N_7544,N_6678,N_6026);
or U7545 (N_7545,N_6314,N_6710);
xor U7546 (N_7546,N_6090,N_6541);
xnor U7547 (N_7547,N_6865,N_6966);
xor U7548 (N_7548,N_6608,N_6878);
nand U7549 (N_7549,N_6251,N_6676);
nor U7550 (N_7550,N_6555,N_6491);
nand U7551 (N_7551,N_6330,N_6484);
xnor U7552 (N_7552,N_6404,N_6094);
nor U7553 (N_7553,N_6006,N_6179);
and U7554 (N_7554,N_6533,N_6462);
nor U7555 (N_7555,N_6751,N_6753);
nand U7556 (N_7556,N_6863,N_6519);
nor U7557 (N_7557,N_6238,N_6527);
xnor U7558 (N_7558,N_6814,N_6374);
xnor U7559 (N_7559,N_6080,N_6961);
and U7560 (N_7560,N_6245,N_6077);
xor U7561 (N_7561,N_6835,N_6662);
nor U7562 (N_7562,N_6838,N_6503);
nand U7563 (N_7563,N_6441,N_6167);
nor U7564 (N_7564,N_6976,N_6975);
xor U7565 (N_7565,N_6274,N_6460);
xnor U7566 (N_7566,N_6154,N_6422);
xnor U7567 (N_7567,N_6278,N_6886);
nand U7568 (N_7568,N_6789,N_6214);
nand U7569 (N_7569,N_6054,N_6866);
xnor U7570 (N_7570,N_6251,N_6555);
or U7571 (N_7571,N_6789,N_6731);
and U7572 (N_7572,N_6330,N_6655);
and U7573 (N_7573,N_6215,N_6095);
nand U7574 (N_7574,N_6108,N_6662);
xor U7575 (N_7575,N_6561,N_6032);
or U7576 (N_7576,N_6974,N_6949);
and U7577 (N_7577,N_6756,N_6238);
nand U7578 (N_7578,N_6161,N_6624);
and U7579 (N_7579,N_6104,N_6002);
nor U7580 (N_7580,N_6319,N_6033);
xnor U7581 (N_7581,N_6990,N_6494);
nand U7582 (N_7582,N_6043,N_6382);
nand U7583 (N_7583,N_6977,N_6445);
nor U7584 (N_7584,N_6456,N_6626);
or U7585 (N_7585,N_6249,N_6490);
or U7586 (N_7586,N_6503,N_6055);
or U7587 (N_7587,N_6489,N_6958);
or U7588 (N_7588,N_6360,N_6843);
nand U7589 (N_7589,N_6120,N_6365);
or U7590 (N_7590,N_6181,N_6471);
nor U7591 (N_7591,N_6729,N_6587);
nor U7592 (N_7592,N_6756,N_6549);
nor U7593 (N_7593,N_6127,N_6857);
nand U7594 (N_7594,N_6160,N_6103);
xnor U7595 (N_7595,N_6632,N_6192);
xnor U7596 (N_7596,N_6352,N_6519);
or U7597 (N_7597,N_6307,N_6016);
or U7598 (N_7598,N_6244,N_6329);
xnor U7599 (N_7599,N_6446,N_6111);
or U7600 (N_7600,N_6360,N_6836);
and U7601 (N_7601,N_6338,N_6322);
nand U7602 (N_7602,N_6008,N_6369);
xnor U7603 (N_7603,N_6504,N_6720);
nand U7604 (N_7604,N_6008,N_6586);
nand U7605 (N_7605,N_6646,N_6030);
or U7606 (N_7606,N_6028,N_6042);
or U7607 (N_7607,N_6482,N_6623);
xor U7608 (N_7608,N_6557,N_6670);
and U7609 (N_7609,N_6443,N_6274);
or U7610 (N_7610,N_6689,N_6150);
and U7611 (N_7611,N_6777,N_6860);
xor U7612 (N_7612,N_6390,N_6353);
xnor U7613 (N_7613,N_6285,N_6847);
or U7614 (N_7614,N_6102,N_6085);
xor U7615 (N_7615,N_6715,N_6518);
xnor U7616 (N_7616,N_6055,N_6876);
xor U7617 (N_7617,N_6253,N_6496);
xnor U7618 (N_7618,N_6443,N_6979);
or U7619 (N_7619,N_6485,N_6991);
nor U7620 (N_7620,N_6344,N_6618);
nor U7621 (N_7621,N_6115,N_6621);
xnor U7622 (N_7622,N_6560,N_6033);
and U7623 (N_7623,N_6860,N_6983);
xnor U7624 (N_7624,N_6038,N_6276);
xnor U7625 (N_7625,N_6356,N_6981);
nand U7626 (N_7626,N_6461,N_6805);
nor U7627 (N_7627,N_6899,N_6559);
nor U7628 (N_7628,N_6086,N_6651);
nor U7629 (N_7629,N_6520,N_6550);
xnor U7630 (N_7630,N_6030,N_6733);
xor U7631 (N_7631,N_6695,N_6888);
or U7632 (N_7632,N_6107,N_6693);
and U7633 (N_7633,N_6609,N_6488);
nor U7634 (N_7634,N_6375,N_6720);
or U7635 (N_7635,N_6116,N_6702);
nand U7636 (N_7636,N_6245,N_6624);
or U7637 (N_7637,N_6109,N_6107);
nand U7638 (N_7638,N_6915,N_6474);
or U7639 (N_7639,N_6404,N_6696);
xnor U7640 (N_7640,N_6717,N_6212);
and U7641 (N_7641,N_6103,N_6651);
or U7642 (N_7642,N_6972,N_6435);
and U7643 (N_7643,N_6986,N_6158);
nor U7644 (N_7644,N_6378,N_6402);
xnor U7645 (N_7645,N_6101,N_6901);
nor U7646 (N_7646,N_6573,N_6442);
and U7647 (N_7647,N_6617,N_6059);
nor U7648 (N_7648,N_6510,N_6061);
xor U7649 (N_7649,N_6295,N_6051);
and U7650 (N_7650,N_6875,N_6233);
nor U7651 (N_7651,N_6736,N_6849);
and U7652 (N_7652,N_6050,N_6314);
and U7653 (N_7653,N_6602,N_6973);
nor U7654 (N_7654,N_6920,N_6235);
xnor U7655 (N_7655,N_6288,N_6886);
or U7656 (N_7656,N_6786,N_6818);
nor U7657 (N_7657,N_6896,N_6029);
and U7658 (N_7658,N_6339,N_6689);
and U7659 (N_7659,N_6534,N_6671);
nand U7660 (N_7660,N_6825,N_6684);
nor U7661 (N_7661,N_6845,N_6933);
xor U7662 (N_7662,N_6110,N_6142);
xor U7663 (N_7663,N_6059,N_6636);
nor U7664 (N_7664,N_6932,N_6643);
and U7665 (N_7665,N_6612,N_6671);
nor U7666 (N_7666,N_6919,N_6105);
nand U7667 (N_7667,N_6786,N_6973);
xor U7668 (N_7668,N_6500,N_6480);
xor U7669 (N_7669,N_6050,N_6265);
nand U7670 (N_7670,N_6642,N_6886);
nand U7671 (N_7671,N_6957,N_6507);
xnor U7672 (N_7672,N_6483,N_6120);
nand U7673 (N_7673,N_6739,N_6837);
nand U7674 (N_7674,N_6579,N_6130);
and U7675 (N_7675,N_6885,N_6203);
and U7676 (N_7676,N_6417,N_6908);
xnor U7677 (N_7677,N_6888,N_6589);
and U7678 (N_7678,N_6275,N_6776);
or U7679 (N_7679,N_6880,N_6061);
nor U7680 (N_7680,N_6260,N_6545);
and U7681 (N_7681,N_6892,N_6125);
xor U7682 (N_7682,N_6488,N_6296);
and U7683 (N_7683,N_6311,N_6190);
or U7684 (N_7684,N_6797,N_6163);
nand U7685 (N_7685,N_6470,N_6558);
or U7686 (N_7686,N_6724,N_6650);
or U7687 (N_7687,N_6905,N_6892);
nand U7688 (N_7688,N_6865,N_6441);
xnor U7689 (N_7689,N_6304,N_6060);
nor U7690 (N_7690,N_6234,N_6232);
or U7691 (N_7691,N_6573,N_6149);
nor U7692 (N_7692,N_6330,N_6408);
nand U7693 (N_7693,N_6000,N_6652);
and U7694 (N_7694,N_6148,N_6577);
nor U7695 (N_7695,N_6010,N_6416);
xnor U7696 (N_7696,N_6881,N_6496);
xnor U7697 (N_7697,N_6689,N_6514);
nor U7698 (N_7698,N_6143,N_6439);
nand U7699 (N_7699,N_6587,N_6281);
or U7700 (N_7700,N_6795,N_6156);
nand U7701 (N_7701,N_6566,N_6785);
or U7702 (N_7702,N_6157,N_6362);
nand U7703 (N_7703,N_6711,N_6620);
nand U7704 (N_7704,N_6185,N_6394);
nand U7705 (N_7705,N_6289,N_6293);
xnor U7706 (N_7706,N_6182,N_6614);
nand U7707 (N_7707,N_6944,N_6150);
nand U7708 (N_7708,N_6856,N_6047);
xor U7709 (N_7709,N_6423,N_6299);
and U7710 (N_7710,N_6733,N_6545);
xnor U7711 (N_7711,N_6425,N_6310);
nor U7712 (N_7712,N_6019,N_6307);
and U7713 (N_7713,N_6035,N_6181);
and U7714 (N_7714,N_6243,N_6221);
and U7715 (N_7715,N_6119,N_6662);
or U7716 (N_7716,N_6811,N_6435);
nand U7717 (N_7717,N_6629,N_6269);
xnor U7718 (N_7718,N_6882,N_6592);
nand U7719 (N_7719,N_6754,N_6162);
xor U7720 (N_7720,N_6646,N_6425);
or U7721 (N_7721,N_6318,N_6959);
nand U7722 (N_7722,N_6867,N_6960);
nor U7723 (N_7723,N_6667,N_6869);
nor U7724 (N_7724,N_6248,N_6009);
nor U7725 (N_7725,N_6942,N_6091);
nor U7726 (N_7726,N_6491,N_6348);
and U7727 (N_7727,N_6904,N_6414);
or U7728 (N_7728,N_6413,N_6571);
nor U7729 (N_7729,N_6135,N_6853);
or U7730 (N_7730,N_6601,N_6296);
xor U7731 (N_7731,N_6846,N_6218);
xnor U7732 (N_7732,N_6933,N_6738);
or U7733 (N_7733,N_6338,N_6330);
xnor U7734 (N_7734,N_6940,N_6910);
or U7735 (N_7735,N_6229,N_6613);
xor U7736 (N_7736,N_6969,N_6689);
nand U7737 (N_7737,N_6190,N_6859);
or U7738 (N_7738,N_6806,N_6371);
nand U7739 (N_7739,N_6664,N_6432);
or U7740 (N_7740,N_6463,N_6781);
nor U7741 (N_7741,N_6365,N_6005);
nand U7742 (N_7742,N_6807,N_6138);
xnor U7743 (N_7743,N_6122,N_6863);
nand U7744 (N_7744,N_6389,N_6697);
and U7745 (N_7745,N_6701,N_6747);
or U7746 (N_7746,N_6465,N_6149);
and U7747 (N_7747,N_6375,N_6133);
and U7748 (N_7748,N_6461,N_6709);
or U7749 (N_7749,N_6687,N_6819);
nor U7750 (N_7750,N_6962,N_6416);
xor U7751 (N_7751,N_6716,N_6375);
nand U7752 (N_7752,N_6223,N_6507);
or U7753 (N_7753,N_6905,N_6586);
xor U7754 (N_7754,N_6201,N_6783);
nor U7755 (N_7755,N_6705,N_6081);
nand U7756 (N_7756,N_6316,N_6317);
or U7757 (N_7757,N_6489,N_6938);
nand U7758 (N_7758,N_6437,N_6892);
or U7759 (N_7759,N_6514,N_6194);
xnor U7760 (N_7760,N_6020,N_6372);
nand U7761 (N_7761,N_6802,N_6221);
xnor U7762 (N_7762,N_6519,N_6479);
nand U7763 (N_7763,N_6235,N_6557);
and U7764 (N_7764,N_6234,N_6585);
nand U7765 (N_7765,N_6480,N_6159);
nor U7766 (N_7766,N_6353,N_6406);
and U7767 (N_7767,N_6847,N_6446);
and U7768 (N_7768,N_6675,N_6403);
nor U7769 (N_7769,N_6939,N_6885);
nand U7770 (N_7770,N_6015,N_6075);
nand U7771 (N_7771,N_6716,N_6811);
xnor U7772 (N_7772,N_6948,N_6150);
nand U7773 (N_7773,N_6724,N_6900);
and U7774 (N_7774,N_6388,N_6105);
and U7775 (N_7775,N_6379,N_6862);
or U7776 (N_7776,N_6517,N_6592);
xnor U7777 (N_7777,N_6449,N_6463);
nand U7778 (N_7778,N_6118,N_6791);
nand U7779 (N_7779,N_6416,N_6644);
nand U7780 (N_7780,N_6190,N_6694);
nand U7781 (N_7781,N_6085,N_6799);
nand U7782 (N_7782,N_6098,N_6068);
and U7783 (N_7783,N_6341,N_6958);
nor U7784 (N_7784,N_6728,N_6321);
nand U7785 (N_7785,N_6611,N_6932);
xor U7786 (N_7786,N_6359,N_6528);
nand U7787 (N_7787,N_6276,N_6178);
nor U7788 (N_7788,N_6458,N_6930);
nand U7789 (N_7789,N_6421,N_6794);
nor U7790 (N_7790,N_6221,N_6416);
xnor U7791 (N_7791,N_6228,N_6943);
and U7792 (N_7792,N_6411,N_6783);
xor U7793 (N_7793,N_6221,N_6717);
and U7794 (N_7794,N_6815,N_6791);
or U7795 (N_7795,N_6858,N_6032);
nand U7796 (N_7796,N_6303,N_6236);
xnor U7797 (N_7797,N_6163,N_6556);
nand U7798 (N_7798,N_6601,N_6915);
nor U7799 (N_7799,N_6518,N_6574);
xor U7800 (N_7800,N_6263,N_6184);
nand U7801 (N_7801,N_6075,N_6956);
nor U7802 (N_7802,N_6163,N_6924);
nand U7803 (N_7803,N_6568,N_6155);
xnor U7804 (N_7804,N_6753,N_6094);
xnor U7805 (N_7805,N_6950,N_6356);
xnor U7806 (N_7806,N_6726,N_6391);
nor U7807 (N_7807,N_6014,N_6049);
and U7808 (N_7808,N_6123,N_6010);
nor U7809 (N_7809,N_6650,N_6905);
nand U7810 (N_7810,N_6016,N_6555);
or U7811 (N_7811,N_6108,N_6517);
or U7812 (N_7812,N_6011,N_6010);
xnor U7813 (N_7813,N_6119,N_6144);
nand U7814 (N_7814,N_6809,N_6754);
and U7815 (N_7815,N_6822,N_6492);
and U7816 (N_7816,N_6074,N_6037);
nor U7817 (N_7817,N_6150,N_6375);
xor U7818 (N_7818,N_6017,N_6014);
and U7819 (N_7819,N_6330,N_6694);
and U7820 (N_7820,N_6812,N_6148);
or U7821 (N_7821,N_6558,N_6641);
nand U7822 (N_7822,N_6879,N_6277);
nor U7823 (N_7823,N_6143,N_6252);
and U7824 (N_7824,N_6871,N_6885);
nor U7825 (N_7825,N_6197,N_6368);
or U7826 (N_7826,N_6576,N_6369);
xnor U7827 (N_7827,N_6796,N_6310);
nand U7828 (N_7828,N_6084,N_6584);
nor U7829 (N_7829,N_6552,N_6416);
nand U7830 (N_7830,N_6105,N_6562);
nand U7831 (N_7831,N_6318,N_6439);
nor U7832 (N_7832,N_6943,N_6462);
xor U7833 (N_7833,N_6917,N_6229);
nor U7834 (N_7834,N_6876,N_6796);
xor U7835 (N_7835,N_6615,N_6101);
or U7836 (N_7836,N_6516,N_6298);
and U7837 (N_7837,N_6677,N_6667);
xnor U7838 (N_7838,N_6478,N_6491);
and U7839 (N_7839,N_6965,N_6204);
xor U7840 (N_7840,N_6017,N_6196);
or U7841 (N_7841,N_6301,N_6564);
nor U7842 (N_7842,N_6160,N_6790);
or U7843 (N_7843,N_6672,N_6620);
or U7844 (N_7844,N_6116,N_6951);
nor U7845 (N_7845,N_6288,N_6003);
nor U7846 (N_7846,N_6830,N_6365);
nand U7847 (N_7847,N_6660,N_6089);
nor U7848 (N_7848,N_6172,N_6254);
nand U7849 (N_7849,N_6805,N_6913);
xor U7850 (N_7850,N_6237,N_6798);
nand U7851 (N_7851,N_6109,N_6853);
nand U7852 (N_7852,N_6216,N_6947);
nand U7853 (N_7853,N_6958,N_6535);
and U7854 (N_7854,N_6377,N_6283);
or U7855 (N_7855,N_6310,N_6269);
nor U7856 (N_7856,N_6096,N_6044);
xnor U7857 (N_7857,N_6958,N_6121);
xnor U7858 (N_7858,N_6380,N_6419);
nor U7859 (N_7859,N_6743,N_6366);
nand U7860 (N_7860,N_6629,N_6156);
and U7861 (N_7861,N_6156,N_6402);
nand U7862 (N_7862,N_6458,N_6030);
nor U7863 (N_7863,N_6834,N_6275);
xnor U7864 (N_7864,N_6982,N_6628);
nand U7865 (N_7865,N_6675,N_6674);
and U7866 (N_7866,N_6777,N_6243);
nand U7867 (N_7867,N_6484,N_6101);
and U7868 (N_7868,N_6433,N_6550);
nand U7869 (N_7869,N_6116,N_6165);
xor U7870 (N_7870,N_6446,N_6692);
nand U7871 (N_7871,N_6660,N_6610);
and U7872 (N_7872,N_6972,N_6644);
or U7873 (N_7873,N_6753,N_6370);
and U7874 (N_7874,N_6424,N_6537);
nand U7875 (N_7875,N_6737,N_6053);
or U7876 (N_7876,N_6841,N_6773);
or U7877 (N_7877,N_6658,N_6735);
nand U7878 (N_7878,N_6205,N_6316);
or U7879 (N_7879,N_6991,N_6871);
nand U7880 (N_7880,N_6157,N_6046);
nand U7881 (N_7881,N_6947,N_6432);
nor U7882 (N_7882,N_6281,N_6870);
nor U7883 (N_7883,N_6398,N_6377);
xnor U7884 (N_7884,N_6110,N_6137);
xor U7885 (N_7885,N_6300,N_6454);
and U7886 (N_7886,N_6710,N_6019);
nand U7887 (N_7887,N_6424,N_6251);
or U7888 (N_7888,N_6775,N_6424);
or U7889 (N_7889,N_6521,N_6491);
xnor U7890 (N_7890,N_6311,N_6336);
nand U7891 (N_7891,N_6697,N_6494);
nor U7892 (N_7892,N_6940,N_6317);
and U7893 (N_7893,N_6268,N_6691);
nand U7894 (N_7894,N_6025,N_6772);
and U7895 (N_7895,N_6725,N_6656);
and U7896 (N_7896,N_6661,N_6782);
nor U7897 (N_7897,N_6418,N_6121);
nand U7898 (N_7898,N_6769,N_6244);
nand U7899 (N_7899,N_6479,N_6129);
or U7900 (N_7900,N_6920,N_6152);
or U7901 (N_7901,N_6843,N_6219);
nor U7902 (N_7902,N_6585,N_6598);
nor U7903 (N_7903,N_6447,N_6390);
nand U7904 (N_7904,N_6098,N_6234);
nor U7905 (N_7905,N_6485,N_6630);
nor U7906 (N_7906,N_6550,N_6272);
and U7907 (N_7907,N_6334,N_6771);
or U7908 (N_7908,N_6555,N_6483);
xor U7909 (N_7909,N_6840,N_6912);
nand U7910 (N_7910,N_6675,N_6894);
or U7911 (N_7911,N_6449,N_6745);
or U7912 (N_7912,N_6073,N_6485);
nor U7913 (N_7913,N_6519,N_6501);
xor U7914 (N_7914,N_6690,N_6653);
and U7915 (N_7915,N_6182,N_6958);
or U7916 (N_7916,N_6122,N_6795);
and U7917 (N_7917,N_6994,N_6272);
or U7918 (N_7918,N_6943,N_6924);
and U7919 (N_7919,N_6055,N_6519);
or U7920 (N_7920,N_6041,N_6743);
or U7921 (N_7921,N_6878,N_6205);
nand U7922 (N_7922,N_6200,N_6287);
nor U7923 (N_7923,N_6960,N_6645);
and U7924 (N_7924,N_6952,N_6470);
or U7925 (N_7925,N_6266,N_6217);
or U7926 (N_7926,N_6172,N_6341);
and U7927 (N_7927,N_6031,N_6110);
nor U7928 (N_7928,N_6478,N_6670);
xor U7929 (N_7929,N_6727,N_6648);
and U7930 (N_7930,N_6261,N_6647);
nor U7931 (N_7931,N_6528,N_6220);
nor U7932 (N_7932,N_6112,N_6514);
xor U7933 (N_7933,N_6693,N_6519);
nand U7934 (N_7934,N_6496,N_6324);
or U7935 (N_7935,N_6895,N_6622);
nand U7936 (N_7936,N_6587,N_6852);
or U7937 (N_7937,N_6852,N_6115);
nor U7938 (N_7938,N_6019,N_6145);
nor U7939 (N_7939,N_6249,N_6315);
nand U7940 (N_7940,N_6991,N_6094);
xor U7941 (N_7941,N_6582,N_6135);
nor U7942 (N_7942,N_6243,N_6495);
nor U7943 (N_7943,N_6908,N_6775);
and U7944 (N_7944,N_6403,N_6762);
nand U7945 (N_7945,N_6600,N_6237);
nand U7946 (N_7946,N_6484,N_6691);
xor U7947 (N_7947,N_6685,N_6723);
nand U7948 (N_7948,N_6429,N_6718);
nand U7949 (N_7949,N_6080,N_6532);
or U7950 (N_7950,N_6198,N_6656);
xnor U7951 (N_7951,N_6051,N_6908);
nor U7952 (N_7952,N_6937,N_6158);
nand U7953 (N_7953,N_6324,N_6915);
nand U7954 (N_7954,N_6549,N_6939);
xnor U7955 (N_7955,N_6613,N_6549);
xnor U7956 (N_7956,N_6589,N_6653);
xnor U7957 (N_7957,N_6489,N_6068);
and U7958 (N_7958,N_6232,N_6085);
or U7959 (N_7959,N_6043,N_6141);
nor U7960 (N_7960,N_6620,N_6481);
nor U7961 (N_7961,N_6614,N_6279);
and U7962 (N_7962,N_6546,N_6181);
nor U7963 (N_7963,N_6243,N_6384);
nor U7964 (N_7964,N_6222,N_6871);
or U7965 (N_7965,N_6053,N_6929);
nor U7966 (N_7966,N_6962,N_6052);
xor U7967 (N_7967,N_6389,N_6965);
xnor U7968 (N_7968,N_6027,N_6969);
xor U7969 (N_7969,N_6627,N_6571);
xnor U7970 (N_7970,N_6603,N_6824);
or U7971 (N_7971,N_6556,N_6743);
and U7972 (N_7972,N_6214,N_6382);
xor U7973 (N_7973,N_6122,N_6062);
nand U7974 (N_7974,N_6678,N_6901);
or U7975 (N_7975,N_6908,N_6646);
nand U7976 (N_7976,N_6539,N_6658);
nor U7977 (N_7977,N_6772,N_6869);
xor U7978 (N_7978,N_6387,N_6746);
nor U7979 (N_7979,N_6674,N_6965);
nand U7980 (N_7980,N_6534,N_6453);
or U7981 (N_7981,N_6435,N_6400);
nand U7982 (N_7982,N_6808,N_6381);
nand U7983 (N_7983,N_6850,N_6745);
or U7984 (N_7984,N_6333,N_6889);
nor U7985 (N_7985,N_6711,N_6982);
and U7986 (N_7986,N_6379,N_6423);
nand U7987 (N_7987,N_6659,N_6119);
or U7988 (N_7988,N_6490,N_6087);
or U7989 (N_7989,N_6044,N_6736);
nand U7990 (N_7990,N_6900,N_6107);
or U7991 (N_7991,N_6138,N_6801);
nor U7992 (N_7992,N_6911,N_6334);
nor U7993 (N_7993,N_6999,N_6760);
and U7994 (N_7994,N_6897,N_6857);
nand U7995 (N_7995,N_6649,N_6530);
and U7996 (N_7996,N_6722,N_6247);
xor U7997 (N_7997,N_6218,N_6775);
and U7998 (N_7998,N_6881,N_6628);
and U7999 (N_7999,N_6366,N_6203);
nor U8000 (N_8000,N_7912,N_7710);
or U8001 (N_8001,N_7743,N_7344);
nor U8002 (N_8002,N_7893,N_7574);
and U8003 (N_8003,N_7214,N_7934);
xnor U8004 (N_8004,N_7484,N_7654);
xor U8005 (N_8005,N_7719,N_7013);
and U8006 (N_8006,N_7303,N_7607);
nor U8007 (N_8007,N_7935,N_7972);
and U8008 (N_8008,N_7491,N_7429);
or U8009 (N_8009,N_7040,N_7694);
xnor U8010 (N_8010,N_7414,N_7921);
nor U8011 (N_8011,N_7968,N_7843);
nor U8012 (N_8012,N_7631,N_7708);
or U8013 (N_8013,N_7307,N_7068);
or U8014 (N_8014,N_7752,N_7197);
and U8015 (N_8015,N_7176,N_7531);
or U8016 (N_8016,N_7350,N_7786);
and U8017 (N_8017,N_7449,N_7021);
xor U8018 (N_8018,N_7092,N_7979);
xnor U8019 (N_8019,N_7846,N_7385);
or U8020 (N_8020,N_7583,N_7560);
nor U8021 (N_8021,N_7777,N_7993);
xnor U8022 (N_8022,N_7219,N_7593);
and U8023 (N_8023,N_7137,N_7440);
or U8024 (N_8024,N_7754,N_7558);
and U8025 (N_8025,N_7139,N_7376);
xnor U8026 (N_8026,N_7693,N_7578);
xnor U8027 (N_8027,N_7923,N_7148);
nand U8028 (N_8028,N_7806,N_7788);
nor U8029 (N_8029,N_7102,N_7157);
xnor U8030 (N_8030,N_7158,N_7546);
nand U8031 (N_8031,N_7625,N_7173);
nand U8032 (N_8032,N_7728,N_7761);
xor U8033 (N_8033,N_7916,N_7868);
nand U8034 (N_8034,N_7146,N_7817);
or U8035 (N_8035,N_7318,N_7741);
or U8036 (N_8036,N_7876,N_7585);
nor U8037 (N_8037,N_7589,N_7084);
nor U8038 (N_8038,N_7857,N_7835);
nand U8039 (N_8039,N_7361,N_7099);
and U8040 (N_8040,N_7644,N_7841);
xor U8041 (N_8041,N_7265,N_7462);
or U8042 (N_8042,N_7579,N_7861);
xor U8043 (N_8043,N_7825,N_7779);
xor U8044 (N_8044,N_7842,N_7679);
or U8045 (N_8045,N_7490,N_7272);
and U8046 (N_8046,N_7186,N_7360);
nand U8047 (N_8047,N_7443,N_7571);
and U8048 (N_8048,N_7594,N_7246);
nor U8049 (N_8049,N_7727,N_7367);
xor U8050 (N_8050,N_7200,N_7280);
nand U8051 (N_8051,N_7346,N_7918);
nand U8052 (N_8052,N_7080,N_7283);
nor U8053 (N_8053,N_7333,N_7807);
nand U8054 (N_8054,N_7420,N_7438);
or U8055 (N_8055,N_7172,N_7536);
and U8056 (N_8056,N_7793,N_7486);
nor U8057 (N_8057,N_7010,N_7960);
or U8058 (N_8058,N_7480,N_7948);
nor U8059 (N_8059,N_7195,N_7522);
nor U8060 (N_8060,N_7833,N_7389);
or U8061 (N_8061,N_7335,N_7903);
or U8062 (N_8062,N_7682,N_7969);
nor U8063 (N_8063,N_7014,N_7117);
or U8064 (N_8064,N_7590,N_7596);
nor U8065 (N_8065,N_7991,N_7945);
nor U8066 (N_8066,N_7009,N_7949);
or U8067 (N_8067,N_7856,N_7669);
xnor U8068 (N_8068,N_7025,N_7123);
nand U8069 (N_8069,N_7844,N_7377);
xnor U8070 (N_8070,N_7416,N_7362);
nand U8071 (N_8071,N_7340,N_7987);
and U8072 (N_8072,N_7038,N_7811);
or U8073 (N_8073,N_7624,N_7971);
nor U8074 (N_8074,N_7943,N_7826);
nand U8075 (N_8075,N_7629,N_7218);
or U8076 (N_8076,N_7904,N_7323);
or U8077 (N_8077,N_7666,N_7412);
nor U8078 (N_8078,N_7518,N_7919);
nor U8079 (N_8079,N_7610,N_7430);
or U8080 (N_8080,N_7959,N_7999);
nand U8081 (N_8081,N_7037,N_7920);
nand U8082 (N_8082,N_7875,N_7707);
or U8083 (N_8083,N_7834,N_7519);
nor U8084 (N_8084,N_7848,N_7715);
and U8085 (N_8085,N_7862,N_7096);
xor U8086 (N_8086,N_7295,N_7570);
and U8087 (N_8087,N_7279,N_7633);
and U8088 (N_8088,N_7882,N_7561);
and U8089 (N_8089,N_7789,N_7300);
and U8090 (N_8090,N_7368,N_7824);
nand U8091 (N_8091,N_7608,N_7083);
xor U8092 (N_8092,N_7077,N_7802);
or U8093 (N_8093,N_7983,N_7758);
or U8094 (N_8094,N_7622,N_7114);
or U8095 (N_8095,N_7641,N_7392);
and U8096 (N_8096,N_7456,N_7426);
nor U8097 (N_8097,N_7100,N_7183);
nor U8098 (N_8098,N_7515,N_7512);
xor U8099 (N_8099,N_7820,N_7556);
or U8100 (N_8100,N_7905,N_7144);
or U8101 (N_8101,N_7963,N_7302);
or U8102 (N_8102,N_7212,N_7384);
nand U8103 (N_8103,N_7529,N_7615);
nand U8104 (N_8104,N_7093,N_7374);
nand U8105 (N_8105,N_7263,N_7926);
xor U8106 (N_8106,N_7364,N_7446);
nand U8107 (N_8107,N_7822,N_7568);
nor U8108 (N_8108,N_7643,N_7181);
xor U8109 (N_8109,N_7165,N_7836);
and U8110 (N_8110,N_7725,N_7626);
xnor U8111 (N_8111,N_7526,N_7692);
and U8112 (N_8112,N_7771,N_7140);
nor U8113 (N_8113,N_7073,N_7899);
nor U8114 (N_8114,N_7517,N_7680);
or U8115 (N_8115,N_7499,N_7854);
nand U8116 (N_8116,N_7913,N_7477);
or U8117 (N_8117,N_7598,N_7026);
nand U8118 (N_8118,N_7248,N_7830);
xnor U8119 (N_8119,N_7717,N_7485);
nand U8120 (N_8120,N_7797,N_7961);
and U8121 (N_8121,N_7884,N_7036);
or U8122 (N_8122,N_7595,N_7940);
nand U8123 (N_8123,N_7506,N_7074);
or U8124 (N_8124,N_7223,N_7031);
nand U8125 (N_8125,N_7434,N_7896);
nand U8126 (N_8126,N_7188,N_7986);
and U8127 (N_8127,N_7316,N_7023);
nand U8128 (N_8128,N_7270,N_7553);
nor U8129 (N_8129,N_7163,N_7184);
nand U8130 (N_8130,N_7070,N_7652);
nand U8131 (N_8131,N_7706,N_7932);
and U8132 (N_8132,N_7818,N_7770);
nand U8133 (N_8133,N_7674,N_7827);
and U8134 (N_8134,N_7287,N_7034);
nor U8135 (N_8135,N_7386,N_7247);
nand U8136 (N_8136,N_7317,N_7466);
xor U8137 (N_8137,N_7790,N_7325);
or U8138 (N_8138,N_7152,N_7394);
and U8139 (N_8139,N_7125,N_7798);
nand U8140 (N_8140,N_7273,N_7575);
and U8141 (N_8141,N_7673,N_7513);
nand U8142 (N_8142,N_7730,N_7768);
xnor U8143 (N_8143,N_7939,N_7813);
or U8144 (N_8144,N_7402,N_7193);
xor U8145 (N_8145,N_7103,N_7775);
nand U8146 (N_8146,N_7609,N_7461);
xnor U8147 (N_8147,N_7177,N_7716);
nand U8148 (N_8148,N_7930,N_7950);
nor U8149 (N_8149,N_7505,N_7168);
and U8150 (N_8150,N_7227,N_7329);
xor U8151 (N_8151,N_7498,N_7545);
xor U8152 (N_8152,N_7003,N_7520);
and U8153 (N_8153,N_7343,N_7105);
xnor U8154 (N_8154,N_7621,N_7753);
xor U8155 (N_8155,N_7524,N_7053);
or U8156 (N_8156,N_7627,N_7783);
and U8157 (N_8157,N_7823,N_7019);
and U8158 (N_8158,N_7723,N_7210);
nor U8159 (N_8159,N_7653,N_7142);
nand U8160 (N_8160,N_7638,N_7665);
nor U8161 (N_8161,N_7981,N_7839);
and U8162 (N_8162,N_7891,N_7687);
nor U8163 (N_8163,N_7769,N_7762);
nor U8164 (N_8164,N_7550,N_7071);
or U8165 (N_8165,N_7668,N_7164);
xnor U8166 (N_8166,N_7879,N_7632);
nand U8167 (N_8167,N_7355,N_7736);
xnor U8168 (N_8168,N_7390,N_7778);
and U8169 (N_8169,N_7130,N_7689);
nand U8170 (N_8170,N_7847,N_7145);
nor U8171 (N_8171,N_7703,N_7591);
xor U8172 (N_8172,N_7814,N_7190);
nand U8173 (N_8173,N_7659,N_7058);
xnor U8174 (N_8174,N_7348,N_7015);
nand U8175 (N_8175,N_7809,N_7675);
or U8176 (N_8176,N_7056,N_7109);
xnor U8177 (N_8177,N_7500,N_7994);
nand U8178 (N_8178,N_7870,N_7584);
nor U8179 (N_8179,N_7880,N_7312);
xnor U8180 (N_8180,N_7564,N_7975);
nand U8181 (N_8181,N_7604,N_7050);
and U8182 (N_8182,N_7088,N_7713);
and U8183 (N_8183,N_7525,N_7027);
or U8184 (N_8184,N_7751,N_7455);
nand U8185 (N_8185,N_7264,N_7042);
nand U8186 (N_8186,N_7510,N_7759);
and U8187 (N_8187,N_7366,N_7239);
nand U8188 (N_8188,N_7309,N_7132);
nand U8189 (N_8189,N_7127,N_7320);
nand U8190 (N_8190,N_7378,N_7143);
nor U8191 (N_8191,N_7840,N_7562);
and U8192 (N_8192,N_7001,N_7232);
or U8193 (N_8193,N_7586,N_7742);
xor U8194 (N_8194,N_7924,N_7557);
nor U8195 (N_8195,N_7268,N_7469);
nor U8196 (N_8196,N_7315,N_7577);
nor U8197 (N_8197,N_7773,N_7634);
nand U8198 (N_8198,N_7569,N_7944);
xor U8199 (N_8199,N_7081,N_7305);
xnor U8200 (N_8200,N_7411,N_7258);
or U8201 (N_8201,N_7685,N_7191);
or U8202 (N_8202,N_7055,N_7982);
and U8203 (N_8203,N_7511,N_7954);
xnor U8204 (N_8204,N_7199,N_7837);
or U8205 (N_8205,N_7478,N_7128);
nand U8206 (N_8206,N_7538,N_7418);
nand U8207 (N_8207,N_7878,N_7410);
and U8208 (N_8208,N_7444,N_7110);
nand U8209 (N_8209,N_7639,N_7792);
xnor U8210 (N_8210,N_7765,N_7358);
and U8211 (N_8211,N_7863,N_7097);
nor U8212 (N_8212,N_7059,N_7205);
and U8213 (N_8213,N_7953,N_7403);
xor U8214 (N_8214,N_7032,N_7787);
or U8215 (N_8215,N_7721,N_7445);
nor U8216 (N_8216,N_7179,N_7463);
or U8217 (N_8217,N_7697,N_7688);
xor U8218 (N_8218,N_7234,N_7311);
nand U8219 (N_8219,N_7475,N_7967);
nand U8220 (N_8220,N_7964,N_7582);
xnor U8221 (N_8221,N_7767,N_7453);
nor U8222 (N_8222,N_7175,N_7541);
nand U8223 (N_8223,N_7829,N_7698);
and U8224 (N_8224,N_7852,N_7061);
nand U8225 (N_8225,N_7313,N_7565);
or U8226 (N_8226,N_7649,N_7098);
or U8227 (N_8227,N_7532,N_7873);
or U8228 (N_8228,N_7763,N_7664);
xor U8229 (N_8229,N_7047,N_7020);
nor U8230 (N_8230,N_7696,N_7756);
nand U8231 (N_8231,N_7187,N_7845);
xnor U8232 (N_8232,N_7211,N_7141);
xor U8233 (N_8233,N_7241,N_7616);
and U8234 (N_8234,N_7508,N_7597);
or U8235 (N_8235,N_7911,N_7867);
nor U8236 (N_8236,N_7111,N_7496);
nand U8237 (N_8237,N_7889,N_7201);
and U8238 (N_8238,N_7740,N_7149);
nor U8239 (N_8239,N_7230,N_7005);
nand U8240 (N_8240,N_7774,N_7894);
or U8241 (N_8241,N_7243,N_7832);
xor U8242 (N_8242,N_7337,N_7611);
or U8243 (N_8243,N_7980,N_7018);
xor U8244 (N_8244,N_7467,N_7291);
or U8245 (N_8245,N_7540,N_7066);
nand U8246 (N_8246,N_7587,N_7474);
or U8247 (N_8247,N_7060,N_7860);
and U8248 (N_8248,N_7720,N_7459);
nand U8249 (N_8249,N_7489,N_7617);
or U8250 (N_8250,N_7075,N_7108);
nor U8251 (N_8251,N_7162,N_7890);
or U8252 (N_8252,N_7791,N_7252);
nand U8253 (N_8253,N_7865,N_7086);
or U8254 (N_8254,N_7220,N_7831);
nand U8255 (N_8255,N_7925,N_7233);
nor U8256 (N_8256,N_7691,N_7282);
xnor U8257 (N_8257,N_7888,N_7330);
nand U8258 (N_8258,N_7734,N_7784);
xnor U8259 (N_8259,N_7922,N_7189);
or U8260 (N_8260,N_7242,N_7749);
nor U8261 (N_8261,N_7819,N_7699);
and U8262 (N_8262,N_7859,N_7648);
nor U8263 (N_8263,N_7079,N_7992);
and U8264 (N_8264,N_7998,N_7549);
and U8265 (N_8265,N_7450,N_7274);
xnor U8266 (N_8266,N_7933,N_7702);
or U8267 (N_8267,N_7421,N_7286);
or U8268 (N_8268,N_7357,N_7222);
nor U8269 (N_8269,N_7359,N_7657);
nor U8270 (N_8270,N_7471,N_7166);
nand U8271 (N_8271,N_7332,N_7507);
nor U8272 (N_8272,N_7231,N_7726);
or U8273 (N_8273,N_7988,N_7129);
or U8274 (N_8274,N_7082,N_7441);
xnor U8275 (N_8275,N_7373,N_7855);
nand U8276 (N_8276,N_7238,N_7658);
and U8277 (N_8277,N_7795,N_7677);
and U8278 (N_8278,N_7120,N_7400);
or U8279 (N_8279,N_7048,N_7937);
nand U8280 (N_8280,N_7245,N_7600);
nor U8281 (N_8281,N_7978,N_7345);
nor U8282 (N_8282,N_7683,N_7324);
nand U8283 (N_8283,N_7602,N_7976);
nand U8284 (N_8284,N_7612,N_7004);
xor U8285 (N_8285,N_7057,N_7065);
or U8286 (N_8286,N_7308,N_7554);
or U8287 (N_8287,N_7016,N_7711);
or U8288 (N_8288,N_7909,N_7559);
nor U8289 (N_8289,N_7801,N_7472);
nor U8290 (N_8290,N_7116,N_7735);
nor U8291 (N_8291,N_7748,N_7393);
or U8292 (N_8292,N_7662,N_7285);
and U8293 (N_8293,N_7365,N_7008);
and U8294 (N_8294,N_7872,N_7113);
or U8295 (N_8295,N_7161,N_7482);
or U8296 (N_8296,N_7528,N_7637);
xor U8297 (N_8297,N_7433,N_7618);
xor U8298 (N_8298,N_7941,N_7134);
or U8299 (N_8299,N_7701,N_7521);
nand U8300 (N_8300,N_7849,N_7257);
nand U8301 (N_8301,N_7704,N_7527);
and U8302 (N_8302,N_7647,N_7497);
nor U8303 (N_8303,N_7372,N_7799);
or U8304 (N_8304,N_7864,N_7995);
xnor U8305 (N_8305,N_7990,N_7881);
or U8306 (N_8306,N_7606,N_7722);
and U8307 (N_8307,N_7292,N_7928);
or U8308 (N_8308,N_7178,N_7089);
nor U8309 (N_8309,N_7906,N_7603);
nand U8310 (N_8310,N_7504,N_7196);
or U8311 (N_8311,N_7493,N_7551);
nand U8312 (N_8312,N_7382,N_7858);
xnor U8313 (N_8313,N_7260,N_7171);
xor U8314 (N_8314,N_7347,N_7821);
xnor U8315 (N_8315,N_7984,N_7996);
and U8316 (N_8316,N_7383,N_7650);
xor U8317 (N_8317,N_7085,N_7000);
or U8318 (N_8318,N_7427,N_7215);
and U8319 (N_8319,N_7428,N_7956);
nand U8320 (N_8320,N_7002,N_7319);
nand U8321 (N_8321,N_7709,N_7090);
and U8322 (N_8322,N_7126,N_7236);
or U8323 (N_8323,N_7576,N_7483);
or U8324 (N_8324,N_7588,N_7503);
xor U8325 (N_8325,N_7022,N_7293);
xnor U8326 (N_8326,N_7501,N_7297);
nand U8327 (N_8327,N_7087,N_7962);
nor U8328 (N_8328,N_7447,N_7388);
nor U8329 (N_8329,N_7910,N_7850);
or U8330 (N_8330,N_7572,N_7476);
or U8331 (N_8331,N_7072,N_7892);
xnor U8332 (N_8332,N_7237,N_7439);
or U8333 (N_8333,N_7636,N_7700);
nor U8334 (N_8334,N_7613,N_7874);
xor U8335 (N_8335,N_7401,N_7045);
or U8336 (N_8336,N_7555,N_7757);
nand U8337 (N_8337,N_7314,N_7064);
nor U8338 (N_8338,N_7473,N_7192);
and U8339 (N_8339,N_7076,N_7250);
nor U8340 (N_8340,N_7049,N_7249);
nor U8341 (N_8341,N_7544,N_7328);
nand U8342 (N_8342,N_7327,N_7408);
nor U8343 (N_8343,N_7776,N_7067);
or U8344 (N_8344,N_7661,N_7255);
and U8345 (N_8345,N_7468,N_7422);
nand U8346 (N_8346,N_7259,N_7380);
and U8347 (N_8347,N_7733,N_7457);
nor U8348 (N_8348,N_7407,N_7448);
nand U8349 (N_8349,N_7646,N_7321);
nand U8350 (N_8350,N_7542,N_7623);
xor U8351 (N_8351,N_7039,N_7567);
or U8352 (N_8352,N_7914,N_7046);
and U8353 (N_8353,N_7017,N_7052);
or U8354 (N_8354,N_7695,N_7078);
nor U8355 (N_8355,N_7262,N_7464);
or U8356 (N_8356,N_7766,N_7780);
nand U8357 (N_8357,N_7011,N_7573);
nand U8358 (N_8358,N_7240,N_7122);
xor U8359 (N_8359,N_7887,N_7395);
nand U8360 (N_8360,N_7620,N_7266);
nor U8361 (N_8361,N_7399,N_7352);
nand U8362 (N_8362,N_7901,N_7041);
nor U8363 (N_8363,N_7739,N_7206);
or U8364 (N_8364,N_7442,N_7261);
nor U8365 (N_8365,N_7946,N_7198);
xnor U8366 (N_8366,N_7533,N_7277);
and U8367 (N_8367,N_7853,N_7229);
nand U8368 (N_8368,N_7936,N_7136);
or U8369 (N_8369,N_7288,N_7547);
nor U8370 (N_8370,N_7724,N_7481);
nor U8371 (N_8371,N_7101,N_7686);
or U8372 (N_8372,N_7488,N_7417);
xnor U8373 (N_8373,N_7470,N_7580);
nand U8374 (N_8374,N_7043,N_7396);
nand U8375 (N_8375,N_7539,N_7131);
and U8376 (N_8376,N_7269,N_7024);
or U8377 (N_8377,N_7885,N_7782);
or U8378 (N_8378,N_7290,N_7718);
nor U8379 (N_8379,N_7635,N_7363);
and U8380 (N_8380,N_7684,N_7007);
or U8381 (N_8381,N_7672,N_7118);
nor U8382 (N_8382,N_7494,N_7299);
xor U8383 (N_8383,N_7938,N_7424);
xor U8384 (N_8384,N_7929,N_7244);
xnor U8385 (N_8385,N_7534,N_7628);
xor U8386 (N_8386,N_7224,N_7465);
or U8387 (N_8387,N_7851,N_7804);
xor U8388 (N_8388,N_7738,N_7810);
and U8389 (N_8389,N_7681,N_7895);
nor U8390 (N_8390,N_7745,N_7454);
xor U8391 (N_8391,N_7062,N_7640);
xnor U8392 (N_8392,N_7326,N_7115);
and U8393 (N_8393,N_7182,N_7712);
nand U8394 (N_8394,N_7398,N_7035);
nand U8395 (N_8395,N_7902,N_7369);
or U8396 (N_8396,N_7705,N_7535);
or U8397 (N_8397,N_7747,N_7306);
xor U8398 (N_8398,N_7581,N_7296);
or U8399 (N_8399,N_7957,N_7808);
or U8400 (N_8400,N_7729,N_7331);
xor U8401 (N_8401,N_7391,N_7235);
and U8402 (N_8402,N_7871,N_7927);
xor U8403 (N_8403,N_7732,N_7977);
and U8404 (N_8404,N_7760,N_7942);
and U8405 (N_8405,N_7275,N_7051);
or U8406 (N_8406,N_7397,N_7671);
xor U8407 (N_8407,N_7154,N_7974);
nor U8408 (N_8408,N_7304,N_7800);
nor U8409 (N_8409,N_7431,N_7155);
and U8410 (N_8410,N_7805,N_7054);
xor U8411 (N_8411,N_7356,N_7530);
nor U8412 (N_8412,N_7256,N_7351);
nor U8413 (N_8413,N_7663,N_7714);
nand U8414 (N_8414,N_7966,N_7651);
and U8415 (N_8415,N_7253,N_7271);
nor U8416 (N_8416,N_7028,N_7915);
xnor U8417 (N_8417,N_7135,N_7336);
and U8418 (N_8418,N_7970,N_7112);
nand U8419 (N_8419,N_7342,N_7353);
nand U8420 (N_8420,N_7869,N_7012);
or U8421 (N_8421,N_7294,N_7413);
or U8422 (N_8422,N_7217,N_7204);
nor U8423 (N_8423,N_7044,N_7772);
nor U8424 (N_8424,N_7094,N_7678);
xnor U8425 (N_8425,N_7670,N_7281);
nor U8426 (N_8426,N_7931,N_7642);
xor U8427 (N_8427,N_7796,N_7655);
xor U8428 (N_8428,N_7592,N_7106);
or U8429 (N_8429,N_7301,N_7381);
and U8430 (N_8430,N_7194,N_7310);
or U8431 (N_8431,N_7552,N_7947);
or U8432 (N_8432,N_7029,N_7121);
and U8433 (N_8433,N_7908,N_7514);
nor U8434 (N_8434,N_7156,N_7322);
nor U8435 (N_8435,N_7150,N_7209);
xor U8436 (N_8436,N_7185,N_7803);
nand U8437 (N_8437,N_7289,N_7660);
and U8438 (N_8438,N_7254,N_7815);
or U8439 (N_8439,N_7460,N_7746);
or U8440 (N_8440,N_7371,N_7151);
xnor U8441 (N_8441,N_7605,N_7202);
nor U8442 (N_8442,N_7812,N_7965);
xor U8443 (N_8443,N_7989,N_7744);
nand U8444 (N_8444,N_7159,N_7069);
nor U8445 (N_8445,N_7458,N_7278);
xnor U8446 (N_8446,N_7415,N_7897);
nand U8447 (N_8447,N_7951,N_7133);
or U8448 (N_8448,N_7731,N_7425);
nor U8449 (N_8449,N_7958,N_7794);
nor U8450 (N_8450,N_7170,N_7107);
or U8451 (N_8451,N_7406,N_7409);
and U8452 (N_8452,N_7341,N_7404);
and U8453 (N_8453,N_7599,N_7630);
nor U8454 (N_8454,N_7267,N_7091);
nor U8455 (N_8455,N_7656,N_7543);
xor U8456 (N_8456,N_7667,N_7276);
and U8457 (N_8457,N_7437,N_7917);
nor U8458 (N_8458,N_7221,N_7284);
or U8459 (N_8459,N_7423,N_7203);
nor U8460 (N_8460,N_7354,N_7523);
and U8461 (N_8461,N_7785,N_7479);
nand U8462 (N_8462,N_7838,N_7492);
and U8463 (N_8463,N_7379,N_7160);
or U8464 (N_8464,N_7452,N_7339);
nor U8465 (N_8465,N_7338,N_7169);
or U8466 (N_8466,N_7566,N_7030);
nand U8467 (N_8467,N_7750,N_7006);
or U8468 (N_8468,N_7167,N_7153);
nand U8469 (N_8469,N_7095,N_7755);
or U8470 (N_8470,N_7487,N_7370);
nor U8471 (N_8471,N_7451,N_7251);
nand U8472 (N_8472,N_7955,N_7298);
nand U8473 (N_8473,N_7866,N_7563);
and U8474 (N_8474,N_7645,N_7207);
or U8475 (N_8475,N_7228,N_7781);
and U8476 (N_8476,N_7334,N_7509);
or U8477 (N_8477,N_7676,N_7213);
nor U8478 (N_8478,N_7537,N_7119);
xor U8479 (N_8479,N_7816,N_7877);
nor U8480 (N_8480,N_7495,N_7502);
nand U8481 (N_8481,N_7973,N_7216);
or U8482 (N_8482,N_7907,N_7619);
nor U8483 (N_8483,N_7828,N_7104);
nand U8484 (N_8484,N_7601,N_7375);
nor U8485 (N_8485,N_7226,N_7886);
xor U8486 (N_8486,N_7033,N_7225);
and U8487 (N_8487,N_7548,N_7952);
xnor U8488 (N_8488,N_7737,N_7883);
and U8489 (N_8489,N_7898,N_7063);
xor U8490 (N_8490,N_7436,N_7900);
nand U8491 (N_8491,N_7432,N_7174);
xnor U8492 (N_8492,N_7419,N_7387);
nor U8493 (N_8493,N_7435,N_7208);
nand U8494 (N_8494,N_7516,N_7997);
nor U8495 (N_8495,N_7614,N_7764);
nor U8496 (N_8496,N_7690,N_7405);
nand U8497 (N_8497,N_7349,N_7180);
xnor U8498 (N_8498,N_7138,N_7124);
nor U8499 (N_8499,N_7147,N_7985);
and U8500 (N_8500,N_7670,N_7498);
nand U8501 (N_8501,N_7548,N_7988);
nand U8502 (N_8502,N_7454,N_7469);
xnor U8503 (N_8503,N_7084,N_7347);
or U8504 (N_8504,N_7742,N_7062);
and U8505 (N_8505,N_7060,N_7075);
nor U8506 (N_8506,N_7501,N_7382);
nand U8507 (N_8507,N_7478,N_7981);
and U8508 (N_8508,N_7496,N_7618);
nor U8509 (N_8509,N_7829,N_7335);
and U8510 (N_8510,N_7126,N_7359);
nor U8511 (N_8511,N_7959,N_7156);
nor U8512 (N_8512,N_7670,N_7152);
or U8513 (N_8513,N_7095,N_7011);
or U8514 (N_8514,N_7773,N_7135);
or U8515 (N_8515,N_7398,N_7642);
nor U8516 (N_8516,N_7634,N_7519);
nor U8517 (N_8517,N_7716,N_7441);
xnor U8518 (N_8518,N_7414,N_7914);
nor U8519 (N_8519,N_7325,N_7080);
and U8520 (N_8520,N_7460,N_7280);
nor U8521 (N_8521,N_7659,N_7184);
and U8522 (N_8522,N_7649,N_7454);
and U8523 (N_8523,N_7673,N_7400);
xnor U8524 (N_8524,N_7857,N_7807);
nor U8525 (N_8525,N_7757,N_7290);
or U8526 (N_8526,N_7042,N_7772);
nand U8527 (N_8527,N_7890,N_7351);
or U8528 (N_8528,N_7657,N_7388);
and U8529 (N_8529,N_7725,N_7648);
xnor U8530 (N_8530,N_7555,N_7661);
nor U8531 (N_8531,N_7299,N_7775);
or U8532 (N_8532,N_7923,N_7820);
nor U8533 (N_8533,N_7742,N_7840);
or U8534 (N_8534,N_7181,N_7553);
xnor U8535 (N_8535,N_7429,N_7908);
and U8536 (N_8536,N_7396,N_7854);
and U8537 (N_8537,N_7383,N_7094);
nor U8538 (N_8538,N_7322,N_7805);
xor U8539 (N_8539,N_7965,N_7491);
nor U8540 (N_8540,N_7424,N_7572);
and U8541 (N_8541,N_7576,N_7195);
nand U8542 (N_8542,N_7522,N_7450);
nand U8543 (N_8543,N_7036,N_7985);
nor U8544 (N_8544,N_7977,N_7794);
xor U8545 (N_8545,N_7492,N_7640);
nand U8546 (N_8546,N_7606,N_7136);
and U8547 (N_8547,N_7180,N_7950);
or U8548 (N_8548,N_7195,N_7053);
nand U8549 (N_8549,N_7586,N_7449);
or U8550 (N_8550,N_7278,N_7211);
and U8551 (N_8551,N_7367,N_7789);
or U8552 (N_8552,N_7611,N_7850);
and U8553 (N_8553,N_7829,N_7862);
or U8554 (N_8554,N_7287,N_7135);
xnor U8555 (N_8555,N_7138,N_7797);
nor U8556 (N_8556,N_7570,N_7404);
xor U8557 (N_8557,N_7346,N_7347);
nand U8558 (N_8558,N_7102,N_7463);
or U8559 (N_8559,N_7063,N_7519);
xnor U8560 (N_8560,N_7710,N_7901);
nand U8561 (N_8561,N_7649,N_7310);
nor U8562 (N_8562,N_7735,N_7791);
and U8563 (N_8563,N_7928,N_7560);
and U8564 (N_8564,N_7344,N_7505);
and U8565 (N_8565,N_7853,N_7702);
or U8566 (N_8566,N_7163,N_7394);
nor U8567 (N_8567,N_7101,N_7140);
or U8568 (N_8568,N_7135,N_7011);
and U8569 (N_8569,N_7068,N_7567);
or U8570 (N_8570,N_7729,N_7597);
nand U8571 (N_8571,N_7548,N_7749);
nand U8572 (N_8572,N_7846,N_7632);
xor U8573 (N_8573,N_7544,N_7998);
nor U8574 (N_8574,N_7610,N_7164);
or U8575 (N_8575,N_7124,N_7219);
nor U8576 (N_8576,N_7073,N_7839);
xnor U8577 (N_8577,N_7230,N_7133);
nand U8578 (N_8578,N_7422,N_7324);
and U8579 (N_8579,N_7058,N_7033);
or U8580 (N_8580,N_7883,N_7110);
nand U8581 (N_8581,N_7193,N_7622);
nand U8582 (N_8582,N_7004,N_7611);
or U8583 (N_8583,N_7489,N_7707);
nor U8584 (N_8584,N_7339,N_7883);
xor U8585 (N_8585,N_7078,N_7073);
or U8586 (N_8586,N_7237,N_7504);
nand U8587 (N_8587,N_7626,N_7234);
or U8588 (N_8588,N_7554,N_7157);
or U8589 (N_8589,N_7633,N_7233);
and U8590 (N_8590,N_7382,N_7534);
or U8591 (N_8591,N_7545,N_7691);
xnor U8592 (N_8592,N_7246,N_7937);
and U8593 (N_8593,N_7652,N_7765);
xor U8594 (N_8594,N_7578,N_7310);
nand U8595 (N_8595,N_7352,N_7844);
xnor U8596 (N_8596,N_7806,N_7560);
nor U8597 (N_8597,N_7025,N_7273);
nor U8598 (N_8598,N_7243,N_7625);
nor U8599 (N_8599,N_7877,N_7625);
or U8600 (N_8600,N_7300,N_7164);
nand U8601 (N_8601,N_7691,N_7879);
and U8602 (N_8602,N_7571,N_7684);
nand U8603 (N_8603,N_7942,N_7491);
nor U8604 (N_8604,N_7162,N_7074);
nand U8605 (N_8605,N_7905,N_7541);
and U8606 (N_8606,N_7622,N_7874);
or U8607 (N_8607,N_7857,N_7997);
nor U8608 (N_8608,N_7248,N_7297);
or U8609 (N_8609,N_7403,N_7203);
and U8610 (N_8610,N_7423,N_7885);
nor U8611 (N_8611,N_7043,N_7120);
and U8612 (N_8612,N_7157,N_7630);
xor U8613 (N_8613,N_7961,N_7021);
xnor U8614 (N_8614,N_7902,N_7357);
nand U8615 (N_8615,N_7926,N_7100);
nand U8616 (N_8616,N_7060,N_7170);
or U8617 (N_8617,N_7657,N_7556);
xor U8618 (N_8618,N_7555,N_7522);
and U8619 (N_8619,N_7666,N_7014);
nor U8620 (N_8620,N_7015,N_7920);
nor U8621 (N_8621,N_7712,N_7715);
and U8622 (N_8622,N_7040,N_7084);
xor U8623 (N_8623,N_7497,N_7420);
or U8624 (N_8624,N_7074,N_7018);
or U8625 (N_8625,N_7117,N_7805);
nand U8626 (N_8626,N_7113,N_7232);
xor U8627 (N_8627,N_7320,N_7314);
xor U8628 (N_8628,N_7083,N_7932);
nand U8629 (N_8629,N_7050,N_7909);
xnor U8630 (N_8630,N_7347,N_7698);
and U8631 (N_8631,N_7893,N_7388);
nand U8632 (N_8632,N_7701,N_7259);
nand U8633 (N_8633,N_7763,N_7336);
nor U8634 (N_8634,N_7260,N_7798);
and U8635 (N_8635,N_7341,N_7322);
nand U8636 (N_8636,N_7931,N_7681);
nand U8637 (N_8637,N_7402,N_7479);
nand U8638 (N_8638,N_7988,N_7104);
nand U8639 (N_8639,N_7280,N_7476);
and U8640 (N_8640,N_7761,N_7916);
nand U8641 (N_8641,N_7305,N_7104);
xor U8642 (N_8642,N_7492,N_7116);
nor U8643 (N_8643,N_7139,N_7649);
nor U8644 (N_8644,N_7341,N_7168);
and U8645 (N_8645,N_7603,N_7040);
nand U8646 (N_8646,N_7156,N_7780);
and U8647 (N_8647,N_7162,N_7962);
nor U8648 (N_8648,N_7843,N_7013);
and U8649 (N_8649,N_7787,N_7553);
and U8650 (N_8650,N_7926,N_7975);
nand U8651 (N_8651,N_7749,N_7135);
nand U8652 (N_8652,N_7329,N_7340);
nand U8653 (N_8653,N_7598,N_7373);
nand U8654 (N_8654,N_7531,N_7372);
and U8655 (N_8655,N_7368,N_7814);
and U8656 (N_8656,N_7143,N_7700);
nor U8657 (N_8657,N_7718,N_7227);
xnor U8658 (N_8658,N_7754,N_7870);
nand U8659 (N_8659,N_7869,N_7832);
xor U8660 (N_8660,N_7514,N_7388);
nor U8661 (N_8661,N_7266,N_7784);
and U8662 (N_8662,N_7770,N_7172);
and U8663 (N_8663,N_7196,N_7591);
nor U8664 (N_8664,N_7505,N_7374);
or U8665 (N_8665,N_7595,N_7026);
nand U8666 (N_8666,N_7443,N_7633);
xor U8667 (N_8667,N_7319,N_7988);
and U8668 (N_8668,N_7797,N_7464);
and U8669 (N_8669,N_7588,N_7650);
xor U8670 (N_8670,N_7465,N_7351);
nand U8671 (N_8671,N_7655,N_7340);
and U8672 (N_8672,N_7470,N_7518);
or U8673 (N_8673,N_7538,N_7720);
nor U8674 (N_8674,N_7580,N_7170);
and U8675 (N_8675,N_7634,N_7915);
xor U8676 (N_8676,N_7869,N_7874);
or U8677 (N_8677,N_7503,N_7358);
nand U8678 (N_8678,N_7872,N_7909);
or U8679 (N_8679,N_7108,N_7122);
and U8680 (N_8680,N_7885,N_7564);
nor U8681 (N_8681,N_7610,N_7780);
nor U8682 (N_8682,N_7641,N_7954);
nor U8683 (N_8683,N_7321,N_7562);
nand U8684 (N_8684,N_7866,N_7338);
xor U8685 (N_8685,N_7972,N_7034);
xnor U8686 (N_8686,N_7392,N_7188);
nor U8687 (N_8687,N_7411,N_7514);
nand U8688 (N_8688,N_7451,N_7535);
xor U8689 (N_8689,N_7884,N_7832);
nor U8690 (N_8690,N_7065,N_7159);
nand U8691 (N_8691,N_7319,N_7065);
and U8692 (N_8692,N_7019,N_7384);
nand U8693 (N_8693,N_7180,N_7790);
or U8694 (N_8694,N_7395,N_7452);
nor U8695 (N_8695,N_7271,N_7776);
xor U8696 (N_8696,N_7669,N_7988);
nor U8697 (N_8697,N_7686,N_7622);
nand U8698 (N_8698,N_7133,N_7426);
and U8699 (N_8699,N_7756,N_7282);
xnor U8700 (N_8700,N_7453,N_7194);
nor U8701 (N_8701,N_7825,N_7026);
xor U8702 (N_8702,N_7090,N_7844);
xor U8703 (N_8703,N_7170,N_7940);
nand U8704 (N_8704,N_7071,N_7877);
and U8705 (N_8705,N_7412,N_7047);
nor U8706 (N_8706,N_7556,N_7116);
or U8707 (N_8707,N_7089,N_7436);
or U8708 (N_8708,N_7700,N_7870);
or U8709 (N_8709,N_7164,N_7798);
nand U8710 (N_8710,N_7667,N_7391);
nor U8711 (N_8711,N_7163,N_7649);
xnor U8712 (N_8712,N_7746,N_7819);
nor U8713 (N_8713,N_7431,N_7708);
nand U8714 (N_8714,N_7025,N_7453);
nand U8715 (N_8715,N_7248,N_7978);
or U8716 (N_8716,N_7363,N_7374);
and U8717 (N_8717,N_7573,N_7397);
nor U8718 (N_8718,N_7184,N_7887);
or U8719 (N_8719,N_7114,N_7922);
or U8720 (N_8720,N_7425,N_7505);
nor U8721 (N_8721,N_7231,N_7284);
nor U8722 (N_8722,N_7569,N_7591);
nand U8723 (N_8723,N_7729,N_7752);
and U8724 (N_8724,N_7092,N_7070);
or U8725 (N_8725,N_7681,N_7975);
or U8726 (N_8726,N_7541,N_7783);
and U8727 (N_8727,N_7734,N_7044);
and U8728 (N_8728,N_7057,N_7578);
and U8729 (N_8729,N_7916,N_7290);
nor U8730 (N_8730,N_7773,N_7265);
nor U8731 (N_8731,N_7040,N_7763);
nor U8732 (N_8732,N_7883,N_7542);
nor U8733 (N_8733,N_7970,N_7999);
nand U8734 (N_8734,N_7937,N_7356);
nand U8735 (N_8735,N_7638,N_7484);
and U8736 (N_8736,N_7076,N_7365);
xor U8737 (N_8737,N_7792,N_7933);
or U8738 (N_8738,N_7412,N_7694);
nand U8739 (N_8739,N_7080,N_7417);
or U8740 (N_8740,N_7386,N_7288);
and U8741 (N_8741,N_7462,N_7313);
or U8742 (N_8742,N_7813,N_7740);
nand U8743 (N_8743,N_7947,N_7423);
nor U8744 (N_8744,N_7116,N_7102);
and U8745 (N_8745,N_7284,N_7714);
nand U8746 (N_8746,N_7553,N_7714);
or U8747 (N_8747,N_7455,N_7701);
nor U8748 (N_8748,N_7530,N_7550);
xnor U8749 (N_8749,N_7792,N_7306);
nand U8750 (N_8750,N_7618,N_7560);
and U8751 (N_8751,N_7363,N_7442);
or U8752 (N_8752,N_7895,N_7534);
nand U8753 (N_8753,N_7697,N_7016);
nor U8754 (N_8754,N_7528,N_7068);
nor U8755 (N_8755,N_7778,N_7102);
nor U8756 (N_8756,N_7692,N_7645);
or U8757 (N_8757,N_7401,N_7023);
nor U8758 (N_8758,N_7081,N_7731);
and U8759 (N_8759,N_7246,N_7104);
or U8760 (N_8760,N_7142,N_7456);
nor U8761 (N_8761,N_7293,N_7728);
and U8762 (N_8762,N_7274,N_7614);
nand U8763 (N_8763,N_7974,N_7152);
xnor U8764 (N_8764,N_7820,N_7480);
or U8765 (N_8765,N_7062,N_7052);
xnor U8766 (N_8766,N_7836,N_7999);
xor U8767 (N_8767,N_7665,N_7181);
nand U8768 (N_8768,N_7413,N_7720);
nor U8769 (N_8769,N_7492,N_7539);
nor U8770 (N_8770,N_7689,N_7262);
nand U8771 (N_8771,N_7318,N_7129);
or U8772 (N_8772,N_7449,N_7438);
and U8773 (N_8773,N_7875,N_7352);
nand U8774 (N_8774,N_7506,N_7299);
and U8775 (N_8775,N_7145,N_7723);
xnor U8776 (N_8776,N_7420,N_7910);
nand U8777 (N_8777,N_7076,N_7918);
nand U8778 (N_8778,N_7079,N_7059);
nand U8779 (N_8779,N_7360,N_7011);
xor U8780 (N_8780,N_7735,N_7833);
and U8781 (N_8781,N_7910,N_7677);
xnor U8782 (N_8782,N_7935,N_7272);
nor U8783 (N_8783,N_7944,N_7370);
xor U8784 (N_8784,N_7901,N_7936);
nand U8785 (N_8785,N_7435,N_7930);
and U8786 (N_8786,N_7554,N_7566);
xnor U8787 (N_8787,N_7488,N_7067);
xnor U8788 (N_8788,N_7664,N_7306);
xor U8789 (N_8789,N_7638,N_7759);
and U8790 (N_8790,N_7142,N_7827);
or U8791 (N_8791,N_7087,N_7973);
and U8792 (N_8792,N_7570,N_7308);
xnor U8793 (N_8793,N_7384,N_7614);
and U8794 (N_8794,N_7698,N_7683);
and U8795 (N_8795,N_7110,N_7337);
nand U8796 (N_8796,N_7549,N_7667);
nand U8797 (N_8797,N_7767,N_7955);
and U8798 (N_8798,N_7451,N_7297);
nor U8799 (N_8799,N_7998,N_7637);
nor U8800 (N_8800,N_7114,N_7334);
nand U8801 (N_8801,N_7076,N_7934);
or U8802 (N_8802,N_7330,N_7913);
and U8803 (N_8803,N_7098,N_7519);
and U8804 (N_8804,N_7339,N_7849);
and U8805 (N_8805,N_7038,N_7774);
nor U8806 (N_8806,N_7617,N_7151);
or U8807 (N_8807,N_7216,N_7279);
nand U8808 (N_8808,N_7980,N_7859);
nand U8809 (N_8809,N_7531,N_7449);
nand U8810 (N_8810,N_7285,N_7634);
and U8811 (N_8811,N_7739,N_7198);
and U8812 (N_8812,N_7283,N_7819);
and U8813 (N_8813,N_7531,N_7885);
xnor U8814 (N_8814,N_7987,N_7703);
nor U8815 (N_8815,N_7025,N_7257);
nor U8816 (N_8816,N_7493,N_7699);
nor U8817 (N_8817,N_7258,N_7172);
xor U8818 (N_8818,N_7631,N_7294);
or U8819 (N_8819,N_7248,N_7576);
nor U8820 (N_8820,N_7949,N_7256);
nor U8821 (N_8821,N_7867,N_7240);
nand U8822 (N_8822,N_7632,N_7507);
and U8823 (N_8823,N_7088,N_7186);
and U8824 (N_8824,N_7959,N_7556);
xnor U8825 (N_8825,N_7742,N_7448);
or U8826 (N_8826,N_7195,N_7499);
nor U8827 (N_8827,N_7067,N_7223);
and U8828 (N_8828,N_7854,N_7828);
and U8829 (N_8829,N_7159,N_7291);
and U8830 (N_8830,N_7660,N_7579);
and U8831 (N_8831,N_7936,N_7071);
xor U8832 (N_8832,N_7210,N_7092);
xnor U8833 (N_8833,N_7134,N_7629);
nand U8834 (N_8834,N_7394,N_7526);
xnor U8835 (N_8835,N_7571,N_7681);
nor U8836 (N_8836,N_7768,N_7219);
xor U8837 (N_8837,N_7166,N_7740);
nand U8838 (N_8838,N_7482,N_7987);
and U8839 (N_8839,N_7406,N_7644);
and U8840 (N_8840,N_7932,N_7277);
xnor U8841 (N_8841,N_7936,N_7762);
nor U8842 (N_8842,N_7335,N_7716);
xor U8843 (N_8843,N_7058,N_7711);
or U8844 (N_8844,N_7888,N_7032);
xor U8845 (N_8845,N_7197,N_7711);
nor U8846 (N_8846,N_7800,N_7400);
and U8847 (N_8847,N_7306,N_7531);
and U8848 (N_8848,N_7469,N_7781);
or U8849 (N_8849,N_7661,N_7168);
nor U8850 (N_8850,N_7254,N_7047);
nand U8851 (N_8851,N_7937,N_7531);
and U8852 (N_8852,N_7137,N_7142);
nor U8853 (N_8853,N_7534,N_7054);
and U8854 (N_8854,N_7583,N_7378);
nand U8855 (N_8855,N_7052,N_7947);
xor U8856 (N_8856,N_7499,N_7627);
and U8857 (N_8857,N_7580,N_7623);
or U8858 (N_8858,N_7033,N_7020);
nor U8859 (N_8859,N_7803,N_7558);
nand U8860 (N_8860,N_7761,N_7495);
or U8861 (N_8861,N_7478,N_7336);
xnor U8862 (N_8862,N_7461,N_7955);
nor U8863 (N_8863,N_7134,N_7099);
nand U8864 (N_8864,N_7079,N_7664);
or U8865 (N_8865,N_7532,N_7521);
nor U8866 (N_8866,N_7815,N_7294);
and U8867 (N_8867,N_7728,N_7454);
nor U8868 (N_8868,N_7601,N_7885);
or U8869 (N_8869,N_7916,N_7753);
nor U8870 (N_8870,N_7839,N_7626);
nand U8871 (N_8871,N_7053,N_7188);
xor U8872 (N_8872,N_7696,N_7097);
or U8873 (N_8873,N_7741,N_7239);
xnor U8874 (N_8874,N_7111,N_7998);
nand U8875 (N_8875,N_7892,N_7403);
xnor U8876 (N_8876,N_7923,N_7643);
xor U8877 (N_8877,N_7772,N_7547);
and U8878 (N_8878,N_7798,N_7696);
xnor U8879 (N_8879,N_7246,N_7968);
or U8880 (N_8880,N_7965,N_7341);
or U8881 (N_8881,N_7857,N_7537);
nor U8882 (N_8882,N_7565,N_7249);
nor U8883 (N_8883,N_7723,N_7134);
nand U8884 (N_8884,N_7006,N_7660);
xor U8885 (N_8885,N_7388,N_7984);
nand U8886 (N_8886,N_7434,N_7217);
or U8887 (N_8887,N_7234,N_7588);
nor U8888 (N_8888,N_7407,N_7072);
nor U8889 (N_8889,N_7182,N_7696);
xnor U8890 (N_8890,N_7707,N_7226);
nand U8891 (N_8891,N_7738,N_7303);
nand U8892 (N_8892,N_7850,N_7161);
nor U8893 (N_8893,N_7086,N_7893);
or U8894 (N_8894,N_7404,N_7618);
nand U8895 (N_8895,N_7376,N_7831);
nand U8896 (N_8896,N_7007,N_7093);
nand U8897 (N_8897,N_7214,N_7546);
or U8898 (N_8898,N_7771,N_7501);
and U8899 (N_8899,N_7790,N_7871);
nor U8900 (N_8900,N_7448,N_7479);
xor U8901 (N_8901,N_7833,N_7114);
nand U8902 (N_8902,N_7808,N_7696);
and U8903 (N_8903,N_7688,N_7801);
xnor U8904 (N_8904,N_7919,N_7046);
or U8905 (N_8905,N_7853,N_7457);
or U8906 (N_8906,N_7640,N_7609);
nor U8907 (N_8907,N_7333,N_7160);
and U8908 (N_8908,N_7790,N_7587);
or U8909 (N_8909,N_7948,N_7821);
or U8910 (N_8910,N_7113,N_7560);
xnor U8911 (N_8911,N_7472,N_7734);
nand U8912 (N_8912,N_7150,N_7743);
and U8913 (N_8913,N_7244,N_7845);
xor U8914 (N_8914,N_7395,N_7728);
and U8915 (N_8915,N_7751,N_7907);
and U8916 (N_8916,N_7402,N_7076);
and U8917 (N_8917,N_7029,N_7906);
xnor U8918 (N_8918,N_7852,N_7738);
and U8919 (N_8919,N_7138,N_7869);
and U8920 (N_8920,N_7496,N_7958);
and U8921 (N_8921,N_7811,N_7339);
or U8922 (N_8922,N_7561,N_7213);
nand U8923 (N_8923,N_7936,N_7106);
or U8924 (N_8924,N_7654,N_7201);
nand U8925 (N_8925,N_7983,N_7577);
xor U8926 (N_8926,N_7154,N_7212);
nand U8927 (N_8927,N_7998,N_7877);
and U8928 (N_8928,N_7091,N_7902);
nand U8929 (N_8929,N_7896,N_7244);
xor U8930 (N_8930,N_7473,N_7505);
or U8931 (N_8931,N_7283,N_7116);
or U8932 (N_8932,N_7862,N_7807);
nor U8933 (N_8933,N_7014,N_7678);
and U8934 (N_8934,N_7899,N_7018);
and U8935 (N_8935,N_7947,N_7746);
or U8936 (N_8936,N_7531,N_7629);
or U8937 (N_8937,N_7228,N_7215);
nor U8938 (N_8938,N_7160,N_7053);
nor U8939 (N_8939,N_7903,N_7496);
and U8940 (N_8940,N_7786,N_7806);
xor U8941 (N_8941,N_7501,N_7169);
nand U8942 (N_8942,N_7142,N_7166);
xor U8943 (N_8943,N_7998,N_7322);
nor U8944 (N_8944,N_7208,N_7698);
nor U8945 (N_8945,N_7081,N_7383);
nor U8946 (N_8946,N_7288,N_7693);
and U8947 (N_8947,N_7132,N_7174);
nor U8948 (N_8948,N_7189,N_7232);
xor U8949 (N_8949,N_7851,N_7538);
or U8950 (N_8950,N_7729,N_7654);
and U8951 (N_8951,N_7948,N_7095);
or U8952 (N_8952,N_7603,N_7568);
and U8953 (N_8953,N_7781,N_7784);
nor U8954 (N_8954,N_7631,N_7285);
and U8955 (N_8955,N_7214,N_7900);
nand U8956 (N_8956,N_7634,N_7730);
nand U8957 (N_8957,N_7883,N_7260);
nor U8958 (N_8958,N_7211,N_7338);
xnor U8959 (N_8959,N_7293,N_7989);
nand U8960 (N_8960,N_7668,N_7702);
xor U8961 (N_8961,N_7562,N_7714);
and U8962 (N_8962,N_7291,N_7878);
nand U8963 (N_8963,N_7961,N_7197);
and U8964 (N_8964,N_7368,N_7303);
nor U8965 (N_8965,N_7717,N_7796);
nor U8966 (N_8966,N_7035,N_7455);
and U8967 (N_8967,N_7680,N_7392);
and U8968 (N_8968,N_7014,N_7714);
nor U8969 (N_8969,N_7282,N_7349);
nand U8970 (N_8970,N_7954,N_7488);
or U8971 (N_8971,N_7932,N_7288);
and U8972 (N_8972,N_7266,N_7540);
or U8973 (N_8973,N_7519,N_7761);
xnor U8974 (N_8974,N_7555,N_7888);
or U8975 (N_8975,N_7660,N_7052);
and U8976 (N_8976,N_7164,N_7804);
nand U8977 (N_8977,N_7094,N_7373);
nor U8978 (N_8978,N_7655,N_7740);
and U8979 (N_8979,N_7465,N_7972);
nor U8980 (N_8980,N_7697,N_7480);
or U8981 (N_8981,N_7018,N_7628);
xor U8982 (N_8982,N_7498,N_7987);
xor U8983 (N_8983,N_7809,N_7462);
xor U8984 (N_8984,N_7095,N_7167);
or U8985 (N_8985,N_7457,N_7081);
nor U8986 (N_8986,N_7477,N_7994);
nand U8987 (N_8987,N_7134,N_7775);
nand U8988 (N_8988,N_7025,N_7416);
and U8989 (N_8989,N_7252,N_7576);
and U8990 (N_8990,N_7392,N_7254);
xnor U8991 (N_8991,N_7132,N_7640);
nor U8992 (N_8992,N_7845,N_7377);
or U8993 (N_8993,N_7456,N_7510);
or U8994 (N_8994,N_7302,N_7320);
xor U8995 (N_8995,N_7585,N_7618);
xor U8996 (N_8996,N_7524,N_7811);
and U8997 (N_8997,N_7788,N_7733);
and U8998 (N_8998,N_7378,N_7775);
xnor U8999 (N_8999,N_7803,N_7965);
xnor U9000 (N_9000,N_8679,N_8430);
nor U9001 (N_9001,N_8800,N_8878);
nor U9002 (N_9002,N_8027,N_8236);
xor U9003 (N_9003,N_8008,N_8605);
and U9004 (N_9004,N_8045,N_8775);
nand U9005 (N_9005,N_8967,N_8603);
and U9006 (N_9006,N_8713,N_8900);
and U9007 (N_9007,N_8639,N_8655);
nor U9008 (N_9008,N_8864,N_8038);
nor U9009 (N_9009,N_8353,N_8745);
nor U9010 (N_9010,N_8442,N_8369);
nand U9011 (N_9011,N_8565,N_8357);
and U9012 (N_9012,N_8462,N_8367);
xnor U9013 (N_9013,N_8464,N_8562);
nand U9014 (N_9014,N_8798,N_8948);
and U9015 (N_9015,N_8450,N_8458);
xnor U9016 (N_9016,N_8057,N_8966);
xor U9017 (N_9017,N_8403,N_8472);
xnor U9018 (N_9018,N_8059,N_8697);
nor U9019 (N_9019,N_8232,N_8742);
nand U9020 (N_9020,N_8041,N_8460);
and U9021 (N_9021,N_8613,N_8972);
and U9022 (N_9022,N_8939,N_8677);
nor U9023 (N_9023,N_8485,N_8456);
nor U9024 (N_9024,N_8769,N_8201);
or U9025 (N_9025,N_8830,N_8061);
nand U9026 (N_9026,N_8991,N_8482);
or U9027 (N_9027,N_8951,N_8902);
nor U9028 (N_9028,N_8424,N_8189);
nand U9029 (N_9029,N_8338,N_8540);
nor U9030 (N_9030,N_8068,N_8223);
and U9031 (N_9031,N_8764,N_8199);
or U9032 (N_9032,N_8203,N_8139);
nand U9033 (N_9033,N_8977,N_8283);
nor U9034 (N_9034,N_8310,N_8543);
or U9035 (N_9035,N_8163,N_8617);
and U9036 (N_9036,N_8166,N_8036);
and U9037 (N_9037,N_8693,N_8842);
or U9038 (N_9038,N_8641,N_8593);
nor U9039 (N_9039,N_8984,N_8720);
nand U9040 (N_9040,N_8893,N_8071);
nand U9041 (N_9041,N_8569,N_8635);
or U9042 (N_9042,N_8894,N_8663);
and U9043 (N_9043,N_8327,N_8858);
nand U9044 (N_9044,N_8585,N_8938);
xnor U9045 (N_9045,N_8123,N_8293);
and U9046 (N_9046,N_8409,N_8446);
and U9047 (N_9047,N_8321,N_8486);
xor U9048 (N_9048,N_8350,N_8457);
xnor U9049 (N_9049,N_8261,N_8561);
nand U9050 (N_9050,N_8471,N_8859);
nand U9051 (N_9051,N_8454,N_8592);
nand U9052 (N_9052,N_8924,N_8640);
or U9053 (N_9053,N_8533,N_8459);
nand U9054 (N_9054,N_8700,N_8684);
and U9055 (N_9055,N_8136,N_8314);
and U9056 (N_9056,N_8699,N_8777);
or U9057 (N_9057,N_8422,N_8807);
or U9058 (N_9058,N_8214,N_8823);
nand U9059 (N_9059,N_8872,N_8668);
or U9060 (N_9060,N_8179,N_8671);
xor U9061 (N_9061,N_8082,N_8771);
and U9062 (N_9062,N_8116,N_8575);
nand U9063 (N_9063,N_8757,N_8297);
or U9064 (N_9064,N_8149,N_8161);
and U9065 (N_9065,N_8867,N_8110);
nand U9066 (N_9066,N_8710,N_8860);
and U9067 (N_9067,N_8755,N_8686);
xnor U9068 (N_9068,N_8352,N_8481);
and U9069 (N_9069,N_8682,N_8219);
xnor U9070 (N_9070,N_8397,N_8672);
or U9071 (N_9071,N_8373,N_8866);
nor U9072 (N_9072,N_8784,N_8174);
nor U9073 (N_9073,N_8616,N_8437);
nand U9074 (N_9074,N_8208,N_8590);
xnor U9075 (N_9075,N_8959,N_8138);
nor U9076 (N_9076,N_8414,N_8928);
or U9077 (N_9077,N_8088,N_8703);
nand U9078 (N_9078,N_8254,N_8105);
and U9079 (N_9079,N_8147,N_8490);
xor U9080 (N_9080,N_8268,N_8505);
nand U9081 (N_9081,N_8191,N_8003);
xor U9082 (N_9082,N_8349,N_8124);
nor U9083 (N_9083,N_8478,N_8384);
nand U9084 (N_9084,N_8553,N_8962);
xnor U9085 (N_9085,N_8760,N_8722);
nor U9086 (N_9086,N_8580,N_8032);
nand U9087 (N_9087,N_8588,N_8887);
nor U9088 (N_9088,N_8625,N_8183);
and U9089 (N_9089,N_8584,N_8224);
nand U9090 (N_9090,N_8670,N_8730);
or U9091 (N_9091,N_8212,N_8066);
and U9092 (N_9092,N_8850,N_8547);
and U9093 (N_9093,N_8521,N_8520);
or U9094 (N_9094,N_8065,N_8111);
or U9095 (N_9095,N_8564,N_8824);
xnor U9096 (N_9096,N_8282,N_8342);
or U9097 (N_9097,N_8549,N_8738);
xor U9098 (N_9098,N_8762,N_8811);
nand U9099 (N_9099,N_8766,N_8341);
nor U9100 (N_9100,N_8740,N_8573);
nand U9101 (N_9101,N_8746,N_8542);
nor U9102 (N_9102,N_8463,N_8048);
nand U9103 (N_9103,N_8455,N_8210);
xnor U9104 (N_9104,N_8748,N_8998);
or U9105 (N_9105,N_8644,N_8904);
nor U9106 (N_9106,N_8218,N_8465);
or U9107 (N_9107,N_8200,N_8133);
nor U9108 (N_9108,N_8243,N_8091);
nor U9109 (N_9109,N_8107,N_8122);
and U9110 (N_9110,N_8954,N_8906);
nand U9111 (N_9111,N_8865,N_8546);
nor U9112 (N_9112,N_8378,N_8031);
and U9113 (N_9113,N_8736,N_8598);
nor U9114 (N_9114,N_8137,N_8674);
and U9115 (N_9115,N_8491,N_8368);
nand U9116 (N_9116,N_8690,N_8918);
nand U9117 (N_9117,N_8932,N_8646);
and U9118 (N_9118,N_8750,N_8789);
xor U9119 (N_9119,N_8175,N_8556);
nand U9120 (N_9120,N_8417,N_8721);
nor U9121 (N_9121,N_8407,N_8198);
xor U9122 (N_9122,N_8099,N_8994);
nor U9123 (N_9123,N_8390,N_8415);
or U9124 (N_9124,N_8381,N_8987);
and U9125 (N_9125,N_8541,N_8899);
and U9126 (N_9126,N_8156,N_8093);
nand U9127 (N_9127,N_8531,N_8770);
nor U9128 (N_9128,N_8386,N_8062);
or U9129 (N_9129,N_8577,N_8474);
nand U9130 (N_9130,N_8204,N_8952);
and U9131 (N_9131,N_8552,N_8120);
nor U9132 (N_9132,N_8050,N_8652);
or U9133 (N_9133,N_8763,N_8279);
and U9134 (N_9134,N_8339,N_8011);
and U9135 (N_9135,N_8944,N_8258);
nand U9136 (N_9136,N_8266,N_8026);
xnor U9137 (N_9137,N_8252,N_8876);
nor U9138 (N_9138,N_8586,N_8963);
xnor U9139 (N_9139,N_8375,N_8265);
and U9140 (N_9140,N_8799,N_8946);
xor U9141 (N_9141,N_8796,N_8854);
or U9142 (N_9142,N_8599,N_8404);
nand U9143 (N_9143,N_8498,N_8097);
and U9144 (N_9144,N_8012,N_8947);
or U9145 (N_9145,N_8309,N_8567);
nor U9146 (N_9146,N_8919,N_8631);
nor U9147 (N_9147,N_8802,N_8018);
nand U9148 (N_9148,N_8995,N_8473);
xnor U9149 (N_9149,N_8233,N_8935);
nand U9150 (N_9150,N_8571,N_8269);
or U9151 (N_9151,N_8634,N_8255);
nand U9152 (N_9152,N_8131,N_8129);
and U9153 (N_9153,N_8080,N_8981);
xor U9154 (N_9154,N_8165,N_8500);
nand U9155 (N_9155,N_8786,N_8595);
or U9156 (N_9156,N_8162,N_8047);
and U9157 (N_9157,N_8790,N_8953);
xor U9158 (N_9158,N_8756,N_8753);
or U9159 (N_9159,N_8544,N_8570);
xnor U9160 (N_9160,N_8436,N_8278);
or U9161 (N_9161,N_8361,N_8379);
nor U9162 (N_9162,N_8461,N_8128);
or U9163 (N_9163,N_8318,N_8666);
xor U9164 (N_9164,N_8364,N_8413);
xor U9165 (N_9165,N_8626,N_8724);
nor U9166 (N_9166,N_8167,N_8661);
or U9167 (N_9167,N_8072,N_8040);
nor U9168 (N_9168,N_8271,N_8615);
and U9169 (N_9169,N_8836,N_8145);
nor U9170 (N_9170,N_8767,N_8073);
nor U9171 (N_9171,N_8717,N_8094);
or U9172 (N_9172,N_8920,N_8832);
nand U9173 (N_9173,N_8237,N_8999);
xnor U9174 (N_9174,N_8095,N_8328);
xor U9175 (N_9175,N_8492,N_8602);
xnor U9176 (N_9176,N_8211,N_8083);
or U9177 (N_9177,N_8007,N_8795);
nand U9178 (N_9178,N_8551,N_8619);
and U9179 (N_9179,N_8209,N_8936);
xor U9180 (N_9180,N_8934,N_8608);
nand U9181 (N_9181,N_8370,N_8805);
and U9182 (N_9182,N_8344,N_8714);
nand U9183 (N_9183,N_8319,N_8525);
nand U9184 (N_9184,N_8362,N_8180);
nand U9185 (N_9185,N_8499,N_8028);
xor U9186 (N_9186,N_8443,N_8827);
and U9187 (N_9187,N_8519,N_8776);
xnor U9188 (N_9188,N_8194,N_8423);
and U9189 (N_9189,N_8197,N_8815);
xor U9190 (N_9190,N_8664,N_8862);
xnor U9191 (N_9191,N_8019,N_8971);
nand U9192 (N_9192,N_8146,N_8432);
nand U9193 (N_9193,N_8705,N_8662);
and U9194 (N_9194,N_8335,N_8964);
or U9195 (N_9195,N_8930,N_8431);
and U9196 (N_9196,N_8067,N_8558);
nand U9197 (N_9197,N_8726,N_8734);
xor U9198 (N_9198,N_8758,N_8659);
nor U9199 (N_9199,N_8821,N_8933);
nor U9200 (N_9200,N_8820,N_8227);
or U9201 (N_9201,N_8250,N_8391);
xnor U9202 (N_9202,N_8522,N_8627);
and U9203 (N_9203,N_8246,N_8704);
xor U9204 (N_9204,N_8060,N_8042);
or U9205 (N_9205,N_8155,N_8121);
nor U9206 (N_9206,N_8629,N_8380);
and U9207 (N_9207,N_8345,N_8915);
nor U9208 (N_9208,N_8125,N_8648);
nand U9209 (N_9209,N_8070,N_8401);
or U9210 (N_9210,N_8809,N_8804);
and U9211 (N_9211,N_8957,N_8256);
nand U9212 (N_9212,N_8911,N_8594);
or U9213 (N_9213,N_8891,N_8468);
nor U9214 (N_9214,N_8618,N_8772);
or U9215 (N_9215,N_8049,N_8645);
nor U9216 (N_9216,N_8510,N_8143);
xor U9217 (N_9217,N_8970,N_8480);
nor U9218 (N_9218,N_8537,N_8851);
xor U9219 (N_9219,N_8728,N_8782);
nor U9220 (N_9220,N_8877,N_8829);
or U9221 (N_9221,N_8150,N_8638);
and U9222 (N_9222,N_8377,N_8992);
nand U9223 (N_9223,N_8419,N_8975);
nor U9224 (N_9224,N_8910,N_8169);
nand U9225 (N_9225,N_8030,N_8515);
and U9226 (N_9226,N_8142,N_8322);
xor U9227 (N_9227,N_8673,N_8117);
or U9228 (N_9228,N_8333,N_8908);
or U9229 (N_9229,N_8834,N_8239);
and U9230 (N_9230,N_8871,N_8284);
and U9231 (N_9231,N_8444,N_8006);
or U9232 (N_9232,N_8536,N_8507);
nor U9233 (N_9233,N_8532,N_8400);
xor U9234 (N_9234,N_8861,N_8325);
and U9235 (N_9235,N_8650,N_8287);
or U9236 (N_9236,N_8574,N_8152);
nand U9237 (N_9237,N_8922,N_8702);
or U9238 (N_9238,N_8441,N_8248);
nand U9239 (N_9239,N_8270,N_8421);
and U9240 (N_9240,N_8363,N_8818);
nand U9241 (N_9241,N_8729,N_8509);
and U9242 (N_9242,N_8304,N_8184);
and U9243 (N_9243,N_8780,N_8604);
and U9244 (N_9244,N_8968,N_8791);
nor U9245 (N_9245,N_8177,N_8759);
or U9246 (N_9246,N_8609,N_8600);
and U9247 (N_9247,N_8418,N_8448);
nor U9248 (N_9248,N_8942,N_8596);
nand U9249 (N_9249,N_8831,N_8043);
nor U9250 (N_9250,N_8225,N_8281);
or U9251 (N_9251,N_8986,N_8399);
and U9252 (N_9252,N_8495,N_8852);
nand U9253 (N_9253,N_8503,N_8579);
nor U9254 (N_9254,N_8601,N_8427);
and U9255 (N_9255,N_8037,N_8921);
nand U9256 (N_9256,N_8181,N_8883);
nand U9257 (N_9257,N_8497,N_8979);
nand U9258 (N_9258,N_8299,N_8909);
or U9259 (N_9259,N_8108,N_8305);
nor U9260 (N_9260,N_8438,N_8242);
and U9261 (N_9261,N_8913,N_8170);
and U9262 (N_9262,N_8451,N_8466);
xnor U9263 (N_9263,N_8220,N_8896);
nor U9264 (N_9264,N_8078,N_8085);
nor U9265 (N_9265,N_8649,N_8405);
nand U9266 (N_9266,N_8317,N_8846);
or U9267 (N_9267,N_8990,N_8694);
nand U9268 (N_9268,N_8044,N_8744);
or U9269 (N_9269,N_8535,N_8127);
and U9270 (N_9270,N_8743,N_8814);
and U9271 (N_9271,N_8336,N_8501);
or U9272 (N_9272,N_8905,N_8803);
nor U9273 (N_9273,N_8857,N_8941);
nor U9274 (N_9274,N_8240,N_8222);
nor U9275 (N_9275,N_8251,N_8692);
nand U9276 (N_9276,N_8015,N_8187);
or U9277 (N_9277,N_8514,N_8768);
or U9278 (N_9278,N_8783,N_8359);
xor U9279 (N_9279,N_8897,N_8229);
nor U9280 (N_9280,N_8000,N_8737);
and U9281 (N_9281,N_8069,N_8812);
nor U9282 (N_9282,N_8965,N_8005);
xor U9283 (N_9283,N_8195,N_8524);
nor U9284 (N_9284,N_8207,N_8192);
nor U9285 (N_9285,N_8315,N_8633);
nand U9286 (N_9286,N_8504,N_8848);
xnor U9287 (N_9287,N_8263,N_8630);
xnor U9288 (N_9288,N_8548,N_8323);
and U9289 (N_9289,N_8410,N_8171);
and U9290 (N_9290,N_8022,N_8013);
xnor U9291 (N_9291,N_8329,N_8695);
and U9292 (N_9292,N_8589,N_8356);
or U9293 (N_9293,N_8993,N_8733);
and U9294 (N_9294,N_8021,N_8628);
nand U9295 (N_9295,N_8973,N_8539);
nand U9296 (N_9296,N_8098,N_8493);
and U9297 (N_9297,N_8063,N_8560);
nor U9298 (N_9298,N_8385,N_8428);
nor U9299 (N_9299,N_8898,N_8833);
xnor U9300 (N_9300,N_8051,N_8676);
xnor U9301 (N_9301,N_8334,N_8518);
and U9302 (N_9302,N_8917,N_8835);
or U9303 (N_9303,N_8653,N_8058);
or U9304 (N_9304,N_8033,N_8190);
nor U9305 (N_9305,N_8716,N_8907);
nand U9306 (N_9306,N_8371,N_8054);
and U9307 (N_9307,N_8453,N_8838);
xnor U9308 (N_9308,N_8837,N_8940);
xor U9309 (N_9309,N_8416,N_8159);
xnor U9310 (N_9310,N_8527,N_8889);
and U9311 (N_9311,N_8508,N_8496);
nor U9312 (N_9312,N_8289,N_8182);
or U9313 (N_9313,N_8985,N_8885);
nor U9314 (N_9314,N_8274,N_8374);
or U9315 (N_9315,N_8193,N_8280);
xor U9316 (N_9316,N_8234,N_8779);
xor U9317 (N_9317,N_8840,N_8228);
nand U9318 (N_9318,N_8119,N_8186);
and U9319 (N_9319,N_8660,N_8004);
and U9320 (N_9320,N_8259,N_8132);
or U9321 (N_9321,N_8020,N_8879);
nand U9322 (N_9322,N_8685,N_8039);
or U9323 (N_9323,N_8286,N_8530);
nand U9324 (N_9324,N_8958,N_8778);
nor U9325 (N_9325,N_8669,N_8106);
nand U9326 (N_9326,N_8387,N_8077);
or U9327 (N_9327,N_8988,N_8412);
nand U9328 (N_9328,N_8882,N_8731);
or U9329 (N_9329,N_8273,N_8402);
or U9330 (N_9330,N_8185,N_8997);
and U9331 (N_9331,N_8024,N_8614);
and U9332 (N_9332,N_8439,N_8135);
nand U9333 (N_9333,N_8153,N_8488);
or U9334 (N_9334,N_8081,N_8253);
and U9335 (N_9335,N_8611,N_8715);
nand U9336 (N_9336,N_8916,N_8092);
nand U9337 (N_9337,N_8974,N_8528);
nor U9338 (N_9338,N_8046,N_8914);
and U9339 (N_9339,N_8711,N_8554);
nand U9340 (N_9340,N_8523,N_8052);
nor U9341 (N_9341,N_8912,N_8816);
nor U9342 (N_9342,N_8406,N_8331);
nor U9343 (N_9343,N_8002,N_8751);
nor U9344 (N_9344,N_8154,N_8076);
and U9345 (N_9345,N_8178,N_8429);
nand U9346 (N_9346,N_8813,N_8213);
or U9347 (N_9347,N_8320,N_8396);
or U9348 (N_9348,N_8806,N_8612);
and U9349 (N_9349,N_8365,N_8732);
and U9350 (N_9350,N_8469,N_8383);
nor U9351 (N_9351,N_8610,N_8324);
nor U9352 (N_9352,N_8134,N_8087);
or U9353 (N_9353,N_8642,N_8215);
or U9354 (N_9354,N_8707,N_8053);
nor U9355 (N_9355,N_8989,N_8727);
nand U9356 (N_9356,N_8392,N_8452);
xnor U9357 (N_9357,N_8825,N_8316);
nand U9358 (N_9358,N_8870,N_8023);
nand U9359 (N_9359,N_8176,N_8637);
xnor U9360 (N_9360,N_8074,N_8582);
and U9361 (N_9361,N_8591,N_8372);
or U9362 (N_9362,N_8657,N_8955);
or U9363 (N_9363,N_8014,N_8376);
or U9364 (N_9364,N_8247,N_8440);
nand U9365 (N_9365,N_8272,N_8343);
nor U9366 (N_9366,N_8797,N_8761);
or U9367 (N_9367,N_8025,N_8346);
xor U9368 (N_9368,N_8148,N_8017);
xnor U9369 (N_9369,N_8785,N_8086);
xor U9370 (N_9370,N_8164,N_8754);
nand U9371 (N_9371,N_8563,N_8445);
nor U9372 (N_9372,N_8494,N_8801);
and U9373 (N_9373,N_8856,N_8517);
nand U9374 (N_9374,N_8822,N_8901);
or U9375 (N_9375,N_8296,N_8658);
xor U9376 (N_9376,N_8793,N_8160);
or U9377 (N_9377,N_8398,N_8839);
and U9378 (N_9378,N_8996,N_8675);
and U9379 (N_9379,N_8622,N_8654);
nor U9380 (N_9380,N_8151,N_8275);
xnor U9381 (N_9381,N_8075,N_8647);
xnor U9382 (N_9382,N_8665,N_8241);
xnor U9383 (N_9383,N_8260,N_8277);
nor U9384 (N_9384,N_8308,N_8526);
and U9385 (N_9385,N_8470,N_8576);
nor U9386 (N_9386,N_8978,N_8113);
and U9387 (N_9387,N_8868,N_8892);
or U9388 (N_9388,N_8348,N_8506);
nor U9389 (N_9389,N_8845,N_8597);
nor U9390 (N_9390,N_8245,N_8792);
xor U9391 (N_9391,N_8606,N_8794);
nand U9392 (N_9392,N_8841,N_8828);
xnor U9393 (N_9393,N_8880,N_8708);
xnor U9394 (N_9394,N_8288,N_8312);
nor U9395 (N_9395,N_8394,N_8354);
xnor U9396 (N_9396,N_8678,N_8489);
xor U9397 (N_9397,N_8667,N_8476);
nor U9398 (N_9398,N_8313,N_8926);
nand U9399 (N_9399,N_8483,N_8292);
and U9400 (N_9400,N_8262,N_8467);
nand U9401 (N_9401,N_8884,N_8035);
or U9402 (N_9402,N_8929,N_8230);
or U9403 (N_9403,N_8114,N_8545);
nor U9404 (N_9404,N_8226,N_8689);
and U9405 (N_9405,N_8960,N_8079);
xor U9406 (N_9406,N_8300,N_8221);
xnor U9407 (N_9407,N_8819,N_8034);
or U9408 (N_9408,N_8687,N_8976);
and U9409 (N_9409,N_8172,N_8555);
or U9410 (N_9410,N_8969,N_8621);
xnor U9411 (N_9411,N_8810,N_8337);
xor U9412 (N_9412,N_8188,N_8290);
nand U9413 (N_9413,N_8311,N_8306);
nand U9414 (N_9414,N_8168,N_8425);
nand U9415 (N_9415,N_8301,N_8843);
nor U9416 (N_9416,N_8607,N_8847);
xor U9417 (N_9417,N_8217,N_8895);
or U9418 (N_9418,N_8084,N_8568);
nor U9419 (N_9419,N_8090,N_8395);
and U9420 (N_9420,N_8477,N_8709);
or U9421 (N_9421,N_8886,N_8249);
and U9422 (N_9422,N_8484,N_8890);
nor U9423 (N_9423,N_8010,N_8511);
nor U9424 (N_9424,N_8408,N_8340);
or U9425 (N_9425,N_8512,N_8096);
and U9426 (N_9426,N_8244,N_8688);
or U9427 (N_9427,N_8389,N_8433);
and U9428 (N_9428,N_8479,N_8844);
xor U9429 (N_9429,N_8583,N_8173);
xnor U9430 (N_9430,N_8937,N_8118);
and U9431 (N_9431,N_8680,N_8719);
and U9432 (N_9432,N_8698,N_8752);
nand U9433 (N_9433,N_8881,N_8620);
nand U9434 (N_9434,N_8202,N_8141);
xnor U9435 (N_9435,N_8347,N_8873);
or U9436 (N_9436,N_8723,N_8559);
nor U9437 (N_9437,N_8624,N_8747);
nor U9438 (N_9438,N_8001,N_8115);
nor U9439 (N_9439,N_8487,N_8449);
nand U9440 (N_9440,N_8765,N_8718);
nand U9441 (N_9441,N_8683,N_8303);
nor U9442 (N_9442,N_8238,N_8869);
nor U9443 (N_9443,N_8875,N_8903);
nor U9444 (N_9444,N_8950,N_8434);
or U9445 (N_9445,N_8330,N_8681);
and U9446 (N_9446,N_8502,N_8888);
nor U9447 (N_9447,N_8696,N_8257);
nand U9448 (N_9448,N_8235,N_8636);
nand U9449 (N_9449,N_8140,N_8513);
nand U9450 (N_9450,N_8817,N_8055);
nor U9451 (N_9451,N_8285,N_8109);
or U9452 (N_9452,N_8643,N_8130);
nand U9453 (N_9453,N_8949,N_8104);
nand U9454 (N_9454,N_8447,N_8298);
nand U9455 (N_9455,N_8863,N_8788);
xor U9456 (N_9456,N_8382,N_8632);
or U9457 (N_9457,N_8196,N_8264);
nand U9458 (N_9458,N_8102,N_8578);
xnor U9459 (N_9459,N_8529,N_8781);
nor U9460 (N_9460,N_8706,N_8064);
xnor U9461 (N_9461,N_8388,N_8029);
and U9462 (N_9462,N_8475,N_8294);
nor U9463 (N_9463,N_8739,N_8931);
nand U9464 (N_9464,N_8849,N_8295);
xnor U9465 (N_9465,N_8712,N_8332);
nor U9466 (N_9466,N_8725,N_8701);
or U9467 (N_9467,N_8009,N_8393);
nor U9468 (N_9468,N_8231,N_8826);
or U9469 (N_9469,N_8360,N_8112);
xnor U9470 (N_9470,N_8534,N_8205);
xor U9471 (N_9471,N_8980,N_8874);
xnor U9472 (N_9472,N_8358,N_8158);
nand U9473 (N_9473,N_8144,N_8557);
nand U9474 (N_9474,N_8426,N_8587);
and U9475 (N_9475,N_8923,N_8581);
or U9476 (N_9476,N_8773,N_8351);
xor U9477 (N_9477,N_8774,N_8656);
nor U9478 (N_9478,N_8420,N_8651);
nor U9479 (N_9479,N_8961,N_8566);
nand U9480 (N_9480,N_8741,N_8157);
and U9481 (N_9481,N_8572,N_8411);
nand U9482 (N_9482,N_8808,N_8307);
or U9483 (N_9483,N_8326,N_8206);
xor U9484 (N_9484,N_8103,N_8016);
nand U9485 (N_9485,N_8302,N_8355);
nand U9486 (N_9486,N_8623,N_8943);
and U9487 (N_9487,N_8276,N_8787);
nand U9488 (N_9488,N_8056,N_8925);
xor U9489 (N_9489,N_8366,N_8749);
nor U9490 (N_9490,N_8267,N_8982);
xnor U9491 (N_9491,N_8927,N_8101);
xor U9492 (N_9492,N_8956,N_8855);
nor U9493 (N_9493,N_8291,N_8983);
or U9494 (N_9494,N_8945,N_8089);
and U9495 (N_9495,N_8126,N_8516);
nor U9496 (N_9496,N_8691,N_8435);
xor U9497 (N_9497,N_8216,N_8735);
nand U9498 (N_9498,N_8100,N_8550);
nor U9499 (N_9499,N_8538,N_8853);
or U9500 (N_9500,N_8488,N_8684);
nor U9501 (N_9501,N_8818,N_8230);
nor U9502 (N_9502,N_8928,N_8229);
or U9503 (N_9503,N_8275,N_8711);
and U9504 (N_9504,N_8021,N_8934);
or U9505 (N_9505,N_8566,N_8755);
and U9506 (N_9506,N_8812,N_8894);
nor U9507 (N_9507,N_8909,N_8010);
or U9508 (N_9508,N_8092,N_8988);
nor U9509 (N_9509,N_8642,N_8832);
xnor U9510 (N_9510,N_8433,N_8261);
nor U9511 (N_9511,N_8286,N_8737);
nand U9512 (N_9512,N_8743,N_8788);
nor U9513 (N_9513,N_8217,N_8257);
xor U9514 (N_9514,N_8129,N_8120);
xnor U9515 (N_9515,N_8310,N_8623);
or U9516 (N_9516,N_8893,N_8624);
and U9517 (N_9517,N_8909,N_8351);
xnor U9518 (N_9518,N_8921,N_8716);
nor U9519 (N_9519,N_8541,N_8067);
nand U9520 (N_9520,N_8635,N_8776);
or U9521 (N_9521,N_8261,N_8121);
and U9522 (N_9522,N_8832,N_8310);
nor U9523 (N_9523,N_8055,N_8326);
and U9524 (N_9524,N_8628,N_8600);
and U9525 (N_9525,N_8908,N_8053);
and U9526 (N_9526,N_8545,N_8122);
or U9527 (N_9527,N_8158,N_8365);
or U9528 (N_9528,N_8062,N_8518);
nand U9529 (N_9529,N_8689,N_8531);
nand U9530 (N_9530,N_8168,N_8745);
xnor U9531 (N_9531,N_8188,N_8000);
nand U9532 (N_9532,N_8598,N_8896);
nand U9533 (N_9533,N_8223,N_8091);
nor U9534 (N_9534,N_8688,N_8389);
nor U9535 (N_9535,N_8323,N_8857);
or U9536 (N_9536,N_8035,N_8647);
nand U9537 (N_9537,N_8528,N_8841);
nand U9538 (N_9538,N_8136,N_8590);
nand U9539 (N_9539,N_8158,N_8602);
nand U9540 (N_9540,N_8422,N_8245);
nand U9541 (N_9541,N_8492,N_8673);
nand U9542 (N_9542,N_8150,N_8695);
nor U9543 (N_9543,N_8590,N_8857);
nor U9544 (N_9544,N_8825,N_8191);
nor U9545 (N_9545,N_8700,N_8521);
and U9546 (N_9546,N_8872,N_8576);
xnor U9547 (N_9547,N_8748,N_8328);
nor U9548 (N_9548,N_8665,N_8071);
xnor U9549 (N_9549,N_8441,N_8895);
and U9550 (N_9550,N_8796,N_8078);
or U9551 (N_9551,N_8489,N_8482);
and U9552 (N_9552,N_8944,N_8597);
nor U9553 (N_9553,N_8615,N_8737);
nor U9554 (N_9554,N_8176,N_8813);
or U9555 (N_9555,N_8462,N_8500);
nand U9556 (N_9556,N_8964,N_8099);
nand U9557 (N_9557,N_8581,N_8224);
xnor U9558 (N_9558,N_8061,N_8080);
and U9559 (N_9559,N_8659,N_8664);
xnor U9560 (N_9560,N_8800,N_8012);
and U9561 (N_9561,N_8496,N_8015);
nand U9562 (N_9562,N_8921,N_8670);
xor U9563 (N_9563,N_8143,N_8751);
nand U9564 (N_9564,N_8757,N_8336);
or U9565 (N_9565,N_8292,N_8921);
nor U9566 (N_9566,N_8274,N_8307);
nor U9567 (N_9567,N_8105,N_8745);
and U9568 (N_9568,N_8101,N_8049);
or U9569 (N_9569,N_8210,N_8190);
and U9570 (N_9570,N_8175,N_8352);
xnor U9571 (N_9571,N_8022,N_8718);
nor U9572 (N_9572,N_8690,N_8041);
nor U9573 (N_9573,N_8148,N_8344);
nand U9574 (N_9574,N_8383,N_8556);
nand U9575 (N_9575,N_8916,N_8528);
nor U9576 (N_9576,N_8959,N_8402);
nand U9577 (N_9577,N_8176,N_8368);
nand U9578 (N_9578,N_8856,N_8559);
or U9579 (N_9579,N_8895,N_8630);
xnor U9580 (N_9580,N_8439,N_8232);
and U9581 (N_9581,N_8113,N_8805);
nor U9582 (N_9582,N_8306,N_8523);
nor U9583 (N_9583,N_8072,N_8840);
or U9584 (N_9584,N_8570,N_8565);
or U9585 (N_9585,N_8131,N_8101);
or U9586 (N_9586,N_8558,N_8555);
nor U9587 (N_9587,N_8731,N_8567);
xnor U9588 (N_9588,N_8842,N_8041);
xnor U9589 (N_9589,N_8162,N_8466);
xor U9590 (N_9590,N_8146,N_8242);
xnor U9591 (N_9591,N_8138,N_8742);
nor U9592 (N_9592,N_8828,N_8074);
xnor U9593 (N_9593,N_8981,N_8272);
or U9594 (N_9594,N_8748,N_8980);
and U9595 (N_9595,N_8711,N_8141);
xor U9596 (N_9596,N_8118,N_8954);
nand U9597 (N_9597,N_8697,N_8801);
nor U9598 (N_9598,N_8167,N_8343);
and U9599 (N_9599,N_8637,N_8594);
nand U9600 (N_9600,N_8021,N_8310);
nor U9601 (N_9601,N_8224,N_8754);
nand U9602 (N_9602,N_8420,N_8060);
and U9603 (N_9603,N_8634,N_8133);
nand U9604 (N_9604,N_8675,N_8772);
xnor U9605 (N_9605,N_8175,N_8644);
nand U9606 (N_9606,N_8821,N_8961);
and U9607 (N_9607,N_8583,N_8227);
xor U9608 (N_9608,N_8636,N_8958);
xnor U9609 (N_9609,N_8029,N_8019);
nand U9610 (N_9610,N_8824,N_8658);
xnor U9611 (N_9611,N_8104,N_8684);
nand U9612 (N_9612,N_8962,N_8708);
nor U9613 (N_9613,N_8868,N_8267);
and U9614 (N_9614,N_8483,N_8926);
nor U9615 (N_9615,N_8914,N_8447);
nor U9616 (N_9616,N_8826,N_8498);
and U9617 (N_9617,N_8115,N_8617);
nand U9618 (N_9618,N_8029,N_8562);
xnor U9619 (N_9619,N_8652,N_8149);
nor U9620 (N_9620,N_8778,N_8772);
and U9621 (N_9621,N_8989,N_8417);
xnor U9622 (N_9622,N_8542,N_8013);
xnor U9623 (N_9623,N_8700,N_8061);
or U9624 (N_9624,N_8259,N_8316);
nor U9625 (N_9625,N_8017,N_8328);
or U9626 (N_9626,N_8650,N_8391);
nor U9627 (N_9627,N_8050,N_8375);
and U9628 (N_9628,N_8491,N_8531);
xor U9629 (N_9629,N_8085,N_8482);
and U9630 (N_9630,N_8573,N_8281);
nor U9631 (N_9631,N_8023,N_8730);
xnor U9632 (N_9632,N_8730,N_8967);
nand U9633 (N_9633,N_8238,N_8141);
xor U9634 (N_9634,N_8480,N_8885);
nor U9635 (N_9635,N_8425,N_8542);
xnor U9636 (N_9636,N_8249,N_8237);
xnor U9637 (N_9637,N_8326,N_8114);
nor U9638 (N_9638,N_8327,N_8138);
xnor U9639 (N_9639,N_8251,N_8932);
and U9640 (N_9640,N_8720,N_8139);
or U9641 (N_9641,N_8609,N_8126);
nor U9642 (N_9642,N_8305,N_8216);
and U9643 (N_9643,N_8404,N_8515);
nor U9644 (N_9644,N_8170,N_8563);
nand U9645 (N_9645,N_8063,N_8798);
nor U9646 (N_9646,N_8665,N_8128);
xnor U9647 (N_9647,N_8999,N_8038);
and U9648 (N_9648,N_8657,N_8910);
or U9649 (N_9649,N_8664,N_8738);
nor U9650 (N_9650,N_8218,N_8297);
nand U9651 (N_9651,N_8754,N_8948);
or U9652 (N_9652,N_8242,N_8522);
nor U9653 (N_9653,N_8454,N_8973);
nand U9654 (N_9654,N_8877,N_8794);
or U9655 (N_9655,N_8820,N_8995);
and U9656 (N_9656,N_8979,N_8185);
or U9657 (N_9657,N_8233,N_8540);
xor U9658 (N_9658,N_8219,N_8880);
nor U9659 (N_9659,N_8700,N_8796);
nor U9660 (N_9660,N_8140,N_8517);
and U9661 (N_9661,N_8879,N_8251);
or U9662 (N_9662,N_8875,N_8122);
and U9663 (N_9663,N_8430,N_8201);
nor U9664 (N_9664,N_8769,N_8374);
nand U9665 (N_9665,N_8360,N_8563);
nor U9666 (N_9666,N_8578,N_8081);
and U9667 (N_9667,N_8563,N_8664);
and U9668 (N_9668,N_8617,N_8932);
nor U9669 (N_9669,N_8943,N_8740);
nand U9670 (N_9670,N_8321,N_8981);
nand U9671 (N_9671,N_8281,N_8422);
nand U9672 (N_9672,N_8406,N_8356);
xor U9673 (N_9673,N_8156,N_8433);
xor U9674 (N_9674,N_8942,N_8969);
xnor U9675 (N_9675,N_8093,N_8215);
and U9676 (N_9676,N_8505,N_8114);
or U9677 (N_9677,N_8009,N_8028);
xor U9678 (N_9678,N_8150,N_8257);
and U9679 (N_9679,N_8280,N_8700);
xor U9680 (N_9680,N_8651,N_8831);
nand U9681 (N_9681,N_8943,N_8734);
or U9682 (N_9682,N_8809,N_8556);
and U9683 (N_9683,N_8549,N_8172);
or U9684 (N_9684,N_8276,N_8918);
and U9685 (N_9685,N_8640,N_8387);
xnor U9686 (N_9686,N_8359,N_8035);
nor U9687 (N_9687,N_8085,N_8214);
xnor U9688 (N_9688,N_8735,N_8881);
xnor U9689 (N_9689,N_8790,N_8004);
and U9690 (N_9690,N_8889,N_8295);
xnor U9691 (N_9691,N_8451,N_8937);
or U9692 (N_9692,N_8090,N_8289);
xnor U9693 (N_9693,N_8935,N_8565);
nand U9694 (N_9694,N_8776,N_8345);
or U9695 (N_9695,N_8111,N_8804);
xnor U9696 (N_9696,N_8453,N_8676);
xnor U9697 (N_9697,N_8644,N_8337);
or U9698 (N_9698,N_8560,N_8634);
and U9699 (N_9699,N_8672,N_8415);
and U9700 (N_9700,N_8390,N_8173);
xor U9701 (N_9701,N_8319,N_8550);
and U9702 (N_9702,N_8736,N_8287);
xnor U9703 (N_9703,N_8423,N_8942);
xor U9704 (N_9704,N_8368,N_8337);
nand U9705 (N_9705,N_8548,N_8994);
or U9706 (N_9706,N_8437,N_8345);
and U9707 (N_9707,N_8599,N_8147);
and U9708 (N_9708,N_8305,N_8061);
nor U9709 (N_9709,N_8872,N_8417);
xnor U9710 (N_9710,N_8492,N_8603);
nand U9711 (N_9711,N_8071,N_8460);
xor U9712 (N_9712,N_8511,N_8774);
and U9713 (N_9713,N_8883,N_8481);
or U9714 (N_9714,N_8090,N_8216);
and U9715 (N_9715,N_8907,N_8232);
and U9716 (N_9716,N_8832,N_8298);
or U9717 (N_9717,N_8579,N_8524);
and U9718 (N_9718,N_8090,N_8036);
nor U9719 (N_9719,N_8239,N_8025);
and U9720 (N_9720,N_8335,N_8430);
or U9721 (N_9721,N_8541,N_8247);
or U9722 (N_9722,N_8176,N_8155);
nand U9723 (N_9723,N_8558,N_8878);
or U9724 (N_9724,N_8102,N_8862);
or U9725 (N_9725,N_8587,N_8049);
or U9726 (N_9726,N_8369,N_8774);
or U9727 (N_9727,N_8126,N_8789);
or U9728 (N_9728,N_8784,N_8990);
nor U9729 (N_9729,N_8780,N_8390);
nor U9730 (N_9730,N_8137,N_8647);
nor U9731 (N_9731,N_8662,N_8580);
nor U9732 (N_9732,N_8125,N_8109);
xnor U9733 (N_9733,N_8731,N_8114);
and U9734 (N_9734,N_8632,N_8710);
nor U9735 (N_9735,N_8786,N_8355);
nor U9736 (N_9736,N_8454,N_8513);
or U9737 (N_9737,N_8228,N_8507);
xnor U9738 (N_9738,N_8894,N_8349);
xnor U9739 (N_9739,N_8666,N_8926);
or U9740 (N_9740,N_8691,N_8239);
and U9741 (N_9741,N_8463,N_8096);
and U9742 (N_9742,N_8046,N_8496);
and U9743 (N_9743,N_8886,N_8198);
and U9744 (N_9744,N_8059,N_8274);
and U9745 (N_9745,N_8498,N_8167);
nor U9746 (N_9746,N_8185,N_8925);
and U9747 (N_9747,N_8636,N_8775);
nor U9748 (N_9748,N_8380,N_8432);
and U9749 (N_9749,N_8358,N_8389);
and U9750 (N_9750,N_8758,N_8400);
or U9751 (N_9751,N_8314,N_8507);
xor U9752 (N_9752,N_8778,N_8836);
or U9753 (N_9753,N_8860,N_8999);
nand U9754 (N_9754,N_8580,N_8571);
nor U9755 (N_9755,N_8357,N_8593);
nor U9756 (N_9756,N_8225,N_8242);
or U9757 (N_9757,N_8826,N_8593);
or U9758 (N_9758,N_8255,N_8003);
or U9759 (N_9759,N_8979,N_8175);
xor U9760 (N_9760,N_8715,N_8785);
nor U9761 (N_9761,N_8906,N_8184);
or U9762 (N_9762,N_8446,N_8306);
or U9763 (N_9763,N_8195,N_8275);
nor U9764 (N_9764,N_8662,N_8605);
nand U9765 (N_9765,N_8824,N_8281);
and U9766 (N_9766,N_8659,N_8346);
or U9767 (N_9767,N_8478,N_8832);
nor U9768 (N_9768,N_8233,N_8361);
and U9769 (N_9769,N_8822,N_8762);
nor U9770 (N_9770,N_8988,N_8851);
or U9771 (N_9771,N_8398,N_8182);
or U9772 (N_9772,N_8405,N_8448);
xnor U9773 (N_9773,N_8954,N_8374);
nand U9774 (N_9774,N_8520,N_8669);
and U9775 (N_9775,N_8928,N_8793);
nor U9776 (N_9776,N_8095,N_8806);
nand U9777 (N_9777,N_8218,N_8778);
and U9778 (N_9778,N_8474,N_8271);
nor U9779 (N_9779,N_8128,N_8735);
nor U9780 (N_9780,N_8548,N_8217);
nor U9781 (N_9781,N_8975,N_8133);
nor U9782 (N_9782,N_8228,N_8368);
nor U9783 (N_9783,N_8553,N_8810);
xnor U9784 (N_9784,N_8581,N_8492);
xnor U9785 (N_9785,N_8562,N_8664);
and U9786 (N_9786,N_8547,N_8722);
xor U9787 (N_9787,N_8809,N_8558);
xor U9788 (N_9788,N_8598,N_8183);
xnor U9789 (N_9789,N_8889,N_8435);
or U9790 (N_9790,N_8818,N_8018);
xor U9791 (N_9791,N_8025,N_8910);
and U9792 (N_9792,N_8738,N_8845);
xor U9793 (N_9793,N_8805,N_8924);
nor U9794 (N_9794,N_8869,N_8384);
nor U9795 (N_9795,N_8430,N_8548);
and U9796 (N_9796,N_8950,N_8316);
xor U9797 (N_9797,N_8287,N_8551);
nand U9798 (N_9798,N_8103,N_8369);
xor U9799 (N_9799,N_8023,N_8995);
nor U9800 (N_9800,N_8660,N_8498);
and U9801 (N_9801,N_8635,N_8134);
nor U9802 (N_9802,N_8122,N_8241);
xnor U9803 (N_9803,N_8908,N_8093);
xnor U9804 (N_9804,N_8323,N_8331);
and U9805 (N_9805,N_8968,N_8571);
nand U9806 (N_9806,N_8847,N_8177);
or U9807 (N_9807,N_8330,N_8103);
or U9808 (N_9808,N_8610,N_8483);
nand U9809 (N_9809,N_8917,N_8987);
xnor U9810 (N_9810,N_8009,N_8672);
xnor U9811 (N_9811,N_8138,N_8109);
and U9812 (N_9812,N_8199,N_8258);
nor U9813 (N_9813,N_8114,N_8617);
xor U9814 (N_9814,N_8549,N_8613);
xor U9815 (N_9815,N_8217,N_8798);
nand U9816 (N_9816,N_8537,N_8985);
nor U9817 (N_9817,N_8357,N_8321);
xnor U9818 (N_9818,N_8922,N_8175);
nor U9819 (N_9819,N_8974,N_8098);
nor U9820 (N_9820,N_8483,N_8841);
xnor U9821 (N_9821,N_8946,N_8818);
nor U9822 (N_9822,N_8999,N_8159);
xor U9823 (N_9823,N_8057,N_8833);
or U9824 (N_9824,N_8761,N_8535);
or U9825 (N_9825,N_8080,N_8103);
nor U9826 (N_9826,N_8718,N_8579);
nor U9827 (N_9827,N_8443,N_8125);
nor U9828 (N_9828,N_8394,N_8595);
nand U9829 (N_9829,N_8413,N_8322);
nand U9830 (N_9830,N_8496,N_8845);
or U9831 (N_9831,N_8771,N_8474);
nor U9832 (N_9832,N_8046,N_8997);
and U9833 (N_9833,N_8968,N_8875);
xor U9834 (N_9834,N_8133,N_8627);
and U9835 (N_9835,N_8945,N_8799);
or U9836 (N_9836,N_8530,N_8302);
xor U9837 (N_9837,N_8078,N_8300);
xor U9838 (N_9838,N_8722,N_8057);
and U9839 (N_9839,N_8847,N_8948);
nand U9840 (N_9840,N_8944,N_8242);
xnor U9841 (N_9841,N_8756,N_8629);
or U9842 (N_9842,N_8156,N_8115);
and U9843 (N_9843,N_8323,N_8900);
and U9844 (N_9844,N_8771,N_8284);
nor U9845 (N_9845,N_8895,N_8197);
xnor U9846 (N_9846,N_8298,N_8164);
nor U9847 (N_9847,N_8631,N_8123);
nand U9848 (N_9848,N_8428,N_8616);
xnor U9849 (N_9849,N_8886,N_8032);
xor U9850 (N_9850,N_8484,N_8513);
and U9851 (N_9851,N_8590,N_8150);
xor U9852 (N_9852,N_8343,N_8836);
xor U9853 (N_9853,N_8745,N_8620);
nor U9854 (N_9854,N_8540,N_8118);
and U9855 (N_9855,N_8821,N_8633);
nor U9856 (N_9856,N_8500,N_8833);
nor U9857 (N_9857,N_8004,N_8739);
nand U9858 (N_9858,N_8546,N_8725);
and U9859 (N_9859,N_8358,N_8227);
nor U9860 (N_9860,N_8687,N_8063);
nand U9861 (N_9861,N_8980,N_8785);
xnor U9862 (N_9862,N_8367,N_8931);
nand U9863 (N_9863,N_8909,N_8163);
nand U9864 (N_9864,N_8266,N_8099);
nor U9865 (N_9865,N_8545,N_8400);
or U9866 (N_9866,N_8722,N_8673);
and U9867 (N_9867,N_8093,N_8710);
nand U9868 (N_9868,N_8347,N_8737);
or U9869 (N_9869,N_8911,N_8478);
or U9870 (N_9870,N_8494,N_8865);
nand U9871 (N_9871,N_8060,N_8477);
or U9872 (N_9872,N_8515,N_8908);
xnor U9873 (N_9873,N_8957,N_8823);
nand U9874 (N_9874,N_8400,N_8553);
nor U9875 (N_9875,N_8422,N_8879);
or U9876 (N_9876,N_8790,N_8049);
and U9877 (N_9877,N_8800,N_8456);
nor U9878 (N_9878,N_8550,N_8414);
and U9879 (N_9879,N_8378,N_8418);
or U9880 (N_9880,N_8486,N_8755);
or U9881 (N_9881,N_8396,N_8775);
or U9882 (N_9882,N_8141,N_8700);
xnor U9883 (N_9883,N_8617,N_8392);
nand U9884 (N_9884,N_8820,N_8827);
nor U9885 (N_9885,N_8635,N_8092);
or U9886 (N_9886,N_8144,N_8695);
xnor U9887 (N_9887,N_8811,N_8260);
and U9888 (N_9888,N_8371,N_8729);
and U9889 (N_9889,N_8236,N_8016);
nand U9890 (N_9890,N_8907,N_8296);
nor U9891 (N_9891,N_8303,N_8116);
nand U9892 (N_9892,N_8504,N_8243);
and U9893 (N_9893,N_8557,N_8474);
and U9894 (N_9894,N_8330,N_8648);
and U9895 (N_9895,N_8541,N_8092);
nand U9896 (N_9896,N_8595,N_8246);
nand U9897 (N_9897,N_8288,N_8425);
nor U9898 (N_9898,N_8532,N_8732);
nand U9899 (N_9899,N_8527,N_8155);
or U9900 (N_9900,N_8614,N_8798);
xnor U9901 (N_9901,N_8282,N_8870);
nand U9902 (N_9902,N_8370,N_8567);
xor U9903 (N_9903,N_8639,N_8596);
and U9904 (N_9904,N_8105,N_8600);
and U9905 (N_9905,N_8215,N_8722);
or U9906 (N_9906,N_8015,N_8345);
or U9907 (N_9907,N_8791,N_8665);
nor U9908 (N_9908,N_8371,N_8591);
nand U9909 (N_9909,N_8407,N_8354);
or U9910 (N_9910,N_8193,N_8620);
xor U9911 (N_9911,N_8159,N_8786);
xnor U9912 (N_9912,N_8117,N_8815);
and U9913 (N_9913,N_8225,N_8297);
xnor U9914 (N_9914,N_8101,N_8023);
nor U9915 (N_9915,N_8629,N_8273);
nand U9916 (N_9916,N_8501,N_8741);
or U9917 (N_9917,N_8851,N_8269);
or U9918 (N_9918,N_8009,N_8678);
nand U9919 (N_9919,N_8171,N_8459);
xnor U9920 (N_9920,N_8999,N_8319);
xnor U9921 (N_9921,N_8250,N_8827);
xnor U9922 (N_9922,N_8345,N_8788);
xor U9923 (N_9923,N_8379,N_8450);
nor U9924 (N_9924,N_8001,N_8037);
nand U9925 (N_9925,N_8979,N_8103);
nor U9926 (N_9926,N_8608,N_8799);
and U9927 (N_9927,N_8186,N_8918);
nor U9928 (N_9928,N_8142,N_8664);
nand U9929 (N_9929,N_8374,N_8201);
and U9930 (N_9930,N_8854,N_8786);
nand U9931 (N_9931,N_8895,N_8774);
or U9932 (N_9932,N_8876,N_8050);
nor U9933 (N_9933,N_8389,N_8770);
and U9934 (N_9934,N_8649,N_8284);
nor U9935 (N_9935,N_8894,N_8260);
nor U9936 (N_9936,N_8416,N_8749);
nor U9937 (N_9937,N_8047,N_8671);
nor U9938 (N_9938,N_8512,N_8152);
or U9939 (N_9939,N_8762,N_8834);
or U9940 (N_9940,N_8768,N_8279);
nand U9941 (N_9941,N_8968,N_8314);
and U9942 (N_9942,N_8919,N_8231);
nor U9943 (N_9943,N_8275,N_8292);
or U9944 (N_9944,N_8449,N_8522);
xor U9945 (N_9945,N_8494,N_8084);
or U9946 (N_9946,N_8267,N_8166);
or U9947 (N_9947,N_8838,N_8329);
nand U9948 (N_9948,N_8907,N_8407);
nand U9949 (N_9949,N_8907,N_8487);
and U9950 (N_9950,N_8946,N_8316);
nand U9951 (N_9951,N_8529,N_8881);
and U9952 (N_9952,N_8432,N_8902);
and U9953 (N_9953,N_8554,N_8875);
nor U9954 (N_9954,N_8198,N_8473);
or U9955 (N_9955,N_8151,N_8838);
nand U9956 (N_9956,N_8909,N_8082);
and U9957 (N_9957,N_8945,N_8926);
nand U9958 (N_9958,N_8364,N_8321);
nor U9959 (N_9959,N_8565,N_8887);
nand U9960 (N_9960,N_8839,N_8022);
and U9961 (N_9961,N_8993,N_8053);
xnor U9962 (N_9962,N_8074,N_8023);
or U9963 (N_9963,N_8701,N_8551);
nor U9964 (N_9964,N_8821,N_8379);
or U9965 (N_9965,N_8458,N_8576);
nand U9966 (N_9966,N_8988,N_8434);
xor U9967 (N_9967,N_8353,N_8332);
xnor U9968 (N_9968,N_8189,N_8908);
and U9969 (N_9969,N_8532,N_8890);
nor U9970 (N_9970,N_8374,N_8040);
nor U9971 (N_9971,N_8367,N_8447);
nor U9972 (N_9972,N_8336,N_8569);
nor U9973 (N_9973,N_8999,N_8529);
nand U9974 (N_9974,N_8863,N_8240);
xor U9975 (N_9975,N_8816,N_8337);
nand U9976 (N_9976,N_8074,N_8880);
nor U9977 (N_9977,N_8149,N_8916);
nor U9978 (N_9978,N_8801,N_8589);
and U9979 (N_9979,N_8444,N_8371);
nor U9980 (N_9980,N_8514,N_8052);
nand U9981 (N_9981,N_8611,N_8431);
and U9982 (N_9982,N_8103,N_8703);
xnor U9983 (N_9983,N_8369,N_8800);
xor U9984 (N_9984,N_8202,N_8282);
nor U9985 (N_9985,N_8986,N_8595);
nor U9986 (N_9986,N_8768,N_8750);
xnor U9987 (N_9987,N_8749,N_8443);
or U9988 (N_9988,N_8178,N_8740);
xnor U9989 (N_9989,N_8040,N_8956);
xor U9990 (N_9990,N_8503,N_8480);
nand U9991 (N_9991,N_8732,N_8449);
xor U9992 (N_9992,N_8351,N_8159);
or U9993 (N_9993,N_8583,N_8391);
and U9994 (N_9994,N_8013,N_8854);
nand U9995 (N_9995,N_8257,N_8793);
xor U9996 (N_9996,N_8102,N_8332);
nand U9997 (N_9997,N_8342,N_8166);
or U9998 (N_9998,N_8186,N_8863);
and U9999 (N_9999,N_8494,N_8245);
nor U10000 (N_10000,N_9627,N_9565);
or U10001 (N_10001,N_9856,N_9870);
nand U10002 (N_10002,N_9062,N_9551);
xor U10003 (N_10003,N_9135,N_9249);
or U10004 (N_10004,N_9746,N_9027);
and U10005 (N_10005,N_9813,N_9507);
nand U10006 (N_10006,N_9344,N_9465);
or U10007 (N_10007,N_9968,N_9660);
nand U10008 (N_10008,N_9191,N_9212);
nor U10009 (N_10009,N_9635,N_9085);
or U10010 (N_10010,N_9791,N_9207);
or U10011 (N_10011,N_9236,N_9313);
or U10012 (N_10012,N_9527,N_9462);
or U10013 (N_10013,N_9431,N_9332);
and U10014 (N_10014,N_9869,N_9484);
nor U10015 (N_10015,N_9524,N_9785);
xnor U10016 (N_10016,N_9984,N_9742);
nor U10017 (N_10017,N_9826,N_9975);
xor U10018 (N_10018,N_9952,N_9908);
xnor U10019 (N_10019,N_9277,N_9563);
nor U10020 (N_10020,N_9807,N_9490);
and U10021 (N_10021,N_9632,N_9081);
xor U10022 (N_10022,N_9594,N_9169);
and U10023 (N_10023,N_9227,N_9156);
xnor U10024 (N_10024,N_9725,N_9113);
or U10025 (N_10025,N_9997,N_9679);
nand U10026 (N_10026,N_9841,N_9699);
or U10027 (N_10027,N_9258,N_9769);
or U10028 (N_10028,N_9314,N_9060);
xnor U10029 (N_10029,N_9363,N_9449);
nand U10030 (N_10030,N_9716,N_9437);
nor U10031 (N_10031,N_9577,N_9711);
nand U10032 (N_10032,N_9015,N_9949);
or U10033 (N_10033,N_9329,N_9357);
and U10034 (N_10034,N_9967,N_9380);
nand U10035 (N_10035,N_9090,N_9630);
or U10036 (N_10036,N_9965,N_9165);
nand U10037 (N_10037,N_9278,N_9100);
nor U10038 (N_10038,N_9487,N_9858);
nor U10039 (N_10039,N_9932,N_9787);
xnor U10040 (N_10040,N_9913,N_9803);
nor U10041 (N_10041,N_9107,N_9886);
and U10042 (N_10042,N_9446,N_9948);
and U10043 (N_10043,N_9904,N_9531);
or U10044 (N_10044,N_9341,N_9804);
and U10045 (N_10045,N_9181,N_9201);
and U10046 (N_10046,N_9405,N_9383);
xor U10047 (N_10047,N_9788,N_9628);
and U10048 (N_10048,N_9440,N_9889);
and U10049 (N_10049,N_9718,N_9571);
nand U10050 (N_10050,N_9280,N_9288);
or U10051 (N_10051,N_9159,N_9194);
or U10052 (N_10052,N_9642,N_9765);
or U10053 (N_10053,N_9110,N_9466);
nor U10054 (N_10054,N_9853,N_9616);
xnor U10055 (N_10055,N_9205,N_9456);
and U10056 (N_10056,N_9365,N_9850);
nand U10057 (N_10057,N_9820,N_9195);
nand U10058 (N_10058,N_9270,N_9663);
and U10059 (N_10059,N_9962,N_9703);
nor U10060 (N_10060,N_9482,N_9115);
nor U10061 (N_10061,N_9108,N_9372);
nor U10062 (N_10062,N_9873,N_9809);
xnor U10063 (N_10063,N_9935,N_9631);
and U10064 (N_10064,N_9289,N_9218);
nand U10065 (N_10065,N_9239,N_9874);
and U10066 (N_10066,N_9155,N_9614);
and U10067 (N_10067,N_9839,N_9384);
or U10068 (N_10068,N_9203,N_9981);
xnor U10069 (N_10069,N_9749,N_9530);
and U10070 (N_10070,N_9512,N_9994);
nand U10071 (N_10071,N_9423,N_9139);
xnor U10072 (N_10072,N_9128,N_9650);
nand U10073 (N_10073,N_9301,N_9297);
nand U10074 (N_10074,N_9596,N_9152);
nand U10075 (N_10075,N_9358,N_9223);
xnor U10076 (N_10076,N_9778,N_9681);
or U10077 (N_10077,N_9247,N_9419);
or U10078 (N_10078,N_9327,N_9202);
and U10079 (N_10079,N_9050,N_9286);
or U10080 (N_10080,N_9417,N_9736);
nand U10081 (N_10081,N_9618,N_9242);
and U10082 (N_10082,N_9306,N_9272);
and U10083 (N_10083,N_9934,N_9665);
nand U10084 (N_10084,N_9883,N_9554);
xor U10085 (N_10085,N_9517,N_9977);
and U10086 (N_10086,N_9351,N_9401);
and U10087 (N_10087,N_9215,N_9941);
or U10088 (N_10088,N_9282,N_9099);
xnor U10089 (N_10089,N_9689,N_9966);
and U10090 (N_10090,N_9399,N_9771);
nor U10091 (N_10091,N_9451,N_9368);
or U10092 (N_10092,N_9309,N_9238);
xor U10093 (N_10093,N_9037,N_9636);
nand U10094 (N_10094,N_9798,N_9498);
nand U10095 (N_10095,N_9117,N_9986);
xnor U10096 (N_10096,N_9269,N_9573);
xnor U10097 (N_10097,N_9416,N_9445);
nor U10098 (N_10098,N_9187,N_9307);
xor U10099 (N_10099,N_9095,N_9486);
xnor U10100 (N_10100,N_9353,N_9865);
xnor U10101 (N_10101,N_9658,N_9067);
nand U10102 (N_10102,N_9453,N_9505);
xor U10103 (N_10103,N_9132,N_9895);
or U10104 (N_10104,N_9519,N_9786);
xor U10105 (N_10105,N_9472,N_9338);
or U10106 (N_10106,N_9342,N_9225);
and U10107 (N_10107,N_9094,N_9056);
nor U10108 (N_10108,N_9386,N_9168);
or U10109 (N_10109,N_9285,N_9035);
nand U10110 (N_10110,N_9963,N_9879);
nor U10111 (N_10111,N_9103,N_9007);
and U10112 (N_10112,N_9295,N_9151);
xnor U10113 (N_10113,N_9240,N_9940);
or U10114 (N_10114,N_9956,N_9750);
nor U10115 (N_10115,N_9694,N_9476);
nor U10116 (N_10116,N_9305,N_9890);
nand U10117 (N_10117,N_9074,N_9544);
xor U10118 (N_10118,N_9481,N_9504);
nand U10119 (N_10119,N_9615,N_9914);
and U10120 (N_10120,N_9370,N_9947);
or U10121 (N_10121,N_9167,N_9082);
nor U10122 (N_10122,N_9292,N_9188);
and U10123 (N_10123,N_9396,N_9672);
and U10124 (N_10124,N_9989,N_9492);
and U10125 (N_10125,N_9773,N_9959);
or U10126 (N_10126,N_9510,N_9591);
and U10127 (N_10127,N_9574,N_9972);
nand U10128 (N_10128,N_9604,N_9724);
nor U10129 (N_10129,N_9092,N_9752);
xor U10130 (N_10130,N_9810,N_9979);
and U10131 (N_10131,N_9146,N_9937);
nand U10132 (N_10132,N_9998,N_9059);
and U10133 (N_10133,N_9147,N_9019);
nand U10134 (N_10134,N_9923,N_9683);
or U10135 (N_10135,N_9232,N_9177);
or U10136 (N_10136,N_9568,N_9933);
xnor U10137 (N_10137,N_9104,N_9707);
nor U10138 (N_10138,N_9776,N_9611);
or U10139 (N_10139,N_9899,N_9164);
nand U10140 (N_10140,N_9815,N_9467);
or U10141 (N_10141,N_9831,N_9267);
nor U10142 (N_10142,N_9084,N_9970);
nand U10143 (N_10143,N_9721,N_9652);
and U10144 (N_10144,N_9153,N_9974);
or U10145 (N_10145,N_9023,N_9184);
or U10146 (N_10146,N_9846,N_9144);
and U10147 (N_10147,N_9252,N_9910);
and U10148 (N_10148,N_9433,N_9730);
xnor U10149 (N_10149,N_9066,N_9311);
nor U10150 (N_10150,N_9073,N_9878);
nor U10151 (N_10151,N_9264,N_9996);
or U10152 (N_10152,N_9545,N_9633);
nor U10153 (N_10153,N_9246,N_9319);
nand U10154 (N_10154,N_9079,N_9720);
nand U10155 (N_10155,N_9045,N_9927);
nor U10156 (N_10156,N_9511,N_9009);
nand U10157 (N_10157,N_9680,N_9822);
and U10158 (N_10158,N_9438,N_9052);
xor U10159 (N_10159,N_9281,N_9101);
xnor U10160 (N_10160,N_9284,N_9584);
xnor U10161 (N_10161,N_9131,N_9158);
xnor U10162 (N_10162,N_9579,N_9180);
nor U10163 (N_10163,N_9142,N_9369);
nand U10164 (N_10164,N_9653,N_9331);
nand U10165 (N_10165,N_9199,N_9421);
nand U10166 (N_10166,N_9091,N_9034);
nand U10167 (N_10167,N_9651,N_9755);
nor U10168 (N_10168,N_9838,N_9706);
xor U10169 (N_10169,N_9414,N_9528);
or U10170 (N_10170,N_9821,N_9671);
xor U10171 (N_10171,N_9640,N_9572);
or U10172 (N_10172,N_9053,N_9439);
nor U10173 (N_10173,N_9213,N_9888);
or U10174 (N_10174,N_9595,N_9335);
nand U10175 (N_10175,N_9061,N_9273);
or U10176 (N_10176,N_9256,N_9569);
xnor U10177 (N_10177,N_9817,N_9560);
nand U10178 (N_10178,N_9794,N_9739);
xor U10179 (N_10179,N_9864,N_9491);
or U10180 (N_10180,N_9120,N_9068);
or U10181 (N_10181,N_9898,N_9536);
nor U10182 (N_10182,N_9474,N_9861);
nor U10183 (N_10183,N_9488,N_9464);
or U10184 (N_10184,N_9759,N_9069);
or U10185 (N_10185,N_9243,N_9597);
xnor U10186 (N_10186,N_9406,N_9014);
or U10187 (N_10187,N_9655,N_9602);
or U10188 (N_10188,N_9471,N_9415);
xor U10189 (N_10189,N_9389,N_9696);
or U10190 (N_10190,N_9772,N_9170);
xnor U10191 (N_10191,N_9008,N_9320);
nor U10192 (N_10192,N_9624,N_9398);
nand U10193 (N_10193,N_9098,N_9182);
or U10194 (N_10194,N_9499,N_9047);
or U10195 (N_10195,N_9782,N_9926);
or U10196 (N_10196,N_9950,N_9983);
and U10197 (N_10197,N_9859,N_9729);
nor U10198 (N_10198,N_9133,N_9478);
and U10199 (N_10199,N_9529,N_9848);
nor U10200 (N_10200,N_9221,N_9620);
nand U10201 (N_10201,N_9876,N_9029);
nand U10202 (N_10202,N_9598,N_9400);
nor U10203 (N_10203,N_9916,N_9764);
xor U10204 (N_10204,N_9121,N_9832);
or U10205 (N_10205,N_9646,N_9578);
nand U10206 (N_10206,N_9352,N_9754);
xor U10207 (N_10207,N_9262,N_9324);
nand U10208 (N_10208,N_9525,N_9961);
and U10209 (N_10209,N_9204,N_9112);
nand U10210 (N_10210,N_9796,N_9172);
nand U10211 (N_10211,N_9662,N_9586);
nor U10212 (N_10212,N_9429,N_9255);
nand U10213 (N_10213,N_9031,N_9617);
nor U10214 (N_10214,N_9290,N_9808);
or U10215 (N_10215,N_9496,N_9402);
or U10216 (N_10216,N_9346,N_9377);
and U10217 (N_10217,N_9509,N_9483);
nand U10218 (N_10218,N_9058,N_9557);
or U10219 (N_10219,N_9388,N_9792);
xnor U10220 (N_10220,N_9013,N_9863);
and U10221 (N_10221,N_9766,N_9493);
nor U10222 (N_10222,N_9534,N_9896);
nor U10223 (N_10223,N_9420,N_9312);
xor U10224 (N_10224,N_9812,N_9622);
nand U10225 (N_10225,N_9245,N_9315);
or U10226 (N_10226,N_9921,N_9828);
nand U10227 (N_10227,N_9669,N_9799);
and U10228 (N_10228,N_9709,N_9522);
and U10229 (N_10229,N_9917,N_9321);
nor U10230 (N_10230,N_9403,N_9366);
or U10231 (N_10231,N_9999,N_9691);
xor U10232 (N_10232,N_9021,N_9945);
or U10233 (N_10233,N_9376,N_9851);
xor U10234 (N_10234,N_9909,N_9452);
nand U10235 (N_10235,N_9392,N_9667);
or U10236 (N_10236,N_9763,N_9459);
and U10237 (N_10237,N_9845,N_9469);
nand U10238 (N_10238,N_9072,N_9230);
and U10239 (N_10239,N_9592,N_9955);
or U10240 (N_10240,N_9849,N_9185);
xor U10241 (N_10241,N_9685,N_9840);
or U10242 (N_10242,N_9770,N_9006);
nand U10243 (N_10243,N_9625,N_9922);
xor U10244 (N_10244,N_9608,N_9779);
xnor U10245 (N_10245,N_9753,N_9978);
and U10246 (N_10246,N_9274,N_9485);
nor U10247 (N_10247,N_9234,N_9233);
nor U10248 (N_10248,N_9263,N_9521);
or U10249 (N_10249,N_9127,N_9715);
nor U10250 (N_10250,N_9378,N_9109);
nand U10251 (N_10251,N_9265,N_9659);
or U10252 (N_10252,N_9546,N_9382);
nand U10253 (N_10253,N_9086,N_9200);
nor U10254 (N_10254,N_9600,N_9116);
and U10255 (N_10255,N_9424,N_9175);
or U10256 (N_10256,N_9244,N_9906);
or U10257 (N_10257,N_9901,N_9192);
nor U10258 (N_10258,N_9470,N_9621);
nor U10259 (N_10259,N_9538,N_9723);
nand U10260 (N_10260,N_9702,N_9783);
and U10261 (N_10261,N_9097,N_9700);
nor U10262 (N_10262,N_9251,N_9830);
nand U10263 (N_10263,N_9229,N_9532);
xor U10264 (N_10264,N_9661,N_9126);
nand U10265 (N_10265,N_9000,N_9426);
nor U10266 (N_10266,N_9427,N_9985);
nand U10267 (N_10267,N_9761,N_9017);
xnor U10268 (N_10268,N_9790,N_9743);
nor U10269 (N_10269,N_9535,N_9668);
nor U10270 (N_10270,N_9219,N_9348);
nand U10271 (N_10271,N_9148,N_9118);
xor U10272 (N_10272,N_9593,N_9196);
nand U10273 (N_10273,N_9198,N_9298);
and U10274 (N_10274,N_9322,N_9973);
xor U10275 (N_10275,N_9078,N_9951);
nor U10276 (N_10276,N_9751,N_9179);
nor U10277 (N_10277,N_9713,N_9789);
or U10278 (N_10278,N_9049,N_9408);
nand U10279 (N_10279,N_9435,N_9842);
and U10280 (N_10280,N_9684,N_9552);
nand U10281 (N_10281,N_9141,N_9434);
or U10282 (N_10282,N_9065,N_9990);
and U10283 (N_10283,N_9137,N_9777);
nand U10284 (N_10284,N_9575,N_9119);
nor U10285 (N_10285,N_9692,N_9268);
or U10286 (N_10286,N_9387,N_9174);
and U10287 (N_10287,N_9220,N_9178);
and U10288 (N_10288,N_9237,N_9728);
nor U10289 (N_10289,N_9217,N_9556);
nand U10290 (N_10290,N_9514,N_9443);
nor U10291 (N_10291,N_9409,N_9800);
nand U10292 (N_10292,N_9025,N_9825);
or U10293 (N_10293,N_9946,N_9183);
xor U10294 (N_10294,N_9964,N_9361);
nor U10295 (N_10295,N_9030,N_9458);
xnor U10296 (N_10296,N_9537,N_9385);
xnor U10297 (N_10297,N_9953,N_9677);
xor U10298 (N_10298,N_9197,N_9980);
nor U10299 (N_10299,N_9939,N_9011);
nand U10300 (N_10300,N_9075,N_9334);
or U10301 (N_10301,N_9461,N_9774);
or U10302 (N_10302,N_9735,N_9762);
xor U10303 (N_10303,N_9516,N_9339);
xor U10304 (N_10304,N_9228,N_9226);
and U10305 (N_10305,N_9515,N_9612);
or U10306 (N_10306,N_9016,N_9882);
or U10307 (N_10307,N_9533,N_9543);
nand U10308 (N_10308,N_9745,N_9374);
or U10309 (N_10309,N_9136,N_9364);
xor U10310 (N_10310,N_9824,N_9040);
nor U10311 (N_10311,N_9125,N_9410);
nor U10312 (N_10312,N_9871,N_9603);
and U10313 (N_10313,N_9077,N_9042);
xnor U10314 (N_10314,N_9930,N_9039);
and U10315 (N_10315,N_9583,N_9971);
or U10316 (N_10316,N_9623,N_9818);
xnor U10317 (N_10317,N_9071,N_9310);
xor U10318 (N_10318,N_9982,N_9737);
xor U10319 (N_10319,N_9371,N_9114);
or U10320 (N_10320,N_9350,N_9958);
nand U10321 (N_10321,N_9308,N_9436);
nor U10322 (N_10322,N_9644,N_9124);
xor U10323 (N_10323,N_9300,N_9649);
and U10324 (N_10324,N_9520,N_9548);
and U10325 (N_10325,N_9589,N_9835);
and U10326 (N_10326,N_9559,N_9678);
or U10327 (N_10327,N_9954,N_9912);
and U10328 (N_10328,N_9570,N_9171);
and U10329 (N_10329,N_9106,N_9638);
or U10330 (N_10330,N_9455,N_9539);
or U10331 (N_10331,N_9734,N_9130);
nand U10332 (N_10332,N_9639,N_9748);
and U10333 (N_10333,N_9872,N_9920);
nor U10334 (N_10334,N_9860,N_9048);
and U10335 (N_10335,N_9843,N_9526);
xnor U10336 (N_10336,N_9494,N_9326);
nand U10337 (N_10337,N_9797,N_9038);
nand U10338 (N_10338,N_9381,N_9957);
and U10339 (N_10339,N_9328,N_9287);
nor U10340 (N_10340,N_9122,N_9688);
xor U10341 (N_10341,N_9855,N_9676);
and U10342 (N_10342,N_9816,N_9606);
xnor U10343 (N_10343,N_9588,N_9299);
nor U10344 (N_10344,N_9732,N_9727);
and U10345 (N_10345,N_9479,N_9102);
or U10346 (N_10346,N_9905,N_9722);
nor U10347 (N_10347,N_9643,N_9362);
nor U10348 (N_10348,N_9944,N_9657);
or U10349 (N_10349,N_9553,N_9211);
nor U10350 (N_10350,N_9626,N_9157);
nand U10351 (N_10351,N_9441,N_9349);
nand U10352 (N_10352,N_9719,N_9540);
nor U10353 (N_10353,N_9897,N_9145);
and U10354 (N_10354,N_9294,N_9189);
xor U10355 (N_10355,N_9744,N_9173);
nor U10356 (N_10356,N_9336,N_9915);
and U10357 (N_10357,N_9991,N_9795);
or U10358 (N_10358,N_9375,N_9430);
nor U10359 (N_10359,N_9654,N_9004);
xor U10360 (N_10360,N_9190,N_9811);
or U10361 (N_10361,N_9036,N_9740);
nor U10362 (N_10362,N_9506,N_9664);
xor U10363 (N_10363,N_9032,N_9609);
and U10364 (N_10364,N_9891,N_9089);
nor U10365 (N_10365,N_9276,N_9176);
and U10366 (N_10366,N_9911,N_9866);
xnor U10367 (N_10367,N_9054,N_9582);
nand U10368 (N_10368,N_9619,N_9444);
or U10369 (N_10369,N_9760,N_9701);
nor U10370 (N_10370,N_9928,N_9717);
or U10371 (N_10371,N_9210,N_9823);
or U10372 (N_10372,N_9931,N_9460);
xor U10373 (N_10373,N_9024,N_9186);
and U10374 (N_10374,N_9995,N_9028);
or U10375 (N_10375,N_9450,N_9634);
nor U10376 (N_10376,N_9356,N_9393);
nor U10377 (N_10377,N_9833,N_9235);
xnor U10378 (N_10378,N_9561,N_9340);
or U10379 (N_10379,N_9836,N_9360);
and U10380 (N_10380,N_9687,N_9637);
or U10381 (N_10381,N_9976,N_9969);
xnor U10382 (N_10382,N_9330,N_9005);
and U10383 (N_10383,N_9063,N_9325);
nand U10384 (N_10384,N_9844,N_9473);
xor U10385 (N_10385,N_9647,N_9022);
nor U10386 (N_10386,N_9026,N_9044);
or U10387 (N_10387,N_9805,N_9599);
or U10388 (N_10388,N_9303,N_9002);
or U10389 (N_10389,N_9283,N_9834);
nand U10390 (N_10390,N_9318,N_9648);
nand U10391 (N_10391,N_9367,N_9518);
nor U10392 (N_10392,N_9222,N_9547);
xnor U10393 (N_10393,N_9576,N_9454);
and U10394 (N_10394,N_9601,N_9610);
or U10395 (N_10395,N_9877,N_9784);
or U10396 (N_10396,N_9166,N_9495);
and U10397 (N_10397,N_9693,N_9682);
nand U10398 (N_10398,N_9379,N_9629);
and U10399 (N_10399,N_9373,N_9412);
nand U10400 (N_10400,N_9162,N_9698);
nand U10401 (N_10401,N_9885,N_9259);
or U10402 (N_10402,N_9670,N_9129);
or U10403 (N_10403,N_9541,N_9988);
or U10404 (N_10404,N_9880,N_9087);
and U10405 (N_10405,N_9775,N_9275);
xnor U10406 (N_10406,N_9550,N_9291);
nand U10407 (N_10407,N_9758,N_9391);
nor U10408 (N_10408,N_9407,N_9001);
and U10409 (N_10409,N_9938,N_9747);
and U10410 (N_10410,N_9253,N_9697);
nor U10411 (N_10411,N_9829,N_9020);
nor U10412 (N_10412,N_9562,N_9867);
xor U10413 (N_10413,N_9343,N_9523);
xnor U10414 (N_10414,N_9271,N_9345);
nor U10415 (N_10415,N_9080,N_9497);
xor U10416 (N_10416,N_9854,N_9802);
nand U10417 (N_10417,N_9111,N_9695);
and U10418 (N_10418,N_9943,N_9852);
xnor U10419 (N_10419,N_9432,N_9590);
or U10420 (N_10420,N_9704,N_9900);
xor U10421 (N_10421,N_9208,N_9302);
nor U10422 (N_10422,N_9881,N_9477);
nand U10423 (N_10423,N_9814,N_9323);
and U10424 (N_10424,N_9404,N_9105);
or U10425 (N_10425,N_9645,N_9801);
and U10426 (N_10426,N_9793,N_9395);
xnor U10427 (N_10427,N_9992,N_9422);
nor U10428 (N_10428,N_9051,N_9480);
or U10429 (N_10429,N_9508,N_9475);
nand U10430 (N_10430,N_9960,N_9206);
and U10431 (N_10431,N_9500,N_9875);
and U10432 (N_10432,N_9018,N_9686);
nor U10433 (N_10433,N_9581,N_9567);
nor U10434 (N_10434,N_9150,N_9731);
or U10435 (N_10435,N_9012,N_9675);
xor U10436 (N_10436,N_9316,N_9304);
xor U10437 (N_10437,N_9260,N_9418);
or U10438 (N_10438,N_9096,N_9907);
nand U10439 (N_10439,N_9241,N_9163);
nor U10440 (N_10440,N_9413,N_9123);
nand U10441 (N_10441,N_9919,N_9705);
nor U10442 (N_10442,N_9138,N_9296);
nor U10443 (N_10443,N_9425,N_9394);
or U10444 (N_10444,N_9549,N_9231);
xor U10445 (N_10445,N_9827,N_9093);
xnor U10446 (N_10446,N_9605,N_9806);
or U10447 (N_10447,N_9250,N_9489);
or U10448 (N_10448,N_9868,N_9411);
nor U10449 (N_10449,N_9354,N_9193);
and U10450 (N_10450,N_9857,N_9143);
and U10451 (N_10451,N_9442,N_9756);
nand U10452 (N_10452,N_9847,N_9580);
nor U10453 (N_10453,N_9738,N_9925);
and U10454 (N_10454,N_9887,N_9149);
nand U10455 (N_10455,N_9448,N_9564);
nand U10456 (N_10456,N_9674,N_9714);
nor U10457 (N_10457,N_9993,N_9587);
xnor U10458 (N_10458,N_9929,N_9741);
nor U10459 (N_10459,N_9666,N_9613);
nand U10460 (N_10460,N_9390,N_9224);
nor U10461 (N_10461,N_9894,N_9248);
xor U10462 (N_10462,N_9733,N_9726);
nand U10463 (N_10463,N_9502,N_9317);
or U10464 (N_10464,N_9542,N_9214);
and U10465 (N_10465,N_9041,N_9903);
nor U10466 (N_10466,N_9892,N_9781);
or U10467 (N_10467,N_9463,N_9585);
nor U10468 (N_10468,N_9293,N_9513);
nand U10469 (N_10469,N_9003,N_9055);
and U10470 (N_10470,N_9918,N_9837);
nor U10471 (N_10471,N_9457,N_9641);
nor U10472 (N_10472,N_9209,N_9862);
nand U10473 (N_10473,N_9266,N_9261);
nand U10474 (N_10474,N_9447,N_9083);
nand U10475 (N_10475,N_9160,N_9501);
nand U10476 (N_10476,N_9936,N_9216);
and U10477 (N_10477,N_9708,N_9161);
nor U10478 (N_10478,N_9088,N_9566);
nor U10479 (N_10479,N_9710,N_9555);
xor U10480 (N_10480,N_9057,N_9757);
and U10481 (N_10481,N_9397,N_9337);
nand U10482 (N_10482,N_9333,N_9070);
nor U10483 (N_10483,N_9033,N_9767);
and U10484 (N_10484,N_9780,N_9428);
nor U10485 (N_10485,N_9893,N_9884);
nor U10486 (N_10486,N_9010,N_9154);
and U10487 (N_10487,N_9690,N_9768);
or U10488 (N_10488,N_9254,N_9046);
nor U10489 (N_10489,N_9076,N_9347);
or U10490 (N_10490,N_9134,N_9355);
and U10491 (N_10491,N_9359,N_9987);
nor U10492 (N_10492,N_9257,N_9673);
xnor U10493 (N_10493,N_9924,N_9607);
nand U10494 (N_10494,N_9819,N_9558);
and U10495 (N_10495,N_9902,N_9942);
nor U10496 (N_10496,N_9656,N_9468);
xnor U10497 (N_10497,N_9712,N_9064);
nor U10498 (N_10498,N_9503,N_9140);
nand U10499 (N_10499,N_9043,N_9279);
and U10500 (N_10500,N_9910,N_9355);
nor U10501 (N_10501,N_9642,N_9054);
or U10502 (N_10502,N_9185,N_9116);
xnor U10503 (N_10503,N_9722,N_9762);
nand U10504 (N_10504,N_9897,N_9068);
nor U10505 (N_10505,N_9206,N_9106);
nor U10506 (N_10506,N_9237,N_9134);
nor U10507 (N_10507,N_9542,N_9490);
nor U10508 (N_10508,N_9047,N_9695);
nor U10509 (N_10509,N_9049,N_9171);
and U10510 (N_10510,N_9926,N_9743);
or U10511 (N_10511,N_9093,N_9233);
nor U10512 (N_10512,N_9384,N_9689);
and U10513 (N_10513,N_9802,N_9545);
xor U10514 (N_10514,N_9602,N_9660);
nor U10515 (N_10515,N_9335,N_9482);
nor U10516 (N_10516,N_9400,N_9094);
and U10517 (N_10517,N_9067,N_9716);
nor U10518 (N_10518,N_9331,N_9280);
xnor U10519 (N_10519,N_9627,N_9286);
nor U10520 (N_10520,N_9370,N_9938);
nor U10521 (N_10521,N_9826,N_9049);
nor U10522 (N_10522,N_9365,N_9299);
or U10523 (N_10523,N_9249,N_9938);
nor U10524 (N_10524,N_9394,N_9766);
or U10525 (N_10525,N_9688,N_9079);
xor U10526 (N_10526,N_9681,N_9772);
xor U10527 (N_10527,N_9173,N_9561);
nor U10528 (N_10528,N_9313,N_9770);
or U10529 (N_10529,N_9449,N_9677);
nand U10530 (N_10530,N_9076,N_9825);
nor U10531 (N_10531,N_9826,N_9883);
or U10532 (N_10532,N_9708,N_9528);
nand U10533 (N_10533,N_9448,N_9815);
nand U10534 (N_10534,N_9662,N_9825);
and U10535 (N_10535,N_9819,N_9915);
xnor U10536 (N_10536,N_9006,N_9259);
nand U10537 (N_10537,N_9778,N_9754);
nor U10538 (N_10538,N_9106,N_9806);
and U10539 (N_10539,N_9675,N_9864);
xor U10540 (N_10540,N_9459,N_9580);
xnor U10541 (N_10541,N_9226,N_9724);
or U10542 (N_10542,N_9509,N_9918);
xor U10543 (N_10543,N_9574,N_9794);
xor U10544 (N_10544,N_9954,N_9123);
or U10545 (N_10545,N_9177,N_9856);
and U10546 (N_10546,N_9094,N_9092);
or U10547 (N_10547,N_9672,N_9133);
nor U10548 (N_10548,N_9187,N_9132);
nor U10549 (N_10549,N_9784,N_9373);
nor U10550 (N_10550,N_9834,N_9585);
and U10551 (N_10551,N_9067,N_9824);
or U10552 (N_10552,N_9672,N_9347);
and U10553 (N_10553,N_9587,N_9126);
and U10554 (N_10554,N_9328,N_9238);
xnor U10555 (N_10555,N_9875,N_9937);
xnor U10556 (N_10556,N_9515,N_9924);
nand U10557 (N_10557,N_9523,N_9411);
nor U10558 (N_10558,N_9574,N_9614);
nor U10559 (N_10559,N_9360,N_9813);
xor U10560 (N_10560,N_9141,N_9547);
and U10561 (N_10561,N_9350,N_9924);
or U10562 (N_10562,N_9234,N_9829);
xor U10563 (N_10563,N_9309,N_9562);
or U10564 (N_10564,N_9608,N_9135);
nand U10565 (N_10565,N_9755,N_9834);
or U10566 (N_10566,N_9553,N_9206);
nor U10567 (N_10567,N_9875,N_9245);
or U10568 (N_10568,N_9578,N_9723);
and U10569 (N_10569,N_9445,N_9365);
and U10570 (N_10570,N_9340,N_9476);
and U10571 (N_10571,N_9742,N_9840);
nor U10572 (N_10572,N_9072,N_9354);
nand U10573 (N_10573,N_9773,N_9647);
nor U10574 (N_10574,N_9998,N_9707);
xnor U10575 (N_10575,N_9353,N_9618);
and U10576 (N_10576,N_9209,N_9794);
nand U10577 (N_10577,N_9104,N_9191);
xor U10578 (N_10578,N_9579,N_9174);
or U10579 (N_10579,N_9610,N_9843);
xnor U10580 (N_10580,N_9592,N_9577);
nand U10581 (N_10581,N_9816,N_9070);
nor U10582 (N_10582,N_9376,N_9685);
nand U10583 (N_10583,N_9081,N_9910);
and U10584 (N_10584,N_9019,N_9388);
nand U10585 (N_10585,N_9244,N_9592);
nand U10586 (N_10586,N_9027,N_9210);
or U10587 (N_10587,N_9131,N_9379);
nand U10588 (N_10588,N_9096,N_9204);
and U10589 (N_10589,N_9306,N_9675);
nor U10590 (N_10590,N_9875,N_9735);
nor U10591 (N_10591,N_9373,N_9575);
nand U10592 (N_10592,N_9180,N_9322);
nor U10593 (N_10593,N_9459,N_9964);
nor U10594 (N_10594,N_9686,N_9066);
nand U10595 (N_10595,N_9892,N_9706);
and U10596 (N_10596,N_9003,N_9401);
xnor U10597 (N_10597,N_9109,N_9271);
xor U10598 (N_10598,N_9527,N_9097);
xnor U10599 (N_10599,N_9363,N_9150);
nand U10600 (N_10600,N_9431,N_9342);
and U10601 (N_10601,N_9812,N_9280);
xor U10602 (N_10602,N_9627,N_9111);
xor U10603 (N_10603,N_9610,N_9212);
xnor U10604 (N_10604,N_9735,N_9512);
and U10605 (N_10605,N_9342,N_9815);
and U10606 (N_10606,N_9470,N_9028);
and U10607 (N_10607,N_9493,N_9629);
nand U10608 (N_10608,N_9990,N_9060);
nor U10609 (N_10609,N_9839,N_9671);
nor U10610 (N_10610,N_9407,N_9315);
or U10611 (N_10611,N_9129,N_9032);
nor U10612 (N_10612,N_9523,N_9209);
or U10613 (N_10613,N_9666,N_9215);
or U10614 (N_10614,N_9148,N_9771);
and U10615 (N_10615,N_9419,N_9603);
nor U10616 (N_10616,N_9989,N_9135);
xor U10617 (N_10617,N_9480,N_9531);
and U10618 (N_10618,N_9754,N_9980);
xor U10619 (N_10619,N_9434,N_9156);
xnor U10620 (N_10620,N_9552,N_9488);
nand U10621 (N_10621,N_9871,N_9383);
nand U10622 (N_10622,N_9964,N_9612);
or U10623 (N_10623,N_9110,N_9718);
xnor U10624 (N_10624,N_9729,N_9116);
nand U10625 (N_10625,N_9651,N_9462);
or U10626 (N_10626,N_9417,N_9330);
nor U10627 (N_10627,N_9815,N_9583);
nand U10628 (N_10628,N_9834,N_9439);
xor U10629 (N_10629,N_9532,N_9976);
xnor U10630 (N_10630,N_9521,N_9608);
xor U10631 (N_10631,N_9563,N_9694);
or U10632 (N_10632,N_9633,N_9315);
and U10633 (N_10633,N_9364,N_9912);
nand U10634 (N_10634,N_9266,N_9940);
xnor U10635 (N_10635,N_9098,N_9348);
nor U10636 (N_10636,N_9268,N_9983);
nor U10637 (N_10637,N_9523,N_9661);
xor U10638 (N_10638,N_9429,N_9502);
and U10639 (N_10639,N_9917,N_9087);
and U10640 (N_10640,N_9761,N_9269);
xor U10641 (N_10641,N_9365,N_9056);
xor U10642 (N_10642,N_9245,N_9706);
nand U10643 (N_10643,N_9678,N_9565);
nand U10644 (N_10644,N_9303,N_9201);
nor U10645 (N_10645,N_9539,N_9278);
xnor U10646 (N_10646,N_9916,N_9863);
nand U10647 (N_10647,N_9964,N_9594);
nor U10648 (N_10648,N_9309,N_9134);
xor U10649 (N_10649,N_9485,N_9442);
nor U10650 (N_10650,N_9534,N_9565);
or U10651 (N_10651,N_9872,N_9560);
xor U10652 (N_10652,N_9658,N_9136);
or U10653 (N_10653,N_9529,N_9009);
and U10654 (N_10654,N_9197,N_9779);
or U10655 (N_10655,N_9532,N_9096);
and U10656 (N_10656,N_9741,N_9715);
nand U10657 (N_10657,N_9197,N_9028);
or U10658 (N_10658,N_9941,N_9389);
nor U10659 (N_10659,N_9531,N_9211);
or U10660 (N_10660,N_9831,N_9291);
or U10661 (N_10661,N_9115,N_9449);
nor U10662 (N_10662,N_9915,N_9281);
nor U10663 (N_10663,N_9649,N_9960);
xor U10664 (N_10664,N_9994,N_9975);
nand U10665 (N_10665,N_9473,N_9740);
xor U10666 (N_10666,N_9248,N_9179);
and U10667 (N_10667,N_9915,N_9376);
nand U10668 (N_10668,N_9527,N_9042);
and U10669 (N_10669,N_9622,N_9660);
or U10670 (N_10670,N_9065,N_9942);
xor U10671 (N_10671,N_9963,N_9431);
nor U10672 (N_10672,N_9194,N_9068);
xnor U10673 (N_10673,N_9889,N_9818);
nand U10674 (N_10674,N_9345,N_9988);
nand U10675 (N_10675,N_9663,N_9897);
xor U10676 (N_10676,N_9311,N_9315);
or U10677 (N_10677,N_9590,N_9389);
nand U10678 (N_10678,N_9404,N_9263);
xnor U10679 (N_10679,N_9252,N_9691);
xor U10680 (N_10680,N_9051,N_9528);
and U10681 (N_10681,N_9493,N_9657);
and U10682 (N_10682,N_9323,N_9171);
nor U10683 (N_10683,N_9013,N_9177);
xor U10684 (N_10684,N_9512,N_9344);
nand U10685 (N_10685,N_9447,N_9788);
nor U10686 (N_10686,N_9325,N_9724);
and U10687 (N_10687,N_9459,N_9549);
or U10688 (N_10688,N_9836,N_9229);
nor U10689 (N_10689,N_9813,N_9468);
nand U10690 (N_10690,N_9063,N_9567);
nor U10691 (N_10691,N_9529,N_9751);
nand U10692 (N_10692,N_9716,N_9652);
xnor U10693 (N_10693,N_9850,N_9781);
xor U10694 (N_10694,N_9614,N_9780);
nand U10695 (N_10695,N_9007,N_9705);
and U10696 (N_10696,N_9435,N_9149);
nor U10697 (N_10697,N_9139,N_9484);
xor U10698 (N_10698,N_9871,N_9690);
xnor U10699 (N_10699,N_9034,N_9750);
xor U10700 (N_10700,N_9334,N_9652);
nand U10701 (N_10701,N_9396,N_9945);
or U10702 (N_10702,N_9067,N_9492);
nor U10703 (N_10703,N_9923,N_9059);
or U10704 (N_10704,N_9665,N_9148);
nand U10705 (N_10705,N_9208,N_9995);
xnor U10706 (N_10706,N_9784,N_9386);
nor U10707 (N_10707,N_9855,N_9207);
and U10708 (N_10708,N_9910,N_9060);
and U10709 (N_10709,N_9157,N_9912);
or U10710 (N_10710,N_9553,N_9834);
nor U10711 (N_10711,N_9088,N_9482);
and U10712 (N_10712,N_9719,N_9265);
nor U10713 (N_10713,N_9072,N_9066);
and U10714 (N_10714,N_9455,N_9480);
and U10715 (N_10715,N_9033,N_9940);
nand U10716 (N_10716,N_9780,N_9896);
xnor U10717 (N_10717,N_9400,N_9709);
xor U10718 (N_10718,N_9786,N_9801);
nand U10719 (N_10719,N_9558,N_9561);
nand U10720 (N_10720,N_9904,N_9414);
nand U10721 (N_10721,N_9952,N_9561);
xnor U10722 (N_10722,N_9373,N_9250);
or U10723 (N_10723,N_9909,N_9877);
xor U10724 (N_10724,N_9301,N_9599);
nand U10725 (N_10725,N_9204,N_9213);
nand U10726 (N_10726,N_9502,N_9924);
nor U10727 (N_10727,N_9804,N_9692);
nand U10728 (N_10728,N_9317,N_9135);
or U10729 (N_10729,N_9494,N_9944);
nor U10730 (N_10730,N_9461,N_9199);
nand U10731 (N_10731,N_9017,N_9648);
nor U10732 (N_10732,N_9938,N_9243);
nand U10733 (N_10733,N_9287,N_9442);
xor U10734 (N_10734,N_9668,N_9031);
and U10735 (N_10735,N_9145,N_9618);
nand U10736 (N_10736,N_9641,N_9515);
nor U10737 (N_10737,N_9103,N_9949);
xor U10738 (N_10738,N_9494,N_9488);
and U10739 (N_10739,N_9466,N_9082);
nand U10740 (N_10740,N_9157,N_9274);
xnor U10741 (N_10741,N_9289,N_9738);
nand U10742 (N_10742,N_9861,N_9033);
nand U10743 (N_10743,N_9084,N_9905);
and U10744 (N_10744,N_9266,N_9570);
xor U10745 (N_10745,N_9412,N_9394);
xor U10746 (N_10746,N_9796,N_9776);
xor U10747 (N_10747,N_9024,N_9399);
and U10748 (N_10748,N_9589,N_9402);
nor U10749 (N_10749,N_9889,N_9834);
xor U10750 (N_10750,N_9159,N_9247);
or U10751 (N_10751,N_9549,N_9917);
or U10752 (N_10752,N_9387,N_9659);
nand U10753 (N_10753,N_9652,N_9821);
or U10754 (N_10754,N_9876,N_9998);
xnor U10755 (N_10755,N_9024,N_9195);
xor U10756 (N_10756,N_9194,N_9302);
or U10757 (N_10757,N_9462,N_9052);
or U10758 (N_10758,N_9380,N_9558);
xor U10759 (N_10759,N_9569,N_9967);
or U10760 (N_10760,N_9062,N_9579);
xor U10761 (N_10761,N_9860,N_9219);
and U10762 (N_10762,N_9833,N_9228);
and U10763 (N_10763,N_9855,N_9121);
xnor U10764 (N_10764,N_9555,N_9664);
and U10765 (N_10765,N_9743,N_9121);
xor U10766 (N_10766,N_9785,N_9513);
or U10767 (N_10767,N_9113,N_9561);
nand U10768 (N_10768,N_9344,N_9905);
nor U10769 (N_10769,N_9842,N_9871);
or U10770 (N_10770,N_9665,N_9513);
nand U10771 (N_10771,N_9403,N_9477);
xnor U10772 (N_10772,N_9305,N_9739);
xnor U10773 (N_10773,N_9961,N_9818);
or U10774 (N_10774,N_9492,N_9887);
nor U10775 (N_10775,N_9380,N_9008);
nor U10776 (N_10776,N_9796,N_9619);
and U10777 (N_10777,N_9240,N_9753);
nand U10778 (N_10778,N_9534,N_9485);
nor U10779 (N_10779,N_9102,N_9930);
xor U10780 (N_10780,N_9778,N_9766);
nor U10781 (N_10781,N_9165,N_9377);
nor U10782 (N_10782,N_9892,N_9412);
nor U10783 (N_10783,N_9000,N_9548);
nor U10784 (N_10784,N_9775,N_9140);
nand U10785 (N_10785,N_9697,N_9854);
or U10786 (N_10786,N_9843,N_9225);
xor U10787 (N_10787,N_9823,N_9198);
nand U10788 (N_10788,N_9874,N_9123);
or U10789 (N_10789,N_9376,N_9825);
nand U10790 (N_10790,N_9244,N_9231);
nand U10791 (N_10791,N_9169,N_9572);
nor U10792 (N_10792,N_9020,N_9768);
xnor U10793 (N_10793,N_9920,N_9955);
nand U10794 (N_10794,N_9797,N_9057);
or U10795 (N_10795,N_9994,N_9022);
nor U10796 (N_10796,N_9347,N_9739);
nor U10797 (N_10797,N_9189,N_9550);
and U10798 (N_10798,N_9839,N_9905);
or U10799 (N_10799,N_9728,N_9932);
or U10800 (N_10800,N_9365,N_9949);
and U10801 (N_10801,N_9053,N_9067);
nand U10802 (N_10802,N_9118,N_9932);
or U10803 (N_10803,N_9785,N_9211);
nand U10804 (N_10804,N_9862,N_9979);
nor U10805 (N_10805,N_9824,N_9366);
nor U10806 (N_10806,N_9952,N_9494);
and U10807 (N_10807,N_9269,N_9689);
nor U10808 (N_10808,N_9541,N_9677);
or U10809 (N_10809,N_9994,N_9435);
and U10810 (N_10810,N_9848,N_9670);
or U10811 (N_10811,N_9600,N_9404);
nor U10812 (N_10812,N_9015,N_9621);
or U10813 (N_10813,N_9879,N_9909);
and U10814 (N_10814,N_9061,N_9828);
xor U10815 (N_10815,N_9243,N_9853);
nor U10816 (N_10816,N_9602,N_9005);
nand U10817 (N_10817,N_9011,N_9184);
xnor U10818 (N_10818,N_9513,N_9672);
and U10819 (N_10819,N_9804,N_9685);
or U10820 (N_10820,N_9775,N_9800);
xnor U10821 (N_10821,N_9606,N_9175);
nor U10822 (N_10822,N_9659,N_9090);
nor U10823 (N_10823,N_9482,N_9340);
xor U10824 (N_10824,N_9324,N_9995);
or U10825 (N_10825,N_9516,N_9999);
nand U10826 (N_10826,N_9724,N_9197);
nand U10827 (N_10827,N_9014,N_9894);
nor U10828 (N_10828,N_9272,N_9697);
nor U10829 (N_10829,N_9845,N_9736);
nand U10830 (N_10830,N_9440,N_9147);
or U10831 (N_10831,N_9268,N_9835);
or U10832 (N_10832,N_9192,N_9554);
nor U10833 (N_10833,N_9292,N_9161);
nor U10834 (N_10834,N_9673,N_9492);
or U10835 (N_10835,N_9837,N_9375);
nor U10836 (N_10836,N_9125,N_9604);
or U10837 (N_10837,N_9968,N_9358);
xnor U10838 (N_10838,N_9410,N_9802);
nand U10839 (N_10839,N_9526,N_9629);
nor U10840 (N_10840,N_9982,N_9834);
or U10841 (N_10841,N_9425,N_9344);
and U10842 (N_10842,N_9581,N_9710);
or U10843 (N_10843,N_9042,N_9088);
and U10844 (N_10844,N_9593,N_9795);
or U10845 (N_10845,N_9794,N_9446);
nor U10846 (N_10846,N_9855,N_9903);
nor U10847 (N_10847,N_9127,N_9964);
nor U10848 (N_10848,N_9030,N_9808);
and U10849 (N_10849,N_9742,N_9601);
and U10850 (N_10850,N_9330,N_9568);
or U10851 (N_10851,N_9612,N_9415);
nand U10852 (N_10852,N_9353,N_9252);
nor U10853 (N_10853,N_9372,N_9475);
or U10854 (N_10854,N_9696,N_9979);
and U10855 (N_10855,N_9013,N_9207);
xnor U10856 (N_10856,N_9076,N_9338);
xnor U10857 (N_10857,N_9806,N_9126);
nand U10858 (N_10858,N_9695,N_9590);
or U10859 (N_10859,N_9239,N_9211);
nand U10860 (N_10860,N_9159,N_9927);
nand U10861 (N_10861,N_9962,N_9980);
nand U10862 (N_10862,N_9440,N_9086);
or U10863 (N_10863,N_9690,N_9006);
and U10864 (N_10864,N_9829,N_9093);
and U10865 (N_10865,N_9992,N_9867);
or U10866 (N_10866,N_9993,N_9973);
nand U10867 (N_10867,N_9283,N_9794);
nand U10868 (N_10868,N_9619,N_9789);
xor U10869 (N_10869,N_9723,N_9143);
or U10870 (N_10870,N_9302,N_9823);
nand U10871 (N_10871,N_9300,N_9797);
nor U10872 (N_10872,N_9984,N_9948);
xnor U10873 (N_10873,N_9013,N_9158);
or U10874 (N_10874,N_9244,N_9882);
and U10875 (N_10875,N_9927,N_9579);
xnor U10876 (N_10876,N_9113,N_9144);
or U10877 (N_10877,N_9069,N_9837);
and U10878 (N_10878,N_9629,N_9236);
xnor U10879 (N_10879,N_9615,N_9433);
or U10880 (N_10880,N_9428,N_9416);
or U10881 (N_10881,N_9580,N_9564);
nand U10882 (N_10882,N_9267,N_9722);
nand U10883 (N_10883,N_9277,N_9945);
nand U10884 (N_10884,N_9290,N_9324);
or U10885 (N_10885,N_9475,N_9160);
or U10886 (N_10886,N_9225,N_9146);
xor U10887 (N_10887,N_9575,N_9234);
nor U10888 (N_10888,N_9779,N_9025);
and U10889 (N_10889,N_9918,N_9752);
or U10890 (N_10890,N_9585,N_9622);
xnor U10891 (N_10891,N_9262,N_9345);
or U10892 (N_10892,N_9211,N_9402);
or U10893 (N_10893,N_9756,N_9859);
xnor U10894 (N_10894,N_9411,N_9034);
or U10895 (N_10895,N_9693,N_9376);
nor U10896 (N_10896,N_9195,N_9222);
nand U10897 (N_10897,N_9352,N_9303);
and U10898 (N_10898,N_9992,N_9406);
or U10899 (N_10899,N_9835,N_9361);
xor U10900 (N_10900,N_9301,N_9475);
and U10901 (N_10901,N_9033,N_9746);
and U10902 (N_10902,N_9845,N_9281);
nand U10903 (N_10903,N_9453,N_9421);
xnor U10904 (N_10904,N_9731,N_9904);
xnor U10905 (N_10905,N_9718,N_9820);
nor U10906 (N_10906,N_9379,N_9875);
nor U10907 (N_10907,N_9168,N_9416);
or U10908 (N_10908,N_9223,N_9827);
and U10909 (N_10909,N_9511,N_9116);
or U10910 (N_10910,N_9310,N_9656);
and U10911 (N_10911,N_9939,N_9292);
and U10912 (N_10912,N_9585,N_9547);
xnor U10913 (N_10913,N_9317,N_9260);
and U10914 (N_10914,N_9558,N_9756);
nand U10915 (N_10915,N_9665,N_9241);
nand U10916 (N_10916,N_9465,N_9984);
and U10917 (N_10917,N_9979,N_9799);
nand U10918 (N_10918,N_9571,N_9419);
and U10919 (N_10919,N_9839,N_9128);
or U10920 (N_10920,N_9713,N_9444);
or U10921 (N_10921,N_9054,N_9970);
xor U10922 (N_10922,N_9693,N_9388);
xnor U10923 (N_10923,N_9394,N_9966);
nor U10924 (N_10924,N_9427,N_9725);
xor U10925 (N_10925,N_9376,N_9871);
xor U10926 (N_10926,N_9573,N_9951);
or U10927 (N_10927,N_9189,N_9623);
nor U10928 (N_10928,N_9390,N_9675);
or U10929 (N_10929,N_9585,N_9774);
nand U10930 (N_10930,N_9457,N_9846);
and U10931 (N_10931,N_9177,N_9062);
nand U10932 (N_10932,N_9082,N_9293);
and U10933 (N_10933,N_9706,N_9344);
nand U10934 (N_10934,N_9161,N_9851);
nand U10935 (N_10935,N_9804,N_9067);
nor U10936 (N_10936,N_9974,N_9417);
xnor U10937 (N_10937,N_9931,N_9117);
nand U10938 (N_10938,N_9382,N_9315);
xnor U10939 (N_10939,N_9670,N_9800);
xor U10940 (N_10940,N_9553,N_9694);
xnor U10941 (N_10941,N_9133,N_9257);
and U10942 (N_10942,N_9648,N_9534);
xnor U10943 (N_10943,N_9427,N_9424);
xnor U10944 (N_10944,N_9934,N_9318);
xor U10945 (N_10945,N_9473,N_9568);
or U10946 (N_10946,N_9956,N_9975);
nand U10947 (N_10947,N_9157,N_9856);
nand U10948 (N_10948,N_9111,N_9200);
or U10949 (N_10949,N_9127,N_9397);
nand U10950 (N_10950,N_9531,N_9866);
or U10951 (N_10951,N_9999,N_9913);
or U10952 (N_10952,N_9923,N_9544);
xnor U10953 (N_10953,N_9918,N_9189);
nand U10954 (N_10954,N_9458,N_9315);
or U10955 (N_10955,N_9001,N_9045);
or U10956 (N_10956,N_9062,N_9961);
and U10957 (N_10957,N_9566,N_9355);
or U10958 (N_10958,N_9489,N_9961);
xnor U10959 (N_10959,N_9421,N_9674);
and U10960 (N_10960,N_9048,N_9143);
and U10961 (N_10961,N_9781,N_9108);
and U10962 (N_10962,N_9099,N_9754);
and U10963 (N_10963,N_9517,N_9596);
and U10964 (N_10964,N_9779,N_9173);
nand U10965 (N_10965,N_9971,N_9505);
and U10966 (N_10966,N_9756,N_9891);
or U10967 (N_10967,N_9548,N_9716);
nor U10968 (N_10968,N_9984,N_9257);
or U10969 (N_10969,N_9108,N_9179);
xnor U10970 (N_10970,N_9305,N_9403);
nor U10971 (N_10971,N_9623,N_9162);
nor U10972 (N_10972,N_9808,N_9579);
nand U10973 (N_10973,N_9566,N_9912);
nor U10974 (N_10974,N_9735,N_9481);
and U10975 (N_10975,N_9744,N_9028);
nand U10976 (N_10976,N_9071,N_9962);
or U10977 (N_10977,N_9646,N_9877);
or U10978 (N_10978,N_9242,N_9766);
nand U10979 (N_10979,N_9844,N_9028);
nand U10980 (N_10980,N_9125,N_9280);
nor U10981 (N_10981,N_9791,N_9531);
or U10982 (N_10982,N_9441,N_9034);
xnor U10983 (N_10983,N_9923,N_9938);
or U10984 (N_10984,N_9027,N_9674);
xnor U10985 (N_10985,N_9495,N_9687);
and U10986 (N_10986,N_9959,N_9626);
nor U10987 (N_10987,N_9180,N_9264);
and U10988 (N_10988,N_9653,N_9192);
nor U10989 (N_10989,N_9816,N_9669);
nor U10990 (N_10990,N_9755,N_9215);
xnor U10991 (N_10991,N_9680,N_9530);
nand U10992 (N_10992,N_9614,N_9298);
xor U10993 (N_10993,N_9067,N_9777);
or U10994 (N_10994,N_9007,N_9443);
xor U10995 (N_10995,N_9639,N_9558);
and U10996 (N_10996,N_9917,N_9028);
nor U10997 (N_10997,N_9470,N_9282);
and U10998 (N_10998,N_9908,N_9235);
and U10999 (N_10999,N_9410,N_9460);
and U11000 (N_11000,N_10546,N_10630);
nor U11001 (N_11001,N_10527,N_10440);
and U11002 (N_11002,N_10183,N_10532);
nor U11003 (N_11003,N_10087,N_10408);
or U11004 (N_11004,N_10148,N_10008);
and U11005 (N_11005,N_10357,N_10940);
nand U11006 (N_11006,N_10102,N_10572);
and U11007 (N_11007,N_10173,N_10376);
or U11008 (N_11008,N_10269,N_10647);
and U11009 (N_11009,N_10800,N_10064);
nor U11010 (N_11010,N_10762,N_10093);
xnor U11011 (N_11011,N_10319,N_10758);
and U11012 (N_11012,N_10878,N_10748);
nor U11013 (N_11013,N_10127,N_10742);
nor U11014 (N_11014,N_10254,N_10709);
or U11015 (N_11015,N_10722,N_10724);
or U11016 (N_11016,N_10455,N_10781);
nand U11017 (N_11017,N_10265,N_10063);
nand U11018 (N_11018,N_10207,N_10753);
nand U11019 (N_11019,N_10578,N_10231);
and U11020 (N_11020,N_10785,N_10418);
and U11021 (N_11021,N_10386,N_10216);
or U11022 (N_11022,N_10035,N_10863);
and U11023 (N_11023,N_10037,N_10689);
or U11024 (N_11024,N_10760,N_10658);
nor U11025 (N_11025,N_10350,N_10112);
nand U11026 (N_11026,N_10680,N_10777);
nor U11027 (N_11027,N_10374,N_10660);
and U11028 (N_11028,N_10019,N_10105);
nor U11029 (N_11029,N_10859,N_10109);
or U11030 (N_11030,N_10021,N_10471);
nand U11031 (N_11031,N_10784,N_10497);
xor U11032 (N_11032,N_10048,N_10429);
or U11033 (N_11033,N_10125,N_10246);
and U11034 (N_11034,N_10168,N_10931);
nand U11035 (N_11035,N_10707,N_10142);
xnor U11036 (N_11036,N_10293,N_10558);
nand U11037 (N_11037,N_10110,N_10239);
and U11038 (N_11038,N_10294,N_10977);
and U11039 (N_11039,N_10022,N_10211);
or U11040 (N_11040,N_10552,N_10477);
and U11041 (N_11041,N_10669,N_10364);
nor U11042 (N_11042,N_10494,N_10208);
and U11043 (N_11043,N_10426,N_10718);
nor U11044 (N_11044,N_10681,N_10803);
nor U11045 (N_11045,N_10519,N_10808);
xor U11046 (N_11046,N_10190,N_10244);
nand U11047 (N_11047,N_10002,N_10621);
nand U11048 (N_11048,N_10619,N_10156);
and U11049 (N_11049,N_10908,N_10320);
or U11050 (N_11050,N_10645,N_10197);
and U11051 (N_11051,N_10007,N_10754);
and U11052 (N_11052,N_10823,N_10170);
nand U11053 (N_11053,N_10475,N_10480);
nor U11054 (N_11054,N_10696,N_10000);
and U11055 (N_11055,N_10833,N_10038);
or U11056 (N_11056,N_10486,N_10143);
nor U11057 (N_11057,N_10034,N_10258);
and U11058 (N_11058,N_10797,N_10330);
and U11059 (N_11059,N_10469,N_10603);
xor U11060 (N_11060,N_10447,N_10739);
nor U11061 (N_11061,N_10529,N_10004);
and U11062 (N_11062,N_10686,N_10778);
or U11063 (N_11063,N_10407,N_10229);
or U11064 (N_11064,N_10904,N_10192);
nor U11065 (N_11065,N_10695,N_10262);
and U11066 (N_11066,N_10981,N_10865);
or U11067 (N_11067,N_10832,N_10139);
and U11068 (N_11068,N_10520,N_10980);
xor U11069 (N_11069,N_10721,N_10371);
nor U11070 (N_11070,N_10014,N_10523);
or U11071 (N_11071,N_10646,N_10678);
and U11072 (N_11072,N_10045,N_10544);
xnor U11073 (N_11073,N_10697,N_10082);
and U11074 (N_11074,N_10047,N_10194);
xnor U11075 (N_11075,N_10868,N_10614);
nor U11076 (N_11076,N_10581,N_10793);
nor U11077 (N_11077,N_10430,N_10242);
nor U11078 (N_11078,N_10343,N_10261);
nand U11079 (N_11079,N_10982,N_10484);
nand U11080 (N_11080,N_10006,N_10056);
and U11081 (N_11081,N_10372,N_10118);
xor U11082 (N_11082,N_10270,N_10310);
nand U11083 (N_11083,N_10297,N_10360);
and U11084 (N_11084,N_10074,N_10932);
or U11085 (N_11085,N_10478,N_10562);
or U11086 (N_11086,N_10235,N_10103);
nand U11087 (N_11087,N_10906,N_10772);
and U11088 (N_11088,N_10026,N_10749);
and U11089 (N_11089,N_10281,N_10234);
nor U11090 (N_11090,N_10589,N_10677);
or U11091 (N_11091,N_10271,N_10584);
and U11092 (N_11092,N_10327,N_10687);
and U11093 (N_11093,N_10060,N_10574);
nand U11094 (N_11094,N_10967,N_10538);
nor U11095 (N_11095,N_10570,N_10607);
nor U11096 (N_11096,N_10406,N_10180);
nor U11097 (N_11097,N_10363,N_10598);
and U11098 (N_11098,N_10691,N_10569);
or U11099 (N_11099,N_10915,N_10959);
and U11100 (N_11100,N_10155,N_10706);
and U11101 (N_11101,N_10567,N_10955);
and U11102 (N_11102,N_10298,N_10062);
xnor U11103 (N_11103,N_10555,N_10198);
and U11104 (N_11104,N_10186,N_10684);
and U11105 (N_11105,N_10759,N_10049);
and U11106 (N_11106,N_10286,N_10126);
xnor U11107 (N_11107,N_10410,N_10487);
and U11108 (N_11108,N_10276,N_10864);
xor U11109 (N_11109,N_10594,N_10307);
nor U11110 (N_11110,N_10903,N_10479);
nand U11111 (N_11111,N_10641,N_10086);
xor U11112 (N_11112,N_10446,N_10413);
or U11113 (N_11113,N_10543,N_10095);
nand U11114 (N_11114,N_10358,N_10934);
nand U11115 (N_11115,N_10354,N_10366);
nor U11116 (N_11116,N_10205,N_10916);
and U11117 (N_11117,N_10287,N_10771);
nand U11118 (N_11118,N_10869,N_10223);
nand U11119 (N_11119,N_10620,N_10811);
xor U11120 (N_11120,N_10114,N_10522);
and U11121 (N_11121,N_10027,N_10667);
nand U11122 (N_11122,N_10020,N_10462);
or U11123 (N_11123,N_10377,N_10801);
nor U11124 (N_11124,N_10767,N_10375);
nand U11125 (N_11125,N_10476,N_10987);
nand U11126 (N_11126,N_10174,N_10542);
nand U11127 (N_11127,N_10514,N_10381);
nor U11128 (N_11128,N_10836,N_10003);
xor U11129 (N_11129,N_10734,N_10819);
nand U11130 (N_11130,N_10837,N_10481);
or U11131 (N_11131,N_10861,N_10495);
nor U11132 (N_11132,N_10453,N_10136);
or U11133 (N_11133,N_10463,N_10666);
and U11134 (N_11134,N_10409,N_10752);
nor U11135 (N_11135,N_10124,N_10556);
nor U11136 (N_11136,N_10338,N_10184);
xnor U11137 (N_11137,N_10090,N_10018);
and U11138 (N_11138,N_10040,N_10296);
xor U11139 (N_11139,N_10444,N_10611);
or U11140 (N_11140,N_10962,N_10346);
and U11141 (N_11141,N_10396,N_10810);
nand U11142 (N_11142,N_10972,N_10617);
xnor U11143 (N_11143,N_10518,N_10873);
and U11144 (N_11144,N_10827,N_10703);
nor U11145 (N_11145,N_10061,N_10998);
xnor U11146 (N_11146,N_10640,N_10858);
or U11147 (N_11147,N_10547,N_10052);
or U11148 (N_11148,N_10822,N_10943);
xor U11149 (N_11149,N_10896,N_10111);
nand U11150 (N_11150,N_10768,N_10786);
nand U11151 (N_11151,N_10253,N_10181);
nor U11152 (N_11152,N_10512,N_10395);
nor U11153 (N_11153,N_10911,N_10421);
or U11154 (N_11154,N_10177,N_10147);
nand U11155 (N_11155,N_10348,N_10965);
nand U11156 (N_11156,N_10704,N_10694);
nand U11157 (N_11157,N_10502,N_10994);
nand U11158 (N_11158,N_10774,N_10732);
nor U11159 (N_11159,N_10989,N_10227);
or U11160 (N_11160,N_10491,N_10648);
nor U11161 (N_11161,N_10952,N_10563);
xnor U11162 (N_11162,N_10437,N_10220);
nand U11163 (N_11163,N_10834,N_10893);
nand U11164 (N_11164,N_10880,N_10013);
or U11165 (N_11165,N_10120,N_10728);
nor U11166 (N_11166,N_10466,N_10405);
nand U11167 (N_11167,N_10399,N_10098);
nor U11168 (N_11168,N_10411,N_10150);
or U11169 (N_11169,N_10830,N_10628);
xnor U11170 (N_11170,N_10971,N_10275);
and U11171 (N_11171,N_10291,N_10775);
nor U11172 (N_11172,N_10166,N_10218);
or U11173 (N_11173,N_10009,N_10137);
xor U11174 (N_11174,N_10664,N_10613);
or U11175 (N_11175,N_10263,N_10368);
nand U11176 (N_11176,N_10794,N_10665);
nand U11177 (N_11177,N_10266,N_10099);
xnor U11178 (N_11178,N_10847,N_10300);
or U11179 (N_11179,N_10590,N_10744);
nor U11180 (N_11180,N_10306,N_10394);
or U11181 (N_11181,N_10993,N_10160);
and U11182 (N_11182,N_10145,N_10738);
or U11183 (N_11183,N_10571,N_10152);
nand U11184 (N_11184,N_10969,N_10023);
xnor U11185 (N_11185,N_10698,N_10461);
nor U11186 (N_11186,N_10663,N_10369);
xor U11187 (N_11187,N_10860,N_10385);
nand U11188 (N_11188,N_10039,N_10073);
nor U11189 (N_11189,N_10610,N_10322);
nor U11190 (N_11190,N_10041,N_10597);
or U11191 (N_11191,N_10890,N_10163);
nand U11192 (N_11192,N_10313,N_10545);
nor U11193 (N_11193,N_10930,N_10116);
or U11194 (N_11194,N_10415,N_10164);
xor U11195 (N_11195,N_10092,N_10737);
xnor U11196 (N_11196,N_10923,N_10154);
and U11197 (N_11197,N_10089,N_10496);
and U11198 (N_11198,N_10755,N_10644);
and U11199 (N_11199,N_10131,N_10731);
nor U11200 (N_11200,N_10909,N_10433);
or U11201 (N_11201,N_10699,N_10146);
or U11202 (N_11202,N_10939,N_10919);
and U11203 (N_11203,N_10920,N_10158);
nor U11204 (N_11204,N_10248,N_10654);
xor U11205 (N_11205,N_10200,N_10420);
nand U11206 (N_11206,N_10895,N_10789);
xnor U11207 (N_11207,N_10540,N_10222);
or U11208 (N_11208,N_10028,N_10284);
nor U11209 (N_11209,N_10889,N_10730);
nor U11210 (N_11210,N_10165,N_10854);
xor U11211 (N_11211,N_10171,N_10252);
and U11212 (N_11212,N_10973,N_10872);
xnor U11213 (N_11213,N_10966,N_10991);
xnor U11214 (N_11214,N_10442,N_10072);
and U11215 (N_11215,N_10285,N_10070);
xnor U11216 (N_11216,N_10844,N_10113);
nand U11217 (N_11217,N_10465,N_10841);
and U11218 (N_11218,N_10199,N_10963);
nor U11219 (N_11219,N_10653,N_10945);
nand U11220 (N_11220,N_10257,N_10389);
and U11221 (N_11221,N_10575,N_10016);
or U11222 (N_11222,N_10970,N_10507);
xor U11223 (N_11223,N_10659,N_10601);
xnor U11224 (N_11224,N_10974,N_10138);
or U11225 (N_11225,N_10428,N_10676);
nor U11226 (N_11226,N_10928,N_10378);
and U11227 (N_11227,N_10080,N_10946);
or U11228 (N_11228,N_10325,N_10999);
xnor U11229 (N_11229,N_10172,N_10729);
nand U11230 (N_11230,N_10712,N_10956);
nor U11231 (N_11231,N_10012,N_10219);
nor U11232 (N_11232,N_10720,N_10826);
and U11233 (N_11233,N_10910,N_10331);
nor U11234 (N_11234,N_10950,N_10247);
and U11235 (N_11235,N_10788,N_10586);
nor U11236 (N_11236,N_10736,N_10879);
xor U11237 (N_11237,N_10067,N_10290);
nand U11238 (N_11238,N_10745,N_10609);
nand U11239 (N_11239,N_10141,N_10875);
xor U11240 (N_11240,N_10240,N_10936);
or U11241 (N_11241,N_10384,N_10651);
nand U11242 (N_11242,N_10935,N_10249);
nand U11243 (N_11243,N_10907,N_10526);
or U11244 (N_11244,N_10710,N_10984);
nor U11245 (N_11245,N_10344,N_10602);
xor U11246 (N_11246,N_10106,N_10929);
xor U11247 (N_11247,N_10783,N_10886);
nor U11248 (N_11248,N_10443,N_10553);
nor U11249 (N_11249,N_10353,N_10288);
nand U11250 (N_11250,N_10500,N_10005);
or U11251 (N_11251,N_10627,N_10191);
nor U11252 (N_11252,N_10888,N_10341);
or U11253 (N_11253,N_10452,N_10282);
or U11254 (N_11254,N_10159,N_10232);
nand U11255 (N_11255,N_10182,N_10355);
and U11256 (N_11256,N_10795,N_10516);
nor U11257 (N_11257,N_10299,N_10506);
nor U11258 (N_11258,N_10900,N_10809);
nand U11259 (N_11259,N_10947,N_10668);
nand U11260 (N_11260,N_10756,N_10457);
or U11261 (N_11261,N_10870,N_10882);
nand U11262 (N_11262,N_10831,N_10960);
xor U11263 (N_11263,N_10599,N_10390);
xor U11264 (N_11264,N_10485,N_10902);
or U11265 (N_11265,N_10046,N_10938);
nand U11266 (N_11266,N_10050,N_10937);
and U11267 (N_11267,N_10855,N_10990);
nand U11268 (N_11268,N_10770,N_10427);
and U11269 (N_11269,N_10577,N_10078);
or U11270 (N_11270,N_10001,N_10515);
xnor U11271 (N_11271,N_10814,N_10069);
nor U11272 (N_11272,N_10798,N_10874);
and U11273 (N_11273,N_10326,N_10656);
xnor U11274 (N_11274,N_10311,N_10820);
nor U11275 (N_11275,N_10539,N_10883);
and U11276 (N_11276,N_10986,N_10054);
and U11277 (N_11277,N_10448,N_10245);
xor U11278 (N_11278,N_10958,N_10107);
or U11279 (N_11279,N_10441,N_10856);
xnor U11280 (N_11280,N_10835,N_10345);
xor U11281 (N_11281,N_10370,N_10436);
or U11282 (N_11282,N_10314,N_10312);
nor U11283 (N_11283,N_10735,N_10482);
nand U11284 (N_11284,N_10334,N_10383);
and U11285 (N_11285,N_10979,N_10812);
or U11286 (N_11286,N_10193,N_10921);
nand U11287 (N_11287,N_10838,N_10179);
or U11288 (N_11288,N_10321,N_10011);
nor U11289 (N_11289,N_10238,N_10782);
and U11290 (N_11290,N_10806,N_10449);
nor U11291 (N_11291,N_10941,N_10277);
and U11292 (N_11292,N_10308,N_10488);
and U11293 (N_11293,N_10079,N_10670);
xor U11294 (N_11294,N_10504,N_10583);
or U11295 (N_11295,N_10853,N_10091);
and U11296 (N_11296,N_10228,N_10828);
nand U11297 (N_11297,N_10280,N_10100);
nor U11298 (N_11298,N_10392,N_10259);
nor U11299 (N_11299,N_10057,N_10029);
or U11300 (N_11300,N_10066,N_10176);
nor U11301 (N_11301,N_10985,N_10650);
or U11302 (N_11302,N_10790,N_10787);
nand U11303 (N_11303,N_10766,N_10434);
and U11304 (N_11304,N_10551,N_10918);
nand U11305 (N_11305,N_10978,N_10051);
nor U11306 (N_11306,N_10588,N_10241);
nor U11307 (N_11307,N_10685,N_10203);
nor U11308 (N_11308,N_10264,N_10279);
and U11309 (N_11309,N_10328,N_10690);
or U11310 (N_11310,N_10533,N_10295);
nand U11311 (N_11311,N_10212,N_10213);
nand U11312 (N_11312,N_10224,N_10133);
nand U11313 (N_11313,N_10451,N_10631);
nand U11314 (N_11314,N_10031,N_10818);
nand U11315 (N_11315,N_10115,N_10323);
nand U11316 (N_11316,N_10422,N_10596);
nand U11317 (N_11317,N_10397,N_10848);
and U11318 (N_11318,N_10424,N_10750);
or U11319 (N_11319,N_10568,N_10713);
nand U11320 (N_11320,N_10391,N_10877);
xnor U11321 (N_11321,N_10682,N_10492);
nand U11322 (N_11322,N_10530,N_10417);
or U11323 (N_11323,N_10195,N_10388);
nand U11324 (N_11324,N_10414,N_10632);
xnor U11325 (N_11325,N_10055,N_10303);
nor U11326 (N_11326,N_10779,N_10187);
nor U11327 (N_11327,N_10460,N_10683);
nor U11328 (N_11328,N_10084,N_10846);
nand U11329 (N_11329,N_10196,N_10802);
or U11330 (N_11330,N_10153,N_10849);
and U11331 (N_11331,N_10128,N_10508);
nor U11332 (N_11332,N_10302,N_10740);
nand U11333 (N_11333,N_10983,N_10309);
nand U11334 (N_11334,N_10315,N_10272);
nor U11335 (N_11335,N_10605,N_10202);
nor U11336 (N_11336,N_10033,N_10764);
xnor U11337 (N_11337,N_10175,N_10693);
nand U11338 (N_11338,N_10995,N_10509);
and U11339 (N_11339,N_10705,N_10379);
xor U11340 (N_11340,N_10083,N_10917);
xor U11341 (N_11341,N_10135,N_10214);
xor U11342 (N_11342,N_10361,N_10733);
or U11343 (N_11343,N_10821,N_10881);
nand U11344 (N_11344,N_10840,N_10565);
and U11345 (N_11345,N_10534,N_10121);
nand U11346 (N_11346,N_10304,N_10301);
nor U11347 (N_11347,N_10839,N_10557);
nand U11348 (N_11348,N_10123,N_10468);
or U11349 (N_11349,N_10961,N_10560);
nor U11350 (N_11350,N_10926,N_10373);
nand U11351 (N_11351,N_10473,N_10209);
nor U11352 (N_11352,N_10824,N_10010);
or U11353 (N_11353,N_10576,N_10897);
nor U11354 (N_11354,N_10503,N_10329);
or U11355 (N_11355,N_10517,N_10513);
and U11356 (N_11356,N_10942,N_10432);
and U11357 (N_11357,N_10852,N_10108);
xor U11358 (N_11358,N_10615,N_10679);
nand U11359 (N_11359,N_10119,N_10167);
nand U11360 (N_11360,N_10042,N_10474);
and U11361 (N_11361,N_10925,N_10425);
or U11362 (N_11362,N_10891,N_10600);
or U11363 (N_11363,N_10727,N_10278);
xnor U11364 (N_11364,N_10161,N_10592);
nor U11365 (N_11365,N_10566,N_10226);
nand U11366 (N_11366,N_10065,N_10580);
and U11367 (N_11367,N_10243,N_10843);
xor U11368 (N_11368,N_10525,N_10454);
and U11369 (N_11369,N_10548,N_10573);
nand U11370 (N_11370,N_10825,N_10256);
nor U11371 (N_11371,N_10725,N_10914);
xnor U11372 (N_11372,N_10899,N_10470);
xor U11373 (N_11373,N_10867,N_10857);
nand U11374 (N_11374,N_10711,N_10715);
nand U11375 (N_11375,N_10719,N_10901);
nor U11376 (N_11376,N_10922,N_10892);
nor U11377 (N_11377,N_10401,N_10804);
or U11378 (N_11378,N_10130,N_10185);
nor U11379 (N_11379,N_10816,N_10524);
or U11380 (N_11380,N_10639,N_10701);
nor U11381 (N_11381,N_10964,N_10351);
xor U11382 (N_11382,N_10535,N_10564);
and U11383 (N_11383,N_10431,N_10493);
and U11384 (N_11384,N_10400,N_10210);
nor U11385 (N_11385,N_10842,N_10799);
and U11386 (N_11386,N_10655,N_10624);
and U11387 (N_11387,N_10324,N_10393);
xor U11388 (N_11388,N_10273,N_10129);
and U11389 (N_11389,N_10692,N_10521);
xor U11390 (N_11390,N_10550,N_10606);
and U11391 (N_11391,N_10635,N_10318);
nand U11392 (N_11392,N_10189,N_10283);
xor U11393 (N_11393,N_10403,N_10537);
xor U11394 (N_11394,N_10075,N_10541);
xnor U11395 (N_11395,N_10757,N_10629);
xor U11396 (N_11396,N_10250,N_10913);
and U11397 (N_11397,N_10531,N_10674);
nand U11398 (N_11398,N_10887,N_10933);
or U11399 (N_11399,N_10673,N_10894);
xnor U11400 (N_11400,N_10510,N_10289);
nand U11401 (N_11401,N_10702,N_10489);
or U11402 (N_11402,N_10215,N_10104);
or U11403 (N_11403,N_10595,N_10671);
nor U11404 (N_11404,N_10268,N_10992);
and U11405 (N_11405,N_10657,N_10043);
nor U11406 (N_11406,N_10976,N_10149);
nor U11407 (N_11407,N_10499,N_10636);
and U11408 (N_11408,N_10968,N_10763);
and U11409 (N_11409,N_10490,N_10380);
xnor U11410 (N_11410,N_10813,N_10032);
or U11411 (N_11411,N_10815,N_10700);
nand U11412 (N_11412,N_10618,N_10483);
xnor U11413 (N_11413,N_10081,N_10132);
nand U11414 (N_11414,N_10367,N_10412);
or U11415 (N_11415,N_10817,N_10217);
nor U11416 (N_11416,N_10162,N_10044);
xor U11417 (N_11417,N_10642,N_10387);
xor U11418 (N_11418,N_10807,N_10498);
xnor U11419 (N_11419,N_10255,N_10140);
xor U11420 (N_11420,N_10957,N_10423);
or U11421 (N_11421,N_10608,N_10638);
and U11422 (N_11422,N_10714,N_10340);
nand U11423 (N_11423,N_10204,N_10450);
and U11424 (N_11424,N_10459,N_10688);
xor U11425 (N_11425,N_10761,N_10267);
xnor U11426 (N_11426,N_10776,N_10251);
xnor U11427 (N_11427,N_10015,N_10662);
or U11428 (N_11428,N_10675,N_10912);
xnor U11429 (N_11429,N_10169,N_10097);
nand U11430 (N_11430,N_10356,N_10456);
nor U11431 (N_11431,N_10206,N_10382);
and U11432 (N_11432,N_10747,N_10404);
nor U11433 (N_11433,N_10997,N_10122);
nor U11434 (N_11434,N_10743,N_10746);
and U11435 (N_11435,N_10464,N_10030);
and U11436 (N_11436,N_10780,N_10511);
and U11437 (N_11437,N_10773,N_10419);
and U11438 (N_11438,N_10845,N_10332);
xor U11439 (N_11439,N_10643,N_10723);
nand U11440 (N_11440,N_10117,N_10649);
and U11441 (N_11441,N_10949,N_10094);
or U11442 (N_11442,N_10866,N_10333);
or U11443 (N_11443,N_10472,N_10096);
xnor U11444 (N_11444,N_10579,N_10829);
and U11445 (N_11445,N_10017,N_10365);
nand U11446 (N_11446,N_10591,N_10604);
xor U11447 (N_11447,N_10292,N_10274);
and U11448 (N_11448,N_10445,N_10726);
nand U11449 (N_11449,N_10549,N_10536);
nor U11450 (N_11450,N_10233,N_10077);
or U11451 (N_11451,N_10230,N_10988);
and U11452 (N_11452,N_10622,N_10975);
xor U11453 (N_11453,N_10501,N_10805);
nand U11454 (N_11454,N_10157,N_10717);
and U11455 (N_11455,N_10791,N_10237);
xnor U11456 (N_11456,N_10898,N_10347);
and U11457 (N_11457,N_10672,N_10036);
xnor U11458 (N_11458,N_10201,N_10612);
nor U11459 (N_11459,N_10221,N_10948);
nor U11460 (N_11460,N_10024,N_10633);
nand U11461 (N_11461,N_10559,N_10339);
nand U11462 (N_11462,N_10769,N_10349);
xor U11463 (N_11463,N_10335,N_10587);
nand U11464 (N_11464,N_10708,N_10336);
xor U11465 (N_11465,N_10071,N_10151);
and U11466 (N_11466,N_10352,N_10661);
nor U11467 (N_11467,N_10884,N_10582);
and U11468 (N_11468,N_10585,N_10085);
or U11469 (N_11469,N_10885,N_10402);
or U11470 (N_11470,N_10134,N_10236);
nor U11471 (N_11471,N_10944,N_10076);
nor U11472 (N_11472,N_10439,N_10554);
and U11473 (N_11473,N_10741,N_10059);
nand U11474 (N_11474,N_10305,N_10751);
xor U11475 (N_11475,N_10458,N_10188);
xnor U11476 (N_11476,N_10058,N_10623);
nor U11477 (N_11477,N_10053,N_10561);
and U11478 (N_11478,N_10593,N_10862);
or U11479 (N_11479,N_10616,N_10144);
xor U11480 (N_11480,N_10362,N_10951);
xnor U11481 (N_11481,N_10416,N_10876);
nor U11482 (N_11482,N_10652,N_10342);
or U11483 (N_11483,N_10317,N_10260);
and U11484 (N_11484,N_10626,N_10438);
xor U11485 (N_11485,N_10954,N_10337);
nand U11486 (N_11486,N_10505,N_10634);
nand U11487 (N_11487,N_10953,N_10716);
xnor U11488 (N_11488,N_10927,N_10905);
and U11489 (N_11489,N_10088,N_10178);
nand U11490 (N_11490,N_10467,N_10101);
or U11491 (N_11491,N_10765,N_10316);
nor U11492 (N_11492,N_10637,N_10850);
xnor U11493 (N_11493,N_10025,N_10796);
nor U11494 (N_11494,N_10359,N_10068);
and U11495 (N_11495,N_10924,N_10528);
or U11496 (N_11496,N_10225,N_10625);
and U11497 (N_11497,N_10435,N_10792);
xnor U11498 (N_11498,N_10851,N_10398);
nor U11499 (N_11499,N_10996,N_10871);
nor U11500 (N_11500,N_10129,N_10128);
nand U11501 (N_11501,N_10283,N_10461);
nor U11502 (N_11502,N_10750,N_10310);
and U11503 (N_11503,N_10499,N_10965);
and U11504 (N_11504,N_10228,N_10764);
xor U11505 (N_11505,N_10223,N_10097);
nand U11506 (N_11506,N_10053,N_10635);
and U11507 (N_11507,N_10914,N_10447);
or U11508 (N_11508,N_10797,N_10229);
nor U11509 (N_11509,N_10797,N_10199);
xor U11510 (N_11510,N_10750,N_10537);
or U11511 (N_11511,N_10794,N_10394);
and U11512 (N_11512,N_10643,N_10596);
and U11513 (N_11513,N_10327,N_10623);
xor U11514 (N_11514,N_10741,N_10000);
nand U11515 (N_11515,N_10676,N_10082);
and U11516 (N_11516,N_10817,N_10096);
nand U11517 (N_11517,N_10017,N_10057);
xor U11518 (N_11518,N_10156,N_10222);
xnor U11519 (N_11519,N_10689,N_10179);
and U11520 (N_11520,N_10669,N_10459);
and U11521 (N_11521,N_10584,N_10635);
nor U11522 (N_11522,N_10359,N_10854);
and U11523 (N_11523,N_10210,N_10410);
xor U11524 (N_11524,N_10973,N_10057);
or U11525 (N_11525,N_10816,N_10696);
nand U11526 (N_11526,N_10217,N_10635);
xnor U11527 (N_11527,N_10944,N_10708);
nor U11528 (N_11528,N_10008,N_10279);
or U11529 (N_11529,N_10003,N_10900);
or U11530 (N_11530,N_10913,N_10561);
nor U11531 (N_11531,N_10377,N_10232);
and U11532 (N_11532,N_10998,N_10040);
xor U11533 (N_11533,N_10445,N_10703);
and U11534 (N_11534,N_10434,N_10850);
nor U11535 (N_11535,N_10046,N_10179);
or U11536 (N_11536,N_10666,N_10187);
and U11537 (N_11537,N_10082,N_10635);
xor U11538 (N_11538,N_10319,N_10223);
and U11539 (N_11539,N_10350,N_10900);
and U11540 (N_11540,N_10362,N_10546);
nand U11541 (N_11541,N_10927,N_10249);
and U11542 (N_11542,N_10205,N_10668);
xnor U11543 (N_11543,N_10633,N_10723);
nand U11544 (N_11544,N_10689,N_10367);
xor U11545 (N_11545,N_10847,N_10145);
xnor U11546 (N_11546,N_10823,N_10286);
nor U11547 (N_11547,N_10102,N_10473);
xnor U11548 (N_11548,N_10705,N_10073);
or U11549 (N_11549,N_10823,N_10429);
nand U11550 (N_11550,N_10511,N_10624);
or U11551 (N_11551,N_10880,N_10206);
and U11552 (N_11552,N_10634,N_10439);
xor U11553 (N_11553,N_10152,N_10060);
nor U11554 (N_11554,N_10141,N_10914);
xnor U11555 (N_11555,N_10471,N_10337);
xnor U11556 (N_11556,N_10219,N_10211);
nand U11557 (N_11557,N_10656,N_10338);
nor U11558 (N_11558,N_10573,N_10770);
nor U11559 (N_11559,N_10580,N_10771);
or U11560 (N_11560,N_10736,N_10214);
or U11561 (N_11561,N_10351,N_10276);
nand U11562 (N_11562,N_10717,N_10557);
and U11563 (N_11563,N_10957,N_10686);
or U11564 (N_11564,N_10547,N_10537);
nand U11565 (N_11565,N_10901,N_10262);
nand U11566 (N_11566,N_10286,N_10647);
xor U11567 (N_11567,N_10422,N_10662);
xnor U11568 (N_11568,N_10989,N_10328);
or U11569 (N_11569,N_10008,N_10367);
nand U11570 (N_11570,N_10650,N_10886);
nand U11571 (N_11571,N_10850,N_10543);
nand U11572 (N_11572,N_10446,N_10206);
or U11573 (N_11573,N_10945,N_10968);
nor U11574 (N_11574,N_10219,N_10510);
nor U11575 (N_11575,N_10085,N_10044);
nor U11576 (N_11576,N_10273,N_10222);
xnor U11577 (N_11577,N_10988,N_10555);
and U11578 (N_11578,N_10641,N_10249);
and U11579 (N_11579,N_10548,N_10520);
xnor U11580 (N_11580,N_10714,N_10037);
xnor U11581 (N_11581,N_10039,N_10840);
nand U11582 (N_11582,N_10475,N_10964);
or U11583 (N_11583,N_10391,N_10061);
xnor U11584 (N_11584,N_10235,N_10515);
or U11585 (N_11585,N_10360,N_10952);
and U11586 (N_11586,N_10446,N_10545);
xnor U11587 (N_11587,N_10893,N_10021);
and U11588 (N_11588,N_10449,N_10451);
nand U11589 (N_11589,N_10639,N_10736);
nand U11590 (N_11590,N_10310,N_10977);
and U11591 (N_11591,N_10926,N_10108);
or U11592 (N_11592,N_10559,N_10418);
and U11593 (N_11593,N_10480,N_10744);
and U11594 (N_11594,N_10814,N_10774);
nor U11595 (N_11595,N_10299,N_10532);
nor U11596 (N_11596,N_10210,N_10795);
nand U11597 (N_11597,N_10133,N_10373);
or U11598 (N_11598,N_10293,N_10441);
nor U11599 (N_11599,N_10440,N_10861);
and U11600 (N_11600,N_10611,N_10389);
nand U11601 (N_11601,N_10535,N_10787);
or U11602 (N_11602,N_10725,N_10422);
nor U11603 (N_11603,N_10361,N_10866);
nand U11604 (N_11604,N_10472,N_10355);
nand U11605 (N_11605,N_10882,N_10199);
or U11606 (N_11606,N_10442,N_10249);
xor U11607 (N_11607,N_10948,N_10285);
xor U11608 (N_11608,N_10292,N_10220);
and U11609 (N_11609,N_10081,N_10950);
or U11610 (N_11610,N_10626,N_10200);
nand U11611 (N_11611,N_10379,N_10006);
and U11612 (N_11612,N_10808,N_10489);
or U11613 (N_11613,N_10113,N_10621);
nand U11614 (N_11614,N_10534,N_10991);
nand U11615 (N_11615,N_10292,N_10656);
xnor U11616 (N_11616,N_10273,N_10520);
and U11617 (N_11617,N_10059,N_10413);
nand U11618 (N_11618,N_10842,N_10816);
xnor U11619 (N_11619,N_10907,N_10758);
nand U11620 (N_11620,N_10536,N_10514);
nor U11621 (N_11621,N_10941,N_10822);
nor U11622 (N_11622,N_10036,N_10634);
or U11623 (N_11623,N_10880,N_10814);
nor U11624 (N_11624,N_10923,N_10725);
or U11625 (N_11625,N_10286,N_10644);
xnor U11626 (N_11626,N_10780,N_10031);
or U11627 (N_11627,N_10076,N_10634);
or U11628 (N_11628,N_10136,N_10860);
or U11629 (N_11629,N_10717,N_10758);
or U11630 (N_11630,N_10355,N_10696);
xor U11631 (N_11631,N_10686,N_10361);
or U11632 (N_11632,N_10465,N_10364);
and U11633 (N_11633,N_10482,N_10117);
nand U11634 (N_11634,N_10759,N_10289);
nor U11635 (N_11635,N_10338,N_10414);
or U11636 (N_11636,N_10803,N_10410);
and U11637 (N_11637,N_10559,N_10766);
nor U11638 (N_11638,N_10042,N_10265);
and U11639 (N_11639,N_10719,N_10986);
nor U11640 (N_11640,N_10091,N_10972);
xor U11641 (N_11641,N_10146,N_10923);
and U11642 (N_11642,N_10410,N_10000);
xnor U11643 (N_11643,N_10604,N_10371);
and U11644 (N_11644,N_10566,N_10329);
xor U11645 (N_11645,N_10058,N_10852);
and U11646 (N_11646,N_10355,N_10561);
nor U11647 (N_11647,N_10460,N_10092);
xor U11648 (N_11648,N_10217,N_10568);
xnor U11649 (N_11649,N_10777,N_10485);
nand U11650 (N_11650,N_10349,N_10197);
and U11651 (N_11651,N_10251,N_10894);
or U11652 (N_11652,N_10131,N_10116);
nor U11653 (N_11653,N_10483,N_10480);
or U11654 (N_11654,N_10464,N_10279);
nand U11655 (N_11655,N_10017,N_10414);
and U11656 (N_11656,N_10424,N_10641);
xnor U11657 (N_11657,N_10944,N_10488);
xnor U11658 (N_11658,N_10870,N_10608);
xnor U11659 (N_11659,N_10004,N_10971);
nor U11660 (N_11660,N_10141,N_10608);
nor U11661 (N_11661,N_10549,N_10986);
nand U11662 (N_11662,N_10303,N_10083);
and U11663 (N_11663,N_10433,N_10100);
nand U11664 (N_11664,N_10276,N_10615);
nand U11665 (N_11665,N_10573,N_10641);
nor U11666 (N_11666,N_10266,N_10361);
nor U11667 (N_11667,N_10500,N_10143);
nor U11668 (N_11668,N_10727,N_10044);
nand U11669 (N_11669,N_10223,N_10689);
nor U11670 (N_11670,N_10573,N_10206);
xor U11671 (N_11671,N_10795,N_10480);
nor U11672 (N_11672,N_10536,N_10709);
and U11673 (N_11673,N_10056,N_10410);
and U11674 (N_11674,N_10033,N_10628);
or U11675 (N_11675,N_10037,N_10976);
xor U11676 (N_11676,N_10385,N_10822);
xnor U11677 (N_11677,N_10880,N_10762);
xnor U11678 (N_11678,N_10913,N_10124);
or U11679 (N_11679,N_10212,N_10484);
or U11680 (N_11680,N_10166,N_10408);
nor U11681 (N_11681,N_10088,N_10118);
and U11682 (N_11682,N_10090,N_10066);
and U11683 (N_11683,N_10273,N_10371);
or U11684 (N_11684,N_10136,N_10661);
or U11685 (N_11685,N_10841,N_10352);
xor U11686 (N_11686,N_10808,N_10713);
xor U11687 (N_11687,N_10639,N_10466);
nand U11688 (N_11688,N_10400,N_10449);
xor U11689 (N_11689,N_10304,N_10924);
xor U11690 (N_11690,N_10302,N_10164);
and U11691 (N_11691,N_10547,N_10092);
xnor U11692 (N_11692,N_10850,N_10577);
and U11693 (N_11693,N_10767,N_10662);
xnor U11694 (N_11694,N_10707,N_10754);
nand U11695 (N_11695,N_10609,N_10446);
or U11696 (N_11696,N_10677,N_10043);
nor U11697 (N_11697,N_10673,N_10724);
or U11698 (N_11698,N_10610,N_10851);
and U11699 (N_11699,N_10645,N_10163);
and U11700 (N_11700,N_10412,N_10365);
or U11701 (N_11701,N_10905,N_10152);
nand U11702 (N_11702,N_10258,N_10080);
or U11703 (N_11703,N_10708,N_10656);
or U11704 (N_11704,N_10256,N_10659);
xnor U11705 (N_11705,N_10351,N_10098);
nand U11706 (N_11706,N_10868,N_10773);
nand U11707 (N_11707,N_10234,N_10245);
and U11708 (N_11708,N_10924,N_10463);
nand U11709 (N_11709,N_10747,N_10649);
nor U11710 (N_11710,N_10765,N_10999);
nand U11711 (N_11711,N_10474,N_10190);
xnor U11712 (N_11712,N_10529,N_10581);
nor U11713 (N_11713,N_10762,N_10278);
nor U11714 (N_11714,N_10419,N_10499);
xor U11715 (N_11715,N_10595,N_10197);
nand U11716 (N_11716,N_10721,N_10870);
nand U11717 (N_11717,N_10394,N_10606);
or U11718 (N_11718,N_10001,N_10525);
nor U11719 (N_11719,N_10133,N_10716);
nand U11720 (N_11720,N_10835,N_10222);
xnor U11721 (N_11721,N_10474,N_10398);
or U11722 (N_11722,N_10194,N_10821);
and U11723 (N_11723,N_10274,N_10269);
nor U11724 (N_11724,N_10351,N_10567);
nor U11725 (N_11725,N_10002,N_10876);
xnor U11726 (N_11726,N_10710,N_10698);
nand U11727 (N_11727,N_10753,N_10038);
nand U11728 (N_11728,N_10152,N_10118);
and U11729 (N_11729,N_10148,N_10874);
and U11730 (N_11730,N_10570,N_10155);
or U11731 (N_11731,N_10349,N_10965);
xor U11732 (N_11732,N_10852,N_10213);
xor U11733 (N_11733,N_10638,N_10094);
xor U11734 (N_11734,N_10085,N_10328);
or U11735 (N_11735,N_10692,N_10311);
or U11736 (N_11736,N_10577,N_10036);
nand U11737 (N_11737,N_10342,N_10425);
and U11738 (N_11738,N_10521,N_10091);
nor U11739 (N_11739,N_10835,N_10831);
and U11740 (N_11740,N_10921,N_10792);
nor U11741 (N_11741,N_10166,N_10806);
and U11742 (N_11742,N_10808,N_10000);
or U11743 (N_11743,N_10561,N_10341);
and U11744 (N_11744,N_10049,N_10668);
nand U11745 (N_11745,N_10435,N_10104);
and U11746 (N_11746,N_10760,N_10357);
nand U11747 (N_11747,N_10927,N_10003);
nand U11748 (N_11748,N_10726,N_10084);
nand U11749 (N_11749,N_10038,N_10214);
xnor U11750 (N_11750,N_10041,N_10044);
xnor U11751 (N_11751,N_10476,N_10861);
and U11752 (N_11752,N_10439,N_10234);
or U11753 (N_11753,N_10364,N_10675);
xor U11754 (N_11754,N_10865,N_10672);
xnor U11755 (N_11755,N_10156,N_10094);
nor U11756 (N_11756,N_10788,N_10622);
nor U11757 (N_11757,N_10522,N_10022);
and U11758 (N_11758,N_10019,N_10814);
xor U11759 (N_11759,N_10108,N_10096);
nor U11760 (N_11760,N_10076,N_10936);
nor U11761 (N_11761,N_10044,N_10999);
xor U11762 (N_11762,N_10770,N_10060);
or U11763 (N_11763,N_10258,N_10284);
nor U11764 (N_11764,N_10631,N_10552);
nand U11765 (N_11765,N_10177,N_10297);
and U11766 (N_11766,N_10409,N_10203);
nor U11767 (N_11767,N_10777,N_10759);
nand U11768 (N_11768,N_10503,N_10584);
and U11769 (N_11769,N_10384,N_10891);
nand U11770 (N_11770,N_10527,N_10351);
xnor U11771 (N_11771,N_10038,N_10163);
xnor U11772 (N_11772,N_10127,N_10209);
or U11773 (N_11773,N_10885,N_10931);
nor U11774 (N_11774,N_10558,N_10656);
nand U11775 (N_11775,N_10983,N_10951);
nand U11776 (N_11776,N_10070,N_10249);
nand U11777 (N_11777,N_10666,N_10098);
xnor U11778 (N_11778,N_10340,N_10000);
nor U11779 (N_11779,N_10936,N_10978);
nand U11780 (N_11780,N_10286,N_10391);
xor U11781 (N_11781,N_10093,N_10824);
nor U11782 (N_11782,N_10280,N_10881);
nor U11783 (N_11783,N_10063,N_10020);
and U11784 (N_11784,N_10921,N_10423);
and U11785 (N_11785,N_10901,N_10356);
xnor U11786 (N_11786,N_10148,N_10654);
or U11787 (N_11787,N_10598,N_10041);
nand U11788 (N_11788,N_10824,N_10912);
nor U11789 (N_11789,N_10034,N_10285);
nand U11790 (N_11790,N_10230,N_10052);
or U11791 (N_11791,N_10148,N_10306);
nor U11792 (N_11792,N_10204,N_10273);
xor U11793 (N_11793,N_10827,N_10194);
or U11794 (N_11794,N_10937,N_10251);
xnor U11795 (N_11795,N_10339,N_10413);
and U11796 (N_11796,N_10028,N_10903);
xnor U11797 (N_11797,N_10278,N_10894);
nand U11798 (N_11798,N_10665,N_10070);
or U11799 (N_11799,N_10482,N_10666);
nand U11800 (N_11800,N_10502,N_10022);
nand U11801 (N_11801,N_10253,N_10961);
nand U11802 (N_11802,N_10279,N_10807);
xnor U11803 (N_11803,N_10428,N_10878);
or U11804 (N_11804,N_10782,N_10047);
and U11805 (N_11805,N_10966,N_10306);
nand U11806 (N_11806,N_10627,N_10474);
and U11807 (N_11807,N_10884,N_10403);
nor U11808 (N_11808,N_10219,N_10193);
xnor U11809 (N_11809,N_10164,N_10842);
and U11810 (N_11810,N_10834,N_10368);
xor U11811 (N_11811,N_10078,N_10561);
xor U11812 (N_11812,N_10004,N_10481);
or U11813 (N_11813,N_10940,N_10941);
nor U11814 (N_11814,N_10601,N_10824);
or U11815 (N_11815,N_10079,N_10939);
or U11816 (N_11816,N_10480,N_10776);
and U11817 (N_11817,N_10233,N_10242);
and U11818 (N_11818,N_10585,N_10639);
and U11819 (N_11819,N_10821,N_10552);
xnor U11820 (N_11820,N_10794,N_10677);
xnor U11821 (N_11821,N_10194,N_10002);
or U11822 (N_11822,N_10834,N_10321);
or U11823 (N_11823,N_10121,N_10573);
nor U11824 (N_11824,N_10199,N_10951);
xor U11825 (N_11825,N_10526,N_10113);
or U11826 (N_11826,N_10816,N_10324);
nor U11827 (N_11827,N_10180,N_10573);
xor U11828 (N_11828,N_10543,N_10026);
xor U11829 (N_11829,N_10476,N_10321);
and U11830 (N_11830,N_10845,N_10509);
or U11831 (N_11831,N_10356,N_10997);
and U11832 (N_11832,N_10941,N_10764);
nand U11833 (N_11833,N_10166,N_10398);
or U11834 (N_11834,N_10846,N_10971);
or U11835 (N_11835,N_10563,N_10133);
xor U11836 (N_11836,N_10864,N_10963);
nand U11837 (N_11837,N_10177,N_10710);
nand U11838 (N_11838,N_10189,N_10316);
nand U11839 (N_11839,N_10142,N_10063);
nor U11840 (N_11840,N_10763,N_10552);
nor U11841 (N_11841,N_10294,N_10970);
nand U11842 (N_11842,N_10428,N_10936);
nor U11843 (N_11843,N_10126,N_10184);
nand U11844 (N_11844,N_10867,N_10208);
nand U11845 (N_11845,N_10223,N_10394);
or U11846 (N_11846,N_10763,N_10862);
nor U11847 (N_11847,N_10300,N_10005);
xor U11848 (N_11848,N_10070,N_10430);
or U11849 (N_11849,N_10855,N_10136);
xor U11850 (N_11850,N_10555,N_10112);
xnor U11851 (N_11851,N_10814,N_10142);
xor U11852 (N_11852,N_10676,N_10851);
xnor U11853 (N_11853,N_10064,N_10665);
nor U11854 (N_11854,N_10782,N_10778);
xnor U11855 (N_11855,N_10892,N_10405);
or U11856 (N_11856,N_10542,N_10402);
or U11857 (N_11857,N_10084,N_10482);
and U11858 (N_11858,N_10290,N_10287);
nand U11859 (N_11859,N_10911,N_10240);
xor U11860 (N_11860,N_10513,N_10185);
xor U11861 (N_11861,N_10622,N_10195);
nand U11862 (N_11862,N_10803,N_10155);
or U11863 (N_11863,N_10594,N_10875);
nand U11864 (N_11864,N_10146,N_10243);
xor U11865 (N_11865,N_10119,N_10479);
nand U11866 (N_11866,N_10686,N_10786);
xnor U11867 (N_11867,N_10323,N_10365);
and U11868 (N_11868,N_10707,N_10734);
xor U11869 (N_11869,N_10455,N_10933);
nor U11870 (N_11870,N_10774,N_10711);
nand U11871 (N_11871,N_10148,N_10433);
nand U11872 (N_11872,N_10648,N_10302);
nor U11873 (N_11873,N_10498,N_10728);
and U11874 (N_11874,N_10712,N_10242);
nand U11875 (N_11875,N_10122,N_10540);
xnor U11876 (N_11876,N_10526,N_10532);
xor U11877 (N_11877,N_10644,N_10106);
nand U11878 (N_11878,N_10440,N_10173);
nand U11879 (N_11879,N_10244,N_10462);
and U11880 (N_11880,N_10876,N_10172);
xnor U11881 (N_11881,N_10318,N_10915);
nor U11882 (N_11882,N_10400,N_10466);
nand U11883 (N_11883,N_10896,N_10803);
and U11884 (N_11884,N_10362,N_10788);
and U11885 (N_11885,N_10580,N_10644);
nand U11886 (N_11886,N_10946,N_10986);
nand U11887 (N_11887,N_10125,N_10953);
nand U11888 (N_11888,N_10940,N_10505);
xor U11889 (N_11889,N_10547,N_10630);
nand U11890 (N_11890,N_10298,N_10128);
or U11891 (N_11891,N_10191,N_10499);
or U11892 (N_11892,N_10279,N_10697);
xor U11893 (N_11893,N_10876,N_10008);
or U11894 (N_11894,N_10364,N_10817);
nand U11895 (N_11895,N_10107,N_10384);
nand U11896 (N_11896,N_10979,N_10647);
and U11897 (N_11897,N_10950,N_10235);
xnor U11898 (N_11898,N_10694,N_10364);
and U11899 (N_11899,N_10654,N_10214);
xnor U11900 (N_11900,N_10913,N_10559);
and U11901 (N_11901,N_10934,N_10815);
nand U11902 (N_11902,N_10074,N_10429);
nor U11903 (N_11903,N_10429,N_10233);
nor U11904 (N_11904,N_10616,N_10443);
xor U11905 (N_11905,N_10307,N_10931);
nor U11906 (N_11906,N_10397,N_10005);
xor U11907 (N_11907,N_10296,N_10557);
xnor U11908 (N_11908,N_10071,N_10867);
or U11909 (N_11909,N_10845,N_10400);
nor U11910 (N_11910,N_10130,N_10324);
nand U11911 (N_11911,N_10320,N_10212);
xor U11912 (N_11912,N_10251,N_10176);
or U11913 (N_11913,N_10403,N_10689);
or U11914 (N_11914,N_10886,N_10215);
or U11915 (N_11915,N_10066,N_10810);
or U11916 (N_11916,N_10218,N_10273);
or U11917 (N_11917,N_10571,N_10584);
nor U11918 (N_11918,N_10333,N_10581);
xor U11919 (N_11919,N_10779,N_10728);
nand U11920 (N_11920,N_10721,N_10925);
xor U11921 (N_11921,N_10747,N_10599);
or U11922 (N_11922,N_10839,N_10965);
nand U11923 (N_11923,N_10615,N_10094);
and U11924 (N_11924,N_10485,N_10162);
nand U11925 (N_11925,N_10853,N_10762);
xor U11926 (N_11926,N_10603,N_10207);
and U11927 (N_11927,N_10432,N_10033);
and U11928 (N_11928,N_10640,N_10597);
and U11929 (N_11929,N_10918,N_10216);
xnor U11930 (N_11930,N_10437,N_10317);
nand U11931 (N_11931,N_10683,N_10693);
nand U11932 (N_11932,N_10893,N_10703);
or U11933 (N_11933,N_10763,N_10087);
nand U11934 (N_11934,N_10504,N_10642);
nor U11935 (N_11935,N_10611,N_10297);
and U11936 (N_11936,N_10390,N_10205);
nor U11937 (N_11937,N_10357,N_10128);
xnor U11938 (N_11938,N_10941,N_10808);
and U11939 (N_11939,N_10994,N_10713);
or U11940 (N_11940,N_10892,N_10834);
and U11941 (N_11941,N_10226,N_10875);
nand U11942 (N_11942,N_10419,N_10366);
and U11943 (N_11943,N_10936,N_10796);
xnor U11944 (N_11944,N_10538,N_10155);
or U11945 (N_11945,N_10512,N_10699);
xor U11946 (N_11946,N_10676,N_10608);
and U11947 (N_11947,N_10272,N_10330);
and U11948 (N_11948,N_10018,N_10864);
xor U11949 (N_11949,N_10704,N_10302);
nor U11950 (N_11950,N_10588,N_10802);
nand U11951 (N_11951,N_10257,N_10368);
xnor U11952 (N_11952,N_10488,N_10378);
and U11953 (N_11953,N_10332,N_10751);
xor U11954 (N_11954,N_10762,N_10783);
nand U11955 (N_11955,N_10770,N_10264);
nand U11956 (N_11956,N_10540,N_10376);
and U11957 (N_11957,N_10805,N_10630);
nand U11958 (N_11958,N_10963,N_10917);
nand U11959 (N_11959,N_10489,N_10033);
or U11960 (N_11960,N_10814,N_10152);
or U11961 (N_11961,N_10038,N_10518);
xnor U11962 (N_11962,N_10498,N_10424);
nand U11963 (N_11963,N_10452,N_10864);
and U11964 (N_11964,N_10797,N_10028);
nor U11965 (N_11965,N_10577,N_10989);
xnor U11966 (N_11966,N_10866,N_10944);
and U11967 (N_11967,N_10529,N_10260);
and U11968 (N_11968,N_10791,N_10332);
xnor U11969 (N_11969,N_10553,N_10343);
nand U11970 (N_11970,N_10442,N_10384);
nor U11971 (N_11971,N_10654,N_10240);
xor U11972 (N_11972,N_10406,N_10638);
nand U11973 (N_11973,N_10504,N_10776);
nand U11974 (N_11974,N_10671,N_10978);
nor U11975 (N_11975,N_10844,N_10706);
xor U11976 (N_11976,N_10170,N_10117);
xor U11977 (N_11977,N_10161,N_10940);
nor U11978 (N_11978,N_10912,N_10736);
and U11979 (N_11979,N_10126,N_10006);
and U11980 (N_11980,N_10756,N_10277);
or U11981 (N_11981,N_10883,N_10206);
nor U11982 (N_11982,N_10003,N_10298);
nor U11983 (N_11983,N_10730,N_10635);
and U11984 (N_11984,N_10912,N_10267);
nand U11985 (N_11985,N_10049,N_10678);
nand U11986 (N_11986,N_10046,N_10398);
nor U11987 (N_11987,N_10817,N_10873);
and U11988 (N_11988,N_10325,N_10171);
and U11989 (N_11989,N_10167,N_10451);
and U11990 (N_11990,N_10347,N_10669);
and U11991 (N_11991,N_10697,N_10505);
nor U11992 (N_11992,N_10162,N_10008);
nor U11993 (N_11993,N_10966,N_10111);
nor U11994 (N_11994,N_10431,N_10484);
xor U11995 (N_11995,N_10512,N_10702);
nor U11996 (N_11996,N_10709,N_10237);
nor U11997 (N_11997,N_10198,N_10447);
and U11998 (N_11998,N_10540,N_10783);
xor U11999 (N_11999,N_10887,N_10780);
or U12000 (N_12000,N_11551,N_11741);
or U12001 (N_12001,N_11698,N_11163);
xnor U12002 (N_12002,N_11338,N_11669);
or U12003 (N_12003,N_11681,N_11813);
nand U12004 (N_12004,N_11168,N_11581);
nor U12005 (N_12005,N_11991,N_11881);
xor U12006 (N_12006,N_11602,N_11816);
nor U12007 (N_12007,N_11738,N_11639);
nor U12008 (N_12008,N_11418,N_11927);
nand U12009 (N_12009,N_11643,N_11729);
xnor U12010 (N_12010,N_11705,N_11178);
nor U12011 (N_12011,N_11277,N_11149);
and U12012 (N_12012,N_11531,N_11518);
xnor U12013 (N_12013,N_11987,N_11345);
or U12014 (N_12014,N_11280,N_11533);
and U12015 (N_12015,N_11295,N_11799);
nor U12016 (N_12016,N_11771,N_11542);
xnor U12017 (N_12017,N_11644,N_11709);
and U12018 (N_12018,N_11624,N_11344);
nand U12019 (N_12019,N_11220,N_11475);
nor U12020 (N_12020,N_11300,N_11895);
xor U12021 (N_12021,N_11066,N_11386);
nor U12022 (N_12022,N_11399,N_11364);
nand U12023 (N_12023,N_11232,N_11155);
or U12024 (N_12024,N_11478,N_11564);
xor U12025 (N_12025,N_11527,N_11853);
nor U12026 (N_12026,N_11350,N_11878);
or U12027 (N_12027,N_11479,N_11875);
nor U12028 (N_12028,N_11710,N_11962);
or U12029 (N_12029,N_11638,N_11578);
nor U12030 (N_12030,N_11309,N_11267);
nor U12031 (N_12031,N_11359,N_11872);
xor U12032 (N_12032,N_11281,N_11038);
xor U12033 (N_12033,N_11867,N_11499);
and U12034 (N_12034,N_11282,N_11413);
nand U12035 (N_12035,N_11563,N_11079);
and U12036 (N_12036,N_11395,N_11166);
and U12037 (N_12037,N_11432,N_11194);
nand U12038 (N_12038,N_11251,N_11071);
nand U12039 (N_12039,N_11834,N_11275);
nand U12040 (N_12040,N_11529,N_11731);
xor U12041 (N_12041,N_11000,N_11798);
nor U12042 (N_12042,N_11102,N_11826);
and U12043 (N_12043,N_11692,N_11468);
nand U12044 (N_12044,N_11934,N_11494);
xnor U12045 (N_12045,N_11704,N_11080);
nor U12046 (N_12046,N_11109,N_11011);
and U12047 (N_12047,N_11185,N_11387);
xnor U12048 (N_12048,N_11752,N_11921);
nand U12049 (N_12049,N_11792,N_11288);
and U12050 (N_12050,N_11258,N_11960);
nand U12051 (N_12051,N_11748,N_11247);
xnor U12052 (N_12052,N_11898,N_11668);
xor U12053 (N_12053,N_11977,N_11595);
nand U12054 (N_12054,N_11158,N_11538);
or U12055 (N_12055,N_11459,N_11957);
and U12056 (N_12056,N_11544,N_11983);
nand U12057 (N_12057,N_11375,N_11981);
xnor U12058 (N_12058,N_11691,N_11125);
and U12059 (N_12059,N_11753,N_11605);
or U12060 (N_12060,N_11706,N_11507);
or U12061 (N_12061,N_11371,N_11808);
nand U12062 (N_12062,N_11008,N_11276);
and U12063 (N_12063,N_11268,N_11296);
xor U12064 (N_12064,N_11539,N_11416);
and U12065 (N_12065,N_11697,N_11683);
nand U12066 (N_12066,N_11606,N_11471);
nor U12067 (N_12067,N_11757,N_11390);
and U12068 (N_12068,N_11336,N_11262);
and U12069 (N_12069,N_11222,N_11716);
or U12070 (N_12070,N_11754,N_11591);
and U12071 (N_12071,N_11391,N_11209);
nor U12072 (N_12072,N_11679,N_11273);
nor U12073 (N_12073,N_11477,N_11961);
and U12074 (N_12074,N_11810,N_11448);
or U12075 (N_12075,N_11920,N_11956);
nor U12076 (N_12076,N_11848,N_11924);
or U12077 (N_12077,N_11649,N_11984);
and U12078 (N_12078,N_11233,N_11690);
xor U12079 (N_12079,N_11728,N_11935);
nor U12080 (N_12080,N_11022,N_11536);
nand U12081 (N_12081,N_11031,N_11851);
xnor U12082 (N_12082,N_11820,N_11381);
nor U12083 (N_12083,N_11549,N_11244);
and U12084 (N_12084,N_11756,N_11883);
nor U12085 (N_12085,N_11594,N_11617);
nor U12086 (N_12086,N_11372,N_11948);
and U12087 (N_12087,N_11772,N_11596);
and U12088 (N_12088,N_11138,N_11737);
xor U12089 (N_12089,N_11331,N_11455);
and U12090 (N_12090,N_11763,N_11714);
or U12091 (N_12091,N_11522,N_11629);
nand U12092 (N_12092,N_11648,N_11365);
or U12093 (N_12093,N_11685,N_11625);
nor U12094 (N_12094,N_11990,N_11446);
or U12095 (N_12095,N_11501,N_11259);
or U12096 (N_12096,N_11909,N_11561);
nand U12097 (N_12097,N_11623,N_11918);
or U12098 (N_12098,N_11192,N_11287);
nor U12099 (N_12099,N_11923,N_11779);
xor U12100 (N_12100,N_11374,N_11767);
or U12101 (N_12101,N_11874,N_11958);
xnor U12102 (N_12102,N_11148,N_11833);
nor U12103 (N_12103,N_11274,N_11318);
or U12104 (N_12104,N_11900,N_11117);
or U12105 (N_12105,N_11089,N_11060);
nor U12106 (N_12106,N_11887,N_11032);
nor U12107 (N_12107,N_11812,N_11963);
nor U12108 (N_12108,N_11165,N_11124);
xnor U12109 (N_12109,N_11310,N_11830);
xor U12110 (N_12110,N_11122,N_11746);
or U12111 (N_12111,N_11204,N_11431);
nand U12112 (N_12112,N_11588,N_11425);
nor U12113 (N_12113,N_11463,N_11469);
nand U12114 (N_12114,N_11755,N_11028);
nand U12115 (N_12115,N_11975,N_11422);
nand U12116 (N_12116,N_11645,N_11540);
and U12117 (N_12117,N_11996,N_11770);
nor U12118 (N_12118,N_11176,N_11559);
nor U12119 (N_12119,N_11968,N_11742);
or U12120 (N_12120,N_11653,N_11328);
nor U12121 (N_12121,N_11511,N_11712);
and U12122 (N_12122,N_11857,N_11067);
nor U12123 (N_12123,N_11910,N_11864);
and U12124 (N_12124,N_11330,N_11440);
xnor U12125 (N_12125,N_11946,N_11264);
xor U12126 (N_12126,N_11238,N_11868);
nor U12127 (N_12127,N_11576,N_11243);
nand U12128 (N_12128,N_11284,N_11674);
and U12129 (N_12129,N_11135,N_11351);
nand U12130 (N_12130,N_11676,N_11804);
or U12131 (N_12131,N_11096,N_11519);
or U12132 (N_12132,N_11419,N_11579);
and U12133 (N_12133,N_11120,N_11686);
and U12134 (N_12134,N_11814,N_11570);
nand U12135 (N_12135,N_11836,N_11959);
xor U12136 (N_12136,N_11435,N_11408);
xnor U12137 (N_12137,N_11670,N_11535);
or U12138 (N_12138,N_11450,N_11907);
nor U12139 (N_12139,N_11411,N_11896);
nand U12140 (N_12140,N_11472,N_11389);
xor U12141 (N_12141,N_11208,N_11634);
nor U12142 (N_12142,N_11307,N_11483);
nor U12143 (N_12143,N_11304,N_11825);
or U12144 (N_12144,N_11270,N_11203);
nand U12145 (N_12145,N_11917,N_11689);
xnor U12146 (N_12146,N_11552,N_11950);
or U12147 (N_12147,N_11018,N_11794);
nor U12148 (N_12148,N_11377,N_11073);
nor U12149 (N_12149,N_11888,N_11778);
nand U12150 (N_12150,N_11156,N_11303);
and U12151 (N_12151,N_11436,N_11157);
xnor U12152 (N_12152,N_11574,N_11662);
nand U12153 (N_12153,N_11914,N_11201);
nand U12154 (N_12154,N_11041,N_11005);
nand U12155 (N_12155,N_11725,N_11903);
xnor U12156 (N_12156,N_11272,N_11530);
nand U12157 (N_12157,N_11837,N_11189);
nor U12158 (N_12158,N_11735,N_11183);
nand U12159 (N_12159,N_11719,N_11140);
nand U12160 (N_12160,N_11932,N_11488);
and U12161 (N_12161,N_11131,N_11765);
or U12162 (N_12162,N_11610,N_11460);
nor U12163 (N_12163,N_11589,N_11327);
xnor U12164 (N_12164,N_11323,N_11911);
xor U12165 (N_12165,N_11392,N_11835);
nand U12166 (N_12166,N_11050,N_11555);
nor U12167 (N_12167,N_11180,N_11760);
and U12168 (N_12168,N_11361,N_11711);
nand U12169 (N_12169,N_11926,N_11401);
or U12170 (N_12170,N_11657,N_11147);
nor U12171 (N_12171,N_11225,N_11029);
nand U12172 (N_12172,N_11791,N_11191);
or U12173 (N_12173,N_11179,N_11046);
nand U12174 (N_12174,N_11199,N_11663);
or U12175 (N_12175,N_11904,N_11249);
and U12176 (N_12176,N_11487,N_11315);
nor U12177 (N_12177,N_11115,N_11116);
or U12178 (N_12178,N_11062,N_11747);
nor U12179 (N_12179,N_11575,N_11154);
nor U12180 (N_12180,N_11906,N_11396);
or U12181 (N_12181,N_11236,N_11177);
nand U12182 (N_12182,N_11023,N_11762);
and U12183 (N_12183,N_11652,N_11495);
nor U12184 (N_12184,N_11072,N_11940);
or U12185 (N_12185,N_11929,N_11491);
or U12186 (N_12186,N_11609,N_11290);
and U12187 (N_12187,N_11466,N_11036);
or U12188 (N_12188,N_11231,N_11811);
or U12189 (N_12189,N_11724,N_11357);
nand U12190 (N_12190,N_11085,N_11912);
xor U12191 (N_12191,N_11127,N_11286);
nor U12192 (N_12192,N_11126,N_11097);
or U12193 (N_12193,N_11997,N_11415);
and U12194 (N_12194,N_11393,N_11133);
nor U12195 (N_12195,N_11894,N_11088);
nand U12196 (N_12196,N_11721,N_11658);
xor U12197 (N_12197,N_11534,N_11618);
xor U12198 (N_12198,N_11458,N_11356);
or U12199 (N_12199,N_11640,N_11103);
nand U12200 (N_12200,N_11931,N_11995);
nor U12201 (N_12201,N_11597,N_11047);
nand U12202 (N_12202,N_11437,N_11449);
nand U12203 (N_12203,N_11426,N_11637);
nand U12204 (N_12204,N_11945,N_11385);
nor U12205 (N_12205,N_11780,N_11806);
nand U12206 (N_12206,N_11938,N_11882);
or U12207 (N_12207,N_11944,N_11665);
xor U12208 (N_12208,N_11279,N_11305);
and U12209 (N_12209,N_11630,N_11604);
or U12210 (N_12210,N_11560,N_11844);
and U12211 (N_12211,N_11420,N_11892);
nand U12212 (N_12212,N_11291,N_11992);
and U12213 (N_12213,N_11383,N_11394);
xnor U12214 (N_12214,N_11334,N_11659);
nor U12215 (N_12215,N_11758,N_11039);
xor U12216 (N_12216,N_11664,N_11819);
and U12217 (N_12217,N_11335,N_11119);
nor U12218 (N_12218,N_11308,N_11212);
xor U12219 (N_12219,N_11366,N_11130);
nor U12220 (N_12220,N_11797,N_11558);
or U12221 (N_12221,N_11615,N_11289);
nand U12222 (N_12222,N_11986,N_11084);
or U12223 (N_12223,N_11150,N_11592);
and U12224 (N_12224,N_11255,N_11726);
or U12225 (N_12225,N_11614,N_11314);
or U12226 (N_12226,N_11207,N_11749);
and U12227 (N_12227,N_11025,N_11769);
or U12228 (N_12228,N_11347,N_11840);
xor U12229 (N_12229,N_11325,N_11058);
or U12230 (N_12230,N_11684,N_11490);
nand U12231 (N_12231,N_11661,N_11734);
and U12232 (N_12232,N_11053,N_11521);
or U12233 (N_12233,N_11456,N_11673);
nand U12234 (N_12234,N_11817,N_11562);
or U12235 (N_12235,N_11173,N_11134);
nor U12236 (N_12236,N_11302,N_11144);
nand U12237 (N_12237,N_11856,N_11573);
nor U12238 (N_12238,N_11197,N_11656);
or U12239 (N_12239,N_11680,N_11342);
nor U12240 (N_12240,N_11877,N_11925);
nor U12241 (N_12241,N_11633,N_11785);
or U12242 (N_12242,N_11108,N_11548);
nand U12243 (N_12243,N_11500,N_11660);
or U12244 (N_12244,N_11332,N_11846);
and U12245 (N_12245,N_11566,N_11568);
and U12246 (N_12246,N_11751,N_11464);
and U12247 (N_12247,N_11441,N_11513);
nor U12248 (N_12248,N_11118,N_11821);
xor U12249 (N_12249,N_11476,N_11526);
nor U12250 (N_12250,N_11405,N_11145);
nor U12251 (N_12251,N_11717,N_11363);
nand U12252 (N_12252,N_11261,N_11482);
or U12253 (N_12253,N_11442,N_11015);
nor U12254 (N_12254,N_11354,N_11498);
xnor U12255 (N_12255,N_11257,N_11107);
nand U12256 (N_12256,N_11254,N_11505);
nand U12257 (N_12257,N_11739,N_11021);
xor U12258 (N_12258,N_11019,N_11245);
xor U12259 (N_12259,N_11326,N_11210);
xnor U12260 (N_12260,N_11790,N_11489);
nand U12261 (N_12261,N_11933,N_11905);
nor U12262 (N_12262,N_11828,N_11452);
nor U12263 (N_12263,N_11265,N_11824);
and U12264 (N_12264,N_11172,N_11626);
nor U12265 (N_12265,N_11317,N_11859);
nor U12266 (N_12266,N_11915,N_11064);
and U12267 (N_12267,N_11226,N_11993);
nand U12268 (N_12268,N_11744,N_11202);
and U12269 (N_12269,N_11211,N_11502);
nand U12270 (N_12270,N_11111,N_11414);
nand U12271 (N_12271,N_11873,N_11473);
and U12272 (N_12272,N_11943,N_11380);
nor U12273 (N_12273,N_11708,N_11044);
and U12274 (N_12274,N_11234,N_11313);
and U12275 (N_12275,N_11321,N_11040);
xor U12276 (N_12276,N_11852,N_11947);
and U12277 (N_12277,N_11515,N_11786);
or U12278 (N_12278,N_11557,N_11299);
or U12279 (N_12279,N_11889,N_11409);
xnor U12280 (N_12280,N_11871,N_11893);
nor U12281 (N_12281,N_11182,N_11775);
xnor U12282 (N_12282,N_11695,N_11913);
and U12283 (N_12283,N_11707,N_11675);
nor U12284 (N_12284,N_11082,N_11567);
nand U12285 (N_12285,N_11620,N_11009);
or U12286 (N_12286,N_11743,N_11965);
nand U12287 (N_12287,N_11546,N_11086);
or U12288 (N_12288,N_11899,N_11042);
nand U12289 (N_12289,N_11964,N_11988);
nor U12290 (N_12290,N_11013,N_11438);
nor U12291 (N_12291,N_11443,N_11402);
or U12292 (N_12292,N_11523,N_11196);
and U12293 (N_12293,N_11901,N_11585);
or U12294 (N_12294,N_11745,N_11727);
nor U12295 (N_12295,N_11693,N_11781);
nor U12296 (N_12296,N_11237,N_11908);
nor U12297 (N_12297,N_11035,N_11492);
nand U12298 (N_12298,N_11167,N_11667);
xor U12299 (N_12299,N_11271,N_11324);
xor U12300 (N_12300,N_11016,N_11001);
xnor U12301 (N_12301,N_11571,N_11121);
nand U12302 (N_12302,N_11517,N_11229);
or U12303 (N_12303,N_11541,N_11666);
or U12304 (N_12304,N_11930,N_11553);
xnor U12305 (N_12305,N_11699,N_11181);
or U12306 (N_12306,N_11362,N_11343);
nand U12307 (N_12307,N_11049,N_11942);
nor U12308 (N_12308,N_11428,N_11355);
nor U12309 (N_12309,N_11230,N_11537);
and U12310 (N_12310,N_11764,N_11235);
nor U12311 (N_12311,N_11429,N_11221);
or U12312 (N_12312,N_11885,N_11104);
xnor U12313 (N_12313,N_11936,N_11481);
and U12314 (N_12314,N_11004,N_11205);
nor U12315 (N_12315,N_11074,N_11353);
or U12316 (N_12316,N_11090,N_11854);
or U12317 (N_12317,N_11136,N_11801);
or U12318 (N_12318,N_11627,N_11520);
nand U12319 (N_12319,N_11789,N_11554);
nand U12320 (N_12320,N_11855,N_11188);
xor U12321 (N_12321,N_11105,N_11723);
nor U12322 (N_12322,N_11916,N_11654);
and U12323 (N_12323,N_11454,N_11101);
or U12324 (N_12324,N_11439,N_11195);
nand U12325 (N_12325,N_11715,N_11075);
and U12326 (N_12326,N_11713,N_11333);
xor U12327 (N_12327,N_11818,N_11922);
and U12328 (N_12328,N_11784,N_11832);
or U12329 (N_12329,N_11974,N_11512);
and U12330 (N_12330,N_11616,N_11151);
or U12331 (N_12331,N_11170,N_11003);
xor U12332 (N_12332,N_11768,N_11051);
nor U12333 (N_12333,N_11349,N_11174);
and U12334 (N_12334,N_11462,N_11341);
and U12335 (N_12335,N_11953,N_11822);
and U12336 (N_12336,N_11774,N_11807);
and U12337 (N_12337,N_11358,N_11582);
nor U12338 (N_12338,N_11897,N_11378);
and U12339 (N_12339,N_11928,N_11382);
and U12340 (N_12340,N_11092,N_11516);
nor U12341 (N_12341,N_11006,N_11860);
or U12342 (N_12342,N_11858,N_11982);
xnor U12343 (N_12343,N_11583,N_11269);
or U12344 (N_12344,N_11651,N_11007);
xor U12345 (N_12345,N_11162,N_11447);
or U12346 (N_12346,N_11186,N_11384);
nor U12347 (N_12347,N_11761,N_11146);
nand U12348 (N_12348,N_11445,N_11219);
and U12349 (N_12349,N_11030,N_11367);
nand U12350 (N_12350,N_11580,N_11532);
and U12351 (N_12351,N_11677,N_11052);
xor U12352 (N_12352,N_11292,N_11622);
xor U12353 (N_12353,N_11503,N_11223);
xor U12354 (N_12354,N_11862,N_11525);
nor U12355 (N_12355,N_11671,N_11973);
or U12356 (N_12356,N_11966,N_11444);
nor U12357 (N_12357,N_11952,N_11421);
xnor U12358 (N_12358,N_11206,N_11024);
nor U12359 (N_12359,N_11619,N_11057);
nor U12360 (N_12360,N_11193,N_11528);
or U12361 (N_12361,N_11607,N_11647);
or U12362 (N_12362,N_11985,N_11218);
nand U12363 (N_12363,N_11484,N_11010);
nor U12364 (N_12364,N_11087,N_11863);
nor U12365 (N_12365,N_11636,N_11400);
nor U12366 (N_12366,N_11750,N_11045);
and U12367 (N_12367,N_11322,N_11027);
nand U12368 (N_12368,N_11672,N_11593);
nand U12369 (N_12369,N_11352,N_11070);
and U12370 (N_12370,N_11083,N_11252);
nand U12371 (N_12371,N_11632,N_11129);
nor U12372 (N_12372,N_11847,N_11843);
and U12373 (N_12373,N_11424,N_11348);
or U12374 (N_12374,N_11506,N_11340);
nand U12375 (N_12375,N_11740,N_11655);
nand U12376 (N_12376,N_11989,N_11687);
nor U12377 (N_12377,N_11621,N_11599);
or U12378 (N_12378,N_11635,N_11720);
nand U12379 (N_12379,N_11081,N_11803);
nand U12380 (N_12380,N_11838,N_11870);
nor U12381 (N_12381,N_11733,N_11410);
or U12382 (N_12382,N_11514,N_11586);
and U12383 (N_12383,N_11628,N_11631);
nand U12384 (N_12384,N_11346,N_11978);
nand U12385 (N_12385,N_11998,N_11078);
and U12386 (N_12386,N_11972,N_11373);
and U12387 (N_12387,N_11971,N_11565);
nor U12388 (N_12388,N_11423,N_11815);
nor U12389 (N_12389,N_11955,N_11161);
or U12390 (N_12390,N_11598,N_11169);
xor U12391 (N_12391,N_11865,N_11246);
xnor U12392 (N_12392,N_11869,N_11248);
and U12393 (N_12393,N_11612,N_11164);
or U12394 (N_12394,N_11298,N_11465);
xor U12395 (N_12395,N_11260,N_11278);
and U12396 (N_12396,N_11091,N_11783);
and U12397 (N_12397,N_11369,N_11970);
xor U12398 (N_12398,N_11608,N_11239);
and U12399 (N_12399,N_11250,N_11433);
nand U12400 (N_12400,N_11611,N_11795);
and U12401 (N_12401,N_11782,N_11879);
nand U12402 (N_12402,N_11153,N_11474);
or U12403 (N_12403,N_11451,N_11880);
and U12404 (N_12404,N_11417,N_11316);
xor U12405 (N_12405,N_11509,N_11601);
nor U12406 (N_12406,N_11099,N_11732);
nor U12407 (N_12407,N_11069,N_11886);
or U12408 (N_12408,N_11379,N_11113);
nor U12409 (N_12409,N_11641,N_11137);
and U12410 (N_12410,N_11954,N_11603);
xnor U12411 (N_12411,N_11823,N_11730);
nor U12412 (N_12412,N_11160,N_11227);
nor U12413 (N_12413,N_11951,N_11510);
xnor U12414 (N_12414,N_11020,N_11702);
or U12415 (N_12415,N_11545,N_11240);
and U12416 (N_12416,N_11068,N_11937);
nand U12417 (N_12417,N_11175,N_11486);
or U12418 (N_12418,N_11123,N_11796);
xnor U12419 (N_12419,N_11829,N_11388);
nand U12420 (N_12420,N_11026,N_11061);
and U12421 (N_12421,N_11547,N_11569);
nor U12422 (N_12422,N_11839,N_11694);
nand U12423 (N_12423,N_11320,N_11600);
xor U12424 (N_12424,N_11736,N_11056);
nand U12425 (N_12425,N_11093,N_11141);
and U12426 (N_12426,N_11397,N_11033);
nand U12427 (N_12427,N_11866,N_11453);
xnor U12428 (N_12428,N_11059,N_11646);
nor U12429 (N_12429,N_11339,N_11017);
xor U12430 (N_12430,N_11171,N_11703);
nor U12431 (N_12431,N_11398,N_11360);
and U12432 (N_12432,N_11048,N_11979);
xor U12433 (N_12433,N_11200,N_11550);
nor U12434 (N_12434,N_11508,N_11682);
or U12435 (N_12435,N_11902,N_11132);
or U12436 (N_12436,N_11480,N_11297);
nand U12437 (N_12437,N_11311,N_11941);
nor U12438 (N_12438,N_11114,N_11831);
nor U12439 (N_12439,N_11301,N_11190);
nand U12440 (N_12440,N_11215,N_11337);
or U12441 (N_12441,N_11577,N_11587);
nand U12442 (N_12442,N_11773,N_11100);
xnor U12443 (N_12443,N_11043,N_11407);
or U12444 (N_12444,N_11994,N_11312);
nor U12445 (N_12445,N_11294,N_11037);
and U12446 (N_12446,N_11406,N_11063);
nor U12447 (N_12447,N_11805,N_11077);
or U12448 (N_12448,N_11696,N_11319);
or U12449 (N_12449,N_11700,N_11143);
or U12450 (N_12450,N_11034,N_11678);
nand U12451 (N_12451,N_11430,N_11461);
or U12452 (N_12452,N_11584,N_11054);
and U12453 (N_12453,N_11827,N_11110);
nand U12454 (N_12454,N_11776,N_11404);
and U12455 (N_12455,N_11939,N_11841);
nor U12456 (N_12456,N_11376,N_11242);
nor U12457 (N_12457,N_11139,N_11787);
nor U12458 (N_12458,N_11434,N_11216);
nor U12459 (N_12459,N_11845,N_11142);
xor U12460 (N_12460,N_11777,N_11403);
nand U12461 (N_12461,N_11504,N_11800);
and U12462 (N_12462,N_11493,N_11224);
nand U12463 (N_12463,N_11228,N_11470);
and U12464 (N_12464,N_11128,N_11650);
and U12465 (N_12465,N_11688,N_11976);
xor U12466 (N_12466,N_11293,N_11980);
xnor U12467 (N_12467,N_11266,N_11967);
nor U12468 (N_12468,N_11217,N_11949);
nand U12469 (N_12469,N_11497,N_11524);
nor U12470 (N_12470,N_11861,N_11809);
nor U12471 (N_12471,N_11368,N_11718);
xnor U12472 (N_12472,N_11722,N_11891);
xor U12473 (N_12473,N_11969,N_11094);
nand U12474 (N_12474,N_11112,N_11543);
xnor U12475 (N_12475,N_11642,N_11412);
nand U12476 (N_12476,N_11842,N_11241);
nand U12477 (N_12477,N_11014,N_11065);
or U12478 (N_12478,N_11802,N_11919);
xnor U12479 (N_12479,N_11214,N_11613);
xnor U12480 (N_12480,N_11590,N_11184);
or U12481 (N_12481,N_11766,N_11572);
xnor U12482 (N_12482,N_11876,N_11098);
nand U12483 (N_12483,N_11457,N_11253);
nor U12484 (N_12484,N_11095,N_11999);
or U12485 (N_12485,N_11427,N_11759);
nand U12486 (N_12486,N_11285,N_11198);
xnor U12487 (N_12487,N_11306,N_11701);
xor U12488 (N_12488,N_11850,N_11788);
nand U12489 (N_12489,N_11055,N_11849);
xor U12490 (N_12490,N_11159,N_11213);
xnor U12491 (N_12491,N_11187,N_11012);
xor U12492 (N_12492,N_11485,N_11496);
or U12493 (N_12493,N_11076,N_11263);
nor U12494 (N_12494,N_11556,N_11884);
or U12495 (N_12495,N_11106,N_11793);
nor U12496 (N_12496,N_11467,N_11256);
and U12497 (N_12497,N_11329,N_11370);
nand U12498 (N_12498,N_11002,N_11890);
nor U12499 (N_12499,N_11283,N_11152);
or U12500 (N_12500,N_11097,N_11717);
and U12501 (N_12501,N_11740,N_11026);
and U12502 (N_12502,N_11069,N_11697);
or U12503 (N_12503,N_11476,N_11519);
nand U12504 (N_12504,N_11754,N_11816);
or U12505 (N_12505,N_11946,N_11766);
nand U12506 (N_12506,N_11979,N_11925);
nand U12507 (N_12507,N_11488,N_11792);
nor U12508 (N_12508,N_11857,N_11622);
and U12509 (N_12509,N_11251,N_11379);
xor U12510 (N_12510,N_11516,N_11385);
nor U12511 (N_12511,N_11219,N_11274);
xnor U12512 (N_12512,N_11690,N_11993);
xnor U12513 (N_12513,N_11691,N_11784);
nor U12514 (N_12514,N_11331,N_11759);
or U12515 (N_12515,N_11920,N_11327);
or U12516 (N_12516,N_11520,N_11822);
nand U12517 (N_12517,N_11660,N_11829);
xnor U12518 (N_12518,N_11990,N_11501);
nor U12519 (N_12519,N_11801,N_11239);
nand U12520 (N_12520,N_11306,N_11873);
or U12521 (N_12521,N_11874,N_11934);
or U12522 (N_12522,N_11438,N_11648);
xnor U12523 (N_12523,N_11137,N_11060);
nand U12524 (N_12524,N_11239,N_11524);
or U12525 (N_12525,N_11649,N_11925);
xnor U12526 (N_12526,N_11165,N_11549);
nor U12527 (N_12527,N_11935,N_11640);
nand U12528 (N_12528,N_11757,N_11881);
and U12529 (N_12529,N_11233,N_11274);
or U12530 (N_12530,N_11527,N_11656);
nor U12531 (N_12531,N_11213,N_11218);
nor U12532 (N_12532,N_11195,N_11143);
nor U12533 (N_12533,N_11548,N_11547);
or U12534 (N_12534,N_11884,N_11409);
or U12535 (N_12535,N_11342,N_11815);
xor U12536 (N_12536,N_11553,N_11320);
and U12537 (N_12537,N_11002,N_11932);
nor U12538 (N_12538,N_11441,N_11780);
nor U12539 (N_12539,N_11413,N_11814);
nand U12540 (N_12540,N_11899,N_11320);
or U12541 (N_12541,N_11369,N_11390);
and U12542 (N_12542,N_11569,N_11966);
and U12543 (N_12543,N_11265,N_11166);
and U12544 (N_12544,N_11888,N_11601);
nand U12545 (N_12545,N_11479,N_11067);
nor U12546 (N_12546,N_11145,N_11649);
and U12547 (N_12547,N_11644,N_11267);
or U12548 (N_12548,N_11472,N_11134);
nor U12549 (N_12549,N_11028,N_11828);
and U12550 (N_12550,N_11692,N_11345);
or U12551 (N_12551,N_11712,N_11437);
nand U12552 (N_12552,N_11397,N_11024);
nand U12553 (N_12553,N_11575,N_11851);
nand U12554 (N_12554,N_11285,N_11846);
or U12555 (N_12555,N_11879,N_11177);
or U12556 (N_12556,N_11751,N_11052);
nor U12557 (N_12557,N_11308,N_11231);
or U12558 (N_12558,N_11931,N_11485);
or U12559 (N_12559,N_11878,N_11415);
xnor U12560 (N_12560,N_11671,N_11994);
nand U12561 (N_12561,N_11803,N_11629);
nor U12562 (N_12562,N_11075,N_11136);
or U12563 (N_12563,N_11878,N_11677);
nor U12564 (N_12564,N_11014,N_11279);
and U12565 (N_12565,N_11535,N_11356);
or U12566 (N_12566,N_11931,N_11494);
or U12567 (N_12567,N_11842,N_11182);
and U12568 (N_12568,N_11417,N_11207);
and U12569 (N_12569,N_11436,N_11814);
and U12570 (N_12570,N_11588,N_11822);
or U12571 (N_12571,N_11966,N_11062);
nand U12572 (N_12572,N_11816,N_11402);
nand U12573 (N_12573,N_11670,N_11095);
nor U12574 (N_12574,N_11071,N_11176);
nor U12575 (N_12575,N_11860,N_11620);
nand U12576 (N_12576,N_11245,N_11273);
and U12577 (N_12577,N_11630,N_11670);
nand U12578 (N_12578,N_11875,N_11822);
nor U12579 (N_12579,N_11577,N_11525);
nor U12580 (N_12580,N_11213,N_11955);
xor U12581 (N_12581,N_11301,N_11748);
xor U12582 (N_12582,N_11480,N_11333);
or U12583 (N_12583,N_11150,N_11363);
xor U12584 (N_12584,N_11946,N_11178);
xor U12585 (N_12585,N_11582,N_11469);
or U12586 (N_12586,N_11018,N_11930);
nor U12587 (N_12587,N_11602,N_11365);
nand U12588 (N_12588,N_11792,N_11455);
xnor U12589 (N_12589,N_11199,N_11776);
xor U12590 (N_12590,N_11816,N_11297);
and U12591 (N_12591,N_11881,N_11184);
xor U12592 (N_12592,N_11767,N_11500);
or U12593 (N_12593,N_11766,N_11624);
and U12594 (N_12594,N_11739,N_11440);
nand U12595 (N_12595,N_11751,N_11317);
nor U12596 (N_12596,N_11295,N_11731);
xnor U12597 (N_12597,N_11148,N_11411);
xnor U12598 (N_12598,N_11144,N_11333);
xor U12599 (N_12599,N_11632,N_11479);
nand U12600 (N_12600,N_11029,N_11927);
and U12601 (N_12601,N_11834,N_11982);
xor U12602 (N_12602,N_11808,N_11732);
nor U12603 (N_12603,N_11694,N_11780);
xnor U12604 (N_12604,N_11432,N_11378);
and U12605 (N_12605,N_11014,N_11467);
nand U12606 (N_12606,N_11418,N_11661);
or U12607 (N_12607,N_11598,N_11399);
nand U12608 (N_12608,N_11304,N_11790);
and U12609 (N_12609,N_11098,N_11561);
nor U12610 (N_12610,N_11374,N_11695);
nand U12611 (N_12611,N_11267,N_11581);
and U12612 (N_12612,N_11872,N_11715);
or U12613 (N_12613,N_11442,N_11597);
nor U12614 (N_12614,N_11920,N_11877);
nor U12615 (N_12615,N_11893,N_11960);
nand U12616 (N_12616,N_11351,N_11342);
xor U12617 (N_12617,N_11231,N_11373);
xnor U12618 (N_12618,N_11157,N_11885);
or U12619 (N_12619,N_11709,N_11423);
and U12620 (N_12620,N_11443,N_11274);
or U12621 (N_12621,N_11860,N_11214);
nor U12622 (N_12622,N_11775,N_11904);
nand U12623 (N_12623,N_11885,N_11225);
or U12624 (N_12624,N_11000,N_11449);
xor U12625 (N_12625,N_11465,N_11791);
or U12626 (N_12626,N_11006,N_11334);
or U12627 (N_12627,N_11139,N_11046);
and U12628 (N_12628,N_11820,N_11678);
and U12629 (N_12629,N_11164,N_11154);
and U12630 (N_12630,N_11812,N_11705);
or U12631 (N_12631,N_11046,N_11616);
nand U12632 (N_12632,N_11917,N_11063);
nor U12633 (N_12633,N_11274,N_11828);
or U12634 (N_12634,N_11361,N_11034);
xor U12635 (N_12635,N_11596,N_11151);
or U12636 (N_12636,N_11374,N_11976);
and U12637 (N_12637,N_11962,N_11182);
or U12638 (N_12638,N_11273,N_11422);
xnor U12639 (N_12639,N_11827,N_11676);
nand U12640 (N_12640,N_11700,N_11545);
nor U12641 (N_12641,N_11028,N_11471);
or U12642 (N_12642,N_11304,N_11991);
or U12643 (N_12643,N_11390,N_11527);
xor U12644 (N_12644,N_11929,N_11639);
and U12645 (N_12645,N_11899,N_11532);
nand U12646 (N_12646,N_11913,N_11334);
nand U12647 (N_12647,N_11974,N_11604);
xnor U12648 (N_12648,N_11073,N_11053);
nand U12649 (N_12649,N_11522,N_11685);
xor U12650 (N_12650,N_11028,N_11146);
nand U12651 (N_12651,N_11711,N_11877);
or U12652 (N_12652,N_11486,N_11604);
nand U12653 (N_12653,N_11762,N_11320);
xor U12654 (N_12654,N_11370,N_11091);
xor U12655 (N_12655,N_11095,N_11689);
xnor U12656 (N_12656,N_11263,N_11259);
nor U12657 (N_12657,N_11028,N_11166);
nor U12658 (N_12658,N_11967,N_11464);
nand U12659 (N_12659,N_11591,N_11683);
nand U12660 (N_12660,N_11765,N_11301);
xor U12661 (N_12661,N_11927,N_11705);
nor U12662 (N_12662,N_11342,N_11045);
and U12663 (N_12663,N_11710,N_11154);
xnor U12664 (N_12664,N_11080,N_11244);
nor U12665 (N_12665,N_11664,N_11056);
nor U12666 (N_12666,N_11397,N_11528);
and U12667 (N_12667,N_11523,N_11468);
and U12668 (N_12668,N_11508,N_11399);
nand U12669 (N_12669,N_11319,N_11492);
xor U12670 (N_12670,N_11406,N_11126);
and U12671 (N_12671,N_11729,N_11377);
xnor U12672 (N_12672,N_11195,N_11995);
or U12673 (N_12673,N_11860,N_11193);
xor U12674 (N_12674,N_11904,N_11611);
nor U12675 (N_12675,N_11031,N_11561);
nor U12676 (N_12676,N_11639,N_11061);
or U12677 (N_12677,N_11823,N_11791);
or U12678 (N_12678,N_11463,N_11342);
and U12679 (N_12679,N_11005,N_11330);
nor U12680 (N_12680,N_11520,N_11760);
or U12681 (N_12681,N_11314,N_11308);
nand U12682 (N_12682,N_11910,N_11648);
and U12683 (N_12683,N_11965,N_11686);
nor U12684 (N_12684,N_11589,N_11762);
xor U12685 (N_12685,N_11153,N_11963);
and U12686 (N_12686,N_11779,N_11025);
nor U12687 (N_12687,N_11453,N_11892);
or U12688 (N_12688,N_11684,N_11699);
nor U12689 (N_12689,N_11220,N_11758);
and U12690 (N_12690,N_11963,N_11429);
nor U12691 (N_12691,N_11142,N_11027);
and U12692 (N_12692,N_11863,N_11354);
nand U12693 (N_12693,N_11543,N_11989);
nand U12694 (N_12694,N_11754,N_11099);
and U12695 (N_12695,N_11845,N_11966);
nor U12696 (N_12696,N_11712,N_11963);
or U12697 (N_12697,N_11516,N_11046);
nand U12698 (N_12698,N_11789,N_11612);
nor U12699 (N_12699,N_11236,N_11479);
nor U12700 (N_12700,N_11893,N_11418);
nand U12701 (N_12701,N_11131,N_11835);
and U12702 (N_12702,N_11308,N_11657);
xnor U12703 (N_12703,N_11651,N_11921);
nor U12704 (N_12704,N_11535,N_11865);
or U12705 (N_12705,N_11819,N_11945);
nand U12706 (N_12706,N_11834,N_11727);
nand U12707 (N_12707,N_11030,N_11405);
xor U12708 (N_12708,N_11749,N_11432);
nor U12709 (N_12709,N_11715,N_11971);
nor U12710 (N_12710,N_11633,N_11466);
or U12711 (N_12711,N_11199,N_11713);
xnor U12712 (N_12712,N_11573,N_11331);
and U12713 (N_12713,N_11609,N_11456);
or U12714 (N_12714,N_11493,N_11500);
and U12715 (N_12715,N_11571,N_11043);
and U12716 (N_12716,N_11773,N_11116);
nand U12717 (N_12717,N_11774,N_11811);
or U12718 (N_12718,N_11566,N_11958);
nor U12719 (N_12719,N_11298,N_11733);
nand U12720 (N_12720,N_11703,N_11177);
nor U12721 (N_12721,N_11377,N_11529);
or U12722 (N_12722,N_11999,N_11607);
and U12723 (N_12723,N_11817,N_11919);
xor U12724 (N_12724,N_11142,N_11815);
nor U12725 (N_12725,N_11789,N_11024);
and U12726 (N_12726,N_11369,N_11729);
or U12727 (N_12727,N_11662,N_11449);
or U12728 (N_12728,N_11101,N_11782);
xor U12729 (N_12729,N_11697,N_11878);
and U12730 (N_12730,N_11189,N_11568);
or U12731 (N_12731,N_11158,N_11456);
and U12732 (N_12732,N_11256,N_11539);
xnor U12733 (N_12733,N_11943,N_11121);
nor U12734 (N_12734,N_11671,N_11025);
and U12735 (N_12735,N_11109,N_11139);
or U12736 (N_12736,N_11053,N_11549);
nor U12737 (N_12737,N_11189,N_11282);
nor U12738 (N_12738,N_11229,N_11486);
xnor U12739 (N_12739,N_11403,N_11452);
or U12740 (N_12740,N_11171,N_11117);
and U12741 (N_12741,N_11711,N_11528);
or U12742 (N_12742,N_11212,N_11703);
or U12743 (N_12743,N_11239,N_11151);
or U12744 (N_12744,N_11859,N_11356);
and U12745 (N_12745,N_11679,N_11389);
xor U12746 (N_12746,N_11960,N_11229);
xnor U12747 (N_12747,N_11310,N_11556);
and U12748 (N_12748,N_11459,N_11847);
nand U12749 (N_12749,N_11725,N_11423);
or U12750 (N_12750,N_11042,N_11630);
nor U12751 (N_12751,N_11065,N_11325);
and U12752 (N_12752,N_11949,N_11399);
xor U12753 (N_12753,N_11336,N_11937);
xor U12754 (N_12754,N_11450,N_11029);
or U12755 (N_12755,N_11470,N_11277);
nand U12756 (N_12756,N_11641,N_11954);
nor U12757 (N_12757,N_11416,N_11972);
and U12758 (N_12758,N_11935,N_11576);
and U12759 (N_12759,N_11393,N_11726);
and U12760 (N_12760,N_11544,N_11752);
nor U12761 (N_12761,N_11908,N_11919);
or U12762 (N_12762,N_11980,N_11771);
and U12763 (N_12763,N_11510,N_11031);
xnor U12764 (N_12764,N_11335,N_11079);
nand U12765 (N_12765,N_11684,N_11934);
nor U12766 (N_12766,N_11384,N_11204);
and U12767 (N_12767,N_11656,N_11664);
or U12768 (N_12768,N_11877,N_11822);
xnor U12769 (N_12769,N_11106,N_11692);
xor U12770 (N_12770,N_11746,N_11884);
or U12771 (N_12771,N_11180,N_11499);
and U12772 (N_12772,N_11560,N_11238);
or U12773 (N_12773,N_11452,N_11194);
or U12774 (N_12774,N_11000,N_11912);
nor U12775 (N_12775,N_11292,N_11208);
xor U12776 (N_12776,N_11744,N_11642);
xor U12777 (N_12777,N_11083,N_11313);
nand U12778 (N_12778,N_11311,N_11849);
xor U12779 (N_12779,N_11201,N_11137);
nand U12780 (N_12780,N_11524,N_11659);
nor U12781 (N_12781,N_11095,N_11172);
nor U12782 (N_12782,N_11111,N_11777);
and U12783 (N_12783,N_11449,N_11718);
xnor U12784 (N_12784,N_11848,N_11881);
nor U12785 (N_12785,N_11178,N_11073);
nand U12786 (N_12786,N_11862,N_11067);
nor U12787 (N_12787,N_11808,N_11969);
and U12788 (N_12788,N_11673,N_11133);
or U12789 (N_12789,N_11905,N_11496);
xor U12790 (N_12790,N_11228,N_11670);
or U12791 (N_12791,N_11474,N_11650);
xor U12792 (N_12792,N_11055,N_11987);
xnor U12793 (N_12793,N_11503,N_11751);
or U12794 (N_12794,N_11710,N_11542);
nand U12795 (N_12795,N_11627,N_11013);
xnor U12796 (N_12796,N_11029,N_11203);
or U12797 (N_12797,N_11909,N_11178);
nor U12798 (N_12798,N_11381,N_11652);
or U12799 (N_12799,N_11331,N_11414);
and U12800 (N_12800,N_11290,N_11923);
nand U12801 (N_12801,N_11022,N_11635);
or U12802 (N_12802,N_11297,N_11690);
and U12803 (N_12803,N_11226,N_11870);
nor U12804 (N_12804,N_11920,N_11965);
xor U12805 (N_12805,N_11061,N_11378);
nor U12806 (N_12806,N_11368,N_11828);
nand U12807 (N_12807,N_11777,N_11326);
xor U12808 (N_12808,N_11746,N_11953);
nor U12809 (N_12809,N_11510,N_11698);
nand U12810 (N_12810,N_11083,N_11059);
nor U12811 (N_12811,N_11595,N_11213);
nand U12812 (N_12812,N_11876,N_11866);
and U12813 (N_12813,N_11783,N_11885);
xnor U12814 (N_12814,N_11102,N_11268);
nor U12815 (N_12815,N_11337,N_11044);
or U12816 (N_12816,N_11588,N_11063);
nand U12817 (N_12817,N_11618,N_11076);
xnor U12818 (N_12818,N_11532,N_11786);
xor U12819 (N_12819,N_11272,N_11081);
and U12820 (N_12820,N_11164,N_11119);
xnor U12821 (N_12821,N_11241,N_11755);
or U12822 (N_12822,N_11087,N_11536);
nor U12823 (N_12823,N_11474,N_11584);
and U12824 (N_12824,N_11782,N_11931);
or U12825 (N_12825,N_11977,N_11031);
nand U12826 (N_12826,N_11934,N_11505);
or U12827 (N_12827,N_11992,N_11216);
or U12828 (N_12828,N_11153,N_11255);
and U12829 (N_12829,N_11887,N_11644);
nand U12830 (N_12830,N_11314,N_11646);
or U12831 (N_12831,N_11325,N_11427);
nor U12832 (N_12832,N_11964,N_11729);
and U12833 (N_12833,N_11417,N_11451);
or U12834 (N_12834,N_11876,N_11115);
or U12835 (N_12835,N_11513,N_11098);
or U12836 (N_12836,N_11570,N_11914);
and U12837 (N_12837,N_11946,N_11953);
xnor U12838 (N_12838,N_11957,N_11295);
nor U12839 (N_12839,N_11178,N_11976);
xor U12840 (N_12840,N_11355,N_11182);
xor U12841 (N_12841,N_11082,N_11476);
nand U12842 (N_12842,N_11327,N_11287);
xor U12843 (N_12843,N_11552,N_11822);
xor U12844 (N_12844,N_11197,N_11266);
nand U12845 (N_12845,N_11363,N_11867);
or U12846 (N_12846,N_11895,N_11181);
xnor U12847 (N_12847,N_11909,N_11802);
nor U12848 (N_12848,N_11173,N_11395);
nor U12849 (N_12849,N_11902,N_11811);
and U12850 (N_12850,N_11343,N_11761);
xor U12851 (N_12851,N_11381,N_11267);
and U12852 (N_12852,N_11257,N_11183);
nor U12853 (N_12853,N_11968,N_11137);
nor U12854 (N_12854,N_11506,N_11483);
xnor U12855 (N_12855,N_11784,N_11513);
nor U12856 (N_12856,N_11779,N_11157);
or U12857 (N_12857,N_11992,N_11999);
nor U12858 (N_12858,N_11652,N_11584);
nand U12859 (N_12859,N_11234,N_11152);
nor U12860 (N_12860,N_11625,N_11284);
nor U12861 (N_12861,N_11471,N_11840);
xor U12862 (N_12862,N_11322,N_11755);
nor U12863 (N_12863,N_11083,N_11632);
nor U12864 (N_12864,N_11469,N_11507);
nor U12865 (N_12865,N_11893,N_11190);
or U12866 (N_12866,N_11528,N_11082);
nor U12867 (N_12867,N_11465,N_11604);
xnor U12868 (N_12868,N_11410,N_11390);
and U12869 (N_12869,N_11377,N_11960);
nor U12870 (N_12870,N_11864,N_11179);
xor U12871 (N_12871,N_11131,N_11431);
and U12872 (N_12872,N_11266,N_11645);
nand U12873 (N_12873,N_11872,N_11983);
nand U12874 (N_12874,N_11965,N_11119);
or U12875 (N_12875,N_11081,N_11380);
nor U12876 (N_12876,N_11182,N_11209);
nor U12877 (N_12877,N_11419,N_11766);
nand U12878 (N_12878,N_11627,N_11891);
xor U12879 (N_12879,N_11906,N_11644);
nor U12880 (N_12880,N_11177,N_11240);
and U12881 (N_12881,N_11732,N_11512);
and U12882 (N_12882,N_11115,N_11420);
and U12883 (N_12883,N_11915,N_11540);
nor U12884 (N_12884,N_11634,N_11274);
or U12885 (N_12885,N_11629,N_11920);
and U12886 (N_12886,N_11193,N_11405);
nand U12887 (N_12887,N_11969,N_11587);
xor U12888 (N_12888,N_11678,N_11969);
nand U12889 (N_12889,N_11446,N_11595);
and U12890 (N_12890,N_11041,N_11069);
and U12891 (N_12891,N_11773,N_11403);
xnor U12892 (N_12892,N_11739,N_11549);
or U12893 (N_12893,N_11187,N_11064);
nor U12894 (N_12894,N_11017,N_11113);
xnor U12895 (N_12895,N_11547,N_11197);
nand U12896 (N_12896,N_11932,N_11285);
xor U12897 (N_12897,N_11532,N_11487);
or U12898 (N_12898,N_11579,N_11744);
and U12899 (N_12899,N_11501,N_11580);
or U12900 (N_12900,N_11685,N_11668);
or U12901 (N_12901,N_11123,N_11004);
nor U12902 (N_12902,N_11579,N_11839);
nand U12903 (N_12903,N_11487,N_11251);
xnor U12904 (N_12904,N_11748,N_11571);
xnor U12905 (N_12905,N_11586,N_11636);
xnor U12906 (N_12906,N_11860,N_11619);
xnor U12907 (N_12907,N_11158,N_11832);
xor U12908 (N_12908,N_11325,N_11254);
xor U12909 (N_12909,N_11688,N_11082);
xnor U12910 (N_12910,N_11258,N_11309);
or U12911 (N_12911,N_11430,N_11198);
nor U12912 (N_12912,N_11312,N_11535);
nand U12913 (N_12913,N_11092,N_11467);
and U12914 (N_12914,N_11270,N_11590);
nand U12915 (N_12915,N_11122,N_11264);
nor U12916 (N_12916,N_11688,N_11920);
and U12917 (N_12917,N_11656,N_11960);
nand U12918 (N_12918,N_11936,N_11782);
nor U12919 (N_12919,N_11565,N_11510);
and U12920 (N_12920,N_11961,N_11607);
or U12921 (N_12921,N_11340,N_11342);
xor U12922 (N_12922,N_11178,N_11671);
or U12923 (N_12923,N_11763,N_11715);
nor U12924 (N_12924,N_11036,N_11905);
or U12925 (N_12925,N_11864,N_11576);
nor U12926 (N_12926,N_11148,N_11126);
xnor U12927 (N_12927,N_11820,N_11198);
nor U12928 (N_12928,N_11654,N_11333);
nor U12929 (N_12929,N_11236,N_11923);
nand U12930 (N_12930,N_11842,N_11027);
nand U12931 (N_12931,N_11403,N_11192);
or U12932 (N_12932,N_11385,N_11103);
xor U12933 (N_12933,N_11014,N_11159);
xnor U12934 (N_12934,N_11027,N_11769);
and U12935 (N_12935,N_11461,N_11271);
xnor U12936 (N_12936,N_11142,N_11983);
and U12937 (N_12937,N_11251,N_11976);
and U12938 (N_12938,N_11659,N_11624);
and U12939 (N_12939,N_11436,N_11586);
or U12940 (N_12940,N_11956,N_11070);
nand U12941 (N_12941,N_11643,N_11953);
xnor U12942 (N_12942,N_11737,N_11345);
and U12943 (N_12943,N_11580,N_11346);
xnor U12944 (N_12944,N_11475,N_11202);
nor U12945 (N_12945,N_11385,N_11723);
nor U12946 (N_12946,N_11649,N_11212);
nor U12947 (N_12947,N_11651,N_11418);
and U12948 (N_12948,N_11418,N_11419);
xor U12949 (N_12949,N_11658,N_11578);
nand U12950 (N_12950,N_11267,N_11128);
xor U12951 (N_12951,N_11213,N_11813);
or U12952 (N_12952,N_11949,N_11524);
nand U12953 (N_12953,N_11371,N_11974);
nand U12954 (N_12954,N_11783,N_11349);
xnor U12955 (N_12955,N_11702,N_11663);
or U12956 (N_12956,N_11118,N_11181);
and U12957 (N_12957,N_11886,N_11824);
or U12958 (N_12958,N_11496,N_11812);
nand U12959 (N_12959,N_11694,N_11822);
and U12960 (N_12960,N_11548,N_11845);
and U12961 (N_12961,N_11894,N_11978);
nor U12962 (N_12962,N_11453,N_11741);
xnor U12963 (N_12963,N_11832,N_11074);
and U12964 (N_12964,N_11311,N_11530);
nand U12965 (N_12965,N_11997,N_11975);
xor U12966 (N_12966,N_11652,N_11970);
xnor U12967 (N_12967,N_11905,N_11610);
and U12968 (N_12968,N_11423,N_11617);
or U12969 (N_12969,N_11595,N_11660);
and U12970 (N_12970,N_11460,N_11107);
xnor U12971 (N_12971,N_11768,N_11782);
nand U12972 (N_12972,N_11748,N_11249);
nor U12973 (N_12973,N_11039,N_11602);
or U12974 (N_12974,N_11043,N_11903);
nand U12975 (N_12975,N_11004,N_11233);
xnor U12976 (N_12976,N_11437,N_11837);
or U12977 (N_12977,N_11962,N_11162);
xnor U12978 (N_12978,N_11157,N_11942);
xor U12979 (N_12979,N_11510,N_11397);
or U12980 (N_12980,N_11005,N_11676);
nor U12981 (N_12981,N_11692,N_11803);
nor U12982 (N_12982,N_11517,N_11756);
and U12983 (N_12983,N_11117,N_11822);
xor U12984 (N_12984,N_11945,N_11402);
and U12985 (N_12985,N_11178,N_11517);
xor U12986 (N_12986,N_11835,N_11041);
nor U12987 (N_12987,N_11680,N_11265);
and U12988 (N_12988,N_11688,N_11652);
or U12989 (N_12989,N_11148,N_11543);
nor U12990 (N_12990,N_11169,N_11770);
nand U12991 (N_12991,N_11892,N_11040);
nand U12992 (N_12992,N_11826,N_11119);
nand U12993 (N_12993,N_11772,N_11536);
xor U12994 (N_12994,N_11069,N_11215);
nor U12995 (N_12995,N_11189,N_11102);
or U12996 (N_12996,N_11622,N_11200);
nor U12997 (N_12997,N_11603,N_11849);
xor U12998 (N_12998,N_11149,N_11336);
and U12999 (N_12999,N_11016,N_11025);
xnor U13000 (N_13000,N_12325,N_12838);
nor U13001 (N_13001,N_12001,N_12361);
nor U13002 (N_13002,N_12317,N_12551);
xnor U13003 (N_13003,N_12622,N_12244);
or U13004 (N_13004,N_12357,N_12349);
or U13005 (N_13005,N_12151,N_12256);
and U13006 (N_13006,N_12889,N_12826);
xor U13007 (N_13007,N_12105,N_12042);
or U13008 (N_13008,N_12350,N_12293);
nor U13009 (N_13009,N_12849,N_12626);
nand U13010 (N_13010,N_12434,N_12462);
and U13011 (N_13011,N_12192,N_12786);
and U13012 (N_13012,N_12916,N_12381);
xnor U13013 (N_13013,N_12323,N_12468);
and U13014 (N_13014,N_12821,N_12473);
nand U13015 (N_13015,N_12047,N_12074);
or U13016 (N_13016,N_12301,N_12960);
and U13017 (N_13017,N_12258,N_12517);
or U13018 (N_13018,N_12255,N_12142);
nor U13019 (N_13019,N_12614,N_12606);
xor U13020 (N_13020,N_12744,N_12898);
and U13021 (N_13021,N_12359,N_12145);
or U13022 (N_13022,N_12809,N_12076);
and U13023 (N_13023,N_12979,N_12190);
and U13024 (N_13024,N_12605,N_12287);
nor U13025 (N_13025,N_12629,N_12312);
nor U13026 (N_13026,N_12432,N_12833);
nand U13027 (N_13027,N_12014,N_12218);
nor U13028 (N_13028,N_12099,N_12379);
xor U13029 (N_13029,N_12199,N_12087);
or U13030 (N_13030,N_12419,N_12686);
xor U13031 (N_13031,N_12777,N_12949);
nor U13032 (N_13032,N_12391,N_12370);
nand U13033 (N_13033,N_12007,N_12846);
nand U13034 (N_13034,N_12822,N_12522);
xor U13035 (N_13035,N_12543,N_12946);
or U13036 (N_13036,N_12263,N_12827);
xor U13037 (N_13037,N_12496,N_12059);
and U13038 (N_13038,N_12611,N_12439);
or U13039 (N_13039,N_12625,N_12913);
and U13040 (N_13040,N_12431,N_12273);
xor U13041 (N_13041,N_12901,N_12937);
xor U13042 (N_13042,N_12637,N_12238);
nor U13043 (N_13043,N_12499,N_12234);
nor U13044 (N_13044,N_12928,N_12912);
or U13045 (N_13045,N_12168,N_12900);
xor U13046 (N_13046,N_12157,N_12340);
and U13047 (N_13047,N_12289,N_12897);
or U13048 (N_13048,N_12167,N_12117);
nand U13049 (N_13049,N_12482,N_12750);
nor U13050 (N_13050,N_12619,N_12436);
nor U13051 (N_13051,N_12682,N_12505);
xor U13052 (N_13052,N_12139,N_12012);
and U13053 (N_13053,N_12861,N_12915);
nand U13054 (N_13054,N_12048,N_12935);
nand U13055 (N_13055,N_12348,N_12518);
xor U13056 (N_13056,N_12698,N_12885);
xnor U13057 (N_13057,N_12623,N_12977);
nand U13058 (N_13058,N_12343,N_12806);
or U13059 (N_13059,N_12557,N_12058);
nor U13060 (N_13060,N_12534,N_12268);
nor U13061 (N_13061,N_12683,N_12320);
nand U13062 (N_13062,N_12975,N_12033);
nor U13063 (N_13063,N_12636,N_12847);
xnor U13064 (N_13064,N_12600,N_12504);
and U13065 (N_13065,N_12651,N_12372);
or U13066 (N_13066,N_12337,N_12174);
nor U13067 (N_13067,N_12415,N_12133);
nor U13068 (N_13068,N_12607,N_12329);
xor U13069 (N_13069,N_12477,N_12851);
xor U13070 (N_13070,N_12333,N_12364);
or U13071 (N_13071,N_12789,N_12144);
nor U13072 (N_13072,N_12107,N_12314);
or U13073 (N_13073,N_12132,N_12004);
xor U13074 (N_13074,N_12705,N_12741);
and U13075 (N_13075,N_12709,N_12321);
and U13076 (N_13076,N_12120,N_12036);
xnor U13077 (N_13077,N_12267,N_12377);
and U13078 (N_13078,N_12580,N_12961);
nor U13079 (N_13079,N_12627,N_12862);
and U13080 (N_13080,N_12128,N_12638);
xnor U13081 (N_13081,N_12888,N_12194);
nor U13082 (N_13082,N_12875,N_12338);
and U13083 (N_13083,N_12054,N_12112);
nor U13084 (N_13084,N_12771,N_12429);
nand U13085 (N_13085,N_12701,N_12583);
nor U13086 (N_13086,N_12540,N_12009);
or U13087 (N_13087,N_12443,N_12383);
or U13088 (N_13088,N_12963,N_12448);
and U13089 (N_13089,N_12511,N_12308);
nor U13090 (N_13090,N_12713,N_12173);
nor U13091 (N_13091,N_12630,N_12566);
xor U13092 (N_13092,N_12965,N_12652);
nand U13093 (N_13093,N_12088,N_12553);
nand U13094 (N_13094,N_12365,N_12689);
or U13095 (N_13095,N_12109,N_12290);
and U13096 (N_13096,N_12219,N_12914);
nor U13097 (N_13097,N_12990,N_12992);
and U13098 (N_13098,N_12988,N_12274);
or U13099 (N_13099,N_12746,N_12114);
or U13100 (N_13100,N_12776,N_12177);
nand U13101 (N_13101,N_12634,N_12596);
and U13102 (N_13102,N_12426,N_12828);
nor U13103 (N_13103,N_12420,N_12457);
nand U13104 (N_13104,N_12989,N_12332);
nand U13105 (N_13105,N_12648,N_12351);
nand U13106 (N_13106,N_12119,N_12011);
nor U13107 (N_13107,N_12208,N_12510);
and U13108 (N_13108,N_12090,N_12401);
and U13109 (N_13109,N_12345,N_12834);
nor U13110 (N_13110,N_12936,N_12277);
nor U13111 (N_13111,N_12118,N_12322);
or U13112 (N_13112,N_12529,N_12156);
and U13113 (N_13113,N_12533,N_12342);
and U13114 (N_13114,N_12164,N_12572);
nor U13115 (N_13115,N_12845,N_12696);
xnor U13116 (N_13116,N_12220,N_12772);
and U13117 (N_13117,N_12062,N_12037);
nand U13118 (N_13118,N_12295,N_12631);
or U13119 (N_13119,N_12418,N_12183);
nand U13120 (N_13120,N_12288,N_12104);
or U13121 (N_13121,N_12876,N_12502);
or U13122 (N_13122,N_12095,N_12739);
nor U13123 (N_13123,N_12163,N_12933);
xnor U13124 (N_13124,N_12591,N_12298);
nand U13125 (N_13125,N_12802,N_12438);
or U13126 (N_13126,N_12593,N_12760);
xnor U13127 (N_13127,N_12675,N_12201);
nor U13128 (N_13128,N_12672,N_12556);
and U13129 (N_13129,N_12236,N_12545);
nor U13130 (N_13130,N_12956,N_12911);
or U13131 (N_13131,N_12718,N_12666);
xnor U13132 (N_13132,N_12774,N_12013);
nand U13133 (N_13133,N_12769,N_12451);
xnor U13134 (N_13134,N_12252,N_12563);
or U13135 (N_13135,N_12228,N_12405);
nand U13136 (N_13136,N_12560,N_12554);
nor U13137 (N_13137,N_12832,N_12435);
and U13138 (N_13138,N_12998,N_12697);
or U13139 (N_13139,N_12526,N_12159);
nor U13140 (N_13140,N_12335,N_12603);
nand U13141 (N_13141,N_12538,N_12138);
nor U13142 (N_13142,N_12407,N_12953);
nand U13143 (N_13143,N_12646,N_12945);
nor U13144 (N_13144,N_12052,N_12130);
xnor U13145 (N_13145,N_12733,N_12680);
nor U13146 (N_13146,N_12261,N_12586);
and U13147 (N_13147,N_12035,N_12209);
xor U13148 (N_13148,N_12836,N_12818);
nand U13149 (N_13149,N_12757,N_12131);
nand U13150 (N_13150,N_12224,N_12588);
nor U13151 (N_13151,N_12985,N_12300);
or U13152 (N_13152,N_12470,N_12654);
nand U13153 (N_13153,N_12795,N_12642);
nor U13154 (N_13154,N_12486,N_12070);
xnor U13155 (N_13155,N_12053,N_12100);
xnor U13156 (N_13156,N_12171,N_12893);
xor U13157 (N_13157,N_12981,N_12356);
xnor U13158 (N_13158,N_12574,N_12924);
and U13159 (N_13159,N_12728,N_12221);
and U13160 (N_13160,N_12223,N_12678);
nand U13161 (N_13161,N_12269,N_12137);
or U13162 (N_13162,N_12284,N_12479);
xnor U13163 (N_13163,N_12200,N_12445);
xnor U13164 (N_13164,N_12080,N_12724);
xor U13165 (N_13165,N_12811,N_12115);
nor U13166 (N_13166,N_12483,N_12206);
xnor U13167 (N_13167,N_12464,N_12480);
and U13168 (N_13168,N_12250,N_12038);
nand U13169 (N_13169,N_12110,N_12794);
and U13170 (N_13170,N_12213,N_12970);
nor U13171 (N_13171,N_12286,N_12463);
nor U13172 (N_13172,N_12406,N_12918);
or U13173 (N_13173,N_12531,N_12010);
or U13174 (N_13174,N_12549,N_12031);
and U13175 (N_13175,N_12082,N_12920);
nand U13176 (N_13176,N_12957,N_12424);
or U13177 (N_13177,N_12804,N_12028);
and U13178 (N_13178,N_12919,N_12925);
nor U13179 (N_13179,N_12140,N_12576);
nand U13180 (N_13180,N_12067,N_12797);
nor U13181 (N_13181,N_12866,N_12461);
nor U13182 (N_13182,N_12389,N_12362);
nor U13183 (N_13183,N_12066,N_12101);
xnor U13184 (N_13184,N_12245,N_12046);
xor U13185 (N_13185,N_12315,N_12952);
nor U13186 (N_13186,N_12753,N_12185);
or U13187 (N_13187,N_12527,N_12495);
xor U13188 (N_13188,N_12968,N_12181);
nor U13189 (N_13189,N_12465,N_12707);
nor U13190 (N_13190,N_12581,N_12254);
nor U13191 (N_13191,N_12454,N_12061);
xnor U13192 (N_13192,N_12870,N_12964);
nor U13193 (N_13193,N_12881,N_12906);
and U13194 (N_13194,N_12650,N_12535);
xor U13195 (N_13195,N_12143,N_12410);
xor U13196 (N_13196,N_12197,N_12512);
xnor U13197 (N_13197,N_12703,N_12417);
and U13198 (N_13198,N_12060,N_12708);
and U13199 (N_13199,N_12765,N_12693);
and U13200 (N_13200,N_12839,N_12716);
xnor U13201 (N_13201,N_12587,N_12318);
or U13202 (N_13202,N_12500,N_12073);
and U13203 (N_13203,N_12819,N_12747);
and U13204 (N_13204,N_12027,N_12779);
and U13205 (N_13205,N_12063,N_12570);
or U13206 (N_13206,N_12302,N_12879);
and U13207 (N_13207,N_12691,N_12649);
or U13208 (N_13208,N_12247,N_12720);
nand U13209 (N_13209,N_12083,N_12153);
nor U13210 (N_13210,N_12316,N_12376);
xnor U13211 (N_13211,N_12475,N_12170);
nand U13212 (N_13212,N_12489,N_12515);
xnor U13213 (N_13213,N_12229,N_12695);
nand U13214 (N_13214,N_12278,N_12514);
xor U13215 (N_13215,N_12902,N_12240);
nand U13216 (N_13216,N_12699,N_12241);
nor U13217 (N_13217,N_12018,N_12559);
xor U13218 (N_13218,N_12840,N_12816);
or U13219 (N_13219,N_12950,N_12266);
nor U13220 (N_13220,N_12971,N_12459);
or U13221 (N_13221,N_12021,N_12657);
or U13222 (N_13222,N_12715,N_12437);
xor U13223 (N_13223,N_12210,N_12422);
and U13224 (N_13224,N_12395,N_12392);
nor U13225 (N_13225,N_12193,N_12442);
nand U13226 (N_13226,N_12921,N_12509);
or U13227 (N_13227,N_12768,N_12353);
and U13228 (N_13228,N_12032,N_12877);
or U13229 (N_13229,N_12141,N_12341);
or U13230 (N_13230,N_12694,N_12265);
or U13231 (N_13231,N_12413,N_12837);
or U13232 (N_13232,N_12668,N_12270);
and U13233 (N_13233,N_12959,N_12677);
xor U13234 (N_13234,N_12766,N_12661);
or U13235 (N_13235,N_12366,N_12815);
or U13236 (N_13236,N_12858,N_12447);
nor U13237 (N_13237,N_12049,N_12859);
or U13238 (N_13238,N_12742,N_12719);
nor U13239 (N_13239,N_12860,N_12191);
xor U13240 (N_13240,N_12934,N_12974);
and U13241 (N_13241,N_12874,N_12712);
or U13242 (N_13242,N_12150,N_12326);
nor U13243 (N_13243,N_12730,N_12179);
xor U13244 (N_13244,N_12855,N_12040);
nor U13245 (N_13245,N_12700,N_12425);
and U13246 (N_13246,N_12122,N_12980);
nand U13247 (N_13247,N_12612,N_12121);
xnor U13248 (N_13248,N_12072,N_12068);
and U13249 (N_13249,N_12490,N_12520);
or U13250 (N_13250,N_12230,N_12260);
xor U13251 (N_13251,N_12441,N_12761);
nand U13252 (N_13252,N_12116,N_12178);
and U13253 (N_13253,N_12643,N_12759);
nor U13254 (N_13254,N_12525,N_12123);
nor U13255 (N_13255,N_12983,N_12079);
nor U13256 (N_13256,N_12069,N_12064);
xnor U13257 (N_13257,N_12334,N_12610);
and U13258 (N_13258,N_12564,N_12613);
nor U13259 (N_13259,N_12594,N_12878);
xor U13260 (N_13260,N_12214,N_12633);
and U13261 (N_13261,N_12235,N_12883);
or U13262 (N_13262,N_12727,N_12667);
nor U13263 (N_13263,N_12722,N_12714);
xor U13264 (N_13264,N_12360,N_12571);
xnor U13265 (N_13265,N_12938,N_12884);
and U13266 (N_13266,N_12873,N_12324);
nor U13267 (N_13267,N_12573,N_12427);
nand U13268 (N_13268,N_12910,N_12831);
nand U13269 (N_13269,N_12215,N_12148);
nand U13270 (N_13270,N_12050,N_12530);
nand U13271 (N_13271,N_12374,N_12103);
or U13272 (N_13272,N_12737,N_12669);
and U13273 (N_13273,N_12907,N_12947);
nor U13274 (N_13274,N_12015,N_12008);
nand U13275 (N_13275,N_12762,N_12909);
or U13276 (N_13276,N_12400,N_12239);
and U13277 (N_13277,N_12841,N_12196);
xor U13278 (N_13278,N_12598,N_12558);
and U13279 (N_13279,N_12555,N_12226);
and U13280 (N_13280,N_12966,N_12257);
xnor U13281 (N_13281,N_12781,N_12955);
nor U13282 (N_13282,N_12787,N_12835);
or U13283 (N_13283,N_12280,N_12702);
and U13284 (N_13284,N_12125,N_12368);
and U13285 (N_13285,N_12721,N_12620);
or U13286 (N_13286,N_12908,N_12641);
or U13287 (N_13287,N_12481,N_12615);
nor U13288 (N_13288,N_12519,N_12084);
nor U13289 (N_13289,N_12198,N_12516);
nand U13290 (N_13290,N_12756,N_12045);
or U13291 (N_13291,N_12217,N_12154);
nor U13292 (N_13292,N_12378,N_12820);
nand U13293 (N_13293,N_12299,N_12801);
xnor U13294 (N_13294,N_12679,N_12710);
nand U13295 (N_13295,N_12182,N_12246);
xor U13296 (N_13296,N_12446,N_12891);
or U13297 (N_13297,N_12390,N_12513);
nand U13298 (N_13298,N_12987,N_12404);
or U13299 (N_13299,N_12307,N_12222);
xor U13300 (N_13300,N_12396,N_12205);
xnor U13301 (N_13301,N_12582,N_12127);
and U13302 (N_13302,N_12954,N_12147);
nand U13303 (N_13303,N_12124,N_12285);
nor U13304 (N_13304,N_12149,N_12291);
or U13305 (N_13305,N_12005,N_12793);
xor U13306 (N_13306,N_12671,N_12386);
nand U13307 (N_13307,N_12880,N_12327);
nand U13308 (N_13308,N_12186,N_12997);
or U13309 (N_13309,N_12621,N_12567);
and U13310 (N_13310,N_12398,N_12373);
or U13311 (N_13311,N_12561,N_12972);
nand U13312 (N_13312,N_12503,N_12547);
and U13313 (N_13313,N_12394,N_12414);
nand U13314 (N_13314,N_12958,N_12764);
and U13315 (N_13315,N_12172,N_12995);
and U13316 (N_13316,N_12725,N_12352);
xnor U13317 (N_13317,N_12294,N_12108);
or U13318 (N_13318,N_12842,N_12225);
nand U13319 (N_13319,N_12097,N_12532);
and U13320 (N_13320,N_12940,N_12111);
and U13321 (N_13321,N_12175,N_12180);
nand U13322 (N_13322,N_12026,N_12830);
nor U13323 (N_13323,N_12262,N_12281);
nand U13324 (N_13324,N_12303,N_12922);
nand U13325 (N_13325,N_12930,N_12590);
xor U13326 (N_13326,N_12458,N_12189);
nand U13327 (N_13327,N_12941,N_12617);
nand U13328 (N_13328,N_12749,N_12663);
xnor U13329 (N_13329,N_12681,N_12272);
nand U13330 (N_13330,N_12863,N_12803);
or U13331 (N_13331,N_12313,N_12670);
nor U13332 (N_13332,N_12020,N_12569);
or U13333 (N_13333,N_12871,N_12639);
xnor U13334 (N_13334,N_12729,N_12339);
or U13335 (N_13335,N_12055,N_12207);
nand U13336 (N_13336,N_12864,N_12973);
nand U13337 (N_13337,N_12812,N_12169);
and U13338 (N_13338,N_12492,N_12310);
and U13339 (N_13339,N_12024,N_12655);
and U13340 (N_13340,N_12264,N_12904);
and U13341 (N_13341,N_12093,N_12754);
xor U13342 (N_13342,N_12599,N_12537);
and U13343 (N_13343,N_12982,N_12685);
nor U13344 (N_13344,N_12051,N_12501);
xor U13345 (N_13345,N_12896,N_12094);
and U13346 (N_13346,N_12917,N_12471);
or U13347 (N_13347,N_12166,N_12640);
nand U13348 (N_13348,N_12408,N_12523);
or U13349 (N_13349,N_12609,N_12986);
nand U13350 (N_13350,N_12616,N_12375);
and U13351 (N_13351,N_12152,N_12430);
and U13352 (N_13352,N_12271,N_12507);
xnor U13353 (N_13353,N_12203,N_12212);
nor U13354 (N_13354,N_12472,N_12296);
nor U13355 (N_13355,N_12738,N_12991);
nand U13356 (N_13356,N_12813,N_12387);
nor U13357 (N_13357,N_12624,N_12363);
or U13358 (N_13358,N_12791,N_12589);
xor U13359 (N_13359,N_12155,N_12943);
nor U13360 (N_13360,N_12452,N_12780);
and U13361 (N_13361,N_12692,N_12211);
nand U13362 (N_13362,N_12595,N_12380);
nand U13363 (N_13363,N_12790,N_12176);
or U13364 (N_13364,N_12478,N_12854);
nand U13365 (N_13365,N_12202,N_12184);
nor U13366 (N_13366,N_12098,N_12276);
nor U13367 (N_13367,N_12544,N_12647);
nand U13368 (N_13368,N_12002,N_12926);
xnor U13369 (N_13369,N_12796,N_12330);
nand U13370 (N_13370,N_12204,N_12449);
and U13371 (N_13371,N_12003,N_12644);
or U13372 (N_13372,N_12493,N_12135);
nand U13373 (N_13373,N_12767,N_12216);
nand U13374 (N_13374,N_12065,N_12344);
nand U13375 (N_13375,N_12126,N_12231);
nand U13376 (N_13376,N_12485,N_12597);
or U13377 (N_13377,N_12041,N_12824);
nor U13378 (N_13378,N_12081,N_12242);
nand U13379 (N_13379,N_12688,N_12160);
nor U13380 (N_13380,N_12528,N_12808);
or U13381 (N_13381,N_12550,N_12487);
nand U13382 (N_13382,N_12592,N_12232);
nor U13383 (N_13383,N_12484,N_12248);
nand U13384 (N_13384,N_12962,N_12102);
xnor U13385 (N_13385,N_12942,N_12731);
nand U13386 (N_13386,N_12664,N_12660);
or U13387 (N_13387,N_12734,N_12195);
xnor U13388 (N_13388,N_12541,N_12034);
and U13389 (N_13389,N_12732,N_12469);
and U13390 (N_13390,N_12019,N_12129);
or U13391 (N_13391,N_12783,N_12676);
or U13392 (N_13392,N_12999,N_12539);
xnor U13393 (N_13393,N_12399,N_12456);
nand U13394 (N_13394,N_12662,N_12984);
nor U13395 (N_13395,N_12711,N_12106);
nor U13396 (N_13396,N_12440,N_12233);
xnor U13397 (N_13397,N_12450,N_12899);
and U13398 (N_13398,N_12187,N_12792);
xor U13399 (N_13399,N_12939,N_12453);
nand U13400 (N_13400,N_12086,N_12577);
nor U13401 (N_13401,N_12706,N_12726);
xor U13402 (N_13402,N_12077,N_12388);
nor U13403 (N_13403,N_12872,N_12944);
nand U13404 (N_13404,N_12402,N_12306);
and U13405 (N_13405,N_12474,N_12367);
xor U13406 (N_13406,N_12844,N_12565);
and U13407 (N_13407,N_12673,N_12584);
and U13408 (N_13408,N_12575,N_12023);
xor U13409 (N_13409,N_12823,N_12096);
nand U13410 (N_13410,N_12134,N_12085);
nor U13411 (N_13411,N_12506,N_12409);
or U13412 (N_13412,N_12929,N_12976);
nand U13413 (N_13413,N_12347,N_12385);
nand U13414 (N_13414,N_12025,N_12868);
and U13415 (N_13415,N_12319,N_12931);
xor U13416 (N_13416,N_12358,N_12416);
nor U13417 (N_13417,N_12817,N_12146);
or U13418 (N_13418,N_12328,N_12632);
and U13419 (N_13419,N_12788,N_12850);
xnor U13420 (N_13420,N_12006,N_12403);
or U13421 (N_13421,N_12887,N_12044);
and U13422 (N_13422,N_12782,N_12656);
nand U13423 (N_13423,N_12016,N_12755);
and U13424 (N_13424,N_12770,N_12336);
nand U13425 (N_13425,N_12071,N_12775);
nor U13426 (N_13426,N_12078,N_12165);
and U13427 (N_13427,N_12807,N_12022);
nand U13428 (N_13428,N_12092,N_12346);
or U13429 (N_13429,N_12029,N_12508);
xor U13430 (N_13430,N_12932,N_12743);
xnor U13431 (N_13431,N_12785,N_12354);
and U13432 (N_13432,N_12665,N_12740);
nor U13433 (N_13433,N_12243,N_12444);
or U13434 (N_13434,N_12865,N_12498);
nor U13435 (N_13435,N_12886,N_12903);
or U13436 (N_13436,N_12996,N_12089);
nand U13437 (N_13437,N_12136,N_12905);
nor U13438 (N_13438,N_12735,N_12039);
or U13439 (N_13439,N_12536,N_12188);
or U13440 (N_13440,N_12856,N_12382);
xnor U13441 (N_13441,N_12857,N_12867);
or U13442 (N_13442,N_12653,N_12494);
xnor U13443 (N_13443,N_12421,N_12784);
and U13444 (N_13444,N_12455,N_12690);
xnor U13445 (N_13445,N_12162,N_12253);
nand U13446 (N_13446,N_12674,N_12292);
xor U13447 (N_13447,N_12978,N_12562);
nand U13448 (N_13448,N_12057,N_12635);
or U13449 (N_13449,N_12311,N_12763);
or U13450 (N_13450,N_12227,N_12282);
xor U13451 (N_13451,N_12748,N_12491);
xnor U13452 (N_13452,N_12800,N_12412);
nand U13453 (N_13453,N_12704,N_12948);
nor U13454 (N_13454,N_12773,N_12923);
and U13455 (N_13455,N_12994,N_12736);
and U13456 (N_13456,N_12161,N_12546);
nor U13457 (N_13457,N_12810,N_12259);
xnor U13458 (N_13458,N_12853,N_12604);
nand U13459 (N_13459,N_12542,N_12331);
nand U13460 (N_13460,N_12758,N_12869);
xor U13461 (N_13461,N_12384,N_12601);
nor U13462 (N_13462,N_12428,N_12467);
xnor U13463 (N_13463,N_12927,N_12397);
xnor U13464 (N_13464,N_12814,N_12552);
or U13465 (N_13465,N_12895,N_12602);
and U13466 (N_13466,N_12618,N_12752);
nand U13467 (N_13467,N_12805,N_12890);
nand U13468 (N_13468,N_12158,N_12305);
nor U13469 (N_13469,N_12488,N_12275);
nand U13470 (N_13470,N_12659,N_12466);
nor U13471 (N_13471,N_12309,N_12825);
or U13472 (N_13472,N_12283,N_12433);
and U13473 (N_13473,N_12371,N_12017);
or U13474 (N_13474,N_12951,N_12113);
and U13475 (N_13475,N_12279,N_12843);
xnor U13476 (N_13476,N_12524,N_12237);
nor U13477 (N_13477,N_12497,N_12369);
nand U13478 (N_13478,N_12969,N_12628);
nand U13479 (N_13479,N_12075,N_12799);
xor U13480 (N_13480,N_12355,N_12829);
nand U13481 (N_13481,N_12894,N_12251);
nor U13482 (N_13482,N_12030,N_12578);
xnor U13483 (N_13483,N_12423,N_12411);
and U13484 (N_13484,N_12579,N_12717);
xor U13485 (N_13485,N_12684,N_12297);
nand U13486 (N_13486,N_12043,N_12852);
or U13487 (N_13487,N_12521,N_12476);
and U13488 (N_13488,N_12882,N_12548);
nand U13489 (N_13489,N_12993,N_12249);
nor U13490 (N_13490,N_12723,N_12393);
nor U13491 (N_13491,N_12687,N_12967);
or U13492 (N_13492,N_12751,N_12568);
or U13493 (N_13493,N_12658,N_12056);
and U13494 (N_13494,N_12585,N_12608);
xnor U13495 (N_13495,N_12778,N_12645);
nor U13496 (N_13496,N_12798,N_12848);
and U13497 (N_13497,N_12000,N_12460);
or U13498 (N_13498,N_12091,N_12304);
and U13499 (N_13499,N_12745,N_12892);
or U13500 (N_13500,N_12662,N_12317);
and U13501 (N_13501,N_12335,N_12970);
and U13502 (N_13502,N_12409,N_12120);
xor U13503 (N_13503,N_12194,N_12930);
nand U13504 (N_13504,N_12587,N_12636);
and U13505 (N_13505,N_12088,N_12783);
nor U13506 (N_13506,N_12177,N_12742);
or U13507 (N_13507,N_12810,N_12296);
xnor U13508 (N_13508,N_12307,N_12681);
nand U13509 (N_13509,N_12004,N_12854);
nor U13510 (N_13510,N_12972,N_12119);
nor U13511 (N_13511,N_12823,N_12365);
nand U13512 (N_13512,N_12348,N_12100);
xnor U13513 (N_13513,N_12414,N_12399);
xnor U13514 (N_13514,N_12705,N_12531);
xnor U13515 (N_13515,N_12488,N_12209);
nand U13516 (N_13516,N_12910,N_12266);
or U13517 (N_13517,N_12411,N_12819);
nor U13518 (N_13518,N_12467,N_12276);
xor U13519 (N_13519,N_12889,N_12253);
xor U13520 (N_13520,N_12024,N_12155);
or U13521 (N_13521,N_12489,N_12360);
nand U13522 (N_13522,N_12459,N_12178);
nor U13523 (N_13523,N_12531,N_12367);
and U13524 (N_13524,N_12525,N_12216);
nand U13525 (N_13525,N_12461,N_12693);
and U13526 (N_13526,N_12841,N_12174);
and U13527 (N_13527,N_12477,N_12906);
nor U13528 (N_13528,N_12591,N_12224);
and U13529 (N_13529,N_12899,N_12192);
and U13530 (N_13530,N_12204,N_12104);
or U13531 (N_13531,N_12294,N_12216);
and U13532 (N_13532,N_12153,N_12545);
or U13533 (N_13533,N_12474,N_12040);
nor U13534 (N_13534,N_12046,N_12306);
and U13535 (N_13535,N_12250,N_12801);
nor U13536 (N_13536,N_12673,N_12860);
and U13537 (N_13537,N_12229,N_12771);
nor U13538 (N_13538,N_12752,N_12942);
xnor U13539 (N_13539,N_12893,N_12620);
nand U13540 (N_13540,N_12342,N_12853);
nand U13541 (N_13541,N_12305,N_12468);
or U13542 (N_13542,N_12164,N_12931);
nor U13543 (N_13543,N_12793,N_12732);
and U13544 (N_13544,N_12756,N_12594);
nor U13545 (N_13545,N_12361,N_12518);
or U13546 (N_13546,N_12825,N_12677);
nor U13547 (N_13547,N_12348,N_12845);
and U13548 (N_13548,N_12699,N_12198);
xor U13549 (N_13549,N_12654,N_12705);
or U13550 (N_13550,N_12331,N_12480);
nor U13551 (N_13551,N_12216,N_12239);
nand U13552 (N_13552,N_12894,N_12212);
or U13553 (N_13553,N_12574,N_12446);
nand U13554 (N_13554,N_12242,N_12391);
nand U13555 (N_13555,N_12547,N_12976);
xor U13556 (N_13556,N_12448,N_12288);
or U13557 (N_13557,N_12457,N_12479);
nand U13558 (N_13558,N_12970,N_12591);
nor U13559 (N_13559,N_12580,N_12533);
or U13560 (N_13560,N_12919,N_12728);
nor U13561 (N_13561,N_12798,N_12008);
and U13562 (N_13562,N_12411,N_12630);
xor U13563 (N_13563,N_12615,N_12575);
or U13564 (N_13564,N_12960,N_12639);
nor U13565 (N_13565,N_12607,N_12515);
and U13566 (N_13566,N_12473,N_12912);
nor U13567 (N_13567,N_12826,N_12835);
nor U13568 (N_13568,N_12080,N_12307);
and U13569 (N_13569,N_12067,N_12928);
or U13570 (N_13570,N_12546,N_12692);
and U13571 (N_13571,N_12009,N_12056);
or U13572 (N_13572,N_12832,N_12468);
nor U13573 (N_13573,N_12935,N_12110);
nand U13574 (N_13574,N_12504,N_12370);
and U13575 (N_13575,N_12746,N_12555);
nand U13576 (N_13576,N_12566,N_12534);
or U13577 (N_13577,N_12737,N_12501);
xor U13578 (N_13578,N_12194,N_12212);
nor U13579 (N_13579,N_12110,N_12370);
xor U13580 (N_13580,N_12306,N_12332);
nor U13581 (N_13581,N_12353,N_12134);
nor U13582 (N_13582,N_12912,N_12238);
xor U13583 (N_13583,N_12398,N_12555);
xor U13584 (N_13584,N_12717,N_12995);
nand U13585 (N_13585,N_12460,N_12952);
or U13586 (N_13586,N_12113,N_12749);
nand U13587 (N_13587,N_12693,N_12899);
nand U13588 (N_13588,N_12470,N_12989);
nor U13589 (N_13589,N_12393,N_12313);
and U13590 (N_13590,N_12945,N_12702);
xor U13591 (N_13591,N_12105,N_12335);
or U13592 (N_13592,N_12741,N_12098);
and U13593 (N_13593,N_12085,N_12025);
nor U13594 (N_13594,N_12996,N_12780);
nor U13595 (N_13595,N_12671,N_12651);
or U13596 (N_13596,N_12930,N_12326);
nor U13597 (N_13597,N_12024,N_12527);
or U13598 (N_13598,N_12618,N_12952);
nand U13599 (N_13599,N_12126,N_12085);
nor U13600 (N_13600,N_12107,N_12205);
and U13601 (N_13601,N_12523,N_12014);
xor U13602 (N_13602,N_12071,N_12639);
nor U13603 (N_13603,N_12232,N_12358);
or U13604 (N_13604,N_12461,N_12616);
or U13605 (N_13605,N_12787,N_12776);
or U13606 (N_13606,N_12798,N_12088);
nand U13607 (N_13607,N_12324,N_12341);
and U13608 (N_13608,N_12583,N_12824);
nor U13609 (N_13609,N_12357,N_12273);
nor U13610 (N_13610,N_12990,N_12492);
xnor U13611 (N_13611,N_12642,N_12395);
xor U13612 (N_13612,N_12977,N_12394);
nand U13613 (N_13613,N_12667,N_12009);
xnor U13614 (N_13614,N_12352,N_12262);
or U13615 (N_13615,N_12587,N_12723);
and U13616 (N_13616,N_12350,N_12753);
nand U13617 (N_13617,N_12229,N_12735);
xnor U13618 (N_13618,N_12366,N_12432);
and U13619 (N_13619,N_12737,N_12906);
or U13620 (N_13620,N_12305,N_12665);
and U13621 (N_13621,N_12111,N_12958);
nor U13622 (N_13622,N_12780,N_12486);
and U13623 (N_13623,N_12893,N_12754);
or U13624 (N_13624,N_12289,N_12421);
xor U13625 (N_13625,N_12202,N_12278);
xnor U13626 (N_13626,N_12515,N_12762);
nor U13627 (N_13627,N_12897,N_12671);
nand U13628 (N_13628,N_12561,N_12299);
and U13629 (N_13629,N_12595,N_12859);
xor U13630 (N_13630,N_12304,N_12433);
and U13631 (N_13631,N_12547,N_12734);
xnor U13632 (N_13632,N_12574,N_12357);
nor U13633 (N_13633,N_12322,N_12195);
or U13634 (N_13634,N_12770,N_12674);
or U13635 (N_13635,N_12950,N_12056);
nor U13636 (N_13636,N_12929,N_12338);
and U13637 (N_13637,N_12989,N_12416);
nand U13638 (N_13638,N_12817,N_12440);
xor U13639 (N_13639,N_12930,N_12377);
or U13640 (N_13640,N_12256,N_12595);
nand U13641 (N_13641,N_12004,N_12092);
and U13642 (N_13642,N_12667,N_12534);
xnor U13643 (N_13643,N_12666,N_12006);
nor U13644 (N_13644,N_12656,N_12295);
or U13645 (N_13645,N_12752,N_12174);
xnor U13646 (N_13646,N_12081,N_12652);
nand U13647 (N_13647,N_12436,N_12459);
xnor U13648 (N_13648,N_12327,N_12368);
xor U13649 (N_13649,N_12007,N_12132);
or U13650 (N_13650,N_12755,N_12270);
or U13651 (N_13651,N_12939,N_12585);
or U13652 (N_13652,N_12967,N_12883);
or U13653 (N_13653,N_12804,N_12825);
xnor U13654 (N_13654,N_12355,N_12522);
xnor U13655 (N_13655,N_12707,N_12634);
or U13656 (N_13656,N_12408,N_12494);
xor U13657 (N_13657,N_12220,N_12616);
and U13658 (N_13658,N_12013,N_12521);
nor U13659 (N_13659,N_12819,N_12532);
nor U13660 (N_13660,N_12924,N_12308);
or U13661 (N_13661,N_12702,N_12898);
or U13662 (N_13662,N_12103,N_12172);
xor U13663 (N_13663,N_12988,N_12329);
xnor U13664 (N_13664,N_12875,N_12666);
and U13665 (N_13665,N_12465,N_12996);
and U13666 (N_13666,N_12644,N_12766);
or U13667 (N_13667,N_12226,N_12624);
nor U13668 (N_13668,N_12370,N_12560);
nand U13669 (N_13669,N_12176,N_12387);
xnor U13670 (N_13670,N_12732,N_12418);
or U13671 (N_13671,N_12880,N_12823);
nor U13672 (N_13672,N_12719,N_12556);
xor U13673 (N_13673,N_12843,N_12035);
nand U13674 (N_13674,N_12648,N_12891);
and U13675 (N_13675,N_12515,N_12615);
xnor U13676 (N_13676,N_12227,N_12117);
or U13677 (N_13677,N_12926,N_12491);
nand U13678 (N_13678,N_12825,N_12812);
and U13679 (N_13679,N_12855,N_12828);
and U13680 (N_13680,N_12986,N_12115);
xnor U13681 (N_13681,N_12447,N_12811);
and U13682 (N_13682,N_12373,N_12568);
and U13683 (N_13683,N_12650,N_12116);
and U13684 (N_13684,N_12582,N_12832);
or U13685 (N_13685,N_12706,N_12157);
nor U13686 (N_13686,N_12889,N_12418);
and U13687 (N_13687,N_12814,N_12336);
and U13688 (N_13688,N_12714,N_12309);
xor U13689 (N_13689,N_12246,N_12613);
nor U13690 (N_13690,N_12152,N_12627);
nand U13691 (N_13691,N_12909,N_12595);
nand U13692 (N_13692,N_12131,N_12348);
nand U13693 (N_13693,N_12249,N_12236);
and U13694 (N_13694,N_12442,N_12762);
or U13695 (N_13695,N_12361,N_12035);
nor U13696 (N_13696,N_12760,N_12242);
nor U13697 (N_13697,N_12264,N_12482);
and U13698 (N_13698,N_12152,N_12779);
or U13699 (N_13699,N_12261,N_12782);
and U13700 (N_13700,N_12705,N_12070);
and U13701 (N_13701,N_12123,N_12165);
xor U13702 (N_13702,N_12636,N_12224);
nand U13703 (N_13703,N_12478,N_12333);
nor U13704 (N_13704,N_12000,N_12177);
xor U13705 (N_13705,N_12427,N_12706);
xnor U13706 (N_13706,N_12859,N_12531);
nand U13707 (N_13707,N_12647,N_12910);
or U13708 (N_13708,N_12739,N_12659);
nor U13709 (N_13709,N_12921,N_12620);
nor U13710 (N_13710,N_12353,N_12303);
nand U13711 (N_13711,N_12157,N_12126);
nor U13712 (N_13712,N_12696,N_12998);
or U13713 (N_13713,N_12525,N_12794);
nand U13714 (N_13714,N_12096,N_12078);
xor U13715 (N_13715,N_12050,N_12852);
nand U13716 (N_13716,N_12062,N_12930);
nand U13717 (N_13717,N_12560,N_12297);
nand U13718 (N_13718,N_12210,N_12798);
or U13719 (N_13719,N_12589,N_12854);
nor U13720 (N_13720,N_12770,N_12964);
nor U13721 (N_13721,N_12909,N_12584);
or U13722 (N_13722,N_12769,N_12404);
xor U13723 (N_13723,N_12401,N_12519);
and U13724 (N_13724,N_12333,N_12932);
and U13725 (N_13725,N_12723,N_12456);
nor U13726 (N_13726,N_12828,N_12341);
or U13727 (N_13727,N_12855,N_12257);
or U13728 (N_13728,N_12968,N_12698);
and U13729 (N_13729,N_12090,N_12669);
and U13730 (N_13730,N_12651,N_12542);
and U13731 (N_13731,N_12781,N_12828);
and U13732 (N_13732,N_12280,N_12145);
or U13733 (N_13733,N_12646,N_12294);
xor U13734 (N_13734,N_12080,N_12055);
xor U13735 (N_13735,N_12206,N_12399);
nand U13736 (N_13736,N_12556,N_12192);
nand U13737 (N_13737,N_12456,N_12779);
nor U13738 (N_13738,N_12098,N_12679);
and U13739 (N_13739,N_12308,N_12720);
nor U13740 (N_13740,N_12797,N_12994);
and U13741 (N_13741,N_12162,N_12297);
nand U13742 (N_13742,N_12769,N_12898);
xnor U13743 (N_13743,N_12658,N_12995);
or U13744 (N_13744,N_12728,N_12741);
nor U13745 (N_13745,N_12522,N_12912);
nand U13746 (N_13746,N_12668,N_12875);
xor U13747 (N_13747,N_12329,N_12794);
nand U13748 (N_13748,N_12125,N_12861);
nor U13749 (N_13749,N_12909,N_12980);
xnor U13750 (N_13750,N_12717,N_12015);
xor U13751 (N_13751,N_12398,N_12564);
nor U13752 (N_13752,N_12596,N_12400);
and U13753 (N_13753,N_12262,N_12887);
nor U13754 (N_13754,N_12678,N_12384);
nand U13755 (N_13755,N_12188,N_12330);
or U13756 (N_13756,N_12030,N_12387);
and U13757 (N_13757,N_12260,N_12964);
or U13758 (N_13758,N_12451,N_12681);
nand U13759 (N_13759,N_12886,N_12728);
and U13760 (N_13760,N_12972,N_12716);
xnor U13761 (N_13761,N_12601,N_12826);
nand U13762 (N_13762,N_12694,N_12806);
and U13763 (N_13763,N_12616,N_12080);
nand U13764 (N_13764,N_12772,N_12311);
or U13765 (N_13765,N_12727,N_12021);
and U13766 (N_13766,N_12125,N_12982);
nor U13767 (N_13767,N_12746,N_12981);
or U13768 (N_13768,N_12634,N_12819);
or U13769 (N_13769,N_12477,N_12393);
and U13770 (N_13770,N_12055,N_12566);
xnor U13771 (N_13771,N_12062,N_12304);
nand U13772 (N_13772,N_12156,N_12729);
nor U13773 (N_13773,N_12794,N_12280);
nor U13774 (N_13774,N_12461,N_12826);
nand U13775 (N_13775,N_12768,N_12226);
or U13776 (N_13776,N_12368,N_12010);
xor U13777 (N_13777,N_12071,N_12980);
xnor U13778 (N_13778,N_12904,N_12036);
or U13779 (N_13779,N_12298,N_12526);
and U13780 (N_13780,N_12916,N_12458);
nor U13781 (N_13781,N_12327,N_12595);
xor U13782 (N_13782,N_12355,N_12662);
or U13783 (N_13783,N_12653,N_12408);
xnor U13784 (N_13784,N_12958,N_12222);
xor U13785 (N_13785,N_12069,N_12843);
xor U13786 (N_13786,N_12979,N_12873);
or U13787 (N_13787,N_12767,N_12049);
and U13788 (N_13788,N_12002,N_12462);
nand U13789 (N_13789,N_12503,N_12039);
xnor U13790 (N_13790,N_12021,N_12266);
nand U13791 (N_13791,N_12683,N_12102);
and U13792 (N_13792,N_12962,N_12562);
nor U13793 (N_13793,N_12445,N_12396);
and U13794 (N_13794,N_12239,N_12887);
or U13795 (N_13795,N_12489,N_12775);
nand U13796 (N_13796,N_12018,N_12519);
or U13797 (N_13797,N_12386,N_12055);
or U13798 (N_13798,N_12368,N_12181);
and U13799 (N_13799,N_12602,N_12227);
and U13800 (N_13800,N_12052,N_12133);
and U13801 (N_13801,N_12039,N_12949);
xor U13802 (N_13802,N_12921,N_12838);
or U13803 (N_13803,N_12205,N_12965);
or U13804 (N_13804,N_12930,N_12004);
nor U13805 (N_13805,N_12350,N_12625);
nor U13806 (N_13806,N_12721,N_12995);
nor U13807 (N_13807,N_12581,N_12334);
nand U13808 (N_13808,N_12133,N_12529);
or U13809 (N_13809,N_12030,N_12039);
and U13810 (N_13810,N_12590,N_12805);
nand U13811 (N_13811,N_12665,N_12401);
or U13812 (N_13812,N_12266,N_12438);
xor U13813 (N_13813,N_12893,N_12322);
and U13814 (N_13814,N_12607,N_12699);
or U13815 (N_13815,N_12619,N_12425);
nor U13816 (N_13816,N_12562,N_12193);
and U13817 (N_13817,N_12590,N_12778);
or U13818 (N_13818,N_12344,N_12751);
or U13819 (N_13819,N_12473,N_12607);
nor U13820 (N_13820,N_12996,N_12662);
nand U13821 (N_13821,N_12336,N_12065);
xor U13822 (N_13822,N_12787,N_12020);
or U13823 (N_13823,N_12827,N_12735);
nor U13824 (N_13824,N_12676,N_12063);
xnor U13825 (N_13825,N_12822,N_12687);
nand U13826 (N_13826,N_12307,N_12888);
or U13827 (N_13827,N_12137,N_12880);
nor U13828 (N_13828,N_12244,N_12856);
and U13829 (N_13829,N_12436,N_12491);
xnor U13830 (N_13830,N_12857,N_12386);
xnor U13831 (N_13831,N_12761,N_12044);
nor U13832 (N_13832,N_12935,N_12847);
and U13833 (N_13833,N_12133,N_12344);
nand U13834 (N_13834,N_12370,N_12204);
and U13835 (N_13835,N_12855,N_12379);
nor U13836 (N_13836,N_12424,N_12274);
xor U13837 (N_13837,N_12158,N_12226);
or U13838 (N_13838,N_12315,N_12193);
nor U13839 (N_13839,N_12851,N_12072);
and U13840 (N_13840,N_12325,N_12657);
or U13841 (N_13841,N_12046,N_12030);
nand U13842 (N_13842,N_12115,N_12405);
or U13843 (N_13843,N_12053,N_12562);
and U13844 (N_13844,N_12351,N_12916);
nand U13845 (N_13845,N_12567,N_12364);
and U13846 (N_13846,N_12231,N_12750);
or U13847 (N_13847,N_12655,N_12231);
xor U13848 (N_13848,N_12440,N_12091);
and U13849 (N_13849,N_12652,N_12388);
nor U13850 (N_13850,N_12316,N_12304);
xnor U13851 (N_13851,N_12214,N_12502);
nor U13852 (N_13852,N_12487,N_12145);
nand U13853 (N_13853,N_12804,N_12480);
or U13854 (N_13854,N_12130,N_12187);
xnor U13855 (N_13855,N_12640,N_12283);
nor U13856 (N_13856,N_12717,N_12194);
nand U13857 (N_13857,N_12167,N_12412);
nor U13858 (N_13858,N_12614,N_12121);
and U13859 (N_13859,N_12919,N_12508);
and U13860 (N_13860,N_12856,N_12516);
xnor U13861 (N_13861,N_12997,N_12976);
or U13862 (N_13862,N_12533,N_12787);
or U13863 (N_13863,N_12403,N_12553);
nand U13864 (N_13864,N_12747,N_12813);
or U13865 (N_13865,N_12625,N_12571);
nor U13866 (N_13866,N_12753,N_12760);
or U13867 (N_13867,N_12570,N_12843);
or U13868 (N_13868,N_12336,N_12945);
and U13869 (N_13869,N_12823,N_12924);
nor U13870 (N_13870,N_12828,N_12697);
or U13871 (N_13871,N_12063,N_12418);
nor U13872 (N_13872,N_12420,N_12528);
or U13873 (N_13873,N_12408,N_12226);
nor U13874 (N_13874,N_12278,N_12157);
nor U13875 (N_13875,N_12049,N_12557);
or U13876 (N_13876,N_12470,N_12960);
nor U13877 (N_13877,N_12812,N_12460);
and U13878 (N_13878,N_12856,N_12302);
nor U13879 (N_13879,N_12853,N_12793);
xor U13880 (N_13880,N_12935,N_12036);
or U13881 (N_13881,N_12509,N_12308);
xor U13882 (N_13882,N_12424,N_12599);
nand U13883 (N_13883,N_12234,N_12118);
nor U13884 (N_13884,N_12595,N_12566);
and U13885 (N_13885,N_12055,N_12913);
nand U13886 (N_13886,N_12075,N_12233);
nor U13887 (N_13887,N_12948,N_12410);
xnor U13888 (N_13888,N_12286,N_12085);
and U13889 (N_13889,N_12236,N_12071);
nand U13890 (N_13890,N_12837,N_12604);
xnor U13891 (N_13891,N_12503,N_12919);
and U13892 (N_13892,N_12218,N_12522);
xnor U13893 (N_13893,N_12466,N_12656);
and U13894 (N_13894,N_12633,N_12252);
or U13895 (N_13895,N_12337,N_12819);
or U13896 (N_13896,N_12559,N_12138);
xor U13897 (N_13897,N_12263,N_12592);
nor U13898 (N_13898,N_12897,N_12927);
and U13899 (N_13899,N_12955,N_12759);
and U13900 (N_13900,N_12035,N_12968);
nand U13901 (N_13901,N_12267,N_12820);
xor U13902 (N_13902,N_12743,N_12643);
and U13903 (N_13903,N_12045,N_12682);
and U13904 (N_13904,N_12153,N_12684);
nand U13905 (N_13905,N_12920,N_12996);
or U13906 (N_13906,N_12478,N_12060);
nor U13907 (N_13907,N_12894,N_12226);
and U13908 (N_13908,N_12970,N_12762);
or U13909 (N_13909,N_12461,N_12956);
and U13910 (N_13910,N_12859,N_12790);
xor U13911 (N_13911,N_12305,N_12070);
nand U13912 (N_13912,N_12185,N_12828);
nor U13913 (N_13913,N_12744,N_12311);
nand U13914 (N_13914,N_12768,N_12075);
or U13915 (N_13915,N_12954,N_12041);
and U13916 (N_13916,N_12914,N_12890);
or U13917 (N_13917,N_12251,N_12324);
or U13918 (N_13918,N_12609,N_12194);
nor U13919 (N_13919,N_12537,N_12214);
nor U13920 (N_13920,N_12332,N_12478);
xnor U13921 (N_13921,N_12474,N_12586);
nand U13922 (N_13922,N_12362,N_12748);
xnor U13923 (N_13923,N_12795,N_12031);
nor U13924 (N_13924,N_12149,N_12281);
nor U13925 (N_13925,N_12756,N_12684);
and U13926 (N_13926,N_12274,N_12203);
nor U13927 (N_13927,N_12809,N_12875);
xnor U13928 (N_13928,N_12919,N_12927);
xnor U13929 (N_13929,N_12344,N_12715);
or U13930 (N_13930,N_12542,N_12436);
and U13931 (N_13931,N_12511,N_12448);
or U13932 (N_13932,N_12994,N_12855);
nor U13933 (N_13933,N_12493,N_12325);
nor U13934 (N_13934,N_12492,N_12502);
nand U13935 (N_13935,N_12163,N_12541);
nor U13936 (N_13936,N_12871,N_12950);
or U13937 (N_13937,N_12619,N_12683);
or U13938 (N_13938,N_12956,N_12658);
xor U13939 (N_13939,N_12929,N_12901);
or U13940 (N_13940,N_12467,N_12307);
xnor U13941 (N_13941,N_12237,N_12711);
nand U13942 (N_13942,N_12157,N_12184);
nand U13943 (N_13943,N_12402,N_12919);
or U13944 (N_13944,N_12575,N_12261);
xnor U13945 (N_13945,N_12277,N_12822);
and U13946 (N_13946,N_12537,N_12616);
or U13947 (N_13947,N_12413,N_12096);
nor U13948 (N_13948,N_12189,N_12723);
xor U13949 (N_13949,N_12151,N_12713);
xnor U13950 (N_13950,N_12411,N_12420);
xor U13951 (N_13951,N_12527,N_12440);
xor U13952 (N_13952,N_12798,N_12315);
xor U13953 (N_13953,N_12355,N_12688);
xnor U13954 (N_13954,N_12670,N_12773);
nor U13955 (N_13955,N_12207,N_12285);
nand U13956 (N_13956,N_12156,N_12935);
or U13957 (N_13957,N_12641,N_12289);
and U13958 (N_13958,N_12944,N_12628);
xor U13959 (N_13959,N_12763,N_12269);
and U13960 (N_13960,N_12860,N_12961);
and U13961 (N_13961,N_12266,N_12778);
or U13962 (N_13962,N_12391,N_12355);
nor U13963 (N_13963,N_12068,N_12538);
nor U13964 (N_13964,N_12347,N_12432);
or U13965 (N_13965,N_12817,N_12219);
xor U13966 (N_13966,N_12656,N_12171);
and U13967 (N_13967,N_12260,N_12393);
and U13968 (N_13968,N_12133,N_12864);
xor U13969 (N_13969,N_12564,N_12753);
nand U13970 (N_13970,N_12076,N_12728);
nand U13971 (N_13971,N_12991,N_12483);
or U13972 (N_13972,N_12341,N_12518);
xor U13973 (N_13973,N_12916,N_12561);
nor U13974 (N_13974,N_12605,N_12871);
xor U13975 (N_13975,N_12702,N_12789);
or U13976 (N_13976,N_12867,N_12676);
and U13977 (N_13977,N_12720,N_12554);
nand U13978 (N_13978,N_12720,N_12151);
nor U13979 (N_13979,N_12306,N_12927);
xnor U13980 (N_13980,N_12744,N_12094);
nand U13981 (N_13981,N_12248,N_12799);
or U13982 (N_13982,N_12591,N_12234);
xor U13983 (N_13983,N_12793,N_12523);
nor U13984 (N_13984,N_12834,N_12074);
xor U13985 (N_13985,N_12614,N_12458);
nor U13986 (N_13986,N_12269,N_12652);
xor U13987 (N_13987,N_12689,N_12461);
nor U13988 (N_13988,N_12297,N_12820);
and U13989 (N_13989,N_12175,N_12838);
and U13990 (N_13990,N_12360,N_12264);
xor U13991 (N_13991,N_12419,N_12104);
or U13992 (N_13992,N_12008,N_12408);
and U13993 (N_13993,N_12435,N_12266);
and U13994 (N_13994,N_12901,N_12576);
and U13995 (N_13995,N_12712,N_12260);
nor U13996 (N_13996,N_12639,N_12347);
nand U13997 (N_13997,N_12753,N_12105);
and U13998 (N_13998,N_12580,N_12211);
nand U13999 (N_13999,N_12671,N_12107);
xnor U14000 (N_14000,N_13440,N_13712);
or U14001 (N_14001,N_13448,N_13290);
xor U14002 (N_14002,N_13112,N_13141);
xnor U14003 (N_14003,N_13518,N_13048);
nand U14004 (N_14004,N_13232,N_13840);
xor U14005 (N_14005,N_13601,N_13709);
xor U14006 (N_14006,N_13167,N_13338);
or U14007 (N_14007,N_13857,N_13435);
nor U14008 (N_14008,N_13864,N_13910);
xnor U14009 (N_14009,N_13230,N_13997);
or U14010 (N_14010,N_13936,N_13198);
or U14011 (N_14011,N_13066,N_13498);
nand U14012 (N_14012,N_13433,N_13137);
or U14013 (N_14013,N_13236,N_13134);
nand U14014 (N_14014,N_13037,N_13256);
or U14015 (N_14015,N_13504,N_13416);
xnor U14016 (N_14016,N_13485,N_13047);
nor U14017 (N_14017,N_13704,N_13662);
nand U14018 (N_14018,N_13104,N_13547);
and U14019 (N_14019,N_13337,N_13725);
and U14020 (N_14020,N_13376,N_13226);
nor U14021 (N_14021,N_13180,N_13564);
or U14022 (N_14022,N_13646,N_13636);
xor U14023 (N_14023,N_13312,N_13332);
or U14024 (N_14024,N_13330,N_13396);
xor U14025 (N_14025,N_13072,N_13943);
nand U14026 (N_14026,N_13912,N_13001);
nand U14027 (N_14027,N_13061,N_13696);
nor U14028 (N_14028,N_13272,N_13701);
nand U14029 (N_14029,N_13475,N_13611);
nand U14030 (N_14030,N_13521,N_13270);
nor U14031 (N_14031,N_13306,N_13838);
nand U14032 (N_14032,N_13217,N_13613);
nand U14033 (N_14033,N_13560,N_13428);
xor U14034 (N_14034,N_13013,N_13251);
nor U14035 (N_14035,N_13426,N_13628);
nor U14036 (N_14036,N_13933,N_13625);
and U14037 (N_14037,N_13220,N_13122);
and U14038 (N_14038,N_13873,N_13827);
or U14039 (N_14039,N_13264,N_13238);
or U14040 (N_14040,N_13216,N_13599);
xor U14041 (N_14041,N_13019,N_13456);
nand U14042 (N_14042,N_13716,N_13576);
nor U14043 (N_14043,N_13310,N_13239);
and U14044 (N_14044,N_13612,N_13170);
xnor U14045 (N_14045,N_13593,N_13073);
nand U14046 (N_14046,N_13993,N_13591);
xnor U14047 (N_14047,N_13637,N_13314);
and U14048 (N_14048,N_13516,N_13252);
or U14049 (N_14049,N_13453,N_13057);
nand U14050 (N_14050,N_13968,N_13004);
or U14051 (N_14051,N_13169,N_13821);
or U14052 (N_14052,N_13941,N_13111);
nor U14053 (N_14053,N_13519,N_13419);
or U14054 (N_14054,N_13010,N_13443);
or U14055 (N_14055,N_13370,N_13710);
or U14056 (N_14056,N_13015,N_13179);
nand U14057 (N_14057,N_13411,N_13438);
xnor U14058 (N_14058,N_13298,N_13157);
xor U14059 (N_14059,N_13746,N_13344);
nand U14060 (N_14060,N_13667,N_13371);
nand U14061 (N_14061,N_13720,N_13598);
nand U14062 (N_14062,N_13178,N_13702);
and U14063 (N_14063,N_13722,N_13724);
xnor U14064 (N_14064,N_13816,N_13621);
or U14065 (N_14065,N_13536,N_13723);
and U14066 (N_14066,N_13647,N_13358);
nor U14067 (N_14067,N_13835,N_13817);
nor U14068 (N_14068,N_13368,N_13932);
nor U14069 (N_14069,N_13302,N_13204);
or U14070 (N_14070,N_13892,N_13695);
or U14071 (N_14071,N_13693,N_13703);
nor U14072 (N_14072,N_13789,N_13249);
nor U14073 (N_14073,N_13118,N_13361);
and U14074 (N_14074,N_13493,N_13886);
or U14075 (N_14075,N_13415,N_13793);
nand U14076 (N_14076,N_13934,N_13904);
nand U14077 (N_14077,N_13096,N_13555);
xor U14078 (N_14078,N_13676,N_13558);
nor U14079 (N_14079,N_13291,N_13138);
or U14080 (N_14080,N_13742,N_13920);
nand U14081 (N_14081,N_13820,N_13758);
or U14082 (N_14082,N_13745,N_13152);
xor U14083 (N_14083,N_13948,N_13786);
nor U14084 (N_14084,N_13201,N_13641);
nor U14085 (N_14085,N_13574,N_13403);
xor U14086 (N_14086,N_13374,N_13327);
and U14087 (N_14087,N_13492,N_13799);
or U14088 (N_14088,N_13382,N_13117);
nor U14089 (N_14089,N_13785,N_13911);
or U14090 (N_14090,N_13577,N_13590);
nand U14091 (N_14091,N_13867,N_13592);
xnor U14092 (N_14092,N_13511,N_13120);
nor U14093 (N_14093,N_13441,N_13014);
nand U14094 (N_14094,N_13992,N_13472);
nand U14095 (N_14095,N_13035,N_13034);
xnor U14096 (N_14096,N_13397,N_13043);
nand U14097 (N_14097,N_13732,N_13285);
nand U14098 (N_14098,N_13607,N_13727);
nand U14099 (N_14099,N_13208,N_13153);
nand U14100 (N_14100,N_13069,N_13770);
nand U14101 (N_14101,N_13622,N_13324);
nand U14102 (N_14102,N_13342,N_13654);
nand U14103 (N_14103,N_13103,N_13868);
and U14104 (N_14104,N_13953,N_13529);
nor U14105 (N_14105,N_13352,N_13533);
or U14106 (N_14106,N_13429,N_13478);
or U14107 (N_14107,N_13460,N_13675);
xor U14108 (N_14108,N_13212,N_13954);
and U14109 (N_14109,N_13802,N_13483);
nand U14110 (N_14110,N_13250,N_13909);
nor U14111 (N_14111,N_13263,N_13186);
and U14112 (N_14112,N_13610,N_13819);
and U14113 (N_14113,N_13549,N_13095);
or U14114 (N_14114,N_13713,N_13000);
nand U14115 (N_14115,N_13174,N_13214);
xor U14116 (N_14116,N_13307,N_13595);
and U14117 (N_14117,N_13060,N_13798);
and U14118 (N_14118,N_13353,N_13931);
and U14119 (N_14119,N_13862,N_13102);
or U14120 (N_14120,N_13020,N_13737);
nand U14121 (N_14121,N_13181,N_13412);
nand U14122 (N_14122,N_13049,N_13050);
nor U14123 (N_14123,N_13804,N_13183);
nand U14124 (N_14124,N_13045,N_13751);
nor U14125 (N_14125,N_13889,N_13557);
nand U14126 (N_14126,N_13237,N_13143);
and U14127 (N_14127,N_13729,N_13063);
and U14128 (N_14128,N_13631,N_13972);
nor U14129 (N_14129,N_13458,N_13017);
or U14130 (N_14130,N_13356,N_13707);
nand U14131 (N_14131,N_13445,N_13869);
and U14132 (N_14132,N_13331,N_13828);
xnor U14133 (N_14133,N_13300,N_13464);
nand U14134 (N_14134,N_13747,N_13147);
and U14135 (N_14135,N_13124,N_13357);
or U14136 (N_14136,N_13373,N_13121);
and U14137 (N_14137,N_13506,N_13618);
nand U14138 (N_14138,N_13148,N_13790);
nor U14139 (N_14139,N_13313,N_13683);
xor U14140 (N_14140,N_13859,N_13594);
and U14141 (N_14141,N_13561,N_13530);
and U14142 (N_14142,N_13552,N_13818);
nand U14143 (N_14143,N_13788,N_13898);
nor U14144 (N_14144,N_13513,N_13490);
or U14145 (N_14145,N_13856,N_13036);
xnor U14146 (N_14146,N_13190,N_13627);
nor U14147 (N_14147,N_13949,N_13774);
xor U14148 (N_14148,N_13345,N_13149);
and U14149 (N_14149,N_13092,N_13109);
nor U14150 (N_14150,N_13056,N_13571);
nand U14151 (N_14151,N_13772,N_13038);
xor U14152 (N_14152,N_13224,N_13455);
nor U14153 (N_14153,N_13466,N_13841);
nand U14154 (N_14154,N_13962,N_13915);
nor U14155 (N_14155,N_13207,N_13024);
nor U14156 (N_14156,N_13741,N_13283);
and U14157 (N_14157,N_13858,N_13215);
xor U14158 (N_14158,N_13273,N_13287);
xor U14159 (N_14159,N_13754,N_13655);
nand U14160 (N_14160,N_13286,N_13971);
xor U14161 (N_14161,N_13379,N_13658);
and U14162 (N_14162,N_13410,N_13219);
and U14163 (N_14163,N_13218,N_13086);
nand U14164 (N_14164,N_13807,N_13903);
nand U14165 (N_14165,N_13003,N_13981);
and U14166 (N_14166,N_13527,N_13814);
or U14167 (N_14167,N_13360,N_13184);
or U14168 (N_14168,N_13284,N_13791);
nor U14169 (N_14169,N_13570,N_13127);
xor U14170 (N_14170,N_13206,N_13914);
nor U14171 (N_14171,N_13517,N_13481);
nand U14172 (N_14172,N_13486,N_13457);
or U14173 (N_14173,N_13765,N_13930);
nor U14174 (N_14174,N_13626,N_13303);
xnor U14175 (N_14175,N_13918,N_13878);
nand U14176 (N_14176,N_13372,N_13580);
or U14177 (N_14177,N_13865,N_13189);
and U14178 (N_14178,N_13294,N_13719);
xnor U14179 (N_14179,N_13267,N_13805);
nand U14180 (N_14180,N_13940,N_13196);
xor U14181 (N_14181,N_13076,N_13105);
xnor U14182 (N_14182,N_13783,N_13497);
xnor U14183 (N_14183,N_13586,N_13512);
or U14184 (N_14184,N_13579,N_13829);
xor U14185 (N_14185,N_13797,N_13008);
xor U14186 (N_14186,N_13334,N_13192);
nand U14187 (N_14187,N_13967,N_13163);
or U14188 (N_14188,N_13896,N_13398);
xor U14189 (N_14189,N_13671,N_13028);
nor U14190 (N_14190,N_13489,N_13359);
nand U14191 (N_14191,N_13444,N_13094);
or U14192 (N_14192,N_13074,N_13587);
nor U14193 (N_14193,N_13316,N_13759);
nor U14194 (N_14194,N_13258,N_13756);
or U14195 (N_14195,N_13053,N_13810);
xor U14196 (N_14196,N_13969,N_13247);
or U14197 (N_14197,N_13325,N_13452);
nand U14198 (N_14198,N_13301,N_13939);
nor U14199 (N_14199,N_13023,N_13439);
nand U14200 (N_14200,N_13150,N_13678);
and U14201 (N_14201,N_13202,N_13479);
nand U14202 (N_14202,N_13950,N_13385);
and U14203 (N_14203,N_13668,N_13826);
or U14204 (N_14204,N_13830,N_13450);
or U14205 (N_14205,N_13211,N_13604);
and U14206 (N_14206,N_13348,N_13566);
and U14207 (N_14207,N_13084,N_13752);
nand U14208 (N_14208,N_13364,N_13917);
or U14209 (N_14209,N_13349,N_13762);
or U14210 (N_14210,N_13743,N_13656);
or U14211 (N_14211,N_13108,N_13554);
xnor U14212 (N_14212,N_13142,N_13381);
xor U14213 (N_14213,N_13899,N_13669);
xnor U14214 (N_14214,N_13488,N_13528);
and U14215 (N_14215,N_13402,N_13383);
and U14216 (N_14216,N_13246,N_13449);
xor U14217 (N_14217,N_13424,N_13494);
or U14218 (N_14218,N_13923,N_13919);
or U14219 (N_14219,N_13694,N_13387);
or U14220 (N_14220,N_13677,N_13400);
xnor U14221 (N_14221,N_13854,N_13843);
nor U14222 (N_14222,N_13225,N_13187);
or U14223 (N_14223,N_13876,N_13659);
xnor U14224 (N_14224,N_13041,N_13687);
nor U14225 (N_14225,N_13796,N_13391);
nand U14226 (N_14226,N_13495,N_13423);
nand U14227 (N_14227,N_13434,N_13699);
xnor U14228 (N_14228,N_13871,N_13781);
or U14229 (N_14229,N_13526,N_13648);
and U14230 (N_14230,N_13366,N_13144);
nand U14231 (N_14231,N_13062,N_13525);
nor U14232 (N_14232,N_13228,N_13085);
nor U14233 (N_14233,N_13308,N_13947);
nor U14234 (N_14234,N_13437,N_13945);
xnor U14235 (N_14235,N_13874,N_13280);
or U14236 (N_14236,N_13227,N_13705);
and U14237 (N_14237,N_13319,N_13395);
and U14238 (N_14238,N_13323,N_13771);
and U14239 (N_14239,N_13907,N_13474);
nand U14240 (N_14240,N_13575,N_13254);
xnor U14241 (N_14241,N_13380,N_13064);
xnor U14242 (N_14242,N_13642,N_13690);
or U14243 (N_14243,N_13900,N_13763);
and U14244 (N_14244,N_13362,N_13089);
nand U14245 (N_14245,N_13059,N_13422);
xor U14246 (N_14246,N_13347,N_13652);
xor U14247 (N_14247,N_13305,N_13970);
nor U14248 (N_14248,N_13906,N_13459);
xnor U14249 (N_14249,N_13735,N_13275);
or U14250 (N_14250,N_13119,N_13235);
and U14251 (N_14251,N_13986,N_13461);
or U14252 (N_14252,N_13293,N_13384);
nand U14253 (N_14253,N_13309,N_13006);
xor U14254 (N_14254,N_13633,N_13018);
or U14255 (N_14255,N_13957,N_13132);
nor U14256 (N_14256,N_13908,N_13768);
nor U14257 (N_14257,N_13688,N_13110);
or U14258 (N_14258,N_13476,N_13133);
nor U14259 (N_14259,N_13617,N_13806);
xnor U14260 (N_14260,N_13209,N_13556);
and U14261 (N_14261,N_13988,N_13418);
nor U14262 (N_14262,N_13711,N_13401);
or U14263 (N_14263,N_13921,N_13650);
nor U14264 (N_14264,N_13087,N_13800);
or U14265 (N_14265,N_13531,N_13213);
or U14266 (N_14266,N_13161,N_13990);
and U14267 (N_14267,N_13255,N_13354);
nand U14268 (N_14268,N_13644,N_13162);
or U14269 (N_14269,N_13421,N_13311);
or U14270 (N_14270,N_13905,N_13794);
nor U14271 (N_14271,N_13075,N_13099);
or U14272 (N_14272,N_13399,N_13692);
and U14273 (N_14273,N_13715,N_13935);
nand U14274 (N_14274,N_13427,N_13825);
xnor U14275 (N_14275,N_13714,N_13893);
nand U14276 (N_14276,N_13801,N_13276);
nor U14277 (N_14277,N_13991,N_13365);
and U14278 (N_14278,N_13158,N_13259);
or U14279 (N_14279,N_13977,N_13507);
or U14280 (N_14280,N_13686,N_13779);
and U14281 (N_14281,N_13545,N_13128);
and U14282 (N_14282,N_13406,N_13866);
or U14283 (N_14283,N_13393,N_13510);
or U14284 (N_14284,N_13965,N_13156);
nor U14285 (N_14285,N_13245,N_13261);
nand U14286 (N_14286,N_13098,N_13262);
nand U14287 (N_14287,N_13113,N_13040);
xor U14288 (N_14288,N_13665,N_13567);
nor U14289 (N_14289,N_13363,N_13462);
nor U14290 (N_14290,N_13346,N_13145);
and U14291 (N_14291,N_13223,N_13585);
nand U14292 (N_14292,N_13279,N_13042);
and U14293 (N_14293,N_13271,N_13375);
or U14294 (N_14294,N_13321,N_13386);
and U14295 (N_14295,N_13776,N_13182);
or U14296 (N_14296,N_13605,N_13740);
nor U14297 (N_14297,N_13634,N_13755);
nor U14298 (N_14298,N_13265,N_13054);
or U14299 (N_14299,N_13568,N_13884);
nor U14300 (N_14300,N_13822,N_13578);
nand U14301 (N_14301,N_13734,N_13975);
nand U14302 (N_14302,N_13787,N_13340);
and U14303 (N_14303,N_13388,N_13295);
xnor U14304 (N_14304,N_13191,N_13292);
nand U14305 (N_14305,N_13088,N_13377);
xnor U14306 (N_14306,N_13199,N_13477);
xnor U14307 (N_14307,N_13680,N_13482);
nand U14308 (N_14308,N_13890,N_13995);
nor U14309 (N_14309,N_13684,N_13846);
nand U14310 (N_14310,N_13322,N_13985);
xnor U14311 (N_14311,N_13509,N_13879);
or U14312 (N_14312,N_13065,N_13185);
xor U14313 (N_14313,N_13135,N_13581);
nand U14314 (N_14314,N_13657,N_13942);
nor U14315 (N_14315,N_13203,N_13436);
nand U14316 (N_14316,N_13480,N_13297);
and U14317 (N_14317,N_13154,N_13012);
or U14318 (N_14318,N_13537,N_13584);
xnor U14319 (N_14319,N_13058,N_13660);
nor U14320 (N_14320,N_13431,N_13863);
xnor U14321 (N_14321,N_13165,N_13620);
and U14322 (N_14322,N_13877,N_13649);
nor U14323 (N_14323,N_13390,N_13335);
xnor U14324 (N_14324,N_13663,N_13522);
or U14325 (N_14325,N_13039,N_13151);
xor U14326 (N_14326,N_13430,N_13274);
xor U14327 (N_14327,N_13955,N_13333);
xor U14328 (N_14328,N_13168,N_13243);
nand U14329 (N_14329,N_13367,N_13093);
xnor U14330 (N_14330,N_13471,N_13160);
and U14331 (N_14331,N_13539,N_13559);
or U14332 (N_14332,N_13176,N_13469);
xnor U14333 (N_14333,N_13125,N_13229);
or U14334 (N_14334,N_13491,N_13304);
or U14335 (N_14335,N_13823,N_13408);
nor U14336 (N_14336,N_13027,N_13999);
nand U14337 (N_14337,N_13775,N_13473);
and U14338 (N_14338,N_13540,N_13425);
nor U14339 (N_14339,N_13257,N_13881);
and U14340 (N_14340,N_13624,N_13523);
xnor U14341 (N_14341,N_13928,N_13922);
nand U14342 (N_14342,N_13760,N_13011);
nand U14343 (N_14343,N_13514,N_13728);
xor U14344 (N_14344,N_13926,N_13639);
or U14345 (N_14345,N_13389,N_13562);
nand U14346 (N_14346,N_13916,N_13812);
nand U14347 (N_14347,N_13080,N_13984);
or U14348 (N_14348,N_13960,N_13832);
and U14349 (N_14349,N_13467,N_13956);
and U14350 (N_14350,N_13336,N_13630);
xor U14351 (N_14351,N_13468,N_13033);
nand U14352 (N_14352,N_13025,N_13414);
or U14353 (N_14353,N_13499,N_13326);
nor U14354 (N_14354,N_13629,N_13572);
and U14355 (N_14355,N_13673,N_13842);
or U14356 (N_14356,N_13546,N_13730);
xnor U14357 (N_14357,N_13753,N_13500);
nor U14358 (N_14358,N_13016,N_13139);
or U14359 (N_14359,N_13277,N_13222);
and U14360 (N_14360,N_13573,N_13851);
nand U14361 (N_14361,N_13689,N_13268);
or U14362 (N_14362,N_13031,N_13068);
or U14363 (N_14363,N_13726,N_13083);
nor U14364 (N_14364,N_13339,N_13937);
nor U14365 (N_14365,N_13974,N_13811);
nor U14366 (N_14366,N_13833,N_13515);
nand U14367 (N_14367,N_13442,N_13155);
nor U14368 (N_14368,N_13927,N_13738);
and U14369 (N_14369,N_13343,N_13731);
and U14370 (N_14370,N_13848,N_13780);
nor U14371 (N_14371,N_13407,N_13897);
and U14372 (N_14372,N_13131,N_13081);
xor U14373 (N_14373,N_13404,N_13792);
nand U14374 (N_14374,N_13685,N_13299);
or U14375 (N_14375,N_13378,N_13417);
nand U14376 (N_14376,N_13318,N_13872);
nor U14377 (N_14377,N_13706,N_13849);
nand U14378 (N_14378,N_13071,N_13761);
nor U14379 (N_14379,N_13924,N_13718);
xnor U14380 (N_14380,N_13803,N_13115);
and U14381 (N_14381,N_13964,N_13808);
and U14382 (N_14382,N_13369,N_13666);
xor U14383 (N_14383,N_13809,N_13508);
nand U14384 (N_14384,N_13670,N_13679);
and U14385 (N_14385,N_13989,N_13766);
or U14386 (N_14386,N_13982,N_13051);
and U14387 (N_14387,N_13895,N_13350);
nor U14388 (N_14388,N_13691,N_13114);
and U14389 (N_14389,N_13623,N_13976);
nand U14390 (N_14390,N_13664,N_13852);
and U14391 (N_14391,N_13861,N_13553);
nor U14392 (N_14392,N_13778,N_13882);
nand U14393 (N_14393,N_13470,N_13005);
and U14394 (N_14394,N_13317,N_13253);
or U14395 (N_14395,N_13983,N_13773);
nand U14396 (N_14396,N_13496,N_13883);
xor U14397 (N_14397,N_13888,N_13231);
nand U14398 (N_14398,N_13248,N_13171);
or U14399 (N_14399,N_13885,N_13260);
xor U14400 (N_14400,N_13195,N_13487);
xor U14401 (N_14401,N_13550,N_13077);
and U14402 (N_14402,N_13543,N_13173);
or U14403 (N_14403,N_13748,N_13606);
and U14404 (N_14404,N_13643,N_13505);
nor U14405 (N_14405,N_13880,N_13503);
nand U14406 (N_14406,N_13315,N_13834);
and U14407 (N_14407,N_13844,N_13681);
nand U14408 (N_14408,N_13355,N_13269);
or U14409 (N_14409,N_13029,N_13698);
or U14410 (N_14410,N_13980,N_13837);
nor U14411 (N_14411,N_13242,N_13538);
xor U14412 (N_14412,N_13172,N_13281);
xor U14413 (N_14413,N_13739,N_13244);
and U14414 (N_14414,N_13405,N_13320);
nand U14415 (N_14415,N_13891,N_13824);
or U14416 (N_14416,N_13901,N_13123);
and U14417 (N_14417,N_13548,N_13597);
xor U14418 (N_14418,N_13420,N_13067);
and U14419 (N_14419,N_13532,N_13409);
nand U14420 (N_14420,N_13030,N_13026);
xnor U14421 (N_14421,N_13855,N_13535);
or U14422 (N_14422,N_13126,N_13749);
nor U14423 (N_14423,N_13845,N_13130);
nor U14424 (N_14424,N_13619,N_13055);
nand U14425 (N_14425,N_13736,N_13784);
and U14426 (N_14426,N_13463,N_13973);
nand U14427 (N_14427,N_13046,N_13288);
xor U14428 (N_14428,N_13328,N_13733);
or U14429 (N_14429,N_13082,N_13501);
nand U14430 (N_14430,N_13240,N_13961);
and U14431 (N_14431,N_13944,N_13524);
or U14432 (N_14432,N_13963,N_13241);
or U14433 (N_14433,N_13853,N_13563);
xnor U14434 (N_14434,N_13465,N_13009);
and U14435 (N_14435,N_13994,N_13782);
nor U14436 (N_14436,N_13166,N_13278);
and U14437 (N_14437,N_13850,N_13987);
nand U14438 (N_14438,N_13777,N_13588);
or U14439 (N_14439,N_13645,N_13002);
or U14440 (N_14440,N_13847,N_13959);
nor U14441 (N_14441,N_13129,N_13769);
or U14442 (N_14442,N_13454,N_13392);
xor U14443 (N_14443,N_13116,N_13413);
xor U14444 (N_14444,N_13329,N_13234);
and U14445 (N_14445,N_13534,N_13600);
or U14446 (N_14446,N_13544,N_13193);
and U14447 (N_14447,N_13582,N_13007);
nor U14448 (N_14448,N_13764,N_13446);
and U14449 (N_14449,N_13674,N_13894);
nor U14450 (N_14450,N_13101,N_13795);
or U14451 (N_14451,N_13870,N_13815);
and U14452 (N_14452,N_13635,N_13032);
xor U14453 (N_14453,N_13164,N_13929);
nand U14454 (N_14454,N_13542,N_13887);
or U14455 (N_14455,N_13233,N_13106);
xnor U14456 (N_14456,N_13602,N_13177);
and U14457 (N_14457,N_13925,N_13266);
and U14458 (N_14458,N_13757,N_13836);
and U14459 (N_14459,N_13136,N_13640);
nor U14460 (N_14460,N_13188,N_13839);
nand U14461 (N_14461,N_13175,N_13551);
nand U14462 (N_14462,N_13351,N_13052);
nand U14463 (N_14463,N_13210,N_13091);
or U14464 (N_14464,N_13565,N_13140);
nand U14465 (N_14465,N_13608,N_13194);
nor U14466 (N_14466,N_13596,N_13541);
xnor U14467 (N_14467,N_13159,N_13717);
xor U14468 (N_14468,N_13682,N_13341);
xnor U14469 (N_14469,N_13197,N_13750);
or U14470 (N_14470,N_13090,N_13913);
or U14471 (N_14471,N_13205,N_13502);
or U14472 (N_14472,N_13744,N_13100);
nand U14473 (N_14473,N_13044,N_13021);
nor U14474 (N_14474,N_13813,N_13200);
xor U14475 (N_14475,N_13938,N_13998);
nor U14476 (N_14476,N_13615,N_13653);
nand U14477 (N_14477,N_13721,N_13979);
or U14478 (N_14478,N_13609,N_13708);
nor U14479 (N_14479,N_13221,N_13107);
nand U14480 (N_14480,N_13902,N_13520);
nor U14481 (N_14481,N_13583,N_13447);
or U14482 (N_14482,N_13661,N_13697);
or U14483 (N_14483,N_13616,N_13638);
and U14484 (N_14484,N_13951,N_13394);
xnor U14485 (N_14485,N_13875,N_13289);
xnor U14486 (N_14486,N_13614,N_13978);
and U14487 (N_14487,N_13296,N_13078);
nand U14488 (N_14488,N_13958,N_13146);
nand U14489 (N_14489,N_13767,N_13700);
nand U14490 (N_14490,N_13651,N_13070);
nor U14491 (N_14491,N_13097,N_13484);
nand U14492 (N_14492,N_13860,N_13022);
or U14493 (N_14493,N_13632,N_13079);
and U14494 (N_14494,N_13966,N_13672);
nand U14495 (N_14495,N_13432,N_13589);
or U14496 (N_14496,N_13952,N_13569);
and U14497 (N_14497,N_13451,N_13603);
and U14498 (N_14498,N_13831,N_13946);
nor U14499 (N_14499,N_13282,N_13996);
and U14500 (N_14500,N_13476,N_13503);
or U14501 (N_14501,N_13129,N_13249);
nor U14502 (N_14502,N_13800,N_13240);
or U14503 (N_14503,N_13765,N_13806);
and U14504 (N_14504,N_13453,N_13324);
and U14505 (N_14505,N_13581,N_13659);
xor U14506 (N_14506,N_13672,N_13617);
and U14507 (N_14507,N_13595,N_13588);
or U14508 (N_14508,N_13817,N_13754);
nand U14509 (N_14509,N_13983,N_13325);
and U14510 (N_14510,N_13560,N_13414);
xnor U14511 (N_14511,N_13489,N_13986);
nand U14512 (N_14512,N_13854,N_13616);
and U14513 (N_14513,N_13360,N_13083);
and U14514 (N_14514,N_13834,N_13125);
xnor U14515 (N_14515,N_13037,N_13430);
or U14516 (N_14516,N_13889,N_13538);
xor U14517 (N_14517,N_13363,N_13663);
nand U14518 (N_14518,N_13783,N_13620);
or U14519 (N_14519,N_13698,N_13324);
nand U14520 (N_14520,N_13061,N_13661);
nor U14521 (N_14521,N_13680,N_13435);
and U14522 (N_14522,N_13325,N_13111);
nor U14523 (N_14523,N_13615,N_13874);
or U14524 (N_14524,N_13704,N_13958);
nor U14525 (N_14525,N_13727,N_13269);
nor U14526 (N_14526,N_13902,N_13674);
or U14527 (N_14527,N_13663,N_13684);
xor U14528 (N_14528,N_13089,N_13118);
nand U14529 (N_14529,N_13030,N_13306);
nor U14530 (N_14530,N_13677,N_13697);
nor U14531 (N_14531,N_13769,N_13069);
xnor U14532 (N_14532,N_13945,N_13359);
nor U14533 (N_14533,N_13762,N_13085);
or U14534 (N_14534,N_13489,N_13557);
xnor U14535 (N_14535,N_13458,N_13463);
xor U14536 (N_14536,N_13887,N_13090);
nand U14537 (N_14537,N_13922,N_13794);
xnor U14538 (N_14538,N_13546,N_13787);
and U14539 (N_14539,N_13810,N_13040);
nor U14540 (N_14540,N_13847,N_13923);
or U14541 (N_14541,N_13690,N_13359);
or U14542 (N_14542,N_13580,N_13597);
xor U14543 (N_14543,N_13220,N_13200);
nand U14544 (N_14544,N_13474,N_13961);
and U14545 (N_14545,N_13837,N_13356);
and U14546 (N_14546,N_13548,N_13926);
xor U14547 (N_14547,N_13572,N_13294);
nand U14548 (N_14548,N_13554,N_13764);
and U14549 (N_14549,N_13555,N_13500);
xor U14550 (N_14550,N_13026,N_13333);
and U14551 (N_14551,N_13334,N_13551);
nand U14552 (N_14552,N_13736,N_13668);
xnor U14553 (N_14553,N_13372,N_13299);
and U14554 (N_14554,N_13059,N_13925);
and U14555 (N_14555,N_13648,N_13557);
xnor U14556 (N_14556,N_13270,N_13318);
nand U14557 (N_14557,N_13992,N_13398);
xnor U14558 (N_14558,N_13158,N_13262);
nand U14559 (N_14559,N_13078,N_13465);
nor U14560 (N_14560,N_13231,N_13338);
nand U14561 (N_14561,N_13731,N_13866);
xor U14562 (N_14562,N_13537,N_13604);
and U14563 (N_14563,N_13502,N_13037);
or U14564 (N_14564,N_13693,N_13999);
xnor U14565 (N_14565,N_13810,N_13018);
xnor U14566 (N_14566,N_13291,N_13218);
nand U14567 (N_14567,N_13461,N_13753);
nand U14568 (N_14568,N_13245,N_13355);
nor U14569 (N_14569,N_13803,N_13109);
nand U14570 (N_14570,N_13422,N_13242);
xnor U14571 (N_14571,N_13615,N_13136);
or U14572 (N_14572,N_13798,N_13005);
nor U14573 (N_14573,N_13981,N_13515);
xnor U14574 (N_14574,N_13913,N_13799);
or U14575 (N_14575,N_13487,N_13483);
and U14576 (N_14576,N_13293,N_13673);
nor U14577 (N_14577,N_13929,N_13008);
and U14578 (N_14578,N_13457,N_13182);
and U14579 (N_14579,N_13245,N_13814);
and U14580 (N_14580,N_13248,N_13903);
and U14581 (N_14581,N_13305,N_13302);
nor U14582 (N_14582,N_13614,N_13314);
nor U14583 (N_14583,N_13595,N_13426);
and U14584 (N_14584,N_13362,N_13959);
nand U14585 (N_14585,N_13411,N_13800);
and U14586 (N_14586,N_13475,N_13214);
and U14587 (N_14587,N_13655,N_13003);
and U14588 (N_14588,N_13606,N_13130);
xnor U14589 (N_14589,N_13941,N_13276);
or U14590 (N_14590,N_13881,N_13982);
nor U14591 (N_14591,N_13470,N_13599);
nor U14592 (N_14592,N_13889,N_13674);
nor U14593 (N_14593,N_13183,N_13359);
nor U14594 (N_14594,N_13974,N_13558);
nor U14595 (N_14595,N_13419,N_13485);
nand U14596 (N_14596,N_13200,N_13920);
nor U14597 (N_14597,N_13691,N_13170);
xnor U14598 (N_14598,N_13981,N_13386);
nand U14599 (N_14599,N_13255,N_13822);
or U14600 (N_14600,N_13553,N_13676);
nor U14601 (N_14601,N_13413,N_13077);
nor U14602 (N_14602,N_13622,N_13188);
nand U14603 (N_14603,N_13265,N_13191);
nand U14604 (N_14604,N_13892,N_13861);
nand U14605 (N_14605,N_13195,N_13282);
xor U14606 (N_14606,N_13729,N_13427);
or U14607 (N_14607,N_13661,N_13885);
nor U14608 (N_14608,N_13601,N_13947);
or U14609 (N_14609,N_13494,N_13275);
nor U14610 (N_14610,N_13289,N_13084);
and U14611 (N_14611,N_13414,N_13562);
and U14612 (N_14612,N_13750,N_13766);
nor U14613 (N_14613,N_13629,N_13495);
nor U14614 (N_14614,N_13338,N_13113);
xor U14615 (N_14615,N_13175,N_13646);
and U14616 (N_14616,N_13015,N_13686);
nor U14617 (N_14617,N_13810,N_13223);
or U14618 (N_14618,N_13886,N_13632);
xnor U14619 (N_14619,N_13057,N_13312);
and U14620 (N_14620,N_13009,N_13954);
nor U14621 (N_14621,N_13961,N_13339);
nor U14622 (N_14622,N_13576,N_13613);
nor U14623 (N_14623,N_13708,N_13801);
and U14624 (N_14624,N_13812,N_13286);
or U14625 (N_14625,N_13583,N_13242);
xnor U14626 (N_14626,N_13393,N_13129);
and U14627 (N_14627,N_13743,N_13505);
nor U14628 (N_14628,N_13559,N_13949);
nor U14629 (N_14629,N_13637,N_13106);
nand U14630 (N_14630,N_13518,N_13999);
nand U14631 (N_14631,N_13447,N_13458);
or U14632 (N_14632,N_13302,N_13026);
xor U14633 (N_14633,N_13698,N_13218);
xor U14634 (N_14634,N_13030,N_13826);
xnor U14635 (N_14635,N_13155,N_13574);
or U14636 (N_14636,N_13191,N_13881);
nor U14637 (N_14637,N_13263,N_13964);
nor U14638 (N_14638,N_13061,N_13743);
nand U14639 (N_14639,N_13152,N_13687);
nand U14640 (N_14640,N_13439,N_13667);
nor U14641 (N_14641,N_13495,N_13692);
nand U14642 (N_14642,N_13776,N_13613);
and U14643 (N_14643,N_13389,N_13403);
and U14644 (N_14644,N_13916,N_13182);
nand U14645 (N_14645,N_13265,N_13890);
xor U14646 (N_14646,N_13107,N_13554);
xnor U14647 (N_14647,N_13071,N_13360);
nand U14648 (N_14648,N_13956,N_13236);
xnor U14649 (N_14649,N_13583,N_13377);
and U14650 (N_14650,N_13037,N_13459);
nor U14651 (N_14651,N_13972,N_13352);
nor U14652 (N_14652,N_13310,N_13645);
xnor U14653 (N_14653,N_13902,N_13189);
or U14654 (N_14654,N_13420,N_13671);
xnor U14655 (N_14655,N_13663,N_13704);
nand U14656 (N_14656,N_13290,N_13087);
and U14657 (N_14657,N_13089,N_13682);
xor U14658 (N_14658,N_13996,N_13470);
nand U14659 (N_14659,N_13877,N_13823);
nor U14660 (N_14660,N_13210,N_13487);
and U14661 (N_14661,N_13313,N_13722);
nand U14662 (N_14662,N_13612,N_13623);
nand U14663 (N_14663,N_13976,N_13493);
and U14664 (N_14664,N_13651,N_13006);
and U14665 (N_14665,N_13996,N_13712);
and U14666 (N_14666,N_13876,N_13594);
or U14667 (N_14667,N_13116,N_13890);
or U14668 (N_14668,N_13458,N_13517);
or U14669 (N_14669,N_13545,N_13155);
or U14670 (N_14670,N_13639,N_13208);
nand U14671 (N_14671,N_13020,N_13106);
xnor U14672 (N_14672,N_13559,N_13197);
xnor U14673 (N_14673,N_13220,N_13162);
and U14674 (N_14674,N_13642,N_13176);
or U14675 (N_14675,N_13521,N_13106);
nand U14676 (N_14676,N_13301,N_13233);
or U14677 (N_14677,N_13926,N_13017);
xnor U14678 (N_14678,N_13916,N_13657);
nand U14679 (N_14679,N_13025,N_13605);
and U14680 (N_14680,N_13943,N_13274);
and U14681 (N_14681,N_13678,N_13892);
nor U14682 (N_14682,N_13925,N_13711);
nand U14683 (N_14683,N_13701,N_13558);
and U14684 (N_14684,N_13056,N_13556);
nor U14685 (N_14685,N_13231,N_13737);
and U14686 (N_14686,N_13356,N_13250);
or U14687 (N_14687,N_13528,N_13297);
and U14688 (N_14688,N_13473,N_13024);
nand U14689 (N_14689,N_13765,N_13115);
nor U14690 (N_14690,N_13287,N_13808);
nor U14691 (N_14691,N_13695,N_13365);
nor U14692 (N_14692,N_13689,N_13656);
nand U14693 (N_14693,N_13377,N_13746);
nor U14694 (N_14694,N_13343,N_13379);
xnor U14695 (N_14695,N_13071,N_13990);
xnor U14696 (N_14696,N_13084,N_13862);
nor U14697 (N_14697,N_13837,N_13281);
nor U14698 (N_14698,N_13839,N_13682);
or U14699 (N_14699,N_13431,N_13039);
and U14700 (N_14700,N_13971,N_13349);
or U14701 (N_14701,N_13680,N_13333);
or U14702 (N_14702,N_13157,N_13484);
nor U14703 (N_14703,N_13771,N_13197);
or U14704 (N_14704,N_13621,N_13676);
or U14705 (N_14705,N_13306,N_13292);
nor U14706 (N_14706,N_13005,N_13413);
xnor U14707 (N_14707,N_13220,N_13941);
nor U14708 (N_14708,N_13941,N_13380);
nand U14709 (N_14709,N_13421,N_13361);
and U14710 (N_14710,N_13436,N_13522);
nor U14711 (N_14711,N_13599,N_13531);
and U14712 (N_14712,N_13104,N_13622);
nor U14713 (N_14713,N_13797,N_13630);
or U14714 (N_14714,N_13808,N_13513);
nand U14715 (N_14715,N_13925,N_13801);
and U14716 (N_14716,N_13887,N_13312);
nor U14717 (N_14717,N_13254,N_13427);
nor U14718 (N_14718,N_13138,N_13319);
nor U14719 (N_14719,N_13340,N_13513);
and U14720 (N_14720,N_13626,N_13958);
and U14721 (N_14721,N_13338,N_13417);
nand U14722 (N_14722,N_13724,N_13776);
or U14723 (N_14723,N_13223,N_13395);
or U14724 (N_14724,N_13239,N_13177);
and U14725 (N_14725,N_13922,N_13861);
xnor U14726 (N_14726,N_13896,N_13865);
and U14727 (N_14727,N_13576,N_13668);
or U14728 (N_14728,N_13081,N_13331);
nand U14729 (N_14729,N_13077,N_13292);
or U14730 (N_14730,N_13236,N_13634);
or U14731 (N_14731,N_13803,N_13402);
and U14732 (N_14732,N_13501,N_13444);
or U14733 (N_14733,N_13348,N_13520);
nor U14734 (N_14734,N_13330,N_13596);
nor U14735 (N_14735,N_13468,N_13844);
xnor U14736 (N_14736,N_13777,N_13336);
or U14737 (N_14737,N_13565,N_13805);
and U14738 (N_14738,N_13743,N_13991);
or U14739 (N_14739,N_13214,N_13788);
xnor U14740 (N_14740,N_13318,N_13300);
or U14741 (N_14741,N_13031,N_13931);
xnor U14742 (N_14742,N_13399,N_13101);
or U14743 (N_14743,N_13860,N_13566);
nand U14744 (N_14744,N_13252,N_13101);
and U14745 (N_14745,N_13894,N_13514);
nand U14746 (N_14746,N_13002,N_13525);
xor U14747 (N_14747,N_13546,N_13784);
nor U14748 (N_14748,N_13871,N_13187);
or U14749 (N_14749,N_13865,N_13116);
xnor U14750 (N_14750,N_13185,N_13071);
nand U14751 (N_14751,N_13935,N_13971);
nand U14752 (N_14752,N_13279,N_13744);
or U14753 (N_14753,N_13562,N_13621);
and U14754 (N_14754,N_13778,N_13238);
xnor U14755 (N_14755,N_13889,N_13083);
nor U14756 (N_14756,N_13174,N_13235);
and U14757 (N_14757,N_13031,N_13368);
or U14758 (N_14758,N_13813,N_13917);
nand U14759 (N_14759,N_13767,N_13901);
xnor U14760 (N_14760,N_13438,N_13531);
and U14761 (N_14761,N_13268,N_13489);
and U14762 (N_14762,N_13697,N_13172);
and U14763 (N_14763,N_13147,N_13762);
and U14764 (N_14764,N_13319,N_13565);
or U14765 (N_14765,N_13037,N_13619);
xnor U14766 (N_14766,N_13511,N_13166);
nor U14767 (N_14767,N_13495,N_13524);
nand U14768 (N_14768,N_13052,N_13445);
or U14769 (N_14769,N_13181,N_13797);
nor U14770 (N_14770,N_13608,N_13846);
nor U14771 (N_14771,N_13385,N_13957);
xnor U14772 (N_14772,N_13825,N_13595);
and U14773 (N_14773,N_13918,N_13311);
nand U14774 (N_14774,N_13437,N_13075);
or U14775 (N_14775,N_13424,N_13254);
or U14776 (N_14776,N_13545,N_13435);
nand U14777 (N_14777,N_13831,N_13726);
and U14778 (N_14778,N_13625,N_13586);
or U14779 (N_14779,N_13257,N_13595);
xor U14780 (N_14780,N_13066,N_13194);
nor U14781 (N_14781,N_13492,N_13171);
and U14782 (N_14782,N_13164,N_13569);
nor U14783 (N_14783,N_13597,N_13761);
or U14784 (N_14784,N_13374,N_13635);
or U14785 (N_14785,N_13970,N_13194);
nand U14786 (N_14786,N_13805,N_13638);
nand U14787 (N_14787,N_13202,N_13006);
or U14788 (N_14788,N_13167,N_13914);
nand U14789 (N_14789,N_13219,N_13131);
nor U14790 (N_14790,N_13606,N_13817);
or U14791 (N_14791,N_13101,N_13086);
or U14792 (N_14792,N_13410,N_13123);
nor U14793 (N_14793,N_13967,N_13890);
xor U14794 (N_14794,N_13013,N_13496);
nor U14795 (N_14795,N_13512,N_13345);
nor U14796 (N_14796,N_13265,N_13776);
or U14797 (N_14797,N_13191,N_13949);
or U14798 (N_14798,N_13382,N_13460);
xnor U14799 (N_14799,N_13879,N_13740);
and U14800 (N_14800,N_13510,N_13444);
nor U14801 (N_14801,N_13463,N_13959);
nor U14802 (N_14802,N_13240,N_13074);
and U14803 (N_14803,N_13734,N_13640);
nor U14804 (N_14804,N_13549,N_13050);
or U14805 (N_14805,N_13641,N_13819);
nor U14806 (N_14806,N_13803,N_13185);
and U14807 (N_14807,N_13345,N_13310);
xnor U14808 (N_14808,N_13570,N_13773);
xor U14809 (N_14809,N_13293,N_13302);
xor U14810 (N_14810,N_13779,N_13087);
nand U14811 (N_14811,N_13710,N_13483);
and U14812 (N_14812,N_13248,N_13765);
and U14813 (N_14813,N_13372,N_13441);
xor U14814 (N_14814,N_13827,N_13703);
nor U14815 (N_14815,N_13836,N_13389);
xor U14816 (N_14816,N_13502,N_13938);
nand U14817 (N_14817,N_13472,N_13913);
xnor U14818 (N_14818,N_13876,N_13247);
and U14819 (N_14819,N_13636,N_13629);
or U14820 (N_14820,N_13853,N_13054);
xnor U14821 (N_14821,N_13168,N_13928);
or U14822 (N_14822,N_13164,N_13901);
or U14823 (N_14823,N_13099,N_13591);
xor U14824 (N_14824,N_13426,N_13428);
or U14825 (N_14825,N_13662,N_13611);
or U14826 (N_14826,N_13968,N_13962);
or U14827 (N_14827,N_13600,N_13545);
and U14828 (N_14828,N_13665,N_13693);
or U14829 (N_14829,N_13388,N_13643);
nand U14830 (N_14830,N_13391,N_13489);
nor U14831 (N_14831,N_13194,N_13244);
nor U14832 (N_14832,N_13419,N_13810);
xnor U14833 (N_14833,N_13129,N_13906);
nor U14834 (N_14834,N_13724,N_13382);
and U14835 (N_14835,N_13268,N_13704);
nand U14836 (N_14836,N_13341,N_13961);
or U14837 (N_14837,N_13496,N_13288);
nor U14838 (N_14838,N_13268,N_13235);
nor U14839 (N_14839,N_13929,N_13925);
and U14840 (N_14840,N_13135,N_13352);
nand U14841 (N_14841,N_13056,N_13716);
and U14842 (N_14842,N_13082,N_13962);
xnor U14843 (N_14843,N_13976,N_13756);
or U14844 (N_14844,N_13938,N_13826);
or U14845 (N_14845,N_13131,N_13539);
xor U14846 (N_14846,N_13361,N_13688);
nor U14847 (N_14847,N_13200,N_13995);
and U14848 (N_14848,N_13067,N_13257);
nand U14849 (N_14849,N_13121,N_13853);
nand U14850 (N_14850,N_13068,N_13654);
or U14851 (N_14851,N_13446,N_13071);
and U14852 (N_14852,N_13286,N_13461);
nand U14853 (N_14853,N_13987,N_13371);
xnor U14854 (N_14854,N_13779,N_13700);
nor U14855 (N_14855,N_13524,N_13702);
or U14856 (N_14856,N_13184,N_13648);
and U14857 (N_14857,N_13494,N_13390);
nand U14858 (N_14858,N_13165,N_13169);
nand U14859 (N_14859,N_13116,N_13319);
nand U14860 (N_14860,N_13646,N_13161);
xnor U14861 (N_14861,N_13615,N_13375);
and U14862 (N_14862,N_13737,N_13563);
nand U14863 (N_14863,N_13272,N_13927);
nand U14864 (N_14864,N_13504,N_13263);
and U14865 (N_14865,N_13639,N_13655);
xor U14866 (N_14866,N_13776,N_13028);
or U14867 (N_14867,N_13705,N_13313);
xor U14868 (N_14868,N_13619,N_13402);
nand U14869 (N_14869,N_13877,N_13644);
and U14870 (N_14870,N_13353,N_13516);
nand U14871 (N_14871,N_13344,N_13395);
xnor U14872 (N_14872,N_13873,N_13781);
nor U14873 (N_14873,N_13149,N_13112);
nor U14874 (N_14874,N_13852,N_13192);
and U14875 (N_14875,N_13499,N_13204);
and U14876 (N_14876,N_13605,N_13913);
nand U14877 (N_14877,N_13388,N_13986);
and U14878 (N_14878,N_13144,N_13216);
or U14879 (N_14879,N_13321,N_13930);
xnor U14880 (N_14880,N_13066,N_13769);
nor U14881 (N_14881,N_13318,N_13331);
nand U14882 (N_14882,N_13942,N_13730);
or U14883 (N_14883,N_13121,N_13343);
nor U14884 (N_14884,N_13314,N_13709);
xor U14885 (N_14885,N_13817,N_13360);
nor U14886 (N_14886,N_13551,N_13994);
and U14887 (N_14887,N_13101,N_13894);
and U14888 (N_14888,N_13502,N_13644);
nor U14889 (N_14889,N_13127,N_13573);
xnor U14890 (N_14890,N_13375,N_13331);
nor U14891 (N_14891,N_13786,N_13356);
xnor U14892 (N_14892,N_13206,N_13784);
nor U14893 (N_14893,N_13499,N_13224);
nor U14894 (N_14894,N_13151,N_13351);
nand U14895 (N_14895,N_13830,N_13777);
nand U14896 (N_14896,N_13073,N_13691);
and U14897 (N_14897,N_13114,N_13834);
and U14898 (N_14898,N_13796,N_13710);
xor U14899 (N_14899,N_13774,N_13868);
nor U14900 (N_14900,N_13799,N_13159);
or U14901 (N_14901,N_13897,N_13953);
and U14902 (N_14902,N_13527,N_13247);
and U14903 (N_14903,N_13864,N_13860);
nand U14904 (N_14904,N_13503,N_13235);
nor U14905 (N_14905,N_13814,N_13115);
nor U14906 (N_14906,N_13108,N_13991);
nor U14907 (N_14907,N_13998,N_13315);
or U14908 (N_14908,N_13295,N_13012);
nor U14909 (N_14909,N_13754,N_13524);
xor U14910 (N_14910,N_13329,N_13503);
nor U14911 (N_14911,N_13213,N_13751);
nor U14912 (N_14912,N_13017,N_13768);
nand U14913 (N_14913,N_13185,N_13395);
nand U14914 (N_14914,N_13453,N_13415);
nand U14915 (N_14915,N_13410,N_13318);
xor U14916 (N_14916,N_13192,N_13452);
and U14917 (N_14917,N_13839,N_13352);
xnor U14918 (N_14918,N_13437,N_13274);
nand U14919 (N_14919,N_13974,N_13014);
or U14920 (N_14920,N_13868,N_13326);
nand U14921 (N_14921,N_13049,N_13965);
nor U14922 (N_14922,N_13377,N_13317);
and U14923 (N_14923,N_13365,N_13927);
xor U14924 (N_14924,N_13930,N_13848);
and U14925 (N_14925,N_13428,N_13917);
nand U14926 (N_14926,N_13175,N_13891);
xnor U14927 (N_14927,N_13567,N_13258);
or U14928 (N_14928,N_13420,N_13715);
nor U14929 (N_14929,N_13441,N_13567);
or U14930 (N_14930,N_13876,N_13120);
and U14931 (N_14931,N_13543,N_13455);
nor U14932 (N_14932,N_13116,N_13326);
xor U14933 (N_14933,N_13441,N_13444);
nor U14934 (N_14934,N_13252,N_13386);
nor U14935 (N_14935,N_13065,N_13745);
xor U14936 (N_14936,N_13652,N_13713);
and U14937 (N_14937,N_13093,N_13627);
nand U14938 (N_14938,N_13612,N_13626);
and U14939 (N_14939,N_13401,N_13777);
and U14940 (N_14940,N_13933,N_13354);
nor U14941 (N_14941,N_13597,N_13787);
nand U14942 (N_14942,N_13058,N_13323);
xor U14943 (N_14943,N_13351,N_13663);
and U14944 (N_14944,N_13324,N_13998);
xor U14945 (N_14945,N_13713,N_13024);
nor U14946 (N_14946,N_13751,N_13139);
xor U14947 (N_14947,N_13582,N_13884);
and U14948 (N_14948,N_13305,N_13836);
nor U14949 (N_14949,N_13622,N_13471);
nand U14950 (N_14950,N_13580,N_13893);
nor U14951 (N_14951,N_13308,N_13109);
nor U14952 (N_14952,N_13339,N_13003);
nor U14953 (N_14953,N_13423,N_13437);
nor U14954 (N_14954,N_13708,N_13849);
and U14955 (N_14955,N_13156,N_13088);
nor U14956 (N_14956,N_13218,N_13239);
xnor U14957 (N_14957,N_13577,N_13505);
xnor U14958 (N_14958,N_13820,N_13227);
nand U14959 (N_14959,N_13687,N_13866);
and U14960 (N_14960,N_13999,N_13724);
xor U14961 (N_14961,N_13822,N_13956);
xnor U14962 (N_14962,N_13560,N_13800);
nand U14963 (N_14963,N_13564,N_13794);
nand U14964 (N_14964,N_13910,N_13132);
xor U14965 (N_14965,N_13294,N_13507);
nor U14966 (N_14966,N_13993,N_13711);
nor U14967 (N_14967,N_13431,N_13002);
and U14968 (N_14968,N_13523,N_13153);
nor U14969 (N_14969,N_13085,N_13113);
nor U14970 (N_14970,N_13082,N_13802);
or U14971 (N_14971,N_13536,N_13092);
xnor U14972 (N_14972,N_13480,N_13886);
or U14973 (N_14973,N_13965,N_13426);
or U14974 (N_14974,N_13287,N_13417);
nor U14975 (N_14975,N_13263,N_13857);
nand U14976 (N_14976,N_13987,N_13857);
nand U14977 (N_14977,N_13512,N_13895);
and U14978 (N_14978,N_13059,N_13747);
nor U14979 (N_14979,N_13534,N_13005);
and U14980 (N_14980,N_13831,N_13987);
xnor U14981 (N_14981,N_13497,N_13872);
xnor U14982 (N_14982,N_13360,N_13233);
nand U14983 (N_14983,N_13401,N_13904);
or U14984 (N_14984,N_13618,N_13334);
nand U14985 (N_14985,N_13227,N_13279);
nor U14986 (N_14986,N_13437,N_13229);
nand U14987 (N_14987,N_13021,N_13759);
or U14988 (N_14988,N_13473,N_13791);
nor U14989 (N_14989,N_13797,N_13948);
and U14990 (N_14990,N_13091,N_13718);
xnor U14991 (N_14991,N_13279,N_13609);
nand U14992 (N_14992,N_13591,N_13959);
and U14993 (N_14993,N_13258,N_13745);
xor U14994 (N_14994,N_13661,N_13269);
or U14995 (N_14995,N_13754,N_13809);
nor U14996 (N_14996,N_13931,N_13520);
nand U14997 (N_14997,N_13786,N_13571);
nand U14998 (N_14998,N_13152,N_13498);
xor U14999 (N_14999,N_13522,N_13495);
and U15000 (N_15000,N_14303,N_14484);
nand U15001 (N_15001,N_14243,N_14857);
or U15002 (N_15002,N_14277,N_14301);
nor U15003 (N_15003,N_14178,N_14693);
nor U15004 (N_15004,N_14330,N_14069);
nor U15005 (N_15005,N_14519,N_14692);
nand U15006 (N_15006,N_14023,N_14767);
or U15007 (N_15007,N_14597,N_14559);
nand U15008 (N_15008,N_14455,N_14502);
xor U15009 (N_15009,N_14247,N_14921);
xor U15010 (N_15010,N_14124,N_14111);
nand U15011 (N_15011,N_14932,N_14497);
nand U15012 (N_15012,N_14593,N_14479);
and U15013 (N_15013,N_14035,N_14586);
xnor U15014 (N_15014,N_14245,N_14065);
and U15015 (N_15015,N_14831,N_14092);
and U15016 (N_15016,N_14902,N_14450);
nand U15017 (N_15017,N_14527,N_14575);
and U15018 (N_15018,N_14025,N_14553);
or U15019 (N_15019,N_14337,N_14003);
nor U15020 (N_15020,N_14581,N_14231);
or U15021 (N_15021,N_14253,N_14409);
xor U15022 (N_15022,N_14151,N_14079);
nand U15023 (N_15023,N_14207,N_14220);
and U15024 (N_15024,N_14747,N_14421);
or U15025 (N_15025,N_14934,N_14127);
nor U15026 (N_15026,N_14839,N_14280);
and U15027 (N_15027,N_14856,N_14953);
xnor U15028 (N_15028,N_14100,N_14487);
xnor U15029 (N_15029,N_14238,N_14590);
or U15030 (N_15030,N_14371,N_14798);
nor U15031 (N_15031,N_14477,N_14877);
or U15032 (N_15032,N_14478,N_14211);
or U15033 (N_15033,N_14853,N_14293);
and U15034 (N_15034,N_14420,N_14465);
or U15035 (N_15035,N_14287,N_14602);
nor U15036 (N_15036,N_14439,N_14369);
nor U15037 (N_15037,N_14876,N_14355);
or U15038 (N_15038,N_14153,N_14097);
and U15039 (N_15039,N_14144,N_14683);
nor U15040 (N_15040,N_14807,N_14631);
or U15041 (N_15041,N_14748,N_14070);
and U15042 (N_15042,N_14942,N_14263);
or U15043 (N_15043,N_14077,N_14691);
xor U15044 (N_15044,N_14805,N_14222);
and U15045 (N_15045,N_14407,N_14979);
and U15046 (N_15046,N_14598,N_14982);
nand U15047 (N_15047,N_14679,N_14733);
nand U15048 (N_15048,N_14370,N_14970);
or U15049 (N_15049,N_14816,N_14917);
and U15050 (N_15050,N_14348,N_14269);
and U15051 (N_15051,N_14678,N_14435);
xnor U15052 (N_15052,N_14039,N_14061);
nand U15053 (N_15053,N_14154,N_14017);
and U15054 (N_15054,N_14570,N_14592);
nand U15055 (N_15055,N_14517,N_14083);
nand U15056 (N_15056,N_14694,N_14413);
and U15057 (N_15057,N_14509,N_14635);
and U15058 (N_15058,N_14501,N_14166);
nor U15059 (N_15059,N_14168,N_14430);
and U15060 (N_15060,N_14295,N_14366);
and U15061 (N_15061,N_14344,N_14399);
or U15062 (N_15062,N_14612,N_14562);
or U15063 (N_15063,N_14302,N_14974);
nand U15064 (N_15064,N_14233,N_14545);
nor U15065 (N_15065,N_14028,N_14822);
xor U15066 (N_15066,N_14493,N_14904);
and U15067 (N_15067,N_14888,N_14076);
nand U15068 (N_15068,N_14216,N_14062);
and U15069 (N_15069,N_14684,N_14986);
or U15070 (N_15070,N_14647,N_14195);
nand U15071 (N_15071,N_14452,N_14563);
and U15072 (N_15072,N_14905,N_14812);
xnor U15073 (N_15073,N_14160,N_14432);
xor U15074 (N_15074,N_14368,N_14008);
nand U15075 (N_15075,N_14978,N_14254);
xnor U15076 (N_15076,N_14043,N_14235);
or U15077 (N_15077,N_14383,N_14965);
nand U15078 (N_15078,N_14447,N_14862);
and U15079 (N_15079,N_14543,N_14882);
and U15080 (N_15080,N_14580,N_14848);
and U15081 (N_15081,N_14777,N_14595);
nor U15082 (N_15082,N_14380,N_14504);
xor U15083 (N_15083,N_14304,N_14041);
nand U15084 (N_15084,N_14448,N_14194);
xor U15085 (N_15085,N_14164,N_14989);
nand U15086 (N_15086,N_14030,N_14653);
nand U15087 (N_15087,N_14252,N_14619);
and U15088 (N_15088,N_14406,N_14012);
nor U15089 (N_15089,N_14819,N_14672);
and U15090 (N_15090,N_14896,N_14997);
or U15091 (N_15091,N_14388,N_14603);
nor U15092 (N_15092,N_14342,N_14656);
nand U15093 (N_15093,N_14762,N_14387);
nand U15094 (N_15094,N_14664,N_14485);
nor U15095 (N_15095,N_14481,N_14845);
and U15096 (N_15096,N_14667,N_14248);
and U15097 (N_15097,N_14752,N_14072);
or U15098 (N_15098,N_14507,N_14713);
nand U15099 (N_15099,N_14405,N_14270);
and U15100 (N_15100,N_14670,N_14494);
or U15101 (N_15101,N_14868,N_14512);
nand U15102 (N_15102,N_14305,N_14101);
xnor U15103 (N_15103,N_14734,N_14751);
nand U15104 (N_15104,N_14939,N_14992);
xor U15105 (N_15105,N_14849,N_14806);
or U15106 (N_15106,N_14310,N_14701);
nand U15107 (N_15107,N_14114,N_14537);
and U15108 (N_15108,N_14396,N_14923);
and U15109 (N_15109,N_14063,N_14514);
nor U15110 (N_15110,N_14459,N_14362);
nor U15111 (N_15111,N_14789,N_14741);
and U15112 (N_15112,N_14056,N_14909);
or U15113 (N_15113,N_14224,N_14709);
and U15114 (N_15114,N_14521,N_14040);
xnor U15115 (N_15115,N_14843,N_14754);
nand U15116 (N_15116,N_14073,N_14900);
nor U15117 (N_15117,N_14744,N_14760);
and U15118 (N_15118,N_14985,N_14662);
and U15119 (N_15119,N_14089,N_14984);
nand U15120 (N_15120,N_14384,N_14577);
xor U15121 (N_15121,N_14453,N_14400);
or U15122 (N_15122,N_14281,N_14784);
nand U15123 (N_15123,N_14532,N_14214);
and U15124 (N_15124,N_14050,N_14356);
or U15125 (N_15125,N_14795,N_14067);
nand U15126 (N_15126,N_14774,N_14139);
and U15127 (N_15127,N_14312,N_14548);
or U15128 (N_15128,N_14429,N_14628);
nor U15129 (N_15129,N_14555,N_14964);
nor U15130 (N_15130,N_14492,N_14772);
and U15131 (N_15131,N_14021,N_14033);
xor U15132 (N_15132,N_14520,N_14757);
nor U15133 (N_15133,N_14606,N_14438);
and U15134 (N_15134,N_14443,N_14726);
nand U15135 (N_15135,N_14018,N_14542);
nor U15136 (N_15136,N_14239,N_14594);
and U15137 (N_15137,N_14945,N_14549);
or U15138 (N_15138,N_14206,N_14949);
or U15139 (N_15139,N_14957,N_14172);
nand U15140 (N_15140,N_14865,N_14193);
xnor U15141 (N_15141,N_14201,N_14320);
xnor U15142 (N_15142,N_14085,N_14522);
or U15143 (N_15143,N_14715,N_14722);
nand U15144 (N_15144,N_14599,N_14758);
or U15145 (N_15145,N_14325,N_14968);
or U15146 (N_15146,N_14318,N_14861);
or U15147 (N_15147,N_14686,N_14756);
nor U15148 (N_15148,N_14274,N_14668);
nand U15149 (N_15149,N_14218,N_14219);
or U15150 (N_15150,N_14319,N_14081);
nand U15151 (N_15151,N_14551,N_14914);
and U15152 (N_15152,N_14908,N_14048);
or U15153 (N_15153,N_14611,N_14288);
xnor U15154 (N_15154,N_14915,N_14711);
nand U15155 (N_15155,N_14350,N_14931);
or U15156 (N_15156,N_14136,N_14966);
nor U15157 (N_15157,N_14360,N_14657);
nand U15158 (N_15158,N_14027,N_14632);
xor U15159 (N_15159,N_14740,N_14137);
or U15160 (N_15160,N_14426,N_14375);
nand U15161 (N_15161,N_14335,N_14437);
or U15162 (N_15162,N_14860,N_14490);
or U15163 (N_15163,N_14541,N_14394);
or U15164 (N_15164,N_14296,N_14090);
or U15165 (N_15165,N_14649,N_14156);
or U15166 (N_15166,N_14317,N_14180);
nand U15167 (N_15167,N_14674,N_14422);
and U15168 (N_15168,N_14122,N_14676);
nand U15169 (N_15169,N_14941,N_14257);
and U15170 (N_15170,N_14859,N_14907);
nor U15171 (N_15171,N_14531,N_14183);
and U15172 (N_15172,N_14182,N_14376);
nand U15173 (N_15173,N_14621,N_14442);
and U15174 (N_15174,N_14217,N_14585);
nand U15175 (N_15175,N_14561,N_14011);
and U15176 (N_15176,N_14334,N_14140);
and U15177 (N_15177,N_14389,N_14044);
xnor U15178 (N_15178,N_14697,N_14624);
nand U15179 (N_15179,N_14835,N_14765);
and U15180 (N_15180,N_14636,N_14724);
xor U15181 (N_15181,N_14264,N_14379);
or U15182 (N_15182,N_14880,N_14745);
xor U15183 (N_15183,N_14866,N_14117);
and U15184 (N_15184,N_14228,N_14052);
nand U15185 (N_15185,N_14644,N_14617);
nor U15186 (N_15186,N_14823,N_14874);
nor U15187 (N_15187,N_14232,N_14457);
nor U15188 (N_15188,N_14495,N_14086);
xor U15189 (N_15189,N_14416,N_14223);
or U15190 (N_15190,N_14605,N_14940);
nor U15191 (N_15191,N_14382,N_14571);
nand U15192 (N_15192,N_14526,N_14212);
and U15193 (N_15193,N_14832,N_14107);
nor U15194 (N_15194,N_14015,N_14339);
and U15195 (N_15195,N_14708,N_14290);
xor U15196 (N_15196,N_14347,N_14392);
and U15197 (N_15197,N_14131,N_14428);
or U15198 (N_15198,N_14273,N_14847);
and U15199 (N_15199,N_14299,N_14503);
and U15200 (N_15200,N_14768,N_14828);
nor U15201 (N_15201,N_14267,N_14630);
and U15202 (N_15202,N_14246,N_14258);
nand U15203 (N_15203,N_14651,N_14129);
nor U15204 (N_15204,N_14262,N_14098);
nor U15205 (N_15205,N_14834,N_14483);
and U15206 (N_15206,N_14471,N_14648);
and U15207 (N_15207,N_14998,N_14564);
and U15208 (N_15208,N_14869,N_14150);
nor U15209 (N_15209,N_14336,N_14391);
nor U15210 (N_15210,N_14118,N_14689);
and U15211 (N_15211,N_14060,N_14759);
nand U15212 (N_15212,N_14738,N_14962);
or U15213 (N_15213,N_14723,N_14002);
and U15214 (N_15214,N_14286,N_14665);
nor U15215 (N_15215,N_14331,N_14746);
or U15216 (N_15216,N_14053,N_14046);
nand U15217 (N_15217,N_14491,N_14196);
nor U15218 (N_15218,N_14547,N_14198);
nor U15219 (N_15219,N_14990,N_14714);
xnor U15220 (N_15220,N_14922,N_14353);
nor U15221 (N_15221,N_14687,N_14627);
nand U15222 (N_15222,N_14121,N_14566);
or U15223 (N_15223,N_14103,N_14778);
or U15224 (N_15224,N_14604,N_14913);
nand U15225 (N_15225,N_14189,N_14016);
xor U15226 (N_15226,N_14327,N_14558);
xor U15227 (N_15227,N_14797,N_14844);
nand U15228 (N_15228,N_14518,N_14276);
nor U15229 (N_15229,N_14059,N_14226);
and U15230 (N_15230,N_14177,N_14538);
nand U15231 (N_15231,N_14176,N_14954);
xor U15232 (N_15232,N_14431,N_14811);
nand U15233 (N_15233,N_14769,N_14725);
and U15234 (N_15234,N_14000,N_14169);
and U15235 (N_15235,N_14074,N_14719);
nor U15236 (N_15236,N_14879,N_14192);
nand U15237 (N_15237,N_14367,N_14316);
or U15238 (N_15238,N_14625,N_14135);
nor U15239 (N_15239,N_14893,N_14474);
or U15240 (N_15240,N_14980,N_14793);
xnor U15241 (N_15241,N_14009,N_14161);
and U15242 (N_15242,N_14326,N_14791);
and U15243 (N_15243,N_14449,N_14550);
or U15244 (N_15244,N_14640,N_14402);
nand U15245 (N_15245,N_14249,N_14582);
xor U15246 (N_15246,N_14434,N_14851);
and U15247 (N_15247,N_14268,N_14956);
nand U15248 (N_15248,N_14799,N_14108);
or U15249 (N_15249,N_14717,N_14162);
or U15250 (N_15250,N_14963,N_14424);
and U15251 (N_15251,N_14814,N_14133);
or U15252 (N_15252,N_14589,N_14467);
nor U15253 (N_15253,N_14781,N_14903);
nor U15254 (N_15254,N_14961,N_14663);
and U15255 (N_15255,N_14846,N_14397);
nand U15256 (N_15256,N_14680,N_14829);
and U15257 (N_15257,N_14842,N_14241);
or U15258 (N_15258,N_14739,N_14933);
or U15259 (N_15259,N_14049,N_14203);
and U15260 (N_15260,N_14324,N_14093);
xnor U15261 (N_15261,N_14813,N_14130);
xor U15262 (N_15262,N_14610,N_14186);
or U15263 (N_15263,N_14138,N_14988);
or U15264 (N_15264,N_14185,N_14250);
and U15265 (N_15265,N_14386,N_14256);
nor U15266 (N_15266,N_14234,N_14584);
xnor U15267 (N_15267,N_14699,N_14489);
or U15268 (N_15268,N_14675,N_14700);
nand U15269 (N_15269,N_14047,N_14261);
and U15270 (N_15270,N_14977,N_14123);
or U15271 (N_15271,N_14889,N_14615);
nand U15272 (N_15272,N_14634,N_14332);
nand U15273 (N_15273,N_14572,N_14125);
and U15274 (N_15274,N_14057,N_14308);
and U15275 (N_15275,N_14006,N_14157);
nor U15276 (N_15276,N_14045,N_14365);
nor U15277 (N_15277,N_14528,N_14706);
or U15278 (N_15278,N_14569,N_14987);
or U15279 (N_15279,N_14535,N_14272);
or U15280 (N_15280,N_14800,N_14445);
and U15281 (N_15281,N_14530,N_14544);
nand U15282 (N_15282,N_14669,N_14929);
or U15283 (N_15283,N_14958,N_14796);
and U15284 (N_15284,N_14613,N_14333);
nand U15285 (N_15285,N_14251,N_14300);
xor U15286 (N_15286,N_14643,N_14973);
nor U15287 (N_15287,N_14529,N_14068);
xor U15288 (N_15288,N_14309,N_14005);
or U15289 (N_15289,N_14322,N_14255);
nor U15290 (N_15290,N_14925,N_14641);
xor U15291 (N_15291,N_14885,N_14788);
nor U15292 (N_15292,N_14480,N_14340);
nor U15293 (N_15293,N_14451,N_14863);
nand U15294 (N_15294,N_14658,N_14213);
nand U15295 (N_15295,N_14034,N_14677);
nor U15296 (N_15296,N_14704,N_14343);
xor U15297 (N_15297,N_14031,N_14080);
xnor U15298 (N_15298,N_14938,N_14568);
nor U15299 (N_15299,N_14901,N_14910);
nor U15300 (N_15300,N_14840,N_14588);
xor U15301 (N_15301,N_14352,N_14583);
nor U15302 (N_15302,N_14596,N_14403);
and U15303 (N_15303,N_14524,N_14496);
xor U15304 (N_15304,N_14415,N_14486);
xnor U15305 (N_15305,N_14463,N_14852);
nor U15306 (N_15306,N_14802,N_14410);
and U15307 (N_15307,N_14533,N_14279);
xor U15308 (N_15308,N_14660,N_14794);
nand U15309 (N_15309,N_14001,N_14505);
or U15310 (N_15310,N_14361,N_14804);
xor U15311 (N_15311,N_14418,N_14064);
or U15312 (N_15312,N_14646,N_14579);
and U15313 (N_15313,N_14109,N_14084);
and U15314 (N_15314,N_14119,N_14513);
and U15315 (N_15315,N_14506,N_14927);
nor U15316 (N_15316,N_14850,N_14082);
nand U15317 (N_15317,N_14508,N_14875);
nor U15318 (N_15318,N_14462,N_14951);
xnor U15319 (N_15319,N_14996,N_14473);
or U15320 (N_15320,N_14833,N_14013);
xnor U15321 (N_15321,N_14237,N_14731);
nand U15322 (N_15322,N_14381,N_14948);
and U15323 (N_15323,N_14094,N_14078);
xnor U15324 (N_15324,N_14995,N_14919);
nand U15325 (N_15325,N_14142,N_14390);
nor U15326 (N_15326,N_14120,N_14215);
and U15327 (N_15327,N_14398,N_14817);
xor U15328 (N_15328,N_14141,N_14600);
or U15329 (N_15329,N_14946,N_14266);
nand U15330 (N_15330,N_14818,N_14753);
xnor U15331 (N_15331,N_14999,N_14099);
and U15332 (N_15332,N_14947,N_14786);
and U15333 (N_15333,N_14766,N_14419);
nor U15334 (N_15334,N_14742,N_14730);
or U15335 (N_15335,N_14688,N_14427);
nor U15336 (N_15336,N_14906,N_14197);
and U15337 (N_15337,N_14042,N_14899);
nand U15338 (N_15338,N_14841,N_14469);
and U15339 (N_15339,N_14510,N_14476);
nand U15340 (N_15340,N_14894,N_14358);
xor U15341 (N_15341,N_14500,N_14696);
nand U15342 (N_15342,N_14878,N_14780);
and U15343 (N_15343,N_14928,N_14695);
or U15344 (N_15344,N_14809,N_14472);
or U15345 (N_15345,N_14618,N_14096);
or U15346 (N_15346,N_14314,N_14468);
nor U15347 (N_15347,N_14897,N_14423);
nor U15348 (N_15348,N_14071,N_14761);
xnor U15349 (N_15349,N_14315,N_14175);
nand U15350 (N_15350,N_14886,N_14773);
xor U15351 (N_15351,N_14411,N_14283);
nor U15352 (N_15352,N_14609,N_14775);
nor U15353 (N_15353,N_14460,N_14208);
xor U15354 (N_15354,N_14626,N_14482);
nor U15355 (N_15355,N_14578,N_14629);
or U15356 (N_15356,N_14075,N_14128);
nor U15357 (N_15357,N_14036,N_14720);
nand U15358 (N_15358,N_14019,N_14952);
or U15359 (N_15359,N_14058,N_14969);
nor U15360 (N_15360,N_14837,N_14158);
xor U15361 (N_15361,N_14149,N_14994);
or U15362 (N_15362,N_14787,N_14095);
nand U15363 (N_15363,N_14464,N_14955);
nand U15364 (N_15364,N_14329,N_14385);
and U15365 (N_15365,N_14191,N_14959);
and U15366 (N_15366,N_14116,N_14622);
and U15367 (N_15367,N_14661,N_14967);
nand U15368 (N_15368,N_14771,N_14895);
and U15369 (N_15369,N_14110,N_14539);
xnor U15370 (N_15370,N_14488,N_14014);
or U15371 (N_15371,N_14446,N_14736);
or U15372 (N_15372,N_14854,N_14858);
nor U15373 (N_15373,N_14440,N_14926);
or U15374 (N_15374,N_14655,N_14716);
nand U15375 (N_15375,N_14587,N_14703);
and U15376 (N_15376,N_14346,N_14637);
or U15377 (N_15377,N_14313,N_14770);
xor U15378 (N_15378,N_14022,N_14971);
xor U15379 (N_15379,N_14685,N_14785);
and U15380 (N_15380,N_14444,N_14032);
nand U15381 (N_15381,N_14912,N_14930);
xor U15382 (N_15382,N_14292,N_14825);
or U15383 (N_15383,N_14810,N_14294);
or U15384 (N_15384,N_14924,N_14475);
xor U15385 (N_15385,N_14433,N_14174);
nand U15386 (N_15386,N_14755,N_14779);
xnor U15387 (N_15387,N_14729,N_14359);
nor U15388 (N_15388,N_14242,N_14827);
nand U15389 (N_15389,N_14323,N_14556);
nor U15390 (N_15390,N_14227,N_14654);
and U15391 (N_15391,N_14782,N_14184);
nand U15392 (N_15392,N_14721,N_14026);
or U15393 (N_15393,N_14534,N_14240);
xor U15394 (N_15394,N_14523,N_14229);
nand U15395 (N_15395,N_14735,N_14458);
or U15396 (N_15396,N_14540,N_14284);
and U15397 (N_15397,N_14712,N_14278);
nand U15398 (N_15398,N_14650,N_14975);
nand U15399 (N_15399,N_14338,N_14608);
nand U15400 (N_15400,N_14821,N_14728);
and U15401 (N_15401,N_14560,N_14652);
and U15402 (N_15402,N_14377,N_14710);
nand U15403 (N_15403,N_14666,N_14616);
nand U15404 (N_15404,N_14285,N_14179);
and U15405 (N_15405,N_14557,N_14937);
xor U15406 (N_15406,N_14554,N_14546);
nand U15407 (N_15407,N_14408,N_14204);
xnor U15408 (N_15408,N_14461,N_14456);
and U15409 (N_15409,N_14004,N_14516);
xor U15410 (N_15410,N_14010,N_14792);
and U15411 (N_15411,N_14698,N_14732);
xor U15412 (N_15412,N_14181,N_14727);
xnor U15413 (N_15413,N_14943,N_14404);
nand U15414 (N_15414,N_14282,N_14188);
and U15415 (N_15415,N_14441,N_14944);
nand U15416 (N_15416,N_14105,N_14134);
nand U15417 (N_15417,N_14871,N_14091);
or U15418 (N_15418,N_14815,N_14037);
or U15419 (N_15419,N_14328,N_14525);
and U15420 (N_15420,N_14132,N_14395);
and U15421 (N_15421,N_14705,N_14088);
or U15422 (N_15422,N_14567,N_14682);
and U15423 (N_15423,N_14354,N_14801);
or U15424 (N_15424,N_14259,N_14870);
nand U15425 (N_15425,N_14112,N_14345);
and U15426 (N_15426,N_14976,N_14466);
and U15427 (N_15427,N_14991,N_14892);
nand U15428 (N_15428,N_14155,N_14436);
nor U15429 (N_15429,N_14872,N_14165);
nor U15430 (N_15430,N_14607,N_14764);
or U15431 (N_15431,N_14104,N_14173);
nor U15432 (N_15432,N_14591,N_14351);
xnor U15433 (N_15433,N_14515,N_14230);
or U15434 (N_15434,N_14265,N_14935);
nor U15435 (N_15435,N_14393,N_14702);
and U15436 (N_15436,N_14645,N_14289);
or U15437 (N_15437,N_14115,N_14024);
or U15438 (N_15438,N_14275,N_14159);
nor U15439 (N_15439,N_14271,N_14749);
nor U15440 (N_15440,N_14087,N_14574);
and U15441 (N_15441,N_14638,N_14573);
nor U15442 (N_15442,N_14614,N_14707);
nor U15443 (N_15443,N_14960,N_14146);
and U15444 (N_15444,N_14855,N_14826);
or U15445 (N_15445,N_14363,N_14864);
xnor U15446 (N_15446,N_14981,N_14565);
or U15447 (N_15447,N_14187,N_14808);
nor U15448 (N_15448,N_14066,N_14113);
nand U15449 (N_15449,N_14051,N_14417);
or U15450 (N_15450,N_14167,N_14210);
nor U15451 (N_15451,N_14200,N_14260);
nor U15452 (N_15452,N_14221,N_14867);
and U15453 (N_15453,N_14836,N_14681);
and U15454 (N_15454,N_14152,N_14244);
nor U15455 (N_15455,N_14126,N_14378);
xnor U15456 (N_15456,N_14936,N_14623);
xor U15457 (N_15457,N_14620,N_14642);
xor U15458 (N_15458,N_14364,N_14950);
or U15459 (N_15459,N_14143,N_14225);
nand U15460 (N_15460,N_14357,N_14803);
xor U15461 (N_15461,N_14890,N_14881);
nand U15462 (N_15462,N_14737,N_14884);
or U15463 (N_15463,N_14321,N_14633);
nand U15464 (N_15464,N_14170,N_14983);
or U15465 (N_15465,N_14147,N_14838);
and U15466 (N_15466,N_14425,N_14536);
and U15467 (N_15467,N_14673,N_14873);
or U15468 (N_15468,N_14038,N_14202);
nand U15469 (N_15469,N_14307,N_14671);
xnor U15470 (N_15470,N_14373,N_14718);
nand U15471 (N_15471,N_14750,N_14690);
and U15472 (N_15472,N_14297,N_14414);
or U15473 (N_15473,N_14911,N_14820);
or U15474 (N_15474,N_14163,N_14029);
nor U15475 (N_15475,N_14763,N_14993);
or U15476 (N_15476,N_14972,N_14401);
nand U15477 (N_15477,N_14106,N_14020);
nor U15478 (N_15478,N_14920,N_14918);
nand U15479 (N_15479,N_14511,N_14470);
nor U15480 (N_15480,N_14659,N_14743);
xor U15481 (N_15481,N_14341,N_14830);
nand U15482 (N_15482,N_14916,N_14498);
and U15483 (N_15483,N_14236,N_14298);
nand U15484 (N_15484,N_14372,N_14887);
xor U15485 (N_15485,N_14055,N_14007);
and U15486 (N_15486,N_14205,N_14102);
and U15487 (N_15487,N_14898,N_14454);
and U15488 (N_15488,N_14171,N_14776);
nand U15489 (N_15489,N_14601,N_14499);
nor U15490 (N_15490,N_14783,N_14145);
or U15491 (N_15491,N_14054,N_14790);
xor U15492 (N_15492,N_14291,N_14824);
nor U15493 (N_15493,N_14552,N_14306);
nand U15494 (N_15494,N_14639,N_14148);
nand U15495 (N_15495,N_14374,N_14311);
nor U15496 (N_15496,N_14576,N_14199);
nor U15497 (N_15497,N_14209,N_14412);
xnor U15498 (N_15498,N_14190,N_14883);
or U15499 (N_15499,N_14349,N_14891);
xnor U15500 (N_15500,N_14230,N_14395);
nor U15501 (N_15501,N_14687,N_14328);
nand U15502 (N_15502,N_14894,N_14233);
or U15503 (N_15503,N_14911,N_14955);
nand U15504 (N_15504,N_14476,N_14497);
xor U15505 (N_15505,N_14535,N_14031);
nor U15506 (N_15506,N_14880,N_14752);
and U15507 (N_15507,N_14724,N_14337);
nor U15508 (N_15508,N_14517,N_14372);
and U15509 (N_15509,N_14020,N_14372);
nor U15510 (N_15510,N_14007,N_14053);
or U15511 (N_15511,N_14634,N_14294);
and U15512 (N_15512,N_14825,N_14195);
or U15513 (N_15513,N_14483,N_14172);
and U15514 (N_15514,N_14243,N_14807);
nand U15515 (N_15515,N_14452,N_14111);
or U15516 (N_15516,N_14119,N_14932);
and U15517 (N_15517,N_14224,N_14702);
and U15518 (N_15518,N_14089,N_14386);
and U15519 (N_15519,N_14568,N_14411);
nand U15520 (N_15520,N_14583,N_14156);
nor U15521 (N_15521,N_14538,N_14949);
nor U15522 (N_15522,N_14578,N_14547);
nand U15523 (N_15523,N_14082,N_14455);
or U15524 (N_15524,N_14490,N_14198);
nand U15525 (N_15525,N_14230,N_14888);
or U15526 (N_15526,N_14236,N_14261);
nand U15527 (N_15527,N_14607,N_14985);
nand U15528 (N_15528,N_14396,N_14047);
xnor U15529 (N_15529,N_14775,N_14033);
nor U15530 (N_15530,N_14848,N_14132);
nand U15531 (N_15531,N_14250,N_14297);
nor U15532 (N_15532,N_14824,N_14512);
and U15533 (N_15533,N_14944,N_14553);
and U15534 (N_15534,N_14387,N_14519);
nor U15535 (N_15535,N_14468,N_14532);
nor U15536 (N_15536,N_14879,N_14997);
xnor U15537 (N_15537,N_14831,N_14842);
nand U15538 (N_15538,N_14025,N_14851);
nor U15539 (N_15539,N_14116,N_14451);
nor U15540 (N_15540,N_14704,N_14852);
or U15541 (N_15541,N_14577,N_14967);
nor U15542 (N_15542,N_14926,N_14697);
and U15543 (N_15543,N_14205,N_14332);
nor U15544 (N_15544,N_14316,N_14002);
and U15545 (N_15545,N_14783,N_14988);
xor U15546 (N_15546,N_14268,N_14758);
nand U15547 (N_15547,N_14929,N_14378);
or U15548 (N_15548,N_14950,N_14136);
and U15549 (N_15549,N_14656,N_14795);
xor U15550 (N_15550,N_14484,N_14910);
or U15551 (N_15551,N_14704,N_14302);
nor U15552 (N_15552,N_14781,N_14396);
xor U15553 (N_15553,N_14660,N_14404);
nor U15554 (N_15554,N_14790,N_14056);
xor U15555 (N_15555,N_14628,N_14182);
nor U15556 (N_15556,N_14910,N_14309);
nand U15557 (N_15557,N_14563,N_14627);
nor U15558 (N_15558,N_14343,N_14766);
or U15559 (N_15559,N_14348,N_14716);
or U15560 (N_15560,N_14425,N_14338);
nand U15561 (N_15561,N_14489,N_14052);
nand U15562 (N_15562,N_14426,N_14455);
nor U15563 (N_15563,N_14815,N_14899);
or U15564 (N_15564,N_14478,N_14639);
and U15565 (N_15565,N_14306,N_14028);
or U15566 (N_15566,N_14478,N_14603);
nor U15567 (N_15567,N_14934,N_14654);
and U15568 (N_15568,N_14690,N_14870);
xnor U15569 (N_15569,N_14693,N_14662);
nor U15570 (N_15570,N_14234,N_14053);
nand U15571 (N_15571,N_14680,N_14209);
xnor U15572 (N_15572,N_14954,N_14754);
nand U15573 (N_15573,N_14179,N_14712);
or U15574 (N_15574,N_14000,N_14082);
nor U15575 (N_15575,N_14154,N_14455);
and U15576 (N_15576,N_14730,N_14033);
or U15577 (N_15577,N_14440,N_14500);
xor U15578 (N_15578,N_14612,N_14835);
nand U15579 (N_15579,N_14744,N_14660);
nand U15580 (N_15580,N_14889,N_14680);
nor U15581 (N_15581,N_14106,N_14808);
xor U15582 (N_15582,N_14615,N_14229);
and U15583 (N_15583,N_14116,N_14931);
nor U15584 (N_15584,N_14340,N_14549);
and U15585 (N_15585,N_14939,N_14502);
nor U15586 (N_15586,N_14720,N_14856);
nor U15587 (N_15587,N_14891,N_14811);
or U15588 (N_15588,N_14735,N_14809);
and U15589 (N_15589,N_14920,N_14687);
xor U15590 (N_15590,N_14872,N_14169);
nand U15591 (N_15591,N_14650,N_14987);
xor U15592 (N_15592,N_14910,N_14011);
and U15593 (N_15593,N_14656,N_14378);
and U15594 (N_15594,N_14160,N_14754);
and U15595 (N_15595,N_14854,N_14930);
nor U15596 (N_15596,N_14476,N_14985);
or U15597 (N_15597,N_14027,N_14675);
xnor U15598 (N_15598,N_14258,N_14582);
nand U15599 (N_15599,N_14313,N_14140);
and U15600 (N_15600,N_14355,N_14762);
nor U15601 (N_15601,N_14686,N_14189);
or U15602 (N_15602,N_14858,N_14338);
nand U15603 (N_15603,N_14039,N_14811);
or U15604 (N_15604,N_14168,N_14374);
nand U15605 (N_15605,N_14386,N_14056);
or U15606 (N_15606,N_14269,N_14195);
nor U15607 (N_15607,N_14765,N_14580);
nand U15608 (N_15608,N_14963,N_14416);
and U15609 (N_15609,N_14438,N_14282);
or U15610 (N_15610,N_14503,N_14900);
nand U15611 (N_15611,N_14884,N_14524);
xor U15612 (N_15612,N_14200,N_14118);
and U15613 (N_15613,N_14715,N_14501);
or U15614 (N_15614,N_14771,N_14858);
xnor U15615 (N_15615,N_14751,N_14886);
and U15616 (N_15616,N_14831,N_14138);
xnor U15617 (N_15617,N_14168,N_14490);
nor U15618 (N_15618,N_14066,N_14313);
and U15619 (N_15619,N_14759,N_14937);
and U15620 (N_15620,N_14331,N_14083);
nand U15621 (N_15621,N_14595,N_14917);
or U15622 (N_15622,N_14689,N_14300);
nand U15623 (N_15623,N_14077,N_14398);
xnor U15624 (N_15624,N_14471,N_14428);
nand U15625 (N_15625,N_14913,N_14783);
and U15626 (N_15626,N_14773,N_14932);
and U15627 (N_15627,N_14987,N_14566);
nor U15628 (N_15628,N_14088,N_14091);
and U15629 (N_15629,N_14262,N_14366);
xor U15630 (N_15630,N_14042,N_14281);
nand U15631 (N_15631,N_14314,N_14961);
or U15632 (N_15632,N_14011,N_14966);
xnor U15633 (N_15633,N_14389,N_14687);
and U15634 (N_15634,N_14955,N_14346);
and U15635 (N_15635,N_14811,N_14967);
and U15636 (N_15636,N_14056,N_14091);
or U15637 (N_15637,N_14306,N_14894);
and U15638 (N_15638,N_14371,N_14240);
xnor U15639 (N_15639,N_14260,N_14513);
xnor U15640 (N_15640,N_14704,N_14713);
xor U15641 (N_15641,N_14949,N_14443);
nor U15642 (N_15642,N_14918,N_14052);
or U15643 (N_15643,N_14096,N_14726);
nor U15644 (N_15644,N_14932,N_14351);
nand U15645 (N_15645,N_14621,N_14937);
or U15646 (N_15646,N_14068,N_14367);
nand U15647 (N_15647,N_14997,N_14523);
or U15648 (N_15648,N_14116,N_14340);
and U15649 (N_15649,N_14352,N_14326);
or U15650 (N_15650,N_14949,N_14357);
nor U15651 (N_15651,N_14698,N_14643);
xor U15652 (N_15652,N_14189,N_14393);
or U15653 (N_15653,N_14638,N_14188);
xnor U15654 (N_15654,N_14346,N_14229);
xor U15655 (N_15655,N_14600,N_14629);
xor U15656 (N_15656,N_14479,N_14164);
xnor U15657 (N_15657,N_14948,N_14243);
and U15658 (N_15658,N_14126,N_14588);
nand U15659 (N_15659,N_14711,N_14073);
nand U15660 (N_15660,N_14483,N_14773);
xor U15661 (N_15661,N_14436,N_14989);
nand U15662 (N_15662,N_14962,N_14337);
nand U15663 (N_15663,N_14393,N_14711);
or U15664 (N_15664,N_14731,N_14598);
nand U15665 (N_15665,N_14848,N_14074);
xnor U15666 (N_15666,N_14643,N_14309);
and U15667 (N_15667,N_14668,N_14554);
nor U15668 (N_15668,N_14283,N_14591);
nand U15669 (N_15669,N_14275,N_14093);
nor U15670 (N_15670,N_14115,N_14815);
nand U15671 (N_15671,N_14958,N_14898);
or U15672 (N_15672,N_14598,N_14195);
xor U15673 (N_15673,N_14578,N_14639);
and U15674 (N_15674,N_14105,N_14743);
and U15675 (N_15675,N_14290,N_14176);
nand U15676 (N_15676,N_14585,N_14947);
nor U15677 (N_15677,N_14872,N_14595);
nand U15678 (N_15678,N_14312,N_14989);
xor U15679 (N_15679,N_14640,N_14829);
or U15680 (N_15680,N_14575,N_14602);
xnor U15681 (N_15681,N_14495,N_14562);
or U15682 (N_15682,N_14979,N_14218);
nand U15683 (N_15683,N_14779,N_14688);
nor U15684 (N_15684,N_14903,N_14321);
and U15685 (N_15685,N_14358,N_14127);
nor U15686 (N_15686,N_14267,N_14125);
nand U15687 (N_15687,N_14256,N_14574);
nor U15688 (N_15688,N_14339,N_14317);
nor U15689 (N_15689,N_14836,N_14796);
nor U15690 (N_15690,N_14502,N_14707);
xnor U15691 (N_15691,N_14767,N_14102);
and U15692 (N_15692,N_14112,N_14963);
and U15693 (N_15693,N_14644,N_14971);
nor U15694 (N_15694,N_14992,N_14048);
xor U15695 (N_15695,N_14334,N_14774);
or U15696 (N_15696,N_14086,N_14718);
and U15697 (N_15697,N_14080,N_14276);
nor U15698 (N_15698,N_14215,N_14464);
or U15699 (N_15699,N_14965,N_14663);
xor U15700 (N_15700,N_14743,N_14563);
nand U15701 (N_15701,N_14005,N_14127);
or U15702 (N_15702,N_14040,N_14617);
nand U15703 (N_15703,N_14814,N_14498);
and U15704 (N_15704,N_14031,N_14908);
nand U15705 (N_15705,N_14309,N_14740);
xnor U15706 (N_15706,N_14682,N_14673);
nor U15707 (N_15707,N_14037,N_14267);
and U15708 (N_15708,N_14568,N_14020);
nand U15709 (N_15709,N_14408,N_14683);
xor U15710 (N_15710,N_14845,N_14555);
nand U15711 (N_15711,N_14011,N_14129);
and U15712 (N_15712,N_14649,N_14134);
xor U15713 (N_15713,N_14879,N_14050);
or U15714 (N_15714,N_14286,N_14202);
or U15715 (N_15715,N_14546,N_14075);
and U15716 (N_15716,N_14812,N_14796);
and U15717 (N_15717,N_14767,N_14862);
xor U15718 (N_15718,N_14527,N_14998);
nor U15719 (N_15719,N_14726,N_14951);
xor U15720 (N_15720,N_14372,N_14485);
or U15721 (N_15721,N_14718,N_14531);
nor U15722 (N_15722,N_14312,N_14838);
or U15723 (N_15723,N_14291,N_14982);
nor U15724 (N_15724,N_14401,N_14789);
or U15725 (N_15725,N_14040,N_14922);
or U15726 (N_15726,N_14273,N_14104);
or U15727 (N_15727,N_14304,N_14308);
and U15728 (N_15728,N_14396,N_14049);
nand U15729 (N_15729,N_14224,N_14498);
nand U15730 (N_15730,N_14513,N_14271);
or U15731 (N_15731,N_14965,N_14507);
xnor U15732 (N_15732,N_14787,N_14404);
xor U15733 (N_15733,N_14686,N_14279);
and U15734 (N_15734,N_14825,N_14655);
nor U15735 (N_15735,N_14535,N_14252);
xor U15736 (N_15736,N_14467,N_14720);
nor U15737 (N_15737,N_14308,N_14622);
and U15738 (N_15738,N_14708,N_14294);
nor U15739 (N_15739,N_14560,N_14976);
nor U15740 (N_15740,N_14206,N_14089);
xor U15741 (N_15741,N_14288,N_14043);
xor U15742 (N_15742,N_14266,N_14909);
nand U15743 (N_15743,N_14737,N_14692);
xnor U15744 (N_15744,N_14647,N_14145);
nand U15745 (N_15745,N_14050,N_14650);
or U15746 (N_15746,N_14519,N_14621);
nor U15747 (N_15747,N_14013,N_14282);
nand U15748 (N_15748,N_14369,N_14110);
xor U15749 (N_15749,N_14747,N_14854);
nand U15750 (N_15750,N_14548,N_14852);
and U15751 (N_15751,N_14528,N_14140);
or U15752 (N_15752,N_14549,N_14222);
xnor U15753 (N_15753,N_14737,N_14300);
nor U15754 (N_15754,N_14666,N_14415);
and U15755 (N_15755,N_14494,N_14683);
nor U15756 (N_15756,N_14935,N_14141);
and U15757 (N_15757,N_14048,N_14137);
nor U15758 (N_15758,N_14336,N_14584);
nor U15759 (N_15759,N_14831,N_14122);
nor U15760 (N_15760,N_14646,N_14312);
nand U15761 (N_15761,N_14325,N_14467);
or U15762 (N_15762,N_14614,N_14836);
nand U15763 (N_15763,N_14151,N_14366);
nand U15764 (N_15764,N_14705,N_14855);
or U15765 (N_15765,N_14727,N_14702);
nand U15766 (N_15766,N_14017,N_14045);
nand U15767 (N_15767,N_14568,N_14620);
or U15768 (N_15768,N_14576,N_14773);
xor U15769 (N_15769,N_14671,N_14635);
xor U15770 (N_15770,N_14803,N_14438);
nor U15771 (N_15771,N_14376,N_14649);
nand U15772 (N_15772,N_14398,N_14703);
and U15773 (N_15773,N_14810,N_14212);
nor U15774 (N_15774,N_14392,N_14407);
xor U15775 (N_15775,N_14881,N_14760);
and U15776 (N_15776,N_14952,N_14845);
xnor U15777 (N_15777,N_14811,N_14215);
xor U15778 (N_15778,N_14276,N_14841);
or U15779 (N_15779,N_14169,N_14972);
nor U15780 (N_15780,N_14676,N_14886);
nor U15781 (N_15781,N_14905,N_14455);
nor U15782 (N_15782,N_14339,N_14862);
or U15783 (N_15783,N_14668,N_14394);
nor U15784 (N_15784,N_14653,N_14863);
or U15785 (N_15785,N_14383,N_14165);
nand U15786 (N_15786,N_14277,N_14390);
or U15787 (N_15787,N_14681,N_14029);
and U15788 (N_15788,N_14355,N_14325);
xnor U15789 (N_15789,N_14262,N_14855);
and U15790 (N_15790,N_14753,N_14081);
or U15791 (N_15791,N_14344,N_14314);
or U15792 (N_15792,N_14511,N_14810);
nand U15793 (N_15793,N_14307,N_14096);
or U15794 (N_15794,N_14390,N_14434);
nand U15795 (N_15795,N_14035,N_14326);
nor U15796 (N_15796,N_14267,N_14488);
and U15797 (N_15797,N_14052,N_14281);
xnor U15798 (N_15798,N_14367,N_14750);
nand U15799 (N_15799,N_14222,N_14873);
or U15800 (N_15800,N_14768,N_14440);
nor U15801 (N_15801,N_14056,N_14896);
xnor U15802 (N_15802,N_14704,N_14446);
nor U15803 (N_15803,N_14109,N_14740);
or U15804 (N_15804,N_14538,N_14888);
nor U15805 (N_15805,N_14443,N_14749);
nand U15806 (N_15806,N_14792,N_14105);
and U15807 (N_15807,N_14386,N_14545);
and U15808 (N_15808,N_14208,N_14057);
or U15809 (N_15809,N_14366,N_14097);
xnor U15810 (N_15810,N_14624,N_14558);
or U15811 (N_15811,N_14273,N_14372);
nor U15812 (N_15812,N_14633,N_14825);
nor U15813 (N_15813,N_14696,N_14184);
and U15814 (N_15814,N_14349,N_14775);
and U15815 (N_15815,N_14758,N_14339);
nor U15816 (N_15816,N_14669,N_14223);
and U15817 (N_15817,N_14281,N_14057);
or U15818 (N_15818,N_14320,N_14672);
and U15819 (N_15819,N_14794,N_14004);
xor U15820 (N_15820,N_14381,N_14095);
nor U15821 (N_15821,N_14908,N_14429);
or U15822 (N_15822,N_14176,N_14900);
and U15823 (N_15823,N_14564,N_14975);
or U15824 (N_15824,N_14248,N_14516);
xor U15825 (N_15825,N_14492,N_14621);
nor U15826 (N_15826,N_14932,N_14568);
or U15827 (N_15827,N_14465,N_14576);
nand U15828 (N_15828,N_14018,N_14357);
nor U15829 (N_15829,N_14883,N_14203);
or U15830 (N_15830,N_14638,N_14689);
or U15831 (N_15831,N_14562,N_14954);
xor U15832 (N_15832,N_14723,N_14294);
and U15833 (N_15833,N_14737,N_14665);
xor U15834 (N_15834,N_14579,N_14125);
xnor U15835 (N_15835,N_14803,N_14129);
and U15836 (N_15836,N_14256,N_14109);
and U15837 (N_15837,N_14298,N_14505);
and U15838 (N_15838,N_14238,N_14587);
xnor U15839 (N_15839,N_14592,N_14094);
and U15840 (N_15840,N_14243,N_14019);
or U15841 (N_15841,N_14821,N_14149);
nor U15842 (N_15842,N_14086,N_14655);
or U15843 (N_15843,N_14433,N_14374);
xnor U15844 (N_15844,N_14130,N_14763);
nor U15845 (N_15845,N_14640,N_14369);
xor U15846 (N_15846,N_14846,N_14013);
nor U15847 (N_15847,N_14852,N_14089);
nor U15848 (N_15848,N_14881,N_14413);
and U15849 (N_15849,N_14881,N_14492);
nor U15850 (N_15850,N_14356,N_14865);
or U15851 (N_15851,N_14347,N_14091);
or U15852 (N_15852,N_14392,N_14487);
nand U15853 (N_15853,N_14954,N_14344);
xor U15854 (N_15854,N_14109,N_14671);
nand U15855 (N_15855,N_14035,N_14367);
and U15856 (N_15856,N_14831,N_14992);
or U15857 (N_15857,N_14381,N_14066);
or U15858 (N_15858,N_14262,N_14518);
xnor U15859 (N_15859,N_14839,N_14939);
and U15860 (N_15860,N_14567,N_14043);
nand U15861 (N_15861,N_14003,N_14805);
or U15862 (N_15862,N_14819,N_14538);
xor U15863 (N_15863,N_14549,N_14105);
nor U15864 (N_15864,N_14468,N_14842);
nor U15865 (N_15865,N_14936,N_14514);
nor U15866 (N_15866,N_14541,N_14696);
nand U15867 (N_15867,N_14047,N_14357);
or U15868 (N_15868,N_14292,N_14482);
xnor U15869 (N_15869,N_14424,N_14389);
and U15870 (N_15870,N_14404,N_14532);
or U15871 (N_15871,N_14711,N_14959);
or U15872 (N_15872,N_14256,N_14105);
nor U15873 (N_15873,N_14217,N_14188);
xor U15874 (N_15874,N_14911,N_14692);
nand U15875 (N_15875,N_14116,N_14318);
or U15876 (N_15876,N_14218,N_14503);
nand U15877 (N_15877,N_14130,N_14116);
and U15878 (N_15878,N_14802,N_14633);
xnor U15879 (N_15879,N_14379,N_14304);
xor U15880 (N_15880,N_14144,N_14938);
xnor U15881 (N_15881,N_14440,N_14711);
nor U15882 (N_15882,N_14634,N_14979);
nor U15883 (N_15883,N_14465,N_14392);
xor U15884 (N_15884,N_14928,N_14549);
nand U15885 (N_15885,N_14899,N_14118);
and U15886 (N_15886,N_14007,N_14213);
nor U15887 (N_15887,N_14517,N_14562);
nor U15888 (N_15888,N_14717,N_14369);
nand U15889 (N_15889,N_14790,N_14012);
nor U15890 (N_15890,N_14148,N_14407);
nand U15891 (N_15891,N_14751,N_14764);
and U15892 (N_15892,N_14128,N_14457);
nor U15893 (N_15893,N_14789,N_14760);
or U15894 (N_15894,N_14469,N_14380);
or U15895 (N_15895,N_14293,N_14083);
and U15896 (N_15896,N_14471,N_14613);
nor U15897 (N_15897,N_14976,N_14500);
and U15898 (N_15898,N_14133,N_14809);
or U15899 (N_15899,N_14457,N_14149);
nor U15900 (N_15900,N_14508,N_14216);
xor U15901 (N_15901,N_14035,N_14495);
xor U15902 (N_15902,N_14854,N_14677);
nor U15903 (N_15903,N_14746,N_14611);
xnor U15904 (N_15904,N_14676,N_14070);
nor U15905 (N_15905,N_14182,N_14392);
or U15906 (N_15906,N_14903,N_14173);
nand U15907 (N_15907,N_14281,N_14904);
nor U15908 (N_15908,N_14441,N_14009);
nor U15909 (N_15909,N_14652,N_14897);
xor U15910 (N_15910,N_14757,N_14376);
nor U15911 (N_15911,N_14650,N_14848);
xnor U15912 (N_15912,N_14135,N_14868);
xnor U15913 (N_15913,N_14936,N_14921);
or U15914 (N_15914,N_14663,N_14816);
nand U15915 (N_15915,N_14239,N_14417);
nor U15916 (N_15916,N_14186,N_14621);
xnor U15917 (N_15917,N_14802,N_14893);
nand U15918 (N_15918,N_14142,N_14348);
nor U15919 (N_15919,N_14728,N_14826);
xor U15920 (N_15920,N_14242,N_14410);
or U15921 (N_15921,N_14115,N_14776);
nor U15922 (N_15922,N_14880,N_14335);
and U15923 (N_15923,N_14182,N_14184);
nand U15924 (N_15924,N_14243,N_14457);
nor U15925 (N_15925,N_14721,N_14416);
nor U15926 (N_15926,N_14763,N_14132);
xnor U15927 (N_15927,N_14631,N_14755);
nor U15928 (N_15928,N_14622,N_14625);
and U15929 (N_15929,N_14724,N_14074);
and U15930 (N_15930,N_14267,N_14190);
or U15931 (N_15931,N_14957,N_14821);
nand U15932 (N_15932,N_14658,N_14596);
nor U15933 (N_15933,N_14730,N_14409);
and U15934 (N_15934,N_14968,N_14301);
nor U15935 (N_15935,N_14897,N_14684);
and U15936 (N_15936,N_14673,N_14854);
and U15937 (N_15937,N_14237,N_14783);
and U15938 (N_15938,N_14260,N_14719);
xor U15939 (N_15939,N_14020,N_14006);
xor U15940 (N_15940,N_14605,N_14119);
nand U15941 (N_15941,N_14073,N_14531);
or U15942 (N_15942,N_14706,N_14026);
or U15943 (N_15943,N_14374,N_14664);
and U15944 (N_15944,N_14287,N_14609);
or U15945 (N_15945,N_14436,N_14008);
nor U15946 (N_15946,N_14998,N_14902);
nand U15947 (N_15947,N_14422,N_14997);
nand U15948 (N_15948,N_14085,N_14489);
nor U15949 (N_15949,N_14832,N_14413);
or U15950 (N_15950,N_14299,N_14947);
and U15951 (N_15951,N_14911,N_14943);
or U15952 (N_15952,N_14778,N_14214);
and U15953 (N_15953,N_14942,N_14525);
xnor U15954 (N_15954,N_14050,N_14845);
or U15955 (N_15955,N_14354,N_14503);
or U15956 (N_15956,N_14312,N_14716);
and U15957 (N_15957,N_14346,N_14170);
xnor U15958 (N_15958,N_14079,N_14833);
nand U15959 (N_15959,N_14210,N_14924);
xor U15960 (N_15960,N_14674,N_14178);
nand U15961 (N_15961,N_14479,N_14772);
or U15962 (N_15962,N_14547,N_14412);
nand U15963 (N_15963,N_14044,N_14509);
nand U15964 (N_15964,N_14290,N_14383);
or U15965 (N_15965,N_14294,N_14794);
or U15966 (N_15966,N_14858,N_14051);
xor U15967 (N_15967,N_14897,N_14958);
xor U15968 (N_15968,N_14372,N_14378);
or U15969 (N_15969,N_14759,N_14588);
nor U15970 (N_15970,N_14228,N_14394);
nand U15971 (N_15971,N_14119,N_14565);
xnor U15972 (N_15972,N_14622,N_14083);
nor U15973 (N_15973,N_14438,N_14357);
nand U15974 (N_15974,N_14643,N_14682);
and U15975 (N_15975,N_14402,N_14427);
nor U15976 (N_15976,N_14993,N_14475);
xor U15977 (N_15977,N_14800,N_14794);
and U15978 (N_15978,N_14950,N_14973);
and U15979 (N_15979,N_14716,N_14466);
and U15980 (N_15980,N_14949,N_14002);
nor U15981 (N_15981,N_14760,N_14182);
and U15982 (N_15982,N_14111,N_14019);
nand U15983 (N_15983,N_14879,N_14970);
nand U15984 (N_15984,N_14230,N_14373);
nand U15985 (N_15985,N_14768,N_14707);
or U15986 (N_15986,N_14291,N_14340);
or U15987 (N_15987,N_14543,N_14485);
nor U15988 (N_15988,N_14227,N_14250);
nand U15989 (N_15989,N_14786,N_14423);
nand U15990 (N_15990,N_14197,N_14236);
or U15991 (N_15991,N_14322,N_14363);
or U15992 (N_15992,N_14187,N_14905);
nor U15993 (N_15993,N_14502,N_14014);
and U15994 (N_15994,N_14454,N_14863);
nand U15995 (N_15995,N_14416,N_14376);
or U15996 (N_15996,N_14190,N_14938);
and U15997 (N_15997,N_14930,N_14195);
or U15998 (N_15998,N_14626,N_14605);
xnor U15999 (N_15999,N_14952,N_14439);
nand U16000 (N_16000,N_15494,N_15561);
and U16001 (N_16001,N_15839,N_15944);
nand U16002 (N_16002,N_15925,N_15688);
nor U16003 (N_16003,N_15308,N_15512);
xnor U16004 (N_16004,N_15201,N_15411);
xor U16005 (N_16005,N_15467,N_15229);
and U16006 (N_16006,N_15193,N_15078);
nand U16007 (N_16007,N_15773,N_15216);
or U16008 (N_16008,N_15838,N_15662);
xor U16009 (N_16009,N_15126,N_15824);
nand U16010 (N_16010,N_15014,N_15405);
nand U16011 (N_16011,N_15421,N_15691);
xor U16012 (N_16012,N_15429,N_15288);
xnor U16013 (N_16013,N_15204,N_15530);
or U16014 (N_16014,N_15721,N_15181);
xor U16015 (N_16015,N_15031,N_15079);
xnor U16016 (N_16016,N_15881,N_15585);
nand U16017 (N_16017,N_15789,N_15784);
xnor U16018 (N_16018,N_15750,N_15792);
nand U16019 (N_16019,N_15987,N_15812);
xor U16020 (N_16020,N_15111,N_15149);
nor U16021 (N_16021,N_15300,N_15960);
xor U16022 (N_16022,N_15811,N_15047);
and U16023 (N_16023,N_15053,N_15403);
and U16024 (N_16024,N_15420,N_15055);
and U16025 (N_16025,N_15356,N_15077);
nand U16026 (N_16026,N_15438,N_15781);
or U16027 (N_16027,N_15909,N_15440);
and U16028 (N_16028,N_15353,N_15970);
xnor U16029 (N_16029,N_15952,N_15097);
nor U16030 (N_16030,N_15820,N_15633);
nand U16031 (N_16031,N_15926,N_15546);
nand U16032 (N_16032,N_15565,N_15091);
and U16033 (N_16033,N_15590,N_15763);
nand U16034 (N_16034,N_15066,N_15674);
or U16035 (N_16035,N_15117,N_15445);
nand U16036 (N_16036,N_15890,N_15070);
and U16037 (N_16037,N_15409,N_15772);
xor U16038 (N_16038,N_15019,N_15101);
nor U16039 (N_16039,N_15904,N_15888);
nor U16040 (N_16040,N_15399,N_15114);
xnor U16041 (N_16041,N_15335,N_15284);
or U16042 (N_16042,N_15912,N_15094);
and U16043 (N_16043,N_15550,N_15397);
nand U16044 (N_16044,N_15365,N_15331);
or U16045 (N_16045,N_15879,N_15206);
or U16046 (N_16046,N_15898,N_15707);
or U16047 (N_16047,N_15068,N_15525);
nor U16048 (N_16048,N_15398,N_15861);
nand U16049 (N_16049,N_15661,N_15786);
and U16050 (N_16050,N_15184,N_15516);
or U16051 (N_16051,N_15532,N_15825);
nand U16052 (N_16052,N_15843,N_15415);
nor U16053 (N_16053,N_15998,N_15367);
xnor U16054 (N_16054,N_15639,N_15473);
nor U16055 (N_16055,N_15606,N_15815);
xnor U16056 (N_16056,N_15627,N_15041);
nor U16057 (N_16057,N_15870,N_15695);
xor U16058 (N_16058,N_15032,N_15779);
nand U16059 (N_16059,N_15947,N_15533);
nor U16060 (N_16060,N_15521,N_15185);
nand U16061 (N_16061,N_15859,N_15673);
nor U16062 (N_16062,N_15587,N_15207);
nor U16063 (N_16063,N_15451,N_15683);
nor U16064 (N_16064,N_15882,N_15938);
and U16065 (N_16065,N_15120,N_15314);
xnor U16066 (N_16066,N_15218,N_15122);
nand U16067 (N_16067,N_15033,N_15214);
nand U16068 (N_16068,N_15575,N_15406);
xor U16069 (N_16069,N_15108,N_15900);
or U16070 (N_16070,N_15359,N_15745);
nand U16071 (N_16071,N_15280,N_15934);
and U16072 (N_16072,N_15630,N_15906);
or U16073 (N_16073,N_15624,N_15013);
and U16074 (N_16074,N_15901,N_15913);
xor U16075 (N_16075,N_15497,N_15829);
nor U16076 (N_16076,N_15488,N_15480);
or U16077 (N_16077,N_15831,N_15294);
xor U16078 (N_16078,N_15188,N_15338);
or U16079 (N_16079,N_15584,N_15486);
or U16080 (N_16080,N_15596,N_15030);
nand U16081 (N_16081,N_15025,N_15166);
or U16082 (N_16082,N_15663,N_15493);
or U16083 (N_16083,N_15866,N_15005);
xnor U16084 (N_16084,N_15891,N_15576);
or U16085 (N_16085,N_15876,N_15400);
xor U16086 (N_16086,N_15387,N_15813);
nand U16087 (N_16087,N_15412,N_15837);
xnor U16088 (N_16088,N_15278,N_15263);
nor U16089 (N_16089,N_15062,N_15833);
and U16090 (N_16090,N_15298,N_15247);
or U16091 (N_16091,N_15463,N_15703);
xor U16092 (N_16092,N_15964,N_15995);
or U16093 (N_16093,N_15694,N_15592);
nor U16094 (N_16094,N_15687,N_15959);
and U16095 (N_16095,N_15170,N_15864);
and U16096 (N_16096,N_15322,N_15408);
nand U16097 (N_16097,N_15747,N_15296);
nor U16098 (N_16098,N_15855,N_15669);
nand U16099 (N_16099,N_15395,N_15049);
nor U16100 (N_16100,N_15375,N_15656);
and U16101 (N_16101,N_15577,N_15963);
nand U16102 (N_16102,N_15857,N_15116);
nand U16103 (N_16103,N_15133,N_15783);
nor U16104 (N_16104,N_15301,N_15740);
xor U16105 (N_16105,N_15716,N_15161);
xnor U16106 (N_16106,N_15137,N_15460);
and U16107 (N_16107,N_15197,N_15290);
xnor U16108 (N_16108,N_15540,N_15629);
and U16109 (N_16109,N_15657,N_15644);
nand U16110 (N_16110,N_15720,N_15761);
nand U16111 (N_16111,N_15416,N_15991);
nor U16112 (N_16112,N_15524,N_15706);
or U16113 (N_16113,N_15834,N_15520);
and U16114 (N_16114,N_15896,N_15977);
and U16115 (N_16115,N_15291,N_15199);
and U16116 (N_16116,N_15292,N_15613);
xor U16117 (N_16117,N_15819,N_15758);
or U16118 (N_16118,N_15954,N_15146);
nand U16119 (N_16119,N_15840,N_15345);
xnor U16120 (N_16120,N_15697,N_15671);
and U16121 (N_16121,N_15121,N_15427);
xnor U16122 (N_16122,N_15087,N_15916);
or U16123 (N_16123,N_15243,N_15203);
or U16124 (N_16124,N_15776,N_15220);
or U16125 (N_16125,N_15164,N_15920);
and U16126 (N_16126,N_15038,N_15690);
or U16127 (N_16127,N_15075,N_15035);
nand U16128 (N_16128,N_15967,N_15564);
nor U16129 (N_16129,N_15435,N_15809);
and U16130 (N_16130,N_15602,N_15414);
or U16131 (N_16131,N_15069,N_15914);
xor U16132 (N_16132,N_15363,N_15702);
nand U16133 (N_16133,N_15794,N_15265);
or U16134 (N_16134,N_15378,N_15887);
or U16135 (N_16135,N_15724,N_15299);
nor U16136 (N_16136,N_15351,N_15154);
nand U16137 (N_16137,N_15060,N_15535);
xnor U16138 (N_16138,N_15717,N_15557);
xnor U16139 (N_16139,N_15793,N_15011);
nor U16140 (N_16140,N_15156,N_15431);
or U16141 (N_16141,N_15975,N_15999);
or U16142 (N_16142,N_15641,N_15869);
nor U16143 (N_16143,N_15935,N_15751);
nand U16144 (N_16144,N_15940,N_15515);
xor U16145 (N_16145,N_15680,N_15919);
and U16146 (N_16146,N_15499,N_15942);
nor U16147 (N_16147,N_15328,N_15692);
or U16148 (N_16148,N_15285,N_15453);
nand U16149 (N_16149,N_15910,N_15709);
nor U16150 (N_16150,N_15895,N_15741);
or U16151 (N_16151,N_15092,N_15130);
or U16152 (N_16152,N_15993,N_15501);
or U16153 (N_16153,N_15281,N_15437);
xnor U16154 (N_16154,N_15517,N_15616);
nor U16155 (N_16155,N_15555,N_15700);
or U16156 (N_16156,N_15797,N_15167);
xnor U16157 (N_16157,N_15685,N_15210);
and U16158 (N_16158,N_15004,N_15917);
or U16159 (N_16159,N_15150,N_15796);
nor U16160 (N_16160,N_15109,N_15932);
and U16161 (N_16161,N_15018,N_15542);
nand U16162 (N_16162,N_15347,N_15127);
xor U16163 (N_16163,N_15523,N_15316);
xnor U16164 (N_16164,N_15178,N_15528);
and U16165 (N_16165,N_15880,N_15817);
xnor U16166 (N_16166,N_15461,N_15286);
nand U16167 (N_16167,N_15737,N_15468);
and U16168 (N_16168,N_15024,N_15478);
nand U16169 (N_16169,N_15956,N_15413);
nand U16170 (N_16170,N_15652,N_15074);
nand U16171 (N_16171,N_15456,N_15832);
or U16172 (N_16172,N_15614,N_15088);
xnor U16173 (N_16173,N_15283,N_15174);
or U16174 (N_16174,N_15370,N_15313);
xor U16175 (N_16175,N_15567,N_15309);
and U16176 (N_16176,N_15790,N_15953);
xor U16177 (N_16177,N_15225,N_15168);
nor U16178 (N_16178,N_15410,N_15679);
nand U16179 (N_16179,N_15958,N_15481);
nor U16180 (N_16180,N_15808,N_15647);
nor U16181 (N_16181,N_15531,N_15572);
nand U16182 (N_16182,N_15989,N_15612);
nand U16183 (N_16183,N_15782,N_15476);
and U16184 (N_16184,N_15886,N_15333);
or U16185 (N_16185,N_15714,N_15444);
nor U16186 (N_16186,N_15250,N_15157);
or U16187 (N_16187,N_15076,N_15093);
and U16188 (N_16188,N_15222,N_15202);
and U16189 (N_16189,N_15102,N_15145);
and U16190 (N_16190,N_15417,N_15899);
and U16191 (N_16191,N_15361,N_15262);
and U16192 (N_16192,N_15021,N_15270);
and U16193 (N_16193,N_15997,N_15279);
nor U16194 (N_16194,N_15244,N_15272);
and U16195 (N_16195,N_15675,N_15386);
nand U16196 (N_16196,N_15195,N_15477);
and U16197 (N_16197,N_15379,N_15100);
xnor U16198 (N_16198,N_15198,N_15148);
or U16199 (N_16199,N_15177,N_15470);
and U16200 (N_16200,N_15115,N_15554);
nor U16201 (N_16201,N_15510,N_15595);
or U16202 (N_16202,N_15664,N_15239);
and U16203 (N_16203,N_15040,N_15332);
nand U16204 (N_16204,N_15046,N_15223);
or U16205 (N_16205,N_15182,N_15604);
nand U16206 (N_16206,N_15189,N_15619);
and U16207 (N_16207,N_15732,N_15504);
nor U16208 (N_16208,N_15736,N_15017);
or U16209 (N_16209,N_15930,N_15814);
or U16210 (N_16210,N_15112,N_15393);
nor U16211 (N_16211,N_15699,N_15259);
nand U16212 (N_16212,N_15205,N_15850);
nand U16213 (N_16213,N_15051,N_15352);
nand U16214 (N_16214,N_15082,N_15563);
nor U16215 (N_16215,N_15329,N_15990);
or U16216 (N_16216,N_15972,N_15095);
and U16217 (N_16217,N_15037,N_15357);
nand U16218 (N_16218,N_15394,N_15067);
nor U16219 (N_16219,N_15893,N_15623);
or U16220 (N_16220,N_15349,N_15951);
xor U16221 (N_16221,N_15933,N_15043);
nand U16222 (N_16222,N_15103,N_15380);
nand U16223 (N_16223,N_15231,N_15509);
nor U16224 (N_16224,N_15518,N_15310);
and U16225 (N_16225,N_15491,N_15358);
or U16226 (N_16226,N_15142,N_15735);
nand U16227 (N_16227,N_15465,N_15443);
nor U16228 (N_16228,N_15396,N_15597);
nand U16229 (N_16229,N_15549,N_15113);
nor U16230 (N_16230,N_15988,N_15625);
or U16231 (N_16231,N_15734,N_15464);
xor U16232 (N_16232,N_15946,N_15192);
and U16233 (N_16233,N_15851,N_15254);
nor U16234 (N_16234,N_15096,N_15754);
or U16235 (N_16235,N_15591,N_15373);
and U16236 (N_16236,N_15209,N_15622);
nor U16237 (N_16237,N_15948,N_15752);
and U16238 (N_16238,N_15511,N_15175);
nor U16239 (N_16239,N_15350,N_15725);
and U16240 (N_16240,N_15158,N_15828);
nor U16241 (N_16241,N_15450,N_15774);
nand U16242 (N_16242,N_15526,N_15325);
xnor U16243 (N_16243,N_15267,N_15760);
nor U16244 (N_16244,N_15010,N_15505);
or U16245 (N_16245,N_15241,N_15666);
or U16246 (N_16246,N_15957,N_15648);
nand U16247 (N_16247,N_15059,N_15344);
and U16248 (N_16248,N_15765,N_15442);
nand U16249 (N_16249,N_15620,N_15682);
or U16250 (N_16250,N_15749,N_15883);
or U16251 (N_16251,N_15578,N_15498);
and U16252 (N_16252,N_15862,N_15224);
nand U16253 (N_16253,N_15728,N_15586);
nor U16254 (N_16254,N_15208,N_15269);
or U16255 (N_16255,N_15892,N_15599);
xnor U16256 (N_16256,N_15570,N_15423);
xor U16257 (N_16257,N_15777,N_15908);
xor U16258 (N_16258,N_15573,N_15449);
and U16259 (N_16259,N_15072,N_15063);
or U16260 (N_16260,N_15655,N_15885);
nand U16261 (N_16261,N_15342,N_15798);
xnor U16262 (N_16262,N_15390,N_15377);
and U16263 (N_16263,N_15791,N_15240);
and U16264 (N_16264,N_15419,N_15807);
xor U16265 (N_16265,N_15810,N_15436);
or U16266 (N_16266,N_15366,N_15023);
xnor U16267 (N_16267,N_15766,N_15971);
or U16268 (N_16268,N_15618,N_15140);
and U16269 (N_16269,N_15303,N_15593);
nand U16270 (N_16270,N_15000,N_15803);
xnor U16271 (N_16271,N_15404,N_15090);
and U16272 (N_16272,N_15343,N_15054);
xnor U16273 (N_16273,N_15950,N_15924);
and U16274 (N_16274,N_15317,N_15677);
and U16275 (N_16275,N_15171,N_15246);
or U16276 (N_16276,N_15994,N_15961);
nand U16277 (N_16277,N_15827,N_15787);
xnor U16278 (N_16278,N_15125,N_15846);
xnor U16279 (N_16279,N_15107,N_15743);
nand U16280 (N_16280,N_15128,N_15490);
nand U16281 (N_16281,N_15764,N_15600);
nor U16282 (N_16282,N_15581,N_15248);
nand U16283 (N_16283,N_15878,N_15098);
or U16284 (N_16284,N_15039,N_15847);
xnor U16285 (N_16285,N_15080,N_15966);
xor U16286 (N_16286,N_15007,N_15141);
nor U16287 (N_16287,N_15275,N_15376);
or U16288 (N_16288,N_15617,N_15806);
or U16289 (N_16289,N_15138,N_15326);
nor U16290 (N_16290,N_15529,N_15191);
and U16291 (N_16291,N_15658,N_15816);
xor U16292 (N_16292,N_15514,N_15731);
nor U16293 (N_16293,N_15605,N_15973);
xnor U16294 (N_16294,N_15854,N_15704);
xnor U16295 (N_16295,N_15462,N_15302);
nor U16296 (N_16296,N_15402,N_15978);
and U16297 (N_16297,N_15943,N_15287);
xnor U16298 (N_16298,N_15962,N_15538);
nand U16299 (N_16299,N_15083,N_15318);
and U16300 (N_16300,N_15253,N_15383);
or U16301 (N_16301,N_15346,N_15718);
and U16302 (N_16302,N_15922,N_15305);
nor U16303 (N_16303,N_15562,N_15196);
or U16304 (N_16304,N_15364,N_15921);
or U16305 (N_16305,N_15756,N_15659);
nor U16306 (N_16306,N_15853,N_15762);
xor U16307 (N_16307,N_15073,N_15136);
and U16308 (N_16308,N_15610,N_15475);
nand U16309 (N_16309,N_15061,N_15266);
nand U16310 (N_16310,N_15670,N_15753);
xnor U16311 (N_16311,N_15455,N_15715);
or U16312 (N_16312,N_15022,N_15238);
and U16313 (N_16313,N_15172,N_15295);
xnor U16314 (N_16314,N_15258,N_15842);
nand U16315 (N_16315,N_15277,N_15980);
nor U16316 (N_16316,N_15923,N_15474);
xnor U16317 (N_16317,N_15110,N_15385);
xor U16318 (N_16318,N_15733,N_15500);
and U16319 (N_16319,N_15874,N_15508);
or U16320 (N_16320,N_15050,N_15643);
and U16321 (N_16321,N_15965,N_15173);
nor U16322 (N_16322,N_15712,N_15746);
nand U16323 (N_16323,N_15482,N_15307);
or U16324 (N_16324,N_15949,N_15492);
nand U16325 (N_16325,N_15058,N_15985);
nor U16326 (N_16326,N_15594,N_15274);
nor U16327 (N_16327,N_15589,N_15582);
nand U16328 (N_16328,N_15057,N_15337);
nor U16329 (N_16329,N_15424,N_15770);
and U16330 (N_16330,N_15566,N_15739);
nand U16331 (N_16331,N_15152,N_15545);
or U16332 (N_16332,N_15865,N_15237);
nor U16333 (N_16333,N_15708,N_15466);
nor U16334 (N_16334,N_15875,N_15696);
or U16335 (N_16335,N_15742,N_15727);
nor U16336 (N_16336,N_15234,N_15162);
nand U16337 (N_16337,N_15496,N_15306);
or U16338 (N_16338,N_15915,N_15608);
and U16339 (N_16339,N_15016,N_15015);
or U16340 (N_16340,N_15179,N_15212);
or U16341 (N_16341,N_15907,N_15800);
xnor U16342 (N_16342,N_15360,N_15849);
and U16343 (N_16343,N_15147,N_15160);
xor U16344 (N_16344,N_15123,N_15354);
or U16345 (N_16345,N_15638,N_15969);
nand U16346 (N_16346,N_15568,N_15982);
nor U16347 (N_16347,N_15836,N_15506);
or U16348 (N_16348,N_15632,N_15844);
and U16349 (N_16349,N_15665,N_15339);
nor U16350 (N_16350,N_15454,N_15249);
nor U16351 (N_16351,N_15502,N_15432);
nand U16352 (N_16352,N_15190,N_15071);
or U16353 (N_16353,N_15027,N_15489);
and U16354 (N_16354,N_15165,N_15522);
xnor U16355 (N_16355,N_15045,N_15775);
and U16356 (N_16356,N_15235,N_15681);
nor U16357 (N_16357,N_15479,N_15228);
nor U16358 (N_16358,N_15183,N_15389);
and U16359 (N_16359,N_15221,N_15541);
nand U16360 (N_16360,N_15089,N_15169);
and U16361 (N_16361,N_15579,N_15304);
nand U16362 (N_16362,N_15085,N_15822);
or U16363 (N_16363,N_15484,N_15628);
and U16364 (N_16364,N_15968,N_15187);
xnor U16365 (N_16365,N_15388,N_15547);
xor U16366 (N_16366,N_15392,N_15571);
xnor U16367 (N_16367,N_15560,N_15544);
xnor U16368 (N_16368,N_15003,N_15780);
xnor U16369 (N_16369,N_15795,N_15336);
nand U16370 (N_16370,N_15646,N_15483);
and U16371 (N_16371,N_15371,N_15227);
and U16372 (N_16372,N_15374,N_15384);
nor U16373 (N_16373,N_15001,N_15654);
nand U16374 (N_16374,N_15748,N_15425);
or U16375 (N_16375,N_15002,N_15348);
nand U16376 (N_16376,N_15028,N_15251);
nor U16377 (N_16377,N_15034,N_15226);
xnor U16378 (N_16378,N_15340,N_15955);
nor U16379 (N_16379,N_15722,N_15799);
xor U16380 (N_16380,N_15452,N_15132);
and U16381 (N_16381,N_15788,N_15559);
xnor U16382 (N_16382,N_15186,N_15230);
or U16383 (N_16383,N_15245,N_15903);
and U16384 (N_16384,N_15293,N_15757);
and U16385 (N_16385,N_15369,N_15042);
xor U16386 (N_16386,N_15979,N_15252);
nor U16387 (N_16387,N_15323,N_15918);
nor U16388 (N_16388,N_15884,N_15312);
nor U16389 (N_16389,N_15268,N_15660);
and U16390 (N_16390,N_15928,N_15315);
xnor U16391 (N_16391,N_15064,N_15826);
or U16392 (N_16392,N_15848,N_15428);
xor U16393 (N_16393,N_15642,N_15433);
and U16394 (N_16394,N_15552,N_15911);
nor U16395 (N_16395,N_15401,N_15992);
and U16396 (N_16396,N_15867,N_15860);
nand U16397 (N_16397,N_15006,N_15008);
nor U16398 (N_16398,N_15835,N_15153);
xor U16399 (N_16399,N_15941,N_15144);
and U16400 (N_16400,N_15905,N_15863);
nor U16401 (N_16401,N_15519,N_15513);
nor U16402 (N_16402,N_15588,N_15672);
nand U16403 (N_16403,N_15667,N_15242);
nor U16404 (N_16404,N_15626,N_15084);
xnor U16405 (N_16405,N_15447,N_15439);
and U16406 (N_16406,N_15105,N_15135);
nor U16407 (N_16407,N_15640,N_15609);
nand U16408 (N_16408,N_15527,N_15536);
nand U16409 (N_16409,N_15407,N_15651);
nor U16410 (N_16410,N_15759,N_15485);
xor U16411 (N_16411,N_15503,N_15897);
xor U16412 (N_16412,N_15583,N_15256);
or U16413 (N_16413,N_15434,N_15634);
xor U16414 (N_16414,N_15200,N_15236);
and U16415 (N_16415,N_15569,N_15580);
or U16416 (N_16416,N_15426,N_15927);
and U16417 (N_16417,N_15355,N_15119);
nand U16418 (N_16418,N_15805,N_15446);
or U16419 (N_16419,N_15289,N_15841);
xnor U16420 (N_16420,N_15163,N_15684);
nor U16421 (N_16421,N_15441,N_15653);
nand U16422 (N_16422,N_15871,N_15539);
xnor U16423 (N_16423,N_15297,N_15845);
nor U16424 (N_16424,N_15372,N_15768);
nor U16425 (N_16425,N_15260,N_15676);
nand U16426 (N_16426,N_15282,N_15459);
nand U16427 (N_16427,N_15730,N_15211);
nor U16428 (N_16428,N_15778,N_15009);
xnor U16429 (N_16429,N_15894,N_15012);
nand U16430 (N_16430,N_15804,N_15558);
nand U16431 (N_16431,N_15986,N_15458);
or U16432 (N_16432,N_15341,N_15710);
nor U16433 (N_16433,N_15607,N_15099);
nand U16434 (N_16434,N_15273,N_15769);
and U16435 (N_16435,N_15457,N_15233);
nor U16436 (N_16436,N_15217,N_15321);
and U16437 (N_16437,N_15086,N_15106);
or U16438 (N_16438,N_15382,N_15487);
xnor U16439 (N_16439,N_15081,N_15151);
nand U16440 (N_16440,N_15711,N_15931);
or U16441 (N_16441,N_15693,N_15723);
xor U16442 (N_16442,N_15311,N_15719);
nand U16443 (N_16443,N_15645,N_15271);
xnor U16444 (N_16444,N_15852,N_15036);
and U16445 (N_16445,N_15155,N_15548);
nor U16446 (N_16446,N_15020,N_15362);
nand U16447 (N_16447,N_15983,N_15194);
or U16448 (N_16448,N_15320,N_15319);
nor U16449 (N_16449,N_15255,N_15104);
nor U16450 (N_16450,N_15422,N_15631);
nor U16451 (N_16451,N_15334,N_15534);
and U16452 (N_16452,N_15771,N_15603);
xnor U16453 (N_16453,N_15937,N_15430);
nand U16454 (N_16454,N_15785,N_15621);
xor U16455 (N_16455,N_15381,N_15598);
nor U16456 (N_16456,N_15368,N_15726);
and U16457 (N_16457,N_15945,N_15929);
nor U16458 (N_16458,N_15637,N_15215);
nor U16459 (N_16459,N_15611,N_15143);
xor U16460 (N_16460,N_15936,N_15495);
and U16461 (N_16461,N_15056,N_15469);
or U16462 (N_16462,N_15219,N_15537);
and U16463 (N_16463,N_15601,N_15974);
and U16464 (N_16464,N_15472,N_15984);
nor U16465 (N_16465,N_15868,N_15129);
nand U16466 (N_16466,N_15755,N_15551);
and U16467 (N_16467,N_15981,N_15902);
xor U16468 (N_16468,N_15877,N_15264);
or U16469 (N_16469,N_15124,N_15821);
or U16470 (N_16470,N_15830,N_15668);
or U16471 (N_16471,N_15801,N_15705);
or U16472 (N_16472,N_15048,N_15213);
xnor U16473 (N_16473,N_15615,N_15713);
nor U16474 (N_16474,N_15976,N_15448);
or U16475 (N_16475,N_15729,N_15391);
xnor U16476 (N_16476,N_15698,N_15276);
and U16477 (N_16477,N_15029,N_15823);
xnor U16478 (N_16478,N_15701,N_15818);
xor U16479 (N_16479,N_15996,N_15939);
and U16480 (N_16480,N_15159,N_15327);
or U16481 (N_16481,N_15689,N_15574);
xor U16482 (N_16482,N_15678,N_15176);
and U16483 (N_16483,N_15257,N_15507);
and U16484 (N_16484,N_15738,N_15065);
nor U16485 (N_16485,N_15872,N_15649);
nor U16486 (N_16486,N_15324,N_15180);
and U16487 (N_16487,N_15635,N_15802);
or U16488 (N_16488,N_15261,N_15232);
nor U16489 (N_16489,N_15889,N_15471);
xor U16490 (N_16490,N_15767,N_15026);
xnor U16491 (N_16491,N_15858,N_15118);
and U16492 (N_16492,N_15556,N_15873);
and U16493 (N_16493,N_15330,N_15131);
and U16494 (N_16494,N_15044,N_15543);
nand U16495 (N_16495,N_15134,N_15553);
nor U16496 (N_16496,N_15856,N_15686);
and U16497 (N_16497,N_15139,N_15744);
and U16498 (N_16498,N_15052,N_15418);
nand U16499 (N_16499,N_15636,N_15650);
or U16500 (N_16500,N_15548,N_15126);
xnor U16501 (N_16501,N_15767,N_15059);
or U16502 (N_16502,N_15852,N_15610);
nand U16503 (N_16503,N_15164,N_15497);
and U16504 (N_16504,N_15613,N_15909);
and U16505 (N_16505,N_15296,N_15496);
and U16506 (N_16506,N_15891,N_15373);
nor U16507 (N_16507,N_15966,N_15933);
or U16508 (N_16508,N_15207,N_15815);
nor U16509 (N_16509,N_15154,N_15247);
nor U16510 (N_16510,N_15070,N_15743);
nor U16511 (N_16511,N_15404,N_15742);
and U16512 (N_16512,N_15415,N_15044);
nand U16513 (N_16513,N_15238,N_15981);
nor U16514 (N_16514,N_15367,N_15531);
and U16515 (N_16515,N_15575,N_15571);
xnor U16516 (N_16516,N_15336,N_15581);
or U16517 (N_16517,N_15583,N_15020);
xnor U16518 (N_16518,N_15891,N_15149);
xnor U16519 (N_16519,N_15337,N_15178);
or U16520 (N_16520,N_15003,N_15697);
nor U16521 (N_16521,N_15484,N_15054);
nor U16522 (N_16522,N_15290,N_15288);
or U16523 (N_16523,N_15919,N_15911);
xor U16524 (N_16524,N_15811,N_15353);
or U16525 (N_16525,N_15203,N_15800);
and U16526 (N_16526,N_15266,N_15020);
and U16527 (N_16527,N_15888,N_15790);
xor U16528 (N_16528,N_15880,N_15690);
or U16529 (N_16529,N_15887,N_15327);
nand U16530 (N_16530,N_15049,N_15116);
or U16531 (N_16531,N_15160,N_15958);
xnor U16532 (N_16532,N_15377,N_15474);
or U16533 (N_16533,N_15706,N_15438);
or U16534 (N_16534,N_15368,N_15709);
nor U16535 (N_16535,N_15515,N_15959);
nor U16536 (N_16536,N_15074,N_15738);
xor U16537 (N_16537,N_15722,N_15042);
nor U16538 (N_16538,N_15443,N_15562);
xor U16539 (N_16539,N_15977,N_15588);
nor U16540 (N_16540,N_15451,N_15518);
nor U16541 (N_16541,N_15366,N_15723);
and U16542 (N_16542,N_15413,N_15481);
and U16543 (N_16543,N_15543,N_15491);
or U16544 (N_16544,N_15020,N_15399);
nor U16545 (N_16545,N_15856,N_15890);
and U16546 (N_16546,N_15520,N_15628);
or U16547 (N_16547,N_15599,N_15468);
nor U16548 (N_16548,N_15233,N_15381);
and U16549 (N_16549,N_15900,N_15690);
nor U16550 (N_16550,N_15789,N_15355);
nor U16551 (N_16551,N_15500,N_15767);
nor U16552 (N_16552,N_15055,N_15156);
nand U16553 (N_16553,N_15542,N_15517);
or U16554 (N_16554,N_15991,N_15891);
or U16555 (N_16555,N_15974,N_15862);
or U16556 (N_16556,N_15718,N_15525);
and U16557 (N_16557,N_15059,N_15227);
nand U16558 (N_16558,N_15473,N_15812);
nand U16559 (N_16559,N_15639,N_15304);
and U16560 (N_16560,N_15081,N_15801);
xor U16561 (N_16561,N_15304,N_15554);
and U16562 (N_16562,N_15212,N_15282);
xnor U16563 (N_16563,N_15744,N_15307);
nand U16564 (N_16564,N_15879,N_15910);
nand U16565 (N_16565,N_15533,N_15134);
and U16566 (N_16566,N_15227,N_15274);
and U16567 (N_16567,N_15995,N_15594);
nor U16568 (N_16568,N_15711,N_15229);
xor U16569 (N_16569,N_15660,N_15909);
xor U16570 (N_16570,N_15050,N_15182);
and U16571 (N_16571,N_15047,N_15924);
or U16572 (N_16572,N_15936,N_15455);
and U16573 (N_16573,N_15492,N_15454);
xnor U16574 (N_16574,N_15617,N_15911);
nand U16575 (N_16575,N_15617,N_15079);
nand U16576 (N_16576,N_15005,N_15540);
xnor U16577 (N_16577,N_15710,N_15709);
nand U16578 (N_16578,N_15059,N_15412);
and U16579 (N_16579,N_15663,N_15651);
or U16580 (N_16580,N_15436,N_15210);
nor U16581 (N_16581,N_15775,N_15772);
nand U16582 (N_16582,N_15753,N_15116);
nor U16583 (N_16583,N_15725,N_15417);
and U16584 (N_16584,N_15967,N_15348);
and U16585 (N_16585,N_15449,N_15476);
or U16586 (N_16586,N_15344,N_15390);
and U16587 (N_16587,N_15172,N_15873);
xor U16588 (N_16588,N_15594,N_15536);
nand U16589 (N_16589,N_15066,N_15212);
and U16590 (N_16590,N_15651,N_15707);
and U16591 (N_16591,N_15418,N_15337);
and U16592 (N_16592,N_15669,N_15431);
nor U16593 (N_16593,N_15844,N_15300);
nor U16594 (N_16594,N_15170,N_15444);
or U16595 (N_16595,N_15780,N_15105);
nor U16596 (N_16596,N_15007,N_15247);
and U16597 (N_16597,N_15424,N_15297);
nand U16598 (N_16598,N_15421,N_15885);
nor U16599 (N_16599,N_15547,N_15736);
or U16600 (N_16600,N_15723,N_15433);
xor U16601 (N_16601,N_15814,N_15134);
nand U16602 (N_16602,N_15350,N_15875);
nand U16603 (N_16603,N_15783,N_15173);
nand U16604 (N_16604,N_15579,N_15451);
and U16605 (N_16605,N_15172,N_15331);
xnor U16606 (N_16606,N_15914,N_15755);
nor U16607 (N_16607,N_15918,N_15781);
xor U16608 (N_16608,N_15116,N_15949);
or U16609 (N_16609,N_15114,N_15676);
nand U16610 (N_16610,N_15644,N_15661);
and U16611 (N_16611,N_15162,N_15720);
and U16612 (N_16612,N_15122,N_15078);
xnor U16613 (N_16613,N_15431,N_15754);
nor U16614 (N_16614,N_15690,N_15520);
nor U16615 (N_16615,N_15504,N_15424);
xnor U16616 (N_16616,N_15832,N_15551);
xor U16617 (N_16617,N_15658,N_15352);
xor U16618 (N_16618,N_15305,N_15242);
or U16619 (N_16619,N_15859,N_15960);
nand U16620 (N_16620,N_15088,N_15547);
xnor U16621 (N_16621,N_15780,N_15014);
nor U16622 (N_16622,N_15596,N_15445);
or U16623 (N_16623,N_15783,N_15184);
or U16624 (N_16624,N_15827,N_15281);
nor U16625 (N_16625,N_15029,N_15870);
or U16626 (N_16626,N_15559,N_15088);
xor U16627 (N_16627,N_15093,N_15286);
nand U16628 (N_16628,N_15370,N_15794);
and U16629 (N_16629,N_15680,N_15264);
nand U16630 (N_16630,N_15473,N_15510);
or U16631 (N_16631,N_15594,N_15358);
xor U16632 (N_16632,N_15237,N_15194);
xor U16633 (N_16633,N_15090,N_15231);
or U16634 (N_16634,N_15178,N_15056);
nor U16635 (N_16635,N_15779,N_15611);
nand U16636 (N_16636,N_15507,N_15017);
xor U16637 (N_16637,N_15106,N_15545);
or U16638 (N_16638,N_15616,N_15003);
nor U16639 (N_16639,N_15591,N_15161);
or U16640 (N_16640,N_15254,N_15315);
xnor U16641 (N_16641,N_15694,N_15213);
and U16642 (N_16642,N_15461,N_15028);
and U16643 (N_16643,N_15310,N_15991);
xor U16644 (N_16644,N_15002,N_15544);
nand U16645 (N_16645,N_15305,N_15698);
or U16646 (N_16646,N_15643,N_15990);
xnor U16647 (N_16647,N_15625,N_15026);
and U16648 (N_16648,N_15837,N_15188);
or U16649 (N_16649,N_15490,N_15695);
and U16650 (N_16650,N_15356,N_15012);
and U16651 (N_16651,N_15134,N_15938);
nor U16652 (N_16652,N_15856,N_15971);
or U16653 (N_16653,N_15565,N_15045);
xor U16654 (N_16654,N_15826,N_15049);
xnor U16655 (N_16655,N_15841,N_15973);
nand U16656 (N_16656,N_15964,N_15508);
xor U16657 (N_16657,N_15283,N_15987);
or U16658 (N_16658,N_15861,N_15073);
xor U16659 (N_16659,N_15382,N_15702);
nor U16660 (N_16660,N_15756,N_15609);
nand U16661 (N_16661,N_15769,N_15340);
and U16662 (N_16662,N_15037,N_15004);
nor U16663 (N_16663,N_15729,N_15067);
or U16664 (N_16664,N_15320,N_15368);
nor U16665 (N_16665,N_15209,N_15513);
nor U16666 (N_16666,N_15729,N_15825);
xor U16667 (N_16667,N_15018,N_15944);
nor U16668 (N_16668,N_15075,N_15918);
and U16669 (N_16669,N_15429,N_15381);
or U16670 (N_16670,N_15313,N_15310);
xnor U16671 (N_16671,N_15087,N_15121);
and U16672 (N_16672,N_15942,N_15342);
and U16673 (N_16673,N_15481,N_15864);
and U16674 (N_16674,N_15594,N_15024);
nor U16675 (N_16675,N_15901,N_15276);
and U16676 (N_16676,N_15167,N_15787);
and U16677 (N_16677,N_15915,N_15005);
xor U16678 (N_16678,N_15429,N_15773);
and U16679 (N_16679,N_15170,N_15200);
or U16680 (N_16680,N_15189,N_15391);
xnor U16681 (N_16681,N_15060,N_15558);
and U16682 (N_16682,N_15613,N_15367);
xor U16683 (N_16683,N_15367,N_15832);
nand U16684 (N_16684,N_15095,N_15590);
or U16685 (N_16685,N_15336,N_15356);
or U16686 (N_16686,N_15629,N_15687);
or U16687 (N_16687,N_15512,N_15147);
nand U16688 (N_16688,N_15448,N_15435);
or U16689 (N_16689,N_15305,N_15298);
nand U16690 (N_16690,N_15751,N_15991);
nand U16691 (N_16691,N_15025,N_15588);
xnor U16692 (N_16692,N_15311,N_15078);
nand U16693 (N_16693,N_15611,N_15901);
or U16694 (N_16694,N_15442,N_15416);
nor U16695 (N_16695,N_15176,N_15540);
and U16696 (N_16696,N_15826,N_15188);
xor U16697 (N_16697,N_15239,N_15078);
or U16698 (N_16698,N_15601,N_15620);
and U16699 (N_16699,N_15805,N_15292);
xor U16700 (N_16700,N_15078,N_15968);
and U16701 (N_16701,N_15009,N_15821);
or U16702 (N_16702,N_15889,N_15112);
nor U16703 (N_16703,N_15723,N_15694);
nor U16704 (N_16704,N_15158,N_15177);
xnor U16705 (N_16705,N_15228,N_15734);
nor U16706 (N_16706,N_15222,N_15804);
nand U16707 (N_16707,N_15775,N_15777);
nand U16708 (N_16708,N_15630,N_15892);
nand U16709 (N_16709,N_15479,N_15951);
xnor U16710 (N_16710,N_15234,N_15875);
or U16711 (N_16711,N_15712,N_15234);
nand U16712 (N_16712,N_15185,N_15240);
or U16713 (N_16713,N_15304,N_15134);
nand U16714 (N_16714,N_15285,N_15326);
or U16715 (N_16715,N_15830,N_15144);
or U16716 (N_16716,N_15825,N_15434);
nor U16717 (N_16717,N_15000,N_15768);
nand U16718 (N_16718,N_15848,N_15855);
nand U16719 (N_16719,N_15423,N_15523);
xnor U16720 (N_16720,N_15671,N_15211);
or U16721 (N_16721,N_15701,N_15631);
nor U16722 (N_16722,N_15208,N_15677);
xor U16723 (N_16723,N_15953,N_15820);
nor U16724 (N_16724,N_15195,N_15094);
xnor U16725 (N_16725,N_15775,N_15950);
nor U16726 (N_16726,N_15080,N_15366);
nor U16727 (N_16727,N_15875,N_15519);
or U16728 (N_16728,N_15883,N_15967);
nor U16729 (N_16729,N_15252,N_15922);
nor U16730 (N_16730,N_15595,N_15252);
or U16731 (N_16731,N_15256,N_15302);
xor U16732 (N_16732,N_15921,N_15992);
or U16733 (N_16733,N_15486,N_15316);
nor U16734 (N_16734,N_15721,N_15122);
and U16735 (N_16735,N_15278,N_15566);
or U16736 (N_16736,N_15551,N_15447);
xor U16737 (N_16737,N_15118,N_15385);
nor U16738 (N_16738,N_15367,N_15195);
and U16739 (N_16739,N_15962,N_15010);
or U16740 (N_16740,N_15482,N_15979);
nor U16741 (N_16741,N_15482,N_15173);
xor U16742 (N_16742,N_15369,N_15300);
nor U16743 (N_16743,N_15666,N_15579);
nor U16744 (N_16744,N_15137,N_15847);
and U16745 (N_16745,N_15865,N_15324);
nor U16746 (N_16746,N_15265,N_15981);
nor U16747 (N_16747,N_15886,N_15588);
and U16748 (N_16748,N_15742,N_15573);
nor U16749 (N_16749,N_15984,N_15700);
and U16750 (N_16750,N_15108,N_15828);
xnor U16751 (N_16751,N_15888,N_15952);
nand U16752 (N_16752,N_15939,N_15477);
xor U16753 (N_16753,N_15176,N_15503);
and U16754 (N_16754,N_15353,N_15102);
and U16755 (N_16755,N_15925,N_15365);
xnor U16756 (N_16756,N_15573,N_15695);
and U16757 (N_16757,N_15576,N_15608);
or U16758 (N_16758,N_15278,N_15793);
nor U16759 (N_16759,N_15797,N_15976);
nor U16760 (N_16760,N_15549,N_15354);
nand U16761 (N_16761,N_15228,N_15251);
xnor U16762 (N_16762,N_15440,N_15007);
or U16763 (N_16763,N_15646,N_15130);
xor U16764 (N_16764,N_15035,N_15808);
nand U16765 (N_16765,N_15051,N_15370);
nor U16766 (N_16766,N_15953,N_15092);
xor U16767 (N_16767,N_15621,N_15997);
or U16768 (N_16768,N_15147,N_15851);
nand U16769 (N_16769,N_15796,N_15497);
xnor U16770 (N_16770,N_15753,N_15609);
and U16771 (N_16771,N_15871,N_15507);
and U16772 (N_16772,N_15501,N_15861);
nor U16773 (N_16773,N_15441,N_15845);
or U16774 (N_16774,N_15100,N_15463);
and U16775 (N_16775,N_15792,N_15308);
nand U16776 (N_16776,N_15663,N_15877);
nor U16777 (N_16777,N_15469,N_15081);
nand U16778 (N_16778,N_15095,N_15126);
or U16779 (N_16779,N_15434,N_15909);
or U16780 (N_16780,N_15976,N_15896);
nand U16781 (N_16781,N_15082,N_15245);
and U16782 (N_16782,N_15232,N_15551);
xnor U16783 (N_16783,N_15912,N_15262);
and U16784 (N_16784,N_15335,N_15433);
xnor U16785 (N_16785,N_15430,N_15083);
xor U16786 (N_16786,N_15023,N_15677);
or U16787 (N_16787,N_15397,N_15302);
nand U16788 (N_16788,N_15026,N_15362);
and U16789 (N_16789,N_15085,N_15267);
nand U16790 (N_16790,N_15044,N_15236);
nor U16791 (N_16791,N_15847,N_15601);
and U16792 (N_16792,N_15357,N_15078);
nand U16793 (N_16793,N_15143,N_15941);
and U16794 (N_16794,N_15655,N_15676);
nor U16795 (N_16795,N_15326,N_15411);
and U16796 (N_16796,N_15536,N_15901);
and U16797 (N_16797,N_15233,N_15043);
xor U16798 (N_16798,N_15259,N_15197);
and U16799 (N_16799,N_15003,N_15242);
xor U16800 (N_16800,N_15473,N_15435);
xor U16801 (N_16801,N_15118,N_15084);
nand U16802 (N_16802,N_15185,N_15313);
nand U16803 (N_16803,N_15586,N_15867);
and U16804 (N_16804,N_15661,N_15200);
nor U16805 (N_16805,N_15914,N_15047);
or U16806 (N_16806,N_15625,N_15326);
nand U16807 (N_16807,N_15093,N_15376);
nand U16808 (N_16808,N_15202,N_15245);
or U16809 (N_16809,N_15074,N_15865);
or U16810 (N_16810,N_15737,N_15775);
or U16811 (N_16811,N_15901,N_15420);
and U16812 (N_16812,N_15399,N_15663);
nor U16813 (N_16813,N_15219,N_15312);
nand U16814 (N_16814,N_15203,N_15720);
nor U16815 (N_16815,N_15565,N_15449);
nor U16816 (N_16816,N_15902,N_15632);
nor U16817 (N_16817,N_15243,N_15557);
xor U16818 (N_16818,N_15476,N_15863);
and U16819 (N_16819,N_15347,N_15433);
nor U16820 (N_16820,N_15309,N_15116);
or U16821 (N_16821,N_15692,N_15091);
nor U16822 (N_16822,N_15202,N_15371);
and U16823 (N_16823,N_15307,N_15806);
xnor U16824 (N_16824,N_15003,N_15130);
xor U16825 (N_16825,N_15202,N_15850);
nand U16826 (N_16826,N_15145,N_15398);
nand U16827 (N_16827,N_15335,N_15365);
nand U16828 (N_16828,N_15967,N_15833);
nand U16829 (N_16829,N_15326,N_15007);
nand U16830 (N_16830,N_15406,N_15597);
xor U16831 (N_16831,N_15485,N_15577);
and U16832 (N_16832,N_15153,N_15814);
nor U16833 (N_16833,N_15214,N_15682);
xnor U16834 (N_16834,N_15581,N_15069);
nor U16835 (N_16835,N_15109,N_15453);
nor U16836 (N_16836,N_15751,N_15994);
or U16837 (N_16837,N_15470,N_15337);
xnor U16838 (N_16838,N_15984,N_15448);
nand U16839 (N_16839,N_15303,N_15078);
xor U16840 (N_16840,N_15936,N_15119);
xor U16841 (N_16841,N_15318,N_15094);
nor U16842 (N_16842,N_15869,N_15176);
xnor U16843 (N_16843,N_15949,N_15764);
or U16844 (N_16844,N_15344,N_15084);
and U16845 (N_16845,N_15964,N_15297);
nor U16846 (N_16846,N_15999,N_15257);
nor U16847 (N_16847,N_15096,N_15807);
nor U16848 (N_16848,N_15331,N_15324);
or U16849 (N_16849,N_15439,N_15621);
and U16850 (N_16850,N_15128,N_15586);
and U16851 (N_16851,N_15134,N_15238);
xnor U16852 (N_16852,N_15946,N_15199);
and U16853 (N_16853,N_15772,N_15512);
nand U16854 (N_16854,N_15272,N_15333);
nand U16855 (N_16855,N_15907,N_15627);
xor U16856 (N_16856,N_15002,N_15132);
or U16857 (N_16857,N_15678,N_15742);
and U16858 (N_16858,N_15680,N_15831);
or U16859 (N_16859,N_15554,N_15814);
and U16860 (N_16860,N_15014,N_15629);
or U16861 (N_16861,N_15968,N_15423);
and U16862 (N_16862,N_15568,N_15064);
or U16863 (N_16863,N_15351,N_15513);
or U16864 (N_16864,N_15535,N_15583);
xnor U16865 (N_16865,N_15279,N_15303);
nor U16866 (N_16866,N_15067,N_15864);
nor U16867 (N_16867,N_15173,N_15799);
or U16868 (N_16868,N_15910,N_15489);
or U16869 (N_16869,N_15290,N_15692);
and U16870 (N_16870,N_15576,N_15834);
or U16871 (N_16871,N_15764,N_15316);
nand U16872 (N_16872,N_15720,N_15403);
nand U16873 (N_16873,N_15471,N_15329);
and U16874 (N_16874,N_15334,N_15750);
nand U16875 (N_16875,N_15104,N_15528);
nand U16876 (N_16876,N_15899,N_15933);
or U16877 (N_16877,N_15857,N_15719);
nor U16878 (N_16878,N_15056,N_15906);
and U16879 (N_16879,N_15159,N_15726);
or U16880 (N_16880,N_15629,N_15634);
nand U16881 (N_16881,N_15369,N_15343);
nor U16882 (N_16882,N_15357,N_15611);
nor U16883 (N_16883,N_15817,N_15879);
or U16884 (N_16884,N_15119,N_15157);
nor U16885 (N_16885,N_15508,N_15205);
nor U16886 (N_16886,N_15866,N_15809);
or U16887 (N_16887,N_15066,N_15737);
and U16888 (N_16888,N_15367,N_15863);
or U16889 (N_16889,N_15604,N_15636);
nor U16890 (N_16890,N_15125,N_15139);
xnor U16891 (N_16891,N_15738,N_15488);
nor U16892 (N_16892,N_15007,N_15796);
xor U16893 (N_16893,N_15210,N_15630);
and U16894 (N_16894,N_15829,N_15281);
and U16895 (N_16895,N_15701,N_15452);
or U16896 (N_16896,N_15020,N_15089);
nand U16897 (N_16897,N_15004,N_15471);
xnor U16898 (N_16898,N_15709,N_15962);
nand U16899 (N_16899,N_15716,N_15612);
or U16900 (N_16900,N_15743,N_15671);
and U16901 (N_16901,N_15231,N_15473);
nand U16902 (N_16902,N_15474,N_15685);
xnor U16903 (N_16903,N_15607,N_15642);
or U16904 (N_16904,N_15902,N_15638);
nor U16905 (N_16905,N_15612,N_15766);
or U16906 (N_16906,N_15749,N_15028);
nand U16907 (N_16907,N_15628,N_15733);
nor U16908 (N_16908,N_15565,N_15217);
and U16909 (N_16909,N_15197,N_15666);
nand U16910 (N_16910,N_15060,N_15763);
nor U16911 (N_16911,N_15275,N_15147);
xor U16912 (N_16912,N_15953,N_15551);
and U16913 (N_16913,N_15738,N_15861);
nor U16914 (N_16914,N_15607,N_15927);
xnor U16915 (N_16915,N_15597,N_15756);
xnor U16916 (N_16916,N_15629,N_15003);
nand U16917 (N_16917,N_15966,N_15982);
and U16918 (N_16918,N_15690,N_15059);
nand U16919 (N_16919,N_15638,N_15720);
or U16920 (N_16920,N_15078,N_15130);
nand U16921 (N_16921,N_15558,N_15153);
nor U16922 (N_16922,N_15223,N_15545);
nor U16923 (N_16923,N_15182,N_15715);
nand U16924 (N_16924,N_15011,N_15742);
nor U16925 (N_16925,N_15591,N_15786);
nand U16926 (N_16926,N_15259,N_15085);
and U16927 (N_16927,N_15745,N_15998);
or U16928 (N_16928,N_15388,N_15211);
nand U16929 (N_16929,N_15403,N_15007);
and U16930 (N_16930,N_15398,N_15143);
nand U16931 (N_16931,N_15876,N_15018);
xnor U16932 (N_16932,N_15943,N_15556);
nor U16933 (N_16933,N_15853,N_15199);
and U16934 (N_16934,N_15220,N_15528);
or U16935 (N_16935,N_15323,N_15467);
nand U16936 (N_16936,N_15118,N_15953);
or U16937 (N_16937,N_15161,N_15352);
or U16938 (N_16938,N_15711,N_15943);
or U16939 (N_16939,N_15366,N_15629);
nor U16940 (N_16940,N_15051,N_15898);
nand U16941 (N_16941,N_15213,N_15373);
and U16942 (N_16942,N_15428,N_15630);
or U16943 (N_16943,N_15197,N_15236);
and U16944 (N_16944,N_15457,N_15447);
xor U16945 (N_16945,N_15833,N_15461);
and U16946 (N_16946,N_15644,N_15996);
nor U16947 (N_16947,N_15203,N_15837);
nor U16948 (N_16948,N_15341,N_15155);
xor U16949 (N_16949,N_15207,N_15447);
xnor U16950 (N_16950,N_15034,N_15865);
xor U16951 (N_16951,N_15061,N_15149);
xor U16952 (N_16952,N_15770,N_15720);
and U16953 (N_16953,N_15380,N_15479);
nand U16954 (N_16954,N_15674,N_15271);
nor U16955 (N_16955,N_15567,N_15631);
xnor U16956 (N_16956,N_15417,N_15807);
or U16957 (N_16957,N_15294,N_15087);
and U16958 (N_16958,N_15353,N_15311);
and U16959 (N_16959,N_15615,N_15136);
xnor U16960 (N_16960,N_15760,N_15130);
nor U16961 (N_16961,N_15775,N_15750);
and U16962 (N_16962,N_15855,N_15578);
nand U16963 (N_16963,N_15778,N_15988);
nor U16964 (N_16964,N_15001,N_15564);
and U16965 (N_16965,N_15154,N_15443);
nand U16966 (N_16966,N_15336,N_15098);
nand U16967 (N_16967,N_15968,N_15739);
nand U16968 (N_16968,N_15445,N_15530);
or U16969 (N_16969,N_15478,N_15543);
or U16970 (N_16970,N_15497,N_15257);
or U16971 (N_16971,N_15153,N_15300);
nor U16972 (N_16972,N_15017,N_15464);
xor U16973 (N_16973,N_15447,N_15647);
or U16974 (N_16974,N_15701,N_15756);
xor U16975 (N_16975,N_15642,N_15919);
and U16976 (N_16976,N_15408,N_15597);
or U16977 (N_16977,N_15888,N_15870);
xnor U16978 (N_16978,N_15839,N_15741);
nand U16979 (N_16979,N_15975,N_15902);
and U16980 (N_16980,N_15168,N_15291);
nand U16981 (N_16981,N_15749,N_15045);
xor U16982 (N_16982,N_15249,N_15947);
nor U16983 (N_16983,N_15796,N_15975);
and U16984 (N_16984,N_15332,N_15084);
and U16985 (N_16985,N_15106,N_15170);
and U16986 (N_16986,N_15005,N_15363);
xor U16987 (N_16987,N_15144,N_15058);
xnor U16988 (N_16988,N_15638,N_15278);
xor U16989 (N_16989,N_15776,N_15801);
nor U16990 (N_16990,N_15781,N_15925);
xnor U16991 (N_16991,N_15835,N_15890);
nand U16992 (N_16992,N_15411,N_15570);
and U16993 (N_16993,N_15775,N_15986);
nand U16994 (N_16994,N_15519,N_15080);
and U16995 (N_16995,N_15594,N_15351);
or U16996 (N_16996,N_15366,N_15196);
nand U16997 (N_16997,N_15389,N_15258);
nand U16998 (N_16998,N_15769,N_15554);
or U16999 (N_16999,N_15488,N_15439);
nand U17000 (N_17000,N_16712,N_16702);
nand U17001 (N_17001,N_16398,N_16346);
nand U17002 (N_17002,N_16030,N_16805);
nor U17003 (N_17003,N_16669,N_16885);
and U17004 (N_17004,N_16825,N_16864);
and U17005 (N_17005,N_16911,N_16692);
nand U17006 (N_17006,N_16948,N_16925);
nand U17007 (N_17007,N_16716,N_16802);
xnor U17008 (N_17008,N_16848,N_16116);
nor U17009 (N_17009,N_16473,N_16021);
or U17010 (N_17010,N_16152,N_16184);
or U17011 (N_17011,N_16672,N_16454);
or U17012 (N_17012,N_16219,N_16409);
or U17013 (N_17013,N_16813,N_16552);
xnor U17014 (N_17014,N_16907,N_16946);
xor U17015 (N_17015,N_16936,N_16545);
or U17016 (N_17016,N_16789,N_16289);
or U17017 (N_17017,N_16452,N_16149);
or U17018 (N_17018,N_16131,N_16018);
nor U17019 (N_17019,N_16102,N_16889);
and U17020 (N_17020,N_16227,N_16698);
or U17021 (N_17021,N_16497,N_16902);
and U17022 (N_17022,N_16017,N_16480);
nor U17023 (N_17023,N_16175,N_16894);
nor U17024 (N_17024,N_16621,N_16042);
xor U17025 (N_17025,N_16496,N_16929);
nor U17026 (N_17026,N_16126,N_16031);
xor U17027 (N_17027,N_16979,N_16281);
nor U17028 (N_17028,N_16533,N_16819);
xor U17029 (N_17029,N_16954,N_16118);
xnor U17030 (N_17030,N_16080,N_16396);
xor U17031 (N_17031,N_16790,N_16650);
nand U17032 (N_17032,N_16603,N_16020);
nor U17033 (N_17033,N_16721,N_16294);
nand U17034 (N_17034,N_16982,N_16345);
nor U17035 (N_17035,N_16958,N_16176);
and U17036 (N_17036,N_16488,N_16104);
nor U17037 (N_17037,N_16292,N_16786);
nor U17038 (N_17038,N_16360,N_16604);
or U17039 (N_17039,N_16170,N_16707);
nand U17040 (N_17040,N_16174,N_16996);
or U17041 (N_17041,N_16185,N_16036);
or U17042 (N_17042,N_16154,N_16522);
nor U17043 (N_17043,N_16583,N_16440);
xnor U17044 (N_17044,N_16781,N_16691);
and U17045 (N_17045,N_16158,N_16964);
xnor U17046 (N_17046,N_16638,N_16852);
xnor U17047 (N_17047,N_16298,N_16746);
and U17048 (N_17048,N_16895,N_16617);
or U17049 (N_17049,N_16771,N_16661);
or U17050 (N_17050,N_16041,N_16785);
xnor U17051 (N_17051,N_16254,N_16849);
and U17052 (N_17052,N_16088,N_16594);
nor U17053 (N_17053,N_16363,N_16323);
nand U17054 (N_17054,N_16508,N_16228);
or U17055 (N_17055,N_16914,N_16288);
nand U17056 (N_17056,N_16013,N_16211);
nor U17057 (N_17057,N_16375,N_16690);
and U17058 (N_17058,N_16348,N_16788);
nand U17059 (N_17059,N_16266,N_16335);
nor U17060 (N_17060,N_16034,N_16942);
xor U17061 (N_17061,N_16535,N_16309);
or U17062 (N_17062,N_16483,N_16207);
and U17063 (N_17063,N_16893,N_16420);
nor U17064 (N_17064,N_16119,N_16862);
nor U17065 (N_17065,N_16833,N_16379);
xor U17066 (N_17066,N_16924,N_16319);
and U17067 (N_17067,N_16386,N_16588);
and U17068 (N_17068,N_16045,N_16332);
and U17069 (N_17069,N_16528,N_16025);
xnor U17070 (N_17070,N_16090,N_16960);
or U17071 (N_17071,N_16740,N_16479);
xor U17072 (N_17072,N_16901,N_16312);
and U17073 (N_17073,N_16441,N_16472);
or U17074 (N_17074,N_16608,N_16793);
nand U17075 (N_17075,N_16730,N_16250);
nand U17076 (N_17076,N_16340,N_16900);
nor U17077 (N_17077,N_16973,N_16745);
xor U17078 (N_17078,N_16518,N_16731);
or U17079 (N_17079,N_16359,N_16869);
nor U17080 (N_17080,N_16205,N_16708);
or U17081 (N_17081,N_16331,N_16634);
nor U17082 (N_17082,N_16172,N_16334);
or U17083 (N_17083,N_16941,N_16394);
xor U17084 (N_17084,N_16823,N_16799);
xor U17085 (N_17085,N_16418,N_16201);
nand U17086 (N_17086,N_16387,N_16007);
and U17087 (N_17087,N_16437,N_16354);
nand U17088 (N_17088,N_16632,N_16792);
nand U17089 (N_17089,N_16426,N_16320);
nor U17090 (N_17090,N_16027,N_16444);
xnor U17091 (N_17091,N_16548,N_16274);
or U17092 (N_17092,N_16024,N_16053);
or U17093 (N_17093,N_16477,N_16878);
nand U17094 (N_17094,N_16882,N_16992);
xnor U17095 (N_17095,N_16871,N_16815);
or U17096 (N_17096,N_16517,N_16407);
and U17097 (N_17097,N_16606,N_16693);
xor U17098 (N_17098,N_16618,N_16405);
and U17099 (N_17099,N_16747,N_16238);
or U17100 (N_17100,N_16188,N_16253);
nor U17101 (N_17101,N_16558,N_16866);
or U17102 (N_17102,N_16100,N_16766);
nor U17103 (N_17103,N_16435,N_16549);
nand U17104 (N_17104,N_16775,N_16416);
nand U17105 (N_17105,N_16757,N_16984);
or U17106 (N_17106,N_16905,N_16797);
or U17107 (N_17107,N_16678,N_16612);
nor U17108 (N_17108,N_16610,N_16989);
xor U17109 (N_17109,N_16986,N_16128);
xor U17110 (N_17110,N_16141,N_16314);
and U17111 (N_17111,N_16808,N_16389);
nor U17112 (N_17112,N_16482,N_16891);
or U17113 (N_17113,N_16400,N_16352);
or U17114 (N_17114,N_16972,N_16003);
and U17115 (N_17115,N_16168,N_16645);
or U17116 (N_17116,N_16868,N_16273);
nor U17117 (N_17117,N_16532,N_16539);
xnor U17118 (N_17118,N_16191,N_16845);
nor U17119 (N_17119,N_16713,N_16888);
xnor U17120 (N_17120,N_16991,N_16153);
nand U17121 (N_17121,N_16530,N_16863);
or U17122 (N_17122,N_16657,N_16415);
or U17123 (N_17123,N_16047,N_16167);
or U17124 (N_17124,N_16806,N_16462);
nor U17125 (N_17125,N_16967,N_16308);
xnor U17126 (N_17126,N_16990,N_16248);
nand U17127 (N_17127,N_16008,N_16046);
xnor U17128 (N_17128,N_16724,N_16132);
and U17129 (N_17129,N_16262,N_16777);
and U17130 (N_17130,N_16146,N_16755);
xnor U17131 (N_17131,N_16822,N_16401);
and U17132 (N_17132,N_16738,N_16589);
nand U17133 (N_17133,N_16322,N_16043);
and U17134 (N_17134,N_16801,N_16255);
or U17135 (N_17135,N_16404,N_16505);
nor U17136 (N_17136,N_16240,N_16210);
and U17137 (N_17137,N_16811,N_16576);
nor U17138 (N_17138,N_16920,N_16422);
nand U17139 (N_17139,N_16198,N_16486);
nand U17140 (N_17140,N_16023,N_16040);
or U17141 (N_17141,N_16867,N_16824);
nor U17142 (N_17142,N_16160,N_16770);
and U17143 (N_17143,N_16209,N_16872);
nor U17144 (N_17144,N_16303,N_16706);
and U17145 (N_17145,N_16668,N_16679);
nand U17146 (N_17146,N_16727,N_16392);
and U17147 (N_17147,N_16892,N_16005);
nand U17148 (N_17148,N_16851,N_16243);
nand U17149 (N_17149,N_16417,N_16778);
nand U17150 (N_17150,N_16935,N_16428);
nand U17151 (N_17151,N_16427,N_16385);
nand U17152 (N_17152,N_16546,N_16192);
nand U17153 (N_17153,N_16101,N_16110);
nand U17154 (N_17154,N_16840,N_16573);
nand U17155 (N_17155,N_16926,N_16699);
xnor U17156 (N_17156,N_16190,N_16411);
and U17157 (N_17157,N_16676,N_16049);
and U17158 (N_17158,N_16212,N_16962);
nand U17159 (N_17159,N_16330,N_16291);
nor U17160 (N_17160,N_16764,N_16710);
xor U17161 (N_17161,N_16999,N_16839);
and U17162 (N_17162,N_16874,N_16602);
or U17163 (N_17163,N_16685,N_16780);
xor U17164 (N_17164,N_16074,N_16510);
xor U17165 (N_17165,N_16696,N_16834);
or U17166 (N_17166,N_16665,N_16082);
xnor U17167 (N_17167,N_16615,N_16803);
xor U17168 (N_17168,N_16313,N_16299);
nor U17169 (N_17169,N_16562,N_16767);
and U17170 (N_17170,N_16062,N_16903);
nand U17171 (N_17171,N_16906,N_16841);
xor U17172 (N_17172,N_16897,N_16137);
or U17173 (N_17173,N_16876,N_16246);
or U17174 (N_17174,N_16861,N_16555);
xnor U17175 (N_17175,N_16870,N_16037);
xor U17176 (N_17176,N_16856,N_16376);
xnor U17177 (N_17177,N_16647,N_16233);
nand U17178 (N_17178,N_16351,N_16732);
nor U17179 (N_17179,N_16952,N_16358);
xor U17180 (N_17180,N_16121,N_16382);
nand U17181 (N_17181,N_16913,N_16859);
nor U17182 (N_17182,N_16270,N_16961);
or U17183 (N_17183,N_16560,N_16709);
nand U17184 (N_17184,N_16195,N_16344);
or U17185 (N_17185,N_16620,N_16827);
and U17186 (N_17186,N_16093,N_16529);
or U17187 (N_17187,N_16231,N_16112);
nand U17188 (N_17188,N_16403,N_16177);
or U17189 (N_17189,N_16078,N_16570);
and U17190 (N_17190,N_16216,N_16758);
and U17191 (N_17191,N_16994,N_16582);
or U17192 (N_17192,N_16276,N_16968);
and U17193 (N_17193,N_16613,N_16879);
xnor U17194 (N_17194,N_16217,N_16066);
nor U17195 (N_17195,N_16927,N_16258);
and U17196 (N_17196,N_16932,N_16912);
and U17197 (N_17197,N_16736,N_16247);
xor U17198 (N_17198,N_16094,N_16467);
xnor U17199 (N_17199,N_16026,N_16846);
nand U17200 (N_17200,N_16221,N_16064);
nor U17201 (N_17201,N_16663,N_16371);
xor U17202 (N_17202,N_16577,N_16259);
xnor U17203 (N_17203,N_16103,N_16627);
xor U17204 (N_17204,N_16855,N_16578);
or U17205 (N_17205,N_16140,N_16616);
nand U17206 (N_17206,N_16596,N_16585);
xnor U17207 (N_17207,N_16593,N_16381);
xnor U17208 (N_17208,N_16832,N_16910);
nor U17209 (N_17209,N_16318,N_16493);
or U17210 (N_17210,N_16329,N_16656);
and U17211 (N_17211,N_16640,N_16949);
nand U17212 (N_17212,N_16630,N_16760);
nor U17213 (N_17213,N_16224,N_16350);
and U17214 (N_17214,N_16223,N_16290);
and U17215 (N_17215,N_16068,N_16114);
nand U17216 (N_17216,N_16215,N_16772);
nand U17217 (N_17217,N_16988,N_16884);
nor U17218 (N_17218,N_16490,N_16938);
nand U17219 (N_17219,N_16711,N_16249);
nand U17220 (N_17220,N_16883,N_16611);
nand U17221 (N_17221,N_16957,N_16470);
xnor U17222 (N_17222,N_16099,N_16844);
nand U17223 (N_17223,N_16085,N_16842);
xor U17224 (N_17224,N_16092,N_16279);
nor U17225 (N_17225,N_16791,N_16537);
xor U17226 (N_17226,N_16642,N_16471);
nor U17227 (N_17227,N_16423,N_16006);
xor U17228 (N_17228,N_16644,N_16333);
and U17229 (N_17229,N_16012,N_16197);
xor U17230 (N_17230,N_16723,N_16076);
nor U17231 (N_17231,N_16511,N_16349);
or U17232 (N_17232,N_16985,N_16795);
xnor U17233 (N_17233,N_16139,N_16326);
nand U17234 (N_17234,N_16993,N_16130);
or U17235 (N_17235,N_16714,N_16787);
or U17236 (N_17236,N_16762,N_16408);
or U17237 (N_17237,N_16214,N_16944);
nor U17238 (N_17238,N_16821,N_16460);
nand U17239 (N_17239,N_16425,N_16365);
and U17240 (N_17240,N_16701,N_16705);
nor U17241 (N_17241,N_16674,N_16029);
or U17242 (N_17242,N_16830,N_16590);
or U17243 (N_17243,N_16783,N_16854);
or U17244 (N_17244,N_16521,N_16495);
nor U17245 (N_17245,N_16252,N_16660);
and U17246 (N_17246,N_16442,N_16180);
and U17247 (N_17247,N_16225,N_16111);
nor U17248 (N_17248,N_16481,N_16337);
xnor U17249 (N_17249,N_16150,N_16166);
nand U17250 (N_17250,N_16636,N_16512);
xnor U17251 (N_17251,N_16304,N_16461);
and U17252 (N_17252,N_16836,N_16937);
and U17253 (N_17253,N_16818,N_16000);
nor U17254 (N_17254,N_16828,N_16151);
and U17255 (N_17255,N_16817,N_16028);
xor U17256 (N_17256,N_16492,N_16305);
nor U17257 (N_17257,N_16487,N_16591);
or U17258 (N_17258,N_16814,N_16402);
xnor U17259 (N_17259,N_16413,N_16380);
or U17260 (N_17260,N_16761,N_16853);
nand U17261 (N_17261,N_16494,N_16523);
nor U17262 (N_17262,N_16136,N_16619);
xor U17263 (N_17263,N_16446,N_16081);
xor U17264 (N_17264,N_16873,N_16953);
nand U17265 (N_17265,N_16296,N_16666);
nor U17266 (N_17266,N_16516,N_16751);
or U17267 (N_17267,N_16229,N_16527);
nand U17268 (N_17268,N_16096,N_16744);
nand U17269 (N_17269,N_16526,N_16235);
and U17270 (N_17270,N_16011,N_16652);
and U17271 (N_17271,N_16919,N_16624);
and U17272 (N_17272,N_16673,N_16586);
nand U17273 (N_17273,N_16129,N_16436);
nand U17274 (N_17274,N_16956,N_16916);
xnor U17275 (N_17275,N_16917,N_16476);
or U17276 (N_17276,N_16393,N_16079);
xnor U17277 (N_17277,N_16733,N_16743);
xnor U17278 (N_17278,N_16779,N_16858);
or U17279 (N_17279,N_16930,N_16980);
nor U17280 (N_17280,N_16391,N_16133);
or U17281 (N_17281,N_16875,N_16559);
or U17282 (N_17282,N_16475,N_16609);
xor U17283 (N_17283,N_16316,N_16366);
nor U17284 (N_17284,N_16580,N_16317);
and U17285 (N_17285,N_16083,N_16943);
or U17286 (N_17286,N_16325,N_16507);
and U17287 (N_17287,N_16186,N_16816);
nor U17288 (N_17288,N_16628,N_16361);
xor U17289 (N_17289,N_16922,N_16084);
and U17290 (N_17290,N_16966,N_16173);
nand U17291 (N_17291,N_16509,N_16412);
nor U17292 (N_17292,N_16383,N_16269);
nor U17293 (N_17293,N_16646,N_16265);
xnor U17294 (N_17294,N_16001,N_16543);
nand U17295 (N_17295,N_16904,N_16339);
nor U17296 (N_17296,N_16500,N_16315);
nand U17297 (N_17297,N_16430,N_16453);
nand U17298 (N_17298,N_16032,N_16338);
xnor U17299 (N_17299,N_16498,N_16410);
xor U17300 (N_17300,N_16321,N_16059);
or U17301 (N_17301,N_16568,N_16311);
nor U17302 (N_17302,N_16502,N_16551);
xnor U17303 (N_17303,N_16057,N_16245);
xnor U17304 (N_17304,N_16242,N_16659);
or U17305 (N_17305,N_16282,N_16419);
or U17306 (N_17306,N_16055,N_16581);
xor U17307 (N_17307,N_16033,N_16695);
nor U17308 (N_17308,N_16633,N_16239);
or U17309 (N_17309,N_16302,N_16896);
and U17310 (N_17310,N_16039,N_16504);
nand U17311 (N_17311,N_16651,N_16561);
or U17312 (N_17312,N_16199,N_16147);
xnor U17313 (N_17313,N_16183,N_16458);
or U17314 (N_17314,N_16089,N_16687);
and U17315 (N_17315,N_16353,N_16865);
and U17316 (N_17316,N_16052,N_16019);
xnor U17317 (N_17317,N_16835,N_16970);
or U17318 (N_17318,N_16002,N_16782);
and U17319 (N_17319,N_16162,N_16800);
nor U17320 (N_17320,N_16424,N_16809);
nor U17321 (N_17321,N_16063,N_16843);
and U17322 (N_17322,N_16449,N_16431);
xnor U17323 (N_17323,N_16432,N_16260);
nand U17324 (N_17324,N_16058,N_16134);
or U17325 (N_17325,N_16915,N_16478);
xor U17326 (N_17326,N_16978,N_16038);
nor U17327 (N_17327,N_16256,N_16571);
nand U17328 (N_17328,N_16234,N_16484);
and U17329 (N_17329,N_16748,N_16395);
or U17330 (N_17330,N_16120,N_16213);
nor U17331 (N_17331,N_16165,N_16794);
nor U17332 (N_17332,N_16127,N_16820);
nor U17333 (N_17333,N_16564,N_16566);
nand U17334 (N_17334,N_16623,N_16754);
xor U17335 (N_17335,N_16688,N_16272);
nor U17336 (N_17336,N_16737,N_16369);
nor U17337 (N_17337,N_16998,N_16065);
nand U17338 (N_17338,N_16784,N_16356);
nand U17339 (N_17339,N_16513,N_16157);
or U17340 (N_17340,N_16464,N_16390);
xnor U17341 (N_17341,N_16880,N_16466);
nand U17342 (N_17342,N_16694,N_16536);
nor U17343 (N_17343,N_16686,N_16734);
xnor U17344 (N_17344,N_16362,N_16069);
nor U17345 (N_17345,N_16718,N_16887);
nor U17346 (N_17346,N_16655,N_16286);
xor U17347 (N_17347,N_16554,N_16977);
xor U17348 (N_17348,N_16773,N_16715);
xor U17349 (N_17349,N_16940,N_16631);
nand U17350 (N_17350,N_16307,N_16343);
nor U17351 (N_17351,N_16206,N_16164);
and U17352 (N_17352,N_16807,N_16251);
nor U17353 (N_17353,N_16899,N_16776);
nand U17354 (N_17354,N_16355,N_16014);
nand U17355 (N_17355,N_16287,N_16107);
xnor U17356 (N_17356,N_16067,N_16468);
nand U17357 (N_17357,N_16341,N_16155);
and U17358 (N_17358,N_16626,N_16531);
nand U17359 (N_17359,N_16939,N_16774);
and U17360 (N_17360,N_16503,N_16293);
nor U17361 (N_17361,N_16399,N_16414);
nand U17362 (N_17362,N_16009,N_16677);
and U17363 (N_17363,N_16056,N_16277);
or U17364 (N_17364,N_16682,N_16268);
nor U17365 (N_17365,N_16347,N_16796);
xor U17366 (N_17366,N_16098,N_16550);
nand U17367 (N_17367,N_16684,N_16106);
and U17368 (N_17368,N_16756,N_16831);
and U17369 (N_17369,N_16742,N_16637);
nand U17370 (N_17370,N_16667,N_16075);
nor U17371 (N_17371,N_16923,N_16597);
and U17372 (N_17372,N_16689,N_16283);
nand U17373 (N_17373,N_16997,N_16144);
xor U17374 (N_17374,N_16443,N_16670);
nand U17375 (N_17375,N_16324,N_16534);
xor U17376 (N_17376,N_16342,N_16377);
or U17377 (N_17377,N_16501,N_16675);
or U17378 (N_17378,N_16931,N_16161);
nand U17379 (N_17379,N_16995,N_16004);
nand U17380 (N_17380,N_16886,N_16951);
and U17381 (N_17381,N_16148,N_16450);
and U17382 (N_17382,N_16373,N_16171);
nand U17383 (N_17383,N_16087,N_16544);
and U17384 (N_17384,N_16438,N_16071);
xor U17385 (N_17385,N_16016,N_16236);
xnor U17386 (N_17386,N_16232,N_16918);
or U17387 (N_17387,N_16048,N_16050);
xnor U17388 (N_17388,N_16122,N_16538);
nor U17389 (N_17389,N_16241,N_16421);
and U17390 (N_17390,N_16921,N_16575);
or U17391 (N_17391,N_16541,N_16086);
and U17392 (N_17392,N_16397,N_16035);
nor U17393 (N_17393,N_16060,N_16750);
and U17394 (N_17394,N_16278,N_16187);
xor U17395 (N_17395,N_16680,N_16178);
xnor U17396 (N_17396,N_16542,N_16722);
nand U17397 (N_17397,N_16182,N_16285);
or U17398 (N_17398,N_16336,N_16181);
or U17399 (N_17399,N_16599,N_16226);
nand U17400 (N_17400,N_16725,N_16681);
nor U17401 (N_17401,N_16653,N_16662);
xor U17402 (N_17402,N_16847,N_16607);
nor U17403 (N_17403,N_16515,N_16955);
xnor U17404 (N_17404,N_16614,N_16565);
xnor U17405 (N_17405,N_16704,N_16933);
or U17406 (N_17406,N_16525,N_16169);
or U17407 (N_17407,N_16456,N_16969);
nor U17408 (N_17408,N_16189,N_16357);
nand U17409 (N_17409,N_16963,N_16113);
and U17410 (N_17410,N_16829,N_16553);
nand U17411 (N_17411,N_16697,N_16569);
or U17412 (N_17412,N_16156,N_16664);
nand U17413 (N_17413,N_16928,N_16474);
nand U17414 (N_17414,N_16439,N_16135);
nor U17415 (N_17415,N_16095,N_16881);
nor U17416 (N_17416,N_16584,N_16179);
and U17417 (N_17417,N_16301,N_16908);
xor U17418 (N_17418,N_16204,N_16196);
nor U17419 (N_17419,N_16200,N_16649);
nand U17420 (N_17420,N_16010,N_16890);
and U17421 (N_17421,N_16448,N_16328);
xnor U17422 (N_17422,N_16909,N_16244);
or U17423 (N_17423,N_16044,N_16054);
or U17424 (N_17424,N_16752,N_16465);
and U17425 (N_17425,N_16202,N_16367);
xnor U17426 (N_17426,N_16451,N_16729);
nand U17427 (N_17427,N_16193,N_16975);
xor U17428 (N_17428,N_16370,N_16717);
xor U17429 (N_17429,N_16768,N_16194);
nand U17430 (N_17430,N_16384,N_16798);
nand U17431 (N_17431,N_16388,N_16284);
or U17432 (N_17432,N_16739,N_16124);
xor U17433 (N_17433,N_16264,N_16295);
and U17434 (N_17434,N_16327,N_16429);
nor U17435 (N_17435,N_16759,N_16519);
nand U17436 (N_17436,N_16947,N_16574);
xnor U17437 (N_17437,N_16579,N_16683);
and U17438 (N_17438,N_16257,N_16524);
and U17439 (N_17439,N_16275,N_16514);
nor U17440 (N_17440,N_16983,N_16860);
xnor U17441 (N_17441,N_16115,N_16300);
or U17442 (N_17442,N_16749,N_16520);
and U17443 (N_17443,N_16719,N_16850);
nor U17444 (N_17444,N_16267,N_16364);
or U17445 (N_17445,N_16105,N_16601);
xnor U17446 (N_17446,N_16837,N_16965);
nand U17447 (N_17447,N_16051,N_16445);
and U17448 (N_17448,N_16648,N_16022);
nand U17449 (N_17449,N_16297,N_16109);
nor U17450 (N_17450,N_16457,N_16263);
or U17451 (N_17451,N_16838,N_16741);
nor U17452 (N_17452,N_16810,N_16898);
and U17453 (N_17453,N_16703,N_16671);
nand U17454 (N_17454,N_16222,N_16804);
nand U17455 (N_17455,N_16812,N_16143);
and U17456 (N_17456,N_16455,N_16629);
or U17457 (N_17457,N_16959,N_16540);
xnor U17458 (N_17458,N_16077,N_16230);
nor U17459 (N_17459,N_16433,N_16974);
nor U17460 (N_17460,N_16271,N_16163);
and U17461 (N_17461,N_16598,N_16987);
xor U17462 (N_17462,N_16261,N_16097);
xnor U17463 (N_17463,N_16635,N_16489);
and U17464 (N_17464,N_16981,N_16203);
or U17465 (N_17465,N_16567,N_16015);
and U17466 (N_17466,N_16070,N_16138);
or U17467 (N_17467,N_16123,N_16857);
nand U17468 (N_17468,N_16218,N_16108);
nor U17469 (N_17469,N_16459,N_16447);
xnor U17470 (N_17470,N_16061,N_16769);
and U17471 (N_17471,N_16826,N_16639);
nor U17472 (N_17472,N_16976,N_16547);
and U17473 (N_17473,N_16280,N_16072);
and U17474 (N_17474,N_16592,N_16726);
or U17475 (N_17475,N_16735,N_16654);
or U17476 (N_17476,N_16658,N_16753);
nor U17477 (N_17477,N_16117,N_16208);
or U17478 (N_17478,N_16145,N_16434);
xnor U17479 (N_17479,N_16310,N_16763);
xnor U17480 (N_17480,N_16159,N_16643);
or U17481 (N_17481,N_16374,N_16934);
nand U17482 (N_17482,N_16728,N_16971);
xnor U17483 (N_17483,N_16622,N_16378);
and U17484 (N_17484,N_16945,N_16469);
xnor U17485 (N_17485,N_16125,N_16950);
and U17486 (N_17486,N_16368,N_16572);
nor U17487 (N_17487,N_16499,N_16625);
or U17488 (N_17488,N_16306,N_16720);
or U17489 (N_17489,N_16142,N_16877);
or U17490 (N_17490,N_16220,N_16406);
and U17491 (N_17491,N_16485,N_16765);
and U17492 (N_17492,N_16563,N_16491);
nand U17493 (N_17493,N_16600,N_16463);
nand U17494 (N_17494,N_16237,N_16587);
and U17495 (N_17495,N_16595,N_16700);
nand U17496 (N_17496,N_16641,N_16556);
xor U17497 (N_17497,N_16605,N_16073);
nand U17498 (N_17498,N_16372,N_16091);
or U17499 (N_17499,N_16506,N_16557);
nand U17500 (N_17500,N_16686,N_16674);
xor U17501 (N_17501,N_16429,N_16110);
or U17502 (N_17502,N_16662,N_16929);
or U17503 (N_17503,N_16324,N_16720);
or U17504 (N_17504,N_16988,N_16114);
xnor U17505 (N_17505,N_16548,N_16137);
xor U17506 (N_17506,N_16685,N_16530);
or U17507 (N_17507,N_16897,N_16596);
or U17508 (N_17508,N_16618,N_16217);
nor U17509 (N_17509,N_16207,N_16240);
nand U17510 (N_17510,N_16073,N_16032);
nor U17511 (N_17511,N_16318,N_16997);
and U17512 (N_17512,N_16071,N_16307);
and U17513 (N_17513,N_16556,N_16011);
xnor U17514 (N_17514,N_16395,N_16701);
or U17515 (N_17515,N_16796,N_16842);
nor U17516 (N_17516,N_16376,N_16755);
xnor U17517 (N_17517,N_16330,N_16324);
nor U17518 (N_17518,N_16038,N_16792);
xnor U17519 (N_17519,N_16927,N_16126);
or U17520 (N_17520,N_16860,N_16533);
xnor U17521 (N_17521,N_16949,N_16931);
nand U17522 (N_17522,N_16524,N_16326);
nor U17523 (N_17523,N_16286,N_16784);
xor U17524 (N_17524,N_16502,N_16343);
or U17525 (N_17525,N_16192,N_16388);
xor U17526 (N_17526,N_16442,N_16518);
and U17527 (N_17527,N_16274,N_16481);
xor U17528 (N_17528,N_16161,N_16489);
xor U17529 (N_17529,N_16123,N_16890);
and U17530 (N_17530,N_16032,N_16743);
xnor U17531 (N_17531,N_16451,N_16340);
or U17532 (N_17532,N_16248,N_16630);
nand U17533 (N_17533,N_16551,N_16022);
and U17534 (N_17534,N_16084,N_16022);
xnor U17535 (N_17535,N_16834,N_16400);
and U17536 (N_17536,N_16171,N_16071);
nand U17537 (N_17537,N_16741,N_16817);
nand U17538 (N_17538,N_16937,N_16397);
or U17539 (N_17539,N_16400,N_16117);
nor U17540 (N_17540,N_16048,N_16019);
nand U17541 (N_17541,N_16341,N_16405);
and U17542 (N_17542,N_16060,N_16762);
nand U17543 (N_17543,N_16069,N_16328);
xor U17544 (N_17544,N_16398,N_16363);
and U17545 (N_17545,N_16012,N_16552);
nor U17546 (N_17546,N_16597,N_16683);
xor U17547 (N_17547,N_16917,N_16811);
xor U17548 (N_17548,N_16601,N_16677);
nor U17549 (N_17549,N_16777,N_16407);
nor U17550 (N_17550,N_16716,N_16382);
and U17551 (N_17551,N_16411,N_16700);
xnor U17552 (N_17552,N_16606,N_16558);
and U17553 (N_17553,N_16052,N_16693);
xnor U17554 (N_17554,N_16012,N_16557);
nand U17555 (N_17555,N_16977,N_16622);
or U17556 (N_17556,N_16116,N_16820);
nand U17557 (N_17557,N_16938,N_16441);
nor U17558 (N_17558,N_16675,N_16607);
xnor U17559 (N_17559,N_16728,N_16950);
and U17560 (N_17560,N_16635,N_16743);
and U17561 (N_17561,N_16052,N_16184);
nand U17562 (N_17562,N_16680,N_16283);
xnor U17563 (N_17563,N_16889,N_16535);
and U17564 (N_17564,N_16968,N_16010);
xor U17565 (N_17565,N_16633,N_16207);
and U17566 (N_17566,N_16754,N_16376);
nand U17567 (N_17567,N_16898,N_16545);
or U17568 (N_17568,N_16724,N_16000);
and U17569 (N_17569,N_16285,N_16111);
or U17570 (N_17570,N_16317,N_16903);
xnor U17571 (N_17571,N_16629,N_16277);
nor U17572 (N_17572,N_16358,N_16455);
xnor U17573 (N_17573,N_16138,N_16763);
or U17574 (N_17574,N_16449,N_16806);
and U17575 (N_17575,N_16042,N_16182);
nand U17576 (N_17576,N_16601,N_16178);
nor U17577 (N_17577,N_16928,N_16857);
xor U17578 (N_17578,N_16681,N_16115);
nand U17579 (N_17579,N_16866,N_16940);
nor U17580 (N_17580,N_16175,N_16673);
nand U17581 (N_17581,N_16649,N_16809);
or U17582 (N_17582,N_16506,N_16712);
and U17583 (N_17583,N_16411,N_16376);
nand U17584 (N_17584,N_16709,N_16767);
or U17585 (N_17585,N_16215,N_16508);
and U17586 (N_17586,N_16698,N_16024);
nor U17587 (N_17587,N_16850,N_16527);
xor U17588 (N_17588,N_16182,N_16094);
xor U17589 (N_17589,N_16865,N_16310);
xor U17590 (N_17590,N_16111,N_16138);
xor U17591 (N_17591,N_16861,N_16892);
nor U17592 (N_17592,N_16225,N_16794);
or U17593 (N_17593,N_16652,N_16965);
nor U17594 (N_17594,N_16593,N_16713);
nand U17595 (N_17595,N_16007,N_16446);
nor U17596 (N_17596,N_16250,N_16130);
or U17597 (N_17597,N_16238,N_16276);
nor U17598 (N_17598,N_16770,N_16003);
xor U17599 (N_17599,N_16306,N_16679);
nor U17600 (N_17600,N_16219,N_16519);
nand U17601 (N_17601,N_16430,N_16556);
nand U17602 (N_17602,N_16097,N_16248);
nor U17603 (N_17603,N_16562,N_16678);
nand U17604 (N_17604,N_16115,N_16560);
and U17605 (N_17605,N_16763,N_16983);
and U17606 (N_17606,N_16626,N_16861);
and U17607 (N_17607,N_16861,N_16297);
nand U17608 (N_17608,N_16612,N_16352);
or U17609 (N_17609,N_16768,N_16138);
nand U17610 (N_17610,N_16040,N_16225);
nand U17611 (N_17611,N_16564,N_16350);
or U17612 (N_17612,N_16748,N_16048);
and U17613 (N_17613,N_16250,N_16986);
xnor U17614 (N_17614,N_16696,N_16333);
nand U17615 (N_17615,N_16714,N_16620);
or U17616 (N_17616,N_16815,N_16584);
or U17617 (N_17617,N_16556,N_16550);
and U17618 (N_17618,N_16808,N_16740);
nor U17619 (N_17619,N_16520,N_16446);
nand U17620 (N_17620,N_16031,N_16515);
xor U17621 (N_17621,N_16831,N_16466);
nand U17622 (N_17622,N_16899,N_16375);
and U17623 (N_17623,N_16835,N_16133);
and U17624 (N_17624,N_16564,N_16360);
and U17625 (N_17625,N_16686,N_16369);
nand U17626 (N_17626,N_16760,N_16066);
xor U17627 (N_17627,N_16791,N_16076);
and U17628 (N_17628,N_16671,N_16369);
xor U17629 (N_17629,N_16798,N_16093);
and U17630 (N_17630,N_16610,N_16892);
nand U17631 (N_17631,N_16017,N_16212);
and U17632 (N_17632,N_16352,N_16700);
nor U17633 (N_17633,N_16855,N_16996);
and U17634 (N_17634,N_16189,N_16578);
and U17635 (N_17635,N_16431,N_16996);
xnor U17636 (N_17636,N_16185,N_16497);
and U17637 (N_17637,N_16543,N_16856);
nor U17638 (N_17638,N_16855,N_16850);
nand U17639 (N_17639,N_16087,N_16747);
or U17640 (N_17640,N_16534,N_16826);
and U17641 (N_17641,N_16763,N_16490);
and U17642 (N_17642,N_16109,N_16153);
nand U17643 (N_17643,N_16086,N_16158);
and U17644 (N_17644,N_16129,N_16626);
nor U17645 (N_17645,N_16736,N_16818);
and U17646 (N_17646,N_16638,N_16510);
or U17647 (N_17647,N_16119,N_16548);
xnor U17648 (N_17648,N_16708,N_16622);
or U17649 (N_17649,N_16226,N_16061);
or U17650 (N_17650,N_16529,N_16495);
or U17651 (N_17651,N_16332,N_16004);
nor U17652 (N_17652,N_16311,N_16619);
xor U17653 (N_17653,N_16283,N_16552);
or U17654 (N_17654,N_16731,N_16369);
or U17655 (N_17655,N_16831,N_16626);
nand U17656 (N_17656,N_16633,N_16583);
or U17657 (N_17657,N_16660,N_16807);
nand U17658 (N_17658,N_16760,N_16756);
nor U17659 (N_17659,N_16565,N_16575);
nand U17660 (N_17660,N_16413,N_16186);
xnor U17661 (N_17661,N_16626,N_16657);
or U17662 (N_17662,N_16750,N_16359);
and U17663 (N_17663,N_16978,N_16246);
nor U17664 (N_17664,N_16687,N_16063);
and U17665 (N_17665,N_16692,N_16328);
nor U17666 (N_17666,N_16105,N_16933);
nand U17667 (N_17667,N_16816,N_16245);
xor U17668 (N_17668,N_16306,N_16406);
and U17669 (N_17669,N_16750,N_16826);
and U17670 (N_17670,N_16997,N_16808);
and U17671 (N_17671,N_16148,N_16947);
and U17672 (N_17672,N_16818,N_16352);
xor U17673 (N_17673,N_16483,N_16027);
or U17674 (N_17674,N_16936,N_16300);
xnor U17675 (N_17675,N_16065,N_16955);
nor U17676 (N_17676,N_16348,N_16298);
and U17677 (N_17677,N_16522,N_16901);
nand U17678 (N_17678,N_16982,N_16564);
xnor U17679 (N_17679,N_16143,N_16297);
xor U17680 (N_17680,N_16316,N_16206);
xnor U17681 (N_17681,N_16173,N_16454);
and U17682 (N_17682,N_16120,N_16655);
xnor U17683 (N_17683,N_16958,N_16720);
xnor U17684 (N_17684,N_16667,N_16741);
nand U17685 (N_17685,N_16745,N_16419);
or U17686 (N_17686,N_16144,N_16275);
nor U17687 (N_17687,N_16895,N_16462);
xor U17688 (N_17688,N_16113,N_16961);
or U17689 (N_17689,N_16635,N_16627);
nand U17690 (N_17690,N_16276,N_16571);
or U17691 (N_17691,N_16061,N_16200);
and U17692 (N_17692,N_16251,N_16953);
xnor U17693 (N_17693,N_16108,N_16163);
xnor U17694 (N_17694,N_16574,N_16660);
nor U17695 (N_17695,N_16007,N_16417);
and U17696 (N_17696,N_16673,N_16917);
nand U17697 (N_17697,N_16169,N_16457);
nor U17698 (N_17698,N_16723,N_16511);
or U17699 (N_17699,N_16587,N_16994);
xor U17700 (N_17700,N_16724,N_16685);
nand U17701 (N_17701,N_16188,N_16444);
nand U17702 (N_17702,N_16251,N_16234);
nor U17703 (N_17703,N_16630,N_16514);
nand U17704 (N_17704,N_16359,N_16482);
and U17705 (N_17705,N_16395,N_16000);
nand U17706 (N_17706,N_16996,N_16426);
and U17707 (N_17707,N_16891,N_16447);
nand U17708 (N_17708,N_16514,N_16310);
nor U17709 (N_17709,N_16237,N_16065);
xor U17710 (N_17710,N_16610,N_16459);
and U17711 (N_17711,N_16563,N_16240);
nand U17712 (N_17712,N_16329,N_16043);
nand U17713 (N_17713,N_16074,N_16529);
and U17714 (N_17714,N_16913,N_16648);
nand U17715 (N_17715,N_16540,N_16131);
or U17716 (N_17716,N_16338,N_16613);
nand U17717 (N_17717,N_16033,N_16612);
or U17718 (N_17718,N_16511,N_16359);
nor U17719 (N_17719,N_16428,N_16790);
xnor U17720 (N_17720,N_16777,N_16815);
xnor U17721 (N_17721,N_16456,N_16661);
nor U17722 (N_17722,N_16681,N_16655);
xor U17723 (N_17723,N_16585,N_16408);
and U17724 (N_17724,N_16541,N_16016);
and U17725 (N_17725,N_16624,N_16821);
nand U17726 (N_17726,N_16535,N_16462);
nor U17727 (N_17727,N_16202,N_16875);
nand U17728 (N_17728,N_16403,N_16539);
and U17729 (N_17729,N_16068,N_16560);
nand U17730 (N_17730,N_16373,N_16192);
xnor U17731 (N_17731,N_16560,N_16396);
and U17732 (N_17732,N_16008,N_16486);
xor U17733 (N_17733,N_16484,N_16700);
and U17734 (N_17734,N_16220,N_16504);
or U17735 (N_17735,N_16524,N_16312);
nand U17736 (N_17736,N_16935,N_16358);
and U17737 (N_17737,N_16455,N_16489);
or U17738 (N_17738,N_16131,N_16397);
xor U17739 (N_17739,N_16064,N_16238);
nor U17740 (N_17740,N_16022,N_16973);
nand U17741 (N_17741,N_16978,N_16984);
nand U17742 (N_17742,N_16293,N_16907);
or U17743 (N_17743,N_16623,N_16162);
and U17744 (N_17744,N_16244,N_16266);
and U17745 (N_17745,N_16463,N_16601);
or U17746 (N_17746,N_16359,N_16464);
or U17747 (N_17747,N_16295,N_16557);
or U17748 (N_17748,N_16546,N_16209);
nor U17749 (N_17749,N_16634,N_16315);
nor U17750 (N_17750,N_16118,N_16623);
nand U17751 (N_17751,N_16736,N_16847);
and U17752 (N_17752,N_16179,N_16359);
xor U17753 (N_17753,N_16542,N_16296);
nand U17754 (N_17754,N_16174,N_16177);
nor U17755 (N_17755,N_16845,N_16048);
nand U17756 (N_17756,N_16619,N_16350);
and U17757 (N_17757,N_16368,N_16740);
or U17758 (N_17758,N_16084,N_16551);
xor U17759 (N_17759,N_16085,N_16062);
or U17760 (N_17760,N_16610,N_16891);
nor U17761 (N_17761,N_16293,N_16249);
or U17762 (N_17762,N_16707,N_16130);
nand U17763 (N_17763,N_16289,N_16950);
or U17764 (N_17764,N_16557,N_16142);
nor U17765 (N_17765,N_16175,N_16378);
nand U17766 (N_17766,N_16969,N_16912);
nor U17767 (N_17767,N_16797,N_16662);
nand U17768 (N_17768,N_16985,N_16050);
and U17769 (N_17769,N_16513,N_16420);
or U17770 (N_17770,N_16298,N_16386);
and U17771 (N_17771,N_16161,N_16562);
nor U17772 (N_17772,N_16432,N_16401);
nor U17773 (N_17773,N_16728,N_16180);
xnor U17774 (N_17774,N_16746,N_16048);
xnor U17775 (N_17775,N_16820,N_16122);
and U17776 (N_17776,N_16444,N_16778);
nand U17777 (N_17777,N_16360,N_16809);
xor U17778 (N_17778,N_16099,N_16828);
and U17779 (N_17779,N_16528,N_16150);
or U17780 (N_17780,N_16450,N_16965);
xnor U17781 (N_17781,N_16653,N_16821);
nand U17782 (N_17782,N_16736,N_16832);
nor U17783 (N_17783,N_16749,N_16925);
or U17784 (N_17784,N_16784,N_16821);
nor U17785 (N_17785,N_16195,N_16127);
xnor U17786 (N_17786,N_16653,N_16473);
nand U17787 (N_17787,N_16428,N_16348);
and U17788 (N_17788,N_16506,N_16667);
nor U17789 (N_17789,N_16117,N_16249);
and U17790 (N_17790,N_16221,N_16890);
nand U17791 (N_17791,N_16900,N_16810);
and U17792 (N_17792,N_16530,N_16942);
or U17793 (N_17793,N_16990,N_16203);
nand U17794 (N_17794,N_16603,N_16928);
nand U17795 (N_17795,N_16942,N_16249);
xnor U17796 (N_17796,N_16417,N_16113);
xor U17797 (N_17797,N_16992,N_16244);
nor U17798 (N_17798,N_16277,N_16410);
nor U17799 (N_17799,N_16512,N_16239);
nor U17800 (N_17800,N_16349,N_16583);
nor U17801 (N_17801,N_16055,N_16290);
xnor U17802 (N_17802,N_16763,N_16974);
and U17803 (N_17803,N_16135,N_16987);
xnor U17804 (N_17804,N_16362,N_16067);
nand U17805 (N_17805,N_16880,N_16796);
and U17806 (N_17806,N_16004,N_16716);
nand U17807 (N_17807,N_16033,N_16799);
xor U17808 (N_17808,N_16836,N_16880);
nor U17809 (N_17809,N_16591,N_16675);
nor U17810 (N_17810,N_16227,N_16642);
xnor U17811 (N_17811,N_16171,N_16297);
xor U17812 (N_17812,N_16225,N_16585);
and U17813 (N_17813,N_16449,N_16627);
and U17814 (N_17814,N_16104,N_16017);
nand U17815 (N_17815,N_16066,N_16356);
xor U17816 (N_17816,N_16939,N_16254);
nor U17817 (N_17817,N_16127,N_16175);
xor U17818 (N_17818,N_16729,N_16707);
nand U17819 (N_17819,N_16993,N_16802);
or U17820 (N_17820,N_16637,N_16059);
nor U17821 (N_17821,N_16093,N_16582);
nor U17822 (N_17822,N_16596,N_16075);
nor U17823 (N_17823,N_16316,N_16523);
or U17824 (N_17824,N_16633,N_16417);
and U17825 (N_17825,N_16001,N_16010);
and U17826 (N_17826,N_16772,N_16673);
or U17827 (N_17827,N_16364,N_16944);
or U17828 (N_17828,N_16194,N_16885);
nand U17829 (N_17829,N_16555,N_16635);
and U17830 (N_17830,N_16031,N_16058);
and U17831 (N_17831,N_16435,N_16951);
and U17832 (N_17832,N_16447,N_16196);
xnor U17833 (N_17833,N_16664,N_16923);
or U17834 (N_17834,N_16098,N_16001);
xor U17835 (N_17835,N_16343,N_16229);
and U17836 (N_17836,N_16883,N_16856);
or U17837 (N_17837,N_16100,N_16450);
xor U17838 (N_17838,N_16355,N_16224);
or U17839 (N_17839,N_16806,N_16767);
nand U17840 (N_17840,N_16780,N_16250);
nand U17841 (N_17841,N_16481,N_16318);
xnor U17842 (N_17842,N_16606,N_16651);
nor U17843 (N_17843,N_16554,N_16559);
and U17844 (N_17844,N_16924,N_16461);
nand U17845 (N_17845,N_16292,N_16584);
nand U17846 (N_17846,N_16904,N_16189);
xnor U17847 (N_17847,N_16779,N_16093);
and U17848 (N_17848,N_16535,N_16315);
or U17849 (N_17849,N_16818,N_16577);
xor U17850 (N_17850,N_16738,N_16022);
nor U17851 (N_17851,N_16490,N_16400);
xor U17852 (N_17852,N_16548,N_16296);
xor U17853 (N_17853,N_16979,N_16483);
and U17854 (N_17854,N_16540,N_16002);
xnor U17855 (N_17855,N_16593,N_16015);
and U17856 (N_17856,N_16355,N_16697);
xor U17857 (N_17857,N_16805,N_16276);
xnor U17858 (N_17858,N_16024,N_16911);
and U17859 (N_17859,N_16486,N_16021);
nor U17860 (N_17860,N_16558,N_16529);
nand U17861 (N_17861,N_16214,N_16491);
and U17862 (N_17862,N_16935,N_16507);
nand U17863 (N_17863,N_16217,N_16834);
and U17864 (N_17864,N_16457,N_16437);
and U17865 (N_17865,N_16359,N_16954);
and U17866 (N_17866,N_16771,N_16593);
xor U17867 (N_17867,N_16740,N_16302);
or U17868 (N_17868,N_16216,N_16658);
nand U17869 (N_17869,N_16321,N_16290);
nor U17870 (N_17870,N_16990,N_16727);
nor U17871 (N_17871,N_16197,N_16298);
nand U17872 (N_17872,N_16094,N_16552);
or U17873 (N_17873,N_16336,N_16150);
and U17874 (N_17874,N_16581,N_16136);
nor U17875 (N_17875,N_16037,N_16217);
xor U17876 (N_17876,N_16548,N_16140);
or U17877 (N_17877,N_16482,N_16524);
and U17878 (N_17878,N_16892,N_16390);
nor U17879 (N_17879,N_16644,N_16009);
xnor U17880 (N_17880,N_16190,N_16405);
and U17881 (N_17881,N_16324,N_16208);
or U17882 (N_17882,N_16361,N_16705);
nor U17883 (N_17883,N_16282,N_16703);
nand U17884 (N_17884,N_16174,N_16765);
and U17885 (N_17885,N_16226,N_16532);
and U17886 (N_17886,N_16539,N_16725);
or U17887 (N_17887,N_16072,N_16449);
nor U17888 (N_17888,N_16087,N_16549);
nand U17889 (N_17889,N_16409,N_16137);
nand U17890 (N_17890,N_16310,N_16748);
nand U17891 (N_17891,N_16367,N_16374);
and U17892 (N_17892,N_16965,N_16429);
or U17893 (N_17893,N_16261,N_16086);
or U17894 (N_17894,N_16129,N_16855);
and U17895 (N_17895,N_16343,N_16862);
xnor U17896 (N_17896,N_16811,N_16135);
nand U17897 (N_17897,N_16779,N_16923);
nor U17898 (N_17898,N_16048,N_16579);
nand U17899 (N_17899,N_16825,N_16192);
nand U17900 (N_17900,N_16263,N_16230);
nor U17901 (N_17901,N_16207,N_16815);
or U17902 (N_17902,N_16782,N_16984);
or U17903 (N_17903,N_16164,N_16022);
xor U17904 (N_17904,N_16267,N_16429);
xnor U17905 (N_17905,N_16742,N_16443);
xnor U17906 (N_17906,N_16628,N_16407);
xor U17907 (N_17907,N_16421,N_16851);
nand U17908 (N_17908,N_16235,N_16875);
nand U17909 (N_17909,N_16985,N_16793);
and U17910 (N_17910,N_16361,N_16579);
xor U17911 (N_17911,N_16310,N_16118);
and U17912 (N_17912,N_16122,N_16472);
nor U17913 (N_17913,N_16326,N_16304);
or U17914 (N_17914,N_16883,N_16447);
or U17915 (N_17915,N_16600,N_16935);
and U17916 (N_17916,N_16617,N_16411);
nor U17917 (N_17917,N_16593,N_16183);
xor U17918 (N_17918,N_16107,N_16743);
or U17919 (N_17919,N_16397,N_16393);
and U17920 (N_17920,N_16742,N_16603);
nand U17921 (N_17921,N_16655,N_16975);
or U17922 (N_17922,N_16205,N_16255);
xor U17923 (N_17923,N_16993,N_16146);
nor U17924 (N_17924,N_16229,N_16437);
and U17925 (N_17925,N_16995,N_16459);
nand U17926 (N_17926,N_16888,N_16287);
or U17927 (N_17927,N_16735,N_16392);
or U17928 (N_17928,N_16435,N_16948);
xor U17929 (N_17929,N_16089,N_16881);
nor U17930 (N_17930,N_16661,N_16358);
or U17931 (N_17931,N_16452,N_16025);
nor U17932 (N_17932,N_16208,N_16445);
or U17933 (N_17933,N_16396,N_16028);
nor U17934 (N_17934,N_16566,N_16644);
nor U17935 (N_17935,N_16077,N_16833);
nand U17936 (N_17936,N_16411,N_16567);
nor U17937 (N_17937,N_16641,N_16447);
nor U17938 (N_17938,N_16535,N_16200);
xnor U17939 (N_17939,N_16243,N_16167);
and U17940 (N_17940,N_16245,N_16677);
nand U17941 (N_17941,N_16944,N_16735);
or U17942 (N_17942,N_16526,N_16902);
and U17943 (N_17943,N_16846,N_16804);
nor U17944 (N_17944,N_16204,N_16689);
nor U17945 (N_17945,N_16873,N_16242);
or U17946 (N_17946,N_16854,N_16430);
nand U17947 (N_17947,N_16903,N_16850);
nor U17948 (N_17948,N_16057,N_16075);
xor U17949 (N_17949,N_16738,N_16389);
xor U17950 (N_17950,N_16018,N_16765);
nor U17951 (N_17951,N_16960,N_16832);
nand U17952 (N_17952,N_16643,N_16420);
or U17953 (N_17953,N_16734,N_16070);
and U17954 (N_17954,N_16969,N_16197);
and U17955 (N_17955,N_16235,N_16595);
or U17956 (N_17956,N_16881,N_16278);
or U17957 (N_17957,N_16996,N_16952);
nor U17958 (N_17958,N_16173,N_16642);
xnor U17959 (N_17959,N_16746,N_16497);
or U17960 (N_17960,N_16672,N_16748);
nor U17961 (N_17961,N_16853,N_16586);
xor U17962 (N_17962,N_16665,N_16719);
or U17963 (N_17963,N_16927,N_16523);
xor U17964 (N_17964,N_16071,N_16454);
or U17965 (N_17965,N_16981,N_16828);
and U17966 (N_17966,N_16258,N_16263);
xnor U17967 (N_17967,N_16392,N_16662);
xnor U17968 (N_17968,N_16425,N_16375);
and U17969 (N_17969,N_16665,N_16611);
nor U17970 (N_17970,N_16338,N_16247);
xor U17971 (N_17971,N_16640,N_16619);
or U17972 (N_17972,N_16461,N_16634);
or U17973 (N_17973,N_16244,N_16357);
and U17974 (N_17974,N_16876,N_16956);
nand U17975 (N_17975,N_16647,N_16482);
xnor U17976 (N_17976,N_16926,N_16861);
and U17977 (N_17977,N_16036,N_16249);
or U17978 (N_17978,N_16499,N_16385);
or U17979 (N_17979,N_16291,N_16225);
and U17980 (N_17980,N_16281,N_16010);
nand U17981 (N_17981,N_16816,N_16132);
nor U17982 (N_17982,N_16694,N_16527);
nor U17983 (N_17983,N_16444,N_16475);
nand U17984 (N_17984,N_16660,N_16051);
and U17985 (N_17985,N_16987,N_16937);
or U17986 (N_17986,N_16583,N_16632);
xor U17987 (N_17987,N_16510,N_16365);
or U17988 (N_17988,N_16293,N_16581);
and U17989 (N_17989,N_16059,N_16946);
nand U17990 (N_17990,N_16128,N_16547);
or U17991 (N_17991,N_16763,N_16087);
nor U17992 (N_17992,N_16732,N_16287);
xnor U17993 (N_17993,N_16114,N_16808);
nand U17994 (N_17994,N_16237,N_16780);
and U17995 (N_17995,N_16613,N_16730);
nor U17996 (N_17996,N_16832,N_16766);
and U17997 (N_17997,N_16540,N_16887);
and U17998 (N_17998,N_16727,N_16286);
xnor U17999 (N_17999,N_16506,N_16538);
and U18000 (N_18000,N_17799,N_17696);
xor U18001 (N_18001,N_17409,N_17869);
or U18002 (N_18002,N_17722,N_17516);
xor U18003 (N_18003,N_17000,N_17442);
nand U18004 (N_18004,N_17660,N_17582);
nand U18005 (N_18005,N_17873,N_17498);
nor U18006 (N_18006,N_17657,N_17644);
nand U18007 (N_18007,N_17710,N_17019);
nand U18008 (N_18008,N_17370,N_17860);
nor U18009 (N_18009,N_17693,N_17268);
nor U18010 (N_18010,N_17899,N_17043);
and U18011 (N_18011,N_17047,N_17173);
or U18012 (N_18012,N_17745,N_17548);
xor U18013 (N_18013,N_17249,N_17880);
or U18014 (N_18014,N_17975,N_17196);
nor U18015 (N_18015,N_17870,N_17280);
nand U18016 (N_18016,N_17385,N_17754);
or U18017 (N_18017,N_17094,N_17484);
or U18018 (N_18018,N_17999,N_17113);
xnor U18019 (N_18019,N_17263,N_17414);
or U18020 (N_18020,N_17248,N_17459);
and U18021 (N_18021,N_17956,N_17401);
nand U18022 (N_18022,N_17957,N_17301);
nor U18023 (N_18023,N_17621,N_17685);
xnor U18024 (N_18024,N_17319,N_17384);
nand U18025 (N_18025,N_17001,N_17131);
nand U18026 (N_18026,N_17018,N_17061);
nand U18027 (N_18027,N_17768,N_17298);
xor U18028 (N_18028,N_17357,N_17228);
nand U18029 (N_18029,N_17328,N_17483);
xnor U18030 (N_18030,N_17290,N_17361);
and U18031 (N_18031,N_17240,N_17063);
xor U18032 (N_18032,N_17239,N_17890);
xnor U18033 (N_18033,N_17372,N_17488);
xnor U18034 (N_18034,N_17500,N_17591);
and U18035 (N_18035,N_17005,N_17129);
nand U18036 (N_18036,N_17503,N_17607);
and U18037 (N_18037,N_17731,N_17403);
or U18038 (N_18038,N_17450,N_17154);
xor U18039 (N_18039,N_17759,N_17358);
or U18040 (N_18040,N_17288,N_17990);
nor U18041 (N_18041,N_17225,N_17284);
nand U18042 (N_18042,N_17969,N_17387);
and U18043 (N_18043,N_17440,N_17623);
or U18044 (N_18044,N_17979,N_17354);
or U18045 (N_18045,N_17160,N_17663);
nor U18046 (N_18046,N_17415,N_17736);
and U18047 (N_18047,N_17097,N_17096);
and U18048 (N_18048,N_17692,N_17310);
and U18049 (N_18049,N_17645,N_17705);
and U18050 (N_18050,N_17261,N_17646);
or U18051 (N_18051,N_17785,N_17479);
nand U18052 (N_18052,N_17793,N_17186);
or U18053 (N_18053,N_17888,N_17057);
nor U18054 (N_18054,N_17404,N_17550);
or U18055 (N_18055,N_17824,N_17017);
nand U18056 (N_18056,N_17152,N_17830);
and U18057 (N_18057,N_17733,N_17523);
and U18058 (N_18058,N_17753,N_17464);
nor U18059 (N_18059,N_17070,N_17991);
nor U18060 (N_18060,N_17165,N_17469);
or U18061 (N_18061,N_17568,N_17948);
nor U18062 (N_18062,N_17105,N_17529);
and U18063 (N_18063,N_17453,N_17737);
and U18064 (N_18064,N_17117,N_17378);
nor U18065 (N_18065,N_17220,N_17161);
xor U18066 (N_18066,N_17671,N_17170);
xor U18067 (N_18067,N_17138,N_17968);
nor U18068 (N_18068,N_17713,N_17934);
or U18069 (N_18069,N_17149,N_17128);
nand U18070 (N_18070,N_17281,N_17262);
nor U18071 (N_18071,N_17087,N_17557);
xnor U18072 (N_18072,N_17997,N_17324);
nand U18073 (N_18073,N_17107,N_17474);
and U18074 (N_18074,N_17933,N_17289);
nand U18075 (N_18075,N_17555,N_17726);
or U18076 (N_18076,N_17583,N_17762);
or U18077 (N_18077,N_17576,N_17283);
nor U18078 (N_18078,N_17126,N_17527);
and U18079 (N_18079,N_17192,N_17156);
xor U18080 (N_18080,N_17536,N_17614);
nor U18081 (N_18081,N_17443,N_17652);
or U18082 (N_18082,N_17006,N_17701);
xor U18083 (N_18083,N_17981,N_17502);
and U18084 (N_18084,N_17028,N_17676);
and U18085 (N_18085,N_17862,N_17859);
nor U18086 (N_18086,N_17137,N_17677);
or U18087 (N_18087,N_17617,N_17511);
nand U18088 (N_18088,N_17509,N_17564);
and U18089 (N_18089,N_17963,N_17100);
nand U18090 (N_18090,N_17702,N_17856);
nor U18091 (N_18091,N_17279,N_17441);
and U18092 (N_18092,N_17510,N_17266);
nor U18093 (N_18093,N_17595,N_17925);
and U18094 (N_18094,N_17827,N_17837);
nor U18095 (N_18095,N_17917,N_17075);
or U18096 (N_18096,N_17081,N_17418);
xnor U18097 (N_18097,N_17789,N_17458);
and U18098 (N_18098,N_17430,N_17219);
or U18099 (N_18099,N_17541,N_17515);
and U18100 (N_18100,N_17364,N_17485);
and U18101 (N_18101,N_17210,N_17417);
and U18102 (N_18102,N_17039,N_17208);
xor U18103 (N_18103,N_17135,N_17727);
or U18104 (N_18104,N_17294,N_17130);
xor U18105 (N_18105,N_17055,N_17237);
nand U18106 (N_18106,N_17233,N_17913);
nor U18107 (N_18107,N_17487,N_17898);
xor U18108 (N_18108,N_17496,N_17601);
or U18109 (N_18109,N_17185,N_17891);
nor U18110 (N_18110,N_17588,N_17569);
nand U18111 (N_18111,N_17446,N_17127);
or U18112 (N_18112,N_17408,N_17034);
nand U18113 (N_18113,N_17932,N_17901);
and U18114 (N_18114,N_17912,N_17903);
nand U18115 (N_18115,N_17629,N_17444);
xnor U18116 (N_18116,N_17780,N_17172);
or U18117 (N_18117,N_17315,N_17313);
and U18118 (N_18118,N_17482,N_17486);
or U18119 (N_18119,N_17157,N_17463);
and U18120 (N_18120,N_17247,N_17504);
nor U18121 (N_18121,N_17435,N_17944);
or U18122 (N_18122,N_17774,N_17594);
nand U18123 (N_18123,N_17814,N_17544);
nand U18124 (N_18124,N_17764,N_17662);
and U18125 (N_18125,N_17893,N_17141);
nand U18126 (N_18126,N_17015,N_17460);
nand U18127 (N_18127,N_17300,N_17600);
or U18128 (N_18128,N_17392,N_17633);
nor U18129 (N_18129,N_17021,N_17335);
nand U18130 (N_18130,N_17982,N_17073);
xor U18131 (N_18131,N_17411,N_17635);
nor U18132 (N_18132,N_17563,N_17794);
and U18133 (N_18133,N_17570,N_17560);
xnor U18134 (N_18134,N_17610,N_17339);
and U18135 (N_18135,N_17145,N_17467);
xor U18136 (N_18136,N_17092,N_17033);
xnor U18137 (N_18137,N_17329,N_17807);
xnor U18138 (N_18138,N_17473,N_17059);
or U18139 (N_18139,N_17743,N_17101);
nand U18140 (N_18140,N_17347,N_17738);
nor U18141 (N_18141,N_17489,N_17532);
nand U18142 (N_18142,N_17278,N_17760);
nor U18143 (N_18143,N_17350,N_17391);
nand U18144 (N_18144,N_17756,N_17769);
and U18145 (N_18145,N_17318,N_17355);
xor U18146 (N_18146,N_17025,N_17535);
xnor U18147 (N_18147,N_17421,N_17342);
or U18148 (N_18148,N_17609,N_17885);
nor U18149 (N_18149,N_17707,N_17656);
xnor U18150 (N_18150,N_17945,N_17124);
or U18151 (N_18151,N_17399,N_17276);
and U18152 (N_18152,N_17184,N_17377);
nand U18153 (N_18153,N_17257,N_17032);
nor U18154 (N_18154,N_17204,N_17465);
or U18155 (N_18155,N_17674,N_17844);
xnor U18156 (N_18156,N_17177,N_17992);
nor U18157 (N_18157,N_17950,N_17665);
nand U18158 (N_18158,N_17200,N_17961);
xnor U18159 (N_18159,N_17007,N_17838);
nor U18160 (N_18160,N_17763,N_17832);
nor U18161 (N_18161,N_17820,N_17784);
nor U18162 (N_18162,N_17734,N_17323);
nor U18163 (N_18163,N_17150,N_17778);
or U18164 (N_18164,N_17714,N_17522);
and U18165 (N_18165,N_17752,N_17212);
xnor U18166 (N_18166,N_17686,N_17238);
or U18167 (N_18167,N_17965,N_17631);
nor U18168 (N_18168,N_17461,N_17809);
and U18169 (N_18169,N_17468,N_17045);
nand U18170 (N_18170,N_17584,N_17777);
and U18171 (N_18171,N_17658,N_17090);
nand U18172 (N_18172,N_17259,N_17513);
or U18173 (N_18173,N_17718,N_17106);
xor U18174 (N_18174,N_17553,N_17915);
xnor U18175 (N_18175,N_17861,N_17938);
xnor U18176 (N_18176,N_17771,N_17454);
xor U18177 (N_18177,N_17427,N_17911);
xnor U18178 (N_18178,N_17626,N_17218);
and U18179 (N_18179,N_17596,N_17840);
nor U18180 (N_18180,N_17179,N_17412);
and U18181 (N_18181,N_17428,N_17751);
xor U18182 (N_18182,N_17659,N_17246);
nand U18183 (N_18183,N_17221,N_17643);
nand U18184 (N_18184,N_17333,N_17910);
nand U18185 (N_18185,N_17103,N_17396);
and U18186 (N_18186,N_17941,N_17872);
nand U18187 (N_18187,N_17041,N_17618);
nand U18188 (N_18188,N_17420,N_17810);
nor U18189 (N_18189,N_17366,N_17419);
xor U18190 (N_18190,N_17080,N_17167);
and U18191 (N_18191,N_17368,N_17802);
nand U18192 (N_18192,N_17766,N_17376);
nor U18193 (N_18193,N_17477,N_17732);
xnor U18194 (N_18194,N_17457,N_17700);
nand U18195 (N_18195,N_17111,N_17209);
and U18196 (N_18196,N_17552,N_17566);
xnor U18197 (N_18197,N_17796,N_17835);
nand U18198 (N_18198,N_17267,N_17972);
nand U18199 (N_18199,N_17985,N_17556);
nor U18200 (N_18200,N_17894,N_17589);
nand U18201 (N_18201,N_17195,N_17542);
nand U18202 (N_18202,N_17749,N_17773);
nor U18203 (N_18203,N_17068,N_17429);
and U18204 (N_18204,N_17162,N_17182);
nor U18205 (N_18205,N_17375,N_17823);
and U18206 (N_18206,N_17148,N_17334);
nor U18207 (N_18207,N_17655,N_17110);
nor U18208 (N_18208,N_17863,N_17451);
nor U18209 (N_18209,N_17940,N_17836);
and U18210 (N_18210,N_17669,N_17035);
or U18211 (N_18211,N_17930,N_17920);
nor U18212 (N_18212,N_17864,N_17675);
or U18213 (N_18213,N_17721,N_17653);
xor U18214 (N_18214,N_17155,N_17987);
or U18215 (N_18215,N_17813,N_17146);
nand U18216 (N_18216,N_17365,N_17374);
xor U18217 (N_18217,N_17272,N_17122);
xnor U18218 (N_18218,N_17853,N_17993);
xor U18219 (N_18219,N_17839,N_17425);
nand U18220 (N_18220,N_17775,N_17264);
and U18221 (N_18221,N_17578,N_17193);
nand U18222 (N_18222,N_17876,N_17943);
nand U18223 (N_18223,N_17250,N_17452);
nor U18224 (N_18224,N_17016,N_17959);
nor U18225 (N_18225,N_17243,N_17724);
nand U18226 (N_18226,N_17747,N_17995);
xor U18227 (N_18227,N_17074,N_17245);
xnor U18228 (N_18228,N_17967,N_17123);
nor U18229 (N_18229,N_17694,N_17038);
nand U18230 (N_18230,N_17014,N_17373);
or U18231 (N_18231,N_17191,N_17388);
nor U18232 (N_18232,N_17439,N_17023);
or U18233 (N_18233,N_17748,N_17302);
or U18234 (N_18234,N_17690,N_17758);
and U18235 (N_18235,N_17586,N_17064);
and U18236 (N_18236,N_17091,N_17303);
and U18237 (N_18237,N_17379,N_17466);
nand U18238 (N_18238,N_17390,N_17892);
and U18239 (N_18239,N_17305,N_17761);
nand U18240 (N_18240,N_17069,N_17808);
or U18241 (N_18241,N_17400,N_17590);
nand U18242 (N_18242,N_17389,N_17306);
nand U18243 (N_18243,N_17791,N_17438);
nor U18244 (N_18244,N_17299,N_17962);
nand U18245 (N_18245,N_17175,N_17121);
nand U18246 (N_18246,N_17190,N_17203);
and U18247 (N_18247,N_17627,N_17201);
or U18248 (N_18248,N_17433,N_17902);
or U18249 (N_18249,N_17188,N_17060);
or U18250 (N_18250,N_17779,N_17490);
nand U18251 (N_18251,N_17304,N_17180);
xnor U18252 (N_18252,N_17554,N_17538);
and U18253 (N_18253,N_17235,N_17765);
nand U18254 (N_18254,N_17592,N_17282);
and U18255 (N_18255,N_17112,N_17682);
and U18256 (N_18256,N_17252,N_17332);
xor U18257 (N_18257,N_17456,N_17801);
and U18258 (N_18258,N_17821,N_17255);
or U18259 (N_18259,N_17013,N_17344);
xor U18260 (N_18260,N_17574,N_17966);
nor U18261 (N_18261,N_17958,N_17345);
xor U18262 (N_18262,N_17786,N_17394);
or U18263 (N_18263,N_17611,N_17683);
and U18264 (N_18264,N_17169,N_17922);
nand U18265 (N_18265,N_17277,N_17816);
and U18266 (N_18266,N_17842,N_17012);
or U18267 (N_18267,N_17942,N_17540);
nand U18268 (N_18268,N_17363,N_17125);
or U18269 (N_18269,N_17848,N_17478);
nand U18270 (N_18270,N_17829,N_17983);
and U18271 (N_18271,N_17581,N_17371);
nand U18272 (N_18272,N_17852,N_17884);
or U18273 (N_18273,N_17622,N_17730);
or U18274 (N_18274,N_17684,N_17935);
nor U18275 (N_18275,N_17508,N_17480);
or U18276 (N_18276,N_17071,N_17077);
or U18277 (N_18277,N_17846,N_17603);
xnor U18278 (N_18278,N_17947,N_17900);
nand U18279 (N_18279,N_17978,N_17229);
and U18280 (N_18280,N_17331,N_17410);
and U18281 (N_18281,N_17954,N_17817);
and U18282 (N_18282,N_17691,N_17905);
or U18283 (N_18283,N_17455,N_17174);
nor U18284 (N_18284,N_17678,N_17253);
or U18285 (N_18285,N_17636,N_17974);
nand U18286 (N_18286,N_17673,N_17918);
xor U18287 (N_18287,N_17072,N_17537);
or U18288 (N_18288,N_17528,N_17189);
nor U18289 (N_18289,N_17316,N_17946);
nand U18290 (N_18290,N_17788,N_17879);
or U18291 (N_18291,N_17049,N_17698);
nand U18292 (N_18292,N_17448,N_17187);
or U18293 (N_18293,N_17326,N_17223);
nand U18294 (N_18294,N_17881,N_17790);
xor U18295 (N_18295,N_17163,N_17531);
or U18296 (N_18296,N_17398,N_17783);
nor U18297 (N_18297,N_17605,N_17649);
or U18298 (N_18298,N_17514,N_17044);
nor U18299 (N_18299,N_17330,N_17360);
or U18300 (N_18300,N_17434,N_17159);
nor U18301 (N_18301,N_17337,N_17803);
and U18302 (N_18302,N_17916,N_17679);
xnor U18303 (N_18303,N_17194,N_17311);
nor U18304 (N_18304,N_17845,N_17549);
and U18305 (N_18305,N_17491,N_17921);
or U18306 (N_18306,N_17133,N_17383);
and U18307 (N_18307,N_17782,N_17964);
and U18308 (N_18308,N_17093,N_17348);
or U18309 (N_18309,N_17492,N_17628);
xnor U18310 (N_18310,N_17031,N_17833);
or U18311 (N_18311,N_17939,N_17613);
and U18312 (N_18312,N_17024,N_17599);
and U18313 (N_18313,N_17099,N_17772);
nand U18314 (N_18314,N_17708,N_17851);
and U18315 (N_18315,N_17606,N_17114);
and U18316 (N_18316,N_17285,N_17571);
nand U18317 (N_18317,N_17367,N_17462);
or U18318 (N_18318,N_17176,N_17040);
nor U18319 (N_18319,N_17781,N_17716);
nor U18320 (N_18320,N_17140,N_17053);
nor U18321 (N_18321,N_17955,N_17270);
and U18322 (N_18322,N_17989,N_17612);
xnor U18323 (N_18323,N_17066,N_17166);
nor U18324 (N_18324,N_17422,N_17501);
and U18325 (N_18325,N_17338,N_17604);
xnor U18326 (N_18326,N_17341,N_17108);
nor U18327 (N_18327,N_17719,N_17914);
xor U18328 (N_18328,N_17648,N_17530);
nor U18329 (N_18329,N_17118,N_17937);
and U18330 (N_18330,N_17996,N_17960);
nand U18331 (N_18331,N_17139,N_17088);
or U18332 (N_18332,N_17630,N_17651);
xnor U18333 (N_18333,N_17661,N_17134);
xnor U18334 (N_18334,N_17020,N_17431);
nor U18335 (N_18335,N_17426,N_17062);
nor U18336 (N_18336,N_17539,N_17798);
and U18337 (N_18337,N_17181,N_17562);
nand U18338 (N_18338,N_17750,N_17739);
nand U18339 (N_18339,N_17882,N_17909);
xor U18340 (N_18340,N_17908,N_17744);
nor U18341 (N_18341,N_17011,N_17380);
nand U18342 (N_18342,N_17065,N_17711);
and U18343 (N_18343,N_17349,N_17317);
or U18344 (N_18344,N_17672,N_17241);
nor U18345 (N_18345,N_17199,N_17896);
nand U18346 (N_18346,N_17976,N_17865);
nor U18347 (N_18347,N_17866,N_17084);
xnor U18348 (N_18348,N_17867,N_17949);
or U18349 (N_18349,N_17561,N_17850);
and U18350 (N_18350,N_17575,N_17886);
nand U18351 (N_18351,N_17076,N_17213);
nand U18352 (N_18352,N_17493,N_17518);
xor U18353 (N_18353,N_17082,N_17356);
nor U18354 (N_18354,N_17688,N_17258);
nand U18355 (N_18355,N_17792,N_17639);
nand U18356 (N_18356,N_17207,N_17214);
nand U18357 (N_18357,N_17254,N_17545);
nand U18358 (N_18358,N_17230,N_17052);
and U18359 (N_18359,N_17265,N_17577);
and U18360 (N_18360,N_17889,N_17022);
xor U18361 (N_18361,N_17825,N_17369);
nor U18362 (N_18362,N_17715,N_17309);
nor U18363 (N_18363,N_17142,N_17353);
nor U18364 (N_18364,N_17907,N_17499);
nand U18365 (N_18365,N_17593,N_17587);
nand U18366 (N_18366,N_17205,N_17815);
or U18367 (N_18367,N_17158,N_17847);
nand U18368 (N_18368,N_17857,N_17116);
xnor U18369 (N_18369,N_17565,N_17704);
and U18370 (N_18370,N_17402,N_17002);
nor U18371 (N_18371,N_17227,N_17470);
nor U18372 (N_18372,N_17036,N_17312);
nor U18373 (N_18373,N_17009,N_17534);
nor U18374 (N_18374,N_17874,N_17897);
nand U18375 (N_18375,N_17260,N_17293);
nand U18376 (N_18376,N_17206,N_17637);
nand U18377 (N_18377,N_17812,N_17115);
nor U18378 (N_18378,N_17244,N_17449);
xnor U18379 (N_18379,N_17931,N_17471);
xnor U18380 (N_18380,N_17078,N_17151);
or U18381 (N_18381,N_17275,N_17927);
xnor U18382 (N_18382,N_17416,N_17620);
and U18383 (N_18383,N_17382,N_17067);
or U18384 (N_18384,N_17362,N_17936);
or U18385 (N_18385,N_17709,N_17296);
or U18386 (N_18386,N_17988,N_17871);
nor U18387 (N_18387,N_17551,N_17811);
xnor U18388 (N_18388,N_17615,N_17198);
and U18389 (N_18389,N_17269,N_17533);
or U18390 (N_18390,N_17314,N_17929);
nor U18391 (N_18391,N_17236,N_17986);
and U18392 (N_18392,N_17834,N_17215);
and U18393 (N_18393,N_17720,N_17977);
nor U18394 (N_18394,N_17095,N_17703);
nor U18395 (N_18395,N_17104,N_17256);
or U18396 (N_18396,N_17980,N_17695);
or U18397 (N_18397,N_17386,N_17232);
nand U18398 (N_18398,N_17346,N_17271);
and U18399 (N_18399,N_17216,N_17297);
nor U18400 (N_18400,N_17699,N_17495);
nor U18401 (N_18401,N_17647,N_17740);
nor U18402 (N_18402,N_17854,N_17211);
xnor U18403 (N_18403,N_17397,N_17004);
nor U18404 (N_18404,N_17475,N_17494);
nand U18405 (N_18405,N_17512,N_17287);
xor U18406 (N_18406,N_17497,N_17234);
xnor U18407 (N_18407,N_17619,N_17447);
xnor U18408 (N_18408,N_17437,N_17804);
or U18409 (N_18409,N_17153,N_17026);
or U18410 (N_18410,N_17144,N_17970);
and U18411 (N_18411,N_17650,N_17806);
and U18412 (N_18412,N_17336,N_17274);
nand U18413 (N_18413,N_17395,N_17680);
nor U18414 (N_18414,N_17767,N_17472);
or U18415 (N_18415,N_17868,N_17003);
xnor U18416 (N_18416,N_17654,N_17424);
xor U18417 (N_18417,N_17998,N_17089);
and U18418 (N_18418,N_17048,N_17325);
and U18419 (N_18419,N_17580,N_17109);
nand U18420 (N_18420,N_17405,N_17086);
and U18421 (N_18421,N_17079,N_17393);
and U18422 (N_18422,N_17143,N_17875);
and U18423 (N_18423,N_17352,N_17855);
and U18424 (N_18424,N_17242,N_17547);
nand U18425 (N_18425,N_17406,N_17805);
or U18426 (N_18426,N_17597,N_17776);
and U18427 (N_18427,N_17602,N_17638);
nor U18428 (N_18428,N_17681,N_17273);
nand U18429 (N_18429,N_17687,N_17413);
xor U18430 (N_18430,N_17445,N_17231);
or U18431 (N_18431,N_17526,N_17971);
or U18432 (N_18432,N_17572,N_17224);
nand U18433 (N_18433,N_17083,N_17476);
nor U18434 (N_18434,N_17828,N_17818);
or U18435 (N_18435,N_17795,N_17735);
xor U18436 (N_18436,N_17178,N_17755);
and U18437 (N_18437,N_17056,N_17926);
nand U18438 (N_18438,N_17291,N_17119);
and U18439 (N_18439,N_17666,N_17340);
and U18440 (N_18440,N_17800,N_17295);
or U18441 (N_18441,N_17843,N_17222);
and U18442 (N_18442,N_17519,N_17973);
and U18443 (N_18443,N_17050,N_17286);
nor U18444 (N_18444,N_17559,N_17668);
or U18445 (N_18445,N_17951,N_17787);
or U18446 (N_18446,N_17624,N_17546);
nor U18447 (N_18447,N_17436,N_17928);
and U18448 (N_18448,N_17521,N_17381);
nor U18449 (N_18449,N_17046,N_17321);
xor U18450 (N_18450,N_17689,N_17984);
or U18451 (N_18451,N_17878,N_17723);
nor U18452 (N_18452,N_17037,N_17481);
or U18453 (N_18453,N_17757,N_17634);
or U18454 (N_18454,N_17407,N_17525);
and U18455 (N_18455,N_17567,N_17320);
xnor U18456 (N_18456,N_17102,N_17168);
or U18457 (N_18457,N_17994,N_17895);
nand U18458 (N_18458,N_17667,N_17505);
or U18459 (N_18459,N_17642,N_17327);
nor U18460 (N_18460,N_17423,N_17027);
xor U18461 (N_18461,N_17608,N_17029);
nor U18462 (N_18462,N_17741,N_17292);
and U18463 (N_18463,N_17217,N_17543);
xor U18464 (N_18464,N_17725,N_17904);
and U18465 (N_18465,N_17051,N_17008);
nand U18466 (N_18466,N_17919,N_17432);
xnor U18467 (N_18467,N_17712,N_17952);
or U18468 (N_18468,N_17506,N_17746);
nor U18469 (N_18469,N_17819,N_17171);
xnor U18470 (N_18470,N_17742,N_17826);
and U18471 (N_18471,N_17849,N_17010);
xnor U18472 (N_18472,N_17164,N_17664);
and U18473 (N_18473,N_17517,N_17085);
or U18474 (N_18474,N_17822,N_17507);
or U18475 (N_18475,N_17359,N_17729);
nand U18476 (N_18476,N_17585,N_17706);
xor U18477 (N_18477,N_17343,N_17030);
and U18478 (N_18478,N_17906,N_17877);
nand U18479 (N_18479,N_17132,N_17058);
nand U18480 (N_18480,N_17120,N_17573);
or U18481 (N_18481,N_17558,N_17924);
xor U18482 (N_18482,N_17858,N_17098);
xor U18483 (N_18483,N_17953,N_17770);
nand U18484 (N_18484,N_17524,N_17923);
nor U18485 (N_18485,N_17841,N_17717);
and U18486 (N_18486,N_17625,N_17308);
nor U18487 (N_18487,N_17042,N_17728);
or U18488 (N_18488,N_17147,N_17883);
or U18489 (N_18489,N_17579,N_17136);
nor U18490 (N_18490,N_17226,N_17520);
or U18491 (N_18491,N_17632,N_17054);
or U18492 (N_18492,N_17697,N_17183);
xor U18493 (N_18493,N_17797,N_17598);
nand U18494 (N_18494,N_17616,N_17307);
or U18495 (N_18495,N_17202,N_17670);
xnor U18496 (N_18496,N_17640,N_17641);
and U18497 (N_18497,N_17251,N_17831);
nor U18498 (N_18498,N_17322,N_17351);
and U18499 (N_18499,N_17197,N_17887);
and U18500 (N_18500,N_17037,N_17022);
or U18501 (N_18501,N_17023,N_17050);
or U18502 (N_18502,N_17196,N_17370);
or U18503 (N_18503,N_17952,N_17220);
nand U18504 (N_18504,N_17604,N_17263);
xnor U18505 (N_18505,N_17664,N_17588);
xnor U18506 (N_18506,N_17311,N_17178);
nand U18507 (N_18507,N_17854,N_17700);
nand U18508 (N_18508,N_17377,N_17167);
nor U18509 (N_18509,N_17654,N_17188);
nor U18510 (N_18510,N_17647,N_17920);
nand U18511 (N_18511,N_17170,N_17438);
nand U18512 (N_18512,N_17924,N_17659);
nand U18513 (N_18513,N_17132,N_17999);
and U18514 (N_18514,N_17351,N_17756);
xnor U18515 (N_18515,N_17192,N_17930);
or U18516 (N_18516,N_17533,N_17896);
nor U18517 (N_18517,N_17365,N_17384);
nor U18518 (N_18518,N_17860,N_17295);
nor U18519 (N_18519,N_17807,N_17884);
xnor U18520 (N_18520,N_17311,N_17689);
or U18521 (N_18521,N_17293,N_17770);
or U18522 (N_18522,N_17578,N_17420);
nor U18523 (N_18523,N_17298,N_17203);
nor U18524 (N_18524,N_17410,N_17060);
xor U18525 (N_18525,N_17720,N_17202);
or U18526 (N_18526,N_17708,N_17188);
nand U18527 (N_18527,N_17609,N_17852);
or U18528 (N_18528,N_17231,N_17855);
and U18529 (N_18529,N_17578,N_17525);
nor U18530 (N_18530,N_17918,N_17484);
and U18531 (N_18531,N_17960,N_17270);
or U18532 (N_18532,N_17753,N_17479);
nand U18533 (N_18533,N_17750,N_17426);
or U18534 (N_18534,N_17846,N_17924);
and U18535 (N_18535,N_17405,N_17477);
nand U18536 (N_18536,N_17565,N_17470);
nand U18537 (N_18537,N_17325,N_17804);
nand U18538 (N_18538,N_17516,N_17732);
xnor U18539 (N_18539,N_17309,N_17484);
and U18540 (N_18540,N_17150,N_17303);
nor U18541 (N_18541,N_17869,N_17647);
xor U18542 (N_18542,N_17267,N_17098);
nand U18543 (N_18543,N_17555,N_17040);
xor U18544 (N_18544,N_17577,N_17437);
nor U18545 (N_18545,N_17145,N_17676);
or U18546 (N_18546,N_17882,N_17032);
or U18547 (N_18547,N_17926,N_17567);
nor U18548 (N_18548,N_17850,N_17128);
nor U18549 (N_18549,N_17311,N_17299);
nand U18550 (N_18550,N_17334,N_17761);
and U18551 (N_18551,N_17064,N_17160);
nor U18552 (N_18552,N_17282,N_17020);
nor U18553 (N_18553,N_17490,N_17859);
nor U18554 (N_18554,N_17533,N_17450);
and U18555 (N_18555,N_17831,N_17937);
nor U18556 (N_18556,N_17931,N_17286);
nand U18557 (N_18557,N_17242,N_17255);
or U18558 (N_18558,N_17706,N_17118);
or U18559 (N_18559,N_17548,N_17841);
nand U18560 (N_18560,N_17003,N_17772);
or U18561 (N_18561,N_17048,N_17104);
nor U18562 (N_18562,N_17825,N_17614);
or U18563 (N_18563,N_17113,N_17323);
xor U18564 (N_18564,N_17242,N_17252);
nand U18565 (N_18565,N_17038,N_17866);
or U18566 (N_18566,N_17159,N_17164);
xor U18567 (N_18567,N_17773,N_17102);
nor U18568 (N_18568,N_17481,N_17347);
nand U18569 (N_18569,N_17572,N_17118);
xnor U18570 (N_18570,N_17115,N_17959);
and U18571 (N_18571,N_17370,N_17449);
and U18572 (N_18572,N_17078,N_17270);
or U18573 (N_18573,N_17344,N_17102);
xor U18574 (N_18574,N_17027,N_17426);
nor U18575 (N_18575,N_17930,N_17967);
nand U18576 (N_18576,N_17887,N_17304);
nor U18577 (N_18577,N_17224,N_17602);
xnor U18578 (N_18578,N_17542,N_17868);
or U18579 (N_18579,N_17775,N_17292);
xnor U18580 (N_18580,N_17016,N_17313);
or U18581 (N_18581,N_17199,N_17553);
nand U18582 (N_18582,N_17822,N_17440);
or U18583 (N_18583,N_17143,N_17310);
nand U18584 (N_18584,N_17309,N_17325);
nand U18585 (N_18585,N_17026,N_17365);
and U18586 (N_18586,N_17486,N_17858);
and U18587 (N_18587,N_17693,N_17948);
or U18588 (N_18588,N_17542,N_17576);
xnor U18589 (N_18589,N_17702,N_17625);
and U18590 (N_18590,N_17482,N_17798);
or U18591 (N_18591,N_17870,N_17969);
or U18592 (N_18592,N_17054,N_17820);
nand U18593 (N_18593,N_17580,N_17459);
xor U18594 (N_18594,N_17160,N_17582);
and U18595 (N_18595,N_17241,N_17582);
and U18596 (N_18596,N_17331,N_17222);
xor U18597 (N_18597,N_17136,N_17147);
or U18598 (N_18598,N_17223,N_17133);
xnor U18599 (N_18599,N_17096,N_17814);
nor U18600 (N_18600,N_17967,N_17434);
and U18601 (N_18601,N_17315,N_17869);
xor U18602 (N_18602,N_17721,N_17325);
nand U18603 (N_18603,N_17963,N_17183);
and U18604 (N_18604,N_17550,N_17191);
xor U18605 (N_18605,N_17008,N_17652);
or U18606 (N_18606,N_17195,N_17345);
xor U18607 (N_18607,N_17836,N_17863);
and U18608 (N_18608,N_17362,N_17923);
nor U18609 (N_18609,N_17036,N_17241);
nor U18610 (N_18610,N_17724,N_17702);
and U18611 (N_18611,N_17088,N_17025);
nor U18612 (N_18612,N_17719,N_17243);
or U18613 (N_18613,N_17295,N_17374);
or U18614 (N_18614,N_17774,N_17705);
nand U18615 (N_18615,N_17487,N_17694);
nor U18616 (N_18616,N_17733,N_17745);
xnor U18617 (N_18617,N_17252,N_17137);
nor U18618 (N_18618,N_17620,N_17616);
and U18619 (N_18619,N_17968,N_17058);
xor U18620 (N_18620,N_17468,N_17611);
nand U18621 (N_18621,N_17189,N_17653);
or U18622 (N_18622,N_17482,N_17531);
and U18623 (N_18623,N_17907,N_17609);
or U18624 (N_18624,N_17462,N_17958);
or U18625 (N_18625,N_17359,N_17409);
or U18626 (N_18626,N_17650,N_17011);
or U18627 (N_18627,N_17788,N_17444);
or U18628 (N_18628,N_17778,N_17640);
xor U18629 (N_18629,N_17848,N_17963);
nand U18630 (N_18630,N_17238,N_17565);
and U18631 (N_18631,N_17415,N_17852);
nor U18632 (N_18632,N_17649,N_17659);
xnor U18633 (N_18633,N_17319,N_17506);
or U18634 (N_18634,N_17307,N_17941);
or U18635 (N_18635,N_17433,N_17510);
or U18636 (N_18636,N_17017,N_17012);
and U18637 (N_18637,N_17853,N_17209);
nand U18638 (N_18638,N_17485,N_17779);
xor U18639 (N_18639,N_17689,N_17509);
or U18640 (N_18640,N_17845,N_17885);
nand U18641 (N_18641,N_17375,N_17580);
nor U18642 (N_18642,N_17119,N_17413);
nor U18643 (N_18643,N_17108,N_17889);
and U18644 (N_18644,N_17754,N_17659);
nand U18645 (N_18645,N_17794,N_17781);
and U18646 (N_18646,N_17081,N_17328);
nor U18647 (N_18647,N_17784,N_17744);
and U18648 (N_18648,N_17024,N_17396);
or U18649 (N_18649,N_17973,N_17017);
nor U18650 (N_18650,N_17804,N_17993);
and U18651 (N_18651,N_17284,N_17662);
or U18652 (N_18652,N_17407,N_17008);
nand U18653 (N_18653,N_17327,N_17691);
nand U18654 (N_18654,N_17345,N_17157);
and U18655 (N_18655,N_17956,N_17887);
nand U18656 (N_18656,N_17658,N_17654);
nand U18657 (N_18657,N_17583,N_17991);
xor U18658 (N_18658,N_17093,N_17916);
nand U18659 (N_18659,N_17835,N_17860);
nor U18660 (N_18660,N_17286,N_17257);
nand U18661 (N_18661,N_17372,N_17601);
xnor U18662 (N_18662,N_17731,N_17900);
xor U18663 (N_18663,N_17333,N_17595);
or U18664 (N_18664,N_17370,N_17651);
xor U18665 (N_18665,N_17121,N_17509);
xnor U18666 (N_18666,N_17471,N_17613);
xor U18667 (N_18667,N_17894,N_17875);
xnor U18668 (N_18668,N_17882,N_17091);
or U18669 (N_18669,N_17407,N_17947);
nor U18670 (N_18670,N_17652,N_17302);
or U18671 (N_18671,N_17027,N_17321);
or U18672 (N_18672,N_17386,N_17332);
and U18673 (N_18673,N_17009,N_17320);
xor U18674 (N_18674,N_17093,N_17900);
nor U18675 (N_18675,N_17996,N_17040);
nand U18676 (N_18676,N_17981,N_17147);
or U18677 (N_18677,N_17542,N_17292);
nand U18678 (N_18678,N_17755,N_17125);
xor U18679 (N_18679,N_17793,N_17851);
or U18680 (N_18680,N_17454,N_17162);
nor U18681 (N_18681,N_17523,N_17806);
nand U18682 (N_18682,N_17530,N_17050);
or U18683 (N_18683,N_17858,N_17119);
nor U18684 (N_18684,N_17882,N_17012);
or U18685 (N_18685,N_17444,N_17648);
nand U18686 (N_18686,N_17098,N_17447);
xnor U18687 (N_18687,N_17684,N_17215);
xnor U18688 (N_18688,N_17816,N_17753);
nand U18689 (N_18689,N_17103,N_17756);
xnor U18690 (N_18690,N_17197,N_17082);
or U18691 (N_18691,N_17690,N_17532);
nand U18692 (N_18692,N_17051,N_17037);
or U18693 (N_18693,N_17374,N_17105);
nor U18694 (N_18694,N_17739,N_17245);
or U18695 (N_18695,N_17067,N_17938);
or U18696 (N_18696,N_17875,N_17394);
or U18697 (N_18697,N_17019,N_17854);
nor U18698 (N_18698,N_17743,N_17628);
nand U18699 (N_18699,N_17653,N_17884);
nand U18700 (N_18700,N_17852,N_17697);
nand U18701 (N_18701,N_17388,N_17570);
and U18702 (N_18702,N_17517,N_17849);
nand U18703 (N_18703,N_17571,N_17232);
or U18704 (N_18704,N_17377,N_17727);
nor U18705 (N_18705,N_17749,N_17959);
or U18706 (N_18706,N_17069,N_17922);
nand U18707 (N_18707,N_17576,N_17660);
or U18708 (N_18708,N_17857,N_17425);
nor U18709 (N_18709,N_17590,N_17440);
and U18710 (N_18710,N_17451,N_17758);
nor U18711 (N_18711,N_17063,N_17566);
nand U18712 (N_18712,N_17811,N_17834);
and U18713 (N_18713,N_17948,N_17214);
and U18714 (N_18714,N_17265,N_17596);
nand U18715 (N_18715,N_17179,N_17107);
or U18716 (N_18716,N_17524,N_17713);
or U18717 (N_18717,N_17089,N_17737);
nand U18718 (N_18718,N_17767,N_17129);
nor U18719 (N_18719,N_17686,N_17786);
and U18720 (N_18720,N_17204,N_17301);
or U18721 (N_18721,N_17954,N_17275);
nand U18722 (N_18722,N_17488,N_17949);
nand U18723 (N_18723,N_17440,N_17164);
or U18724 (N_18724,N_17366,N_17436);
nand U18725 (N_18725,N_17017,N_17019);
nand U18726 (N_18726,N_17060,N_17102);
or U18727 (N_18727,N_17448,N_17968);
xnor U18728 (N_18728,N_17408,N_17890);
nor U18729 (N_18729,N_17219,N_17964);
xnor U18730 (N_18730,N_17159,N_17102);
nand U18731 (N_18731,N_17551,N_17128);
nor U18732 (N_18732,N_17784,N_17868);
and U18733 (N_18733,N_17425,N_17728);
nand U18734 (N_18734,N_17059,N_17290);
or U18735 (N_18735,N_17554,N_17048);
xnor U18736 (N_18736,N_17062,N_17686);
nor U18737 (N_18737,N_17704,N_17836);
and U18738 (N_18738,N_17961,N_17522);
nor U18739 (N_18739,N_17505,N_17067);
or U18740 (N_18740,N_17590,N_17748);
nand U18741 (N_18741,N_17385,N_17331);
or U18742 (N_18742,N_17077,N_17643);
xor U18743 (N_18743,N_17303,N_17055);
nor U18744 (N_18744,N_17241,N_17767);
nor U18745 (N_18745,N_17472,N_17793);
nand U18746 (N_18746,N_17943,N_17848);
xnor U18747 (N_18747,N_17171,N_17216);
xor U18748 (N_18748,N_17478,N_17750);
or U18749 (N_18749,N_17063,N_17284);
and U18750 (N_18750,N_17236,N_17251);
nor U18751 (N_18751,N_17275,N_17278);
or U18752 (N_18752,N_17390,N_17122);
nor U18753 (N_18753,N_17572,N_17004);
xnor U18754 (N_18754,N_17276,N_17470);
or U18755 (N_18755,N_17785,N_17872);
or U18756 (N_18756,N_17582,N_17580);
or U18757 (N_18757,N_17866,N_17064);
and U18758 (N_18758,N_17086,N_17469);
and U18759 (N_18759,N_17904,N_17167);
nand U18760 (N_18760,N_17416,N_17638);
nor U18761 (N_18761,N_17122,N_17072);
xor U18762 (N_18762,N_17593,N_17125);
nand U18763 (N_18763,N_17523,N_17189);
nand U18764 (N_18764,N_17938,N_17773);
nor U18765 (N_18765,N_17212,N_17596);
xor U18766 (N_18766,N_17406,N_17614);
and U18767 (N_18767,N_17160,N_17261);
nand U18768 (N_18768,N_17537,N_17752);
and U18769 (N_18769,N_17290,N_17891);
nand U18770 (N_18770,N_17698,N_17591);
or U18771 (N_18771,N_17056,N_17773);
and U18772 (N_18772,N_17643,N_17717);
nand U18773 (N_18773,N_17694,N_17655);
nand U18774 (N_18774,N_17170,N_17175);
and U18775 (N_18775,N_17389,N_17961);
nand U18776 (N_18776,N_17377,N_17670);
nor U18777 (N_18777,N_17299,N_17805);
and U18778 (N_18778,N_17071,N_17168);
nand U18779 (N_18779,N_17794,N_17612);
nand U18780 (N_18780,N_17694,N_17155);
xnor U18781 (N_18781,N_17861,N_17396);
xor U18782 (N_18782,N_17797,N_17094);
nand U18783 (N_18783,N_17131,N_17782);
nor U18784 (N_18784,N_17236,N_17035);
xor U18785 (N_18785,N_17222,N_17129);
nand U18786 (N_18786,N_17195,N_17153);
or U18787 (N_18787,N_17890,N_17158);
nand U18788 (N_18788,N_17743,N_17820);
nand U18789 (N_18789,N_17681,N_17497);
nor U18790 (N_18790,N_17477,N_17102);
nor U18791 (N_18791,N_17763,N_17030);
xor U18792 (N_18792,N_17594,N_17819);
nor U18793 (N_18793,N_17575,N_17356);
and U18794 (N_18794,N_17600,N_17007);
nor U18795 (N_18795,N_17475,N_17437);
xnor U18796 (N_18796,N_17728,N_17345);
xor U18797 (N_18797,N_17292,N_17796);
nand U18798 (N_18798,N_17570,N_17927);
and U18799 (N_18799,N_17429,N_17328);
nand U18800 (N_18800,N_17647,N_17714);
and U18801 (N_18801,N_17276,N_17574);
nand U18802 (N_18802,N_17961,N_17668);
and U18803 (N_18803,N_17176,N_17136);
xnor U18804 (N_18804,N_17371,N_17321);
or U18805 (N_18805,N_17678,N_17979);
nor U18806 (N_18806,N_17507,N_17523);
xor U18807 (N_18807,N_17593,N_17486);
nor U18808 (N_18808,N_17042,N_17018);
or U18809 (N_18809,N_17761,N_17050);
and U18810 (N_18810,N_17592,N_17392);
nor U18811 (N_18811,N_17408,N_17746);
or U18812 (N_18812,N_17938,N_17186);
nand U18813 (N_18813,N_17710,N_17484);
or U18814 (N_18814,N_17463,N_17297);
or U18815 (N_18815,N_17226,N_17395);
or U18816 (N_18816,N_17944,N_17993);
xor U18817 (N_18817,N_17404,N_17998);
xnor U18818 (N_18818,N_17994,N_17885);
or U18819 (N_18819,N_17299,N_17675);
and U18820 (N_18820,N_17741,N_17115);
nor U18821 (N_18821,N_17590,N_17551);
xor U18822 (N_18822,N_17527,N_17210);
xor U18823 (N_18823,N_17625,N_17942);
or U18824 (N_18824,N_17157,N_17410);
nor U18825 (N_18825,N_17581,N_17613);
nand U18826 (N_18826,N_17096,N_17629);
and U18827 (N_18827,N_17198,N_17121);
nor U18828 (N_18828,N_17387,N_17800);
or U18829 (N_18829,N_17743,N_17967);
xnor U18830 (N_18830,N_17989,N_17068);
nor U18831 (N_18831,N_17426,N_17625);
xor U18832 (N_18832,N_17578,N_17509);
and U18833 (N_18833,N_17760,N_17349);
nor U18834 (N_18834,N_17641,N_17859);
nand U18835 (N_18835,N_17228,N_17784);
nand U18836 (N_18836,N_17413,N_17438);
nor U18837 (N_18837,N_17860,N_17185);
nor U18838 (N_18838,N_17759,N_17554);
or U18839 (N_18839,N_17958,N_17336);
and U18840 (N_18840,N_17405,N_17275);
or U18841 (N_18841,N_17491,N_17681);
and U18842 (N_18842,N_17031,N_17283);
nor U18843 (N_18843,N_17355,N_17883);
or U18844 (N_18844,N_17118,N_17773);
nor U18845 (N_18845,N_17949,N_17070);
and U18846 (N_18846,N_17607,N_17956);
nand U18847 (N_18847,N_17927,N_17184);
or U18848 (N_18848,N_17034,N_17909);
or U18849 (N_18849,N_17094,N_17687);
nand U18850 (N_18850,N_17126,N_17594);
xnor U18851 (N_18851,N_17774,N_17128);
and U18852 (N_18852,N_17914,N_17974);
and U18853 (N_18853,N_17336,N_17111);
nor U18854 (N_18854,N_17479,N_17247);
or U18855 (N_18855,N_17777,N_17896);
and U18856 (N_18856,N_17479,N_17802);
or U18857 (N_18857,N_17028,N_17918);
nor U18858 (N_18858,N_17410,N_17414);
and U18859 (N_18859,N_17322,N_17198);
xnor U18860 (N_18860,N_17417,N_17725);
or U18861 (N_18861,N_17626,N_17405);
and U18862 (N_18862,N_17752,N_17476);
or U18863 (N_18863,N_17879,N_17829);
nor U18864 (N_18864,N_17110,N_17062);
and U18865 (N_18865,N_17214,N_17390);
xor U18866 (N_18866,N_17732,N_17699);
or U18867 (N_18867,N_17001,N_17389);
xor U18868 (N_18868,N_17859,N_17771);
nand U18869 (N_18869,N_17564,N_17652);
nand U18870 (N_18870,N_17361,N_17079);
and U18871 (N_18871,N_17159,N_17667);
xnor U18872 (N_18872,N_17797,N_17589);
nor U18873 (N_18873,N_17590,N_17705);
xor U18874 (N_18874,N_17685,N_17044);
or U18875 (N_18875,N_17042,N_17596);
nand U18876 (N_18876,N_17063,N_17904);
and U18877 (N_18877,N_17775,N_17809);
nor U18878 (N_18878,N_17599,N_17094);
nand U18879 (N_18879,N_17382,N_17039);
and U18880 (N_18880,N_17797,N_17707);
and U18881 (N_18881,N_17682,N_17851);
nand U18882 (N_18882,N_17575,N_17790);
nor U18883 (N_18883,N_17145,N_17149);
and U18884 (N_18884,N_17124,N_17383);
nor U18885 (N_18885,N_17201,N_17319);
and U18886 (N_18886,N_17883,N_17774);
nand U18887 (N_18887,N_17426,N_17519);
nor U18888 (N_18888,N_17790,N_17563);
nor U18889 (N_18889,N_17711,N_17512);
nand U18890 (N_18890,N_17823,N_17137);
or U18891 (N_18891,N_17307,N_17264);
and U18892 (N_18892,N_17011,N_17451);
and U18893 (N_18893,N_17262,N_17025);
nor U18894 (N_18894,N_17450,N_17201);
xnor U18895 (N_18895,N_17543,N_17602);
nand U18896 (N_18896,N_17370,N_17114);
and U18897 (N_18897,N_17511,N_17539);
nand U18898 (N_18898,N_17842,N_17607);
nand U18899 (N_18899,N_17541,N_17164);
xor U18900 (N_18900,N_17123,N_17638);
nand U18901 (N_18901,N_17090,N_17322);
xnor U18902 (N_18902,N_17857,N_17871);
xnor U18903 (N_18903,N_17056,N_17677);
or U18904 (N_18904,N_17049,N_17210);
nand U18905 (N_18905,N_17379,N_17039);
nor U18906 (N_18906,N_17879,N_17894);
nor U18907 (N_18907,N_17027,N_17585);
nor U18908 (N_18908,N_17230,N_17511);
nand U18909 (N_18909,N_17750,N_17530);
nor U18910 (N_18910,N_17089,N_17327);
nand U18911 (N_18911,N_17389,N_17041);
nand U18912 (N_18912,N_17937,N_17952);
nand U18913 (N_18913,N_17632,N_17334);
xor U18914 (N_18914,N_17552,N_17197);
and U18915 (N_18915,N_17541,N_17198);
xnor U18916 (N_18916,N_17586,N_17330);
nor U18917 (N_18917,N_17609,N_17133);
xnor U18918 (N_18918,N_17470,N_17531);
or U18919 (N_18919,N_17288,N_17224);
nand U18920 (N_18920,N_17061,N_17857);
or U18921 (N_18921,N_17784,N_17412);
xnor U18922 (N_18922,N_17627,N_17664);
or U18923 (N_18923,N_17259,N_17331);
and U18924 (N_18924,N_17490,N_17151);
or U18925 (N_18925,N_17639,N_17906);
xor U18926 (N_18926,N_17810,N_17960);
and U18927 (N_18927,N_17030,N_17797);
xnor U18928 (N_18928,N_17057,N_17332);
and U18929 (N_18929,N_17282,N_17155);
xnor U18930 (N_18930,N_17050,N_17593);
xor U18931 (N_18931,N_17368,N_17187);
or U18932 (N_18932,N_17591,N_17757);
nand U18933 (N_18933,N_17381,N_17360);
or U18934 (N_18934,N_17360,N_17763);
and U18935 (N_18935,N_17292,N_17506);
and U18936 (N_18936,N_17291,N_17744);
nand U18937 (N_18937,N_17404,N_17346);
nand U18938 (N_18938,N_17148,N_17098);
nor U18939 (N_18939,N_17673,N_17203);
nor U18940 (N_18940,N_17132,N_17072);
or U18941 (N_18941,N_17684,N_17758);
nand U18942 (N_18942,N_17119,N_17137);
and U18943 (N_18943,N_17811,N_17067);
nand U18944 (N_18944,N_17607,N_17085);
or U18945 (N_18945,N_17182,N_17915);
and U18946 (N_18946,N_17976,N_17022);
or U18947 (N_18947,N_17782,N_17603);
xor U18948 (N_18948,N_17778,N_17431);
and U18949 (N_18949,N_17934,N_17055);
nor U18950 (N_18950,N_17738,N_17122);
nand U18951 (N_18951,N_17835,N_17382);
xnor U18952 (N_18952,N_17310,N_17788);
and U18953 (N_18953,N_17915,N_17927);
or U18954 (N_18954,N_17381,N_17145);
nor U18955 (N_18955,N_17043,N_17248);
and U18956 (N_18956,N_17649,N_17002);
xnor U18957 (N_18957,N_17580,N_17280);
nor U18958 (N_18958,N_17865,N_17433);
or U18959 (N_18959,N_17972,N_17662);
nor U18960 (N_18960,N_17089,N_17911);
xor U18961 (N_18961,N_17488,N_17569);
xor U18962 (N_18962,N_17170,N_17816);
nor U18963 (N_18963,N_17729,N_17460);
or U18964 (N_18964,N_17784,N_17764);
nand U18965 (N_18965,N_17239,N_17315);
nand U18966 (N_18966,N_17841,N_17668);
or U18967 (N_18967,N_17072,N_17206);
nor U18968 (N_18968,N_17950,N_17362);
nor U18969 (N_18969,N_17593,N_17461);
xor U18970 (N_18970,N_17190,N_17237);
and U18971 (N_18971,N_17168,N_17824);
and U18972 (N_18972,N_17758,N_17180);
nor U18973 (N_18973,N_17926,N_17492);
nand U18974 (N_18974,N_17700,N_17831);
nor U18975 (N_18975,N_17977,N_17808);
or U18976 (N_18976,N_17428,N_17337);
nor U18977 (N_18977,N_17454,N_17577);
xor U18978 (N_18978,N_17591,N_17522);
or U18979 (N_18979,N_17228,N_17724);
nand U18980 (N_18980,N_17691,N_17362);
or U18981 (N_18981,N_17500,N_17631);
or U18982 (N_18982,N_17905,N_17006);
or U18983 (N_18983,N_17509,N_17573);
and U18984 (N_18984,N_17247,N_17287);
nor U18985 (N_18985,N_17171,N_17653);
nor U18986 (N_18986,N_17255,N_17672);
xnor U18987 (N_18987,N_17055,N_17473);
or U18988 (N_18988,N_17109,N_17923);
xor U18989 (N_18989,N_17775,N_17383);
or U18990 (N_18990,N_17717,N_17576);
and U18991 (N_18991,N_17651,N_17734);
or U18992 (N_18992,N_17122,N_17927);
nand U18993 (N_18993,N_17892,N_17154);
nor U18994 (N_18994,N_17033,N_17647);
or U18995 (N_18995,N_17861,N_17129);
nand U18996 (N_18996,N_17283,N_17869);
nand U18997 (N_18997,N_17603,N_17594);
nor U18998 (N_18998,N_17751,N_17695);
nor U18999 (N_18999,N_17552,N_17594);
nor U19000 (N_19000,N_18027,N_18783);
xnor U19001 (N_19001,N_18011,N_18670);
xor U19002 (N_19002,N_18804,N_18141);
or U19003 (N_19003,N_18662,N_18581);
xor U19004 (N_19004,N_18533,N_18404);
nand U19005 (N_19005,N_18177,N_18343);
or U19006 (N_19006,N_18288,N_18787);
or U19007 (N_19007,N_18201,N_18120);
and U19008 (N_19008,N_18644,N_18504);
nor U19009 (N_19009,N_18016,N_18843);
or U19010 (N_19010,N_18164,N_18582);
nand U19011 (N_19011,N_18736,N_18926);
xor U19012 (N_19012,N_18964,N_18517);
xor U19013 (N_19013,N_18388,N_18538);
xor U19014 (N_19014,N_18544,N_18985);
xor U19015 (N_19015,N_18317,N_18309);
nand U19016 (N_19016,N_18116,N_18329);
or U19017 (N_19017,N_18932,N_18520);
nor U19018 (N_19018,N_18879,N_18398);
and U19019 (N_19019,N_18363,N_18725);
or U19020 (N_19020,N_18383,N_18527);
and U19021 (N_19021,N_18434,N_18456);
or U19022 (N_19022,N_18933,N_18962);
or U19023 (N_19023,N_18245,N_18026);
and U19024 (N_19024,N_18441,N_18983);
nor U19025 (N_19025,N_18485,N_18679);
or U19026 (N_19026,N_18753,N_18058);
nor U19027 (N_19027,N_18945,N_18439);
or U19028 (N_19028,N_18483,N_18209);
nand U19029 (N_19029,N_18336,N_18091);
nor U19030 (N_19030,N_18493,N_18134);
nor U19031 (N_19031,N_18350,N_18673);
xnor U19032 (N_19032,N_18816,N_18811);
and U19033 (N_19033,N_18303,N_18478);
and U19034 (N_19034,N_18198,N_18488);
xnor U19035 (N_19035,N_18023,N_18427);
or U19036 (N_19036,N_18664,N_18676);
and U19037 (N_19037,N_18081,N_18376);
or U19038 (N_19038,N_18524,N_18796);
and U19039 (N_19039,N_18819,N_18460);
xor U19040 (N_19040,N_18642,N_18684);
nand U19041 (N_19041,N_18829,N_18998);
nor U19042 (N_19042,N_18745,N_18692);
nand U19043 (N_19043,N_18609,N_18698);
and U19044 (N_19044,N_18824,N_18680);
nand U19045 (N_19045,N_18121,N_18557);
nand U19046 (N_19046,N_18860,N_18916);
or U19047 (N_19047,N_18778,N_18211);
nand U19048 (N_19048,N_18085,N_18279);
nor U19049 (N_19049,N_18165,N_18827);
xnor U19050 (N_19050,N_18506,N_18666);
nand U19051 (N_19051,N_18794,N_18661);
or U19052 (N_19052,N_18740,N_18019);
or U19053 (N_19053,N_18853,N_18625);
or U19054 (N_19054,N_18175,N_18627);
and U19055 (N_19055,N_18668,N_18179);
or U19056 (N_19056,N_18088,N_18244);
and U19057 (N_19057,N_18210,N_18115);
and U19058 (N_19058,N_18521,N_18462);
nand U19059 (N_19059,N_18415,N_18872);
nand U19060 (N_19060,N_18021,N_18813);
or U19061 (N_19061,N_18820,N_18486);
nand U19062 (N_19062,N_18311,N_18381);
xnor U19063 (N_19063,N_18906,N_18910);
nand U19064 (N_19064,N_18247,N_18845);
and U19065 (N_19065,N_18312,N_18480);
nor U19066 (N_19066,N_18821,N_18596);
nand U19067 (N_19067,N_18534,N_18632);
and U19068 (N_19068,N_18864,N_18737);
xor U19069 (N_19069,N_18575,N_18633);
and U19070 (N_19070,N_18730,N_18743);
and U19071 (N_19071,N_18638,N_18428);
or U19072 (N_19072,N_18856,N_18254);
nand U19073 (N_19073,N_18050,N_18178);
nand U19074 (N_19074,N_18759,N_18919);
nor U19075 (N_19075,N_18941,N_18555);
or U19076 (N_19076,N_18571,N_18358);
nor U19077 (N_19077,N_18189,N_18808);
and U19078 (N_19078,N_18681,N_18741);
and U19079 (N_19079,N_18265,N_18216);
xnor U19080 (N_19080,N_18780,N_18482);
or U19081 (N_19081,N_18589,N_18903);
nand U19082 (N_19082,N_18977,N_18747);
or U19083 (N_19083,N_18257,N_18971);
and U19084 (N_19084,N_18733,N_18296);
and U19085 (N_19085,N_18731,N_18767);
xor U19086 (N_19086,N_18286,N_18242);
xor U19087 (N_19087,N_18539,N_18657);
or U19088 (N_19088,N_18547,N_18142);
xnor U19089 (N_19089,N_18861,N_18444);
nand U19090 (N_19090,N_18801,N_18776);
xor U19091 (N_19091,N_18908,N_18221);
or U19092 (N_19092,N_18621,N_18931);
nand U19093 (N_19093,N_18701,N_18569);
xnor U19094 (N_19094,N_18674,N_18708);
nand U19095 (N_19095,N_18693,N_18966);
nand U19096 (N_19096,N_18848,N_18825);
and U19097 (N_19097,N_18454,N_18641);
xnor U19098 (N_19098,N_18526,N_18938);
xnor U19099 (N_19099,N_18618,N_18915);
nor U19100 (N_19100,N_18890,N_18576);
and U19101 (N_19101,N_18013,N_18503);
nand U19102 (N_19102,N_18306,N_18893);
xnor U19103 (N_19103,N_18552,N_18899);
nor U19104 (N_19104,N_18416,N_18519);
nor U19105 (N_19105,N_18280,N_18368);
xor U19106 (N_19106,N_18509,N_18898);
xnor U19107 (N_19107,N_18402,N_18430);
xnor U19108 (N_19108,N_18671,N_18422);
xor U19109 (N_19109,N_18390,N_18974);
nor U19110 (N_19110,N_18408,N_18994);
xor U19111 (N_19111,N_18573,N_18624);
or U19112 (N_19112,N_18742,N_18315);
nor U19113 (N_19113,N_18342,N_18446);
and U19114 (N_19114,N_18989,N_18849);
or U19115 (N_19115,N_18648,N_18393);
and U19116 (N_19116,N_18991,N_18362);
or U19117 (N_19117,N_18590,N_18719);
and U19118 (N_19118,N_18025,N_18639);
xnor U19119 (N_19119,N_18194,N_18647);
xnor U19120 (N_19120,N_18772,N_18006);
and U19121 (N_19121,N_18489,N_18651);
or U19122 (N_19122,N_18001,N_18087);
and U19123 (N_19123,N_18696,N_18499);
or U19124 (N_19124,N_18225,N_18316);
xnor U19125 (N_19125,N_18578,N_18751);
xor U19126 (N_19126,N_18040,N_18927);
xor U19127 (N_19127,N_18514,N_18954);
and U19128 (N_19128,N_18513,N_18223);
or U19129 (N_19129,N_18395,N_18443);
or U19130 (N_19130,N_18895,N_18150);
xor U19131 (N_19131,N_18432,N_18873);
xnor U19132 (N_19132,N_18044,N_18119);
xor U19133 (N_19133,N_18337,N_18355);
nor U19134 (N_19134,N_18293,N_18135);
nand U19135 (N_19135,N_18756,N_18429);
nand U19136 (N_19136,N_18789,N_18323);
nand U19137 (N_19137,N_18604,N_18146);
nand U19138 (N_19138,N_18961,N_18384);
xor U19139 (N_19139,N_18271,N_18586);
xnor U19140 (N_19140,N_18407,N_18273);
nand U19141 (N_19141,N_18837,N_18038);
nor U19142 (N_19142,N_18066,N_18435);
xor U19143 (N_19143,N_18577,N_18433);
or U19144 (N_19144,N_18803,N_18188);
nor U19145 (N_19145,N_18344,N_18351);
xnor U19146 (N_19146,N_18191,N_18213);
xnor U19147 (N_19147,N_18440,N_18907);
nand U19148 (N_19148,N_18685,N_18340);
xnor U19149 (N_19149,N_18852,N_18243);
and U19150 (N_19150,N_18453,N_18735);
or U19151 (N_19151,N_18494,N_18152);
or U19152 (N_19152,N_18187,N_18339);
xnor U19153 (N_19153,N_18729,N_18531);
or U19154 (N_19154,N_18774,N_18208);
xnor U19155 (N_19155,N_18410,N_18237);
xnor U19156 (N_19156,N_18313,N_18380);
nand U19157 (N_19157,N_18654,N_18965);
and U19158 (N_19158,N_18667,N_18892);
nor U19159 (N_19159,N_18232,N_18960);
nand U19160 (N_19160,N_18944,N_18098);
xor U19161 (N_19161,N_18739,N_18413);
nand U19162 (N_19162,N_18062,N_18274);
and U19163 (N_19163,N_18036,N_18703);
nand U19164 (N_19164,N_18832,N_18836);
or U19165 (N_19165,N_18212,N_18151);
and U19166 (N_19166,N_18417,N_18112);
nor U19167 (N_19167,N_18227,N_18046);
and U19168 (N_19168,N_18951,N_18762);
and U19169 (N_19169,N_18356,N_18282);
or U19170 (N_19170,N_18377,N_18181);
nor U19171 (N_19171,N_18871,N_18963);
and U19172 (N_19172,N_18010,N_18567);
nand U19173 (N_19173,N_18196,N_18511);
and U19174 (N_19174,N_18634,N_18136);
or U19175 (N_19175,N_18782,N_18706);
or U19176 (N_19176,N_18660,N_18455);
and U19177 (N_19177,N_18496,N_18705);
and U19178 (N_19178,N_18847,N_18267);
or U19179 (N_19179,N_18790,N_18822);
or U19180 (N_19180,N_18487,N_18260);
and U19181 (N_19181,N_18952,N_18394);
nand U19182 (N_19182,N_18291,N_18240);
nor U19183 (N_19183,N_18277,N_18992);
or U19184 (N_19184,N_18366,N_18055);
nand U19185 (N_19185,N_18409,N_18838);
or U19186 (N_19186,N_18616,N_18217);
nand U19187 (N_19187,N_18490,N_18839);
xnor U19188 (N_19188,N_18656,N_18302);
nor U19189 (N_19189,N_18607,N_18653);
nand U19190 (N_19190,N_18357,N_18970);
nand U19191 (N_19191,N_18599,N_18828);
or U19192 (N_19192,N_18158,N_18878);
and U19193 (N_19193,N_18349,N_18285);
nand U19194 (N_19194,N_18470,N_18094);
nor U19195 (N_19195,N_18972,N_18124);
nand U19196 (N_19196,N_18688,N_18846);
or U19197 (N_19197,N_18724,N_18758);
or U19198 (N_19198,N_18909,N_18558);
and U19199 (N_19199,N_18610,N_18224);
nand U19200 (N_19200,N_18076,N_18185);
nand U19201 (N_19201,N_18981,N_18414);
and U19202 (N_19202,N_18773,N_18449);
and U19203 (N_19203,N_18765,N_18020);
nand U19204 (N_19204,N_18823,N_18600);
nand U19205 (N_19205,N_18457,N_18949);
and U19206 (N_19206,N_18426,N_18379);
nand U19207 (N_19207,N_18205,N_18170);
or U19208 (N_19208,N_18831,N_18920);
or U19209 (N_19209,N_18580,N_18370);
and U19210 (N_19210,N_18548,N_18817);
or U19211 (N_19211,N_18047,N_18882);
xnor U19212 (N_19212,N_18419,N_18437);
xor U19213 (N_19213,N_18508,N_18850);
xnor U19214 (N_19214,N_18163,N_18318);
nand U19215 (N_19215,N_18431,N_18943);
nor U19216 (N_19216,N_18396,N_18833);
nand U19217 (N_19217,N_18250,N_18620);
nand U19218 (N_19218,N_18445,N_18955);
and U19219 (N_19219,N_18206,N_18921);
xnor U19220 (N_19220,N_18234,N_18566);
xor U19221 (N_19221,N_18631,N_18870);
and U19222 (N_19222,N_18078,N_18934);
nor U19223 (N_19223,N_18014,N_18229);
nor U19224 (N_19224,N_18345,N_18348);
nor U19225 (N_19225,N_18866,N_18925);
and U19226 (N_19226,N_18630,N_18806);
xnor U19227 (N_19227,N_18308,N_18704);
xor U19228 (N_19228,N_18769,N_18721);
or U19229 (N_19229,N_18148,N_18809);
xor U19230 (N_19230,N_18144,N_18008);
and U19231 (N_19231,N_18155,N_18770);
xor U19232 (N_19232,N_18570,N_18325);
nor U19233 (N_19233,N_18476,N_18771);
nor U19234 (N_19234,N_18738,N_18039);
or U19235 (N_19235,N_18272,N_18195);
and U19236 (N_19236,N_18611,N_18602);
and U19237 (N_19237,N_18334,N_18262);
nand U19238 (N_19238,N_18045,N_18830);
nor U19239 (N_19239,N_18518,N_18710);
and U19240 (N_19240,N_18593,N_18574);
or U19241 (N_19241,N_18623,N_18310);
nor U19242 (N_19242,N_18301,N_18074);
and U19243 (N_19243,N_18711,N_18425);
and U19244 (N_19244,N_18424,N_18750);
nor U19245 (N_19245,N_18775,N_18193);
xnor U19246 (N_19246,N_18184,N_18143);
xor U19247 (N_19247,N_18412,N_18619);
and U19248 (N_19248,N_18126,N_18712);
nor U19249 (N_19249,N_18643,N_18640);
nor U19250 (N_19250,N_18421,N_18876);
nor U19251 (N_19251,N_18727,N_18652);
nand U19252 (N_19252,N_18507,N_18810);
xor U19253 (N_19253,N_18251,N_18929);
nor U19254 (N_19254,N_18510,N_18516);
nand U19255 (N_19255,N_18902,N_18473);
or U19256 (N_19256,N_18592,N_18065);
and U19257 (N_19257,N_18248,N_18687);
xnor U19258 (N_19258,N_18889,N_18060);
nor U19259 (N_19259,N_18857,N_18788);
xnor U19260 (N_19260,N_18057,N_18884);
and U19261 (N_19261,N_18754,N_18442);
and U19262 (N_19262,N_18474,N_18333);
or U19263 (N_19263,N_18099,N_18874);
xor U19264 (N_19264,N_18628,N_18495);
or U19265 (N_19265,N_18694,N_18560);
xnor U19266 (N_19266,N_18761,N_18713);
and U19267 (N_19267,N_18691,N_18103);
nand U19268 (N_19268,N_18936,N_18969);
xor U19269 (N_19269,N_18826,N_18764);
or U19270 (N_19270,N_18137,N_18595);
xor U19271 (N_19271,N_18988,N_18689);
or U19272 (N_19272,N_18629,N_18392);
nor U19273 (N_19273,N_18400,N_18858);
xor U19274 (N_19274,N_18975,N_18423);
xor U19275 (N_19275,N_18268,N_18197);
or U19276 (N_19276,N_18022,N_18451);
nor U19277 (N_19277,N_18079,N_18881);
or U19278 (N_19278,N_18075,N_18591);
xnor U19279 (N_19279,N_18284,N_18766);
and U19280 (N_19280,N_18117,N_18341);
nand U19281 (N_19281,N_18695,N_18028);
nand U19282 (N_19282,N_18805,N_18880);
or U19283 (N_19283,N_18814,N_18258);
and U19284 (N_19284,N_18732,N_18397);
or U19285 (N_19285,N_18319,N_18726);
nand U19286 (N_19286,N_18452,N_18886);
nand U19287 (N_19287,N_18785,N_18097);
and U19288 (N_19288,N_18447,N_18073);
and U19289 (N_19289,N_18253,N_18374);
and U19290 (N_19290,N_18791,N_18465);
nor U19291 (N_19291,N_18525,N_18024);
and U19292 (N_19292,N_18228,N_18061);
xnor U19293 (N_19293,N_18162,N_18448);
nand U19294 (N_19294,N_18562,N_18862);
nand U19295 (N_19295,N_18096,N_18798);
nand U19296 (N_19296,N_18905,N_18584);
and U19297 (N_19297,N_18130,N_18338);
or U19298 (N_19298,N_18053,N_18314);
xor U19299 (N_19299,N_18923,N_18655);
xnor U19300 (N_19300,N_18387,N_18249);
xnor U19301 (N_19301,N_18145,N_18501);
or U19302 (N_19302,N_18266,N_18515);
nor U19303 (N_19303,N_18588,N_18542);
xor U19304 (N_19304,N_18035,N_18608);
and U19305 (N_19305,N_18378,N_18298);
xnor U19306 (N_19306,N_18901,N_18347);
and U19307 (N_19307,N_18222,N_18867);
and U19308 (N_19308,N_18259,N_18976);
nor U19309 (N_19309,N_18138,N_18233);
nand U19310 (N_19310,N_18669,N_18009);
xor U19311 (N_19311,N_18252,N_18637);
nand U19312 (N_19312,N_18948,N_18219);
nand U19313 (N_19313,N_18612,N_18289);
and U19314 (N_19314,N_18064,N_18320);
or U19315 (N_19315,N_18479,N_18118);
xnor U19316 (N_19316,N_18156,N_18942);
nor U19317 (N_19317,N_18399,N_18322);
or U19318 (N_19318,N_18054,N_18202);
nor U19319 (N_19319,N_18161,N_18947);
and U19320 (N_19320,N_18799,N_18231);
xnor U19321 (N_19321,N_18481,N_18458);
xor U19322 (N_19322,N_18784,N_18459);
xnor U19323 (N_19323,N_18069,N_18572);
xor U19324 (N_19324,N_18031,N_18709);
nor U19325 (N_19325,N_18002,N_18418);
xor U19326 (N_19326,N_18995,N_18017);
nor U19327 (N_19327,N_18468,N_18800);
and U19328 (N_19328,N_18101,N_18614);
and U19329 (N_19329,N_18270,N_18967);
and U19330 (N_19330,N_18420,N_18080);
nand U19331 (N_19331,N_18030,N_18760);
and U19332 (N_19332,N_18911,N_18361);
and U19333 (N_19333,N_18186,N_18918);
and U19334 (N_19334,N_18937,N_18549);
nand U19335 (N_19335,N_18505,N_18786);
nor U19336 (N_19336,N_18546,N_18382);
xor U19337 (N_19337,N_18720,N_18110);
or U19338 (N_19338,N_18950,N_18568);
xnor U19339 (N_19339,N_18939,N_18835);
nor U19340 (N_19340,N_18070,N_18579);
or U19341 (N_19341,N_18149,N_18049);
nand U19342 (N_19342,N_18553,N_18968);
or U19343 (N_19343,N_18018,N_18131);
and U19344 (N_19344,N_18072,N_18700);
nand U19345 (N_19345,N_18467,N_18894);
xnor U19346 (N_19346,N_18658,N_18176);
or U19347 (N_19347,N_18946,N_18752);
and U19348 (N_19348,N_18042,N_18649);
nor U19349 (N_19349,N_18897,N_18841);
or U19350 (N_19350,N_18084,N_18613);
nand U19351 (N_19351,N_18757,N_18812);
and U19352 (N_19352,N_18535,N_18389);
and U19353 (N_19353,N_18294,N_18763);
or U19354 (N_19354,N_18559,N_18359);
and U19355 (N_19355,N_18617,N_18471);
or U19356 (N_19356,N_18003,N_18093);
nor U19357 (N_19357,N_18167,N_18300);
or U19358 (N_19358,N_18012,N_18168);
or U19359 (N_19359,N_18364,N_18083);
nor U19360 (N_19360,N_18904,N_18048);
nand U19361 (N_19361,N_18900,N_18041);
nand U19362 (N_19362,N_18331,N_18500);
and U19363 (N_19363,N_18215,N_18755);
and U19364 (N_19364,N_18565,N_18436);
xnor U19365 (N_19365,N_18089,N_18463);
nor U19366 (N_19366,N_18818,N_18957);
nand U19367 (N_19367,N_18635,N_18207);
and U19368 (N_19368,N_18438,N_18597);
and U19369 (N_19369,N_18385,N_18748);
nor U19370 (N_19370,N_18353,N_18241);
or U19371 (N_19371,N_18256,N_18716);
nand U19372 (N_19372,N_18472,N_18842);
xnor U19373 (N_19373,N_18722,N_18497);
or U19374 (N_19374,N_18004,N_18204);
and U19375 (N_19375,N_18797,N_18157);
or U19376 (N_19376,N_18563,N_18113);
nand U19377 (N_19377,N_18914,N_18615);
or U19378 (N_19378,N_18645,N_18863);
nor U19379 (N_19379,N_18464,N_18492);
or U19380 (N_19380,N_18768,N_18498);
and U19381 (N_19381,N_18594,N_18160);
nand U19382 (N_19382,N_18677,N_18132);
xor U19383 (N_19383,N_18530,N_18032);
or U19384 (N_19384,N_18522,N_18159);
xnor U19385 (N_19385,N_18281,N_18840);
xor U19386 (N_19386,N_18122,N_18877);
nand U19387 (N_19387,N_18978,N_18128);
nand U19388 (N_19388,N_18690,N_18461);
nand U19389 (N_19389,N_18283,N_18190);
xnor U19390 (N_19390,N_18622,N_18744);
or U19391 (N_19391,N_18226,N_18545);
xnor U19392 (N_19392,N_18749,N_18891);
or U19393 (N_19393,N_18127,N_18887);
nor U19394 (N_19394,N_18238,N_18111);
nor U19395 (N_19395,N_18537,N_18883);
or U19396 (N_19396,N_18105,N_18855);
or U19397 (N_19397,N_18295,N_18529);
and U19398 (N_19398,N_18106,N_18154);
xnor U19399 (N_19399,N_18990,N_18051);
xor U19400 (N_19400,N_18125,N_18854);
or U19401 (N_19401,N_18005,N_18214);
nor U19402 (N_19402,N_18104,N_18912);
nor U19403 (N_19403,N_18913,N_18372);
nand U19404 (N_19404,N_18781,N_18140);
and U19405 (N_19405,N_18200,N_18255);
nand U19406 (N_19406,N_18056,N_18007);
and U19407 (N_19407,N_18746,N_18261);
xor U19408 (N_19408,N_18403,N_18092);
or U19409 (N_19409,N_18411,N_18987);
or U19410 (N_19410,N_18807,N_18365);
xor U19411 (N_19411,N_18466,N_18536);
xnor U19412 (N_19412,N_18802,N_18292);
nor U19413 (N_19413,N_18587,N_18139);
and U19414 (N_19414,N_18779,N_18728);
nor U19415 (N_19415,N_18199,N_18332);
nand U19416 (N_19416,N_18077,N_18606);
xor U19417 (N_19417,N_18000,N_18406);
and U19418 (N_19418,N_18450,N_18956);
or U19419 (N_19419,N_18375,N_18702);
or U19420 (N_19420,N_18391,N_18714);
xnor U19421 (N_19421,N_18675,N_18636);
nor U19422 (N_19422,N_18598,N_18626);
nand U19423 (N_19423,N_18583,N_18371);
nor U19424 (N_19424,N_18102,N_18304);
and U19425 (N_19425,N_18328,N_18230);
nor U19426 (N_19426,N_18996,N_18153);
nor U19427 (N_19427,N_18979,N_18953);
and U19428 (N_19428,N_18236,N_18182);
nor U19429 (N_19429,N_18917,N_18930);
nand U19430 (N_19430,N_18556,N_18665);
nand U19431 (N_19431,N_18367,N_18043);
nor U19432 (N_19432,N_18090,N_18940);
nor U19433 (N_19433,N_18603,N_18373);
and U19434 (N_19434,N_18174,N_18352);
or U19435 (N_19435,N_18707,N_18795);
xor U19436 (N_19436,N_18100,N_18169);
and U19437 (N_19437,N_18299,N_18678);
or U19438 (N_19438,N_18235,N_18109);
nand U19439 (N_19439,N_18346,N_18475);
nor U19440 (N_19440,N_18203,N_18859);
xor U19441 (N_19441,N_18068,N_18123);
and U19442 (N_19442,N_18239,N_18269);
or U19443 (N_19443,N_18997,N_18183);
nand U19444 (N_19444,N_18792,N_18147);
nor U19445 (N_19445,N_18063,N_18360);
nor U19446 (N_19446,N_18082,N_18512);
nand U19447 (N_19447,N_18885,N_18037);
and U19448 (N_19448,N_18305,N_18980);
or U19449 (N_19449,N_18896,N_18192);
or U19450 (N_19450,N_18999,N_18844);
or U19451 (N_19451,N_18650,N_18924);
and U19452 (N_19452,N_18034,N_18129);
xnor U19453 (N_19453,N_18523,N_18834);
nor U19454 (N_19454,N_18324,N_18564);
nand U19455 (N_19455,N_18663,N_18477);
xnor U19456 (N_19456,N_18699,N_18540);
nand U19457 (N_19457,N_18793,N_18264);
or U19458 (N_19458,N_18561,N_18386);
xor U19459 (N_19459,N_18484,N_18297);
or U19460 (N_19460,N_18554,N_18180);
nand U19461 (N_19461,N_18682,N_18528);
xnor U19462 (N_19462,N_18734,N_18986);
nand U19463 (N_19463,N_18029,N_18697);
xnor U19464 (N_19464,N_18290,N_18601);
nor U19465 (N_19465,N_18815,N_18851);
xnor U19466 (N_19466,N_18715,N_18973);
xor U19467 (N_19467,N_18033,N_18133);
nand U19468 (N_19468,N_18777,N_18659);
or U19469 (N_19469,N_18307,N_18172);
or U19470 (N_19470,N_18071,N_18246);
nor U19471 (N_19471,N_18086,N_18646);
xnor U19472 (N_19472,N_18059,N_18718);
or U19473 (N_19473,N_18491,N_18585);
nand U19474 (N_19474,N_18723,N_18327);
xnor U19475 (N_19475,N_18166,N_18868);
nand U19476 (N_19476,N_18405,N_18321);
xnor U19477 (N_19477,N_18330,N_18984);
nand U19478 (N_19478,N_18095,N_18275);
xor U19479 (N_19479,N_18171,N_18469);
nor U19480 (N_19480,N_18401,N_18015);
nand U19481 (N_19481,N_18605,N_18276);
xnor U19482 (N_19482,N_18287,N_18683);
or U19483 (N_19483,N_18052,N_18263);
nor U19484 (N_19484,N_18173,N_18672);
nand U19485 (N_19485,N_18335,N_18543);
nand U19486 (N_19486,N_18220,N_18278);
xor U19487 (N_19487,N_18922,N_18686);
or U19488 (N_19488,N_18108,N_18369);
nand U19489 (N_19489,N_18993,N_18928);
nor U19490 (N_19490,N_18532,N_18541);
xnor U19491 (N_19491,N_18959,N_18114);
nor U19492 (N_19492,N_18982,N_18107);
nand U19493 (N_19493,N_18326,N_18869);
nor U19494 (N_19494,N_18354,N_18717);
and U19495 (N_19495,N_18888,N_18935);
and U19496 (N_19496,N_18958,N_18550);
or U19497 (N_19497,N_18067,N_18551);
and U19498 (N_19498,N_18875,N_18502);
and U19499 (N_19499,N_18865,N_18218);
nand U19500 (N_19500,N_18171,N_18366);
or U19501 (N_19501,N_18094,N_18201);
nand U19502 (N_19502,N_18827,N_18993);
xor U19503 (N_19503,N_18623,N_18366);
xnor U19504 (N_19504,N_18305,N_18287);
nor U19505 (N_19505,N_18352,N_18658);
xnor U19506 (N_19506,N_18284,N_18447);
nor U19507 (N_19507,N_18357,N_18058);
xnor U19508 (N_19508,N_18122,N_18074);
xnor U19509 (N_19509,N_18127,N_18423);
or U19510 (N_19510,N_18421,N_18488);
and U19511 (N_19511,N_18908,N_18938);
xnor U19512 (N_19512,N_18973,N_18884);
nor U19513 (N_19513,N_18114,N_18196);
and U19514 (N_19514,N_18557,N_18115);
or U19515 (N_19515,N_18145,N_18143);
nand U19516 (N_19516,N_18859,N_18073);
or U19517 (N_19517,N_18418,N_18951);
nor U19518 (N_19518,N_18073,N_18264);
nand U19519 (N_19519,N_18213,N_18470);
and U19520 (N_19520,N_18621,N_18272);
or U19521 (N_19521,N_18434,N_18619);
and U19522 (N_19522,N_18617,N_18558);
nand U19523 (N_19523,N_18521,N_18041);
xnor U19524 (N_19524,N_18516,N_18609);
or U19525 (N_19525,N_18768,N_18177);
or U19526 (N_19526,N_18788,N_18664);
or U19527 (N_19527,N_18856,N_18852);
or U19528 (N_19528,N_18846,N_18141);
xor U19529 (N_19529,N_18060,N_18389);
xnor U19530 (N_19530,N_18498,N_18516);
nor U19531 (N_19531,N_18719,N_18002);
or U19532 (N_19532,N_18383,N_18585);
xor U19533 (N_19533,N_18277,N_18212);
and U19534 (N_19534,N_18845,N_18362);
xor U19535 (N_19535,N_18607,N_18497);
or U19536 (N_19536,N_18652,N_18442);
and U19537 (N_19537,N_18777,N_18448);
nand U19538 (N_19538,N_18826,N_18223);
xnor U19539 (N_19539,N_18450,N_18908);
nand U19540 (N_19540,N_18817,N_18704);
or U19541 (N_19541,N_18376,N_18939);
and U19542 (N_19542,N_18773,N_18795);
nand U19543 (N_19543,N_18456,N_18137);
nor U19544 (N_19544,N_18072,N_18770);
or U19545 (N_19545,N_18925,N_18655);
nand U19546 (N_19546,N_18363,N_18948);
and U19547 (N_19547,N_18771,N_18001);
and U19548 (N_19548,N_18719,N_18827);
nand U19549 (N_19549,N_18412,N_18840);
nand U19550 (N_19550,N_18016,N_18965);
and U19551 (N_19551,N_18665,N_18969);
nor U19552 (N_19552,N_18357,N_18225);
and U19553 (N_19553,N_18650,N_18510);
nand U19554 (N_19554,N_18545,N_18369);
xnor U19555 (N_19555,N_18293,N_18048);
nor U19556 (N_19556,N_18928,N_18522);
or U19557 (N_19557,N_18250,N_18464);
xor U19558 (N_19558,N_18330,N_18531);
xor U19559 (N_19559,N_18372,N_18359);
nand U19560 (N_19560,N_18892,N_18975);
and U19561 (N_19561,N_18395,N_18125);
nand U19562 (N_19562,N_18209,N_18899);
xor U19563 (N_19563,N_18595,N_18489);
xnor U19564 (N_19564,N_18485,N_18304);
or U19565 (N_19565,N_18178,N_18550);
nor U19566 (N_19566,N_18548,N_18607);
nand U19567 (N_19567,N_18470,N_18961);
or U19568 (N_19568,N_18663,N_18099);
nand U19569 (N_19569,N_18438,N_18758);
nand U19570 (N_19570,N_18879,N_18843);
nor U19571 (N_19571,N_18228,N_18767);
or U19572 (N_19572,N_18225,N_18852);
and U19573 (N_19573,N_18484,N_18797);
nand U19574 (N_19574,N_18531,N_18204);
and U19575 (N_19575,N_18744,N_18505);
and U19576 (N_19576,N_18363,N_18828);
nor U19577 (N_19577,N_18951,N_18459);
nor U19578 (N_19578,N_18321,N_18427);
nand U19579 (N_19579,N_18450,N_18134);
or U19580 (N_19580,N_18915,N_18864);
nor U19581 (N_19581,N_18410,N_18665);
nor U19582 (N_19582,N_18679,N_18536);
nor U19583 (N_19583,N_18722,N_18994);
nand U19584 (N_19584,N_18867,N_18513);
nor U19585 (N_19585,N_18087,N_18310);
and U19586 (N_19586,N_18095,N_18361);
or U19587 (N_19587,N_18674,N_18201);
or U19588 (N_19588,N_18513,N_18865);
or U19589 (N_19589,N_18517,N_18429);
nand U19590 (N_19590,N_18277,N_18432);
and U19591 (N_19591,N_18882,N_18117);
xor U19592 (N_19592,N_18857,N_18354);
nand U19593 (N_19593,N_18835,N_18096);
nand U19594 (N_19594,N_18247,N_18426);
nand U19595 (N_19595,N_18768,N_18132);
or U19596 (N_19596,N_18296,N_18622);
nor U19597 (N_19597,N_18764,N_18368);
nor U19598 (N_19598,N_18279,N_18129);
and U19599 (N_19599,N_18751,N_18869);
and U19600 (N_19600,N_18509,N_18386);
xnor U19601 (N_19601,N_18538,N_18873);
or U19602 (N_19602,N_18954,N_18563);
or U19603 (N_19603,N_18795,N_18233);
nor U19604 (N_19604,N_18551,N_18718);
or U19605 (N_19605,N_18501,N_18813);
or U19606 (N_19606,N_18854,N_18981);
and U19607 (N_19607,N_18254,N_18298);
or U19608 (N_19608,N_18758,N_18006);
nor U19609 (N_19609,N_18632,N_18855);
xor U19610 (N_19610,N_18991,N_18313);
nor U19611 (N_19611,N_18145,N_18839);
and U19612 (N_19612,N_18297,N_18609);
nor U19613 (N_19613,N_18194,N_18161);
and U19614 (N_19614,N_18483,N_18045);
nor U19615 (N_19615,N_18720,N_18448);
nand U19616 (N_19616,N_18315,N_18014);
and U19617 (N_19617,N_18541,N_18286);
and U19618 (N_19618,N_18894,N_18300);
xnor U19619 (N_19619,N_18614,N_18277);
or U19620 (N_19620,N_18334,N_18501);
xor U19621 (N_19621,N_18369,N_18121);
nor U19622 (N_19622,N_18472,N_18850);
nand U19623 (N_19623,N_18933,N_18773);
nor U19624 (N_19624,N_18945,N_18794);
nor U19625 (N_19625,N_18883,N_18060);
or U19626 (N_19626,N_18962,N_18837);
nor U19627 (N_19627,N_18035,N_18383);
xnor U19628 (N_19628,N_18873,N_18264);
or U19629 (N_19629,N_18843,N_18807);
nor U19630 (N_19630,N_18560,N_18190);
nor U19631 (N_19631,N_18239,N_18804);
or U19632 (N_19632,N_18394,N_18226);
and U19633 (N_19633,N_18388,N_18787);
and U19634 (N_19634,N_18238,N_18949);
nor U19635 (N_19635,N_18739,N_18076);
or U19636 (N_19636,N_18279,N_18708);
xor U19637 (N_19637,N_18062,N_18348);
or U19638 (N_19638,N_18932,N_18741);
and U19639 (N_19639,N_18522,N_18717);
or U19640 (N_19640,N_18978,N_18971);
xor U19641 (N_19641,N_18689,N_18418);
xor U19642 (N_19642,N_18741,N_18671);
and U19643 (N_19643,N_18002,N_18084);
nand U19644 (N_19644,N_18628,N_18345);
nor U19645 (N_19645,N_18639,N_18398);
or U19646 (N_19646,N_18603,N_18278);
nand U19647 (N_19647,N_18266,N_18916);
xor U19648 (N_19648,N_18044,N_18221);
nor U19649 (N_19649,N_18916,N_18672);
xor U19650 (N_19650,N_18833,N_18295);
nand U19651 (N_19651,N_18057,N_18162);
xnor U19652 (N_19652,N_18621,N_18509);
nand U19653 (N_19653,N_18936,N_18025);
nor U19654 (N_19654,N_18484,N_18547);
or U19655 (N_19655,N_18457,N_18878);
xor U19656 (N_19656,N_18585,N_18957);
or U19657 (N_19657,N_18706,N_18209);
and U19658 (N_19658,N_18918,N_18484);
nand U19659 (N_19659,N_18686,N_18213);
nand U19660 (N_19660,N_18253,N_18680);
nand U19661 (N_19661,N_18570,N_18660);
xnor U19662 (N_19662,N_18491,N_18395);
nand U19663 (N_19663,N_18029,N_18159);
or U19664 (N_19664,N_18841,N_18609);
xor U19665 (N_19665,N_18203,N_18496);
nand U19666 (N_19666,N_18930,N_18747);
or U19667 (N_19667,N_18403,N_18580);
and U19668 (N_19668,N_18775,N_18365);
nand U19669 (N_19669,N_18147,N_18408);
nor U19670 (N_19670,N_18735,N_18042);
or U19671 (N_19671,N_18002,N_18897);
nand U19672 (N_19672,N_18295,N_18654);
xor U19673 (N_19673,N_18033,N_18793);
xor U19674 (N_19674,N_18633,N_18913);
nor U19675 (N_19675,N_18248,N_18359);
nand U19676 (N_19676,N_18098,N_18471);
and U19677 (N_19677,N_18503,N_18765);
nand U19678 (N_19678,N_18284,N_18850);
nand U19679 (N_19679,N_18842,N_18962);
and U19680 (N_19680,N_18341,N_18026);
and U19681 (N_19681,N_18980,N_18920);
xnor U19682 (N_19682,N_18115,N_18446);
nor U19683 (N_19683,N_18587,N_18704);
nor U19684 (N_19684,N_18573,N_18306);
nor U19685 (N_19685,N_18407,N_18507);
nand U19686 (N_19686,N_18353,N_18698);
xor U19687 (N_19687,N_18024,N_18741);
or U19688 (N_19688,N_18836,N_18192);
nor U19689 (N_19689,N_18923,N_18769);
or U19690 (N_19690,N_18747,N_18759);
nand U19691 (N_19691,N_18789,N_18718);
xor U19692 (N_19692,N_18880,N_18091);
or U19693 (N_19693,N_18842,N_18086);
nor U19694 (N_19694,N_18706,N_18211);
nor U19695 (N_19695,N_18182,N_18072);
xnor U19696 (N_19696,N_18705,N_18189);
nand U19697 (N_19697,N_18708,N_18705);
xnor U19698 (N_19698,N_18246,N_18988);
and U19699 (N_19699,N_18057,N_18487);
xor U19700 (N_19700,N_18756,N_18821);
or U19701 (N_19701,N_18229,N_18143);
xnor U19702 (N_19702,N_18033,N_18045);
nand U19703 (N_19703,N_18423,N_18243);
nor U19704 (N_19704,N_18241,N_18505);
nor U19705 (N_19705,N_18524,N_18871);
nor U19706 (N_19706,N_18083,N_18187);
or U19707 (N_19707,N_18930,N_18811);
or U19708 (N_19708,N_18854,N_18489);
or U19709 (N_19709,N_18571,N_18667);
or U19710 (N_19710,N_18480,N_18445);
and U19711 (N_19711,N_18811,N_18911);
or U19712 (N_19712,N_18837,N_18926);
xor U19713 (N_19713,N_18359,N_18883);
nand U19714 (N_19714,N_18517,N_18622);
and U19715 (N_19715,N_18265,N_18762);
nand U19716 (N_19716,N_18626,N_18660);
nor U19717 (N_19717,N_18276,N_18131);
xor U19718 (N_19718,N_18351,N_18128);
nor U19719 (N_19719,N_18584,N_18274);
nor U19720 (N_19720,N_18365,N_18461);
nor U19721 (N_19721,N_18114,N_18038);
or U19722 (N_19722,N_18848,N_18574);
nand U19723 (N_19723,N_18436,N_18574);
nor U19724 (N_19724,N_18152,N_18538);
xnor U19725 (N_19725,N_18839,N_18089);
nand U19726 (N_19726,N_18643,N_18832);
and U19727 (N_19727,N_18081,N_18065);
or U19728 (N_19728,N_18248,N_18188);
nor U19729 (N_19729,N_18283,N_18390);
and U19730 (N_19730,N_18056,N_18390);
nor U19731 (N_19731,N_18392,N_18636);
nand U19732 (N_19732,N_18087,N_18995);
and U19733 (N_19733,N_18044,N_18849);
and U19734 (N_19734,N_18008,N_18670);
or U19735 (N_19735,N_18165,N_18193);
xor U19736 (N_19736,N_18182,N_18501);
and U19737 (N_19737,N_18884,N_18491);
and U19738 (N_19738,N_18094,N_18285);
xnor U19739 (N_19739,N_18067,N_18700);
and U19740 (N_19740,N_18892,N_18515);
xnor U19741 (N_19741,N_18988,N_18623);
xnor U19742 (N_19742,N_18123,N_18031);
nand U19743 (N_19743,N_18257,N_18150);
xor U19744 (N_19744,N_18689,N_18516);
nor U19745 (N_19745,N_18031,N_18647);
nor U19746 (N_19746,N_18768,N_18007);
xnor U19747 (N_19747,N_18773,N_18511);
nor U19748 (N_19748,N_18055,N_18192);
and U19749 (N_19749,N_18325,N_18143);
or U19750 (N_19750,N_18027,N_18460);
xnor U19751 (N_19751,N_18211,N_18584);
nor U19752 (N_19752,N_18988,N_18942);
or U19753 (N_19753,N_18621,N_18584);
nand U19754 (N_19754,N_18201,N_18163);
nor U19755 (N_19755,N_18174,N_18302);
and U19756 (N_19756,N_18539,N_18253);
or U19757 (N_19757,N_18944,N_18341);
and U19758 (N_19758,N_18275,N_18948);
and U19759 (N_19759,N_18289,N_18199);
nand U19760 (N_19760,N_18218,N_18313);
nor U19761 (N_19761,N_18588,N_18285);
nor U19762 (N_19762,N_18778,N_18367);
and U19763 (N_19763,N_18820,N_18631);
nor U19764 (N_19764,N_18487,N_18504);
nand U19765 (N_19765,N_18030,N_18648);
xnor U19766 (N_19766,N_18496,N_18703);
and U19767 (N_19767,N_18455,N_18092);
or U19768 (N_19768,N_18618,N_18365);
xor U19769 (N_19769,N_18158,N_18811);
xnor U19770 (N_19770,N_18615,N_18598);
nor U19771 (N_19771,N_18587,N_18685);
nor U19772 (N_19772,N_18489,N_18120);
and U19773 (N_19773,N_18216,N_18737);
nor U19774 (N_19774,N_18364,N_18436);
nor U19775 (N_19775,N_18846,N_18801);
nand U19776 (N_19776,N_18420,N_18360);
xor U19777 (N_19777,N_18080,N_18561);
nand U19778 (N_19778,N_18349,N_18034);
nand U19779 (N_19779,N_18653,N_18610);
or U19780 (N_19780,N_18840,N_18885);
xnor U19781 (N_19781,N_18862,N_18522);
nand U19782 (N_19782,N_18414,N_18182);
or U19783 (N_19783,N_18796,N_18369);
or U19784 (N_19784,N_18039,N_18467);
and U19785 (N_19785,N_18847,N_18404);
nor U19786 (N_19786,N_18277,N_18708);
or U19787 (N_19787,N_18223,N_18884);
nand U19788 (N_19788,N_18783,N_18528);
and U19789 (N_19789,N_18639,N_18948);
nor U19790 (N_19790,N_18830,N_18052);
nand U19791 (N_19791,N_18134,N_18891);
or U19792 (N_19792,N_18363,N_18634);
and U19793 (N_19793,N_18011,N_18596);
and U19794 (N_19794,N_18801,N_18475);
xor U19795 (N_19795,N_18749,N_18775);
xor U19796 (N_19796,N_18268,N_18362);
and U19797 (N_19797,N_18357,N_18893);
xor U19798 (N_19798,N_18146,N_18549);
or U19799 (N_19799,N_18892,N_18104);
xnor U19800 (N_19800,N_18234,N_18027);
or U19801 (N_19801,N_18037,N_18657);
nor U19802 (N_19802,N_18079,N_18239);
and U19803 (N_19803,N_18080,N_18678);
nor U19804 (N_19804,N_18319,N_18423);
or U19805 (N_19805,N_18577,N_18395);
or U19806 (N_19806,N_18895,N_18434);
nor U19807 (N_19807,N_18147,N_18523);
nor U19808 (N_19808,N_18625,N_18623);
xor U19809 (N_19809,N_18648,N_18731);
or U19810 (N_19810,N_18636,N_18275);
or U19811 (N_19811,N_18907,N_18811);
or U19812 (N_19812,N_18197,N_18831);
or U19813 (N_19813,N_18750,N_18956);
xnor U19814 (N_19814,N_18933,N_18697);
and U19815 (N_19815,N_18315,N_18413);
or U19816 (N_19816,N_18301,N_18482);
or U19817 (N_19817,N_18193,N_18872);
or U19818 (N_19818,N_18388,N_18488);
nand U19819 (N_19819,N_18795,N_18619);
and U19820 (N_19820,N_18828,N_18744);
nand U19821 (N_19821,N_18715,N_18853);
or U19822 (N_19822,N_18248,N_18733);
or U19823 (N_19823,N_18447,N_18260);
nand U19824 (N_19824,N_18345,N_18263);
or U19825 (N_19825,N_18203,N_18865);
nor U19826 (N_19826,N_18959,N_18262);
xor U19827 (N_19827,N_18392,N_18046);
or U19828 (N_19828,N_18886,N_18430);
xnor U19829 (N_19829,N_18433,N_18853);
or U19830 (N_19830,N_18077,N_18336);
nor U19831 (N_19831,N_18962,N_18443);
xnor U19832 (N_19832,N_18775,N_18133);
nand U19833 (N_19833,N_18148,N_18992);
xor U19834 (N_19834,N_18464,N_18689);
xnor U19835 (N_19835,N_18753,N_18326);
nor U19836 (N_19836,N_18012,N_18200);
nand U19837 (N_19837,N_18001,N_18307);
xor U19838 (N_19838,N_18642,N_18632);
nor U19839 (N_19839,N_18988,N_18237);
nor U19840 (N_19840,N_18279,N_18480);
nand U19841 (N_19841,N_18439,N_18782);
nand U19842 (N_19842,N_18581,N_18081);
xnor U19843 (N_19843,N_18640,N_18481);
xnor U19844 (N_19844,N_18423,N_18934);
nor U19845 (N_19845,N_18110,N_18326);
nor U19846 (N_19846,N_18320,N_18889);
nor U19847 (N_19847,N_18875,N_18244);
nand U19848 (N_19848,N_18284,N_18760);
xnor U19849 (N_19849,N_18741,N_18182);
and U19850 (N_19850,N_18856,N_18793);
nor U19851 (N_19851,N_18520,N_18922);
nor U19852 (N_19852,N_18669,N_18841);
xnor U19853 (N_19853,N_18034,N_18384);
nor U19854 (N_19854,N_18535,N_18725);
nand U19855 (N_19855,N_18204,N_18746);
nand U19856 (N_19856,N_18848,N_18663);
xnor U19857 (N_19857,N_18503,N_18816);
and U19858 (N_19858,N_18104,N_18775);
nand U19859 (N_19859,N_18967,N_18307);
and U19860 (N_19860,N_18148,N_18447);
xnor U19861 (N_19861,N_18062,N_18387);
and U19862 (N_19862,N_18269,N_18326);
and U19863 (N_19863,N_18209,N_18186);
nor U19864 (N_19864,N_18371,N_18170);
nand U19865 (N_19865,N_18265,N_18330);
or U19866 (N_19866,N_18896,N_18219);
nand U19867 (N_19867,N_18833,N_18182);
xnor U19868 (N_19868,N_18021,N_18007);
xor U19869 (N_19869,N_18714,N_18395);
nand U19870 (N_19870,N_18918,N_18564);
and U19871 (N_19871,N_18174,N_18808);
and U19872 (N_19872,N_18070,N_18153);
and U19873 (N_19873,N_18598,N_18034);
nor U19874 (N_19874,N_18509,N_18212);
or U19875 (N_19875,N_18302,N_18487);
xnor U19876 (N_19876,N_18667,N_18723);
or U19877 (N_19877,N_18783,N_18385);
and U19878 (N_19878,N_18055,N_18853);
or U19879 (N_19879,N_18011,N_18237);
nor U19880 (N_19880,N_18541,N_18949);
nor U19881 (N_19881,N_18534,N_18069);
and U19882 (N_19882,N_18019,N_18273);
and U19883 (N_19883,N_18620,N_18155);
and U19884 (N_19884,N_18287,N_18708);
or U19885 (N_19885,N_18053,N_18018);
nor U19886 (N_19886,N_18934,N_18960);
xor U19887 (N_19887,N_18175,N_18385);
xnor U19888 (N_19888,N_18808,N_18596);
xor U19889 (N_19889,N_18823,N_18129);
nand U19890 (N_19890,N_18259,N_18333);
nand U19891 (N_19891,N_18211,N_18726);
nand U19892 (N_19892,N_18423,N_18673);
nand U19893 (N_19893,N_18485,N_18077);
xnor U19894 (N_19894,N_18763,N_18050);
xor U19895 (N_19895,N_18809,N_18175);
and U19896 (N_19896,N_18463,N_18231);
or U19897 (N_19897,N_18114,N_18968);
or U19898 (N_19898,N_18315,N_18615);
or U19899 (N_19899,N_18606,N_18036);
or U19900 (N_19900,N_18799,N_18181);
and U19901 (N_19901,N_18104,N_18895);
nor U19902 (N_19902,N_18452,N_18792);
or U19903 (N_19903,N_18035,N_18909);
and U19904 (N_19904,N_18168,N_18422);
nor U19905 (N_19905,N_18991,N_18469);
and U19906 (N_19906,N_18649,N_18290);
nand U19907 (N_19907,N_18327,N_18633);
or U19908 (N_19908,N_18757,N_18298);
xor U19909 (N_19909,N_18027,N_18570);
or U19910 (N_19910,N_18701,N_18899);
nor U19911 (N_19911,N_18982,N_18786);
nor U19912 (N_19912,N_18683,N_18351);
xor U19913 (N_19913,N_18859,N_18173);
nand U19914 (N_19914,N_18005,N_18746);
nand U19915 (N_19915,N_18656,N_18983);
xnor U19916 (N_19916,N_18350,N_18777);
xor U19917 (N_19917,N_18936,N_18637);
nand U19918 (N_19918,N_18798,N_18642);
nor U19919 (N_19919,N_18019,N_18481);
xnor U19920 (N_19920,N_18916,N_18189);
or U19921 (N_19921,N_18136,N_18250);
xor U19922 (N_19922,N_18065,N_18797);
and U19923 (N_19923,N_18124,N_18786);
nand U19924 (N_19924,N_18414,N_18796);
and U19925 (N_19925,N_18539,N_18004);
and U19926 (N_19926,N_18569,N_18660);
nand U19927 (N_19927,N_18629,N_18620);
or U19928 (N_19928,N_18603,N_18907);
nand U19929 (N_19929,N_18085,N_18863);
and U19930 (N_19930,N_18036,N_18946);
xor U19931 (N_19931,N_18191,N_18852);
nand U19932 (N_19932,N_18502,N_18658);
or U19933 (N_19933,N_18972,N_18294);
nand U19934 (N_19934,N_18784,N_18750);
nor U19935 (N_19935,N_18747,N_18306);
xnor U19936 (N_19936,N_18923,N_18320);
xnor U19937 (N_19937,N_18348,N_18829);
and U19938 (N_19938,N_18912,N_18481);
xnor U19939 (N_19939,N_18780,N_18267);
xnor U19940 (N_19940,N_18309,N_18462);
xor U19941 (N_19941,N_18099,N_18462);
nand U19942 (N_19942,N_18026,N_18320);
nor U19943 (N_19943,N_18715,N_18271);
nor U19944 (N_19944,N_18442,N_18445);
nor U19945 (N_19945,N_18175,N_18304);
nand U19946 (N_19946,N_18051,N_18432);
nor U19947 (N_19947,N_18937,N_18324);
and U19948 (N_19948,N_18562,N_18928);
or U19949 (N_19949,N_18206,N_18048);
nor U19950 (N_19950,N_18154,N_18350);
nor U19951 (N_19951,N_18559,N_18991);
and U19952 (N_19952,N_18649,N_18208);
or U19953 (N_19953,N_18290,N_18789);
nand U19954 (N_19954,N_18374,N_18533);
or U19955 (N_19955,N_18848,N_18512);
and U19956 (N_19956,N_18449,N_18489);
nand U19957 (N_19957,N_18441,N_18150);
nor U19958 (N_19958,N_18724,N_18404);
nor U19959 (N_19959,N_18030,N_18045);
and U19960 (N_19960,N_18851,N_18025);
or U19961 (N_19961,N_18513,N_18551);
and U19962 (N_19962,N_18519,N_18396);
or U19963 (N_19963,N_18799,N_18443);
nor U19964 (N_19964,N_18753,N_18339);
xnor U19965 (N_19965,N_18926,N_18600);
or U19966 (N_19966,N_18837,N_18587);
and U19967 (N_19967,N_18150,N_18910);
xor U19968 (N_19968,N_18319,N_18897);
xnor U19969 (N_19969,N_18901,N_18554);
and U19970 (N_19970,N_18888,N_18917);
or U19971 (N_19971,N_18856,N_18036);
and U19972 (N_19972,N_18554,N_18804);
nand U19973 (N_19973,N_18333,N_18298);
nor U19974 (N_19974,N_18510,N_18697);
and U19975 (N_19975,N_18768,N_18764);
nand U19976 (N_19976,N_18990,N_18368);
and U19977 (N_19977,N_18657,N_18805);
xnor U19978 (N_19978,N_18195,N_18990);
or U19979 (N_19979,N_18328,N_18249);
xnor U19980 (N_19980,N_18714,N_18656);
xnor U19981 (N_19981,N_18657,N_18447);
nand U19982 (N_19982,N_18893,N_18197);
and U19983 (N_19983,N_18736,N_18491);
or U19984 (N_19984,N_18239,N_18999);
or U19985 (N_19985,N_18613,N_18816);
xor U19986 (N_19986,N_18371,N_18878);
or U19987 (N_19987,N_18806,N_18736);
or U19988 (N_19988,N_18336,N_18074);
nor U19989 (N_19989,N_18007,N_18539);
xor U19990 (N_19990,N_18092,N_18322);
and U19991 (N_19991,N_18541,N_18897);
and U19992 (N_19992,N_18228,N_18324);
xor U19993 (N_19993,N_18560,N_18231);
xnor U19994 (N_19994,N_18533,N_18279);
nor U19995 (N_19995,N_18820,N_18134);
nor U19996 (N_19996,N_18069,N_18145);
xor U19997 (N_19997,N_18035,N_18978);
and U19998 (N_19998,N_18144,N_18681);
and U19999 (N_19999,N_18669,N_18811);
nand U20000 (N_20000,N_19945,N_19468);
or U20001 (N_20001,N_19132,N_19479);
nor U20002 (N_20002,N_19183,N_19587);
or U20003 (N_20003,N_19210,N_19403);
xor U20004 (N_20004,N_19886,N_19645);
nor U20005 (N_20005,N_19292,N_19834);
xor U20006 (N_20006,N_19955,N_19541);
nand U20007 (N_20007,N_19111,N_19303);
nor U20008 (N_20008,N_19428,N_19972);
xnor U20009 (N_20009,N_19413,N_19340);
nor U20010 (N_20010,N_19768,N_19685);
or U20011 (N_20011,N_19454,N_19996);
nor U20012 (N_20012,N_19257,N_19734);
or U20013 (N_20013,N_19166,N_19534);
nand U20014 (N_20014,N_19379,N_19982);
xor U20015 (N_20015,N_19284,N_19633);
or U20016 (N_20016,N_19854,N_19044);
nand U20017 (N_20017,N_19953,N_19372);
or U20018 (N_20018,N_19314,N_19163);
xor U20019 (N_20019,N_19349,N_19752);
xnor U20020 (N_20020,N_19997,N_19255);
xnor U20021 (N_20021,N_19200,N_19009);
and U20022 (N_20022,N_19198,N_19550);
nor U20023 (N_20023,N_19794,N_19072);
or U20024 (N_20024,N_19502,N_19557);
and U20025 (N_20025,N_19141,N_19853);
xor U20026 (N_20026,N_19302,N_19617);
nand U20027 (N_20027,N_19388,N_19704);
nand U20028 (N_20028,N_19983,N_19737);
xor U20029 (N_20029,N_19783,N_19173);
nand U20030 (N_20030,N_19220,N_19805);
or U20031 (N_20031,N_19197,N_19059);
and U20032 (N_20032,N_19596,N_19207);
or U20033 (N_20033,N_19934,N_19247);
nor U20034 (N_20034,N_19532,N_19750);
and U20035 (N_20035,N_19337,N_19298);
xnor U20036 (N_20036,N_19018,N_19491);
and U20037 (N_20037,N_19150,N_19760);
xnor U20038 (N_20038,N_19265,N_19246);
or U20039 (N_20039,N_19892,N_19762);
xor U20040 (N_20040,N_19126,N_19850);
xnor U20041 (N_20041,N_19208,N_19722);
and U20042 (N_20042,N_19660,N_19415);
xnor U20043 (N_20043,N_19114,N_19082);
and U20044 (N_20044,N_19444,N_19273);
and U20045 (N_20045,N_19217,N_19679);
nand U20046 (N_20046,N_19013,N_19909);
xor U20047 (N_20047,N_19090,N_19672);
nor U20048 (N_20048,N_19578,N_19089);
nand U20049 (N_20049,N_19295,N_19668);
xor U20050 (N_20050,N_19731,N_19925);
and U20051 (N_20051,N_19555,N_19772);
and U20052 (N_20052,N_19418,N_19494);
xnor U20053 (N_20053,N_19188,N_19865);
or U20054 (N_20054,N_19702,N_19205);
nor U20055 (N_20055,N_19168,N_19981);
nand U20056 (N_20056,N_19612,N_19887);
or U20057 (N_20057,N_19308,N_19736);
or U20058 (N_20058,N_19359,N_19355);
or U20059 (N_20059,N_19583,N_19800);
nand U20060 (N_20060,N_19562,N_19228);
xnor U20061 (N_20061,N_19261,N_19875);
and U20062 (N_20062,N_19705,N_19860);
xnor U20063 (N_20063,N_19781,N_19135);
and U20064 (N_20064,N_19918,N_19121);
and U20065 (N_20065,N_19919,N_19021);
and U20066 (N_20066,N_19726,N_19976);
or U20067 (N_20067,N_19361,N_19701);
or U20068 (N_20068,N_19463,N_19180);
or U20069 (N_20069,N_19290,N_19231);
nor U20070 (N_20070,N_19944,N_19739);
nor U20071 (N_20071,N_19658,N_19835);
nand U20072 (N_20072,N_19586,N_19015);
xor U20073 (N_20073,N_19977,N_19024);
nand U20074 (N_20074,N_19263,N_19923);
nand U20075 (N_20075,N_19962,N_19108);
nor U20076 (N_20076,N_19951,N_19878);
nand U20077 (N_20077,N_19427,N_19482);
and U20078 (N_20078,N_19033,N_19998);
and U20079 (N_20079,N_19565,N_19052);
nand U20080 (N_20080,N_19942,N_19629);
and U20081 (N_20081,N_19793,N_19443);
or U20082 (N_20082,N_19464,N_19395);
nor U20083 (N_20083,N_19819,N_19515);
xnor U20084 (N_20084,N_19661,N_19085);
xor U20085 (N_20085,N_19821,N_19226);
nand U20086 (N_20086,N_19788,N_19936);
and U20087 (N_20087,N_19954,N_19215);
nor U20088 (N_20088,N_19456,N_19709);
nor U20089 (N_20089,N_19185,N_19352);
or U20090 (N_20090,N_19124,N_19136);
and U20091 (N_20091,N_19461,N_19434);
nand U20092 (N_20092,N_19467,N_19792);
or U20093 (N_20093,N_19902,N_19797);
nor U20094 (N_20094,N_19852,N_19880);
and U20095 (N_20095,N_19016,N_19432);
nor U20096 (N_20096,N_19607,N_19785);
xor U20097 (N_20097,N_19761,N_19022);
xor U20098 (N_20098,N_19759,N_19256);
nor U20099 (N_20099,N_19802,N_19182);
and U20100 (N_20100,N_19234,N_19581);
xnor U20101 (N_20101,N_19070,N_19632);
nor U20102 (N_20102,N_19161,N_19569);
and U20103 (N_20103,N_19410,N_19639);
or U20104 (N_20104,N_19662,N_19659);
nand U20105 (N_20105,N_19552,N_19963);
nand U20106 (N_20106,N_19333,N_19566);
and U20107 (N_20107,N_19094,N_19286);
nor U20108 (N_20108,N_19548,N_19080);
nand U20109 (N_20109,N_19667,N_19398);
or U20110 (N_20110,N_19677,N_19237);
nor U20111 (N_20111,N_19779,N_19368);
and U20112 (N_20112,N_19353,N_19754);
and U20113 (N_20113,N_19956,N_19331);
and U20114 (N_20114,N_19079,N_19683);
and U20115 (N_20115,N_19949,N_19064);
and U20116 (N_20116,N_19882,N_19966);
nor U20117 (N_20117,N_19282,N_19585);
nor U20118 (N_20118,N_19699,N_19145);
nand U20119 (N_20119,N_19350,N_19157);
nor U20120 (N_20120,N_19253,N_19698);
and U20121 (N_20121,N_19526,N_19155);
or U20122 (N_20122,N_19023,N_19749);
nor U20123 (N_20123,N_19572,N_19961);
xor U20124 (N_20124,N_19299,N_19538);
xor U20125 (N_20125,N_19988,N_19728);
and U20126 (N_20126,N_19965,N_19676);
nand U20127 (N_20127,N_19174,N_19610);
nor U20128 (N_20128,N_19003,N_19127);
nor U20129 (N_20129,N_19602,N_19710);
xnor U20130 (N_20130,N_19268,N_19866);
nor U20131 (N_20131,N_19219,N_19034);
xor U20132 (N_20132,N_19230,N_19686);
xor U20133 (N_20133,N_19561,N_19780);
or U20134 (N_20134,N_19575,N_19623);
xor U20135 (N_20135,N_19641,N_19312);
and U20136 (N_20136,N_19830,N_19424);
or U20137 (N_20137,N_19849,N_19339);
nor U20138 (N_20138,N_19836,N_19688);
or U20139 (N_20139,N_19385,N_19628);
nor U20140 (N_20140,N_19964,N_19861);
xnor U20141 (N_20141,N_19730,N_19289);
nor U20142 (N_20142,N_19099,N_19375);
and U20143 (N_20143,N_19839,N_19871);
nand U20144 (N_20144,N_19175,N_19986);
and U20145 (N_20145,N_19540,N_19650);
or U20146 (N_20146,N_19605,N_19043);
and U20147 (N_20147,N_19036,N_19576);
nor U20148 (N_20148,N_19462,N_19521);
xnor U20149 (N_20149,N_19181,N_19249);
and U20150 (N_20150,N_19810,N_19908);
and U20151 (N_20151,N_19321,N_19322);
nor U20152 (N_20152,N_19159,N_19429);
and U20153 (N_20153,N_19513,N_19275);
nor U20154 (N_20154,N_19573,N_19259);
nand U20155 (N_20155,N_19813,N_19422);
and U20156 (N_20156,N_19828,N_19334);
or U20157 (N_20157,N_19451,N_19738);
nand U20158 (N_20158,N_19401,N_19338);
or U20159 (N_20159,N_19713,N_19518);
or U20160 (N_20160,N_19382,N_19179);
or U20161 (N_20161,N_19656,N_19251);
xnor U20162 (N_20162,N_19031,N_19791);
xnor U20163 (N_20163,N_19915,N_19267);
or U20164 (N_20164,N_19390,N_19869);
xnor U20165 (N_20165,N_19535,N_19397);
nor U20166 (N_20166,N_19019,N_19984);
xnor U20167 (N_20167,N_19320,N_19077);
nor U20168 (N_20168,N_19829,N_19847);
and U20169 (N_20169,N_19905,N_19670);
nand U20170 (N_20170,N_19296,N_19663);
and U20171 (N_20171,N_19364,N_19103);
xnor U20172 (N_20172,N_19503,N_19510);
or U20173 (N_20173,N_19664,N_19500);
xor U20174 (N_20174,N_19883,N_19508);
and U20175 (N_20175,N_19947,N_19735);
or U20176 (N_20176,N_19118,N_19276);
nor U20177 (N_20177,N_19050,N_19439);
and U20178 (N_20178,N_19804,N_19154);
xnor U20179 (N_20179,N_19362,N_19343);
xor U20180 (N_20180,N_19357,N_19638);
nand U20181 (N_20181,N_19164,N_19876);
nor U20182 (N_20182,N_19477,N_19973);
or U20183 (N_20183,N_19140,N_19771);
xor U20184 (N_20184,N_19556,N_19038);
or U20185 (N_20185,N_19724,N_19098);
or U20186 (N_20186,N_19509,N_19392);
nor U20187 (N_20187,N_19472,N_19841);
or U20188 (N_20188,N_19096,N_19584);
xnor U20189 (N_20189,N_19851,N_19943);
or U20190 (N_20190,N_19842,N_19974);
nand U20191 (N_20191,N_19990,N_19536);
nand U20192 (N_20192,N_19864,N_19067);
or U20193 (N_20193,N_19279,N_19405);
nor U20194 (N_20194,N_19590,N_19476);
nand U20195 (N_20195,N_19245,N_19727);
nand U20196 (N_20196,N_19811,N_19931);
xor U20197 (N_20197,N_19137,N_19926);
and U20198 (N_20198,N_19458,N_19862);
and U20199 (N_20199,N_19304,N_19631);
nor U20200 (N_20200,N_19913,N_19907);
and U20201 (N_20201,N_19191,N_19957);
or U20202 (N_20202,N_19520,N_19789);
xnor U20203 (N_20203,N_19172,N_19642);
or U20204 (N_20204,N_19606,N_19158);
and U20205 (N_20205,N_19233,N_19655);
nor U20206 (N_20206,N_19795,N_19592);
nor U20207 (N_20207,N_19845,N_19653);
nand U20208 (N_20208,N_19113,N_19809);
xor U20209 (N_20209,N_19348,N_19032);
and U20210 (N_20210,N_19707,N_19687);
nand U20211 (N_20211,N_19053,N_19591);
nand U20212 (N_20212,N_19884,N_19732);
nor U20213 (N_20213,N_19048,N_19525);
xnor U20214 (N_20214,N_19470,N_19342);
or U20215 (N_20215,N_19719,N_19474);
nand U20216 (N_20216,N_19714,N_19595);
or U20217 (N_20217,N_19857,N_19840);
nor U20218 (N_20218,N_19782,N_19622);
or U20219 (N_20219,N_19978,N_19076);
nor U20220 (N_20220,N_19717,N_19489);
and U20221 (N_20221,N_19529,N_19035);
nand U20222 (N_20222,N_19351,N_19316);
or U20223 (N_20223,N_19012,N_19356);
and U20224 (N_20224,N_19287,N_19579);
nand U20225 (N_20225,N_19652,N_19643);
and U20226 (N_20226,N_19042,N_19407);
xor U20227 (N_20227,N_19488,N_19547);
or U20228 (N_20228,N_19380,N_19450);
nor U20229 (N_20229,N_19818,N_19893);
nor U20230 (N_20230,N_19167,N_19758);
or U20231 (N_20231,N_19325,N_19029);
xnor U20232 (N_20232,N_19896,N_19537);
nand U20233 (N_20233,N_19083,N_19317);
nand U20234 (N_20234,N_19311,N_19729);
nand U20235 (N_20235,N_19305,N_19120);
xnor U20236 (N_20236,N_19859,N_19678);
nor U20237 (N_20237,N_19618,N_19421);
nand U20238 (N_20238,N_19143,N_19153);
xor U20239 (N_20239,N_19326,N_19162);
and U20240 (N_20240,N_19335,N_19027);
xnor U20241 (N_20241,N_19360,N_19692);
and U20242 (N_20242,N_19236,N_19946);
nand U20243 (N_20243,N_19545,N_19874);
nand U20244 (N_20244,N_19673,N_19769);
nand U20245 (N_20245,N_19748,N_19657);
and U20246 (N_20246,N_19318,N_19110);
or U20247 (N_20247,N_19506,N_19193);
nor U20248 (N_20248,N_19512,N_19554);
and U20249 (N_20249,N_19481,N_19697);
nand U20250 (N_20250,N_19466,N_19131);
nand U20251 (N_20251,N_19254,N_19374);
or U20252 (N_20252,N_19235,N_19144);
nand U20253 (N_20253,N_19092,N_19056);
or U20254 (N_20254,N_19693,N_19914);
nand U20255 (N_20255,N_19574,N_19531);
or U20256 (N_20256,N_19347,N_19553);
or U20257 (N_20257,N_19097,N_19453);
nor U20258 (N_20258,N_19309,N_19478);
or U20259 (N_20259,N_19039,N_19227);
and U20260 (N_20260,N_19796,N_19930);
nor U20261 (N_20261,N_19078,N_19720);
nand U20262 (N_20262,N_19209,N_19649);
nor U20263 (N_20263,N_19929,N_19549);
and U20264 (N_20264,N_19437,N_19958);
nor U20265 (N_20265,N_19993,N_19912);
or U20266 (N_20266,N_19533,N_19061);
or U20267 (N_20267,N_19696,N_19903);
or U20268 (N_20268,N_19002,N_19423);
xnor U20269 (N_20269,N_19066,N_19812);
xnor U20270 (N_20270,N_19204,N_19411);
or U20271 (N_20271,N_19123,N_19634);
xnor U20272 (N_20272,N_19329,N_19751);
or U20273 (N_20273,N_19074,N_19952);
and U20274 (N_20274,N_19640,N_19928);
or U20275 (N_20275,N_19045,N_19196);
and U20276 (N_20276,N_19753,N_19774);
xnor U20277 (N_20277,N_19560,N_19277);
and U20278 (N_20278,N_19222,N_19313);
or U20279 (N_20279,N_19480,N_19968);
xor U20280 (N_20280,N_19611,N_19848);
and U20281 (N_20281,N_19384,N_19142);
xnor U20282 (N_20282,N_19877,N_19189);
nor U20283 (N_20283,N_19544,N_19274);
and U20284 (N_20284,N_19571,N_19199);
or U20285 (N_20285,N_19101,N_19773);
xnor U20286 (N_20286,N_19890,N_19358);
nand U20287 (N_20287,N_19694,N_19715);
nor U20288 (N_20288,N_19281,N_19307);
and U20289 (N_20289,N_19497,N_19250);
nand U20290 (N_20290,N_19264,N_19597);
nor U20291 (N_20291,N_19558,N_19551);
or U20292 (N_20292,N_19582,N_19069);
and U20293 (N_20293,N_19646,N_19833);
and U20294 (N_20294,N_19486,N_19937);
xnor U20295 (N_20295,N_19654,N_19522);
and U20296 (N_20296,N_19490,N_19473);
and U20297 (N_20297,N_19455,N_19897);
or U20298 (N_20298,N_19396,N_19703);
nor U20299 (N_20299,N_19487,N_19495);
nand U20300 (N_20300,N_19496,N_19378);
and U20301 (N_20301,N_19169,N_19899);
xnor U20302 (N_20302,N_19160,N_19283);
nor U20303 (N_20303,N_19243,N_19589);
nor U20304 (N_20304,N_19916,N_19995);
and U20305 (N_20305,N_19075,N_19394);
xor U20306 (N_20306,N_19093,N_19449);
or U20307 (N_20307,N_19746,N_19383);
or U20308 (N_20308,N_19542,N_19346);
nand U20309 (N_20309,N_19888,N_19431);
nand U20310 (N_20310,N_19336,N_19402);
xor U20311 (N_20311,N_19680,N_19294);
nor U20312 (N_20312,N_19469,N_19400);
xor U20313 (N_20313,N_19608,N_19178);
nor U20314 (N_20314,N_19425,N_19820);
or U20315 (N_20315,N_19637,N_19156);
nand U20316 (N_20316,N_19365,N_19087);
nor U20317 (N_20317,N_19095,N_19505);
and U20318 (N_20318,N_19546,N_19224);
xnor U20319 (N_20319,N_19370,N_19635);
or U20320 (N_20320,N_19519,N_19814);
and U20321 (N_20321,N_19058,N_19125);
and U20322 (N_20322,N_19146,N_19386);
xnor U20323 (N_20323,N_19613,N_19872);
and U20324 (N_20324,N_19856,N_19242);
or U20325 (N_20325,N_19288,N_19970);
xor U20326 (N_20326,N_19784,N_19524);
or U20327 (N_20327,N_19969,N_19285);
xnor U20328 (N_20328,N_19008,N_19328);
and U20329 (N_20329,N_19239,N_19102);
or U20330 (N_20330,N_19808,N_19559);
and U20331 (N_20331,N_19614,N_19999);
nand U20332 (N_20332,N_19567,N_19006);
nand U20333 (N_20333,N_19898,N_19741);
xnor U20334 (N_20334,N_19776,N_19327);
and U20335 (N_20335,N_19221,N_19081);
xnor U20336 (N_20336,N_19763,N_19873);
or U20337 (N_20337,N_19938,N_19507);
nor U20338 (N_20338,N_19615,N_19684);
nor U20339 (N_20339,N_19436,N_19134);
or U20340 (N_20340,N_19319,N_19733);
nand U20341 (N_20341,N_19803,N_19742);
nor U20342 (N_20342,N_19927,N_19528);
or U20343 (N_20343,N_19723,N_19112);
nor U20344 (N_20344,N_19147,N_19412);
or U20345 (N_20345,N_19924,N_19939);
nor U20346 (N_20346,N_19922,N_19084);
and U20347 (N_20347,N_19933,N_19248);
nand U20348 (N_20348,N_19300,N_19743);
or U20349 (N_20349,N_19363,N_19492);
nor U20350 (N_20350,N_19941,N_19543);
or U20351 (N_20351,N_19297,N_19600);
nand U20352 (N_20352,N_19889,N_19910);
or U20353 (N_20353,N_19895,N_19801);
or U20354 (N_20354,N_19671,N_19238);
nor U20355 (N_20355,N_19354,N_19594);
and U20356 (N_20356,N_19511,N_19212);
nor U20357 (N_20357,N_19211,N_19271);
and U20358 (N_20358,N_19620,N_19109);
and U20359 (N_20359,N_19756,N_19483);
nand U20360 (N_20360,N_19991,N_19460);
nor U20361 (N_20361,N_19960,N_19901);
nand U20362 (N_20362,N_19417,N_19900);
and U20363 (N_20363,N_19106,N_19516);
nand U20364 (N_20364,N_19065,N_19409);
or U20365 (N_20365,N_19420,N_19433);
nand U20366 (N_20366,N_19149,N_19831);
or U20367 (N_20367,N_19823,N_19619);
nand U20368 (N_20368,N_19201,N_19570);
or U20369 (N_20369,N_19391,N_19152);
xor U20370 (N_20370,N_19000,N_19604);
nand U20371 (N_20371,N_19005,N_19278);
nand U20372 (N_20372,N_19139,N_19721);
xnor U20373 (N_20373,N_19030,N_19959);
and U20374 (N_20374,N_19894,N_19445);
nor U20375 (N_20375,N_19539,N_19116);
nand U20376 (N_20376,N_19517,N_19475);
or U20377 (N_20377,N_19689,N_19523);
xor U20378 (N_20378,N_19681,N_19007);
xnor U20379 (N_20379,N_19203,N_19122);
nor U20380 (N_20380,N_19186,N_19225);
nand U20381 (N_20381,N_19240,N_19695);
or U20382 (N_20382,N_19406,N_19244);
nand U20383 (N_20383,N_19117,N_19987);
nand U20384 (N_20384,N_19014,N_19040);
or U20385 (N_20385,N_19301,N_19588);
nand U20386 (N_20386,N_19807,N_19419);
and U20387 (N_20387,N_19745,N_19806);
or U20388 (N_20388,N_19148,N_19371);
or U20389 (N_20389,N_19129,N_19017);
nand U20390 (N_20390,N_19989,N_19344);
nor U20391 (N_20391,N_19971,N_19055);
nand U20392 (N_20392,N_19435,N_19115);
nor U20393 (N_20393,N_19377,N_19992);
xor U20394 (N_20394,N_19270,N_19330);
nor U20395 (N_20395,N_19202,N_19879);
xnor U20396 (N_20396,N_19315,N_19332);
nand U20397 (N_20397,N_19151,N_19471);
nand U20398 (N_20398,N_19091,N_19025);
or U20399 (N_20399,N_19194,N_19786);
nor U20400 (N_20400,N_19184,N_19950);
nor U20401 (N_20401,N_19119,N_19980);
nor U20402 (N_20402,N_19843,N_19485);
or U20403 (N_20403,N_19767,N_19817);
or U20404 (N_20404,N_19948,N_19057);
xnor U20405 (N_20405,N_19493,N_19846);
or U20406 (N_20406,N_19940,N_19967);
and U20407 (N_20407,N_19501,N_19904);
and U20408 (N_20408,N_19373,N_19601);
nand U20409 (N_20409,N_19430,N_19280);
and U20410 (N_20410,N_19844,N_19447);
nor U20411 (N_20411,N_19564,N_19858);
xnor U20412 (N_20412,N_19816,N_19393);
xor U20413 (N_20413,N_19881,N_19366);
and U20414 (N_20414,N_19190,N_19465);
nand U20415 (N_20415,N_19577,N_19624);
nor U20416 (N_20416,N_19177,N_19815);
nand U20417 (N_20417,N_19711,N_19716);
nand U20418 (N_20418,N_19855,N_19306);
or U20419 (N_20419,N_19291,N_19051);
nand U20420 (N_20420,N_19665,N_19504);
and U20421 (N_20421,N_19647,N_19975);
and U20422 (N_20422,N_19917,N_19037);
and U20423 (N_20423,N_19138,N_19935);
nor U20424 (N_20424,N_19324,N_19060);
nor U20425 (N_20425,N_19921,N_19499);
nand U20426 (N_20426,N_19293,N_19046);
or U20427 (N_20427,N_19630,N_19459);
or U20428 (N_20428,N_19764,N_19609);
or U20429 (N_20429,N_19775,N_19438);
or U20430 (N_20430,N_19130,N_19985);
xnor U20431 (N_20431,N_19825,N_19269);
nor U20432 (N_20432,N_19086,N_19798);
or U20433 (N_20433,N_19616,N_19062);
xnor U20434 (N_20434,N_19778,N_19744);
or U20435 (N_20435,N_19484,N_19165);
nor U20436 (N_20436,N_19376,N_19691);
or U20437 (N_20437,N_19626,N_19206);
nor U20438 (N_20438,N_19563,N_19049);
nand U20439 (N_20439,N_19260,N_19568);
or U20440 (N_20440,N_19644,N_19389);
nand U20441 (N_20441,N_19310,N_19195);
nand U20442 (N_20442,N_19932,N_19448);
xor U20443 (N_20443,N_19011,N_19004);
and U20444 (N_20444,N_19787,N_19621);
xnor U20445 (N_20445,N_19527,N_19041);
nor U20446 (N_20446,N_19399,N_19128);
nand U20447 (N_20447,N_19187,N_19837);
and U20448 (N_20448,N_19867,N_19669);
nor U20449 (N_20449,N_19258,N_19765);
xor U20450 (N_20450,N_19911,N_19530);
and U20451 (N_20451,N_19107,N_19100);
xor U20452 (N_20452,N_19367,N_19891);
or U20453 (N_20453,N_19223,N_19028);
nor U20454 (N_20454,N_19416,N_19826);
and U20455 (N_20455,N_19442,N_19369);
or U20456 (N_20456,N_19001,N_19648);
nand U20457 (N_20457,N_19192,N_19026);
or U20458 (N_20458,N_19414,N_19906);
nand U20459 (N_20459,N_19229,N_19381);
or U20460 (N_20460,N_19708,N_19105);
nand U20461 (N_20461,N_19822,N_19682);
nor U20462 (N_20462,N_19440,N_19088);
and U20463 (N_20463,N_19020,N_19718);
or U20464 (N_20464,N_19047,N_19700);
nand U20465 (N_20465,N_19498,N_19747);
and U20466 (N_20466,N_19218,N_19133);
xnor U20467 (N_20467,N_19593,N_19827);
and U20468 (N_20468,N_19071,N_19799);
nor U20469 (N_20469,N_19636,N_19262);
and U20470 (N_20470,N_19068,N_19063);
xnor U20471 (N_20471,N_19777,N_19441);
xor U20472 (N_20472,N_19266,N_19868);
nor U20473 (N_20473,N_19666,N_19674);
nand U20474 (N_20474,N_19832,N_19979);
or U20475 (N_20475,N_19790,N_19073);
or U20476 (N_20476,N_19625,N_19725);
xnor U20477 (N_20477,N_19426,N_19404);
and U20478 (N_20478,N_19408,N_19706);
nand U20479 (N_20479,N_19252,N_19171);
or U20480 (N_20480,N_19387,N_19214);
or U20481 (N_20481,N_19740,N_19010);
nor U20482 (N_20482,N_19755,N_19452);
or U20483 (N_20483,N_19766,N_19690);
nand U20484 (N_20484,N_19824,N_19457);
and U20485 (N_20485,N_19598,N_19712);
and U20486 (N_20486,N_19341,N_19627);
nand U20487 (N_20487,N_19770,N_19272);
nor U20488 (N_20488,N_19863,N_19054);
nor U20489 (N_20489,N_19603,N_19870);
nand U20490 (N_20490,N_19446,N_19213);
nor U20491 (N_20491,N_19651,N_19885);
or U20492 (N_20492,N_19599,N_19176);
and U20493 (N_20493,N_19994,N_19323);
and U20494 (N_20494,N_19104,N_19838);
xnor U20495 (N_20495,N_19241,N_19675);
nor U20496 (N_20496,N_19920,N_19757);
xor U20497 (N_20497,N_19232,N_19345);
and U20498 (N_20498,N_19580,N_19216);
nand U20499 (N_20499,N_19170,N_19514);
nor U20500 (N_20500,N_19244,N_19337);
nand U20501 (N_20501,N_19236,N_19396);
xnor U20502 (N_20502,N_19771,N_19926);
or U20503 (N_20503,N_19932,N_19267);
or U20504 (N_20504,N_19609,N_19684);
xnor U20505 (N_20505,N_19598,N_19411);
or U20506 (N_20506,N_19605,N_19256);
or U20507 (N_20507,N_19124,N_19282);
and U20508 (N_20508,N_19819,N_19553);
nand U20509 (N_20509,N_19641,N_19192);
nor U20510 (N_20510,N_19728,N_19019);
or U20511 (N_20511,N_19070,N_19130);
or U20512 (N_20512,N_19036,N_19785);
xor U20513 (N_20513,N_19147,N_19361);
or U20514 (N_20514,N_19522,N_19253);
and U20515 (N_20515,N_19482,N_19401);
nand U20516 (N_20516,N_19520,N_19909);
or U20517 (N_20517,N_19166,N_19961);
and U20518 (N_20518,N_19190,N_19378);
xnor U20519 (N_20519,N_19357,N_19180);
nand U20520 (N_20520,N_19260,N_19795);
nand U20521 (N_20521,N_19782,N_19251);
and U20522 (N_20522,N_19757,N_19754);
or U20523 (N_20523,N_19548,N_19379);
nand U20524 (N_20524,N_19770,N_19595);
or U20525 (N_20525,N_19071,N_19078);
and U20526 (N_20526,N_19050,N_19732);
or U20527 (N_20527,N_19754,N_19479);
nor U20528 (N_20528,N_19792,N_19082);
xor U20529 (N_20529,N_19491,N_19929);
and U20530 (N_20530,N_19883,N_19388);
or U20531 (N_20531,N_19612,N_19042);
nor U20532 (N_20532,N_19878,N_19815);
nor U20533 (N_20533,N_19561,N_19134);
and U20534 (N_20534,N_19956,N_19202);
nor U20535 (N_20535,N_19744,N_19788);
xnor U20536 (N_20536,N_19662,N_19984);
nand U20537 (N_20537,N_19515,N_19463);
or U20538 (N_20538,N_19415,N_19879);
and U20539 (N_20539,N_19796,N_19562);
xor U20540 (N_20540,N_19442,N_19874);
or U20541 (N_20541,N_19884,N_19350);
nand U20542 (N_20542,N_19980,N_19304);
and U20543 (N_20543,N_19295,N_19263);
xnor U20544 (N_20544,N_19499,N_19243);
nor U20545 (N_20545,N_19418,N_19701);
nand U20546 (N_20546,N_19684,N_19944);
or U20547 (N_20547,N_19696,N_19480);
nand U20548 (N_20548,N_19739,N_19286);
xor U20549 (N_20549,N_19537,N_19148);
or U20550 (N_20550,N_19943,N_19859);
and U20551 (N_20551,N_19935,N_19706);
xnor U20552 (N_20552,N_19412,N_19349);
xnor U20553 (N_20553,N_19119,N_19568);
nand U20554 (N_20554,N_19023,N_19523);
nand U20555 (N_20555,N_19673,N_19795);
nor U20556 (N_20556,N_19222,N_19679);
or U20557 (N_20557,N_19601,N_19089);
nand U20558 (N_20558,N_19177,N_19080);
nand U20559 (N_20559,N_19277,N_19402);
xor U20560 (N_20560,N_19435,N_19736);
or U20561 (N_20561,N_19423,N_19169);
nor U20562 (N_20562,N_19117,N_19806);
nor U20563 (N_20563,N_19218,N_19744);
or U20564 (N_20564,N_19163,N_19958);
or U20565 (N_20565,N_19901,N_19685);
nor U20566 (N_20566,N_19522,N_19421);
and U20567 (N_20567,N_19398,N_19935);
nor U20568 (N_20568,N_19657,N_19782);
and U20569 (N_20569,N_19546,N_19202);
nor U20570 (N_20570,N_19287,N_19125);
nor U20571 (N_20571,N_19512,N_19031);
nand U20572 (N_20572,N_19131,N_19670);
nand U20573 (N_20573,N_19607,N_19661);
xor U20574 (N_20574,N_19031,N_19422);
xnor U20575 (N_20575,N_19408,N_19499);
and U20576 (N_20576,N_19407,N_19741);
nor U20577 (N_20577,N_19584,N_19915);
and U20578 (N_20578,N_19720,N_19513);
or U20579 (N_20579,N_19981,N_19731);
nand U20580 (N_20580,N_19414,N_19940);
nor U20581 (N_20581,N_19548,N_19777);
nand U20582 (N_20582,N_19376,N_19605);
or U20583 (N_20583,N_19721,N_19003);
nor U20584 (N_20584,N_19330,N_19277);
or U20585 (N_20585,N_19514,N_19768);
or U20586 (N_20586,N_19691,N_19163);
xnor U20587 (N_20587,N_19511,N_19232);
xnor U20588 (N_20588,N_19248,N_19657);
nand U20589 (N_20589,N_19154,N_19113);
nor U20590 (N_20590,N_19375,N_19646);
and U20591 (N_20591,N_19631,N_19453);
xnor U20592 (N_20592,N_19092,N_19980);
and U20593 (N_20593,N_19099,N_19610);
xor U20594 (N_20594,N_19651,N_19305);
or U20595 (N_20595,N_19251,N_19654);
nor U20596 (N_20596,N_19908,N_19629);
xnor U20597 (N_20597,N_19138,N_19492);
or U20598 (N_20598,N_19517,N_19213);
or U20599 (N_20599,N_19167,N_19374);
xnor U20600 (N_20600,N_19370,N_19323);
xnor U20601 (N_20601,N_19350,N_19608);
or U20602 (N_20602,N_19277,N_19069);
nand U20603 (N_20603,N_19259,N_19042);
or U20604 (N_20604,N_19994,N_19282);
and U20605 (N_20605,N_19203,N_19209);
xnor U20606 (N_20606,N_19783,N_19913);
nor U20607 (N_20607,N_19662,N_19138);
nor U20608 (N_20608,N_19648,N_19083);
xnor U20609 (N_20609,N_19246,N_19009);
or U20610 (N_20610,N_19141,N_19194);
and U20611 (N_20611,N_19752,N_19060);
or U20612 (N_20612,N_19579,N_19337);
xnor U20613 (N_20613,N_19131,N_19758);
or U20614 (N_20614,N_19090,N_19290);
xnor U20615 (N_20615,N_19556,N_19932);
and U20616 (N_20616,N_19423,N_19575);
or U20617 (N_20617,N_19560,N_19271);
and U20618 (N_20618,N_19883,N_19331);
nor U20619 (N_20619,N_19616,N_19590);
xnor U20620 (N_20620,N_19257,N_19836);
nand U20621 (N_20621,N_19030,N_19540);
nand U20622 (N_20622,N_19551,N_19862);
or U20623 (N_20623,N_19455,N_19804);
nor U20624 (N_20624,N_19881,N_19667);
or U20625 (N_20625,N_19347,N_19922);
nor U20626 (N_20626,N_19403,N_19341);
xor U20627 (N_20627,N_19974,N_19789);
nor U20628 (N_20628,N_19178,N_19408);
nor U20629 (N_20629,N_19085,N_19127);
or U20630 (N_20630,N_19942,N_19539);
nor U20631 (N_20631,N_19354,N_19960);
and U20632 (N_20632,N_19408,N_19044);
and U20633 (N_20633,N_19341,N_19908);
xor U20634 (N_20634,N_19873,N_19793);
nor U20635 (N_20635,N_19557,N_19771);
or U20636 (N_20636,N_19267,N_19854);
xnor U20637 (N_20637,N_19688,N_19802);
and U20638 (N_20638,N_19780,N_19219);
nand U20639 (N_20639,N_19407,N_19323);
or U20640 (N_20640,N_19821,N_19248);
nor U20641 (N_20641,N_19164,N_19968);
or U20642 (N_20642,N_19507,N_19875);
xnor U20643 (N_20643,N_19171,N_19887);
nor U20644 (N_20644,N_19145,N_19542);
and U20645 (N_20645,N_19816,N_19087);
xor U20646 (N_20646,N_19891,N_19800);
nand U20647 (N_20647,N_19793,N_19256);
and U20648 (N_20648,N_19008,N_19117);
and U20649 (N_20649,N_19473,N_19595);
or U20650 (N_20650,N_19537,N_19305);
nand U20651 (N_20651,N_19015,N_19404);
or U20652 (N_20652,N_19116,N_19468);
and U20653 (N_20653,N_19747,N_19907);
and U20654 (N_20654,N_19967,N_19377);
nand U20655 (N_20655,N_19541,N_19702);
xor U20656 (N_20656,N_19326,N_19226);
or U20657 (N_20657,N_19947,N_19742);
xnor U20658 (N_20658,N_19495,N_19843);
xnor U20659 (N_20659,N_19475,N_19471);
xor U20660 (N_20660,N_19901,N_19820);
or U20661 (N_20661,N_19381,N_19384);
nor U20662 (N_20662,N_19596,N_19194);
xnor U20663 (N_20663,N_19044,N_19851);
nor U20664 (N_20664,N_19173,N_19942);
and U20665 (N_20665,N_19715,N_19638);
nand U20666 (N_20666,N_19138,N_19640);
or U20667 (N_20667,N_19891,N_19412);
and U20668 (N_20668,N_19335,N_19948);
nand U20669 (N_20669,N_19594,N_19089);
or U20670 (N_20670,N_19302,N_19200);
nor U20671 (N_20671,N_19737,N_19700);
nor U20672 (N_20672,N_19537,N_19848);
and U20673 (N_20673,N_19484,N_19985);
nand U20674 (N_20674,N_19862,N_19990);
and U20675 (N_20675,N_19809,N_19972);
nand U20676 (N_20676,N_19990,N_19315);
nand U20677 (N_20677,N_19764,N_19958);
nor U20678 (N_20678,N_19121,N_19252);
and U20679 (N_20679,N_19823,N_19967);
and U20680 (N_20680,N_19800,N_19345);
or U20681 (N_20681,N_19463,N_19646);
and U20682 (N_20682,N_19473,N_19617);
and U20683 (N_20683,N_19529,N_19903);
or U20684 (N_20684,N_19726,N_19776);
nor U20685 (N_20685,N_19924,N_19356);
nand U20686 (N_20686,N_19315,N_19092);
xnor U20687 (N_20687,N_19754,N_19423);
nand U20688 (N_20688,N_19790,N_19852);
or U20689 (N_20689,N_19686,N_19740);
nor U20690 (N_20690,N_19745,N_19742);
and U20691 (N_20691,N_19865,N_19694);
xnor U20692 (N_20692,N_19429,N_19462);
or U20693 (N_20693,N_19889,N_19801);
nand U20694 (N_20694,N_19455,N_19336);
or U20695 (N_20695,N_19722,N_19108);
nor U20696 (N_20696,N_19312,N_19723);
or U20697 (N_20697,N_19070,N_19377);
xor U20698 (N_20698,N_19006,N_19443);
xor U20699 (N_20699,N_19089,N_19350);
or U20700 (N_20700,N_19448,N_19459);
or U20701 (N_20701,N_19375,N_19796);
or U20702 (N_20702,N_19185,N_19806);
nand U20703 (N_20703,N_19880,N_19091);
nand U20704 (N_20704,N_19805,N_19409);
or U20705 (N_20705,N_19913,N_19778);
and U20706 (N_20706,N_19614,N_19770);
xnor U20707 (N_20707,N_19090,N_19634);
nand U20708 (N_20708,N_19541,N_19506);
or U20709 (N_20709,N_19811,N_19652);
xnor U20710 (N_20710,N_19472,N_19422);
xnor U20711 (N_20711,N_19982,N_19847);
xnor U20712 (N_20712,N_19191,N_19934);
and U20713 (N_20713,N_19177,N_19912);
and U20714 (N_20714,N_19505,N_19026);
xor U20715 (N_20715,N_19533,N_19116);
and U20716 (N_20716,N_19108,N_19012);
nand U20717 (N_20717,N_19526,N_19442);
nor U20718 (N_20718,N_19165,N_19657);
nand U20719 (N_20719,N_19097,N_19526);
xnor U20720 (N_20720,N_19300,N_19460);
and U20721 (N_20721,N_19822,N_19755);
xor U20722 (N_20722,N_19294,N_19243);
nand U20723 (N_20723,N_19558,N_19718);
and U20724 (N_20724,N_19002,N_19021);
nand U20725 (N_20725,N_19313,N_19511);
xor U20726 (N_20726,N_19813,N_19776);
xor U20727 (N_20727,N_19779,N_19141);
xor U20728 (N_20728,N_19669,N_19444);
nor U20729 (N_20729,N_19611,N_19758);
nand U20730 (N_20730,N_19645,N_19406);
xor U20731 (N_20731,N_19186,N_19519);
and U20732 (N_20732,N_19288,N_19829);
nor U20733 (N_20733,N_19812,N_19223);
and U20734 (N_20734,N_19480,N_19545);
xnor U20735 (N_20735,N_19188,N_19617);
xor U20736 (N_20736,N_19063,N_19182);
and U20737 (N_20737,N_19535,N_19646);
or U20738 (N_20738,N_19274,N_19427);
nor U20739 (N_20739,N_19288,N_19812);
xor U20740 (N_20740,N_19199,N_19011);
xor U20741 (N_20741,N_19448,N_19849);
and U20742 (N_20742,N_19557,N_19206);
nor U20743 (N_20743,N_19385,N_19293);
or U20744 (N_20744,N_19538,N_19911);
and U20745 (N_20745,N_19123,N_19623);
nor U20746 (N_20746,N_19025,N_19413);
and U20747 (N_20747,N_19146,N_19718);
nor U20748 (N_20748,N_19304,N_19910);
xor U20749 (N_20749,N_19442,N_19097);
xor U20750 (N_20750,N_19036,N_19381);
and U20751 (N_20751,N_19749,N_19939);
or U20752 (N_20752,N_19969,N_19520);
or U20753 (N_20753,N_19853,N_19354);
or U20754 (N_20754,N_19380,N_19824);
or U20755 (N_20755,N_19143,N_19192);
nand U20756 (N_20756,N_19050,N_19270);
nor U20757 (N_20757,N_19993,N_19779);
xnor U20758 (N_20758,N_19460,N_19437);
or U20759 (N_20759,N_19297,N_19896);
or U20760 (N_20760,N_19474,N_19645);
nor U20761 (N_20761,N_19229,N_19147);
xor U20762 (N_20762,N_19238,N_19865);
nand U20763 (N_20763,N_19230,N_19890);
nand U20764 (N_20764,N_19188,N_19236);
nor U20765 (N_20765,N_19216,N_19331);
nor U20766 (N_20766,N_19974,N_19915);
xnor U20767 (N_20767,N_19204,N_19070);
and U20768 (N_20768,N_19968,N_19447);
nand U20769 (N_20769,N_19026,N_19697);
nor U20770 (N_20770,N_19292,N_19437);
and U20771 (N_20771,N_19243,N_19255);
nor U20772 (N_20772,N_19883,N_19423);
nand U20773 (N_20773,N_19307,N_19999);
nor U20774 (N_20774,N_19763,N_19776);
nor U20775 (N_20775,N_19358,N_19401);
nor U20776 (N_20776,N_19246,N_19677);
nor U20777 (N_20777,N_19408,N_19345);
xnor U20778 (N_20778,N_19378,N_19739);
nand U20779 (N_20779,N_19687,N_19160);
xnor U20780 (N_20780,N_19806,N_19622);
nor U20781 (N_20781,N_19839,N_19783);
and U20782 (N_20782,N_19093,N_19385);
and U20783 (N_20783,N_19970,N_19370);
xnor U20784 (N_20784,N_19097,N_19020);
and U20785 (N_20785,N_19373,N_19194);
or U20786 (N_20786,N_19201,N_19694);
nand U20787 (N_20787,N_19677,N_19682);
and U20788 (N_20788,N_19682,N_19142);
nor U20789 (N_20789,N_19582,N_19120);
nand U20790 (N_20790,N_19660,N_19192);
xor U20791 (N_20791,N_19222,N_19617);
nand U20792 (N_20792,N_19357,N_19876);
and U20793 (N_20793,N_19571,N_19028);
nand U20794 (N_20794,N_19235,N_19680);
or U20795 (N_20795,N_19040,N_19420);
xor U20796 (N_20796,N_19376,N_19471);
nor U20797 (N_20797,N_19157,N_19334);
nand U20798 (N_20798,N_19607,N_19266);
and U20799 (N_20799,N_19368,N_19900);
nand U20800 (N_20800,N_19032,N_19415);
nor U20801 (N_20801,N_19994,N_19697);
or U20802 (N_20802,N_19686,N_19681);
nand U20803 (N_20803,N_19130,N_19721);
nand U20804 (N_20804,N_19746,N_19968);
nor U20805 (N_20805,N_19957,N_19029);
or U20806 (N_20806,N_19895,N_19747);
or U20807 (N_20807,N_19795,N_19298);
nand U20808 (N_20808,N_19586,N_19482);
or U20809 (N_20809,N_19462,N_19558);
and U20810 (N_20810,N_19679,N_19800);
xnor U20811 (N_20811,N_19772,N_19805);
nand U20812 (N_20812,N_19086,N_19077);
nor U20813 (N_20813,N_19884,N_19896);
nor U20814 (N_20814,N_19958,N_19793);
nand U20815 (N_20815,N_19450,N_19714);
and U20816 (N_20816,N_19893,N_19662);
and U20817 (N_20817,N_19460,N_19200);
and U20818 (N_20818,N_19314,N_19105);
and U20819 (N_20819,N_19371,N_19329);
nor U20820 (N_20820,N_19741,N_19004);
xnor U20821 (N_20821,N_19781,N_19235);
or U20822 (N_20822,N_19660,N_19842);
or U20823 (N_20823,N_19725,N_19706);
or U20824 (N_20824,N_19787,N_19982);
or U20825 (N_20825,N_19916,N_19311);
or U20826 (N_20826,N_19186,N_19409);
nor U20827 (N_20827,N_19098,N_19140);
nor U20828 (N_20828,N_19805,N_19581);
nor U20829 (N_20829,N_19568,N_19696);
nand U20830 (N_20830,N_19855,N_19325);
or U20831 (N_20831,N_19990,N_19108);
or U20832 (N_20832,N_19023,N_19534);
nor U20833 (N_20833,N_19782,N_19801);
or U20834 (N_20834,N_19721,N_19695);
nor U20835 (N_20835,N_19296,N_19843);
or U20836 (N_20836,N_19023,N_19941);
or U20837 (N_20837,N_19408,N_19837);
xor U20838 (N_20838,N_19970,N_19001);
and U20839 (N_20839,N_19217,N_19396);
nand U20840 (N_20840,N_19382,N_19922);
nand U20841 (N_20841,N_19610,N_19077);
and U20842 (N_20842,N_19525,N_19742);
or U20843 (N_20843,N_19475,N_19438);
nand U20844 (N_20844,N_19752,N_19551);
nor U20845 (N_20845,N_19689,N_19902);
or U20846 (N_20846,N_19169,N_19717);
nand U20847 (N_20847,N_19206,N_19227);
nand U20848 (N_20848,N_19056,N_19285);
nor U20849 (N_20849,N_19573,N_19019);
xnor U20850 (N_20850,N_19781,N_19017);
nand U20851 (N_20851,N_19531,N_19287);
xnor U20852 (N_20852,N_19109,N_19893);
and U20853 (N_20853,N_19618,N_19756);
and U20854 (N_20854,N_19644,N_19314);
or U20855 (N_20855,N_19018,N_19341);
xnor U20856 (N_20856,N_19362,N_19784);
nor U20857 (N_20857,N_19254,N_19783);
nand U20858 (N_20858,N_19980,N_19965);
or U20859 (N_20859,N_19386,N_19764);
nor U20860 (N_20860,N_19342,N_19900);
nor U20861 (N_20861,N_19321,N_19763);
nor U20862 (N_20862,N_19441,N_19351);
nand U20863 (N_20863,N_19657,N_19641);
xnor U20864 (N_20864,N_19238,N_19321);
or U20865 (N_20865,N_19508,N_19229);
nand U20866 (N_20866,N_19231,N_19470);
or U20867 (N_20867,N_19015,N_19139);
nor U20868 (N_20868,N_19192,N_19907);
xnor U20869 (N_20869,N_19088,N_19037);
xor U20870 (N_20870,N_19392,N_19824);
and U20871 (N_20871,N_19890,N_19319);
nand U20872 (N_20872,N_19859,N_19126);
xnor U20873 (N_20873,N_19342,N_19019);
nand U20874 (N_20874,N_19174,N_19492);
and U20875 (N_20875,N_19054,N_19549);
xnor U20876 (N_20876,N_19948,N_19243);
nand U20877 (N_20877,N_19346,N_19954);
and U20878 (N_20878,N_19685,N_19362);
xnor U20879 (N_20879,N_19188,N_19175);
nand U20880 (N_20880,N_19533,N_19568);
and U20881 (N_20881,N_19371,N_19557);
and U20882 (N_20882,N_19035,N_19551);
and U20883 (N_20883,N_19987,N_19286);
and U20884 (N_20884,N_19283,N_19586);
nor U20885 (N_20885,N_19438,N_19824);
or U20886 (N_20886,N_19746,N_19609);
nand U20887 (N_20887,N_19985,N_19548);
nand U20888 (N_20888,N_19527,N_19736);
nand U20889 (N_20889,N_19665,N_19080);
xnor U20890 (N_20890,N_19391,N_19959);
or U20891 (N_20891,N_19897,N_19251);
nand U20892 (N_20892,N_19655,N_19443);
nand U20893 (N_20893,N_19855,N_19440);
nor U20894 (N_20894,N_19689,N_19120);
xor U20895 (N_20895,N_19663,N_19007);
and U20896 (N_20896,N_19143,N_19009);
xnor U20897 (N_20897,N_19516,N_19450);
nand U20898 (N_20898,N_19849,N_19403);
nor U20899 (N_20899,N_19264,N_19212);
nand U20900 (N_20900,N_19340,N_19318);
nor U20901 (N_20901,N_19885,N_19300);
or U20902 (N_20902,N_19494,N_19472);
nand U20903 (N_20903,N_19545,N_19897);
xor U20904 (N_20904,N_19161,N_19295);
and U20905 (N_20905,N_19232,N_19767);
nand U20906 (N_20906,N_19684,N_19368);
nand U20907 (N_20907,N_19394,N_19868);
xnor U20908 (N_20908,N_19269,N_19519);
nor U20909 (N_20909,N_19166,N_19778);
nand U20910 (N_20910,N_19290,N_19339);
nor U20911 (N_20911,N_19731,N_19447);
or U20912 (N_20912,N_19211,N_19522);
xnor U20913 (N_20913,N_19585,N_19444);
nor U20914 (N_20914,N_19710,N_19423);
nor U20915 (N_20915,N_19089,N_19256);
nor U20916 (N_20916,N_19592,N_19477);
nor U20917 (N_20917,N_19072,N_19443);
xor U20918 (N_20918,N_19588,N_19741);
nand U20919 (N_20919,N_19894,N_19154);
or U20920 (N_20920,N_19019,N_19593);
or U20921 (N_20921,N_19200,N_19029);
or U20922 (N_20922,N_19071,N_19314);
nor U20923 (N_20923,N_19321,N_19849);
and U20924 (N_20924,N_19865,N_19544);
nand U20925 (N_20925,N_19316,N_19333);
nand U20926 (N_20926,N_19662,N_19982);
or U20927 (N_20927,N_19011,N_19745);
xnor U20928 (N_20928,N_19873,N_19326);
or U20929 (N_20929,N_19739,N_19805);
xor U20930 (N_20930,N_19511,N_19098);
nand U20931 (N_20931,N_19876,N_19428);
or U20932 (N_20932,N_19403,N_19982);
xor U20933 (N_20933,N_19811,N_19974);
or U20934 (N_20934,N_19456,N_19966);
and U20935 (N_20935,N_19075,N_19692);
and U20936 (N_20936,N_19661,N_19631);
nand U20937 (N_20937,N_19106,N_19237);
or U20938 (N_20938,N_19877,N_19165);
nor U20939 (N_20939,N_19421,N_19974);
nor U20940 (N_20940,N_19989,N_19832);
nor U20941 (N_20941,N_19813,N_19736);
nor U20942 (N_20942,N_19958,N_19456);
or U20943 (N_20943,N_19196,N_19770);
xnor U20944 (N_20944,N_19377,N_19733);
or U20945 (N_20945,N_19156,N_19644);
nor U20946 (N_20946,N_19975,N_19492);
xor U20947 (N_20947,N_19036,N_19081);
and U20948 (N_20948,N_19129,N_19505);
or U20949 (N_20949,N_19587,N_19720);
xor U20950 (N_20950,N_19227,N_19212);
nor U20951 (N_20951,N_19677,N_19070);
and U20952 (N_20952,N_19037,N_19406);
nor U20953 (N_20953,N_19960,N_19390);
xnor U20954 (N_20954,N_19452,N_19480);
xnor U20955 (N_20955,N_19862,N_19417);
or U20956 (N_20956,N_19315,N_19197);
and U20957 (N_20957,N_19123,N_19299);
xnor U20958 (N_20958,N_19704,N_19279);
and U20959 (N_20959,N_19906,N_19293);
nor U20960 (N_20960,N_19028,N_19077);
xor U20961 (N_20961,N_19837,N_19046);
nor U20962 (N_20962,N_19311,N_19322);
and U20963 (N_20963,N_19862,N_19233);
or U20964 (N_20964,N_19013,N_19487);
nor U20965 (N_20965,N_19290,N_19561);
nand U20966 (N_20966,N_19991,N_19643);
xnor U20967 (N_20967,N_19740,N_19424);
nand U20968 (N_20968,N_19562,N_19971);
or U20969 (N_20969,N_19355,N_19256);
nor U20970 (N_20970,N_19033,N_19199);
and U20971 (N_20971,N_19932,N_19791);
and U20972 (N_20972,N_19743,N_19431);
and U20973 (N_20973,N_19194,N_19237);
xnor U20974 (N_20974,N_19872,N_19866);
nor U20975 (N_20975,N_19082,N_19710);
or U20976 (N_20976,N_19294,N_19794);
and U20977 (N_20977,N_19446,N_19903);
nor U20978 (N_20978,N_19871,N_19214);
nor U20979 (N_20979,N_19049,N_19211);
and U20980 (N_20980,N_19181,N_19415);
and U20981 (N_20981,N_19270,N_19630);
or U20982 (N_20982,N_19994,N_19174);
nand U20983 (N_20983,N_19736,N_19598);
xor U20984 (N_20984,N_19182,N_19861);
xnor U20985 (N_20985,N_19351,N_19245);
nor U20986 (N_20986,N_19559,N_19778);
and U20987 (N_20987,N_19449,N_19652);
or U20988 (N_20988,N_19254,N_19739);
nand U20989 (N_20989,N_19816,N_19853);
nor U20990 (N_20990,N_19224,N_19148);
nand U20991 (N_20991,N_19273,N_19718);
nand U20992 (N_20992,N_19909,N_19097);
xnor U20993 (N_20993,N_19931,N_19643);
nand U20994 (N_20994,N_19525,N_19510);
nand U20995 (N_20995,N_19921,N_19831);
nor U20996 (N_20996,N_19837,N_19923);
or U20997 (N_20997,N_19900,N_19009);
nand U20998 (N_20998,N_19836,N_19429);
or U20999 (N_20999,N_19750,N_19630);
nand U21000 (N_21000,N_20258,N_20277);
and U21001 (N_21001,N_20122,N_20235);
nor U21002 (N_21002,N_20095,N_20520);
and U21003 (N_21003,N_20852,N_20367);
or U21004 (N_21004,N_20265,N_20603);
xor U21005 (N_21005,N_20755,N_20771);
or U21006 (N_21006,N_20613,N_20287);
nor U21007 (N_21007,N_20250,N_20271);
and U21008 (N_21008,N_20004,N_20849);
nand U21009 (N_21009,N_20928,N_20704);
xnor U21010 (N_21010,N_20042,N_20665);
or U21011 (N_21011,N_20306,N_20978);
xnor U21012 (N_21012,N_20161,N_20406);
or U21013 (N_21013,N_20407,N_20888);
xor U21014 (N_21014,N_20365,N_20024);
nor U21015 (N_21015,N_20997,N_20001);
xnor U21016 (N_21016,N_20386,N_20632);
nand U21017 (N_21017,N_20991,N_20425);
nor U21018 (N_21018,N_20240,N_20896);
nor U21019 (N_21019,N_20804,N_20033);
nand U21020 (N_21020,N_20319,N_20430);
nor U21021 (N_21021,N_20730,N_20171);
nor U21022 (N_21022,N_20090,N_20492);
xor U21023 (N_21023,N_20213,N_20894);
xnor U21024 (N_21024,N_20950,N_20146);
nand U21025 (N_21025,N_20253,N_20854);
xor U21026 (N_21026,N_20708,N_20673);
nand U21027 (N_21027,N_20035,N_20156);
xnor U21028 (N_21028,N_20121,N_20479);
nor U21029 (N_21029,N_20263,N_20155);
xnor U21030 (N_21030,N_20356,N_20393);
xor U21031 (N_21031,N_20858,N_20984);
nor U21032 (N_21032,N_20985,N_20521);
nor U21033 (N_21033,N_20838,N_20623);
nor U21034 (N_21034,N_20802,N_20916);
and U21035 (N_21035,N_20812,N_20329);
nor U21036 (N_21036,N_20792,N_20591);
nor U21037 (N_21037,N_20504,N_20296);
nor U21038 (N_21038,N_20311,N_20816);
nand U21039 (N_21039,N_20421,N_20501);
xnor U21040 (N_21040,N_20625,N_20480);
and U21041 (N_21041,N_20357,N_20691);
xor U21042 (N_21042,N_20220,N_20210);
nand U21043 (N_21043,N_20962,N_20526);
nand U21044 (N_21044,N_20661,N_20557);
nand U21045 (N_21045,N_20998,N_20655);
nand U21046 (N_21046,N_20688,N_20494);
nor U21047 (N_21047,N_20843,N_20954);
nor U21048 (N_21048,N_20731,N_20151);
nand U21049 (N_21049,N_20284,N_20753);
or U21050 (N_21050,N_20461,N_20199);
or U21051 (N_21051,N_20579,N_20604);
nand U21052 (N_21052,N_20460,N_20869);
xor U21053 (N_21053,N_20911,N_20019);
nand U21054 (N_21054,N_20369,N_20021);
nand U21055 (N_21055,N_20509,N_20270);
xnor U21056 (N_21056,N_20580,N_20044);
or U21057 (N_21057,N_20405,N_20295);
nand U21058 (N_21058,N_20674,N_20723);
nor U21059 (N_21059,N_20178,N_20535);
and U21060 (N_21060,N_20262,N_20115);
nand U21061 (N_21061,N_20765,N_20397);
or U21062 (N_21062,N_20966,N_20681);
or U21063 (N_21063,N_20427,N_20760);
nand U21064 (N_21064,N_20261,N_20154);
nand U21065 (N_21065,N_20117,N_20193);
nor U21066 (N_21066,N_20182,N_20464);
xor U21067 (N_21067,N_20370,N_20990);
xnor U21068 (N_21068,N_20441,N_20190);
and U21069 (N_21069,N_20634,N_20401);
nor U21070 (N_21070,N_20725,N_20077);
and U21071 (N_21071,N_20545,N_20546);
and U21072 (N_21072,N_20818,N_20813);
or U21073 (N_21073,N_20629,N_20498);
nand U21074 (N_21074,N_20388,N_20690);
nor U21075 (N_21075,N_20744,N_20943);
nand U21076 (N_21076,N_20646,N_20880);
nor U21077 (N_21077,N_20018,N_20946);
nand U21078 (N_21078,N_20354,N_20003);
xnor U21079 (N_21079,N_20639,N_20570);
xor U21080 (N_21080,N_20882,N_20039);
nor U21081 (N_21081,N_20915,N_20067);
and U21082 (N_21082,N_20842,N_20640);
nand U21083 (N_21083,N_20617,N_20175);
or U21084 (N_21084,N_20951,N_20703);
and U21085 (N_21085,N_20973,N_20531);
nand U21086 (N_21086,N_20543,N_20170);
nand U21087 (N_21087,N_20566,N_20736);
xor U21088 (N_21088,N_20958,N_20833);
nor U21089 (N_21089,N_20884,N_20508);
or U21090 (N_21090,N_20205,N_20351);
or U21091 (N_21091,N_20599,N_20685);
or U21092 (N_21092,N_20582,N_20255);
nor U21093 (N_21093,N_20132,N_20874);
and U21094 (N_21094,N_20358,N_20469);
xnor U21095 (N_21095,N_20721,N_20794);
nand U21096 (N_21096,N_20123,N_20179);
nor U21097 (N_21097,N_20457,N_20831);
and U21098 (N_21098,N_20947,N_20314);
nand U21099 (N_21099,N_20815,N_20519);
xnor U21100 (N_21100,N_20791,N_20030);
or U21101 (N_21101,N_20658,N_20248);
or U21102 (N_21102,N_20717,N_20124);
or U21103 (N_21103,N_20993,N_20638);
nand U21104 (N_21104,N_20740,N_20739);
nor U21105 (N_21105,N_20201,N_20800);
and U21106 (N_21106,N_20374,N_20017);
nor U21107 (N_21107,N_20128,N_20168);
and U21108 (N_21108,N_20805,N_20411);
nand U21109 (N_21109,N_20610,N_20169);
xnor U21110 (N_21110,N_20260,N_20288);
xor U21111 (N_21111,N_20559,N_20062);
nand U21112 (N_21112,N_20780,N_20699);
or U21113 (N_21113,N_20225,N_20893);
or U21114 (N_21114,N_20490,N_20249);
and U21115 (N_21115,N_20470,N_20147);
or U21116 (N_21116,N_20862,N_20131);
nand U21117 (N_21117,N_20575,N_20848);
nor U21118 (N_21118,N_20477,N_20788);
and U21119 (N_21119,N_20701,N_20502);
or U21120 (N_21120,N_20987,N_20034);
nand U21121 (N_21121,N_20663,N_20207);
nand U21122 (N_21122,N_20204,N_20925);
nor U21123 (N_21123,N_20627,N_20049);
or U21124 (N_21124,N_20085,N_20025);
and U21125 (N_21125,N_20056,N_20809);
xor U21126 (N_21126,N_20432,N_20404);
nor U21127 (N_21127,N_20586,N_20098);
nand U21128 (N_21128,N_20403,N_20105);
xnor U21129 (N_21129,N_20415,N_20851);
xnor U21130 (N_21130,N_20114,N_20961);
xnor U21131 (N_21131,N_20408,N_20172);
xor U21132 (N_21132,N_20014,N_20530);
or U21133 (N_21133,N_20980,N_20279);
xor U21134 (N_21134,N_20960,N_20944);
or U21135 (N_21135,N_20387,N_20402);
and U21136 (N_21136,N_20410,N_20165);
nand U21137 (N_21137,N_20054,N_20899);
nand U21138 (N_21138,N_20895,N_20633);
and U21139 (N_21139,N_20724,N_20601);
nor U21140 (N_21140,N_20138,N_20338);
xor U21141 (N_21141,N_20865,N_20619);
and U21142 (N_21142,N_20481,N_20359);
nand U21143 (N_21143,N_20116,N_20992);
and U21144 (N_21144,N_20472,N_20709);
and U21145 (N_21145,N_20636,N_20221);
nand U21146 (N_21146,N_20873,N_20215);
or U21147 (N_21147,N_20227,N_20819);
nand U21148 (N_21148,N_20229,N_20289);
xnor U21149 (N_21149,N_20549,N_20103);
and U21150 (N_21150,N_20259,N_20891);
and U21151 (N_21151,N_20841,N_20918);
nor U21152 (N_21152,N_20824,N_20418);
or U21153 (N_21153,N_20883,N_20676);
and U21154 (N_21154,N_20251,N_20879);
xor U21155 (N_21155,N_20994,N_20737);
and U21156 (N_21156,N_20206,N_20308);
and U21157 (N_21157,N_20560,N_20316);
and U21158 (N_21158,N_20878,N_20621);
and U21159 (N_21159,N_20125,N_20332);
nor U21160 (N_21160,N_20533,N_20912);
and U21161 (N_21161,N_20588,N_20798);
and U21162 (N_21162,N_20423,N_20107);
and U21163 (N_21163,N_20705,N_20196);
nor U21164 (N_21164,N_20257,N_20064);
xnor U21165 (N_21165,N_20456,N_20145);
xor U21166 (N_21166,N_20438,N_20647);
xnor U21167 (N_21167,N_20007,N_20746);
and U21168 (N_21168,N_20963,N_20949);
or U21169 (N_21169,N_20795,N_20551);
xnor U21170 (N_21170,N_20174,N_20194);
xor U21171 (N_21171,N_20965,N_20563);
and U21172 (N_21172,N_20377,N_20109);
and U21173 (N_21173,N_20675,N_20136);
and U21174 (N_21174,N_20821,N_20217);
nand U21175 (N_21175,N_20304,N_20781);
xnor U21176 (N_21176,N_20431,N_20719);
nand U21177 (N_21177,N_20399,N_20784);
nor U21178 (N_21178,N_20529,N_20930);
and U21179 (N_21179,N_20097,N_20935);
and U21180 (N_21180,N_20597,N_20075);
nand U21181 (N_21181,N_20614,N_20010);
nand U21182 (N_21182,N_20167,N_20157);
and U21183 (N_21183,N_20129,N_20600);
or U21184 (N_21184,N_20900,N_20073);
nand U21185 (N_21185,N_20137,N_20409);
and U21186 (N_21186,N_20330,N_20327);
nand U21187 (N_21187,N_20528,N_20828);
xor U21188 (N_21188,N_20484,N_20714);
or U21189 (N_21189,N_20023,N_20513);
or U21190 (N_21190,N_20786,N_20086);
or U21191 (N_21191,N_20626,N_20483);
xnor U21192 (N_21192,N_20198,N_20995);
nand U21193 (N_21193,N_20274,N_20364);
xnor U21194 (N_21194,N_20444,N_20555);
nor U21195 (N_21195,N_20986,N_20102);
or U21196 (N_21196,N_20981,N_20176);
nor U21197 (N_21197,N_20081,N_20602);
or U21198 (N_21198,N_20923,N_20245);
nor U21199 (N_21199,N_20343,N_20320);
nor U21200 (N_21200,N_20452,N_20803);
nor U21201 (N_21201,N_20130,N_20334);
or U21202 (N_21202,N_20910,N_20875);
nand U21203 (N_21203,N_20148,N_20202);
nand U21204 (N_21204,N_20488,N_20941);
nor U21205 (N_21205,N_20106,N_20996);
and U21206 (N_21206,N_20362,N_20463);
xnor U21207 (N_21207,N_20808,N_20897);
or U21208 (N_21208,N_20341,N_20904);
nand U21209 (N_21209,N_20061,N_20337);
or U21210 (N_21210,N_20173,N_20127);
nor U21211 (N_21211,N_20133,N_20903);
nor U21212 (N_21212,N_20416,N_20301);
and U21213 (N_21213,N_20635,N_20696);
nor U21214 (N_21214,N_20671,N_20135);
nand U21215 (N_21215,N_20028,N_20777);
nand U21216 (N_21216,N_20518,N_20378);
or U21217 (N_21217,N_20593,N_20066);
xnor U21218 (N_21218,N_20983,N_20219);
nand U21219 (N_21219,N_20368,N_20389);
nor U21220 (N_21220,N_20697,N_20534);
xnor U21221 (N_21221,N_20055,N_20269);
nand U21222 (N_21222,N_20398,N_20385);
or U21223 (N_21223,N_20391,N_20434);
nand U21224 (N_21224,N_20268,N_20743);
or U21225 (N_21225,N_20298,N_20226);
or U21226 (N_21226,N_20952,N_20544);
or U21227 (N_21227,N_20796,N_20829);
or U21228 (N_21228,N_20845,N_20793);
nand U21229 (N_21229,N_20074,N_20203);
xnor U21230 (N_21230,N_20233,N_20093);
xnor U21231 (N_21231,N_20554,N_20473);
nand U21232 (N_21232,N_20458,N_20454);
xnor U21233 (N_21233,N_20342,N_20037);
or U21234 (N_21234,N_20956,N_20113);
or U21235 (N_21235,N_20487,N_20373);
nor U21236 (N_21236,N_20380,N_20547);
and U21237 (N_21237,N_20797,N_20905);
nor U21238 (N_21238,N_20767,N_20119);
and U21239 (N_21239,N_20015,N_20336);
nand U21240 (N_21240,N_20187,N_20682);
and U21241 (N_21241,N_20971,N_20111);
nand U21242 (N_21242,N_20325,N_20293);
and U21243 (N_21243,N_20244,N_20009);
nand U21244 (N_21244,N_20936,N_20331);
xnor U21245 (N_21245,N_20817,N_20283);
nor U21246 (N_21246,N_20550,N_20340);
and U21247 (N_21247,N_20678,N_20726);
or U21248 (N_21248,N_20143,N_20867);
or U21249 (N_21249,N_20525,N_20556);
nand U21250 (N_21250,N_20729,N_20092);
or U21251 (N_21251,N_20641,N_20192);
nand U21252 (N_21252,N_20058,N_20945);
xor U21253 (N_21253,N_20710,N_20578);
nor U21254 (N_21254,N_20861,N_20906);
nand U21255 (N_21255,N_20242,N_20745);
nor U21256 (N_21256,N_20186,N_20063);
and U21257 (N_21257,N_20188,N_20762);
and U21258 (N_21258,N_20008,N_20939);
xor U21259 (N_21259,N_20027,N_20363);
or U21260 (N_21260,N_20738,N_20022);
nand U21261 (N_21261,N_20934,N_20307);
or U21262 (N_21262,N_20615,N_20439);
or U21263 (N_21263,N_20517,N_20382);
and U21264 (N_21264,N_20419,N_20209);
nor U21265 (N_21265,N_20384,N_20768);
or U21266 (N_21266,N_20637,N_20505);
and U21267 (N_21267,N_20564,N_20216);
and U21268 (N_21268,N_20511,N_20806);
nand U21269 (N_21269,N_20853,N_20751);
nand U21270 (N_21270,N_20101,N_20392);
xor U21271 (N_21271,N_20069,N_20686);
nand U21272 (N_21272,N_20970,N_20353);
or U21273 (N_21273,N_20785,N_20496);
or U21274 (N_21274,N_20955,N_20761);
nand U21275 (N_21275,N_20072,N_20715);
and U21276 (N_21276,N_20592,N_20989);
and U21277 (N_21277,N_20653,N_20038);
and U21278 (N_21278,N_20292,N_20720);
and U21279 (N_21279,N_20065,N_20390);
and U21280 (N_21280,N_20503,N_20512);
nor U21281 (N_21281,N_20026,N_20413);
nor U21282 (N_21282,N_20727,N_20344);
nor U21283 (N_21283,N_20442,N_20012);
and U21284 (N_21284,N_20576,N_20747);
xnor U21285 (N_21285,N_20648,N_20266);
nand U21286 (N_21286,N_20857,N_20684);
xnor U21287 (N_21287,N_20628,N_20013);
xor U21288 (N_21288,N_20752,N_20222);
nand U21289 (N_21289,N_20810,N_20732);
nor U21290 (N_21290,N_20567,N_20881);
nor U21291 (N_21291,N_20087,N_20666);
nor U21292 (N_21292,N_20913,N_20158);
or U21293 (N_21293,N_20664,N_20677);
and U21294 (N_21294,N_20863,N_20153);
xor U21295 (N_21295,N_20449,N_20361);
or U21296 (N_21296,N_20999,N_20396);
xnor U21297 (N_21297,N_20532,N_20223);
and U21298 (N_21298,N_20376,N_20185);
nor U21299 (N_21299,N_20975,N_20749);
or U21300 (N_21300,N_20820,N_20741);
and U21301 (N_21301,N_20823,N_20687);
nor U21302 (N_21302,N_20937,N_20609);
nand U21303 (N_21303,N_20281,N_20352);
and U21304 (N_21304,N_20197,N_20247);
nor U21305 (N_21305,N_20914,N_20428);
and U21306 (N_21306,N_20596,N_20537);
or U21307 (N_21307,N_20887,N_20126);
nor U21308 (N_21308,N_20450,N_20683);
xnor U21309 (N_21309,N_20921,N_20830);
nor U21310 (N_21310,N_20006,N_20650);
nor U21311 (N_21311,N_20902,N_20680);
and U21312 (N_21312,N_20150,N_20968);
nand U21313 (N_21313,N_20290,N_20080);
nor U21314 (N_21314,N_20079,N_20548);
nor U21315 (N_21315,N_20889,N_20754);
nand U21316 (N_21316,N_20144,N_20670);
nand U21317 (N_21317,N_20318,N_20275);
nor U21318 (N_21318,N_20349,N_20224);
nand U21319 (N_21319,N_20585,N_20139);
nand U21320 (N_21320,N_20510,N_20618);
or U21321 (N_21321,N_20569,N_20451);
and U21322 (N_21322,N_20909,N_20595);
nor U21323 (N_21323,N_20466,N_20246);
nand U21324 (N_21324,N_20475,N_20099);
xor U21325 (N_21325,N_20573,N_20982);
xor U21326 (N_21326,N_20572,N_20486);
or U21327 (N_21327,N_20459,N_20908);
and U21328 (N_21328,N_20612,N_20890);
xor U21329 (N_21329,N_20507,N_20850);
and U21330 (N_21330,N_20668,N_20834);
and U21331 (N_21331,N_20032,N_20787);
or U21332 (N_21332,N_20482,N_20395);
nand U21333 (N_21333,N_20825,N_20571);
xor U21334 (N_21334,N_20541,N_20345);
xor U21335 (N_21335,N_20043,N_20931);
and U21336 (N_21336,N_20807,N_20231);
or U21337 (N_21337,N_20907,N_20651);
nand U21338 (N_21338,N_20538,N_20429);
nor U21339 (N_21339,N_20256,N_20149);
and U21340 (N_21340,N_20558,N_20278);
nand U21341 (N_21341,N_20321,N_20748);
or U21342 (N_21342,N_20181,N_20514);
and U21343 (N_21343,N_20052,N_20104);
xnor U21344 (N_21344,N_20642,N_20814);
nor U21345 (N_21345,N_20422,N_20191);
and U21346 (N_21346,N_20622,N_20238);
or U21347 (N_21347,N_20577,N_20346);
or U21348 (N_21348,N_20323,N_20587);
nor U21349 (N_21349,N_20412,N_20214);
or U21350 (N_21350,N_20654,N_20299);
nor U21351 (N_21351,N_20379,N_20047);
nand U21352 (N_21352,N_20177,N_20826);
or U21353 (N_21353,N_20424,N_20722);
nand U21354 (N_21354,N_20005,N_20692);
nand U21355 (N_21355,N_20649,N_20478);
or U21356 (N_21356,N_20164,N_20076);
nor U21357 (N_21357,N_20059,N_20134);
nand U21358 (N_21358,N_20051,N_20462);
nand U21359 (N_21359,N_20166,N_20071);
nand U21360 (N_21360,N_20660,N_20522);
or U21361 (N_21361,N_20228,N_20088);
and U21362 (N_21362,N_20892,N_20426);
or U21363 (N_21363,N_20964,N_20309);
and U21364 (N_21364,N_20162,N_20300);
or U21365 (N_21365,N_20734,N_20789);
and U21366 (N_21366,N_20212,N_20078);
and U21367 (N_21367,N_20180,N_20118);
or U21368 (N_21368,N_20790,N_20467);
and U21369 (N_21369,N_20801,N_20757);
xnor U21370 (N_21370,N_20016,N_20839);
and U21371 (N_21371,N_20057,N_20272);
and U21372 (N_21372,N_20772,N_20972);
xor U21373 (N_21373,N_20565,N_20195);
nand U21374 (N_21374,N_20868,N_20835);
or U21375 (N_21375,N_20089,N_20285);
or U21376 (N_21376,N_20112,N_20957);
or U21377 (N_21377,N_20783,N_20583);
and U21378 (N_21378,N_20920,N_20437);
and U21379 (N_21379,N_20000,N_20568);
nand U21380 (N_21380,N_20620,N_20707);
or U21381 (N_21381,N_20305,N_20698);
nand U21382 (N_21382,N_20236,N_20590);
xnor U21383 (N_21383,N_20840,N_20630);
nand U21384 (N_21384,N_20455,N_20313);
nand U21385 (N_21385,N_20712,N_20775);
or U21386 (N_21386,N_20657,N_20264);
nor U21387 (N_21387,N_20953,N_20927);
nor U21388 (N_21388,N_20417,N_20976);
and U21389 (N_21389,N_20499,N_20495);
nor U21390 (N_21390,N_20769,N_20083);
nor U21391 (N_21391,N_20324,N_20297);
xor U21392 (N_21392,N_20924,N_20445);
xor U21393 (N_21393,N_20885,N_20594);
nor U21394 (N_21394,N_20326,N_20782);
or U21395 (N_21395,N_20096,N_20694);
and U21396 (N_21396,N_20711,N_20652);
or U21397 (N_21397,N_20624,N_20211);
and U21398 (N_21398,N_20254,N_20218);
xnor U21399 (N_21399,N_20239,N_20506);
and U21400 (N_21400,N_20866,N_20750);
nor U21401 (N_21401,N_20872,N_20433);
xnor U21402 (N_21402,N_20184,N_20766);
nor U21403 (N_21403,N_20539,N_20159);
nand U21404 (N_21404,N_20643,N_20333);
xnor U21405 (N_21405,N_20312,N_20689);
and U21406 (N_21406,N_20447,N_20029);
nor U21407 (N_21407,N_20045,N_20347);
and U21408 (N_21408,N_20383,N_20877);
or U21409 (N_21409,N_20366,N_20700);
and U21410 (N_21410,N_20758,N_20756);
nor U21411 (N_21411,N_20303,N_20561);
nor U21412 (N_21412,N_20847,N_20152);
xor U21413 (N_21413,N_20082,N_20230);
nor U21414 (N_21414,N_20917,N_20855);
or U21415 (N_21415,N_20315,N_20969);
xnor U21416 (N_21416,N_20764,N_20371);
xnor U21417 (N_21417,N_20471,N_20662);
or U21418 (N_21418,N_20611,N_20110);
and U21419 (N_21419,N_20523,N_20120);
nand U21420 (N_21420,N_20474,N_20606);
or U21421 (N_21421,N_20497,N_20317);
and U21422 (N_21422,N_20667,N_20919);
xor U21423 (N_21423,N_20036,N_20348);
xnor U21424 (N_21424,N_20713,N_20942);
nand U21425 (N_21425,N_20053,N_20443);
or U21426 (N_21426,N_20836,N_20672);
nand U21427 (N_21427,N_20616,N_20048);
or U21428 (N_21428,N_20864,N_20773);
nand U21429 (N_21429,N_20381,N_20468);
or U21430 (N_21430,N_20142,N_20926);
nand U21431 (N_21431,N_20898,N_20659);
and U21432 (N_21432,N_20967,N_20959);
or U21433 (N_21433,N_20932,N_20453);
nand U21434 (N_21434,N_20273,N_20693);
nand U21435 (N_21435,N_20644,N_20716);
nor U21436 (N_21436,N_20607,N_20774);
nor U21437 (N_21437,N_20695,N_20811);
nand U21438 (N_21438,N_20493,N_20189);
nor U21439 (N_21439,N_20581,N_20524);
or U21440 (N_21440,N_20322,N_20584);
nor U21441 (N_21441,N_20735,N_20234);
and U21442 (N_21442,N_20728,N_20988);
xnor U21443 (N_21443,N_20294,N_20733);
and U21444 (N_21444,N_20310,N_20163);
nand U21445 (N_21445,N_20141,N_20286);
nand U21446 (N_21446,N_20068,N_20400);
or U21447 (N_21447,N_20489,N_20679);
nand U21448 (N_21448,N_20328,N_20933);
nor U21449 (N_21449,N_20465,N_20856);
or U21450 (N_21450,N_20491,N_20901);
xnor U21451 (N_21451,N_20394,N_20208);
nand U21452 (N_21452,N_20832,N_20871);
xor U21453 (N_21453,N_20335,N_20435);
xor U21454 (N_21454,N_20360,N_20020);
or U21455 (N_21455,N_20476,N_20589);
and U21456 (N_21456,N_20100,N_20669);
or U21457 (N_21457,N_20631,N_20200);
xnor U21458 (N_21458,N_20436,N_20237);
or U21459 (N_21459,N_20031,N_20350);
xor U21460 (N_21460,N_20060,N_20448);
nor U21461 (N_21461,N_20183,N_20355);
or U21462 (N_21462,N_20243,N_20553);
or U21463 (N_21463,N_20799,N_20375);
xor U21464 (N_21464,N_20718,N_20050);
and U21465 (N_21465,N_20656,N_20778);
nand U21466 (N_21466,N_20948,N_20372);
nor U21467 (N_21467,N_20414,N_20974);
nand U21468 (N_21468,N_20094,N_20108);
and U21469 (N_21469,N_20860,N_20859);
nor U21470 (N_21470,N_20779,N_20552);
nand U21471 (N_21471,N_20267,N_20562);
and U21472 (N_21472,N_20241,N_20500);
or U21473 (N_21473,N_20515,N_20922);
or U21474 (N_21474,N_20046,N_20140);
and U21475 (N_21475,N_20002,N_20979);
or U21476 (N_21476,N_20776,N_20091);
or U21477 (N_21477,N_20598,N_20706);
nand U21478 (N_21478,N_20232,N_20742);
or U21479 (N_21479,N_20763,N_20070);
and U21480 (N_21480,N_20608,N_20540);
and U21481 (N_21481,N_20302,N_20870);
or U21482 (N_21482,N_20420,N_20929);
xor U21483 (N_21483,N_20940,N_20886);
and U21484 (N_21484,N_20160,N_20282);
xor U21485 (N_21485,N_20770,N_20339);
xor U21486 (N_21486,N_20536,N_20011);
xor U21487 (N_21487,N_20485,N_20040);
and U21488 (N_21488,N_20280,N_20542);
nand U21489 (N_21489,N_20276,N_20527);
nand U21490 (N_21490,N_20977,N_20446);
nor U21491 (N_21491,N_20252,N_20876);
and U21492 (N_21492,N_20822,N_20516);
xor U21493 (N_21493,N_20291,N_20041);
nand U21494 (N_21494,N_20938,N_20759);
xnor U21495 (N_21495,N_20702,N_20574);
or U21496 (N_21496,N_20645,N_20440);
nand U21497 (N_21497,N_20084,N_20837);
and U21498 (N_21498,N_20846,N_20827);
nand U21499 (N_21499,N_20844,N_20605);
nor U21500 (N_21500,N_20617,N_20159);
xnor U21501 (N_21501,N_20664,N_20925);
xnor U21502 (N_21502,N_20432,N_20681);
nor U21503 (N_21503,N_20652,N_20309);
or U21504 (N_21504,N_20568,N_20523);
nand U21505 (N_21505,N_20117,N_20843);
nand U21506 (N_21506,N_20087,N_20897);
nor U21507 (N_21507,N_20904,N_20008);
xnor U21508 (N_21508,N_20967,N_20159);
nand U21509 (N_21509,N_20745,N_20177);
and U21510 (N_21510,N_20873,N_20441);
nor U21511 (N_21511,N_20294,N_20813);
and U21512 (N_21512,N_20930,N_20232);
nand U21513 (N_21513,N_20587,N_20960);
xnor U21514 (N_21514,N_20942,N_20001);
nor U21515 (N_21515,N_20262,N_20749);
nor U21516 (N_21516,N_20916,N_20196);
nor U21517 (N_21517,N_20901,N_20141);
nand U21518 (N_21518,N_20222,N_20972);
or U21519 (N_21519,N_20383,N_20948);
or U21520 (N_21520,N_20490,N_20035);
and U21521 (N_21521,N_20839,N_20696);
xnor U21522 (N_21522,N_20287,N_20234);
nor U21523 (N_21523,N_20680,N_20835);
and U21524 (N_21524,N_20955,N_20597);
xor U21525 (N_21525,N_20562,N_20683);
or U21526 (N_21526,N_20558,N_20069);
xnor U21527 (N_21527,N_20325,N_20703);
and U21528 (N_21528,N_20905,N_20665);
and U21529 (N_21529,N_20973,N_20019);
xnor U21530 (N_21530,N_20822,N_20286);
xor U21531 (N_21531,N_20314,N_20641);
and U21532 (N_21532,N_20539,N_20151);
xnor U21533 (N_21533,N_20915,N_20035);
nand U21534 (N_21534,N_20941,N_20880);
nand U21535 (N_21535,N_20846,N_20505);
or U21536 (N_21536,N_20787,N_20816);
or U21537 (N_21537,N_20418,N_20037);
nor U21538 (N_21538,N_20056,N_20667);
nand U21539 (N_21539,N_20409,N_20863);
xnor U21540 (N_21540,N_20891,N_20361);
and U21541 (N_21541,N_20974,N_20427);
and U21542 (N_21542,N_20831,N_20081);
nor U21543 (N_21543,N_20511,N_20148);
nand U21544 (N_21544,N_20304,N_20648);
or U21545 (N_21545,N_20796,N_20977);
or U21546 (N_21546,N_20089,N_20755);
or U21547 (N_21547,N_20497,N_20630);
nand U21548 (N_21548,N_20718,N_20017);
xor U21549 (N_21549,N_20237,N_20500);
xor U21550 (N_21550,N_20741,N_20887);
or U21551 (N_21551,N_20176,N_20722);
or U21552 (N_21552,N_20726,N_20438);
nand U21553 (N_21553,N_20199,N_20660);
or U21554 (N_21554,N_20528,N_20456);
and U21555 (N_21555,N_20477,N_20401);
xnor U21556 (N_21556,N_20434,N_20542);
or U21557 (N_21557,N_20736,N_20239);
or U21558 (N_21558,N_20785,N_20699);
or U21559 (N_21559,N_20307,N_20571);
xor U21560 (N_21560,N_20698,N_20279);
xor U21561 (N_21561,N_20468,N_20493);
xnor U21562 (N_21562,N_20740,N_20009);
nor U21563 (N_21563,N_20212,N_20270);
nand U21564 (N_21564,N_20599,N_20402);
and U21565 (N_21565,N_20422,N_20343);
nand U21566 (N_21566,N_20193,N_20986);
or U21567 (N_21567,N_20679,N_20742);
nand U21568 (N_21568,N_20147,N_20294);
or U21569 (N_21569,N_20481,N_20863);
and U21570 (N_21570,N_20801,N_20804);
nand U21571 (N_21571,N_20350,N_20547);
nor U21572 (N_21572,N_20688,N_20813);
nor U21573 (N_21573,N_20842,N_20693);
nor U21574 (N_21574,N_20922,N_20652);
nor U21575 (N_21575,N_20743,N_20155);
xor U21576 (N_21576,N_20090,N_20699);
xor U21577 (N_21577,N_20664,N_20733);
or U21578 (N_21578,N_20378,N_20878);
xor U21579 (N_21579,N_20944,N_20296);
nand U21580 (N_21580,N_20043,N_20171);
xor U21581 (N_21581,N_20312,N_20151);
nor U21582 (N_21582,N_20597,N_20728);
or U21583 (N_21583,N_20930,N_20306);
and U21584 (N_21584,N_20375,N_20911);
and U21585 (N_21585,N_20885,N_20392);
xnor U21586 (N_21586,N_20268,N_20185);
nor U21587 (N_21587,N_20208,N_20953);
and U21588 (N_21588,N_20539,N_20190);
or U21589 (N_21589,N_20666,N_20213);
or U21590 (N_21590,N_20626,N_20998);
nor U21591 (N_21591,N_20846,N_20702);
nand U21592 (N_21592,N_20661,N_20321);
or U21593 (N_21593,N_20851,N_20193);
nand U21594 (N_21594,N_20279,N_20113);
nand U21595 (N_21595,N_20841,N_20971);
nor U21596 (N_21596,N_20754,N_20944);
nor U21597 (N_21597,N_20277,N_20692);
and U21598 (N_21598,N_20105,N_20525);
xnor U21599 (N_21599,N_20029,N_20055);
and U21600 (N_21600,N_20206,N_20353);
nand U21601 (N_21601,N_20653,N_20624);
nor U21602 (N_21602,N_20859,N_20962);
nor U21603 (N_21603,N_20287,N_20263);
nor U21604 (N_21604,N_20060,N_20177);
or U21605 (N_21605,N_20713,N_20139);
or U21606 (N_21606,N_20676,N_20847);
and U21607 (N_21607,N_20267,N_20907);
or U21608 (N_21608,N_20147,N_20067);
or U21609 (N_21609,N_20727,N_20027);
nor U21610 (N_21610,N_20335,N_20420);
xnor U21611 (N_21611,N_20695,N_20668);
and U21612 (N_21612,N_20734,N_20648);
or U21613 (N_21613,N_20257,N_20317);
or U21614 (N_21614,N_20551,N_20078);
xor U21615 (N_21615,N_20078,N_20780);
xnor U21616 (N_21616,N_20441,N_20354);
nor U21617 (N_21617,N_20315,N_20345);
nand U21618 (N_21618,N_20443,N_20098);
nor U21619 (N_21619,N_20997,N_20741);
nor U21620 (N_21620,N_20554,N_20748);
xnor U21621 (N_21621,N_20778,N_20292);
nor U21622 (N_21622,N_20758,N_20260);
nand U21623 (N_21623,N_20640,N_20320);
and U21624 (N_21624,N_20668,N_20154);
nor U21625 (N_21625,N_20889,N_20386);
nand U21626 (N_21626,N_20171,N_20416);
or U21627 (N_21627,N_20100,N_20999);
and U21628 (N_21628,N_20677,N_20483);
and U21629 (N_21629,N_20496,N_20620);
xor U21630 (N_21630,N_20297,N_20829);
and U21631 (N_21631,N_20322,N_20437);
and U21632 (N_21632,N_20280,N_20971);
or U21633 (N_21633,N_20269,N_20599);
and U21634 (N_21634,N_20399,N_20502);
or U21635 (N_21635,N_20544,N_20164);
or U21636 (N_21636,N_20297,N_20409);
nor U21637 (N_21637,N_20545,N_20738);
nand U21638 (N_21638,N_20653,N_20722);
and U21639 (N_21639,N_20636,N_20696);
nor U21640 (N_21640,N_20451,N_20444);
nor U21641 (N_21641,N_20920,N_20316);
nor U21642 (N_21642,N_20010,N_20669);
or U21643 (N_21643,N_20669,N_20653);
and U21644 (N_21644,N_20294,N_20379);
or U21645 (N_21645,N_20481,N_20829);
or U21646 (N_21646,N_20741,N_20487);
xor U21647 (N_21647,N_20833,N_20443);
or U21648 (N_21648,N_20413,N_20732);
or U21649 (N_21649,N_20688,N_20955);
and U21650 (N_21650,N_20054,N_20664);
nor U21651 (N_21651,N_20312,N_20753);
and U21652 (N_21652,N_20630,N_20617);
or U21653 (N_21653,N_20900,N_20460);
nand U21654 (N_21654,N_20765,N_20983);
nor U21655 (N_21655,N_20564,N_20561);
nor U21656 (N_21656,N_20955,N_20524);
nand U21657 (N_21657,N_20303,N_20571);
nand U21658 (N_21658,N_20531,N_20617);
or U21659 (N_21659,N_20918,N_20003);
or U21660 (N_21660,N_20283,N_20443);
or U21661 (N_21661,N_20845,N_20523);
or U21662 (N_21662,N_20365,N_20965);
and U21663 (N_21663,N_20392,N_20039);
and U21664 (N_21664,N_20670,N_20187);
and U21665 (N_21665,N_20425,N_20209);
or U21666 (N_21666,N_20741,N_20281);
or U21667 (N_21667,N_20227,N_20758);
nand U21668 (N_21668,N_20660,N_20165);
and U21669 (N_21669,N_20509,N_20343);
or U21670 (N_21670,N_20537,N_20977);
nor U21671 (N_21671,N_20206,N_20092);
or U21672 (N_21672,N_20969,N_20677);
or U21673 (N_21673,N_20948,N_20227);
nand U21674 (N_21674,N_20380,N_20531);
xor U21675 (N_21675,N_20124,N_20835);
nor U21676 (N_21676,N_20812,N_20693);
nand U21677 (N_21677,N_20333,N_20467);
nand U21678 (N_21678,N_20529,N_20653);
nor U21679 (N_21679,N_20980,N_20145);
xor U21680 (N_21680,N_20297,N_20092);
or U21681 (N_21681,N_20626,N_20220);
nor U21682 (N_21682,N_20909,N_20590);
nor U21683 (N_21683,N_20549,N_20164);
nor U21684 (N_21684,N_20137,N_20549);
xor U21685 (N_21685,N_20625,N_20086);
nand U21686 (N_21686,N_20164,N_20200);
nor U21687 (N_21687,N_20354,N_20944);
and U21688 (N_21688,N_20913,N_20886);
nand U21689 (N_21689,N_20924,N_20079);
nand U21690 (N_21690,N_20289,N_20109);
or U21691 (N_21691,N_20446,N_20082);
and U21692 (N_21692,N_20024,N_20332);
and U21693 (N_21693,N_20357,N_20593);
and U21694 (N_21694,N_20622,N_20716);
nand U21695 (N_21695,N_20707,N_20035);
nor U21696 (N_21696,N_20357,N_20639);
nand U21697 (N_21697,N_20751,N_20007);
and U21698 (N_21698,N_20643,N_20350);
and U21699 (N_21699,N_20908,N_20946);
and U21700 (N_21700,N_20545,N_20615);
nand U21701 (N_21701,N_20860,N_20741);
nor U21702 (N_21702,N_20404,N_20494);
nor U21703 (N_21703,N_20318,N_20641);
or U21704 (N_21704,N_20353,N_20661);
nand U21705 (N_21705,N_20121,N_20402);
nor U21706 (N_21706,N_20064,N_20851);
nand U21707 (N_21707,N_20512,N_20465);
and U21708 (N_21708,N_20547,N_20117);
and U21709 (N_21709,N_20073,N_20977);
nand U21710 (N_21710,N_20503,N_20686);
nand U21711 (N_21711,N_20636,N_20857);
nand U21712 (N_21712,N_20487,N_20846);
and U21713 (N_21713,N_20309,N_20013);
and U21714 (N_21714,N_20283,N_20654);
xor U21715 (N_21715,N_20276,N_20545);
and U21716 (N_21716,N_20738,N_20664);
xnor U21717 (N_21717,N_20504,N_20638);
and U21718 (N_21718,N_20255,N_20299);
nor U21719 (N_21719,N_20457,N_20970);
or U21720 (N_21720,N_20627,N_20069);
xnor U21721 (N_21721,N_20791,N_20105);
nor U21722 (N_21722,N_20778,N_20285);
or U21723 (N_21723,N_20933,N_20002);
or U21724 (N_21724,N_20225,N_20633);
or U21725 (N_21725,N_20748,N_20871);
or U21726 (N_21726,N_20377,N_20710);
and U21727 (N_21727,N_20503,N_20459);
nand U21728 (N_21728,N_20337,N_20671);
xor U21729 (N_21729,N_20407,N_20541);
nor U21730 (N_21730,N_20385,N_20490);
nand U21731 (N_21731,N_20029,N_20536);
or U21732 (N_21732,N_20937,N_20646);
nor U21733 (N_21733,N_20117,N_20415);
and U21734 (N_21734,N_20808,N_20768);
nand U21735 (N_21735,N_20336,N_20790);
and U21736 (N_21736,N_20749,N_20560);
nor U21737 (N_21737,N_20579,N_20238);
nand U21738 (N_21738,N_20108,N_20200);
xor U21739 (N_21739,N_20003,N_20009);
xnor U21740 (N_21740,N_20621,N_20260);
xor U21741 (N_21741,N_20891,N_20894);
xnor U21742 (N_21742,N_20651,N_20831);
and U21743 (N_21743,N_20269,N_20483);
nor U21744 (N_21744,N_20985,N_20720);
or U21745 (N_21745,N_20302,N_20156);
and U21746 (N_21746,N_20824,N_20996);
nand U21747 (N_21747,N_20633,N_20709);
or U21748 (N_21748,N_20753,N_20279);
nor U21749 (N_21749,N_20559,N_20319);
nor U21750 (N_21750,N_20790,N_20553);
xor U21751 (N_21751,N_20050,N_20516);
and U21752 (N_21752,N_20429,N_20830);
or U21753 (N_21753,N_20805,N_20892);
nand U21754 (N_21754,N_20614,N_20969);
xnor U21755 (N_21755,N_20924,N_20598);
or U21756 (N_21756,N_20625,N_20177);
nor U21757 (N_21757,N_20324,N_20644);
and U21758 (N_21758,N_20702,N_20930);
and U21759 (N_21759,N_20324,N_20538);
nor U21760 (N_21760,N_20669,N_20672);
xor U21761 (N_21761,N_20895,N_20852);
nand U21762 (N_21762,N_20533,N_20808);
and U21763 (N_21763,N_20253,N_20357);
xor U21764 (N_21764,N_20598,N_20517);
nand U21765 (N_21765,N_20154,N_20931);
or U21766 (N_21766,N_20627,N_20562);
xor U21767 (N_21767,N_20147,N_20289);
nand U21768 (N_21768,N_20565,N_20572);
xor U21769 (N_21769,N_20754,N_20699);
nor U21770 (N_21770,N_20945,N_20744);
and U21771 (N_21771,N_20161,N_20665);
nor U21772 (N_21772,N_20036,N_20974);
xor U21773 (N_21773,N_20141,N_20672);
xor U21774 (N_21774,N_20461,N_20503);
nand U21775 (N_21775,N_20905,N_20415);
xor U21776 (N_21776,N_20475,N_20072);
xnor U21777 (N_21777,N_20718,N_20880);
nand U21778 (N_21778,N_20446,N_20007);
nor U21779 (N_21779,N_20959,N_20281);
nor U21780 (N_21780,N_20766,N_20261);
xor U21781 (N_21781,N_20144,N_20162);
nor U21782 (N_21782,N_20663,N_20460);
or U21783 (N_21783,N_20728,N_20075);
nand U21784 (N_21784,N_20327,N_20918);
nor U21785 (N_21785,N_20181,N_20613);
nand U21786 (N_21786,N_20819,N_20067);
nor U21787 (N_21787,N_20725,N_20749);
and U21788 (N_21788,N_20654,N_20204);
xnor U21789 (N_21789,N_20195,N_20062);
and U21790 (N_21790,N_20588,N_20160);
or U21791 (N_21791,N_20471,N_20035);
and U21792 (N_21792,N_20332,N_20957);
nand U21793 (N_21793,N_20949,N_20866);
nand U21794 (N_21794,N_20598,N_20725);
nand U21795 (N_21795,N_20580,N_20147);
xor U21796 (N_21796,N_20950,N_20445);
nand U21797 (N_21797,N_20014,N_20402);
nor U21798 (N_21798,N_20807,N_20923);
or U21799 (N_21799,N_20635,N_20813);
nand U21800 (N_21800,N_20562,N_20338);
and U21801 (N_21801,N_20869,N_20980);
nor U21802 (N_21802,N_20083,N_20147);
nand U21803 (N_21803,N_20115,N_20168);
and U21804 (N_21804,N_20154,N_20678);
nor U21805 (N_21805,N_20019,N_20312);
and U21806 (N_21806,N_20486,N_20553);
or U21807 (N_21807,N_20232,N_20666);
nand U21808 (N_21808,N_20688,N_20807);
xnor U21809 (N_21809,N_20781,N_20505);
and U21810 (N_21810,N_20180,N_20999);
nor U21811 (N_21811,N_20918,N_20575);
and U21812 (N_21812,N_20841,N_20395);
nor U21813 (N_21813,N_20735,N_20561);
or U21814 (N_21814,N_20552,N_20228);
nor U21815 (N_21815,N_20291,N_20730);
xnor U21816 (N_21816,N_20363,N_20580);
nor U21817 (N_21817,N_20060,N_20002);
or U21818 (N_21818,N_20886,N_20512);
nand U21819 (N_21819,N_20878,N_20673);
xnor U21820 (N_21820,N_20486,N_20484);
xnor U21821 (N_21821,N_20870,N_20641);
nor U21822 (N_21822,N_20904,N_20021);
or U21823 (N_21823,N_20231,N_20035);
nor U21824 (N_21824,N_20241,N_20011);
nor U21825 (N_21825,N_20632,N_20483);
nand U21826 (N_21826,N_20461,N_20613);
nand U21827 (N_21827,N_20616,N_20881);
and U21828 (N_21828,N_20820,N_20756);
nand U21829 (N_21829,N_20610,N_20848);
or U21830 (N_21830,N_20842,N_20599);
and U21831 (N_21831,N_20349,N_20795);
or U21832 (N_21832,N_20197,N_20753);
nor U21833 (N_21833,N_20139,N_20134);
nand U21834 (N_21834,N_20745,N_20812);
and U21835 (N_21835,N_20838,N_20224);
nand U21836 (N_21836,N_20206,N_20739);
xor U21837 (N_21837,N_20396,N_20204);
or U21838 (N_21838,N_20773,N_20084);
and U21839 (N_21839,N_20186,N_20324);
nor U21840 (N_21840,N_20341,N_20013);
nand U21841 (N_21841,N_20476,N_20654);
xor U21842 (N_21842,N_20981,N_20207);
and U21843 (N_21843,N_20268,N_20020);
or U21844 (N_21844,N_20749,N_20490);
nand U21845 (N_21845,N_20351,N_20373);
xnor U21846 (N_21846,N_20043,N_20310);
nor U21847 (N_21847,N_20207,N_20024);
nor U21848 (N_21848,N_20116,N_20293);
nor U21849 (N_21849,N_20440,N_20132);
nor U21850 (N_21850,N_20646,N_20029);
and U21851 (N_21851,N_20650,N_20612);
nor U21852 (N_21852,N_20281,N_20752);
nor U21853 (N_21853,N_20235,N_20702);
or U21854 (N_21854,N_20868,N_20888);
nand U21855 (N_21855,N_20217,N_20948);
or U21856 (N_21856,N_20243,N_20561);
nand U21857 (N_21857,N_20193,N_20022);
nand U21858 (N_21858,N_20390,N_20275);
or U21859 (N_21859,N_20468,N_20519);
and U21860 (N_21860,N_20705,N_20049);
nand U21861 (N_21861,N_20569,N_20457);
nand U21862 (N_21862,N_20942,N_20823);
and U21863 (N_21863,N_20799,N_20712);
nand U21864 (N_21864,N_20936,N_20587);
and U21865 (N_21865,N_20509,N_20474);
xor U21866 (N_21866,N_20714,N_20993);
and U21867 (N_21867,N_20150,N_20809);
nand U21868 (N_21868,N_20605,N_20135);
and U21869 (N_21869,N_20061,N_20560);
or U21870 (N_21870,N_20190,N_20264);
nor U21871 (N_21871,N_20300,N_20460);
and U21872 (N_21872,N_20738,N_20641);
nor U21873 (N_21873,N_20043,N_20191);
xnor U21874 (N_21874,N_20280,N_20365);
xnor U21875 (N_21875,N_20777,N_20620);
or U21876 (N_21876,N_20781,N_20432);
or U21877 (N_21877,N_20971,N_20620);
and U21878 (N_21878,N_20746,N_20242);
nor U21879 (N_21879,N_20577,N_20327);
and U21880 (N_21880,N_20002,N_20871);
nor U21881 (N_21881,N_20828,N_20091);
xnor U21882 (N_21882,N_20073,N_20388);
xnor U21883 (N_21883,N_20273,N_20513);
or U21884 (N_21884,N_20731,N_20786);
nor U21885 (N_21885,N_20237,N_20719);
nand U21886 (N_21886,N_20950,N_20843);
nor U21887 (N_21887,N_20776,N_20862);
and U21888 (N_21888,N_20231,N_20229);
nand U21889 (N_21889,N_20034,N_20123);
xnor U21890 (N_21890,N_20095,N_20370);
and U21891 (N_21891,N_20572,N_20174);
nand U21892 (N_21892,N_20872,N_20801);
nand U21893 (N_21893,N_20285,N_20747);
xor U21894 (N_21894,N_20783,N_20694);
nand U21895 (N_21895,N_20429,N_20629);
nand U21896 (N_21896,N_20399,N_20247);
nor U21897 (N_21897,N_20904,N_20465);
nor U21898 (N_21898,N_20867,N_20577);
nand U21899 (N_21899,N_20893,N_20978);
and U21900 (N_21900,N_20858,N_20167);
or U21901 (N_21901,N_20121,N_20320);
xnor U21902 (N_21902,N_20843,N_20558);
or U21903 (N_21903,N_20956,N_20273);
xnor U21904 (N_21904,N_20980,N_20057);
xor U21905 (N_21905,N_20352,N_20847);
nor U21906 (N_21906,N_20995,N_20210);
xnor U21907 (N_21907,N_20190,N_20505);
nor U21908 (N_21908,N_20301,N_20567);
xnor U21909 (N_21909,N_20228,N_20242);
nor U21910 (N_21910,N_20417,N_20126);
nor U21911 (N_21911,N_20786,N_20049);
nor U21912 (N_21912,N_20400,N_20451);
and U21913 (N_21913,N_20456,N_20344);
or U21914 (N_21914,N_20263,N_20335);
nor U21915 (N_21915,N_20831,N_20908);
nand U21916 (N_21916,N_20418,N_20034);
nor U21917 (N_21917,N_20577,N_20628);
nor U21918 (N_21918,N_20275,N_20752);
and U21919 (N_21919,N_20260,N_20003);
or U21920 (N_21920,N_20279,N_20193);
xnor U21921 (N_21921,N_20666,N_20010);
and U21922 (N_21922,N_20694,N_20482);
xor U21923 (N_21923,N_20449,N_20671);
xnor U21924 (N_21924,N_20554,N_20448);
or U21925 (N_21925,N_20103,N_20039);
xnor U21926 (N_21926,N_20766,N_20926);
and U21927 (N_21927,N_20153,N_20927);
nand U21928 (N_21928,N_20636,N_20771);
or U21929 (N_21929,N_20408,N_20773);
nor U21930 (N_21930,N_20361,N_20253);
nand U21931 (N_21931,N_20984,N_20621);
and U21932 (N_21932,N_20340,N_20706);
nand U21933 (N_21933,N_20039,N_20264);
or U21934 (N_21934,N_20914,N_20639);
nor U21935 (N_21935,N_20242,N_20872);
nor U21936 (N_21936,N_20557,N_20645);
and U21937 (N_21937,N_20916,N_20912);
or U21938 (N_21938,N_20648,N_20067);
xor U21939 (N_21939,N_20584,N_20822);
nor U21940 (N_21940,N_20555,N_20813);
nor U21941 (N_21941,N_20496,N_20898);
xor U21942 (N_21942,N_20052,N_20386);
nor U21943 (N_21943,N_20599,N_20778);
nand U21944 (N_21944,N_20217,N_20162);
nand U21945 (N_21945,N_20415,N_20551);
and U21946 (N_21946,N_20159,N_20062);
xnor U21947 (N_21947,N_20081,N_20167);
nand U21948 (N_21948,N_20532,N_20007);
xor U21949 (N_21949,N_20686,N_20188);
or U21950 (N_21950,N_20232,N_20978);
or U21951 (N_21951,N_20327,N_20210);
nand U21952 (N_21952,N_20023,N_20689);
nor U21953 (N_21953,N_20263,N_20493);
nand U21954 (N_21954,N_20847,N_20455);
nand U21955 (N_21955,N_20458,N_20629);
nor U21956 (N_21956,N_20953,N_20049);
or U21957 (N_21957,N_20108,N_20952);
and U21958 (N_21958,N_20589,N_20144);
xor U21959 (N_21959,N_20661,N_20087);
or U21960 (N_21960,N_20853,N_20031);
nor U21961 (N_21961,N_20122,N_20325);
xor U21962 (N_21962,N_20397,N_20724);
nand U21963 (N_21963,N_20375,N_20391);
or U21964 (N_21964,N_20369,N_20351);
or U21965 (N_21965,N_20399,N_20377);
or U21966 (N_21966,N_20040,N_20121);
or U21967 (N_21967,N_20493,N_20986);
nand U21968 (N_21968,N_20266,N_20080);
xnor U21969 (N_21969,N_20842,N_20817);
xor U21970 (N_21970,N_20097,N_20558);
or U21971 (N_21971,N_20804,N_20863);
nand U21972 (N_21972,N_20109,N_20766);
or U21973 (N_21973,N_20720,N_20136);
or U21974 (N_21974,N_20493,N_20013);
or U21975 (N_21975,N_20723,N_20875);
or U21976 (N_21976,N_20643,N_20844);
nor U21977 (N_21977,N_20588,N_20388);
xnor U21978 (N_21978,N_20259,N_20827);
and U21979 (N_21979,N_20608,N_20866);
or U21980 (N_21980,N_20942,N_20386);
and U21981 (N_21981,N_20479,N_20100);
nand U21982 (N_21982,N_20187,N_20496);
or U21983 (N_21983,N_20337,N_20390);
or U21984 (N_21984,N_20148,N_20988);
xnor U21985 (N_21985,N_20975,N_20452);
xnor U21986 (N_21986,N_20819,N_20324);
and U21987 (N_21987,N_20368,N_20345);
nand U21988 (N_21988,N_20699,N_20929);
and U21989 (N_21989,N_20903,N_20301);
xor U21990 (N_21990,N_20250,N_20899);
or U21991 (N_21991,N_20593,N_20396);
nor U21992 (N_21992,N_20057,N_20427);
or U21993 (N_21993,N_20255,N_20225);
nor U21994 (N_21994,N_20151,N_20383);
and U21995 (N_21995,N_20814,N_20393);
nand U21996 (N_21996,N_20120,N_20109);
or U21997 (N_21997,N_20093,N_20946);
nor U21998 (N_21998,N_20028,N_20472);
xnor U21999 (N_21999,N_20621,N_20486);
or U22000 (N_22000,N_21405,N_21996);
nor U22001 (N_22001,N_21085,N_21223);
and U22002 (N_22002,N_21566,N_21845);
or U22003 (N_22003,N_21635,N_21306);
and U22004 (N_22004,N_21354,N_21895);
nor U22005 (N_22005,N_21005,N_21203);
or U22006 (N_22006,N_21418,N_21370);
or U22007 (N_22007,N_21360,N_21526);
nand U22008 (N_22008,N_21151,N_21626);
nand U22009 (N_22009,N_21609,N_21014);
nor U22010 (N_22010,N_21066,N_21857);
or U22011 (N_22011,N_21596,N_21995);
nand U22012 (N_22012,N_21255,N_21813);
and U22013 (N_22013,N_21077,N_21161);
and U22014 (N_22014,N_21422,N_21467);
or U22015 (N_22015,N_21664,N_21634);
xnor U22016 (N_22016,N_21887,N_21239);
and U22017 (N_22017,N_21309,N_21891);
xor U22018 (N_22018,N_21070,N_21362);
nor U22019 (N_22019,N_21440,N_21160);
nor U22020 (N_22020,N_21677,N_21436);
nand U22021 (N_22021,N_21329,N_21952);
and U22022 (N_22022,N_21695,N_21682);
xor U22023 (N_22023,N_21134,N_21285);
or U22024 (N_22024,N_21651,N_21120);
and U22025 (N_22025,N_21031,N_21923);
nor U22026 (N_22026,N_21508,N_21139);
and U22027 (N_22027,N_21372,N_21876);
nand U22028 (N_22028,N_21979,N_21571);
nor U22029 (N_22029,N_21614,N_21126);
nand U22030 (N_22030,N_21373,N_21658);
or U22031 (N_22031,N_21649,N_21495);
and U22032 (N_22032,N_21917,N_21017);
nand U22033 (N_22033,N_21251,N_21043);
and U22034 (N_22034,N_21249,N_21283);
nor U22035 (N_22035,N_21789,N_21915);
nor U22036 (N_22036,N_21831,N_21096);
xnor U22037 (N_22037,N_21276,N_21844);
nand U22038 (N_22038,N_21815,N_21273);
or U22039 (N_22039,N_21140,N_21812);
or U22040 (N_22040,N_21259,N_21368);
or U22041 (N_22041,N_21172,N_21729);
nand U22042 (N_22042,N_21501,N_21973);
xnor U22043 (N_22043,N_21704,N_21650);
nand U22044 (N_22044,N_21879,N_21702);
nand U22045 (N_22045,N_21036,N_21564);
xnor U22046 (N_22046,N_21409,N_21696);
xor U22047 (N_22047,N_21859,N_21921);
nor U22048 (N_22048,N_21234,N_21950);
xnor U22049 (N_22049,N_21709,N_21594);
nor U22050 (N_22050,N_21671,N_21047);
and U22051 (N_22051,N_21459,N_21209);
or U22052 (N_22052,N_21665,N_21836);
nor U22053 (N_22053,N_21647,N_21728);
nand U22054 (N_22054,N_21941,N_21439);
nand U22055 (N_22055,N_21050,N_21073);
xnor U22056 (N_22056,N_21646,N_21639);
xor U22057 (N_22057,N_21780,N_21617);
and U22058 (N_22058,N_21456,N_21114);
nor U22059 (N_22059,N_21260,N_21178);
or U22060 (N_22060,N_21358,N_21156);
nor U22061 (N_22061,N_21794,N_21547);
nand U22062 (N_22062,N_21998,N_21592);
and U22063 (N_22063,N_21783,N_21972);
xor U22064 (N_22064,N_21074,N_21407);
or U22065 (N_22065,N_21618,N_21854);
and U22066 (N_22066,N_21154,N_21423);
nand U22067 (N_22067,N_21980,N_21174);
nor U22068 (N_22068,N_21642,N_21821);
nand U22069 (N_22069,N_21153,N_21475);
nand U22070 (N_22070,N_21395,N_21236);
nor U22071 (N_22071,N_21393,N_21039);
nor U22072 (N_22072,N_21613,N_21137);
nand U22073 (N_22073,N_21379,N_21712);
or U22074 (N_22074,N_21450,N_21270);
xor U22075 (N_22075,N_21796,N_21697);
or U22076 (N_22076,N_21324,N_21898);
or U22077 (N_22077,N_21412,N_21991);
nand U22078 (N_22078,N_21662,N_21371);
or U22079 (N_22079,N_21869,N_21563);
nor U22080 (N_22080,N_21850,N_21997);
nand U22081 (N_22081,N_21896,N_21319);
and U22082 (N_22082,N_21262,N_21087);
nand U22083 (N_22083,N_21714,N_21477);
and U22084 (N_22084,N_21337,N_21336);
xor U22085 (N_22085,N_21745,N_21725);
xor U22086 (N_22086,N_21121,N_21802);
nand U22087 (N_22087,N_21690,N_21252);
nand U22088 (N_22088,N_21335,N_21338);
nand U22089 (N_22089,N_21130,N_21949);
nor U22090 (N_22090,N_21737,N_21870);
xor U22091 (N_22091,N_21318,N_21633);
nor U22092 (N_22092,N_21602,N_21075);
xor U22093 (N_22093,N_21380,N_21930);
nand U22094 (N_22094,N_21814,N_21981);
xor U22095 (N_22095,N_21128,N_21012);
and U22096 (N_22096,N_21211,N_21663);
xnor U22097 (N_22097,N_21044,N_21914);
nand U22098 (N_22098,N_21288,N_21631);
xor U22099 (N_22099,N_21470,N_21103);
xnor U22100 (N_22100,N_21546,N_21305);
and U22101 (N_22101,N_21512,N_21046);
nand U22102 (N_22102,N_21686,N_21080);
xnor U22103 (N_22103,N_21945,N_21514);
xor U22104 (N_22104,N_21599,N_21519);
and U22105 (N_22105,N_21157,N_21143);
xnor U22106 (N_22106,N_21183,N_21976);
or U22107 (N_22107,N_21769,N_21782);
xor U22108 (N_22108,N_21570,N_21747);
xnor U22109 (N_22109,N_21559,N_21109);
xor U22110 (N_22110,N_21127,N_21629);
or U22111 (N_22111,N_21445,N_21805);
nor U22112 (N_22112,N_21927,N_21448);
nor U22113 (N_22113,N_21576,N_21684);
and U22114 (N_22114,N_21403,N_21701);
nor U22115 (N_22115,N_21391,N_21460);
and U22116 (N_22116,N_21138,N_21466);
and U22117 (N_22117,N_21839,N_21163);
and U22118 (N_22118,N_21986,N_21186);
nand U22119 (N_22119,N_21556,N_21600);
or U22120 (N_22120,N_21834,N_21291);
xnor U22121 (N_22121,N_21027,N_21451);
or U22122 (N_22122,N_21759,N_21369);
or U22123 (N_22123,N_21426,N_21666);
or U22124 (N_22124,N_21455,N_21652);
nor U22125 (N_22125,N_21253,N_21773);
xor U22126 (N_22126,N_21698,N_21971);
or U22127 (N_22127,N_21196,N_21034);
xnor U22128 (N_22128,N_21885,N_21575);
xnor U22129 (N_22129,N_21832,N_21830);
nand U22130 (N_22130,N_21731,N_21615);
and U22131 (N_22131,N_21611,N_21461);
or U22132 (N_22132,N_21889,N_21404);
nor U22133 (N_22133,N_21934,N_21800);
nor U22134 (N_22134,N_21543,N_21265);
nor U22135 (N_22135,N_21348,N_21608);
nand U22136 (N_22136,N_21607,N_21962);
nor U22137 (N_22137,N_21676,N_21940);
nor U22138 (N_22138,N_21026,N_21837);
nand U22139 (N_22139,N_21829,N_21217);
or U22140 (N_22140,N_21988,N_21261);
and U22141 (N_22141,N_21037,N_21804);
or U22142 (N_22142,N_21577,N_21247);
nor U22143 (N_22143,N_21180,N_21194);
xnor U22144 (N_22144,N_21287,N_21447);
xor U22145 (N_22145,N_21587,N_21079);
nand U22146 (N_22146,N_21340,N_21586);
or U22147 (N_22147,N_21785,N_21119);
and U22148 (N_22148,N_21562,N_21084);
and U22149 (N_22149,N_21415,N_21732);
and U22150 (N_22150,N_21421,N_21707);
xor U22151 (N_22151,N_21625,N_21083);
nor U22152 (N_22152,N_21071,N_21757);
nor U22153 (N_22153,N_21237,N_21187);
or U22154 (N_22154,N_21946,N_21484);
or U22155 (N_22155,N_21189,N_21510);
xnor U22156 (N_22156,N_21227,N_21573);
xor U22157 (N_22157,N_21094,N_21271);
or U22158 (N_22158,N_21443,N_21820);
or U22159 (N_22159,N_21622,N_21903);
xnor U22160 (N_22160,N_21905,N_21347);
xnor U22161 (N_22161,N_21656,N_21788);
nand U22162 (N_22162,N_21330,N_21533);
or U22163 (N_22163,N_21230,N_21411);
and U22164 (N_22164,N_21063,N_21406);
xor U22165 (N_22165,N_21595,N_21678);
nor U22166 (N_22166,N_21739,N_21766);
nor U22167 (N_22167,N_21169,N_21221);
xnor U22168 (N_22168,N_21758,N_21425);
and U22169 (N_22169,N_21250,N_21922);
xnor U22170 (N_22170,N_21359,N_21520);
and U22171 (N_22171,N_21301,N_21717);
and U22172 (N_22172,N_21811,N_21779);
nor U22173 (N_22173,N_21515,N_21517);
nand U22174 (N_22174,N_21888,N_21052);
nand U22175 (N_22175,N_21053,N_21144);
or U22176 (N_22176,N_21760,N_21700);
xor U22177 (N_22177,N_21269,N_21502);
nand U22178 (N_22178,N_21177,N_21378);
and U22179 (N_22179,N_21056,N_21878);
nor U22180 (N_22180,N_21244,N_21176);
xor U22181 (N_22181,N_21100,N_21105);
nand U22182 (N_22182,N_21058,N_21929);
nor U22183 (N_22183,N_21155,N_21961);
nand U22184 (N_22184,N_21699,N_21382);
or U22185 (N_22185,N_21703,N_21568);
nor U22186 (N_22186,N_21541,N_21803);
nor U22187 (N_22187,N_21311,N_21538);
or U22188 (N_22188,N_21689,N_21532);
or U22189 (N_22189,N_21746,N_21343);
nor U22190 (N_22190,N_21809,N_21478);
nand U22191 (N_22191,N_21110,N_21229);
nand U22192 (N_22192,N_21748,N_21585);
nand U22193 (N_22193,N_21706,N_21088);
nor U22194 (N_22194,N_21363,N_21220);
nor U22195 (N_22195,N_21936,N_21106);
nor U22196 (N_22196,N_21278,N_21580);
nor U22197 (N_22197,N_21414,N_21091);
nand U22198 (N_22198,N_21463,N_21241);
xor U22199 (N_22199,N_21715,N_21694);
nand U22200 (N_22200,N_21353,N_21672);
xnor U22201 (N_22201,N_21429,N_21295);
nand U22202 (N_22202,N_21375,N_21292);
nand U22203 (N_22203,N_21632,N_21300);
and U22204 (N_22204,N_21589,N_21384);
nor U22205 (N_22205,N_21205,N_21420);
xor U22206 (N_22206,N_21736,N_21925);
nand U22207 (N_22207,N_21392,N_21750);
nor U22208 (N_22208,N_21781,N_21245);
or U22209 (N_22209,N_21705,N_21493);
nor U22210 (N_22210,N_21494,N_21135);
nand U22211 (N_22211,N_21603,N_21294);
or U22212 (N_22212,N_21487,N_21619);
nand U22213 (N_22213,N_21204,N_21624);
or U22214 (N_22214,N_21835,N_21383);
nor U22215 (N_22215,N_21640,N_21099);
xnor U22216 (N_22216,N_21910,N_21457);
xnor U22217 (N_22217,N_21281,N_21932);
or U22218 (N_22218,N_21002,N_21808);
nor U22219 (N_22219,N_21317,N_21442);
and U22220 (N_22220,N_21033,N_21637);
nand U22221 (N_22221,N_21025,N_21509);
and U22222 (N_22222,N_21356,N_21978);
nor U22223 (N_22223,N_21072,N_21472);
xnor U22224 (N_22224,N_21849,N_21536);
or U22225 (N_22225,N_21955,N_21819);
xnor U22226 (N_22226,N_21385,N_21345);
and U22227 (N_22227,N_21313,N_21778);
nand U22228 (N_22228,N_21770,N_21334);
xnor U22229 (N_22229,N_21496,N_21268);
xor U22230 (N_22230,N_21145,N_21024);
nor U22231 (N_22231,N_21605,N_21673);
xnor U22232 (N_22232,N_21790,N_21965);
xor U22233 (N_22233,N_21352,N_21065);
and U22234 (N_22234,N_21549,N_21350);
and U22235 (N_22235,N_21282,N_21848);
nand U22236 (N_22236,N_21167,N_21868);
nor U22237 (N_22237,N_21093,N_21503);
xor U22238 (N_22238,N_21873,N_21967);
nor U22239 (N_22239,N_21798,N_21817);
and U22240 (N_22240,N_21751,N_21427);
xnor U22241 (N_22241,N_21799,N_21332);
nor U22242 (N_22242,N_21786,N_21628);
xnor U22243 (N_22243,N_21713,N_21222);
or U22244 (N_22244,N_21431,N_21659);
and U22245 (N_22245,N_21825,N_21548);
xnor U22246 (N_22246,N_21584,N_21302);
or U22247 (N_22247,N_21557,N_21990);
and U22248 (N_22248,N_21553,N_21567);
or U22249 (N_22249,N_21018,N_21013);
nand U22250 (N_22250,N_21544,N_21009);
xor U22251 (N_22251,N_21818,N_21851);
or U22252 (N_22252,N_21207,N_21476);
and U22253 (N_22253,N_21298,N_21938);
xor U22254 (N_22254,N_21752,N_21777);
nand U22255 (N_22255,N_21593,N_21826);
xor U22256 (N_22256,N_21726,N_21048);
and U22257 (N_22257,N_21446,N_21645);
nand U22258 (N_22258,N_21529,N_21092);
nor U22259 (N_22259,N_21911,N_21492);
nor U22260 (N_22260,N_21215,N_21734);
nand U22261 (N_22261,N_21118,N_21606);
or U22262 (N_22262,N_21892,N_21792);
nor U22263 (N_22263,N_21377,N_21454);
nand U22264 (N_22264,N_21045,N_21289);
nor U22265 (N_22265,N_21522,N_21148);
nor U22266 (N_22266,N_21333,N_21987);
and U22267 (N_22267,N_21200,N_21937);
and U22268 (N_22268,N_21280,N_21485);
nor U22269 (N_22269,N_21860,N_21504);
xnor U22270 (N_22270,N_21231,N_21149);
nor U22271 (N_22271,N_21897,N_21078);
or U22272 (N_22272,N_21875,N_21569);
or U22273 (N_22273,N_21001,N_21474);
nand U22274 (N_22274,N_21060,N_21560);
or U22275 (N_22275,N_21668,N_21660);
or U22276 (N_22276,N_21399,N_21108);
or U22277 (N_22277,N_21213,N_21840);
and U22278 (N_22278,N_21195,N_21993);
nand U22279 (N_22279,N_21267,N_21146);
nand U22280 (N_22280,N_21181,N_21555);
nand U22281 (N_22281,N_21344,N_21774);
or U22282 (N_22282,N_21081,N_21190);
nand U22283 (N_22283,N_21513,N_21428);
xnor U22284 (N_22284,N_21490,N_21051);
nor U22285 (N_22285,N_21743,N_21871);
nor U22286 (N_22286,N_21627,N_21807);
nor U22287 (N_22287,N_21068,N_21964);
and U22288 (N_22288,N_21389,N_21537);
and U22289 (N_22289,N_21685,N_21491);
or U22290 (N_22290,N_21064,N_21824);
nand U22291 (N_22291,N_21322,N_21740);
xnor U22292 (N_22292,N_21303,N_21000);
and U22293 (N_22293,N_21008,N_21424);
xnor U22294 (N_22294,N_21376,N_21838);
or U22295 (N_22295,N_21432,N_21994);
nor U22296 (N_22296,N_21097,N_21020);
or U22297 (N_22297,N_21801,N_21902);
and U22298 (N_22298,N_21880,N_21441);
and U22299 (N_22299,N_21710,N_21674);
nand U22300 (N_22300,N_21644,N_21939);
and U22301 (N_22301,N_21687,N_21386);
nor U22302 (N_22302,N_21920,N_21098);
and U22303 (N_22303,N_21974,N_21655);
nor U22304 (N_22304,N_21775,N_21489);
nor U22305 (N_22305,N_21419,N_21597);
or U22306 (N_22306,N_21842,N_21744);
xor U22307 (N_22307,N_21693,N_21396);
and U22308 (N_22308,N_21095,N_21718);
nor U22309 (N_22309,N_21133,N_21540);
nand U22310 (N_22310,N_21591,N_21787);
nand U22311 (N_22311,N_21351,N_21999);
xor U22312 (N_22312,N_21565,N_21248);
or U22313 (N_22313,N_21225,N_21458);
nand U22314 (N_22314,N_21667,N_21164);
and U22315 (N_22315,N_21956,N_21604);
xnor U22316 (N_22316,N_21681,N_21772);
xor U22317 (N_22317,N_21327,N_21122);
xor U22318 (N_22318,N_21661,N_21192);
xor U22319 (N_22319,N_21874,N_21886);
nand U22320 (N_22320,N_21453,N_21968);
xnor U22321 (N_22321,N_21756,N_21669);
nor U22322 (N_22322,N_21581,N_21928);
and U22323 (N_22323,N_21795,N_21086);
nor U22324 (N_22324,N_21198,N_21969);
nand U22325 (N_22325,N_21171,N_21111);
or U22326 (N_22326,N_21483,N_21574);
or U22327 (N_22327,N_21708,N_21308);
and U22328 (N_22328,N_21947,N_21076);
and U22329 (N_22329,N_21833,N_21355);
xnor U22330 (N_22330,N_21730,N_21400);
nand U22331 (N_22331,N_21480,N_21958);
and U22332 (N_22332,N_21004,N_21444);
nor U22333 (N_22333,N_21894,N_21312);
nand U22334 (N_22334,N_21107,N_21688);
or U22335 (N_22335,N_21638,N_21471);
nand U22336 (N_22336,N_21523,N_21497);
or U22337 (N_22337,N_21721,N_21901);
and U22338 (N_22338,N_21913,N_21410);
nor U22339 (N_22339,N_21683,N_21716);
nand U22340 (N_22340,N_21212,N_21957);
xnor U22341 (N_22341,N_21738,N_21102);
nand U22342 (N_22342,N_21636,N_21256);
nor U22343 (N_22343,N_21680,N_21881);
xor U22344 (N_22344,N_21791,N_21742);
or U22345 (N_22345,N_21904,N_21551);
and U22346 (N_22346,N_21719,N_21284);
xor U22347 (N_22347,N_21365,N_21062);
or U22348 (N_22348,N_21473,N_21188);
nor U22349 (N_22349,N_21132,N_21919);
xnor U22350 (N_22350,N_21054,N_21518);
and U22351 (N_22351,N_21893,N_21197);
nor U22352 (N_22352,N_21724,N_21019);
nand U22353 (N_22353,N_21435,N_21055);
xor U22354 (N_22354,N_21847,N_21907);
and U22355 (N_22355,N_21290,N_21390);
nand U22356 (N_22356,N_21028,N_21768);
or U22357 (N_22357,N_21011,N_21884);
xor U22358 (N_22358,N_21679,N_21479);
and U22359 (N_22359,N_21129,N_21315);
or U22360 (N_22360,N_21158,N_21583);
and U22361 (N_22361,N_21464,N_21550);
nand U22362 (N_22362,N_21654,N_21210);
xnor U22363 (N_22363,N_21170,N_21113);
or U22364 (N_22364,N_21883,N_21416);
xor U22365 (N_22365,N_21089,N_21711);
and U22366 (N_22366,N_21310,N_21528);
nor U22367 (N_22367,N_21326,N_21462);
and U22368 (N_22368,N_21727,N_21116);
and U22369 (N_22369,N_21675,N_21042);
xor U22370 (N_22370,N_21951,N_21413);
xor U22371 (N_22371,N_21816,N_21588);
nand U22372 (N_22372,N_21316,N_21612);
and U22373 (N_22373,N_21691,N_21006);
or U22374 (N_22374,N_21733,N_21437);
xnor U22375 (N_22375,N_21765,N_21924);
xor U22376 (N_22376,N_21810,N_21346);
and U22377 (N_22377,N_21219,N_21754);
nor U22378 (N_22378,N_21499,N_21401);
or U22379 (N_22379,N_21159,N_21992);
and U22380 (N_22380,N_21926,N_21349);
nor U22381 (N_22381,N_21124,N_21741);
xnor U22382 (N_22382,N_21216,N_21856);
xnor U22383 (N_22383,N_21342,N_21038);
nand U22384 (N_22384,N_21266,N_21417);
and U22385 (N_22385,N_21616,N_21906);
nand U22386 (N_22386,N_21242,N_21465);
nor U22387 (N_22387,N_21202,N_21822);
nand U22388 (N_22388,N_21142,N_21381);
nor U22389 (N_22389,N_21610,N_21975);
nand U22390 (N_22390,N_21908,N_21960);
or U22391 (N_22391,N_21147,N_21843);
or U22392 (N_22392,N_21361,N_21648);
xor U22393 (N_22393,N_21535,N_21125);
nor U22394 (N_22394,N_21985,N_21506);
nor U22395 (N_22395,N_21264,N_21670);
or U22396 (N_22396,N_21516,N_21433);
and U22397 (N_22397,N_21325,N_21846);
or U22398 (N_22398,N_21657,N_21112);
nor U22399 (N_22399,N_21175,N_21486);
and U22400 (N_22400,N_21982,N_21806);
xnor U22401 (N_22401,N_21184,N_21866);
nor U22402 (N_22402,N_21530,N_21235);
xor U22403 (N_22403,N_21943,N_21722);
xnor U22404 (N_22404,N_21304,N_21763);
and U22405 (N_22405,N_21141,N_21942);
nor U22406 (N_22406,N_21131,N_21468);
nand U22407 (N_22407,N_21021,N_21507);
nand U22408 (N_22408,N_21542,N_21953);
or U22409 (N_22409,N_21224,N_21023);
and U22410 (N_22410,N_21558,N_21525);
or U22411 (N_22411,N_21218,N_21214);
or U22412 (N_22412,N_21449,N_21314);
nor U22413 (N_22413,N_21983,N_21539);
nand U22414 (N_22414,N_21279,N_21341);
and U22415 (N_22415,N_21150,N_21293);
or U22416 (N_22416,N_21374,N_21331);
nor U22417 (N_22417,N_21959,N_21601);
and U22418 (N_22418,N_21552,N_21166);
or U22419 (N_22419,N_21388,N_21090);
or U22420 (N_22420,N_21165,N_21545);
nand U22421 (N_22421,N_21022,N_21398);
or U22422 (N_22422,N_21771,N_21841);
and U22423 (N_22423,N_21862,N_21286);
or U22424 (N_22424,N_21032,N_21339);
nand U22425 (N_22425,N_21041,N_21357);
or U22426 (N_22426,N_21630,N_21828);
xor U22427 (N_22427,N_21179,N_21935);
xor U22428 (N_22428,N_21853,N_21944);
or U22429 (N_22429,N_21057,N_21500);
or U22430 (N_22430,N_21397,N_21452);
and U22431 (N_22431,N_21877,N_21793);
nand U22432 (N_22432,N_21865,N_21572);
or U22433 (N_22433,N_21233,N_21641);
and U22434 (N_22434,N_21069,N_21394);
xnor U22435 (N_22435,N_21598,N_21931);
nor U22436 (N_22436,N_21970,N_21067);
nand U22437 (N_22437,N_21438,N_21900);
xnor U22438 (N_22438,N_21182,N_21299);
nor U22439 (N_22439,N_21890,N_21623);
nand U22440 (N_22440,N_21366,N_21199);
or U22441 (N_22441,N_21582,N_21984);
or U22442 (N_22442,N_21328,N_21408);
nand U22443 (N_22443,N_21867,N_21257);
or U22444 (N_22444,N_21482,N_21954);
xnor U22445 (N_22445,N_21367,N_21753);
or U22446 (N_22446,N_21320,N_21061);
or U22447 (N_22447,N_21864,N_21402);
and U22448 (N_22448,N_21643,N_21872);
nand U22449 (N_22449,N_21797,N_21755);
or U22450 (N_22450,N_21554,N_21007);
xor U22451 (N_22451,N_21827,N_21232);
or U22452 (N_22452,N_21933,N_21240);
xnor U22453 (N_22453,N_21162,N_21272);
nor U22454 (N_22454,N_21297,N_21498);
and U22455 (N_22455,N_21505,N_21010);
nand U22456 (N_22456,N_21123,N_21246);
nor U22457 (N_22457,N_21561,N_21321);
or U22458 (N_22458,N_21040,N_21620);
nor U22459 (N_22459,N_21916,N_21208);
or U22460 (N_22460,N_21136,N_21228);
xor U22461 (N_22461,N_21521,N_21201);
xor U22462 (N_22462,N_21059,N_21749);
or U22463 (N_22463,N_21117,N_21590);
nor U22464 (N_22464,N_21579,N_21761);
or U22465 (N_22465,N_21621,N_21764);
or U22466 (N_22466,N_21323,N_21277);
or U22467 (N_22467,N_21511,N_21852);
and U22468 (N_22468,N_21296,N_21735);
nand U22469 (N_22469,N_21254,N_21168);
and U22470 (N_22470,N_21948,N_21152);
nor U22471 (N_22471,N_21434,N_21527);
or U22472 (N_22472,N_21918,N_21966);
xnor U22473 (N_22473,N_21029,N_21692);
nor U22474 (N_22474,N_21430,N_21307);
nand U22475 (N_22475,N_21653,N_21524);
and U22476 (N_22476,N_21963,N_21115);
nor U22477 (N_22477,N_21082,N_21274);
or U22478 (N_22478,N_21015,N_21855);
and U22479 (N_22479,N_21899,N_21578);
nand U22480 (N_22480,N_21258,N_21030);
nand U22481 (N_22481,N_21912,N_21909);
nand U22482 (N_22482,N_21469,N_21767);
nand U22483 (N_22483,N_21823,N_21784);
and U22484 (N_22484,N_21989,N_21035);
xor U22485 (N_22485,N_21191,N_21364);
xor U22486 (N_22486,N_21387,N_21882);
nand U22487 (N_22487,N_21003,N_21101);
and U22488 (N_22488,N_21861,N_21173);
and U22489 (N_22489,N_21226,N_21776);
and U22490 (N_22490,N_21185,N_21762);
and U22491 (N_22491,N_21977,N_21104);
or U22492 (N_22492,N_21206,N_21238);
nor U22493 (N_22493,N_21243,N_21275);
nor U22494 (N_22494,N_21488,N_21016);
nand U22495 (N_22495,N_21049,N_21723);
and U22496 (N_22496,N_21263,N_21534);
nand U22497 (N_22497,N_21720,N_21858);
or U22498 (N_22498,N_21531,N_21863);
nand U22499 (N_22499,N_21193,N_21481);
nand U22500 (N_22500,N_21794,N_21866);
and U22501 (N_22501,N_21893,N_21761);
nor U22502 (N_22502,N_21944,N_21447);
nand U22503 (N_22503,N_21189,N_21670);
xnor U22504 (N_22504,N_21185,N_21316);
xor U22505 (N_22505,N_21017,N_21444);
nand U22506 (N_22506,N_21327,N_21345);
and U22507 (N_22507,N_21201,N_21106);
nor U22508 (N_22508,N_21214,N_21381);
xnor U22509 (N_22509,N_21200,N_21290);
xnor U22510 (N_22510,N_21694,N_21264);
or U22511 (N_22511,N_21138,N_21349);
and U22512 (N_22512,N_21372,N_21882);
or U22513 (N_22513,N_21243,N_21056);
xor U22514 (N_22514,N_21286,N_21107);
nor U22515 (N_22515,N_21811,N_21583);
or U22516 (N_22516,N_21753,N_21566);
nand U22517 (N_22517,N_21491,N_21236);
or U22518 (N_22518,N_21224,N_21807);
and U22519 (N_22519,N_21583,N_21597);
nand U22520 (N_22520,N_21172,N_21208);
or U22521 (N_22521,N_21943,N_21553);
or U22522 (N_22522,N_21626,N_21746);
nand U22523 (N_22523,N_21241,N_21840);
xor U22524 (N_22524,N_21814,N_21124);
xnor U22525 (N_22525,N_21968,N_21038);
or U22526 (N_22526,N_21021,N_21763);
nor U22527 (N_22527,N_21128,N_21888);
or U22528 (N_22528,N_21692,N_21815);
nand U22529 (N_22529,N_21150,N_21374);
nor U22530 (N_22530,N_21091,N_21799);
nor U22531 (N_22531,N_21418,N_21110);
xor U22532 (N_22532,N_21052,N_21440);
and U22533 (N_22533,N_21020,N_21782);
nor U22534 (N_22534,N_21698,N_21305);
nand U22535 (N_22535,N_21962,N_21382);
and U22536 (N_22536,N_21764,N_21628);
nor U22537 (N_22537,N_21485,N_21055);
nand U22538 (N_22538,N_21093,N_21346);
xor U22539 (N_22539,N_21501,N_21339);
xor U22540 (N_22540,N_21932,N_21927);
nor U22541 (N_22541,N_21036,N_21113);
nor U22542 (N_22542,N_21260,N_21633);
and U22543 (N_22543,N_21333,N_21812);
nand U22544 (N_22544,N_21414,N_21718);
nor U22545 (N_22545,N_21969,N_21100);
and U22546 (N_22546,N_21626,N_21775);
nand U22547 (N_22547,N_21602,N_21953);
xor U22548 (N_22548,N_21133,N_21701);
nor U22549 (N_22549,N_21058,N_21341);
and U22550 (N_22550,N_21103,N_21328);
nand U22551 (N_22551,N_21017,N_21785);
and U22552 (N_22552,N_21454,N_21786);
or U22553 (N_22553,N_21934,N_21290);
xor U22554 (N_22554,N_21495,N_21567);
or U22555 (N_22555,N_21158,N_21217);
xor U22556 (N_22556,N_21465,N_21924);
and U22557 (N_22557,N_21792,N_21224);
and U22558 (N_22558,N_21953,N_21844);
and U22559 (N_22559,N_21832,N_21772);
xor U22560 (N_22560,N_21284,N_21897);
and U22561 (N_22561,N_21889,N_21019);
nand U22562 (N_22562,N_21084,N_21716);
or U22563 (N_22563,N_21609,N_21448);
and U22564 (N_22564,N_21128,N_21380);
and U22565 (N_22565,N_21404,N_21758);
or U22566 (N_22566,N_21420,N_21295);
and U22567 (N_22567,N_21894,N_21213);
nand U22568 (N_22568,N_21734,N_21200);
nand U22569 (N_22569,N_21383,N_21983);
nor U22570 (N_22570,N_21891,N_21457);
or U22571 (N_22571,N_21166,N_21794);
nor U22572 (N_22572,N_21485,N_21486);
xor U22573 (N_22573,N_21997,N_21909);
and U22574 (N_22574,N_21313,N_21097);
or U22575 (N_22575,N_21357,N_21979);
or U22576 (N_22576,N_21765,N_21635);
nor U22577 (N_22577,N_21155,N_21376);
nor U22578 (N_22578,N_21945,N_21909);
xnor U22579 (N_22579,N_21520,N_21558);
xor U22580 (N_22580,N_21528,N_21117);
and U22581 (N_22581,N_21758,N_21849);
and U22582 (N_22582,N_21692,N_21540);
and U22583 (N_22583,N_21388,N_21340);
and U22584 (N_22584,N_21340,N_21289);
nand U22585 (N_22585,N_21568,N_21271);
and U22586 (N_22586,N_21555,N_21285);
or U22587 (N_22587,N_21582,N_21204);
nand U22588 (N_22588,N_21372,N_21157);
nand U22589 (N_22589,N_21363,N_21009);
and U22590 (N_22590,N_21292,N_21615);
or U22591 (N_22591,N_21385,N_21346);
nand U22592 (N_22592,N_21767,N_21676);
nand U22593 (N_22593,N_21142,N_21113);
and U22594 (N_22594,N_21896,N_21728);
and U22595 (N_22595,N_21447,N_21551);
nor U22596 (N_22596,N_21083,N_21461);
or U22597 (N_22597,N_21348,N_21985);
nand U22598 (N_22598,N_21137,N_21851);
or U22599 (N_22599,N_21934,N_21364);
nand U22600 (N_22600,N_21154,N_21865);
or U22601 (N_22601,N_21075,N_21860);
or U22602 (N_22602,N_21298,N_21588);
nand U22603 (N_22603,N_21156,N_21273);
xor U22604 (N_22604,N_21116,N_21659);
or U22605 (N_22605,N_21183,N_21424);
nand U22606 (N_22606,N_21314,N_21442);
nor U22607 (N_22607,N_21784,N_21597);
nor U22608 (N_22608,N_21782,N_21055);
nand U22609 (N_22609,N_21174,N_21143);
nand U22610 (N_22610,N_21555,N_21306);
nor U22611 (N_22611,N_21820,N_21533);
and U22612 (N_22612,N_21244,N_21064);
nor U22613 (N_22613,N_21759,N_21483);
nand U22614 (N_22614,N_21802,N_21666);
xnor U22615 (N_22615,N_21867,N_21764);
or U22616 (N_22616,N_21985,N_21451);
xnor U22617 (N_22617,N_21466,N_21121);
nand U22618 (N_22618,N_21632,N_21522);
nor U22619 (N_22619,N_21360,N_21470);
or U22620 (N_22620,N_21341,N_21391);
nor U22621 (N_22621,N_21982,N_21773);
nand U22622 (N_22622,N_21470,N_21429);
and U22623 (N_22623,N_21843,N_21165);
nor U22624 (N_22624,N_21840,N_21331);
and U22625 (N_22625,N_21957,N_21662);
and U22626 (N_22626,N_21217,N_21044);
nor U22627 (N_22627,N_21555,N_21148);
nand U22628 (N_22628,N_21625,N_21809);
or U22629 (N_22629,N_21131,N_21071);
and U22630 (N_22630,N_21064,N_21716);
nor U22631 (N_22631,N_21167,N_21432);
nor U22632 (N_22632,N_21148,N_21002);
or U22633 (N_22633,N_21045,N_21083);
or U22634 (N_22634,N_21906,N_21826);
nor U22635 (N_22635,N_21805,N_21498);
or U22636 (N_22636,N_21551,N_21472);
and U22637 (N_22637,N_21388,N_21017);
or U22638 (N_22638,N_21545,N_21168);
nor U22639 (N_22639,N_21189,N_21540);
and U22640 (N_22640,N_21862,N_21832);
nor U22641 (N_22641,N_21122,N_21512);
xnor U22642 (N_22642,N_21960,N_21501);
nand U22643 (N_22643,N_21538,N_21553);
and U22644 (N_22644,N_21783,N_21326);
and U22645 (N_22645,N_21678,N_21826);
nor U22646 (N_22646,N_21502,N_21091);
or U22647 (N_22647,N_21702,N_21299);
nor U22648 (N_22648,N_21150,N_21250);
or U22649 (N_22649,N_21231,N_21540);
and U22650 (N_22650,N_21881,N_21532);
nor U22651 (N_22651,N_21049,N_21464);
nor U22652 (N_22652,N_21694,N_21917);
and U22653 (N_22653,N_21766,N_21043);
or U22654 (N_22654,N_21377,N_21112);
nand U22655 (N_22655,N_21696,N_21945);
xnor U22656 (N_22656,N_21015,N_21050);
and U22657 (N_22657,N_21462,N_21769);
nor U22658 (N_22658,N_21878,N_21264);
xor U22659 (N_22659,N_21686,N_21771);
nand U22660 (N_22660,N_21892,N_21599);
or U22661 (N_22661,N_21460,N_21890);
xor U22662 (N_22662,N_21511,N_21831);
or U22663 (N_22663,N_21321,N_21697);
nand U22664 (N_22664,N_21529,N_21078);
nand U22665 (N_22665,N_21074,N_21925);
xnor U22666 (N_22666,N_21249,N_21707);
nor U22667 (N_22667,N_21394,N_21105);
or U22668 (N_22668,N_21505,N_21895);
or U22669 (N_22669,N_21302,N_21077);
nor U22670 (N_22670,N_21158,N_21577);
and U22671 (N_22671,N_21419,N_21131);
nand U22672 (N_22672,N_21765,N_21078);
or U22673 (N_22673,N_21221,N_21859);
nor U22674 (N_22674,N_21508,N_21772);
xor U22675 (N_22675,N_21749,N_21133);
and U22676 (N_22676,N_21637,N_21058);
xor U22677 (N_22677,N_21686,N_21152);
and U22678 (N_22678,N_21160,N_21331);
and U22679 (N_22679,N_21734,N_21525);
and U22680 (N_22680,N_21611,N_21712);
nand U22681 (N_22681,N_21273,N_21714);
nor U22682 (N_22682,N_21876,N_21357);
or U22683 (N_22683,N_21811,N_21599);
or U22684 (N_22684,N_21578,N_21751);
nand U22685 (N_22685,N_21057,N_21031);
or U22686 (N_22686,N_21537,N_21035);
xnor U22687 (N_22687,N_21681,N_21051);
nor U22688 (N_22688,N_21469,N_21159);
and U22689 (N_22689,N_21350,N_21703);
xnor U22690 (N_22690,N_21435,N_21602);
nor U22691 (N_22691,N_21911,N_21147);
nand U22692 (N_22692,N_21440,N_21788);
and U22693 (N_22693,N_21034,N_21083);
nand U22694 (N_22694,N_21986,N_21913);
xor U22695 (N_22695,N_21398,N_21759);
nand U22696 (N_22696,N_21214,N_21756);
nand U22697 (N_22697,N_21102,N_21048);
or U22698 (N_22698,N_21584,N_21726);
or U22699 (N_22699,N_21910,N_21255);
and U22700 (N_22700,N_21105,N_21233);
nor U22701 (N_22701,N_21430,N_21279);
or U22702 (N_22702,N_21088,N_21540);
nand U22703 (N_22703,N_21154,N_21137);
nand U22704 (N_22704,N_21328,N_21357);
xnor U22705 (N_22705,N_21447,N_21267);
and U22706 (N_22706,N_21749,N_21588);
and U22707 (N_22707,N_21413,N_21570);
nor U22708 (N_22708,N_21500,N_21697);
nor U22709 (N_22709,N_21453,N_21608);
and U22710 (N_22710,N_21977,N_21031);
and U22711 (N_22711,N_21419,N_21614);
or U22712 (N_22712,N_21236,N_21803);
nand U22713 (N_22713,N_21714,N_21361);
xor U22714 (N_22714,N_21735,N_21408);
and U22715 (N_22715,N_21600,N_21752);
or U22716 (N_22716,N_21790,N_21703);
nand U22717 (N_22717,N_21688,N_21378);
xor U22718 (N_22718,N_21287,N_21539);
or U22719 (N_22719,N_21557,N_21067);
xnor U22720 (N_22720,N_21449,N_21843);
xnor U22721 (N_22721,N_21704,N_21226);
and U22722 (N_22722,N_21843,N_21461);
nand U22723 (N_22723,N_21317,N_21792);
xnor U22724 (N_22724,N_21738,N_21844);
and U22725 (N_22725,N_21126,N_21556);
nand U22726 (N_22726,N_21698,N_21567);
nor U22727 (N_22727,N_21099,N_21769);
xnor U22728 (N_22728,N_21859,N_21136);
xor U22729 (N_22729,N_21639,N_21998);
xnor U22730 (N_22730,N_21233,N_21974);
nand U22731 (N_22731,N_21745,N_21211);
nor U22732 (N_22732,N_21714,N_21161);
and U22733 (N_22733,N_21773,N_21949);
nor U22734 (N_22734,N_21528,N_21332);
xnor U22735 (N_22735,N_21744,N_21483);
xnor U22736 (N_22736,N_21309,N_21027);
and U22737 (N_22737,N_21069,N_21906);
nor U22738 (N_22738,N_21655,N_21760);
xor U22739 (N_22739,N_21490,N_21139);
nand U22740 (N_22740,N_21451,N_21251);
nor U22741 (N_22741,N_21960,N_21761);
nor U22742 (N_22742,N_21468,N_21459);
nand U22743 (N_22743,N_21527,N_21907);
or U22744 (N_22744,N_21537,N_21426);
nor U22745 (N_22745,N_21339,N_21675);
xnor U22746 (N_22746,N_21777,N_21173);
and U22747 (N_22747,N_21660,N_21896);
xor U22748 (N_22748,N_21163,N_21329);
or U22749 (N_22749,N_21289,N_21748);
or U22750 (N_22750,N_21110,N_21046);
nor U22751 (N_22751,N_21729,N_21556);
or U22752 (N_22752,N_21432,N_21943);
and U22753 (N_22753,N_21927,N_21189);
nor U22754 (N_22754,N_21510,N_21284);
xnor U22755 (N_22755,N_21734,N_21245);
or U22756 (N_22756,N_21933,N_21548);
and U22757 (N_22757,N_21011,N_21929);
or U22758 (N_22758,N_21879,N_21063);
or U22759 (N_22759,N_21822,N_21650);
nand U22760 (N_22760,N_21512,N_21919);
xnor U22761 (N_22761,N_21642,N_21634);
nand U22762 (N_22762,N_21030,N_21292);
and U22763 (N_22763,N_21369,N_21529);
and U22764 (N_22764,N_21338,N_21588);
nor U22765 (N_22765,N_21830,N_21342);
and U22766 (N_22766,N_21094,N_21328);
or U22767 (N_22767,N_21976,N_21420);
nand U22768 (N_22768,N_21927,N_21510);
nand U22769 (N_22769,N_21586,N_21018);
xor U22770 (N_22770,N_21431,N_21876);
nor U22771 (N_22771,N_21667,N_21274);
xor U22772 (N_22772,N_21847,N_21358);
or U22773 (N_22773,N_21084,N_21325);
nand U22774 (N_22774,N_21350,N_21119);
or U22775 (N_22775,N_21860,N_21495);
or U22776 (N_22776,N_21925,N_21860);
or U22777 (N_22777,N_21243,N_21231);
and U22778 (N_22778,N_21998,N_21171);
and U22779 (N_22779,N_21998,N_21294);
nor U22780 (N_22780,N_21630,N_21463);
xnor U22781 (N_22781,N_21709,N_21063);
and U22782 (N_22782,N_21771,N_21586);
xor U22783 (N_22783,N_21445,N_21705);
nand U22784 (N_22784,N_21890,N_21183);
nand U22785 (N_22785,N_21352,N_21511);
nand U22786 (N_22786,N_21882,N_21412);
xor U22787 (N_22787,N_21951,N_21004);
or U22788 (N_22788,N_21425,N_21283);
nor U22789 (N_22789,N_21491,N_21956);
and U22790 (N_22790,N_21469,N_21781);
nand U22791 (N_22791,N_21587,N_21411);
and U22792 (N_22792,N_21271,N_21635);
or U22793 (N_22793,N_21022,N_21524);
xnor U22794 (N_22794,N_21863,N_21927);
nor U22795 (N_22795,N_21514,N_21363);
and U22796 (N_22796,N_21191,N_21077);
and U22797 (N_22797,N_21086,N_21098);
nand U22798 (N_22798,N_21028,N_21275);
xnor U22799 (N_22799,N_21159,N_21266);
nor U22800 (N_22800,N_21350,N_21474);
xnor U22801 (N_22801,N_21450,N_21362);
nor U22802 (N_22802,N_21443,N_21235);
xor U22803 (N_22803,N_21779,N_21551);
or U22804 (N_22804,N_21596,N_21395);
xor U22805 (N_22805,N_21885,N_21520);
nor U22806 (N_22806,N_21875,N_21735);
xor U22807 (N_22807,N_21699,N_21542);
nor U22808 (N_22808,N_21528,N_21103);
nor U22809 (N_22809,N_21997,N_21212);
nor U22810 (N_22810,N_21421,N_21309);
nor U22811 (N_22811,N_21459,N_21526);
nand U22812 (N_22812,N_21982,N_21041);
nand U22813 (N_22813,N_21595,N_21277);
and U22814 (N_22814,N_21402,N_21018);
nand U22815 (N_22815,N_21496,N_21108);
nor U22816 (N_22816,N_21722,N_21288);
or U22817 (N_22817,N_21094,N_21668);
nor U22818 (N_22818,N_21977,N_21112);
and U22819 (N_22819,N_21417,N_21093);
nor U22820 (N_22820,N_21102,N_21798);
nand U22821 (N_22821,N_21566,N_21569);
or U22822 (N_22822,N_21551,N_21713);
and U22823 (N_22823,N_21877,N_21432);
xor U22824 (N_22824,N_21321,N_21054);
xnor U22825 (N_22825,N_21320,N_21431);
nor U22826 (N_22826,N_21867,N_21280);
or U22827 (N_22827,N_21007,N_21059);
and U22828 (N_22828,N_21584,N_21201);
or U22829 (N_22829,N_21207,N_21490);
or U22830 (N_22830,N_21426,N_21614);
nand U22831 (N_22831,N_21919,N_21176);
nand U22832 (N_22832,N_21057,N_21992);
nor U22833 (N_22833,N_21321,N_21685);
or U22834 (N_22834,N_21365,N_21494);
nor U22835 (N_22835,N_21715,N_21024);
xnor U22836 (N_22836,N_21396,N_21277);
xor U22837 (N_22837,N_21879,N_21178);
and U22838 (N_22838,N_21682,N_21630);
and U22839 (N_22839,N_21604,N_21975);
and U22840 (N_22840,N_21977,N_21299);
and U22841 (N_22841,N_21178,N_21530);
nand U22842 (N_22842,N_21523,N_21047);
and U22843 (N_22843,N_21527,N_21942);
and U22844 (N_22844,N_21758,N_21766);
nand U22845 (N_22845,N_21603,N_21666);
nand U22846 (N_22846,N_21764,N_21652);
xor U22847 (N_22847,N_21476,N_21157);
nand U22848 (N_22848,N_21394,N_21834);
xnor U22849 (N_22849,N_21510,N_21459);
or U22850 (N_22850,N_21357,N_21400);
nor U22851 (N_22851,N_21713,N_21384);
or U22852 (N_22852,N_21126,N_21816);
xor U22853 (N_22853,N_21429,N_21111);
nor U22854 (N_22854,N_21415,N_21337);
nand U22855 (N_22855,N_21369,N_21139);
or U22856 (N_22856,N_21390,N_21323);
or U22857 (N_22857,N_21513,N_21218);
xor U22858 (N_22858,N_21859,N_21545);
nor U22859 (N_22859,N_21371,N_21773);
nor U22860 (N_22860,N_21832,N_21040);
nor U22861 (N_22861,N_21736,N_21381);
nand U22862 (N_22862,N_21655,N_21389);
xor U22863 (N_22863,N_21488,N_21165);
xnor U22864 (N_22864,N_21404,N_21658);
nand U22865 (N_22865,N_21323,N_21589);
xor U22866 (N_22866,N_21834,N_21440);
nor U22867 (N_22867,N_21784,N_21373);
nand U22868 (N_22868,N_21847,N_21382);
and U22869 (N_22869,N_21101,N_21932);
nand U22870 (N_22870,N_21210,N_21464);
xnor U22871 (N_22871,N_21709,N_21427);
xor U22872 (N_22872,N_21928,N_21213);
and U22873 (N_22873,N_21501,N_21365);
and U22874 (N_22874,N_21671,N_21545);
nor U22875 (N_22875,N_21397,N_21134);
nand U22876 (N_22876,N_21935,N_21207);
xnor U22877 (N_22877,N_21254,N_21446);
nor U22878 (N_22878,N_21210,N_21437);
nor U22879 (N_22879,N_21336,N_21086);
and U22880 (N_22880,N_21187,N_21859);
and U22881 (N_22881,N_21249,N_21025);
nor U22882 (N_22882,N_21476,N_21086);
nor U22883 (N_22883,N_21835,N_21746);
and U22884 (N_22884,N_21879,N_21635);
or U22885 (N_22885,N_21835,N_21714);
nand U22886 (N_22886,N_21657,N_21734);
and U22887 (N_22887,N_21435,N_21582);
and U22888 (N_22888,N_21862,N_21983);
nor U22889 (N_22889,N_21519,N_21414);
nor U22890 (N_22890,N_21012,N_21785);
and U22891 (N_22891,N_21283,N_21882);
nor U22892 (N_22892,N_21571,N_21434);
xor U22893 (N_22893,N_21006,N_21117);
and U22894 (N_22894,N_21698,N_21259);
xor U22895 (N_22895,N_21973,N_21976);
nand U22896 (N_22896,N_21878,N_21369);
nor U22897 (N_22897,N_21334,N_21056);
or U22898 (N_22898,N_21868,N_21464);
and U22899 (N_22899,N_21604,N_21362);
xnor U22900 (N_22900,N_21290,N_21194);
xnor U22901 (N_22901,N_21461,N_21406);
xor U22902 (N_22902,N_21196,N_21116);
nor U22903 (N_22903,N_21852,N_21065);
xor U22904 (N_22904,N_21312,N_21148);
xor U22905 (N_22905,N_21091,N_21027);
nand U22906 (N_22906,N_21708,N_21241);
or U22907 (N_22907,N_21418,N_21156);
nor U22908 (N_22908,N_21588,N_21378);
nand U22909 (N_22909,N_21850,N_21472);
nor U22910 (N_22910,N_21925,N_21906);
nand U22911 (N_22911,N_21631,N_21657);
and U22912 (N_22912,N_21854,N_21119);
xnor U22913 (N_22913,N_21693,N_21002);
nor U22914 (N_22914,N_21836,N_21125);
nor U22915 (N_22915,N_21098,N_21021);
and U22916 (N_22916,N_21920,N_21614);
or U22917 (N_22917,N_21456,N_21920);
nand U22918 (N_22918,N_21664,N_21760);
or U22919 (N_22919,N_21037,N_21959);
nor U22920 (N_22920,N_21318,N_21231);
nand U22921 (N_22921,N_21249,N_21841);
and U22922 (N_22922,N_21249,N_21868);
nor U22923 (N_22923,N_21145,N_21702);
xor U22924 (N_22924,N_21731,N_21268);
xor U22925 (N_22925,N_21745,N_21507);
nor U22926 (N_22926,N_21998,N_21320);
nand U22927 (N_22927,N_21295,N_21793);
nor U22928 (N_22928,N_21830,N_21306);
xor U22929 (N_22929,N_21302,N_21024);
and U22930 (N_22930,N_21539,N_21000);
nor U22931 (N_22931,N_21488,N_21830);
and U22932 (N_22932,N_21780,N_21650);
nand U22933 (N_22933,N_21966,N_21260);
nand U22934 (N_22934,N_21336,N_21322);
and U22935 (N_22935,N_21945,N_21568);
xnor U22936 (N_22936,N_21971,N_21194);
or U22937 (N_22937,N_21861,N_21087);
nand U22938 (N_22938,N_21682,N_21832);
and U22939 (N_22939,N_21159,N_21853);
nand U22940 (N_22940,N_21980,N_21457);
and U22941 (N_22941,N_21436,N_21540);
xor U22942 (N_22942,N_21945,N_21027);
nand U22943 (N_22943,N_21619,N_21514);
nand U22944 (N_22944,N_21762,N_21647);
nor U22945 (N_22945,N_21794,N_21441);
nor U22946 (N_22946,N_21398,N_21865);
nor U22947 (N_22947,N_21817,N_21044);
or U22948 (N_22948,N_21855,N_21883);
or U22949 (N_22949,N_21452,N_21069);
nand U22950 (N_22950,N_21136,N_21848);
and U22951 (N_22951,N_21266,N_21074);
or U22952 (N_22952,N_21598,N_21713);
nand U22953 (N_22953,N_21992,N_21539);
or U22954 (N_22954,N_21053,N_21533);
nand U22955 (N_22955,N_21431,N_21730);
nand U22956 (N_22956,N_21119,N_21339);
nor U22957 (N_22957,N_21638,N_21550);
nand U22958 (N_22958,N_21764,N_21533);
xnor U22959 (N_22959,N_21224,N_21091);
nor U22960 (N_22960,N_21347,N_21066);
xnor U22961 (N_22961,N_21528,N_21538);
xnor U22962 (N_22962,N_21433,N_21507);
and U22963 (N_22963,N_21673,N_21438);
or U22964 (N_22964,N_21562,N_21108);
nand U22965 (N_22965,N_21761,N_21126);
xnor U22966 (N_22966,N_21577,N_21411);
nor U22967 (N_22967,N_21658,N_21618);
nor U22968 (N_22968,N_21716,N_21557);
xnor U22969 (N_22969,N_21082,N_21527);
nand U22970 (N_22970,N_21864,N_21256);
or U22971 (N_22971,N_21329,N_21906);
nand U22972 (N_22972,N_21920,N_21411);
and U22973 (N_22973,N_21894,N_21476);
xnor U22974 (N_22974,N_21504,N_21653);
nor U22975 (N_22975,N_21053,N_21500);
xnor U22976 (N_22976,N_21911,N_21448);
nand U22977 (N_22977,N_21921,N_21951);
xnor U22978 (N_22978,N_21985,N_21244);
and U22979 (N_22979,N_21030,N_21518);
nand U22980 (N_22980,N_21050,N_21215);
xor U22981 (N_22981,N_21817,N_21285);
or U22982 (N_22982,N_21728,N_21246);
nor U22983 (N_22983,N_21197,N_21098);
and U22984 (N_22984,N_21639,N_21735);
nor U22985 (N_22985,N_21094,N_21220);
xor U22986 (N_22986,N_21476,N_21362);
and U22987 (N_22987,N_21789,N_21550);
nand U22988 (N_22988,N_21765,N_21688);
nand U22989 (N_22989,N_21222,N_21333);
nand U22990 (N_22990,N_21959,N_21691);
nand U22991 (N_22991,N_21338,N_21833);
nand U22992 (N_22992,N_21222,N_21535);
xnor U22993 (N_22993,N_21229,N_21551);
and U22994 (N_22994,N_21519,N_21495);
nor U22995 (N_22995,N_21302,N_21936);
xor U22996 (N_22996,N_21561,N_21734);
nor U22997 (N_22997,N_21109,N_21691);
or U22998 (N_22998,N_21776,N_21927);
xor U22999 (N_22999,N_21641,N_21933);
or U23000 (N_23000,N_22536,N_22755);
xor U23001 (N_23001,N_22740,N_22587);
xnor U23002 (N_23002,N_22836,N_22796);
nor U23003 (N_23003,N_22676,N_22935);
xnor U23004 (N_23004,N_22177,N_22631);
or U23005 (N_23005,N_22593,N_22060);
xor U23006 (N_23006,N_22698,N_22293);
and U23007 (N_23007,N_22961,N_22973);
and U23008 (N_23008,N_22366,N_22799);
nand U23009 (N_23009,N_22339,N_22699);
nor U23010 (N_23010,N_22861,N_22294);
xor U23011 (N_23011,N_22925,N_22263);
or U23012 (N_23012,N_22847,N_22137);
or U23013 (N_23013,N_22282,N_22471);
xor U23014 (N_23014,N_22360,N_22659);
nand U23015 (N_23015,N_22543,N_22645);
nor U23016 (N_23016,N_22426,N_22002);
xnor U23017 (N_23017,N_22354,N_22250);
xor U23018 (N_23018,N_22639,N_22946);
xnor U23019 (N_23019,N_22364,N_22310);
and U23020 (N_23020,N_22095,N_22372);
xor U23021 (N_23021,N_22759,N_22598);
nand U23022 (N_23022,N_22008,N_22292);
nand U23023 (N_23023,N_22070,N_22915);
and U23024 (N_23024,N_22254,N_22724);
and U23025 (N_23025,N_22790,N_22452);
nand U23026 (N_23026,N_22937,N_22330);
xor U23027 (N_23027,N_22741,N_22169);
or U23028 (N_23028,N_22154,N_22136);
nor U23029 (N_23029,N_22821,N_22375);
and U23030 (N_23030,N_22986,N_22465);
or U23031 (N_23031,N_22180,N_22212);
and U23032 (N_23032,N_22057,N_22781);
and U23033 (N_23033,N_22004,N_22776);
nand U23034 (N_23034,N_22408,N_22072);
and U23035 (N_23035,N_22810,N_22114);
and U23036 (N_23036,N_22491,N_22677);
and U23037 (N_23037,N_22457,N_22572);
or U23038 (N_23038,N_22409,N_22966);
and U23039 (N_23039,N_22780,N_22644);
nand U23040 (N_23040,N_22851,N_22733);
and U23041 (N_23041,N_22145,N_22184);
or U23042 (N_23042,N_22804,N_22530);
nor U23043 (N_23043,N_22005,N_22082);
nand U23044 (N_23044,N_22344,N_22248);
or U23045 (N_23045,N_22256,N_22305);
and U23046 (N_23046,N_22022,N_22141);
nand U23047 (N_23047,N_22328,N_22853);
and U23048 (N_23048,N_22130,N_22738);
nand U23049 (N_23049,N_22565,N_22884);
nor U23050 (N_23050,N_22578,N_22885);
nor U23051 (N_23051,N_22561,N_22899);
nor U23052 (N_23052,N_22800,N_22168);
xnor U23053 (N_23053,N_22674,N_22811);
nand U23054 (N_23054,N_22868,N_22507);
nand U23055 (N_23055,N_22871,N_22945);
or U23056 (N_23056,N_22307,N_22031);
and U23057 (N_23057,N_22662,N_22846);
or U23058 (N_23058,N_22591,N_22812);
nand U23059 (N_23059,N_22721,N_22842);
nor U23060 (N_23060,N_22423,N_22048);
xor U23061 (N_23061,N_22497,N_22350);
nand U23062 (N_23062,N_22577,N_22160);
and U23063 (N_23063,N_22316,N_22019);
xor U23064 (N_23064,N_22343,N_22594);
nand U23065 (N_23065,N_22287,N_22444);
xnor U23066 (N_23066,N_22210,N_22189);
nor U23067 (N_23067,N_22296,N_22102);
xor U23068 (N_23068,N_22261,N_22486);
nand U23069 (N_23069,N_22119,N_22363);
and U23070 (N_23070,N_22245,N_22955);
nand U23071 (N_23071,N_22762,N_22187);
and U23072 (N_23072,N_22605,N_22246);
nor U23073 (N_23073,N_22506,N_22630);
nand U23074 (N_23074,N_22850,N_22402);
nor U23075 (N_23075,N_22616,N_22394);
nand U23076 (N_23076,N_22147,N_22708);
or U23077 (N_23077,N_22167,N_22705);
or U23078 (N_23078,N_22151,N_22528);
nand U23079 (N_23079,N_22224,N_22648);
and U23080 (N_23080,N_22007,N_22139);
nor U23081 (N_23081,N_22678,N_22833);
nor U23082 (N_23082,N_22932,N_22106);
and U23083 (N_23083,N_22424,N_22830);
and U23084 (N_23084,N_22280,N_22032);
nor U23085 (N_23085,N_22844,N_22001);
nor U23086 (N_23086,N_22138,N_22226);
or U23087 (N_23087,N_22175,N_22434);
xnor U23088 (N_23088,N_22767,N_22182);
or U23089 (N_23089,N_22231,N_22099);
xor U23090 (N_23090,N_22901,N_22928);
nor U23091 (N_23091,N_22620,N_22914);
nand U23092 (N_23092,N_22275,N_22750);
xor U23093 (N_23093,N_22550,N_22100);
or U23094 (N_23094,N_22916,N_22181);
or U23095 (N_23095,N_22907,N_22390);
xnor U23096 (N_23096,N_22012,N_22586);
xnor U23097 (N_23097,N_22291,N_22027);
xor U23098 (N_23098,N_22317,N_22352);
or U23099 (N_23099,N_22065,N_22987);
nor U23100 (N_23100,N_22793,N_22969);
nand U23101 (N_23101,N_22612,N_22502);
xor U23102 (N_23102,N_22321,N_22618);
and U23103 (N_23103,N_22055,N_22123);
nand U23104 (N_23104,N_22803,N_22641);
xor U23105 (N_23105,N_22039,N_22558);
xor U23106 (N_23106,N_22746,N_22101);
and U23107 (N_23107,N_22232,N_22534);
and U23108 (N_23108,N_22881,N_22362);
or U23109 (N_23109,N_22888,N_22877);
and U23110 (N_23110,N_22237,N_22125);
nand U23111 (N_23111,N_22588,N_22655);
nand U23112 (N_23112,N_22475,N_22814);
nor U23113 (N_23113,N_22758,N_22879);
xor U23114 (N_23114,N_22538,N_22064);
xnor U23115 (N_23115,N_22459,N_22445);
xnor U23116 (N_23116,N_22665,N_22951);
or U23117 (N_23117,N_22131,N_22546);
xnor U23118 (N_23118,N_22451,N_22427);
and U23119 (N_23119,N_22503,N_22301);
or U23120 (N_23120,N_22036,N_22400);
nand U23121 (N_23121,N_22404,N_22826);
or U23122 (N_23122,N_22069,N_22893);
nand U23123 (N_23123,N_22132,N_22815);
nor U23124 (N_23124,N_22133,N_22957);
nand U23125 (N_23125,N_22083,N_22495);
or U23126 (N_23126,N_22026,N_22809);
nor U23127 (N_23127,N_22300,N_22660);
or U23128 (N_23128,N_22824,N_22202);
or U23129 (N_23129,N_22331,N_22933);
xor U23130 (N_23130,N_22149,N_22508);
or U23131 (N_23131,N_22025,N_22201);
or U23132 (N_23132,N_22993,N_22832);
nor U23133 (N_23133,N_22085,N_22484);
and U23134 (N_23134,N_22575,N_22302);
xnor U23135 (N_23135,N_22863,N_22489);
nor U23136 (N_23136,N_22121,N_22112);
and U23137 (N_23137,N_22635,N_22053);
xnor U23138 (N_23138,N_22990,N_22430);
or U23139 (N_23139,N_22941,N_22162);
or U23140 (N_23140,N_22600,N_22329);
xnor U23141 (N_23141,N_22673,N_22663);
nand U23142 (N_23142,N_22773,N_22393);
xor U23143 (N_23143,N_22870,N_22801);
nand U23144 (N_23144,N_22756,N_22564);
nand U23145 (N_23145,N_22178,N_22273);
or U23146 (N_23146,N_22757,N_22000);
or U23147 (N_23147,N_22116,N_22991);
nand U23148 (N_23148,N_22238,N_22348);
nor U23149 (N_23149,N_22504,N_22897);
or U23150 (N_23150,N_22333,N_22105);
nand U23151 (N_23151,N_22524,N_22340);
nor U23152 (N_23152,N_22488,N_22358);
xnor U23153 (N_23153,N_22140,N_22266);
nor U23154 (N_23154,N_22643,N_22518);
and U23155 (N_23155,N_22819,N_22513);
or U23156 (N_23156,N_22255,N_22464);
and U23157 (N_23157,N_22764,N_22415);
and U23158 (N_23158,N_22742,N_22373);
nor U23159 (N_23159,N_22163,N_22029);
and U23160 (N_23160,N_22240,N_22532);
nand U23161 (N_23161,N_22274,N_22469);
and U23162 (N_23162,N_22713,N_22938);
nand U23163 (N_23163,N_22999,N_22158);
or U23164 (N_23164,N_22176,N_22629);
nor U23165 (N_23165,N_22454,N_22703);
or U23166 (N_23166,N_22370,N_22671);
nand U23167 (N_23167,N_22067,N_22632);
xor U23168 (N_23168,N_22148,N_22712);
or U23169 (N_23169,N_22230,N_22802);
or U23170 (N_23170,N_22769,N_22690);
xnor U23171 (N_23171,N_22664,N_22384);
nor U23172 (N_23172,N_22869,N_22483);
nor U23173 (N_23173,N_22622,N_22604);
xnor U23174 (N_23174,N_22535,N_22144);
xnor U23175 (N_23175,N_22979,N_22960);
nand U23176 (N_23176,N_22342,N_22956);
nor U23177 (N_23177,N_22997,N_22429);
xor U23178 (N_23178,N_22944,N_22247);
or U23179 (N_23179,N_22816,N_22397);
nand U23180 (N_23180,N_22942,N_22792);
xor U23181 (N_23181,N_22921,N_22959);
or U23182 (N_23182,N_22953,N_22428);
nor U23183 (N_23183,N_22596,N_22720);
nor U23184 (N_23184,N_22441,N_22468);
nor U23185 (N_23185,N_22225,N_22267);
or U23186 (N_23186,N_22889,N_22438);
xor U23187 (N_23187,N_22368,N_22650);
nand U23188 (N_23188,N_22988,N_22418);
xnor U23189 (N_23189,N_22840,N_22875);
nor U23190 (N_23190,N_22992,N_22276);
nand U23191 (N_23191,N_22490,N_22539);
and U23192 (N_23192,N_22728,N_22387);
or U23193 (N_23193,N_22551,N_22496);
xor U23194 (N_23194,N_22311,N_22243);
or U23195 (N_23195,N_22115,N_22695);
or U23196 (N_23196,N_22980,N_22874);
xnor U23197 (N_23197,N_22549,N_22073);
xor U23198 (N_23198,N_22798,N_22545);
xor U23199 (N_23199,N_22760,N_22474);
nor U23200 (N_23200,N_22878,N_22396);
nand U23201 (N_23201,N_22011,N_22285);
xnor U23202 (N_23202,N_22215,N_22841);
xor U23203 (N_23203,N_22078,N_22185);
and U23204 (N_23204,N_22608,N_22463);
nand U23205 (N_23205,N_22763,N_22930);
nand U23206 (N_23206,N_22559,N_22753);
or U23207 (N_23207,N_22477,N_22929);
xnor U23208 (N_23208,N_22332,N_22466);
and U23209 (N_23209,N_22380,N_22817);
and U23210 (N_23210,N_22272,N_22737);
nor U23211 (N_23211,N_22376,N_22258);
or U23212 (N_23212,N_22827,N_22236);
or U23213 (N_23213,N_22917,N_22270);
or U23214 (N_23214,N_22193,N_22873);
xnor U23215 (N_23215,N_22717,N_22883);
xor U23216 (N_23216,N_22795,N_22222);
and U23217 (N_23217,N_22656,N_22843);
xor U23218 (N_23218,N_22919,N_22056);
nand U23219 (N_23219,N_22059,N_22621);
xor U23220 (N_23220,N_22096,N_22924);
nor U23221 (N_23221,N_22747,N_22820);
nand U23222 (N_23222,N_22661,N_22574);
xnor U23223 (N_23223,N_22831,N_22511);
and U23224 (N_23224,N_22619,N_22218);
or U23225 (N_23225,N_22521,N_22510);
xnor U23226 (N_23226,N_22865,N_22568);
xnor U23227 (N_23227,N_22326,N_22412);
xnor U23228 (N_23228,N_22052,N_22436);
nor U23229 (N_23229,N_22098,N_22848);
or U23230 (N_23230,N_22628,N_22239);
xor U23231 (N_23231,N_22213,N_22950);
nand U23232 (N_23232,N_22075,N_22582);
nor U23233 (N_23233,N_22963,N_22388);
nand U23234 (N_23234,N_22922,N_22516);
xor U23235 (N_23235,N_22704,N_22111);
or U23236 (N_23236,N_22345,N_22003);
or U23237 (N_23237,N_22164,N_22037);
or U23238 (N_23238,N_22143,N_22611);
and U23239 (N_23239,N_22567,N_22736);
xnor U23240 (N_23240,N_22904,N_22092);
nand U23241 (N_23241,N_22702,N_22856);
xnor U23242 (N_23242,N_22894,N_22447);
and U23243 (N_23243,N_22962,N_22989);
or U23244 (N_23244,N_22006,N_22573);
nand U23245 (N_23245,N_22241,N_22470);
and U23246 (N_23246,N_22607,N_22386);
nand U23247 (N_23247,N_22015,N_22571);
or U23248 (N_23248,N_22768,N_22984);
or U23249 (N_23249,N_22725,N_22808);
or U23250 (N_23250,N_22689,N_22028);
or U23251 (N_23251,N_22857,N_22279);
nand U23252 (N_23252,N_22207,N_22152);
xor U23253 (N_23253,N_22204,N_22336);
xor U23254 (N_23254,N_22651,N_22385);
and U23255 (N_23255,N_22739,N_22383);
xnor U23256 (N_23256,N_22880,N_22837);
and U23257 (N_23257,N_22347,N_22968);
xnor U23258 (N_23258,N_22481,N_22014);
nor U23259 (N_23259,N_22638,N_22566);
xnor U23260 (N_23260,N_22359,N_22195);
and U23261 (N_23261,N_22560,N_22669);
and U23262 (N_23262,N_22188,N_22420);
or U23263 (N_23263,N_22867,N_22043);
or U23264 (N_23264,N_22887,N_22244);
xnor U23265 (N_23265,N_22493,N_22972);
or U23266 (N_23266,N_22784,N_22533);
xor U23267 (N_23267,N_22127,N_22634);
nor U23268 (N_23268,N_22107,N_22110);
and U23269 (N_23269,N_22823,N_22526);
or U23270 (N_23270,N_22860,N_22646);
and U23271 (N_23271,N_22617,N_22200);
nor U23272 (N_23272,N_22858,N_22268);
nand U23273 (N_23273,N_22190,N_22835);
nand U23274 (N_23274,N_22461,N_22044);
nand U23275 (N_23275,N_22688,N_22892);
xor U23276 (N_23276,N_22995,N_22734);
xnor U23277 (N_23277,N_22088,N_22401);
or U23278 (N_23278,N_22023,N_22338);
xor U23279 (N_23279,N_22286,N_22652);
and U23280 (N_23280,N_22097,N_22264);
nor U23281 (N_23281,N_22174,N_22304);
nand U23282 (N_23282,N_22374,N_22233);
and U23283 (N_23283,N_22260,N_22985);
and U23284 (N_23284,N_22649,N_22437);
xnor U23285 (N_23285,N_22122,N_22080);
xnor U23286 (N_23286,N_22277,N_22523);
and U23287 (N_23287,N_22996,N_22895);
and U23288 (N_23288,N_22675,N_22252);
xnor U23289 (N_23289,N_22208,N_22449);
or U23290 (N_23290,N_22849,N_22654);
nand U23291 (N_23291,N_22642,N_22353);
and U23292 (N_23292,N_22967,N_22253);
xnor U23293 (N_23293,N_22113,N_22242);
and U23294 (N_23294,N_22766,N_22633);
and U23295 (N_23295,N_22442,N_22902);
xor U23296 (N_23296,N_22789,N_22805);
and U23297 (N_23297,N_22203,N_22179);
and U23298 (N_23298,N_22234,N_22118);
nand U23299 (N_23299,N_22308,N_22357);
nand U23300 (N_23300,N_22797,N_22926);
nor U23301 (N_23301,N_22129,N_22024);
nand U23302 (N_23302,N_22235,N_22791);
and U23303 (N_23303,N_22977,N_22525);
or U23304 (N_23304,N_22920,N_22900);
nand U23305 (N_23305,N_22682,N_22278);
and U23306 (N_23306,N_22727,N_22687);
nand U23307 (N_23307,N_22965,N_22171);
nand U23308 (N_23308,N_22975,N_22487);
nand U23309 (N_23309,N_22192,N_22787);
nand U23310 (N_23310,N_22686,N_22680);
or U23311 (N_23311,N_22084,N_22752);
or U23312 (N_23312,N_22597,N_22379);
and U23313 (N_23313,N_22954,N_22948);
nor U23314 (N_23314,N_22392,N_22462);
nand U23315 (N_23315,N_22439,N_22367);
xor U23316 (N_23316,N_22864,N_22505);
nand U23317 (N_23317,N_22498,N_22569);
nor U23318 (N_23318,N_22089,N_22081);
and U23319 (N_23319,N_22949,N_22636);
and U23320 (N_23320,N_22405,N_22198);
xnor U23321 (N_23321,N_22807,N_22288);
xnor U23322 (N_23322,N_22613,N_22299);
nand U23323 (N_23323,N_22522,N_22398);
and U23324 (N_23324,N_22480,N_22431);
nor U23325 (N_23325,N_22666,N_22590);
nand U23326 (N_23326,N_22681,N_22982);
nand U23327 (N_23327,N_22834,N_22346);
and U23328 (N_23328,N_22603,N_22259);
nor U23329 (N_23329,N_22940,N_22295);
or U23330 (N_23330,N_22411,N_22492);
nor U23331 (N_23331,N_22749,N_22369);
nand U23332 (N_23332,N_22319,N_22016);
nand U23333 (N_23333,N_22381,N_22693);
and U23334 (N_23334,N_22156,N_22013);
and U23335 (N_23335,N_22548,N_22614);
nor U23336 (N_23336,N_22045,N_22970);
xnor U23337 (N_23337,N_22606,N_22407);
nand U23338 (N_23338,N_22335,N_22217);
and U23339 (N_23339,N_22077,N_22456);
nor U23340 (N_23340,N_22049,N_22087);
nor U23341 (N_23341,N_22166,N_22010);
and U23342 (N_23342,N_22838,N_22563);
or U23343 (N_23343,N_22391,N_22269);
xor U23344 (N_23344,N_22509,N_22748);
or U23345 (N_23345,N_22153,N_22589);
nand U23346 (N_23346,N_22958,N_22806);
nand U23347 (N_23347,N_22537,N_22128);
or U23348 (N_23348,N_22126,N_22135);
nand U23349 (N_23349,N_22581,N_22774);
nand U23350 (N_23350,N_22284,N_22050);
nor U23351 (N_23351,N_22668,N_22324);
nor U23352 (N_23352,N_22934,N_22772);
nand U23353 (N_23353,N_22094,N_22104);
or U23354 (N_23354,N_22079,N_22785);
nand U23355 (N_23355,N_22124,N_22592);
nor U23356 (N_23356,N_22034,N_22964);
nand U23357 (N_23357,N_22601,N_22432);
nor U23358 (N_23358,N_22570,N_22718);
or U23359 (N_23359,N_22761,N_22378);
nand U23360 (N_23360,N_22898,N_22421);
and U23361 (N_23361,N_22891,N_22786);
xor U23362 (N_23362,N_22356,N_22625);
nor U23363 (N_23363,N_22637,N_22183);
xnor U23364 (N_23364,N_22556,N_22170);
and U23365 (N_23365,N_22251,N_22199);
nor U23366 (N_23366,N_22211,N_22765);
and U23367 (N_23367,N_22908,N_22839);
and U23368 (N_23368,N_22165,N_22209);
nand U23369 (N_23369,N_22595,N_22685);
xnor U23370 (N_23370,N_22265,N_22658);
nand U23371 (N_23371,N_22672,N_22271);
or U23372 (N_23372,N_22882,N_22779);
nor U23373 (N_23373,N_22365,N_22822);
or U23374 (N_23374,N_22377,N_22455);
nor U23375 (N_23375,N_22794,N_22544);
and U23376 (N_23376,N_22910,N_22419);
and U23377 (N_23377,N_22998,N_22872);
nor U23378 (N_23378,N_22696,N_22219);
nand U23379 (N_23379,N_22947,N_22476);
nor U23380 (N_23380,N_22541,N_22227);
nor U23381 (N_23381,N_22416,N_22775);
nor U23382 (N_23382,N_22825,N_22066);
or U23383 (N_23383,N_22290,N_22038);
or U23384 (N_23384,N_22691,N_22062);
nand U23385 (N_23385,N_22417,N_22303);
xnor U23386 (N_23386,N_22667,N_22460);
nand U23387 (N_23387,N_22479,N_22726);
and U23388 (N_23388,N_22323,N_22220);
and U23389 (N_23389,N_22754,N_22912);
xnor U23390 (N_23390,N_22086,N_22206);
nor U23391 (N_23391,N_22422,N_22197);
nor U23392 (N_23392,N_22697,N_22467);
and U23393 (N_23393,N_22076,N_22494);
or U23394 (N_23394,N_22146,N_22745);
xnor U23395 (N_23395,N_22018,N_22257);
nand U23396 (N_23396,N_22214,N_22579);
or U23397 (N_23397,N_22196,N_22042);
and U23398 (N_23398,N_22722,N_22172);
nand U23399 (N_23399,N_22054,N_22229);
and U23400 (N_23400,N_22120,N_22450);
nand U23401 (N_23401,N_22191,N_22046);
nand U23402 (N_23402,N_22657,N_22927);
nand U23403 (N_23403,N_22297,N_22653);
or U23404 (N_23404,N_22283,N_22473);
nand U23405 (N_23405,N_22173,N_22035);
and U23406 (N_23406,N_22909,N_22710);
and U23407 (N_23407,N_22472,N_22599);
xnor U23408 (N_23408,N_22281,N_22517);
nand U23409 (N_23409,N_22159,N_22782);
and U23410 (N_23410,N_22626,N_22161);
nand U23411 (N_23411,N_22583,N_22553);
xnor U23412 (N_23412,N_22425,N_22009);
xor U23413 (N_23413,N_22435,N_22216);
nor U23414 (N_23414,N_22389,N_22584);
or U23415 (N_23415,N_22047,N_22478);
or U23416 (N_23416,N_22828,N_22074);
nor U23417 (N_23417,N_22443,N_22142);
and U23418 (N_23418,N_22555,N_22406);
or U23419 (N_23419,N_22647,N_22715);
or U23420 (N_23420,N_22512,N_22731);
nand U23421 (N_23421,N_22349,N_22051);
xor U23422 (N_23422,N_22931,N_22707);
nor U23423 (N_23423,N_22552,N_22071);
nand U23424 (N_23424,N_22783,N_22923);
nand U23425 (N_23425,N_22514,N_22205);
nand U23426 (N_23426,N_22771,N_22554);
and U23427 (N_23427,N_22744,N_22318);
xnor U23428 (N_23428,N_22542,N_22557);
nand U23429 (N_23429,N_22906,N_22627);
or U23430 (N_23430,N_22482,N_22221);
and U23431 (N_23431,N_22770,N_22499);
and U23432 (N_23432,N_22440,N_22320);
nor U23433 (N_23433,N_22157,N_22041);
or U23434 (N_23434,N_22063,N_22529);
nor U23435 (N_23435,N_22943,N_22090);
xnor U23436 (N_23436,N_22413,N_22520);
nand U23437 (N_23437,N_22615,N_22640);
xnor U23438 (N_23438,N_22709,N_22433);
and U23439 (N_23439,N_22446,N_22751);
or U23440 (N_23440,N_22306,N_22194);
or U23441 (N_23441,N_22859,N_22058);
nand U23442 (N_23442,N_22976,N_22971);
and U23443 (N_23443,N_22679,N_22918);
and U23444 (N_23444,N_22983,N_22716);
nor U23445 (N_23445,N_22289,N_22351);
xor U23446 (N_23446,N_22134,N_22108);
xnor U23447 (N_23447,N_22361,N_22315);
nor U23448 (N_23448,N_22355,N_22706);
and U23449 (N_23449,N_22093,N_22610);
or U23450 (N_23450,N_22322,N_22371);
and U23451 (N_23451,N_22735,N_22911);
and U23452 (N_23452,N_22314,N_22890);
and U23453 (N_23453,N_22730,N_22030);
xnor U23454 (N_23454,N_22325,N_22684);
nand U23455 (N_23455,N_22701,N_22547);
or U23456 (N_23456,N_22341,N_22453);
nand U23457 (N_23457,N_22994,N_22519);
or U23458 (N_23458,N_22501,N_22981);
xnor U23459 (N_23459,N_22939,N_22410);
and U23460 (N_23460,N_22458,N_22852);
or U23461 (N_23461,N_22515,N_22414);
nand U23462 (N_23462,N_22714,N_22540);
nand U23463 (N_23463,N_22448,N_22818);
or U23464 (N_23464,N_22403,N_22866);
nand U23465 (N_23465,N_22813,N_22103);
or U23466 (N_23466,N_22862,N_22936);
nand U23467 (N_23467,N_22854,N_22562);
and U23468 (N_23468,N_22312,N_22623);
or U23469 (N_23469,N_22576,N_22732);
or U23470 (N_23470,N_22109,N_22585);
nand U23471 (N_23471,N_22694,N_22334);
or U23472 (N_23472,N_22778,N_22974);
nand U23473 (N_23473,N_22223,N_22021);
and U23474 (N_23474,N_22743,N_22855);
xor U23475 (N_23475,N_22903,N_22228);
and U23476 (N_23476,N_22327,N_22531);
xnor U23477 (N_23477,N_22905,N_22609);
nor U23478 (N_23478,N_22624,N_22845);
nand U23479 (N_23479,N_22952,N_22117);
nor U23480 (N_23480,N_22313,N_22091);
and U23481 (N_23481,N_22723,N_22670);
or U23482 (N_23482,N_22068,N_22683);
nand U23483 (N_23483,N_22886,N_22382);
or U23484 (N_23484,N_22298,N_22913);
nand U23485 (N_23485,N_22700,N_22150);
nor U23486 (N_23486,N_22033,N_22017);
and U23487 (N_23487,N_22337,N_22186);
and U23488 (N_23488,N_22876,N_22580);
nor U23489 (N_23489,N_22788,N_22040);
xor U23490 (N_23490,N_22485,N_22399);
or U23491 (N_23491,N_22020,N_22500);
nand U23492 (N_23492,N_22692,N_22729);
nor U23493 (N_23493,N_22309,N_22719);
and U23494 (N_23494,N_22777,N_22249);
nor U23495 (N_23495,N_22061,N_22262);
nor U23496 (N_23496,N_22602,N_22829);
or U23497 (N_23497,N_22978,N_22527);
and U23498 (N_23498,N_22395,N_22711);
nand U23499 (N_23499,N_22155,N_22896);
nand U23500 (N_23500,N_22387,N_22536);
or U23501 (N_23501,N_22812,N_22624);
or U23502 (N_23502,N_22426,N_22579);
nand U23503 (N_23503,N_22963,N_22419);
and U23504 (N_23504,N_22273,N_22882);
and U23505 (N_23505,N_22043,N_22190);
nor U23506 (N_23506,N_22773,N_22780);
nor U23507 (N_23507,N_22488,N_22185);
nor U23508 (N_23508,N_22339,N_22648);
or U23509 (N_23509,N_22313,N_22083);
nand U23510 (N_23510,N_22692,N_22246);
and U23511 (N_23511,N_22610,N_22333);
xnor U23512 (N_23512,N_22059,N_22675);
and U23513 (N_23513,N_22465,N_22177);
xor U23514 (N_23514,N_22998,N_22623);
and U23515 (N_23515,N_22767,N_22800);
nand U23516 (N_23516,N_22317,N_22350);
nor U23517 (N_23517,N_22972,N_22164);
and U23518 (N_23518,N_22592,N_22338);
nor U23519 (N_23519,N_22312,N_22013);
xor U23520 (N_23520,N_22800,N_22518);
nor U23521 (N_23521,N_22394,N_22107);
and U23522 (N_23522,N_22627,N_22556);
or U23523 (N_23523,N_22609,N_22344);
nor U23524 (N_23524,N_22168,N_22006);
or U23525 (N_23525,N_22543,N_22632);
or U23526 (N_23526,N_22428,N_22858);
nand U23527 (N_23527,N_22653,N_22673);
nor U23528 (N_23528,N_22843,N_22403);
nand U23529 (N_23529,N_22142,N_22340);
nor U23530 (N_23530,N_22450,N_22614);
nor U23531 (N_23531,N_22581,N_22481);
nand U23532 (N_23532,N_22412,N_22111);
and U23533 (N_23533,N_22512,N_22457);
or U23534 (N_23534,N_22860,N_22827);
nand U23535 (N_23535,N_22594,N_22097);
nor U23536 (N_23536,N_22181,N_22159);
nor U23537 (N_23537,N_22770,N_22507);
nand U23538 (N_23538,N_22875,N_22020);
nor U23539 (N_23539,N_22515,N_22116);
xnor U23540 (N_23540,N_22948,N_22401);
nand U23541 (N_23541,N_22717,N_22139);
xor U23542 (N_23542,N_22351,N_22223);
xor U23543 (N_23543,N_22664,N_22258);
xor U23544 (N_23544,N_22183,N_22252);
nor U23545 (N_23545,N_22175,N_22663);
or U23546 (N_23546,N_22172,N_22490);
xnor U23547 (N_23547,N_22595,N_22257);
nor U23548 (N_23548,N_22785,N_22879);
nor U23549 (N_23549,N_22892,N_22261);
nor U23550 (N_23550,N_22353,N_22733);
nor U23551 (N_23551,N_22359,N_22987);
or U23552 (N_23552,N_22817,N_22540);
or U23553 (N_23553,N_22572,N_22292);
nor U23554 (N_23554,N_22381,N_22256);
xor U23555 (N_23555,N_22002,N_22005);
nor U23556 (N_23556,N_22521,N_22941);
and U23557 (N_23557,N_22704,N_22964);
nand U23558 (N_23558,N_22257,N_22484);
xnor U23559 (N_23559,N_22817,N_22937);
nand U23560 (N_23560,N_22280,N_22446);
and U23561 (N_23561,N_22090,N_22828);
xor U23562 (N_23562,N_22109,N_22077);
nor U23563 (N_23563,N_22426,N_22918);
nor U23564 (N_23564,N_22403,N_22544);
nor U23565 (N_23565,N_22240,N_22849);
or U23566 (N_23566,N_22782,N_22922);
nand U23567 (N_23567,N_22888,N_22328);
nor U23568 (N_23568,N_22967,N_22122);
nor U23569 (N_23569,N_22973,N_22579);
and U23570 (N_23570,N_22113,N_22193);
nand U23571 (N_23571,N_22972,N_22027);
or U23572 (N_23572,N_22431,N_22589);
and U23573 (N_23573,N_22073,N_22432);
or U23574 (N_23574,N_22654,N_22153);
xor U23575 (N_23575,N_22197,N_22801);
nor U23576 (N_23576,N_22916,N_22680);
nor U23577 (N_23577,N_22919,N_22538);
nor U23578 (N_23578,N_22539,N_22737);
nand U23579 (N_23579,N_22637,N_22572);
nor U23580 (N_23580,N_22191,N_22725);
nor U23581 (N_23581,N_22352,N_22407);
and U23582 (N_23582,N_22758,N_22235);
and U23583 (N_23583,N_22986,N_22816);
and U23584 (N_23584,N_22742,N_22300);
nor U23585 (N_23585,N_22314,N_22799);
nor U23586 (N_23586,N_22113,N_22350);
nand U23587 (N_23587,N_22050,N_22557);
and U23588 (N_23588,N_22895,N_22900);
or U23589 (N_23589,N_22970,N_22474);
nor U23590 (N_23590,N_22562,N_22571);
nand U23591 (N_23591,N_22513,N_22079);
or U23592 (N_23592,N_22901,N_22387);
or U23593 (N_23593,N_22970,N_22978);
and U23594 (N_23594,N_22748,N_22964);
xnor U23595 (N_23595,N_22088,N_22915);
nor U23596 (N_23596,N_22402,N_22909);
nand U23597 (N_23597,N_22939,N_22174);
or U23598 (N_23598,N_22591,N_22283);
xnor U23599 (N_23599,N_22412,N_22062);
xnor U23600 (N_23600,N_22141,N_22920);
nor U23601 (N_23601,N_22831,N_22923);
xnor U23602 (N_23602,N_22052,N_22217);
or U23603 (N_23603,N_22424,N_22502);
or U23604 (N_23604,N_22778,N_22054);
and U23605 (N_23605,N_22899,N_22346);
xnor U23606 (N_23606,N_22345,N_22479);
and U23607 (N_23607,N_22351,N_22669);
nand U23608 (N_23608,N_22640,N_22912);
or U23609 (N_23609,N_22106,N_22032);
or U23610 (N_23610,N_22508,N_22736);
nand U23611 (N_23611,N_22507,N_22757);
nand U23612 (N_23612,N_22292,N_22591);
or U23613 (N_23613,N_22731,N_22966);
or U23614 (N_23614,N_22158,N_22368);
and U23615 (N_23615,N_22484,N_22037);
xor U23616 (N_23616,N_22573,N_22214);
nor U23617 (N_23617,N_22284,N_22979);
nand U23618 (N_23618,N_22238,N_22436);
nand U23619 (N_23619,N_22193,N_22254);
and U23620 (N_23620,N_22245,N_22674);
xnor U23621 (N_23621,N_22463,N_22291);
and U23622 (N_23622,N_22482,N_22340);
and U23623 (N_23623,N_22626,N_22015);
and U23624 (N_23624,N_22387,N_22319);
or U23625 (N_23625,N_22792,N_22245);
nand U23626 (N_23626,N_22266,N_22771);
nor U23627 (N_23627,N_22840,N_22369);
and U23628 (N_23628,N_22949,N_22077);
and U23629 (N_23629,N_22475,N_22360);
and U23630 (N_23630,N_22173,N_22352);
and U23631 (N_23631,N_22374,N_22232);
xnor U23632 (N_23632,N_22227,N_22158);
nand U23633 (N_23633,N_22252,N_22977);
xnor U23634 (N_23634,N_22027,N_22365);
nand U23635 (N_23635,N_22604,N_22873);
xnor U23636 (N_23636,N_22327,N_22514);
and U23637 (N_23637,N_22661,N_22643);
and U23638 (N_23638,N_22055,N_22878);
nand U23639 (N_23639,N_22581,N_22637);
nand U23640 (N_23640,N_22876,N_22954);
and U23641 (N_23641,N_22002,N_22069);
nand U23642 (N_23642,N_22421,N_22415);
xnor U23643 (N_23643,N_22112,N_22819);
xnor U23644 (N_23644,N_22501,N_22991);
and U23645 (N_23645,N_22598,N_22930);
and U23646 (N_23646,N_22985,N_22207);
or U23647 (N_23647,N_22337,N_22742);
and U23648 (N_23648,N_22099,N_22566);
or U23649 (N_23649,N_22261,N_22076);
xor U23650 (N_23650,N_22340,N_22990);
and U23651 (N_23651,N_22826,N_22146);
and U23652 (N_23652,N_22590,N_22348);
nand U23653 (N_23653,N_22958,N_22083);
or U23654 (N_23654,N_22842,N_22679);
xnor U23655 (N_23655,N_22362,N_22661);
nand U23656 (N_23656,N_22675,N_22890);
or U23657 (N_23657,N_22785,N_22886);
or U23658 (N_23658,N_22868,N_22409);
nand U23659 (N_23659,N_22198,N_22706);
nor U23660 (N_23660,N_22838,N_22658);
and U23661 (N_23661,N_22037,N_22222);
and U23662 (N_23662,N_22071,N_22419);
nor U23663 (N_23663,N_22473,N_22516);
nor U23664 (N_23664,N_22087,N_22616);
nor U23665 (N_23665,N_22389,N_22138);
nand U23666 (N_23666,N_22747,N_22106);
nand U23667 (N_23667,N_22617,N_22609);
or U23668 (N_23668,N_22269,N_22871);
and U23669 (N_23669,N_22962,N_22185);
nor U23670 (N_23670,N_22341,N_22983);
nand U23671 (N_23671,N_22868,N_22914);
nor U23672 (N_23672,N_22188,N_22661);
nor U23673 (N_23673,N_22480,N_22788);
or U23674 (N_23674,N_22281,N_22219);
xnor U23675 (N_23675,N_22860,N_22120);
xor U23676 (N_23676,N_22321,N_22975);
nor U23677 (N_23677,N_22093,N_22324);
xor U23678 (N_23678,N_22638,N_22308);
nand U23679 (N_23679,N_22188,N_22298);
or U23680 (N_23680,N_22307,N_22576);
or U23681 (N_23681,N_22151,N_22106);
nand U23682 (N_23682,N_22612,N_22777);
xnor U23683 (N_23683,N_22942,N_22687);
xor U23684 (N_23684,N_22016,N_22716);
nand U23685 (N_23685,N_22330,N_22096);
or U23686 (N_23686,N_22900,N_22632);
nor U23687 (N_23687,N_22684,N_22490);
xnor U23688 (N_23688,N_22896,N_22578);
nor U23689 (N_23689,N_22568,N_22178);
or U23690 (N_23690,N_22447,N_22317);
nand U23691 (N_23691,N_22306,N_22043);
and U23692 (N_23692,N_22365,N_22565);
or U23693 (N_23693,N_22907,N_22763);
nor U23694 (N_23694,N_22980,N_22707);
xor U23695 (N_23695,N_22816,N_22894);
xnor U23696 (N_23696,N_22704,N_22092);
or U23697 (N_23697,N_22310,N_22751);
and U23698 (N_23698,N_22990,N_22900);
and U23699 (N_23699,N_22793,N_22650);
nor U23700 (N_23700,N_22679,N_22284);
nor U23701 (N_23701,N_22683,N_22224);
nor U23702 (N_23702,N_22526,N_22818);
xnor U23703 (N_23703,N_22584,N_22964);
or U23704 (N_23704,N_22283,N_22543);
or U23705 (N_23705,N_22186,N_22090);
and U23706 (N_23706,N_22612,N_22554);
or U23707 (N_23707,N_22067,N_22432);
nor U23708 (N_23708,N_22753,N_22198);
nor U23709 (N_23709,N_22116,N_22946);
nor U23710 (N_23710,N_22120,N_22739);
nor U23711 (N_23711,N_22582,N_22156);
xor U23712 (N_23712,N_22747,N_22619);
xor U23713 (N_23713,N_22253,N_22526);
and U23714 (N_23714,N_22889,N_22733);
or U23715 (N_23715,N_22727,N_22891);
and U23716 (N_23716,N_22143,N_22882);
nor U23717 (N_23717,N_22260,N_22843);
xor U23718 (N_23718,N_22753,N_22097);
nor U23719 (N_23719,N_22772,N_22392);
and U23720 (N_23720,N_22733,N_22124);
xor U23721 (N_23721,N_22098,N_22694);
nand U23722 (N_23722,N_22031,N_22296);
nor U23723 (N_23723,N_22954,N_22990);
nand U23724 (N_23724,N_22317,N_22309);
or U23725 (N_23725,N_22455,N_22391);
nand U23726 (N_23726,N_22413,N_22326);
nand U23727 (N_23727,N_22637,N_22937);
xnor U23728 (N_23728,N_22495,N_22373);
nand U23729 (N_23729,N_22161,N_22032);
xor U23730 (N_23730,N_22063,N_22181);
nor U23731 (N_23731,N_22663,N_22714);
nand U23732 (N_23732,N_22912,N_22650);
xnor U23733 (N_23733,N_22674,N_22626);
and U23734 (N_23734,N_22191,N_22929);
or U23735 (N_23735,N_22823,N_22925);
and U23736 (N_23736,N_22266,N_22259);
nand U23737 (N_23737,N_22128,N_22213);
nor U23738 (N_23738,N_22521,N_22434);
xnor U23739 (N_23739,N_22271,N_22559);
nor U23740 (N_23740,N_22998,N_22259);
nand U23741 (N_23741,N_22920,N_22510);
nand U23742 (N_23742,N_22315,N_22342);
xnor U23743 (N_23743,N_22620,N_22995);
or U23744 (N_23744,N_22508,N_22350);
or U23745 (N_23745,N_22692,N_22030);
xnor U23746 (N_23746,N_22735,N_22956);
or U23747 (N_23747,N_22620,N_22289);
and U23748 (N_23748,N_22188,N_22384);
and U23749 (N_23749,N_22360,N_22230);
or U23750 (N_23750,N_22018,N_22087);
nand U23751 (N_23751,N_22694,N_22470);
xor U23752 (N_23752,N_22809,N_22623);
nor U23753 (N_23753,N_22345,N_22202);
and U23754 (N_23754,N_22786,N_22283);
xor U23755 (N_23755,N_22365,N_22452);
xor U23756 (N_23756,N_22554,N_22459);
nor U23757 (N_23757,N_22640,N_22286);
nand U23758 (N_23758,N_22558,N_22319);
xnor U23759 (N_23759,N_22604,N_22188);
or U23760 (N_23760,N_22718,N_22395);
or U23761 (N_23761,N_22794,N_22605);
nand U23762 (N_23762,N_22570,N_22574);
xor U23763 (N_23763,N_22419,N_22559);
and U23764 (N_23764,N_22975,N_22263);
xnor U23765 (N_23765,N_22575,N_22226);
and U23766 (N_23766,N_22824,N_22519);
nand U23767 (N_23767,N_22013,N_22930);
and U23768 (N_23768,N_22147,N_22076);
and U23769 (N_23769,N_22861,N_22599);
and U23770 (N_23770,N_22873,N_22785);
xor U23771 (N_23771,N_22614,N_22825);
and U23772 (N_23772,N_22438,N_22728);
nand U23773 (N_23773,N_22721,N_22681);
nor U23774 (N_23774,N_22035,N_22776);
nor U23775 (N_23775,N_22362,N_22605);
and U23776 (N_23776,N_22929,N_22112);
nor U23777 (N_23777,N_22825,N_22352);
and U23778 (N_23778,N_22271,N_22445);
and U23779 (N_23779,N_22898,N_22082);
and U23780 (N_23780,N_22652,N_22810);
and U23781 (N_23781,N_22030,N_22576);
nand U23782 (N_23782,N_22922,N_22662);
and U23783 (N_23783,N_22410,N_22648);
or U23784 (N_23784,N_22034,N_22056);
and U23785 (N_23785,N_22562,N_22416);
nor U23786 (N_23786,N_22813,N_22451);
nand U23787 (N_23787,N_22466,N_22349);
and U23788 (N_23788,N_22223,N_22091);
nand U23789 (N_23789,N_22984,N_22740);
xnor U23790 (N_23790,N_22951,N_22615);
nor U23791 (N_23791,N_22434,N_22546);
and U23792 (N_23792,N_22271,N_22314);
xor U23793 (N_23793,N_22155,N_22718);
and U23794 (N_23794,N_22008,N_22635);
and U23795 (N_23795,N_22895,N_22609);
or U23796 (N_23796,N_22133,N_22233);
nand U23797 (N_23797,N_22324,N_22050);
and U23798 (N_23798,N_22840,N_22609);
nand U23799 (N_23799,N_22291,N_22621);
nor U23800 (N_23800,N_22676,N_22284);
xor U23801 (N_23801,N_22863,N_22368);
and U23802 (N_23802,N_22673,N_22867);
nor U23803 (N_23803,N_22971,N_22701);
xnor U23804 (N_23804,N_22690,N_22548);
and U23805 (N_23805,N_22012,N_22062);
and U23806 (N_23806,N_22339,N_22204);
nor U23807 (N_23807,N_22720,N_22601);
or U23808 (N_23808,N_22880,N_22851);
or U23809 (N_23809,N_22293,N_22279);
xor U23810 (N_23810,N_22907,N_22531);
xnor U23811 (N_23811,N_22519,N_22225);
or U23812 (N_23812,N_22039,N_22071);
or U23813 (N_23813,N_22313,N_22017);
or U23814 (N_23814,N_22063,N_22137);
xnor U23815 (N_23815,N_22942,N_22961);
nand U23816 (N_23816,N_22609,N_22241);
or U23817 (N_23817,N_22778,N_22932);
nor U23818 (N_23818,N_22319,N_22699);
nor U23819 (N_23819,N_22824,N_22804);
xor U23820 (N_23820,N_22594,N_22980);
nand U23821 (N_23821,N_22081,N_22155);
nor U23822 (N_23822,N_22559,N_22459);
or U23823 (N_23823,N_22844,N_22060);
or U23824 (N_23824,N_22901,N_22062);
or U23825 (N_23825,N_22599,N_22595);
nand U23826 (N_23826,N_22955,N_22333);
or U23827 (N_23827,N_22375,N_22852);
nor U23828 (N_23828,N_22029,N_22252);
nor U23829 (N_23829,N_22142,N_22892);
and U23830 (N_23830,N_22576,N_22540);
and U23831 (N_23831,N_22751,N_22775);
or U23832 (N_23832,N_22252,N_22378);
and U23833 (N_23833,N_22346,N_22150);
and U23834 (N_23834,N_22667,N_22885);
and U23835 (N_23835,N_22754,N_22364);
or U23836 (N_23836,N_22732,N_22022);
or U23837 (N_23837,N_22113,N_22439);
xor U23838 (N_23838,N_22616,N_22558);
nor U23839 (N_23839,N_22109,N_22973);
or U23840 (N_23840,N_22732,N_22240);
nand U23841 (N_23841,N_22470,N_22293);
nand U23842 (N_23842,N_22694,N_22589);
xor U23843 (N_23843,N_22894,N_22703);
or U23844 (N_23844,N_22435,N_22082);
or U23845 (N_23845,N_22039,N_22771);
nand U23846 (N_23846,N_22026,N_22530);
nor U23847 (N_23847,N_22733,N_22219);
or U23848 (N_23848,N_22300,N_22835);
and U23849 (N_23849,N_22281,N_22004);
xnor U23850 (N_23850,N_22953,N_22666);
nor U23851 (N_23851,N_22587,N_22164);
and U23852 (N_23852,N_22033,N_22438);
xor U23853 (N_23853,N_22430,N_22690);
xnor U23854 (N_23854,N_22869,N_22818);
nand U23855 (N_23855,N_22264,N_22530);
nor U23856 (N_23856,N_22284,N_22636);
and U23857 (N_23857,N_22649,N_22191);
xnor U23858 (N_23858,N_22338,N_22352);
nand U23859 (N_23859,N_22434,N_22444);
or U23860 (N_23860,N_22026,N_22396);
nand U23861 (N_23861,N_22739,N_22434);
and U23862 (N_23862,N_22629,N_22092);
and U23863 (N_23863,N_22848,N_22368);
nand U23864 (N_23864,N_22366,N_22012);
nand U23865 (N_23865,N_22372,N_22120);
and U23866 (N_23866,N_22162,N_22286);
nand U23867 (N_23867,N_22304,N_22789);
nor U23868 (N_23868,N_22956,N_22830);
nor U23869 (N_23869,N_22856,N_22965);
or U23870 (N_23870,N_22913,N_22514);
nand U23871 (N_23871,N_22155,N_22306);
or U23872 (N_23872,N_22649,N_22417);
nand U23873 (N_23873,N_22383,N_22546);
xnor U23874 (N_23874,N_22645,N_22538);
nand U23875 (N_23875,N_22938,N_22117);
xnor U23876 (N_23876,N_22570,N_22134);
xor U23877 (N_23877,N_22798,N_22237);
nand U23878 (N_23878,N_22626,N_22320);
nand U23879 (N_23879,N_22888,N_22889);
nor U23880 (N_23880,N_22117,N_22095);
nand U23881 (N_23881,N_22201,N_22595);
xnor U23882 (N_23882,N_22478,N_22528);
and U23883 (N_23883,N_22979,N_22558);
or U23884 (N_23884,N_22833,N_22639);
or U23885 (N_23885,N_22284,N_22519);
and U23886 (N_23886,N_22660,N_22894);
xor U23887 (N_23887,N_22670,N_22908);
nor U23888 (N_23888,N_22746,N_22199);
xnor U23889 (N_23889,N_22938,N_22373);
and U23890 (N_23890,N_22130,N_22979);
and U23891 (N_23891,N_22942,N_22909);
and U23892 (N_23892,N_22550,N_22380);
nor U23893 (N_23893,N_22048,N_22888);
or U23894 (N_23894,N_22270,N_22914);
nand U23895 (N_23895,N_22562,N_22573);
or U23896 (N_23896,N_22356,N_22467);
nor U23897 (N_23897,N_22148,N_22727);
nand U23898 (N_23898,N_22301,N_22417);
or U23899 (N_23899,N_22127,N_22058);
and U23900 (N_23900,N_22686,N_22945);
xnor U23901 (N_23901,N_22886,N_22109);
or U23902 (N_23902,N_22721,N_22546);
xnor U23903 (N_23903,N_22446,N_22232);
and U23904 (N_23904,N_22546,N_22566);
or U23905 (N_23905,N_22614,N_22827);
and U23906 (N_23906,N_22159,N_22491);
or U23907 (N_23907,N_22329,N_22642);
or U23908 (N_23908,N_22701,N_22842);
or U23909 (N_23909,N_22796,N_22181);
nand U23910 (N_23910,N_22836,N_22956);
nand U23911 (N_23911,N_22697,N_22809);
or U23912 (N_23912,N_22005,N_22654);
xnor U23913 (N_23913,N_22742,N_22659);
xor U23914 (N_23914,N_22891,N_22966);
nand U23915 (N_23915,N_22072,N_22674);
nor U23916 (N_23916,N_22524,N_22645);
xor U23917 (N_23917,N_22590,N_22063);
nor U23918 (N_23918,N_22618,N_22970);
and U23919 (N_23919,N_22398,N_22548);
and U23920 (N_23920,N_22620,N_22892);
nand U23921 (N_23921,N_22661,N_22393);
nand U23922 (N_23922,N_22381,N_22810);
nand U23923 (N_23923,N_22457,N_22179);
or U23924 (N_23924,N_22622,N_22885);
nand U23925 (N_23925,N_22346,N_22013);
nand U23926 (N_23926,N_22106,N_22382);
xor U23927 (N_23927,N_22175,N_22802);
nand U23928 (N_23928,N_22401,N_22720);
nand U23929 (N_23929,N_22094,N_22585);
nor U23930 (N_23930,N_22436,N_22574);
xnor U23931 (N_23931,N_22789,N_22963);
xnor U23932 (N_23932,N_22812,N_22568);
or U23933 (N_23933,N_22384,N_22007);
nand U23934 (N_23934,N_22029,N_22386);
and U23935 (N_23935,N_22694,N_22565);
or U23936 (N_23936,N_22906,N_22730);
nand U23937 (N_23937,N_22547,N_22628);
or U23938 (N_23938,N_22112,N_22561);
nor U23939 (N_23939,N_22975,N_22210);
nand U23940 (N_23940,N_22162,N_22648);
xor U23941 (N_23941,N_22074,N_22763);
and U23942 (N_23942,N_22851,N_22922);
nand U23943 (N_23943,N_22477,N_22444);
or U23944 (N_23944,N_22794,N_22104);
and U23945 (N_23945,N_22574,N_22242);
nand U23946 (N_23946,N_22365,N_22219);
nand U23947 (N_23947,N_22646,N_22290);
nor U23948 (N_23948,N_22879,N_22979);
or U23949 (N_23949,N_22793,N_22949);
xnor U23950 (N_23950,N_22662,N_22659);
nand U23951 (N_23951,N_22388,N_22275);
and U23952 (N_23952,N_22919,N_22962);
or U23953 (N_23953,N_22137,N_22842);
nand U23954 (N_23954,N_22477,N_22503);
or U23955 (N_23955,N_22354,N_22570);
nor U23956 (N_23956,N_22389,N_22756);
and U23957 (N_23957,N_22412,N_22073);
xor U23958 (N_23958,N_22037,N_22862);
xor U23959 (N_23959,N_22374,N_22532);
xnor U23960 (N_23960,N_22395,N_22335);
nor U23961 (N_23961,N_22301,N_22376);
nor U23962 (N_23962,N_22762,N_22339);
nor U23963 (N_23963,N_22685,N_22689);
and U23964 (N_23964,N_22137,N_22634);
nor U23965 (N_23965,N_22461,N_22610);
xor U23966 (N_23966,N_22426,N_22871);
nor U23967 (N_23967,N_22875,N_22390);
and U23968 (N_23968,N_22906,N_22927);
nand U23969 (N_23969,N_22171,N_22482);
or U23970 (N_23970,N_22031,N_22908);
nand U23971 (N_23971,N_22220,N_22864);
nor U23972 (N_23972,N_22553,N_22320);
or U23973 (N_23973,N_22916,N_22441);
nor U23974 (N_23974,N_22952,N_22832);
nor U23975 (N_23975,N_22112,N_22614);
nand U23976 (N_23976,N_22150,N_22064);
or U23977 (N_23977,N_22917,N_22165);
nand U23978 (N_23978,N_22704,N_22492);
and U23979 (N_23979,N_22315,N_22157);
nand U23980 (N_23980,N_22265,N_22393);
and U23981 (N_23981,N_22061,N_22284);
or U23982 (N_23982,N_22107,N_22928);
nor U23983 (N_23983,N_22427,N_22935);
nand U23984 (N_23984,N_22611,N_22676);
and U23985 (N_23985,N_22974,N_22171);
and U23986 (N_23986,N_22933,N_22516);
xnor U23987 (N_23987,N_22379,N_22294);
nor U23988 (N_23988,N_22863,N_22852);
and U23989 (N_23989,N_22609,N_22493);
xor U23990 (N_23990,N_22888,N_22825);
nor U23991 (N_23991,N_22847,N_22305);
or U23992 (N_23992,N_22260,N_22662);
or U23993 (N_23993,N_22476,N_22924);
and U23994 (N_23994,N_22278,N_22715);
nor U23995 (N_23995,N_22269,N_22706);
nor U23996 (N_23996,N_22217,N_22292);
and U23997 (N_23997,N_22248,N_22678);
nand U23998 (N_23998,N_22908,N_22772);
xnor U23999 (N_23999,N_22881,N_22073);
nor U24000 (N_24000,N_23903,N_23487);
or U24001 (N_24001,N_23003,N_23490);
and U24002 (N_24002,N_23025,N_23662);
or U24003 (N_24003,N_23779,N_23952);
nor U24004 (N_24004,N_23657,N_23872);
xor U24005 (N_24005,N_23471,N_23883);
xnor U24006 (N_24006,N_23301,N_23243);
and U24007 (N_24007,N_23240,N_23459);
xnor U24008 (N_24008,N_23644,N_23632);
nand U24009 (N_24009,N_23922,N_23848);
or U24010 (N_24010,N_23699,N_23043);
nor U24011 (N_24011,N_23492,N_23843);
xor U24012 (N_24012,N_23207,N_23065);
nor U24013 (N_24013,N_23723,N_23517);
nor U24014 (N_24014,N_23735,N_23098);
nand U24015 (N_24015,N_23920,N_23849);
or U24016 (N_24016,N_23675,N_23069);
and U24017 (N_24017,N_23093,N_23483);
nor U24018 (N_24018,N_23289,N_23606);
nor U24019 (N_24019,N_23361,N_23695);
nand U24020 (N_24020,N_23727,N_23740);
and U24021 (N_24021,N_23323,N_23251);
xnor U24022 (N_24022,N_23124,N_23566);
nand U24023 (N_24023,N_23269,N_23890);
and U24024 (N_24024,N_23180,N_23198);
or U24025 (N_24025,N_23529,N_23930);
nor U24026 (N_24026,N_23878,N_23295);
nor U24027 (N_24027,N_23297,N_23881);
and U24028 (N_24028,N_23232,N_23418);
and U24029 (N_24029,N_23283,N_23537);
or U24030 (N_24030,N_23976,N_23480);
nor U24031 (N_24031,N_23082,N_23504);
nor U24032 (N_24032,N_23742,N_23173);
or U24033 (N_24033,N_23118,N_23507);
and U24034 (N_24034,N_23114,N_23332);
nor U24035 (N_24035,N_23542,N_23470);
nor U24036 (N_24036,N_23640,N_23137);
and U24037 (N_24037,N_23970,N_23163);
nand U24038 (N_24038,N_23816,N_23979);
and U24039 (N_24039,N_23564,N_23687);
and U24040 (N_24040,N_23485,N_23033);
or U24041 (N_24041,N_23312,N_23782);
and U24042 (N_24042,N_23191,N_23176);
and U24043 (N_24043,N_23619,N_23886);
xnor U24044 (N_24044,N_23255,N_23135);
or U24045 (N_24045,N_23122,N_23860);
and U24046 (N_24046,N_23372,N_23447);
or U24047 (N_24047,N_23998,N_23253);
nor U24048 (N_24048,N_23407,N_23293);
and U24049 (N_24049,N_23831,N_23128);
nand U24050 (N_24050,N_23009,N_23916);
and U24051 (N_24051,N_23776,N_23246);
nand U24052 (N_24052,N_23428,N_23808);
or U24053 (N_24053,N_23494,N_23693);
and U24054 (N_24054,N_23557,N_23469);
nor U24055 (N_24055,N_23919,N_23968);
and U24056 (N_24056,N_23969,N_23142);
nor U24057 (N_24057,N_23584,N_23261);
nor U24058 (N_24058,N_23309,N_23245);
xor U24059 (N_24059,N_23604,N_23885);
or U24060 (N_24060,N_23086,N_23263);
nand U24061 (N_24061,N_23343,N_23132);
or U24062 (N_24062,N_23649,N_23368);
and U24063 (N_24063,N_23822,N_23214);
nand U24064 (N_24064,N_23873,N_23024);
or U24065 (N_24065,N_23169,N_23404);
or U24066 (N_24066,N_23146,N_23461);
nor U24067 (N_24067,N_23053,N_23268);
nand U24068 (N_24068,N_23195,N_23586);
nor U24069 (N_24069,N_23398,N_23907);
xor U24070 (N_24070,N_23204,N_23123);
and U24071 (N_24071,N_23598,N_23955);
nand U24072 (N_24072,N_23452,N_23905);
or U24073 (N_24073,N_23220,N_23829);
or U24074 (N_24074,N_23642,N_23565);
nand U24075 (N_24075,N_23219,N_23030);
or U24076 (N_24076,N_23582,N_23613);
nor U24077 (N_24077,N_23560,N_23753);
nor U24078 (N_24078,N_23274,N_23850);
xor U24079 (N_24079,N_23547,N_23441);
nand U24080 (N_24080,N_23096,N_23999);
nand U24081 (N_24081,N_23451,N_23838);
nand U24082 (N_24082,N_23310,N_23091);
xnor U24083 (N_24083,N_23868,N_23071);
and U24084 (N_24084,N_23771,N_23789);
nor U24085 (N_24085,N_23997,N_23089);
xor U24086 (N_24086,N_23062,N_23541);
or U24087 (N_24087,N_23972,N_23202);
xor U24088 (N_24088,N_23174,N_23320);
xnor U24089 (N_24089,N_23798,N_23936);
nand U24090 (N_24090,N_23403,N_23530);
and U24091 (N_24091,N_23935,N_23410);
nand U24092 (N_24092,N_23574,N_23884);
nand U24093 (N_24093,N_23104,N_23570);
or U24094 (N_24094,N_23773,N_23830);
xor U24095 (N_24095,N_23326,N_23190);
nor U24096 (N_24096,N_23419,N_23421);
xnor U24097 (N_24097,N_23651,N_23673);
or U24098 (N_24098,N_23627,N_23569);
xor U24099 (N_24099,N_23327,N_23159);
or U24100 (N_24100,N_23317,N_23197);
and U24101 (N_24101,N_23505,N_23050);
and U24102 (N_24102,N_23577,N_23305);
or U24103 (N_24103,N_23778,N_23988);
xnor U24104 (N_24104,N_23439,N_23097);
nor U24105 (N_24105,N_23286,N_23933);
and U24106 (N_24106,N_23856,N_23691);
nand U24107 (N_24107,N_23654,N_23580);
and U24108 (N_24108,N_23506,N_23993);
xor U24109 (N_24109,N_23084,N_23514);
nand U24110 (N_24110,N_23801,N_23397);
xor U24111 (N_24111,N_23608,N_23425);
and U24112 (N_24112,N_23593,N_23623);
or U24113 (N_24113,N_23626,N_23717);
nor U24114 (N_24114,N_23085,N_23351);
or U24115 (N_24115,N_23304,N_23511);
or U24116 (N_24116,N_23661,N_23802);
nand U24117 (N_24117,N_23591,N_23746);
nor U24118 (N_24118,N_23681,N_23959);
and U24119 (N_24119,N_23170,N_23156);
and U24120 (N_24120,N_23700,N_23119);
nand U24121 (N_24121,N_23684,N_23667);
and U24122 (N_24122,N_23756,N_23852);
or U24123 (N_24123,N_23821,N_23815);
nor U24124 (N_24124,N_23339,N_23012);
nor U24125 (N_24125,N_23215,N_23844);
and U24126 (N_24126,N_23949,N_23045);
xnor U24127 (N_24127,N_23680,N_23005);
and U24128 (N_24128,N_23719,N_23656);
and U24129 (N_24129,N_23736,N_23165);
and U24130 (N_24130,N_23520,N_23303);
nor U24131 (N_24131,N_23110,N_23076);
xnor U24132 (N_24132,N_23787,N_23278);
nor U24133 (N_24133,N_23276,N_23185);
or U24134 (N_24134,N_23247,N_23502);
nand U24135 (N_24135,N_23677,N_23704);
and U24136 (N_24136,N_23252,N_23855);
nand U24137 (N_24137,N_23229,N_23763);
xnor U24138 (N_24138,N_23874,N_23200);
nand U24139 (N_24139,N_23558,N_23774);
and U24140 (N_24140,N_23664,N_23395);
nor U24141 (N_24141,N_23356,N_23328);
or U24142 (N_24142,N_23536,N_23857);
xor U24143 (N_24143,N_23929,N_23411);
nor U24144 (N_24144,N_23038,N_23401);
nor U24145 (N_24145,N_23047,N_23585);
and U24146 (N_24146,N_23650,N_23548);
or U24147 (N_24147,N_23747,N_23039);
or U24148 (N_24148,N_23319,N_23168);
nand U24149 (N_24149,N_23184,N_23277);
nand U24150 (N_24150,N_23781,N_23175);
nand U24151 (N_24151,N_23383,N_23694);
nor U24152 (N_24152,N_23543,N_23942);
and U24153 (N_24153,N_23898,N_23400);
and U24154 (N_24154,N_23550,N_23408);
and U24155 (N_24155,N_23688,N_23218);
xor U24156 (N_24156,N_23051,N_23369);
or U24157 (N_24157,N_23436,N_23912);
xnor U24158 (N_24158,N_23768,N_23015);
nand U24159 (N_24159,N_23551,N_23824);
nor U24160 (N_24160,N_23417,N_23029);
xnor U24161 (N_24161,N_23671,N_23177);
nand U24162 (N_24162,N_23162,N_23630);
nand U24163 (N_24163,N_23239,N_23980);
nor U24164 (N_24164,N_23178,N_23875);
xnor U24165 (N_24165,N_23475,N_23499);
or U24166 (N_24166,N_23112,N_23237);
and U24167 (N_24167,N_23224,N_23008);
nand U24168 (N_24168,N_23948,N_23234);
xnor U24169 (N_24169,N_23192,N_23772);
nand U24170 (N_24170,N_23796,N_23462);
and U24171 (N_24171,N_23722,N_23702);
nor U24172 (N_24172,N_23805,N_23841);
xnor U24173 (N_24173,N_23108,N_23526);
and U24174 (N_24174,N_23040,N_23612);
nor U24175 (N_24175,N_23944,N_23423);
xnor U24176 (N_24176,N_23555,N_23420);
and U24177 (N_24177,N_23209,N_23187);
and U24178 (N_24178,N_23669,N_23960);
and U24179 (N_24179,N_23910,N_23906);
nand U24180 (N_24180,N_23064,N_23016);
or U24181 (N_24181,N_23095,N_23587);
nand U24182 (N_24182,N_23019,N_23412);
nor U24183 (N_24183,N_23895,N_23458);
xnor U24184 (N_24184,N_23834,N_23380);
xor U24185 (N_24185,N_23892,N_23641);
xnor U24186 (N_24186,N_23576,N_23761);
or U24187 (N_24187,N_23974,N_23610);
or U24188 (N_24188,N_23055,N_23329);
nand U24189 (N_24189,N_23210,N_23167);
nor U24190 (N_24190,N_23666,N_23186);
or U24191 (N_24191,N_23058,N_23140);
nor U24192 (N_24192,N_23357,N_23041);
nand U24193 (N_24193,N_23867,N_23100);
or U24194 (N_24194,N_23981,N_23638);
and U24195 (N_24195,N_23963,N_23048);
nor U24196 (N_24196,N_23429,N_23007);
or U24197 (N_24197,N_23049,N_23896);
nand U24198 (N_24198,N_23424,N_23990);
and U24199 (N_24199,N_23248,N_23618);
nor U24200 (N_24200,N_23535,N_23553);
xor U24201 (N_24201,N_23864,N_23059);
xnor U24202 (N_24202,N_23628,N_23663);
nor U24203 (N_24203,N_23827,N_23670);
and U24204 (N_24204,N_23172,N_23958);
nand U24205 (N_24205,N_23105,N_23915);
xor U24206 (N_24206,N_23217,N_23296);
or U24207 (N_24207,N_23353,N_23189);
nor U24208 (N_24208,N_23338,N_23571);
nor U24209 (N_24209,N_23692,N_23938);
nor U24210 (N_24210,N_23943,N_23706);
nand U24211 (N_24211,N_23000,N_23316);
or U24212 (N_24212,N_23645,N_23399);
nand U24213 (N_24213,N_23525,N_23031);
nor U24214 (N_24214,N_23596,N_23106);
and U24215 (N_24215,N_23486,N_23705);
xnor U24216 (N_24216,N_23738,N_23812);
or U24217 (N_24217,N_23624,N_23523);
xnor U24218 (N_24218,N_23531,N_23054);
nand U24219 (N_24219,N_23897,N_23762);
or U24220 (N_24220,N_23063,N_23734);
nor U24221 (N_24221,N_23396,N_23080);
xnor U24222 (N_24222,N_23804,N_23083);
or U24223 (N_24223,N_23710,N_23902);
xnor U24224 (N_24224,N_23921,N_23876);
or U24225 (N_24225,N_23951,N_23166);
nand U24226 (N_24226,N_23730,N_23386);
and U24227 (N_24227,N_23973,N_23911);
nand U24228 (N_24228,N_23044,N_23371);
xnor U24229 (N_24229,N_23674,N_23602);
or U24230 (N_24230,N_23346,N_23340);
xor U24231 (N_24231,N_23904,N_23465);
nand U24232 (N_24232,N_23780,N_23367);
or U24233 (N_24233,N_23479,N_23767);
xnor U24234 (N_24234,N_23021,N_23010);
xnor U24235 (N_24235,N_23837,N_23101);
or U24236 (N_24236,N_23299,N_23803);
xnor U24237 (N_24237,N_23442,N_23621);
nand U24238 (N_24238,N_23559,N_23111);
xor U24239 (N_24239,N_23561,N_23046);
or U24240 (N_24240,N_23818,N_23467);
or U24241 (N_24241,N_23254,N_23307);
nor U24242 (N_24242,N_23264,N_23540);
and U24243 (N_24243,N_23201,N_23018);
or U24244 (N_24244,N_23785,N_23438);
and U24245 (N_24245,N_23836,N_23790);
or U24246 (N_24246,N_23057,N_23179);
or U24247 (N_24247,N_23134,N_23924);
and U24248 (N_24248,N_23810,N_23847);
nor U24249 (N_24249,N_23472,N_23481);
and U24250 (N_24250,N_23279,N_23151);
and U24251 (N_24251,N_23394,N_23409);
and U24252 (N_24252,N_23879,N_23311);
nand U24253 (N_24253,N_23594,N_23145);
or U24254 (N_24254,N_23182,N_23643);
xnor U24255 (N_24255,N_23127,N_23701);
nand U24256 (N_24256,N_23568,N_23599);
and U24257 (N_24257,N_23149,N_23588);
and U24258 (N_24258,N_23950,N_23249);
and U24259 (N_24259,N_23658,N_23287);
nor U24260 (N_24260,N_23171,N_23877);
nor U24261 (N_24261,N_23258,N_23391);
and U24262 (N_24262,N_23652,N_23527);
and U24263 (N_24263,N_23769,N_23784);
or U24264 (N_24264,N_23230,N_23282);
or U24265 (N_24265,N_23298,N_23109);
and U24266 (N_24266,N_23927,N_23291);
nand U24267 (N_24267,N_23116,N_23744);
and U24268 (N_24268,N_23378,N_23545);
xnor U24269 (N_24269,N_23679,N_23552);
nand U24270 (N_24270,N_23639,N_23528);
and U24271 (N_24271,N_23379,N_23724);
xnor U24272 (N_24272,N_23267,N_23607);
nor U24273 (N_24273,N_23799,N_23842);
or U24274 (N_24274,N_23113,N_23631);
or U24275 (N_24275,N_23617,N_23614);
or U24276 (N_24276,N_23795,N_23503);
or U24277 (N_24277,N_23260,N_23355);
nor U24278 (N_24278,N_23444,N_23636);
nand U24279 (N_24279,N_23665,N_23611);
xor U24280 (N_24280,N_23102,N_23103);
or U24281 (N_24281,N_23579,N_23759);
xor U24282 (N_24282,N_23042,N_23389);
and U24283 (N_24283,N_23382,N_23928);
and U24284 (N_24284,N_23971,N_23074);
nor U24285 (N_24285,N_23061,N_23004);
and U24286 (N_24286,N_23713,N_23225);
xor U24287 (N_24287,N_23073,N_23148);
xor U24288 (N_24288,N_23139,N_23956);
and U24289 (N_24289,N_23066,N_23908);
nand U24290 (N_24290,N_23257,N_23750);
and U24291 (N_24291,N_23512,N_23463);
nand U24292 (N_24292,N_23228,N_23342);
and U24293 (N_24293,N_23280,N_23017);
or U24294 (N_24294,N_23572,N_23385);
xor U24295 (N_24295,N_23181,N_23306);
and U24296 (N_24296,N_23402,N_23205);
nand U24297 (N_24297,N_23414,N_23115);
nor U24298 (N_24298,N_23256,N_23720);
or U24299 (N_24299,N_23581,N_23333);
nor U24300 (N_24300,N_23242,N_23600);
xnor U24301 (N_24301,N_23646,N_23538);
or U24302 (N_24302,N_23213,N_23851);
nand U24303 (N_24303,N_23496,N_23698);
or U24304 (N_24304,N_23390,N_23788);
and U24305 (N_24305,N_23211,N_23913);
nor U24306 (N_24306,N_23996,N_23318);
and U24307 (N_24307,N_23947,N_23144);
or U24308 (N_24308,N_23862,N_23154);
or U24309 (N_24309,N_23986,N_23544);
or U24310 (N_24310,N_23077,N_23393);
nor U24311 (N_24311,N_23573,N_23133);
nand U24312 (N_24312,N_23743,N_23359);
xnor U24313 (N_24313,N_23622,N_23322);
nor U24314 (N_24314,N_23806,N_23381);
and U24315 (N_24315,N_23739,N_23894);
or U24316 (N_24316,N_23648,N_23482);
xor U24317 (N_24317,N_23770,N_23629);
xor U24318 (N_24318,N_23079,N_23075);
nand U24319 (N_24319,N_23023,N_23453);
nor U24320 (N_24320,N_23160,N_23995);
and U24321 (N_24321,N_23521,N_23203);
nor U24322 (N_24322,N_23989,N_23957);
or U24323 (N_24323,N_23099,N_23491);
xnor U24324 (N_24324,N_23011,N_23931);
and U24325 (N_24325,N_23766,N_23783);
xor U24326 (N_24326,N_23493,N_23013);
nand U24327 (N_24327,N_23865,N_23984);
xor U24328 (N_24328,N_23757,N_23647);
nor U24329 (N_24329,N_23388,N_23620);
nor U24330 (N_24330,N_23854,N_23953);
nor U24331 (N_24331,N_23497,N_23792);
nand U24332 (N_24332,N_23152,N_23001);
nor U24333 (N_24333,N_23216,N_23072);
xor U24334 (N_24334,N_23899,N_23501);
nand U24335 (N_24335,N_23370,N_23052);
or U24336 (N_24336,N_23888,N_23440);
nand U24337 (N_24337,N_23697,N_23590);
nor U24338 (N_24338,N_23364,N_23431);
xnor U24339 (N_24339,N_23188,N_23509);
nand U24340 (N_24340,N_23288,N_23349);
or U24341 (N_24341,N_23285,N_23302);
nor U24342 (N_24342,N_23334,N_23078);
xor U24343 (N_24343,N_23835,N_23433);
and U24344 (N_24344,N_23158,N_23194);
nor U24345 (N_24345,N_23961,N_23982);
nand U24346 (N_24346,N_23721,N_23157);
nor U24347 (N_24347,N_23718,N_23519);
or U24348 (N_24348,N_23056,N_23889);
and U24349 (N_24349,N_23498,N_23833);
and U24350 (N_24350,N_23513,N_23153);
and U24351 (N_24351,N_23235,N_23826);
xnor U24352 (N_24352,N_23765,N_23726);
xnor U24353 (N_24353,N_23917,N_23703);
xnor U24354 (N_24354,N_23406,N_23978);
nor U24355 (N_24355,N_23366,N_23869);
nor U24356 (N_24356,N_23358,N_23094);
and U24357 (N_24357,N_23820,N_23655);
or U24358 (N_24358,N_23478,N_23616);
nor U24359 (N_24359,N_23236,N_23081);
and U24360 (N_24360,N_23934,N_23231);
nand U24361 (N_24361,N_23026,N_23244);
and U24362 (N_24362,N_23846,N_23716);
and U24363 (N_24363,N_23136,N_23087);
nand U24364 (N_24364,N_23227,N_23374);
nor U24365 (N_24365,N_23965,N_23634);
xnor U24366 (N_24366,N_23589,N_23281);
or U24367 (N_24367,N_23208,N_23221);
xnor U24368 (N_24368,N_23678,N_23430);
nand U24369 (N_24369,N_23672,N_23653);
and U24370 (N_24370,N_23567,N_23575);
nor U24371 (N_24371,N_23344,N_23308);
xnor U24372 (N_24372,N_23696,N_23454);
nand U24373 (N_24373,N_23271,N_23335);
xnor U24374 (N_24374,N_23384,N_23712);
nor U24375 (N_24375,N_23828,N_23807);
nor U24376 (N_24376,N_23377,N_23484);
nor U24377 (N_24377,N_23445,N_23866);
xnor U24378 (N_24378,N_23635,N_23450);
nor U24379 (N_24379,N_23615,N_23825);
xor U24380 (N_24380,N_23745,N_23354);
nand U24381 (N_24381,N_23284,N_23549);
nand U24382 (N_24382,N_23983,N_23732);
nor U24383 (N_24383,N_23609,N_23443);
and U24384 (N_24384,N_23130,N_23273);
or U24385 (N_24385,N_23977,N_23068);
or U24386 (N_24386,N_23918,N_23832);
and U24387 (N_24387,N_23362,N_23376);
and U24388 (N_24388,N_23754,N_23595);
xor U24389 (N_24389,N_23633,N_23238);
xnor U24390 (N_24390,N_23707,N_23416);
or U24391 (N_24391,N_23006,N_23887);
or U24392 (N_24392,N_23129,N_23562);
nand U24393 (N_24393,N_23262,N_23809);
nor U24394 (N_24394,N_23964,N_23427);
nand U24395 (N_24395,N_23660,N_23233);
and U24396 (N_24396,N_23413,N_23121);
or U24397 (N_24397,N_23597,N_23314);
xor U24398 (N_24398,N_23985,N_23516);
nand U24399 (N_24399,N_23090,N_23415);
nor U24400 (N_24400,N_23926,N_23117);
and U24401 (N_24401,N_23345,N_23914);
and U24402 (N_24402,N_23088,N_23728);
xor U24403 (N_24403,N_23532,N_23435);
nand U24404 (N_24404,N_23468,N_23449);
nand U24405 (N_24405,N_23975,N_23556);
and U24406 (N_24406,N_23932,N_23554);
and U24407 (N_24407,N_23592,N_23966);
and U24408 (N_24408,N_23477,N_23464);
and U24409 (N_24409,N_23941,N_23473);
nand U24410 (N_24410,N_23455,N_23987);
or U24411 (N_24411,N_23199,N_23777);
nor U24412 (N_24412,N_23027,N_23294);
xor U24413 (N_24413,N_23020,N_23028);
xnor U24414 (N_24414,N_23786,N_23092);
nor U24415 (N_24415,N_23515,N_23032);
and U24416 (N_24416,N_23925,N_23222);
xnor U24417 (N_24417,N_23155,N_23432);
or U24418 (N_24418,N_23495,N_23070);
nand U24419 (N_24419,N_23290,N_23206);
or U24420 (N_24420,N_23563,N_23714);
xor U24421 (N_24421,N_23275,N_23946);
xnor U24422 (N_24422,N_23360,N_23711);
xnor U24423 (N_24423,N_23534,N_23321);
or U24424 (N_24424,N_23797,N_23466);
or U24425 (N_24425,N_23161,N_23882);
nand U24426 (N_24426,N_23325,N_23668);
and U24427 (N_24427,N_23347,N_23752);
and U24428 (N_24428,N_23845,N_23751);
nor U24429 (N_24429,N_23539,N_23315);
and U24430 (N_24430,N_23813,N_23682);
and U24431 (N_24431,N_23143,N_23270);
xor U24432 (N_24432,N_23939,N_23373);
and U24433 (N_24433,N_23689,N_23625);
and U24434 (N_24434,N_23223,N_23300);
nand U24435 (N_24435,N_23880,N_23764);
xor U24436 (N_24436,N_23794,N_23060);
or U24437 (N_24437,N_23035,N_23755);
and U24438 (N_24438,N_23002,N_23446);
and U24439 (N_24439,N_23266,N_23337);
xnor U24440 (N_24440,N_23448,N_23690);
xnor U24441 (N_24441,N_23226,N_23954);
nand U24442 (N_24442,N_23476,N_23488);
xor U24443 (N_24443,N_23405,N_23375);
nand U24444 (N_24444,N_23731,N_23861);
xor U24445 (N_24445,N_23272,N_23265);
nand U24446 (N_24446,N_23605,N_23729);
nand U24447 (N_24447,N_23758,N_23034);
nor U24448 (N_24448,N_23749,N_23363);
or U24449 (N_24449,N_23352,N_23870);
xnor U24450 (N_24450,N_23292,N_23715);
nand U24451 (N_24451,N_23489,N_23241);
and U24452 (N_24452,N_23811,N_23387);
nand U24453 (N_24453,N_23067,N_23331);
nand U24454 (N_24454,N_23500,N_23365);
and U24455 (N_24455,N_23150,N_23457);
nand U24456 (N_24456,N_23725,N_23819);
or U24457 (N_24457,N_23183,N_23709);
nand U24458 (N_24458,N_23791,N_23456);
and U24459 (N_24459,N_23893,N_23259);
nor U24460 (N_24460,N_23324,N_23422);
or U24461 (N_24461,N_23676,N_23683);
xor U24462 (N_24462,N_23107,N_23637);
xor U24463 (N_24463,N_23037,N_23871);
xnor U24464 (N_24464,N_23760,N_23900);
nor U24465 (N_24465,N_23126,N_23348);
nand U24466 (N_24466,N_23250,N_23800);
nand U24467 (N_24467,N_23336,N_23022);
or U24468 (N_24468,N_23937,N_23546);
and U24469 (N_24469,N_23603,N_23601);
nor U24470 (N_24470,N_23992,N_23793);
or U24471 (N_24471,N_23522,N_23994);
or U24472 (N_24472,N_23533,N_23120);
nand U24473 (N_24473,N_23141,N_23125);
or U24474 (N_24474,N_23147,N_23708);
xor U24475 (N_24475,N_23460,N_23859);
nor U24476 (N_24476,N_23131,N_23840);
xnor U24477 (N_24477,N_23583,N_23518);
xor U24478 (N_24478,N_23014,N_23962);
and U24479 (N_24479,N_23524,N_23510);
nand U24480 (N_24480,N_23164,N_23036);
xnor U24481 (N_24481,N_23330,N_23686);
nor U24482 (N_24482,N_23350,N_23858);
nor U24483 (N_24483,N_23923,N_23196);
nor U24484 (N_24484,N_23748,N_23909);
nor U24485 (N_24485,N_23659,N_23891);
nor U24486 (N_24486,N_23901,N_23508);
and U24487 (N_24487,N_23741,N_23945);
xor U24488 (N_24488,N_23434,N_23823);
xor U24489 (N_24489,N_23474,N_23193);
xnor U24490 (N_24490,N_23853,N_23817);
nand U24491 (N_24491,N_23863,N_23685);
nor U24492 (N_24492,N_23341,N_23991);
or U24493 (N_24493,N_23733,N_23737);
or U24494 (N_24494,N_23313,N_23426);
or U24495 (N_24495,N_23212,N_23775);
xnor U24496 (N_24496,N_23578,N_23814);
xor U24497 (N_24497,N_23138,N_23940);
or U24498 (N_24498,N_23967,N_23839);
or U24499 (N_24499,N_23437,N_23392);
nor U24500 (N_24500,N_23279,N_23828);
nand U24501 (N_24501,N_23690,N_23467);
or U24502 (N_24502,N_23309,N_23259);
or U24503 (N_24503,N_23331,N_23087);
nor U24504 (N_24504,N_23669,N_23978);
nand U24505 (N_24505,N_23471,N_23151);
or U24506 (N_24506,N_23727,N_23307);
xor U24507 (N_24507,N_23169,N_23933);
nor U24508 (N_24508,N_23393,N_23634);
nor U24509 (N_24509,N_23530,N_23940);
nor U24510 (N_24510,N_23082,N_23434);
nor U24511 (N_24511,N_23448,N_23202);
or U24512 (N_24512,N_23403,N_23803);
and U24513 (N_24513,N_23131,N_23328);
and U24514 (N_24514,N_23920,N_23818);
xnor U24515 (N_24515,N_23850,N_23490);
nand U24516 (N_24516,N_23866,N_23459);
nand U24517 (N_24517,N_23768,N_23946);
nor U24518 (N_24518,N_23296,N_23643);
or U24519 (N_24519,N_23846,N_23802);
or U24520 (N_24520,N_23176,N_23991);
xor U24521 (N_24521,N_23251,N_23257);
nand U24522 (N_24522,N_23226,N_23307);
nand U24523 (N_24523,N_23945,N_23339);
and U24524 (N_24524,N_23376,N_23745);
nand U24525 (N_24525,N_23559,N_23863);
xor U24526 (N_24526,N_23666,N_23668);
xor U24527 (N_24527,N_23077,N_23928);
xor U24528 (N_24528,N_23286,N_23861);
or U24529 (N_24529,N_23959,N_23083);
nor U24530 (N_24530,N_23342,N_23082);
and U24531 (N_24531,N_23442,N_23938);
xor U24532 (N_24532,N_23344,N_23298);
and U24533 (N_24533,N_23424,N_23429);
nand U24534 (N_24534,N_23574,N_23398);
nand U24535 (N_24535,N_23460,N_23672);
nor U24536 (N_24536,N_23556,N_23088);
and U24537 (N_24537,N_23178,N_23519);
nand U24538 (N_24538,N_23146,N_23468);
xnor U24539 (N_24539,N_23391,N_23183);
or U24540 (N_24540,N_23707,N_23781);
nand U24541 (N_24541,N_23102,N_23345);
xor U24542 (N_24542,N_23105,N_23340);
and U24543 (N_24543,N_23208,N_23268);
and U24544 (N_24544,N_23245,N_23128);
and U24545 (N_24545,N_23825,N_23258);
or U24546 (N_24546,N_23694,N_23022);
or U24547 (N_24547,N_23277,N_23789);
and U24548 (N_24548,N_23289,N_23165);
nor U24549 (N_24549,N_23317,N_23085);
and U24550 (N_24550,N_23654,N_23809);
xor U24551 (N_24551,N_23081,N_23988);
and U24552 (N_24552,N_23532,N_23157);
nand U24553 (N_24553,N_23017,N_23845);
nor U24554 (N_24554,N_23691,N_23378);
and U24555 (N_24555,N_23265,N_23991);
nand U24556 (N_24556,N_23394,N_23763);
nor U24557 (N_24557,N_23833,N_23468);
xnor U24558 (N_24558,N_23325,N_23496);
nand U24559 (N_24559,N_23727,N_23491);
or U24560 (N_24560,N_23970,N_23765);
nand U24561 (N_24561,N_23539,N_23001);
xor U24562 (N_24562,N_23371,N_23832);
or U24563 (N_24563,N_23110,N_23125);
and U24564 (N_24564,N_23139,N_23766);
nand U24565 (N_24565,N_23168,N_23948);
xor U24566 (N_24566,N_23680,N_23762);
and U24567 (N_24567,N_23854,N_23976);
and U24568 (N_24568,N_23231,N_23342);
xor U24569 (N_24569,N_23091,N_23506);
and U24570 (N_24570,N_23051,N_23194);
xor U24571 (N_24571,N_23987,N_23612);
nand U24572 (N_24572,N_23422,N_23773);
and U24573 (N_24573,N_23973,N_23979);
xor U24574 (N_24574,N_23809,N_23102);
nand U24575 (N_24575,N_23444,N_23735);
and U24576 (N_24576,N_23938,N_23276);
nor U24577 (N_24577,N_23985,N_23538);
xor U24578 (N_24578,N_23472,N_23080);
and U24579 (N_24579,N_23119,N_23298);
xor U24580 (N_24580,N_23176,N_23444);
nor U24581 (N_24581,N_23084,N_23123);
nor U24582 (N_24582,N_23246,N_23781);
or U24583 (N_24583,N_23220,N_23365);
or U24584 (N_24584,N_23019,N_23719);
xor U24585 (N_24585,N_23082,N_23511);
nor U24586 (N_24586,N_23776,N_23675);
xnor U24587 (N_24587,N_23631,N_23542);
nand U24588 (N_24588,N_23840,N_23782);
xor U24589 (N_24589,N_23279,N_23303);
and U24590 (N_24590,N_23725,N_23926);
or U24591 (N_24591,N_23995,N_23377);
xor U24592 (N_24592,N_23471,N_23253);
xor U24593 (N_24593,N_23448,N_23365);
xor U24594 (N_24594,N_23255,N_23464);
and U24595 (N_24595,N_23034,N_23339);
nand U24596 (N_24596,N_23084,N_23907);
or U24597 (N_24597,N_23448,N_23226);
nor U24598 (N_24598,N_23840,N_23978);
or U24599 (N_24599,N_23807,N_23654);
xor U24600 (N_24600,N_23466,N_23736);
or U24601 (N_24601,N_23805,N_23818);
xor U24602 (N_24602,N_23338,N_23907);
or U24603 (N_24603,N_23912,N_23753);
xor U24604 (N_24604,N_23735,N_23677);
xor U24605 (N_24605,N_23402,N_23947);
and U24606 (N_24606,N_23120,N_23843);
or U24607 (N_24607,N_23253,N_23749);
xnor U24608 (N_24608,N_23095,N_23072);
nor U24609 (N_24609,N_23133,N_23148);
xor U24610 (N_24610,N_23372,N_23608);
xnor U24611 (N_24611,N_23558,N_23865);
nand U24612 (N_24612,N_23316,N_23469);
or U24613 (N_24613,N_23656,N_23037);
or U24614 (N_24614,N_23693,N_23576);
nor U24615 (N_24615,N_23205,N_23707);
xor U24616 (N_24616,N_23385,N_23217);
nor U24617 (N_24617,N_23909,N_23742);
xor U24618 (N_24618,N_23653,N_23202);
nor U24619 (N_24619,N_23000,N_23835);
xor U24620 (N_24620,N_23743,N_23954);
or U24621 (N_24621,N_23728,N_23592);
xnor U24622 (N_24622,N_23336,N_23471);
xnor U24623 (N_24623,N_23977,N_23300);
and U24624 (N_24624,N_23896,N_23847);
nand U24625 (N_24625,N_23992,N_23306);
or U24626 (N_24626,N_23679,N_23967);
xnor U24627 (N_24627,N_23471,N_23165);
or U24628 (N_24628,N_23956,N_23165);
or U24629 (N_24629,N_23257,N_23290);
xor U24630 (N_24630,N_23315,N_23028);
or U24631 (N_24631,N_23477,N_23642);
xor U24632 (N_24632,N_23874,N_23897);
nor U24633 (N_24633,N_23671,N_23560);
or U24634 (N_24634,N_23856,N_23728);
and U24635 (N_24635,N_23733,N_23155);
nand U24636 (N_24636,N_23779,N_23817);
nand U24637 (N_24637,N_23650,N_23796);
xnor U24638 (N_24638,N_23950,N_23000);
nor U24639 (N_24639,N_23206,N_23962);
and U24640 (N_24640,N_23159,N_23164);
xnor U24641 (N_24641,N_23647,N_23946);
nor U24642 (N_24642,N_23208,N_23811);
or U24643 (N_24643,N_23718,N_23556);
nand U24644 (N_24644,N_23638,N_23825);
nor U24645 (N_24645,N_23845,N_23387);
xnor U24646 (N_24646,N_23074,N_23804);
xnor U24647 (N_24647,N_23824,N_23686);
nand U24648 (N_24648,N_23898,N_23228);
xnor U24649 (N_24649,N_23524,N_23144);
nand U24650 (N_24650,N_23387,N_23030);
and U24651 (N_24651,N_23882,N_23026);
or U24652 (N_24652,N_23786,N_23467);
xnor U24653 (N_24653,N_23698,N_23033);
nor U24654 (N_24654,N_23999,N_23801);
nor U24655 (N_24655,N_23343,N_23341);
and U24656 (N_24656,N_23660,N_23219);
or U24657 (N_24657,N_23839,N_23233);
or U24658 (N_24658,N_23952,N_23408);
and U24659 (N_24659,N_23653,N_23976);
and U24660 (N_24660,N_23806,N_23533);
nand U24661 (N_24661,N_23242,N_23711);
nand U24662 (N_24662,N_23014,N_23038);
nand U24663 (N_24663,N_23956,N_23481);
xnor U24664 (N_24664,N_23575,N_23411);
or U24665 (N_24665,N_23698,N_23609);
nor U24666 (N_24666,N_23673,N_23772);
nand U24667 (N_24667,N_23620,N_23370);
xor U24668 (N_24668,N_23615,N_23486);
xor U24669 (N_24669,N_23273,N_23150);
nand U24670 (N_24670,N_23858,N_23881);
or U24671 (N_24671,N_23648,N_23938);
or U24672 (N_24672,N_23482,N_23788);
xnor U24673 (N_24673,N_23318,N_23293);
nor U24674 (N_24674,N_23885,N_23969);
and U24675 (N_24675,N_23632,N_23098);
nand U24676 (N_24676,N_23978,N_23098);
and U24677 (N_24677,N_23446,N_23284);
and U24678 (N_24678,N_23531,N_23873);
nor U24679 (N_24679,N_23738,N_23971);
and U24680 (N_24680,N_23146,N_23694);
nor U24681 (N_24681,N_23581,N_23322);
xnor U24682 (N_24682,N_23832,N_23559);
nor U24683 (N_24683,N_23170,N_23232);
nor U24684 (N_24684,N_23735,N_23401);
nand U24685 (N_24685,N_23925,N_23879);
and U24686 (N_24686,N_23569,N_23380);
nand U24687 (N_24687,N_23351,N_23837);
nand U24688 (N_24688,N_23199,N_23170);
xor U24689 (N_24689,N_23962,N_23698);
or U24690 (N_24690,N_23142,N_23396);
nand U24691 (N_24691,N_23659,N_23725);
xor U24692 (N_24692,N_23190,N_23218);
nor U24693 (N_24693,N_23496,N_23324);
nor U24694 (N_24694,N_23617,N_23914);
or U24695 (N_24695,N_23583,N_23828);
or U24696 (N_24696,N_23674,N_23795);
or U24697 (N_24697,N_23272,N_23541);
or U24698 (N_24698,N_23786,N_23957);
nor U24699 (N_24699,N_23652,N_23547);
nor U24700 (N_24700,N_23556,N_23483);
xor U24701 (N_24701,N_23750,N_23624);
nor U24702 (N_24702,N_23781,N_23334);
or U24703 (N_24703,N_23235,N_23593);
nor U24704 (N_24704,N_23397,N_23721);
xnor U24705 (N_24705,N_23153,N_23933);
and U24706 (N_24706,N_23104,N_23279);
nand U24707 (N_24707,N_23561,N_23197);
xor U24708 (N_24708,N_23826,N_23251);
and U24709 (N_24709,N_23612,N_23230);
nand U24710 (N_24710,N_23620,N_23745);
or U24711 (N_24711,N_23001,N_23424);
nor U24712 (N_24712,N_23691,N_23624);
nand U24713 (N_24713,N_23111,N_23129);
nor U24714 (N_24714,N_23609,N_23702);
or U24715 (N_24715,N_23967,N_23881);
and U24716 (N_24716,N_23070,N_23443);
or U24717 (N_24717,N_23838,N_23094);
nor U24718 (N_24718,N_23440,N_23076);
or U24719 (N_24719,N_23735,N_23038);
nor U24720 (N_24720,N_23660,N_23515);
or U24721 (N_24721,N_23917,N_23248);
nand U24722 (N_24722,N_23712,N_23813);
xnor U24723 (N_24723,N_23597,N_23940);
nor U24724 (N_24724,N_23049,N_23997);
xnor U24725 (N_24725,N_23466,N_23493);
nor U24726 (N_24726,N_23896,N_23300);
nor U24727 (N_24727,N_23035,N_23968);
nand U24728 (N_24728,N_23928,N_23087);
nor U24729 (N_24729,N_23698,N_23632);
or U24730 (N_24730,N_23990,N_23773);
xor U24731 (N_24731,N_23575,N_23998);
nand U24732 (N_24732,N_23662,N_23934);
or U24733 (N_24733,N_23306,N_23964);
or U24734 (N_24734,N_23283,N_23010);
or U24735 (N_24735,N_23417,N_23892);
and U24736 (N_24736,N_23843,N_23611);
nor U24737 (N_24737,N_23182,N_23325);
xor U24738 (N_24738,N_23312,N_23906);
nor U24739 (N_24739,N_23344,N_23779);
or U24740 (N_24740,N_23659,N_23713);
nand U24741 (N_24741,N_23766,N_23218);
and U24742 (N_24742,N_23543,N_23682);
nand U24743 (N_24743,N_23437,N_23506);
xor U24744 (N_24744,N_23053,N_23146);
xor U24745 (N_24745,N_23052,N_23578);
xnor U24746 (N_24746,N_23878,N_23707);
nor U24747 (N_24747,N_23461,N_23496);
and U24748 (N_24748,N_23019,N_23643);
nor U24749 (N_24749,N_23612,N_23602);
or U24750 (N_24750,N_23046,N_23878);
xor U24751 (N_24751,N_23940,N_23274);
nand U24752 (N_24752,N_23371,N_23527);
nand U24753 (N_24753,N_23145,N_23040);
or U24754 (N_24754,N_23747,N_23333);
xor U24755 (N_24755,N_23784,N_23033);
nor U24756 (N_24756,N_23964,N_23737);
nand U24757 (N_24757,N_23031,N_23560);
xnor U24758 (N_24758,N_23247,N_23386);
or U24759 (N_24759,N_23148,N_23524);
xor U24760 (N_24760,N_23682,N_23852);
nor U24761 (N_24761,N_23216,N_23955);
and U24762 (N_24762,N_23913,N_23100);
and U24763 (N_24763,N_23178,N_23288);
or U24764 (N_24764,N_23863,N_23132);
nand U24765 (N_24765,N_23829,N_23466);
and U24766 (N_24766,N_23775,N_23995);
and U24767 (N_24767,N_23137,N_23356);
and U24768 (N_24768,N_23102,N_23415);
nor U24769 (N_24769,N_23736,N_23226);
nor U24770 (N_24770,N_23966,N_23809);
and U24771 (N_24771,N_23071,N_23673);
and U24772 (N_24772,N_23299,N_23238);
xor U24773 (N_24773,N_23465,N_23788);
nor U24774 (N_24774,N_23792,N_23115);
nor U24775 (N_24775,N_23771,N_23447);
nand U24776 (N_24776,N_23247,N_23083);
nand U24777 (N_24777,N_23701,N_23703);
or U24778 (N_24778,N_23422,N_23545);
xor U24779 (N_24779,N_23280,N_23798);
nand U24780 (N_24780,N_23368,N_23378);
nor U24781 (N_24781,N_23595,N_23071);
and U24782 (N_24782,N_23136,N_23180);
nand U24783 (N_24783,N_23036,N_23633);
or U24784 (N_24784,N_23087,N_23700);
or U24785 (N_24785,N_23964,N_23490);
or U24786 (N_24786,N_23065,N_23186);
or U24787 (N_24787,N_23418,N_23010);
or U24788 (N_24788,N_23356,N_23209);
and U24789 (N_24789,N_23431,N_23298);
nand U24790 (N_24790,N_23575,N_23062);
nand U24791 (N_24791,N_23914,N_23222);
xnor U24792 (N_24792,N_23237,N_23132);
xor U24793 (N_24793,N_23632,N_23658);
and U24794 (N_24794,N_23850,N_23896);
nor U24795 (N_24795,N_23846,N_23028);
and U24796 (N_24796,N_23250,N_23419);
nand U24797 (N_24797,N_23772,N_23153);
xor U24798 (N_24798,N_23107,N_23570);
and U24799 (N_24799,N_23169,N_23413);
or U24800 (N_24800,N_23032,N_23991);
nand U24801 (N_24801,N_23936,N_23996);
nor U24802 (N_24802,N_23756,N_23438);
xor U24803 (N_24803,N_23696,N_23782);
xnor U24804 (N_24804,N_23948,N_23027);
or U24805 (N_24805,N_23332,N_23487);
xor U24806 (N_24806,N_23209,N_23568);
xor U24807 (N_24807,N_23299,N_23467);
or U24808 (N_24808,N_23078,N_23431);
and U24809 (N_24809,N_23595,N_23978);
xnor U24810 (N_24810,N_23319,N_23078);
or U24811 (N_24811,N_23574,N_23529);
nor U24812 (N_24812,N_23067,N_23206);
nor U24813 (N_24813,N_23386,N_23865);
and U24814 (N_24814,N_23289,N_23124);
nor U24815 (N_24815,N_23304,N_23049);
nor U24816 (N_24816,N_23605,N_23040);
and U24817 (N_24817,N_23855,N_23188);
or U24818 (N_24818,N_23879,N_23144);
and U24819 (N_24819,N_23126,N_23340);
xnor U24820 (N_24820,N_23096,N_23985);
or U24821 (N_24821,N_23598,N_23117);
nand U24822 (N_24822,N_23006,N_23226);
or U24823 (N_24823,N_23669,N_23658);
or U24824 (N_24824,N_23579,N_23694);
nand U24825 (N_24825,N_23524,N_23806);
nand U24826 (N_24826,N_23176,N_23570);
xor U24827 (N_24827,N_23658,N_23136);
and U24828 (N_24828,N_23983,N_23401);
xnor U24829 (N_24829,N_23234,N_23863);
and U24830 (N_24830,N_23688,N_23735);
nand U24831 (N_24831,N_23962,N_23583);
nand U24832 (N_24832,N_23218,N_23308);
and U24833 (N_24833,N_23156,N_23447);
nor U24834 (N_24834,N_23988,N_23133);
or U24835 (N_24835,N_23429,N_23854);
nor U24836 (N_24836,N_23536,N_23444);
nor U24837 (N_24837,N_23761,N_23274);
or U24838 (N_24838,N_23014,N_23219);
nor U24839 (N_24839,N_23728,N_23534);
xnor U24840 (N_24840,N_23977,N_23633);
nor U24841 (N_24841,N_23446,N_23256);
nor U24842 (N_24842,N_23602,N_23925);
or U24843 (N_24843,N_23990,N_23101);
and U24844 (N_24844,N_23079,N_23540);
and U24845 (N_24845,N_23984,N_23546);
xor U24846 (N_24846,N_23924,N_23508);
nand U24847 (N_24847,N_23802,N_23531);
nand U24848 (N_24848,N_23289,N_23753);
or U24849 (N_24849,N_23312,N_23182);
and U24850 (N_24850,N_23894,N_23972);
and U24851 (N_24851,N_23140,N_23466);
and U24852 (N_24852,N_23973,N_23234);
nor U24853 (N_24853,N_23311,N_23412);
nand U24854 (N_24854,N_23067,N_23730);
xnor U24855 (N_24855,N_23697,N_23790);
and U24856 (N_24856,N_23978,N_23424);
nor U24857 (N_24857,N_23135,N_23207);
or U24858 (N_24858,N_23457,N_23093);
nand U24859 (N_24859,N_23935,N_23136);
nor U24860 (N_24860,N_23198,N_23211);
nor U24861 (N_24861,N_23673,N_23099);
and U24862 (N_24862,N_23817,N_23193);
and U24863 (N_24863,N_23986,N_23014);
and U24864 (N_24864,N_23351,N_23378);
nor U24865 (N_24865,N_23790,N_23592);
xor U24866 (N_24866,N_23685,N_23079);
nand U24867 (N_24867,N_23923,N_23429);
nand U24868 (N_24868,N_23817,N_23783);
nand U24869 (N_24869,N_23265,N_23726);
and U24870 (N_24870,N_23470,N_23957);
or U24871 (N_24871,N_23250,N_23077);
or U24872 (N_24872,N_23831,N_23035);
nand U24873 (N_24873,N_23558,N_23590);
nor U24874 (N_24874,N_23550,N_23981);
nor U24875 (N_24875,N_23562,N_23568);
and U24876 (N_24876,N_23223,N_23052);
or U24877 (N_24877,N_23428,N_23770);
or U24878 (N_24878,N_23791,N_23234);
xnor U24879 (N_24879,N_23780,N_23751);
nor U24880 (N_24880,N_23640,N_23335);
nor U24881 (N_24881,N_23519,N_23847);
and U24882 (N_24882,N_23194,N_23576);
xnor U24883 (N_24883,N_23931,N_23899);
nor U24884 (N_24884,N_23399,N_23909);
xnor U24885 (N_24885,N_23720,N_23268);
nor U24886 (N_24886,N_23433,N_23263);
xnor U24887 (N_24887,N_23368,N_23927);
nor U24888 (N_24888,N_23151,N_23566);
and U24889 (N_24889,N_23842,N_23423);
or U24890 (N_24890,N_23057,N_23804);
nor U24891 (N_24891,N_23625,N_23432);
or U24892 (N_24892,N_23830,N_23851);
and U24893 (N_24893,N_23725,N_23006);
nand U24894 (N_24894,N_23793,N_23497);
nor U24895 (N_24895,N_23581,N_23725);
nand U24896 (N_24896,N_23483,N_23368);
nor U24897 (N_24897,N_23707,N_23885);
and U24898 (N_24898,N_23925,N_23080);
nand U24899 (N_24899,N_23155,N_23992);
or U24900 (N_24900,N_23378,N_23946);
and U24901 (N_24901,N_23486,N_23120);
and U24902 (N_24902,N_23835,N_23118);
nor U24903 (N_24903,N_23730,N_23338);
nand U24904 (N_24904,N_23792,N_23694);
and U24905 (N_24905,N_23346,N_23571);
or U24906 (N_24906,N_23337,N_23715);
xnor U24907 (N_24907,N_23689,N_23301);
nor U24908 (N_24908,N_23753,N_23406);
xnor U24909 (N_24909,N_23963,N_23455);
or U24910 (N_24910,N_23516,N_23884);
xnor U24911 (N_24911,N_23873,N_23800);
nand U24912 (N_24912,N_23300,N_23260);
or U24913 (N_24913,N_23304,N_23361);
or U24914 (N_24914,N_23616,N_23323);
nand U24915 (N_24915,N_23063,N_23715);
and U24916 (N_24916,N_23799,N_23333);
or U24917 (N_24917,N_23634,N_23542);
or U24918 (N_24918,N_23509,N_23363);
xnor U24919 (N_24919,N_23429,N_23922);
or U24920 (N_24920,N_23299,N_23375);
and U24921 (N_24921,N_23143,N_23021);
or U24922 (N_24922,N_23313,N_23571);
nor U24923 (N_24923,N_23213,N_23880);
nor U24924 (N_24924,N_23447,N_23713);
and U24925 (N_24925,N_23550,N_23163);
and U24926 (N_24926,N_23586,N_23270);
nand U24927 (N_24927,N_23762,N_23284);
xnor U24928 (N_24928,N_23325,N_23281);
and U24929 (N_24929,N_23459,N_23449);
xor U24930 (N_24930,N_23462,N_23007);
or U24931 (N_24931,N_23473,N_23726);
nand U24932 (N_24932,N_23851,N_23175);
and U24933 (N_24933,N_23080,N_23096);
nor U24934 (N_24934,N_23305,N_23506);
or U24935 (N_24935,N_23942,N_23511);
nand U24936 (N_24936,N_23395,N_23519);
or U24937 (N_24937,N_23706,N_23424);
nand U24938 (N_24938,N_23532,N_23258);
nand U24939 (N_24939,N_23955,N_23963);
or U24940 (N_24940,N_23340,N_23579);
nand U24941 (N_24941,N_23196,N_23236);
xor U24942 (N_24942,N_23945,N_23634);
nor U24943 (N_24943,N_23522,N_23029);
nor U24944 (N_24944,N_23842,N_23437);
nor U24945 (N_24945,N_23584,N_23703);
or U24946 (N_24946,N_23762,N_23034);
nor U24947 (N_24947,N_23333,N_23102);
xnor U24948 (N_24948,N_23945,N_23677);
or U24949 (N_24949,N_23377,N_23028);
and U24950 (N_24950,N_23188,N_23076);
nand U24951 (N_24951,N_23709,N_23051);
or U24952 (N_24952,N_23442,N_23503);
or U24953 (N_24953,N_23103,N_23096);
xor U24954 (N_24954,N_23045,N_23844);
nor U24955 (N_24955,N_23549,N_23556);
nand U24956 (N_24956,N_23247,N_23040);
nand U24957 (N_24957,N_23124,N_23719);
nor U24958 (N_24958,N_23838,N_23218);
nand U24959 (N_24959,N_23394,N_23610);
nand U24960 (N_24960,N_23599,N_23807);
nor U24961 (N_24961,N_23662,N_23891);
nand U24962 (N_24962,N_23847,N_23131);
nor U24963 (N_24963,N_23512,N_23872);
xor U24964 (N_24964,N_23335,N_23194);
and U24965 (N_24965,N_23090,N_23255);
and U24966 (N_24966,N_23809,N_23986);
or U24967 (N_24967,N_23207,N_23405);
nor U24968 (N_24968,N_23562,N_23518);
xor U24969 (N_24969,N_23656,N_23562);
xor U24970 (N_24970,N_23357,N_23347);
or U24971 (N_24971,N_23066,N_23702);
and U24972 (N_24972,N_23486,N_23009);
and U24973 (N_24973,N_23987,N_23147);
and U24974 (N_24974,N_23723,N_23703);
nor U24975 (N_24975,N_23496,N_23372);
nand U24976 (N_24976,N_23668,N_23484);
xnor U24977 (N_24977,N_23008,N_23951);
nand U24978 (N_24978,N_23809,N_23627);
nor U24979 (N_24979,N_23480,N_23105);
nand U24980 (N_24980,N_23545,N_23394);
or U24981 (N_24981,N_23835,N_23557);
and U24982 (N_24982,N_23436,N_23066);
nor U24983 (N_24983,N_23832,N_23740);
or U24984 (N_24984,N_23658,N_23965);
nand U24985 (N_24985,N_23639,N_23339);
and U24986 (N_24986,N_23213,N_23254);
or U24987 (N_24987,N_23315,N_23788);
nand U24988 (N_24988,N_23744,N_23838);
nor U24989 (N_24989,N_23459,N_23414);
xor U24990 (N_24990,N_23601,N_23270);
nor U24991 (N_24991,N_23703,N_23142);
xnor U24992 (N_24992,N_23303,N_23792);
and U24993 (N_24993,N_23345,N_23904);
nor U24994 (N_24994,N_23326,N_23828);
nor U24995 (N_24995,N_23981,N_23379);
or U24996 (N_24996,N_23581,N_23756);
or U24997 (N_24997,N_23131,N_23426);
or U24998 (N_24998,N_23404,N_23102);
or U24999 (N_24999,N_23554,N_23795);
nand U25000 (N_25000,N_24079,N_24025);
and U25001 (N_25001,N_24236,N_24456);
nand U25002 (N_25002,N_24747,N_24218);
and U25003 (N_25003,N_24563,N_24568);
or U25004 (N_25004,N_24889,N_24624);
xnor U25005 (N_25005,N_24217,N_24420);
nand U25006 (N_25006,N_24931,N_24907);
or U25007 (N_25007,N_24520,N_24390);
xor U25008 (N_25008,N_24799,N_24460);
nand U25009 (N_25009,N_24119,N_24559);
and U25010 (N_25010,N_24816,N_24776);
nor U25011 (N_25011,N_24637,N_24922);
nor U25012 (N_25012,N_24955,N_24906);
xnor U25013 (N_25013,N_24346,N_24329);
xnor U25014 (N_25014,N_24232,N_24483);
nand U25015 (N_25015,N_24485,N_24519);
or U25016 (N_25016,N_24598,N_24846);
xnor U25017 (N_25017,N_24844,N_24579);
nand U25018 (N_25018,N_24547,N_24748);
or U25019 (N_25019,N_24599,N_24773);
nor U25020 (N_25020,N_24060,N_24479);
and U25021 (N_25021,N_24214,N_24762);
or U25022 (N_25022,N_24076,N_24139);
nor U25023 (N_25023,N_24379,N_24251);
nand U25024 (N_25024,N_24399,N_24198);
xor U25025 (N_25025,N_24199,N_24444);
xnor U25026 (N_25026,N_24265,N_24695);
and U25027 (N_25027,N_24133,N_24652);
nand U25028 (N_25028,N_24136,N_24496);
xnor U25029 (N_25029,N_24848,N_24521);
nor U25030 (N_25030,N_24101,N_24548);
nor U25031 (N_25031,N_24942,N_24877);
nand U25032 (N_25032,N_24336,N_24266);
nand U25033 (N_25033,N_24711,N_24604);
and U25034 (N_25034,N_24663,N_24386);
xnor U25035 (N_25035,N_24036,N_24808);
and U25036 (N_25036,N_24222,N_24059);
or U25037 (N_25037,N_24699,N_24007);
nand U25038 (N_25038,N_24583,N_24756);
or U25039 (N_25039,N_24032,N_24845);
or U25040 (N_25040,N_24304,N_24971);
and U25041 (N_25041,N_24383,N_24960);
nand U25042 (N_25042,N_24967,N_24099);
xor U25043 (N_25043,N_24913,N_24991);
nand U25044 (N_25044,N_24350,N_24226);
xnor U25045 (N_25045,N_24785,N_24154);
nor U25046 (N_25046,N_24487,N_24687);
xnor U25047 (N_25047,N_24979,N_24162);
xor U25048 (N_25048,N_24309,N_24412);
or U25049 (N_25049,N_24855,N_24543);
nor U25050 (N_25050,N_24504,N_24181);
nor U25051 (N_25051,N_24393,N_24900);
nand U25052 (N_25052,N_24333,N_24859);
nand U25053 (N_25053,N_24603,N_24433);
nand U25054 (N_25054,N_24580,N_24084);
and U25055 (N_25055,N_24153,N_24308);
nand U25056 (N_25056,N_24499,N_24657);
nand U25057 (N_25057,N_24155,N_24052);
and U25058 (N_25058,N_24502,N_24010);
nor U25059 (N_25059,N_24753,N_24377);
nor U25060 (N_25060,N_24676,N_24810);
and U25061 (N_25061,N_24680,N_24622);
or U25062 (N_25062,N_24229,N_24966);
and U25063 (N_25063,N_24722,N_24372);
nand U25064 (N_25064,N_24546,N_24490);
nand U25065 (N_25065,N_24754,N_24696);
xor U25066 (N_25066,N_24020,N_24213);
or U25067 (N_25067,N_24220,N_24981);
xnor U25068 (N_25068,N_24190,N_24817);
or U25069 (N_25069,N_24999,N_24946);
xor U25070 (N_25070,N_24736,N_24164);
and U25071 (N_25071,N_24638,N_24518);
xor U25072 (N_25072,N_24741,N_24920);
nor U25073 (N_25073,N_24283,N_24883);
and U25074 (N_25074,N_24876,N_24495);
nand U25075 (N_25075,N_24879,N_24128);
or U25076 (N_25076,N_24047,N_24361);
and U25077 (N_25077,N_24488,N_24468);
xor U25078 (N_25078,N_24448,N_24550);
or U25079 (N_25079,N_24824,N_24608);
or U25080 (N_25080,N_24726,N_24111);
nand U25081 (N_25081,N_24963,N_24642);
and U25082 (N_25082,N_24807,N_24031);
or U25083 (N_25083,N_24268,N_24918);
xnor U25084 (N_25084,N_24057,N_24985);
nor U25085 (N_25085,N_24443,N_24789);
nor U25086 (N_25086,N_24328,N_24898);
or U25087 (N_25087,N_24183,N_24078);
nor U25088 (N_25088,N_24203,N_24860);
nor U25089 (N_25089,N_24277,N_24391);
xor U25090 (N_25090,N_24506,N_24639);
or U25091 (N_25091,N_24800,N_24558);
nand U25092 (N_25092,N_24760,N_24668);
or U25093 (N_25093,N_24843,N_24110);
nor U25094 (N_25094,N_24742,N_24175);
nor U25095 (N_25095,N_24780,N_24046);
nor U25096 (N_25096,N_24288,N_24146);
nor U25097 (N_25097,N_24787,N_24949);
nand U25098 (N_25098,N_24893,N_24545);
or U25099 (N_25099,N_24995,N_24834);
and U25100 (N_25100,N_24919,N_24435);
or U25101 (N_25101,N_24738,N_24027);
nand U25102 (N_25102,N_24278,N_24511);
and U25103 (N_25103,N_24744,N_24818);
xor U25104 (N_25104,N_24500,N_24730);
nor U25105 (N_25105,N_24231,N_24235);
nor U25106 (N_25106,N_24196,N_24739);
xor U25107 (N_25107,N_24087,N_24835);
nand U25108 (N_25108,N_24318,N_24296);
nand U25109 (N_25109,N_24857,N_24168);
or U25110 (N_25110,N_24873,N_24063);
nand U25111 (N_25111,N_24248,N_24163);
nor U25112 (N_25112,N_24928,N_24575);
and U25113 (N_25113,N_24396,N_24180);
nand U25114 (N_25114,N_24238,N_24453);
nand U25115 (N_25115,N_24147,N_24690);
xnor U25116 (N_25116,N_24825,N_24040);
or U25117 (N_25117,N_24797,N_24142);
or U25118 (N_25118,N_24974,N_24927);
nor U25119 (N_25119,N_24150,N_24082);
nor U25120 (N_25120,N_24132,N_24322);
nor U25121 (N_25121,N_24300,N_24659);
nor U25122 (N_25122,N_24707,N_24182);
and U25123 (N_25123,N_24677,N_24184);
nor U25124 (N_25124,N_24746,N_24279);
and U25125 (N_25125,N_24679,N_24821);
or U25126 (N_25126,N_24426,N_24571);
or U25127 (N_25127,N_24786,N_24578);
nand U25128 (N_25128,N_24704,N_24529);
xor U25129 (N_25129,N_24752,N_24457);
xor U25130 (N_25130,N_24778,N_24104);
nand U25131 (N_25131,N_24282,N_24023);
and U25132 (N_25132,N_24206,N_24887);
nor U25133 (N_25133,N_24640,N_24703);
or U25134 (N_25134,N_24643,N_24339);
xnor U25135 (N_25135,N_24874,N_24655);
and U25136 (N_25136,N_24992,N_24621);
or U25137 (N_25137,N_24498,N_24536);
xor U25138 (N_25138,N_24437,N_24597);
nor U25139 (N_25139,N_24173,N_24714);
and U25140 (N_25140,N_24713,N_24839);
or U25141 (N_25141,N_24853,N_24523);
nor U25142 (N_25142,N_24812,N_24374);
nand U25143 (N_25143,N_24630,N_24472);
nand U25144 (N_25144,N_24033,N_24872);
nor U25145 (N_25145,N_24403,N_24856);
nand U25146 (N_25146,N_24418,N_24968);
nand U25147 (N_25147,N_24256,N_24708);
xor U25148 (N_25148,N_24765,N_24298);
nand U25149 (N_25149,N_24130,N_24179);
nor U25150 (N_25150,N_24187,N_24455);
xor U25151 (N_25151,N_24494,N_24775);
or U25152 (N_25152,N_24075,N_24449);
xnor U25153 (N_25153,N_24021,N_24351);
and U25154 (N_25154,N_24434,N_24745);
and U25155 (N_25155,N_24662,N_24683);
xnor U25156 (N_25156,N_24569,N_24570);
nand U25157 (N_25157,N_24096,N_24410);
or U25158 (N_25158,N_24541,N_24178);
and U25159 (N_25159,N_24343,N_24505);
xor U25160 (N_25160,N_24287,N_24359);
nand U25161 (N_25161,N_24552,N_24826);
nand U25162 (N_25162,N_24273,N_24295);
nand U25163 (N_25163,N_24000,N_24737);
nand U25164 (N_25164,N_24152,N_24596);
and U25165 (N_25165,N_24881,N_24861);
and U25166 (N_25166,N_24670,N_24530);
xor U25167 (N_25167,N_24194,N_24743);
xor U25168 (N_25168,N_24688,N_24782);
or U25169 (N_25169,N_24385,N_24332);
xnor U25170 (N_25170,N_24016,N_24719);
and U25171 (N_25171,N_24117,N_24779);
and U25172 (N_25172,N_24042,N_24461);
xor U25173 (N_25173,N_24958,N_24145);
or U25174 (N_25174,N_24066,N_24689);
nor U25175 (N_25175,N_24327,N_24430);
xor U25176 (N_25176,N_24069,N_24088);
nor U25177 (N_25177,N_24606,N_24935);
or U25178 (N_25178,N_24041,N_24253);
or U25179 (N_25179,N_24431,N_24647);
nor U25180 (N_25180,N_24769,N_24950);
and U25181 (N_25181,N_24909,N_24636);
and U25182 (N_25182,N_24901,N_24944);
or U25183 (N_25183,N_24885,N_24667);
nor U25184 (N_25184,N_24212,N_24090);
xor U25185 (N_25185,N_24467,N_24915);
xnor U25186 (N_25186,N_24009,N_24055);
nand U25187 (N_25187,N_24865,N_24890);
nor U25188 (N_25188,N_24718,N_24126);
and U25189 (N_25189,N_24029,N_24904);
xor U25190 (N_25190,N_24665,N_24252);
or U25191 (N_25191,N_24698,N_24131);
nor U25192 (N_25192,N_24788,N_24367);
and U25193 (N_25193,N_24177,N_24650);
and U25194 (N_25194,N_24097,N_24709);
nor U25195 (N_25195,N_24053,N_24225);
and U25196 (N_25196,N_24802,N_24849);
xor U25197 (N_25197,N_24261,N_24581);
nand U25198 (N_25198,N_24422,N_24982);
or U25199 (N_25199,N_24589,N_24340);
and U25200 (N_25200,N_24532,N_24534);
nor U25201 (N_25201,N_24983,N_24602);
nand U25202 (N_25202,N_24034,N_24167);
xnor U25203 (N_25203,N_24715,N_24930);
nor U25204 (N_25204,N_24100,N_24089);
and U25205 (N_25205,N_24115,N_24289);
or U25206 (N_25206,N_24701,N_24691);
xnor U25207 (N_25207,N_24735,N_24413);
and U25208 (N_25208,N_24867,N_24174);
and U25209 (N_25209,N_24989,N_24056);
nand U25210 (N_25210,N_24980,N_24903);
nand U25211 (N_25211,N_24121,N_24317);
xnor U25212 (N_25212,N_24245,N_24347);
xor U25213 (N_25213,N_24671,N_24093);
and U25214 (N_25214,N_24204,N_24564);
or U25215 (N_25215,N_24037,N_24940);
nor U25216 (N_25216,N_24555,N_24415);
and U25217 (N_25217,N_24706,N_24666);
or U25218 (N_25218,N_24116,N_24628);
xor U25219 (N_25219,N_24124,N_24244);
or U25220 (N_25220,N_24697,N_24869);
or U25221 (N_25221,N_24573,N_24134);
nand U25222 (N_25222,N_24629,N_24215);
nand U25223 (N_25223,N_24712,N_24939);
nor U25224 (N_25224,N_24355,N_24961);
and U25225 (N_25225,N_24384,N_24401);
or U25226 (N_25226,N_24127,N_24358);
nor U25227 (N_25227,N_24072,N_24414);
or U25228 (N_25228,N_24006,N_24407);
and U25229 (N_25229,N_24122,N_24591);
or U25230 (N_25230,N_24705,N_24243);
nand U25231 (N_25231,N_24623,N_24423);
and U25232 (N_25232,N_24299,N_24686);
xor U25233 (N_25233,N_24917,N_24463);
nand U25234 (N_25234,N_24725,N_24549);
or U25235 (N_25235,N_24613,N_24970);
nand U25236 (N_25236,N_24230,N_24454);
and U25237 (N_25237,N_24284,N_24450);
nand U25238 (N_25238,N_24445,N_24137);
xor U25239 (N_25239,N_24424,N_24442);
or U25240 (N_25240,N_24319,N_24905);
and U25241 (N_25241,N_24428,N_24896);
nor U25242 (N_25242,N_24345,N_24934);
or U25243 (N_25243,N_24929,N_24984);
nor U25244 (N_25244,N_24969,N_24395);
xor U25245 (N_25245,N_24071,N_24517);
and U25246 (N_25246,N_24158,N_24674);
or U25247 (N_25247,N_24313,N_24176);
xnor U25248 (N_25248,N_24717,N_24723);
xor U25249 (N_25249,N_24470,N_24798);
nand U25250 (N_25250,N_24790,N_24216);
nand U25251 (N_25251,N_24392,N_24321);
nand U25252 (N_25252,N_24975,N_24616);
nor U25253 (N_25253,N_24833,N_24143);
or U25254 (N_25254,N_24664,N_24397);
or U25255 (N_25255,N_24610,N_24125);
nor U25256 (N_25256,N_24702,N_24469);
nand U25257 (N_25257,N_24354,N_24886);
nand U25258 (N_25258,N_24440,N_24476);
or U25259 (N_25259,N_24378,N_24951);
nand U25260 (N_25260,N_24525,N_24830);
and U25261 (N_25261,N_24774,N_24429);
or U25262 (N_25262,N_24405,N_24382);
and U25263 (N_25263,N_24672,N_24977);
nand U25264 (N_25264,N_24813,N_24740);
or U25265 (N_25265,N_24172,N_24768);
or U25266 (N_25266,N_24312,N_24409);
xnor U25267 (N_25267,N_24334,N_24827);
nor U25268 (N_25268,N_24223,N_24112);
xnor U25269 (N_25269,N_24030,N_24540);
nand U25270 (N_25270,N_24751,N_24478);
or U25271 (N_25271,N_24406,N_24039);
and U25272 (N_25272,N_24263,N_24987);
and U25273 (N_25273,N_24882,N_24400);
nand U25274 (N_25274,N_24588,N_24627);
nand U25275 (N_25275,N_24866,N_24280);
xor U25276 (N_25276,N_24054,N_24700);
nor U25277 (N_25277,N_24526,N_24065);
xnor U25278 (N_25278,N_24556,N_24480);
nand U25279 (N_25279,N_24446,N_24763);
or U25280 (N_25280,N_24362,N_24542);
nand U25281 (N_25281,N_24720,N_24149);
nor U25282 (N_25282,N_24258,N_24048);
and U25283 (N_25283,N_24993,N_24038);
and U25284 (N_25284,N_24475,N_24024);
or U25285 (N_25285,N_24380,N_24432);
xor U25286 (N_25286,N_24281,N_24310);
nor U25287 (N_25287,N_24938,N_24749);
and U25288 (N_25288,N_24294,N_24863);
and U25289 (N_25289,N_24408,N_24260);
or U25290 (N_25290,N_24693,N_24019);
nand U25291 (N_25291,N_24911,N_24233);
or U25292 (N_25292,N_24916,N_24341);
xor U25293 (N_25293,N_24962,N_24398);
and U25294 (N_25294,N_24612,N_24095);
and U25295 (N_25295,N_24394,N_24211);
nand U25296 (N_25296,N_24489,N_24574);
nor U25297 (N_25297,N_24513,N_24533);
or U25298 (N_25298,N_24794,N_24978);
or U25299 (N_25299,N_24767,N_24441);
or U25300 (N_25300,N_24360,N_24822);
nand U25301 (N_25301,N_24803,N_24107);
or U25302 (N_25302,N_24208,N_24871);
nor U25303 (N_25303,N_24365,N_24477);
and U25304 (N_25304,N_24957,N_24972);
and U25305 (N_25305,N_24337,N_24854);
nand U25306 (N_25306,N_24750,N_24815);
xor U25307 (N_25307,N_24675,N_24535);
nor U25308 (N_25308,N_24017,N_24649);
nand U25309 (N_25309,N_24419,N_24926);
or U25310 (N_25310,N_24820,N_24381);
xor U25311 (N_25311,N_24274,N_24338);
xnor U25312 (N_25312,N_24584,N_24207);
or U25313 (N_25313,N_24986,N_24595);
nand U25314 (N_25314,N_24895,N_24811);
xnor U25315 (N_25315,N_24988,N_24388);
xor U25316 (N_25316,N_24402,N_24404);
nand U25317 (N_25317,N_24796,N_24503);
or U25318 (N_25318,N_24561,N_24587);
and U25319 (N_25319,N_24241,N_24114);
or U25320 (N_25320,N_24912,N_24936);
or U25321 (N_25321,N_24452,N_24755);
nor U25322 (N_25322,N_24050,N_24086);
and U25323 (N_25323,N_24614,N_24366);
and U25324 (N_25324,N_24259,N_24538);
nor U25325 (N_25325,N_24925,N_24899);
nor U25326 (N_25326,N_24759,N_24320);
nor U25327 (N_25327,N_24493,N_24043);
nand U25328 (N_25328,N_24528,N_24766);
xnor U25329 (N_25329,N_24976,N_24497);
or U25330 (N_25330,N_24140,N_24996);
xnor U25331 (N_25331,N_24847,N_24080);
nor U25332 (N_25332,N_24937,N_24305);
nand U25333 (N_25333,N_24837,N_24344);
nor U25334 (N_25334,N_24908,N_24159);
or U25335 (N_25335,N_24836,N_24537);
and U25336 (N_25336,N_24269,N_24829);
and U25337 (N_25337,N_24501,N_24648);
or U25338 (N_25338,N_24221,N_24094);
xor U25339 (N_25339,N_24692,N_24293);
nor U25340 (N_25340,N_24716,N_24840);
nor U25341 (N_25341,N_24777,N_24474);
nand U25342 (N_25342,N_24678,N_24427);
nand U25343 (N_25343,N_24921,N_24436);
and U25344 (N_25344,N_24466,N_24161);
and U25345 (N_25345,N_24932,N_24831);
xnor U25346 (N_25346,N_24369,N_24077);
and U25347 (N_25347,N_24586,N_24144);
and U25348 (N_25348,N_24291,N_24660);
and U25349 (N_25349,N_24531,N_24838);
nand U25350 (N_25350,N_24192,N_24209);
nor U25351 (N_25351,N_24108,N_24013);
and U25352 (N_25352,N_24633,N_24758);
nand U25353 (N_25353,N_24102,N_24870);
or U25354 (N_25354,N_24492,N_24105);
and U25355 (N_25355,N_24770,N_24626);
nor U25356 (N_25356,N_24109,N_24539);
nand U25357 (N_25357,N_24619,N_24370);
nand U25358 (N_25358,N_24193,N_24510);
or U25359 (N_25359,N_24471,N_24828);
or U25360 (N_25360,N_24814,N_24673);
or U25361 (N_25361,N_24416,N_24092);
xnor U25362 (N_25362,N_24314,N_24651);
xor U25363 (N_25363,N_24933,N_24353);
and U25364 (N_25364,N_24884,N_24389);
xnor U25365 (N_25365,N_24601,N_24731);
xnor U25366 (N_25366,N_24809,N_24959);
nor U25367 (N_25367,N_24324,N_24465);
xnor U25368 (N_25368,N_24953,N_24880);
and U25369 (N_25369,N_24275,N_24868);
xnor U25370 (N_25370,N_24894,N_24438);
and U25371 (N_25371,N_24364,N_24311);
or U25372 (N_25372,N_24507,N_24074);
xor U25373 (N_25373,N_24166,N_24165);
xor U25374 (N_25374,N_24615,N_24286);
nand U25375 (N_25375,N_24611,N_24473);
nand U25376 (N_25376,N_24335,N_24348);
nand U25377 (N_25377,N_24491,N_24990);
xnor U25378 (N_25378,N_24635,N_24325);
xor U25379 (N_25379,N_24734,N_24594);
xor U25380 (N_25380,N_24315,N_24878);
nor U25381 (N_25381,N_24710,N_24018);
nand U25382 (N_25382,N_24262,N_24061);
nor U25383 (N_25383,N_24160,N_24656);
nor U25384 (N_25384,N_24795,N_24948);
nand U25385 (N_25385,N_24451,N_24783);
and U25386 (N_25386,N_24120,N_24947);
nor U25387 (N_25387,N_24285,N_24001);
or U25388 (N_25388,N_24417,N_24342);
or U25389 (N_25389,N_24512,N_24439);
nand U25390 (N_25390,N_24205,N_24290);
nor U25391 (N_25391,N_24242,N_24026);
or U25392 (N_25392,N_24585,N_24793);
and U25393 (N_25393,N_24234,N_24562);
nor U25394 (N_25394,N_24250,N_24051);
xor U25395 (N_25395,N_24842,N_24508);
or U25396 (N_25396,N_24669,N_24484);
and U25397 (N_25397,N_24577,N_24851);
nor U25398 (N_25398,N_24352,N_24732);
xnor U25399 (N_25399,N_24157,N_24368);
and U25400 (N_25400,N_24085,N_24965);
and U25401 (N_25401,N_24188,N_24875);
or U25402 (N_25402,N_24910,N_24576);
xor U25403 (N_25403,N_24482,N_24219);
or U25404 (N_25404,N_24363,N_24070);
nand U25405 (N_25405,N_24002,N_24761);
nand U25406 (N_25406,N_24565,N_24135);
or U25407 (N_25407,N_24553,N_24098);
nand U25408 (N_25408,N_24004,N_24527);
or U25409 (N_25409,N_24850,N_24447);
xor U25410 (N_25410,N_24864,N_24197);
nand U25411 (N_25411,N_24681,N_24271);
nand U25412 (N_25412,N_24330,N_24113);
or U25413 (N_25413,N_24301,N_24923);
xnor U25414 (N_25414,N_24654,N_24727);
and U25415 (N_25415,N_24247,N_24185);
nand U25416 (N_25416,N_24103,N_24973);
xor U25417 (N_25417,N_24356,N_24228);
nor U25418 (N_25418,N_24943,N_24592);
or U25419 (N_25419,N_24156,N_24852);
nand U25420 (N_25420,N_24272,N_24994);
or U25421 (N_25421,N_24653,N_24631);
nor U25422 (N_25422,N_24516,N_24891);
nor U25423 (N_25423,N_24632,N_24486);
nand U25424 (N_25424,N_24841,N_24306);
or U25425 (N_25425,N_24118,N_24224);
or U25426 (N_25426,N_24641,N_24645);
and U25427 (N_25427,N_24902,N_24522);
nor U25428 (N_25428,N_24141,N_24590);
nand U25429 (N_25429,N_24897,N_24003);
and U25430 (N_25430,N_24421,N_24249);
or U25431 (N_25431,N_24801,N_24728);
nand U25432 (N_25432,N_24123,N_24035);
and U25433 (N_25433,N_24805,N_24292);
or U25434 (N_25434,N_24239,N_24357);
nand U25435 (N_25435,N_24600,N_24459);
and U25436 (N_25436,N_24129,N_24264);
or U25437 (N_25437,N_24998,N_24151);
nor U25438 (N_25438,N_24685,N_24169);
nor U25439 (N_25439,N_24375,N_24832);
nor U25440 (N_25440,N_24582,N_24862);
nor U25441 (N_25441,N_24609,N_24551);
nand U25442 (N_25442,N_24515,N_24022);
or U25443 (N_25443,N_24138,N_24646);
nor U25444 (N_25444,N_24411,N_24952);
and U25445 (N_25445,N_24326,N_24011);
nor U25446 (N_25446,N_24189,N_24171);
xor U25447 (N_25447,N_24297,N_24764);
nand U25448 (N_25448,N_24081,N_24964);
nand U25449 (N_25449,N_24349,N_24307);
or U25450 (N_25450,N_24888,N_24956);
xnor U25451 (N_25451,N_24464,N_24781);
and U25452 (N_25452,N_24661,N_24012);
or U25453 (N_25453,N_24557,N_24892);
xnor U25454 (N_25454,N_24544,N_24554);
nor U25455 (N_25455,N_24791,N_24148);
and U25456 (N_25456,N_24387,N_24567);
xor U25457 (N_25457,N_24806,N_24634);
or U25458 (N_25458,N_24458,N_24724);
and U25459 (N_25459,N_24858,N_24625);
or U25460 (N_25460,N_24083,N_24607);
and U25461 (N_25461,N_24804,N_24049);
nor U25462 (N_25462,N_24593,N_24772);
xor U25463 (N_25463,N_24267,N_24015);
or U25464 (N_25464,N_24620,N_24210);
or U25465 (N_25465,N_24784,N_24658);
and U25466 (N_25466,N_24823,N_24373);
and U25467 (N_25467,N_24302,N_24276);
nor U25468 (N_25468,N_24201,N_24514);
and U25469 (N_25469,N_24462,N_24064);
nand U25470 (N_25470,N_24941,N_24091);
nand U25471 (N_25471,N_24331,N_24067);
and U25472 (N_25472,N_24371,N_24240);
xnor U25473 (N_25473,N_24694,N_24254);
and U25474 (N_25474,N_24014,N_24605);
xnor U25475 (N_25475,N_24246,N_24684);
nor U25476 (N_25476,N_24195,N_24425);
nor U25477 (N_25477,N_24068,N_24819);
or U25478 (N_25478,N_24062,N_24044);
and U25479 (N_25479,N_24005,N_24376);
xnor U25480 (N_25480,N_24729,N_24237);
nor U25481 (N_25481,N_24058,N_24028);
nand U25482 (N_25482,N_24924,N_24202);
xnor U25483 (N_25483,N_24524,N_24721);
nor U25484 (N_25484,N_24792,N_24191);
xnor U25485 (N_25485,N_24566,N_24303);
and U25486 (N_25486,N_24617,N_24045);
or U25487 (N_25487,N_24771,N_24997);
or U25488 (N_25488,N_24316,N_24618);
or U25489 (N_25489,N_24106,N_24227);
nor U25490 (N_25490,N_24945,N_24200);
nor U25491 (N_25491,N_24757,N_24954);
or U25492 (N_25492,N_24008,N_24572);
and U25493 (N_25493,N_24255,N_24186);
xor U25494 (N_25494,N_24323,N_24682);
nor U25495 (N_25495,N_24481,N_24914);
and U25496 (N_25496,N_24170,N_24270);
nor U25497 (N_25497,N_24073,N_24644);
xnor U25498 (N_25498,N_24509,N_24733);
nand U25499 (N_25499,N_24257,N_24560);
or U25500 (N_25500,N_24157,N_24802);
or U25501 (N_25501,N_24743,N_24096);
or U25502 (N_25502,N_24485,N_24870);
nand U25503 (N_25503,N_24729,N_24274);
and U25504 (N_25504,N_24743,N_24407);
nand U25505 (N_25505,N_24885,N_24035);
xor U25506 (N_25506,N_24391,N_24227);
nor U25507 (N_25507,N_24889,N_24600);
xnor U25508 (N_25508,N_24544,N_24994);
and U25509 (N_25509,N_24334,N_24757);
and U25510 (N_25510,N_24887,N_24012);
and U25511 (N_25511,N_24498,N_24683);
xor U25512 (N_25512,N_24030,N_24286);
nand U25513 (N_25513,N_24678,N_24218);
or U25514 (N_25514,N_24264,N_24955);
or U25515 (N_25515,N_24957,N_24217);
or U25516 (N_25516,N_24423,N_24935);
nand U25517 (N_25517,N_24784,N_24915);
and U25518 (N_25518,N_24615,N_24022);
nor U25519 (N_25519,N_24177,N_24762);
xor U25520 (N_25520,N_24007,N_24369);
nor U25521 (N_25521,N_24142,N_24172);
nor U25522 (N_25522,N_24642,N_24383);
nor U25523 (N_25523,N_24600,N_24181);
nand U25524 (N_25524,N_24101,N_24605);
or U25525 (N_25525,N_24590,N_24012);
nor U25526 (N_25526,N_24951,N_24687);
and U25527 (N_25527,N_24852,N_24331);
nor U25528 (N_25528,N_24583,N_24676);
xor U25529 (N_25529,N_24130,N_24837);
and U25530 (N_25530,N_24512,N_24194);
nor U25531 (N_25531,N_24627,N_24458);
and U25532 (N_25532,N_24634,N_24306);
or U25533 (N_25533,N_24500,N_24350);
and U25534 (N_25534,N_24411,N_24442);
or U25535 (N_25535,N_24520,N_24769);
or U25536 (N_25536,N_24724,N_24409);
and U25537 (N_25537,N_24861,N_24646);
nor U25538 (N_25538,N_24564,N_24575);
or U25539 (N_25539,N_24991,N_24200);
nand U25540 (N_25540,N_24182,N_24620);
nand U25541 (N_25541,N_24112,N_24738);
nand U25542 (N_25542,N_24942,N_24011);
or U25543 (N_25543,N_24849,N_24124);
or U25544 (N_25544,N_24808,N_24773);
and U25545 (N_25545,N_24077,N_24295);
nand U25546 (N_25546,N_24096,N_24048);
and U25547 (N_25547,N_24555,N_24501);
and U25548 (N_25548,N_24110,N_24331);
nor U25549 (N_25549,N_24138,N_24902);
nor U25550 (N_25550,N_24036,N_24169);
nor U25551 (N_25551,N_24511,N_24175);
or U25552 (N_25552,N_24766,N_24737);
or U25553 (N_25553,N_24538,N_24370);
xor U25554 (N_25554,N_24441,N_24766);
xnor U25555 (N_25555,N_24061,N_24342);
xnor U25556 (N_25556,N_24380,N_24424);
nor U25557 (N_25557,N_24137,N_24921);
nor U25558 (N_25558,N_24010,N_24054);
nand U25559 (N_25559,N_24983,N_24628);
nand U25560 (N_25560,N_24659,N_24735);
or U25561 (N_25561,N_24856,N_24395);
nor U25562 (N_25562,N_24325,N_24215);
and U25563 (N_25563,N_24743,N_24829);
and U25564 (N_25564,N_24283,N_24470);
or U25565 (N_25565,N_24053,N_24647);
xnor U25566 (N_25566,N_24991,N_24739);
or U25567 (N_25567,N_24684,N_24161);
xnor U25568 (N_25568,N_24976,N_24934);
nand U25569 (N_25569,N_24794,N_24589);
or U25570 (N_25570,N_24593,N_24443);
nor U25571 (N_25571,N_24521,N_24755);
and U25572 (N_25572,N_24520,N_24978);
nor U25573 (N_25573,N_24323,N_24916);
nand U25574 (N_25574,N_24203,N_24815);
or U25575 (N_25575,N_24799,N_24911);
nand U25576 (N_25576,N_24571,N_24963);
nor U25577 (N_25577,N_24742,N_24756);
nand U25578 (N_25578,N_24962,N_24541);
nor U25579 (N_25579,N_24744,N_24759);
and U25580 (N_25580,N_24392,N_24458);
or U25581 (N_25581,N_24467,N_24494);
nand U25582 (N_25582,N_24165,N_24919);
nor U25583 (N_25583,N_24431,N_24974);
nor U25584 (N_25584,N_24408,N_24697);
nor U25585 (N_25585,N_24581,N_24373);
nand U25586 (N_25586,N_24429,N_24434);
nand U25587 (N_25587,N_24972,N_24984);
and U25588 (N_25588,N_24620,N_24892);
or U25589 (N_25589,N_24538,N_24699);
xor U25590 (N_25590,N_24664,N_24049);
xor U25591 (N_25591,N_24474,N_24101);
xor U25592 (N_25592,N_24856,N_24181);
or U25593 (N_25593,N_24677,N_24394);
nand U25594 (N_25594,N_24011,N_24283);
or U25595 (N_25595,N_24484,N_24291);
xor U25596 (N_25596,N_24774,N_24346);
or U25597 (N_25597,N_24433,N_24076);
and U25598 (N_25598,N_24605,N_24565);
and U25599 (N_25599,N_24044,N_24069);
nand U25600 (N_25600,N_24323,N_24340);
nand U25601 (N_25601,N_24068,N_24485);
nand U25602 (N_25602,N_24951,N_24228);
or U25603 (N_25603,N_24536,N_24104);
xnor U25604 (N_25604,N_24558,N_24339);
nand U25605 (N_25605,N_24827,N_24830);
nor U25606 (N_25606,N_24078,N_24184);
or U25607 (N_25607,N_24931,N_24220);
nand U25608 (N_25608,N_24802,N_24148);
xnor U25609 (N_25609,N_24395,N_24524);
and U25610 (N_25610,N_24783,N_24763);
nand U25611 (N_25611,N_24670,N_24579);
nand U25612 (N_25612,N_24734,N_24054);
or U25613 (N_25613,N_24709,N_24351);
xor U25614 (N_25614,N_24848,N_24843);
nor U25615 (N_25615,N_24016,N_24907);
and U25616 (N_25616,N_24257,N_24139);
or U25617 (N_25617,N_24550,N_24822);
nand U25618 (N_25618,N_24105,N_24630);
and U25619 (N_25619,N_24176,N_24089);
nor U25620 (N_25620,N_24719,N_24092);
xor U25621 (N_25621,N_24346,N_24278);
and U25622 (N_25622,N_24039,N_24745);
nor U25623 (N_25623,N_24692,N_24951);
xnor U25624 (N_25624,N_24224,N_24530);
xnor U25625 (N_25625,N_24996,N_24084);
or U25626 (N_25626,N_24976,N_24469);
xnor U25627 (N_25627,N_24893,N_24934);
and U25628 (N_25628,N_24136,N_24031);
xor U25629 (N_25629,N_24881,N_24585);
xor U25630 (N_25630,N_24943,N_24846);
xnor U25631 (N_25631,N_24984,N_24686);
and U25632 (N_25632,N_24507,N_24887);
and U25633 (N_25633,N_24577,N_24439);
or U25634 (N_25634,N_24921,N_24004);
xor U25635 (N_25635,N_24775,N_24053);
or U25636 (N_25636,N_24351,N_24935);
xnor U25637 (N_25637,N_24491,N_24622);
or U25638 (N_25638,N_24523,N_24166);
nor U25639 (N_25639,N_24950,N_24585);
and U25640 (N_25640,N_24059,N_24390);
nor U25641 (N_25641,N_24956,N_24450);
nand U25642 (N_25642,N_24865,N_24078);
xor U25643 (N_25643,N_24766,N_24564);
and U25644 (N_25644,N_24732,N_24026);
nand U25645 (N_25645,N_24931,N_24411);
nor U25646 (N_25646,N_24601,N_24269);
xnor U25647 (N_25647,N_24048,N_24848);
or U25648 (N_25648,N_24304,N_24616);
nor U25649 (N_25649,N_24316,N_24917);
nor U25650 (N_25650,N_24122,N_24538);
and U25651 (N_25651,N_24166,N_24634);
and U25652 (N_25652,N_24507,N_24526);
or U25653 (N_25653,N_24503,N_24968);
or U25654 (N_25654,N_24059,N_24796);
and U25655 (N_25655,N_24534,N_24879);
and U25656 (N_25656,N_24647,N_24889);
nor U25657 (N_25657,N_24110,N_24170);
nor U25658 (N_25658,N_24412,N_24864);
nor U25659 (N_25659,N_24294,N_24917);
and U25660 (N_25660,N_24182,N_24639);
or U25661 (N_25661,N_24232,N_24678);
xor U25662 (N_25662,N_24570,N_24178);
xor U25663 (N_25663,N_24285,N_24579);
nand U25664 (N_25664,N_24418,N_24403);
xnor U25665 (N_25665,N_24684,N_24128);
xnor U25666 (N_25666,N_24536,N_24474);
nand U25667 (N_25667,N_24310,N_24594);
xnor U25668 (N_25668,N_24436,N_24429);
and U25669 (N_25669,N_24878,N_24033);
nand U25670 (N_25670,N_24709,N_24683);
or U25671 (N_25671,N_24516,N_24156);
or U25672 (N_25672,N_24011,N_24506);
nand U25673 (N_25673,N_24541,N_24457);
nand U25674 (N_25674,N_24662,N_24913);
or U25675 (N_25675,N_24068,N_24975);
nor U25676 (N_25676,N_24627,N_24964);
nand U25677 (N_25677,N_24898,N_24979);
or U25678 (N_25678,N_24441,N_24361);
nor U25679 (N_25679,N_24399,N_24129);
nand U25680 (N_25680,N_24303,N_24021);
xor U25681 (N_25681,N_24863,N_24363);
or U25682 (N_25682,N_24597,N_24586);
xor U25683 (N_25683,N_24378,N_24481);
or U25684 (N_25684,N_24287,N_24255);
nor U25685 (N_25685,N_24697,N_24467);
nor U25686 (N_25686,N_24294,N_24758);
and U25687 (N_25687,N_24513,N_24358);
nand U25688 (N_25688,N_24026,N_24443);
nand U25689 (N_25689,N_24714,N_24804);
and U25690 (N_25690,N_24811,N_24408);
nand U25691 (N_25691,N_24496,N_24944);
xnor U25692 (N_25692,N_24507,N_24150);
and U25693 (N_25693,N_24394,N_24519);
nor U25694 (N_25694,N_24497,N_24699);
nor U25695 (N_25695,N_24768,N_24312);
and U25696 (N_25696,N_24246,N_24471);
and U25697 (N_25697,N_24292,N_24239);
nor U25698 (N_25698,N_24444,N_24926);
xnor U25699 (N_25699,N_24109,N_24497);
nor U25700 (N_25700,N_24911,N_24893);
nand U25701 (N_25701,N_24285,N_24687);
or U25702 (N_25702,N_24992,N_24735);
and U25703 (N_25703,N_24052,N_24583);
or U25704 (N_25704,N_24036,N_24465);
or U25705 (N_25705,N_24321,N_24028);
nand U25706 (N_25706,N_24454,N_24947);
nand U25707 (N_25707,N_24583,N_24644);
and U25708 (N_25708,N_24951,N_24408);
or U25709 (N_25709,N_24619,N_24250);
and U25710 (N_25710,N_24528,N_24550);
xnor U25711 (N_25711,N_24512,N_24163);
xnor U25712 (N_25712,N_24374,N_24654);
xnor U25713 (N_25713,N_24448,N_24050);
xor U25714 (N_25714,N_24208,N_24253);
or U25715 (N_25715,N_24483,N_24531);
xor U25716 (N_25716,N_24514,N_24456);
nor U25717 (N_25717,N_24746,N_24183);
or U25718 (N_25718,N_24027,N_24566);
nand U25719 (N_25719,N_24827,N_24669);
xor U25720 (N_25720,N_24276,N_24294);
and U25721 (N_25721,N_24865,N_24145);
nor U25722 (N_25722,N_24750,N_24985);
xnor U25723 (N_25723,N_24259,N_24587);
and U25724 (N_25724,N_24838,N_24633);
and U25725 (N_25725,N_24806,N_24603);
and U25726 (N_25726,N_24411,N_24678);
xor U25727 (N_25727,N_24318,N_24747);
nor U25728 (N_25728,N_24262,N_24764);
and U25729 (N_25729,N_24039,N_24432);
nor U25730 (N_25730,N_24875,N_24167);
nor U25731 (N_25731,N_24569,N_24068);
nor U25732 (N_25732,N_24723,N_24143);
nand U25733 (N_25733,N_24984,N_24090);
or U25734 (N_25734,N_24108,N_24838);
and U25735 (N_25735,N_24431,N_24441);
nor U25736 (N_25736,N_24236,N_24048);
nor U25737 (N_25737,N_24563,N_24669);
xnor U25738 (N_25738,N_24519,N_24307);
or U25739 (N_25739,N_24574,N_24146);
or U25740 (N_25740,N_24081,N_24196);
or U25741 (N_25741,N_24863,N_24427);
and U25742 (N_25742,N_24725,N_24912);
nand U25743 (N_25743,N_24271,N_24808);
or U25744 (N_25744,N_24719,N_24099);
nor U25745 (N_25745,N_24328,N_24567);
nand U25746 (N_25746,N_24818,N_24645);
xor U25747 (N_25747,N_24722,N_24076);
and U25748 (N_25748,N_24077,N_24804);
and U25749 (N_25749,N_24571,N_24069);
and U25750 (N_25750,N_24161,N_24514);
nor U25751 (N_25751,N_24598,N_24563);
nand U25752 (N_25752,N_24722,N_24632);
or U25753 (N_25753,N_24415,N_24178);
and U25754 (N_25754,N_24903,N_24421);
and U25755 (N_25755,N_24621,N_24991);
or U25756 (N_25756,N_24556,N_24911);
or U25757 (N_25757,N_24256,N_24241);
xor U25758 (N_25758,N_24152,N_24782);
xor U25759 (N_25759,N_24710,N_24771);
nor U25760 (N_25760,N_24532,N_24267);
or U25761 (N_25761,N_24001,N_24137);
nand U25762 (N_25762,N_24897,N_24710);
nand U25763 (N_25763,N_24888,N_24147);
xnor U25764 (N_25764,N_24413,N_24553);
and U25765 (N_25765,N_24417,N_24246);
xnor U25766 (N_25766,N_24111,N_24037);
or U25767 (N_25767,N_24695,N_24486);
and U25768 (N_25768,N_24872,N_24942);
or U25769 (N_25769,N_24417,N_24613);
or U25770 (N_25770,N_24398,N_24749);
xor U25771 (N_25771,N_24831,N_24025);
nand U25772 (N_25772,N_24200,N_24792);
or U25773 (N_25773,N_24265,N_24139);
nand U25774 (N_25774,N_24970,N_24060);
or U25775 (N_25775,N_24149,N_24983);
and U25776 (N_25776,N_24446,N_24018);
nand U25777 (N_25777,N_24459,N_24942);
or U25778 (N_25778,N_24124,N_24380);
or U25779 (N_25779,N_24713,N_24152);
nand U25780 (N_25780,N_24139,N_24658);
nand U25781 (N_25781,N_24659,N_24195);
nor U25782 (N_25782,N_24039,N_24459);
nand U25783 (N_25783,N_24007,N_24396);
xor U25784 (N_25784,N_24525,N_24474);
and U25785 (N_25785,N_24834,N_24082);
nand U25786 (N_25786,N_24334,N_24777);
xor U25787 (N_25787,N_24774,N_24197);
or U25788 (N_25788,N_24353,N_24786);
or U25789 (N_25789,N_24169,N_24039);
xor U25790 (N_25790,N_24709,N_24431);
and U25791 (N_25791,N_24456,N_24616);
nand U25792 (N_25792,N_24046,N_24970);
xnor U25793 (N_25793,N_24711,N_24654);
xnor U25794 (N_25794,N_24804,N_24770);
xor U25795 (N_25795,N_24584,N_24516);
xor U25796 (N_25796,N_24027,N_24432);
and U25797 (N_25797,N_24297,N_24620);
nor U25798 (N_25798,N_24624,N_24362);
and U25799 (N_25799,N_24820,N_24175);
nand U25800 (N_25800,N_24654,N_24398);
or U25801 (N_25801,N_24699,N_24361);
nor U25802 (N_25802,N_24809,N_24250);
xnor U25803 (N_25803,N_24392,N_24380);
nand U25804 (N_25804,N_24182,N_24216);
xnor U25805 (N_25805,N_24675,N_24730);
and U25806 (N_25806,N_24913,N_24148);
xor U25807 (N_25807,N_24867,N_24983);
xnor U25808 (N_25808,N_24071,N_24905);
nor U25809 (N_25809,N_24779,N_24573);
nand U25810 (N_25810,N_24463,N_24290);
nand U25811 (N_25811,N_24396,N_24721);
or U25812 (N_25812,N_24943,N_24502);
or U25813 (N_25813,N_24260,N_24805);
and U25814 (N_25814,N_24583,N_24959);
or U25815 (N_25815,N_24042,N_24105);
and U25816 (N_25816,N_24745,N_24716);
and U25817 (N_25817,N_24956,N_24785);
nand U25818 (N_25818,N_24011,N_24915);
and U25819 (N_25819,N_24359,N_24692);
and U25820 (N_25820,N_24384,N_24275);
xor U25821 (N_25821,N_24006,N_24626);
or U25822 (N_25822,N_24905,N_24621);
xor U25823 (N_25823,N_24320,N_24605);
and U25824 (N_25824,N_24121,N_24663);
and U25825 (N_25825,N_24103,N_24311);
or U25826 (N_25826,N_24052,N_24977);
xnor U25827 (N_25827,N_24784,N_24476);
nor U25828 (N_25828,N_24797,N_24555);
or U25829 (N_25829,N_24711,N_24513);
and U25830 (N_25830,N_24925,N_24656);
nand U25831 (N_25831,N_24280,N_24129);
or U25832 (N_25832,N_24123,N_24186);
nor U25833 (N_25833,N_24486,N_24560);
nor U25834 (N_25834,N_24569,N_24027);
nand U25835 (N_25835,N_24103,N_24273);
nor U25836 (N_25836,N_24157,N_24425);
or U25837 (N_25837,N_24193,N_24351);
nand U25838 (N_25838,N_24795,N_24947);
xor U25839 (N_25839,N_24420,N_24807);
nor U25840 (N_25840,N_24358,N_24663);
and U25841 (N_25841,N_24421,N_24334);
and U25842 (N_25842,N_24190,N_24624);
xor U25843 (N_25843,N_24695,N_24456);
nor U25844 (N_25844,N_24243,N_24757);
nor U25845 (N_25845,N_24547,N_24795);
or U25846 (N_25846,N_24299,N_24629);
nand U25847 (N_25847,N_24970,N_24007);
nor U25848 (N_25848,N_24412,N_24529);
or U25849 (N_25849,N_24245,N_24148);
nand U25850 (N_25850,N_24651,N_24167);
nor U25851 (N_25851,N_24936,N_24032);
xnor U25852 (N_25852,N_24055,N_24050);
nand U25853 (N_25853,N_24980,N_24680);
nand U25854 (N_25854,N_24017,N_24167);
and U25855 (N_25855,N_24762,N_24577);
nor U25856 (N_25856,N_24624,N_24205);
and U25857 (N_25857,N_24904,N_24514);
nor U25858 (N_25858,N_24074,N_24001);
or U25859 (N_25859,N_24918,N_24604);
nand U25860 (N_25860,N_24238,N_24365);
nor U25861 (N_25861,N_24558,N_24182);
or U25862 (N_25862,N_24312,N_24986);
nand U25863 (N_25863,N_24434,N_24634);
xnor U25864 (N_25864,N_24382,N_24907);
xor U25865 (N_25865,N_24542,N_24271);
xor U25866 (N_25866,N_24164,N_24782);
and U25867 (N_25867,N_24349,N_24864);
nor U25868 (N_25868,N_24439,N_24872);
xor U25869 (N_25869,N_24083,N_24124);
and U25870 (N_25870,N_24564,N_24324);
xnor U25871 (N_25871,N_24867,N_24863);
or U25872 (N_25872,N_24291,N_24990);
and U25873 (N_25873,N_24133,N_24979);
and U25874 (N_25874,N_24974,N_24126);
and U25875 (N_25875,N_24760,N_24335);
nor U25876 (N_25876,N_24637,N_24214);
nor U25877 (N_25877,N_24204,N_24005);
or U25878 (N_25878,N_24471,N_24146);
or U25879 (N_25879,N_24510,N_24191);
or U25880 (N_25880,N_24302,N_24043);
xor U25881 (N_25881,N_24419,N_24720);
or U25882 (N_25882,N_24118,N_24971);
nand U25883 (N_25883,N_24128,N_24380);
nor U25884 (N_25884,N_24832,N_24039);
xor U25885 (N_25885,N_24594,N_24073);
xor U25886 (N_25886,N_24992,N_24917);
nor U25887 (N_25887,N_24840,N_24140);
or U25888 (N_25888,N_24943,N_24080);
or U25889 (N_25889,N_24801,N_24117);
or U25890 (N_25890,N_24564,N_24997);
nand U25891 (N_25891,N_24750,N_24902);
nand U25892 (N_25892,N_24415,N_24980);
or U25893 (N_25893,N_24433,N_24683);
nor U25894 (N_25894,N_24324,N_24913);
nor U25895 (N_25895,N_24181,N_24583);
or U25896 (N_25896,N_24037,N_24989);
xor U25897 (N_25897,N_24835,N_24825);
or U25898 (N_25898,N_24605,N_24431);
and U25899 (N_25899,N_24772,N_24219);
nor U25900 (N_25900,N_24040,N_24185);
nand U25901 (N_25901,N_24011,N_24526);
xnor U25902 (N_25902,N_24457,N_24051);
or U25903 (N_25903,N_24545,N_24632);
or U25904 (N_25904,N_24027,N_24831);
and U25905 (N_25905,N_24867,N_24779);
nor U25906 (N_25906,N_24708,N_24373);
xor U25907 (N_25907,N_24475,N_24682);
nor U25908 (N_25908,N_24593,N_24188);
nor U25909 (N_25909,N_24289,N_24039);
xor U25910 (N_25910,N_24893,N_24928);
and U25911 (N_25911,N_24697,N_24791);
or U25912 (N_25912,N_24921,N_24453);
xnor U25913 (N_25913,N_24418,N_24757);
nand U25914 (N_25914,N_24387,N_24902);
nand U25915 (N_25915,N_24098,N_24326);
xnor U25916 (N_25916,N_24924,N_24082);
nor U25917 (N_25917,N_24899,N_24303);
nor U25918 (N_25918,N_24367,N_24646);
and U25919 (N_25919,N_24803,N_24427);
nand U25920 (N_25920,N_24240,N_24407);
and U25921 (N_25921,N_24586,N_24968);
and U25922 (N_25922,N_24655,N_24448);
nor U25923 (N_25923,N_24867,N_24521);
nand U25924 (N_25924,N_24657,N_24385);
nand U25925 (N_25925,N_24285,N_24861);
nand U25926 (N_25926,N_24774,N_24778);
nand U25927 (N_25927,N_24885,N_24134);
xnor U25928 (N_25928,N_24829,N_24893);
nor U25929 (N_25929,N_24017,N_24385);
or U25930 (N_25930,N_24818,N_24542);
and U25931 (N_25931,N_24930,N_24633);
nor U25932 (N_25932,N_24691,N_24173);
and U25933 (N_25933,N_24350,N_24499);
nand U25934 (N_25934,N_24391,N_24328);
and U25935 (N_25935,N_24132,N_24937);
and U25936 (N_25936,N_24476,N_24790);
or U25937 (N_25937,N_24122,N_24578);
or U25938 (N_25938,N_24064,N_24497);
or U25939 (N_25939,N_24587,N_24683);
nor U25940 (N_25940,N_24090,N_24435);
and U25941 (N_25941,N_24538,N_24900);
xor U25942 (N_25942,N_24064,N_24442);
or U25943 (N_25943,N_24079,N_24538);
nor U25944 (N_25944,N_24264,N_24122);
nand U25945 (N_25945,N_24219,N_24574);
nand U25946 (N_25946,N_24913,N_24503);
xor U25947 (N_25947,N_24424,N_24533);
xnor U25948 (N_25948,N_24037,N_24182);
and U25949 (N_25949,N_24512,N_24188);
nor U25950 (N_25950,N_24985,N_24484);
nand U25951 (N_25951,N_24728,N_24151);
nor U25952 (N_25952,N_24971,N_24080);
nor U25953 (N_25953,N_24998,N_24910);
nor U25954 (N_25954,N_24311,N_24953);
or U25955 (N_25955,N_24384,N_24994);
xnor U25956 (N_25956,N_24080,N_24136);
nand U25957 (N_25957,N_24010,N_24915);
xor U25958 (N_25958,N_24058,N_24852);
or U25959 (N_25959,N_24967,N_24030);
nand U25960 (N_25960,N_24691,N_24708);
nor U25961 (N_25961,N_24685,N_24901);
and U25962 (N_25962,N_24699,N_24029);
or U25963 (N_25963,N_24145,N_24803);
and U25964 (N_25964,N_24527,N_24248);
or U25965 (N_25965,N_24126,N_24896);
or U25966 (N_25966,N_24588,N_24748);
or U25967 (N_25967,N_24745,N_24437);
nor U25968 (N_25968,N_24024,N_24450);
and U25969 (N_25969,N_24958,N_24823);
nor U25970 (N_25970,N_24736,N_24052);
xnor U25971 (N_25971,N_24357,N_24314);
and U25972 (N_25972,N_24382,N_24349);
xnor U25973 (N_25973,N_24142,N_24967);
and U25974 (N_25974,N_24051,N_24886);
or U25975 (N_25975,N_24572,N_24393);
xnor U25976 (N_25976,N_24141,N_24527);
nand U25977 (N_25977,N_24446,N_24187);
xor U25978 (N_25978,N_24752,N_24846);
nor U25979 (N_25979,N_24385,N_24760);
and U25980 (N_25980,N_24047,N_24559);
nor U25981 (N_25981,N_24583,N_24992);
and U25982 (N_25982,N_24931,N_24218);
and U25983 (N_25983,N_24492,N_24498);
nor U25984 (N_25984,N_24125,N_24496);
and U25985 (N_25985,N_24455,N_24936);
or U25986 (N_25986,N_24247,N_24216);
nor U25987 (N_25987,N_24845,N_24482);
nor U25988 (N_25988,N_24746,N_24987);
or U25989 (N_25989,N_24349,N_24007);
or U25990 (N_25990,N_24622,N_24147);
nor U25991 (N_25991,N_24835,N_24714);
xor U25992 (N_25992,N_24527,N_24005);
or U25993 (N_25993,N_24562,N_24278);
nand U25994 (N_25994,N_24471,N_24791);
and U25995 (N_25995,N_24631,N_24973);
xor U25996 (N_25996,N_24066,N_24912);
xor U25997 (N_25997,N_24806,N_24117);
xor U25998 (N_25998,N_24766,N_24672);
or U25999 (N_25999,N_24770,N_24189);
nor U26000 (N_26000,N_25724,N_25874);
nor U26001 (N_26001,N_25095,N_25030);
xor U26002 (N_26002,N_25422,N_25259);
nand U26003 (N_26003,N_25691,N_25521);
and U26004 (N_26004,N_25170,N_25167);
or U26005 (N_26005,N_25336,N_25296);
xnor U26006 (N_26006,N_25859,N_25300);
nor U26007 (N_26007,N_25380,N_25599);
and U26008 (N_26008,N_25585,N_25538);
and U26009 (N_26009,N_25733,N_25184);
and U26010 (N_26010,N_25061,N_25718);
nor U26011 (N_26011,N_25710,N_25877);
nand U26012 (N_26012,N_25965,N_25734);
xnor U26013 (N_26013,N_25835,N_25530);
and U26014 (N_26014,N_25009,N_25889);
and U26015 (N_26015,N_25754,N_25858);
and U26016 (N_26016,N_25892,N_25515);
or U26017 (N_26017,N_25563,N_25635);
nand U26018 (N_26018,N_25345,N_25326);
and U26019 (N_26019,N_25478,N_25152);
nor U26020 (N_26020,N_25216,N_25493);
or U26021 (N_26021,N_25987,N_25607);
nor U26022 (N_26022,N_25140,N_25284);
nand U26023 (N_26023,N_25533,N_25525);
nor U26024 (N_26024,N_25143,N_25731);
xor U26025 (N_26025,N_25065,N_25670);
xor U26026 (N_26026,N_25562,N_25435);
or U26027 (N_26027,N_25011,N_25904);
nand U26028 (N_26028,N_25667,N_25163);
or U26029 (N_26029,N_25505,N_25319);
and U26030 (N_26030,N_25348,N_25648);
nand U26031 (N_26031,N_25194,N_25437);
or U26032 (N_26032,N_25334,N_25841);
xor U26033 (N_26033,N_25104,N_25765);
xor U26034 (N_26034,N_25328,N_25499);
nand U26035 (N_26035,N_25470,N_25487);
xor U26036 (N_26036,N_25134,N_25202);
or U26037 (N_26037,N_25130,N_25898);
nand U26038 (N_26038,N_25294,N_25662);
xnor U26039 (N_26039,N_25679,N_25112);
and U26040 (N_26040,N_25629,N_25798);
xor U26041 (N_26041,N_25050,N_25091);
nor U26042 (N_26042,N_25744,N_25467);
xnor U26043 (N_26043,N_25206,N_25366);
nor U26044 (N_26044,N_25368,N_25213);
nand U26045 (N_26045,N_25456,N_25769);
or U26046 (N_26046,N_25389,N_25409);
nand U26047 (N_26047,N_25753,N_25094);
nand U26048 (N_26048,N_25469,N_25702);
xnor U26049 (N_26049,N_25388,N_25245);
and U26050 (N_26050,N_25557,N_25018);
xnor U26051 (N_26051,N_25875,N_25711);
nor U26052 (N_26052,N_25866,N_25196);
or U26053 (N_26053,N_25846,N_25806);
or U26054 (N_26054,N_25021,N_25773);
nand U26055 (N_26055,N_25375,N_25592);
and U26056 (N_26056,N_25414,N_25998);
xor U26057 (N_26057,N_25964,N_25688);
and U26058 (N_26058,N_25325,N_25291);
and U26059 (N_26059,N_25192,N_25709);
and U26060 (N_26060,N_25158,N_25567);
and U26061 (N_26061,N_25074,N_25545);
nand U26062 (N_26062,N_25920,N_25070);
nor U26063 (N_26063,N_25132,N_25238);
nand U26064 (N_26064,N_25102,N_25115);
and U26065 (N_26065,N_25003,N_25539);
or U26066 (N_26066,N_25771,N_25799);
and U26067 (N_26067,N_25796,N_25522);
and U26068 (N_26068,N_25742,N_25556);
nor U26069 (N_26069,N_25031,N_25048);
nor U26070 (N_26070,N_25634,N_25869);
nor U26071 (N_26071,N_25621,N_25982);
and U26072 (N_26072,N_25717,N_25929);
xor U26073 (N_26073,N_25298,N_25615);
xor U26074 (N_26074,N_25647,N_25075);
nor U26075 (N_26075,N_25708,N_25304);
nand U26076 (N_26076,N_25190,N_25921);
nand U26077 (N_26077,N_25623,N_25950);
nor U26078 (N_26078,N_25772,N_25138);
nor U26079 (N_26079,N_25884,N_25800);
and U26080 (N_26080,N_25079,N_25549);
or U26081 (N_26081,N_25820,N_25098);
or U26082 (N_26082,N_25992,N_25241);
or U26083 (N_26083,N_25459,N_25767);
nor U26084 (N_26084,N_25077,N_25504);
and U26085 (N_26085,N_25093,N_25593);
nor U26086 (N_26086,N_25637,N_25330);
nor U26087 (N_26087,N_25084,N_25523);
nand U26088 (N_26088,N_25855,N_25028);
xnor U26089 (N_26089,N_25736,N_25879);
nor U26090 (N_26090,N_25208,N_25945);
or U26091 (N_26091,N_25489,N_25661);
or U26092 (N_26092,N_25517,N_25922);
nor U26093 (N_26093,N_25377,N_25531);
or U26094 (N_26094,N_25264,N_25816);
xor U26095 (N_26095,N_25417,N_25177);
nor U26096 (N_26096,N_25566,N_25344);
and U26097 (N_26097,N_25963,N_25935);
and U26098 (N_26098,N_25195,N_25280);
nor U26099 (N_26099,N_25595,N_25324);
xor U26100 (N_26100,N_25838,N_25949);
xnor U26101 (N_26101,N_25401,N_25979);
nor U26102 (N_26102,N_25385,N_25418);
xnor U26103 (N_26103,N_25883,N_25760);
or U26104 (N_26104,N_25870,N_25354);
nor U26105 (N_26105,N_25958,N_25750);
or U26106 (N_26106,N_25681,N_25761);
nor U26107 (N_26107,N_25780,N_25911);
nand U26108 (N_26108,N_25970,N_25316);
nor U26109 (N_26109,N_25865,N_25698);
xnor U26110 (N_26110,N_25671,N_25775);
xor U26111 (N_26111,N_25453,N_25236);
and U26112 (N_26112,N_25747,N_25495);
nand U26113 (N_26113,N_25980,N_25864);
and U26114 (N_26114,N_25237,N_25179);
nor U26115 (N_26115,N_25613,N_25416);
or U26116 (N_26116,N_25056,N_25932);
or U26117 (N_26117,N_25830,N_25117);
nor U26118 (N_26118,N_25103,N_25540);
and U26119 (N_26119,N_25854,N_25477);
nand U26120 (N_26120,N_25069,N_25390);
xor U26121 (N_26121,N_25451,N_25692);
xor U26122 (N_26122,N_25146,N_25063);
nor U26123 (N_26123,N_25087,N_25497);
and U26124 (N_26124,N_25106,N_25827);
xor U26125 (N_26125,N_25359,N_25730);
and U26126 (N_26126,N_25008,N_25329);
nor U26127 (N_26127,N_25720,N_25412);
or U26128 (N_26128,N_25758,N_25831);
nand U26129 (N_26129,N_25252,N_25608);
nand U26130 (N_26130,N_25673,N_25349);
and U26131 (N_26131,N_25514,N_25555);
nor U26132 (N_26132,N_25356,N_25966);
and U26133 (N_26133,N_25430,N_25253);
nor U26134 (N_26134,N_25161,N_25936);
and U26135 (N_26135,N_25790,N_25047);
nand U26136 (N_26136,N_25728,N_25628);
or U26137 (N_26137,N_25974,N_25223);
or U26138 (N_26138,N_25981,N_25491);
nor U26139 (N_26139,N_25054,N_25032);
or U26140 (N_26140,N_25492,N_25352);
and U26141 (N_26141,N_25783,N_25488);
or U26142 (N_26142,N_25732,N_25686);
nand U26143 (N_26143,N_25513,N_25664);
nand U26144 (N_26144,N_25258,N_25971);
nor U26145 (N_26145,N_25066,N_25942);
xnor U26146 (N_26146,N_25441,N_25128);
nand U26147 (N_26147,N_25885,N_25895);
nand U26148 (N_26148,N_25727,N_25270);
and U26149 (N_26149,N_25712,N_25089);
nor U26150 (N_26150,N_25458,N_25049);
or U26151 (N_26151,N_25397,N_25410);
nand U26152 (N_26152,N_25343,N_25872);
nand U26153 (N_26153,N_25244,N_25861);
nor U26154 (N_26154,N_25697,N_25466);
nor U26155 (N_26155,N_25645,N_25649);
and U26156 (N_26156,N_25439,N_25153);
xnor U26157 (N_26157,N_25240,N_25174);
and U26158 (N_26158,N_25494,N_25528);
nor U26159 (N_26159,N_25255,N_25078);
nor U26160 (N_26160,N_25626,N_25577);
and U26161 (N_26161,N_25405,N_25293);
nand U26162 (N_26162,N_25185,N_25023);
nor U26163 (N_26163,N_25215,N_25756);
and U26164 (N_26164,N_25341,N_25485);
xor U26165 (N_26165,N_25684,N_25526);
nor U26166 (N_26166,N_25694,N_25496);
nand U26167 (N_26167,N_25845,N_25057);
xnor U26168 (N_26168,N_25081,N_25852);
nand U26169 (N_26169,N_25612,N_25794);
and U26170 (N_26170,N_25660,N_25480);
xor U26171 (N_26171,N_25440,N_25689);
and U26172 (N_26172,N_25310,N_25071);
nand U26173 (N_26173,N_25891,N_25604);
or U26174 (N_26174,N_25373,N_25224);
nand U26175 (N_26175,N_25781,N_25658);
xnor U26176 (N_26176,N_25524,N_25640);
or U26177 (N_26177,N_25239,N_25824);
and U26178 (N_26178,N_25187,N_25007);
and U26179 (N_26179,N_25803,N_25901);
or U26180 (N_26180,N_25541,N_25961);
nor U26181 (N_26181,N_25229,N_25120);
and U26182 (N_26182,N_25165,N_25465);
xor U26183 (N_26183,N_25766,N_25666);
nand U26184 (N_26184,N_25299,N_25535);
nor U26185 (N_26185,N_25676,N_25108);
nand U26186 (N_26186,N_25878,N_25933);
or U26187 (N_26187,N_25848,N_25403);
and U26188 (N_26188,N_25124,N_25737);
xnor U26189 (N_26189,N_25818,N_25999);
nor U26190 (N_26190,N_25231,N_25996);
nor U26191 (N_26191,N_25729,N_25272);
and U26192 (N_26192,N_25100,N_25320);
and U26193 (N_26193,N_25129,N_25481);
nor U26194 (N_26194,N_25941,N_25110);
xor U26195 (N_26195,N_25082,N_25819);
xnor U26196 (N_26196,N_25012,N_25886);
nand U26197 (N_26197,N_25695,N_25572);
xnor U26198 (N_26198,N_25991,N_25644);
nand U26199 (N_26199,N_25683,N_25425);
nand U26200 (N_26200,N_25203,N_25150);
nor U26201 (N_26201,N_25723,N_25111);
and U26202 (N_26202,N_25839,N_25751);
or U26203 (N_26203,N_25035,N_25601);
or U26204 (N_26204,N_25943,N_25828);
or U26205 (N_26205,N_25279,N_25764);
and U26206 (N_26206,N_25887,N_25972);
and U26207 (N_26207,N_25387,N_25770);
xor U26208 (N_26208,N_25234,N_25903);
or U26209 (N_26209,N_25669,N_25520);
and U26210 (N_26210,N_25083,N_25639);
xnor U26211 (N_26211,N_25821,N_25990);
or U26212 (N_26212,N_25043,N_25583);
xnor U26213 (N_26213,N_25289,N_25871);
nor U26214 (N_26214,N_25940,N_25778);
xor U26215 (N_26215,N_25927,N_25307);
and U26216 (N_26216,N_25518,N_25757);
xnor U26217 (N_26217,N_25713,N_25804);
or U26218 (N_26218,N_25641,N_25169);
xor U26219 (N_26219,N_25141,N_25810);
and U26220 (N_26220,N_25292,N_25114);
or U26221 (N_26221,N_25479,N_25997);
nand U26222 (N_26222,N_25873,N_25896);
nor U26223 (N_26223,N_25396,N_25986);
or U26224 (N_26224,N_25832,N_25550);
nand U26225 (N_26225,N_25912,N_25598);
and U26226 (N_26226,N_25014,N_25516);
or U26227 (N_26227,N_25571,N_25579);
or U26228 (N_26228,N_25725,N_25947);
xor U26229 (N_26229,N_25755,N_25653);
or U26230 (N_26230,N_25789,N_25622);
or U26231 (N_26231,N_25249,N_25088);
nand U26232 (N_26232,N_25446,N_25250);
or U26233 (N_26233,N_25907,N_25149);
nand U26234 (N_26234,N_25954,N_25286);
xor U26235 (N_26235,N_25256,N_25536);
and U26236 (N_26236,N_25837,N_25529);
xnor U26237 (N_26237,N_25876,N_25045);
or U26238 (N_26238,N_25842,N_25145);
nand U26239 (N_26239,N_25118,N_25969);
xnor U26240 (N_26240,N_25263,N_25242);
or U26241 (N_26241,N_25133,N_25315);
nand U26242 (N_26242,N_25716,N_25897);
nor U26243 (N_26243,N_25421,N_25016);
and U26244 (N_26244,N_25144,N_25784);
xor U26245 (N_26245,N_25276,N_25415);
nand U26246 (N_26246,N_25445,N_25603);
or U26247 (N_26247,N_25680,N_25059);
nand U26248 (N_26248,N_25125,N_25218);
and U26249 (N_26249,N_25551,N_25693);
or U26250 (N_26250,N_25452,N_25109);
xor U26251 (N_26251,N_25973,N_25285);
nand U26252 (N_26252,N_25266,N_25925);
xor U26253 (N_26253,N_25856,N_25400);
or U26254 (N_26254,N_25714,N_25696);
or U26255 (N_26255,N_25092,N_25701);
and U26256 (N_26256,N_25312,N_25956);
or U26257 (N_26257,N_25323,N_25247);
nand U26258 (N_26258,N_25394,N_25155);
or U26259 (N_26259,N_25355,N_25271);
xor U26260 (N_26260,N_25162,N_25472);
nor U26261 (N_26261,N_25321,N_25937);
or U26262 (N_26262,N_25426,N_25166);
nor U26263 (N_26263,N_25086,N_25748);
nand U26264 (N_26264,N_25543,N_25833);
xnor U26265 (N_26265,N_25657,N_25025);
nor U26266 (N_26266,N_25034,N_25802);
or U26267 (N_26267,N_25220,N_25829);
xnor U26268 (N_26268,N_25914,N_25880);
nand U26269 (N_26269,N_25610,N_25857);
nand U26270 (N_26270,N_25137,N_25651);
nor U26271 (N_26271,N_25340,N_25962);
or U26272 (N_26272,N_25243,N_25339);
xnor U26273 (N_26273,N_25602,N_25046);
nand U26274 (N_26274,N_25282,N_25423);
xnor U26275 (N_26275,N_25314,N_25519);
or U26276 (N_26276,N_25331,N_25559);
and U26277 (N_26277,N_25073,N_25309);
and U26278 (N_26278,N_25532,N_25361);
and U26279 (N_26279,N_25262,N_25791);
nand U26280 (N_26280,N_25995,N_25844);
nor U26281 (N_26281,N_25906,N_25159);
nand U26282 (N_26282,N_25917,N_25589);
nand U26283 (N_26283,N_25370,N_25863);
nor U26284 (N_26284,N_25044,N_25588);
nand U26285 (N_26285,N_25656,N_25506);
and U26286 (N_26286,N_25722,N_25448);
xnor U26287 (N_26287,N_25851,N_25631);
nand U26288 (N_26288,N_25450,N_25338);
xnor U26289 (N_26289,N_25042,N_25500);
or U26290 (N_26290,N_25745,N_25616);
xor U26291 (N_26291,N_25399,N_25189);
xnor U26292 (N_26292,N_25611,N_25706);
nor U26293 (N_26293,N_25147,N_25617);
and U26294 (N_26294,N_25668,N_25391);
and U26295 (N_26295,N_25502,N_25449);
xnor U26296 (N_26296,N_25212,N_25490);
or U26297 (N_26297,N_25899,N_25978);
xor U26298 (N_26298,N_25575,N_25834);
or U26299 (N_26299,N_25303,N_25076);
nor U26300 (N_26300,N_25953,N_25010);
nand U26301 (N_26301,N_25739,N_25232);
and U26302 (N_26302,N_25297,N_25759);
nor U26303 (N_26303,N_25173,N_25672);
or U26304 (N_26304,N_25454,N_25197);
and U26305 (N_26305,N_25547,N_25560);
or U26306 (N_26306,N_25570,N_25428);
or U26307 (N_26307,N_25113,N_25946);
nand U26308 (N_26308,N_25384,N_25378);
xnor U26309 (N_26309,N_25994,N_25290);
and U26310 (N_26310,N_25278,N_25952);
nand U26311 (N_26311,N_25743,N_25636);
nand U26312 (N_26312,N_25815,N_25357);
nor U26313 (N_26313,N_25893,N_25029);
and U26314 (N_26314,N_25882,N_25156);
nor U26315 (N_26315,N_25843,N_25580);
and U26316 (N_26316,N_25287,N_25116);
xnor U26317 (N_26317,N_25792,N_25552);
xor U26318 (N_26318,N_25386,N_25546);
nand U26319 (N_26319,N_25609,N_25948);
or U26320 (N_26320,N_25062,N_25383);
or U26321 (N_26321,N_25433,N_25230);
nor U26322 (N_26322,N_25568,N_25139);
nand U26323 (N_26323,N_25786,N_25442);
and U26324 (N_26324,N_25726,N_25652);
xor U26325 (N_26325,N_25191,N_25429);
and U26326 (N_26326,N_25040,N_25928);
or U26327 (N_26327,N_25126,N_25017);
xor U26328 (N_26328,N_25944,N_25248);
nand U26329 (N_26329,N_25890,N_25811);
xnor U26330 (N_26330,N_25814,N_25703);
xor U26331 (N_26331,N_25227,N_25763);
nor U26332 (N_26332,N_25705,N_25420);
xor U26333 (N_26333,N_25160,N_25350);
nor U26334 (N_26334,N_25317,N_25096);
nand U26335 (N_26335,N_25374,N_25569);
xor U26336 (N_26336,N_25026,N_25413);
and U26337 (N_26337,N_25951,N_25822);
xnor U26338 (N_26338,N_25038,N_25265);
and U26339 (N_26339,N_25938,N_25905);
and U26340 (N_26340,N_25406,N_25659);
and U26341 (N_26341,N_25346,N_25544);
nand U26342 (N_26342,N_25807,N_25372);
or U26343 (N_26343,N_25431,N_25826);
nand U26344 (N_26344,N_25351,N_25825);
or U26345 (N_26345,N_25584,N_25131);
xor U26346 (N_26346,N_25119,N_25989);
or U26347 (N_26347,N_25643,N_25360);
nor U26348 (N_26348,N_25172,N_25273);
xnor U26349 (N_26349,N_25793,N_25840);
xor U26350 (N_26350,N_25900,N_25204);
and U26351 (N_26351,N_25438,N_25715);
nor U26352 (N_26352,N_25700,N_25633);
nor U26353 (N_26353,N_25000,N_25561);
nor U26354 (N_26354,N_25738,N_25004);
nand U26355 (N_26355,N_25455,N_25655);
nand U26356 (N_26356,N_25198,N_25483);
nor U26357 (N_26357,N_25565,N_25746);
xnor U26358 (N_26358,N_25573,N_25457);
xor U26359 (N_26359,N_25207,N_25808);
xor U26360 (N_26360,N_25868,N_25288);
xnor U26361 (N_26361,N_25019,N_25306);
nand U26362 (N_26362,N_25685,N_25337);
nor U26363 (N_26363,N_25823,N_25085);
and U26364 (N_26364,N_25376,N_25122);
nand U26365 (N_26365,N_25395,N_25217);
nor U26366 (N_26366,N_25182,N_25148);
xor U26367 (N_26367,N_25301,N_25600);
nand U26368 (N_26368,N_25408,N_25614);
nor U26369 (N_26369,N_25578,N_25507);
xor U26370 (N_26370,N_25053,N_25022);
xor U26371 (N_26371,N_25762,N_25931);
nand U26372 (N_26372,N_25178,N_25365);
nor U26373 (N_26373,N_25548,N_25027);
nand U26374 (N_26374,N_25847,N_25960);
nor U26375 (N_26375,N_25327,N_25967);
nand U26376 (N_26376,N_25427,N_25353);
or U26377 (N_26377,N_25001,N_25606);
xor U26378 (N_26378,N_25369,N_25537);
xnor U26379 (N_26379,N_25055,N_25630);
nand U26380 (N_26380,N_25785,N_25176);
xnor U26381 (N_26381,N_25930,N_25926);
and U26382 (N_26382,N_25015,N_25473);
nand U26383 (N_26383,N_25175,N_25432);
nand U26384 (N_26384,N_25939,N_25068);
or U26385 (N_26385,N_25419,N_25582);
or U26386 (N_26386,N_25006,N_25959);
xor U26387 (N_26387,N_25381,N_25955);
xnor U26388 (N_26388,N_25690,N_25041);
xor U26389 (N_26389,N_25512,N_25654);
xor U26390 (N_26390,N_25157,N_25460);
nor U26391 (N_26391,N_25210,N_25181);
or U26392 (N_26392,N_25051,N_25581);
nor U26393 (N_26393,N_25260,N_25476);
nor U26394 (N_26394,N_25154,N_25254);
or U26395 (N_26395,N_25919,N_25168);
or U26396 (N_26396,N_25067,N_25558);
or U26397 (N_26397,N_25699,N_25020);
xnor U26398 (N_26398,N_25809,N_25058);
or U26399 (N_26399,N_25463,N_25977);
or U26400 (N_26400,N_25127,N_25881);
xor U26401 (N_26401,N_25576,N_25090);
nor U26402 (N_26402,N_25261,N_25107);
xor U26403 (N_26403,N_25302,N_25382);
xor U26404 (N_26404,N_25591,N_25362);
nor U26405 (N_26405,N_25779,N_25590);
xnor U26406 (N_26406,N_25342,N_25674);
nor U26407 (N_26407,N_25618,N_25164);
xnor U26408 (N_26408,N_25510,N_25976);
xor U26409 (N_26409,N_25788,N_25902);
and U26410 (N_26410,N_25404,N_25214);
nor U26411 (N_26411,N_25393,N_25975);
nand U26412 (N_26412,N_25632,N_25251);
nand U26413 (N_26413,N_25620,N_25246);
xor U26414 (N_26414,N_25867,N_25205);
or U26415 (N_26415,N_25013,N_25984);
nand U26416 (N_26416,N_25295,N_25910);
or U26417 (N_26417,N_25527,N_25121);
nand U26418 (N_26418,N_25484,N_25036);
and U26419 (N_26419,N_25188,N_25183);
and U26420 (N_26420,N_25675,N_25392);
and U26421 (N_26421,N_25924,N_25219);
nor U26422 (N_26422,N_25060,N_25735);
nor U26423 (N_26423,N_25915,N_25267);
and U26424 (N_26424,N_25988,N_25311);
or U26425 (N_26425,N_25574,N_25983);
nand U26426 (N_26426,N_25482,N_25151);
or U26427 (N_26427,N_25554,N_25471);
xor U26428 (N_26428,N_25918,N_25913);
nor U26429 (N_26429,N_25646,N_25687);
nor U26430 (N_26430,N_25707,N_25436);
xor U26431 (N_26431,N_25222,N_25850);
or U26432 (N_26432,N_25367,N_25663);
and U26433 (N_26433,N_25801,N_25752);
xnor U26434 (N_26434,N_25269,N_25358);
nand U26435 (N_26435,N_25627,N_25605);
xor U26436 (N_26436,N_25511,N_25171);
or U26437 (N_26437,N_25587,N_25677);
nor U26438 (N_26438,N_25281,N_25812);
nand U26439 (N_26439,N_25235,N_25642);
nor U26440 (N_26440,N_25625,N_25862);
or U26441 (N_26441,N_25749,N_25638);
or U26442 (N_26442,N_25849,N_25424);
xnor U26443 (N_26443,N_25553,N_25719);
and U26444 (N_26444,N_25072,N_25508);
nand U26445 (N_26445,N_25277,N_25624);
nor U26446 (N_26446,N_25444,N_25542);
xor U26447 (N_26447,N_25860,N_25135);
or U26448 (N_26448,N_25002,N_25201);
nor U26449 (N_26449,N_25468,N_25411);
nor U26450 (N_26450,N_25209,N_25274);
nand U26451 (N_26451,N_25193,N_25464);
nand U26452 (N_26452,N_25402,N_25039);
and U26453 (N_26453,N_25475,N_25462);
xor U26454 (N_26454,N_25318,N_25509);
and U26455 (N_26455,N_25136,N_25371);
xnor U26456 (N_26456,N_25909,N_25741);
or U26457 (N_26457,N_25123,N_25097);
xor U26458 (N_26458,N_25805,N_25665);
or U26459 (N_26459,N_25777,N_25787);
nand U26460 (N_26460,N_25443,N_25033);
nor U26461 (N_26461,N_25257,N_25461);
nor U26462 (N_26462,N_25682,N_25005);
or U26463 (N_26463,N_25968,N_25916);
nor U26464 (N_26464,N_25678,N_25853);
nand U26465 (N_26465,N_25597,N_25934);
and U26466 (N_26466,N_25534,N_25985);
nand U26467 (N_26467,N_25797,N_25721);
nor U26468 (N_26468,N_25619,N_25398);
nand U26469 (N_26469,N_25186,N_25305);
xor U26470 (N_26470,N_25498,N_25322);
nor U26471 (N_26471,N_25586,N_25776);
nor U26472 (N_26472,N_25379,N_25813);
nor U26473 (N_26473,N_25228,N_25283);
xor U26474 (N_26474,N_25596,N_25447);
nor U26475 (N_26475,N_25774,N_25768);
or U26476 (N_26476,N_25888,N_25313);
nand U26477 (N_26477,N_25740,N_25024);
nor U26478 (N_26478,N_25064,N_25795);
nand U26479 (N_26479,N_25364,N_25347);
xor U26480 (N_26480,N_25308,N_25434);
nor U26481 (N_26481,N_25052,N_25486);
and U26482 (N_26482,N_25037,N_25200);
nand U26483 (N_26483,N_25503,N_25105);
or U26484 (N_26484,N_25225,N_25817);
or U26485 (N_26485,N_25923,N_25101);
nand U26486 (N_26486,N_25908,N_25564);
nand U26487 (N_26487,N_25199,N_25957);
nand U26488 (N_26488,N_25704,N_25782);
or U26489 (N_26489,N_25332,N_25221);
xor U26490 (N_26490,N_25180,N_25211);
or U26491 (N_26491,N_25894,N_25333);
xnor U26492 (N_26492,N_25226,N_25142);
xor U26493 (N_26493,N_25501,N_25275);
or U26494 (N_26494,N_25099,N_25474);
xor U26495 (N_26495,N_25080,N_25650);
nand U26496 (N_26496,N_25268,N_25233);
or U26497 (N_26497,N_25335,N_25993);
or U26498 (N_26498,N_25407,N_25594);
nand U26499 (N_26499,N_25836,N_25363);
and U26500 (N_26500,N_25832,N_25245);
and U26501 (N_26501,N_25160,N_25413);
and U26502 (N_26502,N_25573,N_25782);
or U26503 (N_26503,N_25388,N_25675);
or U26504 (N_26504,N_25040,N_25937);
nand U26505 (N_26505,N_25809,N_25336);
nor U26506 (N_26506,N_25318,N_25582);
and U26507 (N_26507,N_25969,N_25270);
nand U26508 (N_26508,N_25319,N_25327);
or U26509 (N_26509,N_25409,N_25847);
xor U26510 (N_26510,N_25539,N_25367);
nor U26511 (N_26511,N_25239,N_25676);
nor U26512 (N_26512,N_25100,N_25744);
or U26513 (N_26513,N_25649,N_25979);
and U26514 (N_26514,N_25066,N_25101);
xnor U26515 (N_26515,N_25296,N_25643);
nand U26516 (N_26516,N_25630,N_25809);
or U26517 (N_26517,N_25097,N_25502);
and U26518 (N_26518,N_25762,N_25753);
nand U26519 (N_26519,N_25796,N_25252);
or U26520 (N_26520,N_25367,N_25680);
nand U26521 (N_26521,N_25440,N_25294);
nor U26522 (N_26522,N_25175,N_25049);
nand U26523 (N_26523,N_25111,N_25600);
xnor U26524 (N_26524,N_25344,N_25657);
nor U26525 (N_26525,N_25665,N_25530);
nor U26526 (N_26526,N_25629,N_25604);
or U26527 (N_26527,N_25542,N_25224);
xor U26528 (N_26528,N_25902,N_25591);
nand U26529 (N_26529,N_25745,N_25087);
nand U26530 (N_26530,N_25820,N_25218);
or U26531 (N_26531,N_25241,N_25473);
nand U26532 (N_26532,N_25486,N_25571);
nand U26533 (N_26533,N_25709,N_25496);
nand U26534 (N_26534,N_25857,N_25157);
nand U26535 (N_26535,N_25042,N_25268);
or U26536 (N_26536,N_25028,N_25362);
or U26537 (N_26537,N_25930,N_25992);
nor U26538 (N_26538,N_25036,N_25696);
xor U26539 (N_26539,N_25805,N_25643);
and U26540 (N_26540,N_25466,N_25798);
xor U26541 (N_26541,N_25957,N_25470);
xnor U26542 (N_26542,N_25206,N_25108);
and U26543 (N_26543,N_25605,N_25347);
nor U26544 (N_26544,N_25496,N_25689);
and U26545 (N_26545,N_25072,N_25655);
xor U26546 (N_26546,N_25001,N_25266);
nor U26547 (N_26547,N_25258,N_25140);
or U26548 (N_26548,N_25343,N_25736);
nand U26549 (N_26549,N_25524,N_25450);
nor U26550 (N_26550,N_25867,N_25596);
and U26551 (N_26551,N_25105,N_25471);
and U26552 (N_26552,N_25979,N_25671);
and U26553 (N_26553,N_25332,N_25874);
and U26554 (N_26554,N_25583,N_25676);
xor U26555 (N_26555,N_25023,N_25646);
or U26556 (N_26556,N_25989,N_25925);
nor U26557 (N_26557,N_25945,N_25355);
xnor U26558 (N_26558,N_25827,N_25403);
nand U26559 (N_26559,N_25814,N_25121);
nor U26560 (N_26560,N_25575,N_25732);
xnor U26561 (N_26561,N_25784,N_25415);
nor U26562 (N_26562,N_25350,N_25032);
nor U26563 (N_26563,N_25112,N_25486);
nand U26564 (N_26564,N_25439,N_25451);
nand U26565 (N_26565,N_25843,N_25822);
and U26566 (N_26566,N_25548,N_25668);
nand U26567 (N_26567,N_25212,N_25620);
or U26568 (N_26568,N_25694,N_25950);
and U26569 (N_26569,N_25841,N_25285);
nor U26570 (N_26570,N_25845,N_25419);
xnor U26571 (N_26571,N_25740,N_25493);
and U26572 (N_26572,N_25746,N_25536);
nor U26573 (N_26573,N_25971,N_25914);
or U26574 (N_26574,N_25792,N_25875);
xor U26575 (N_26575,N_25824,N_25646);
or U26576 (N_26576,N_25023,N_25908);
and U26577 (N_26577,N_25164,N_25966);
or U26578 (N_26578,N_25528,N_25935);
xor U26579 (N_26579,N_25251,N_25443);
nor U26580 (N_26580,N_25459,N_25293);
xnor U26581 (N_26581,N_25721,N_25954);
xor U26582 (N_26582,N_25767,N_25232);
xor U26583 (N_26583,N_25466,N_25403);
nand U26584 (N_26584,N_25538,N_25953);
nand U26585 (N_26585,N_25627,N_25654);
nor U26586 (N_26586,N_25930,N_25637);
nor U26587 (N_26587,N_25567,N_25558);
nand U26588 (N_26588,N_25168,N_25008);
xor U26589 (N_26589,N_25506,N_25268);
and U26590 (N_26590,N_25853,N_25077);
nor U26591 (N_26591,N_25121,N_25573);
xor U26592 (N_26592,N_25223,N_25132);
xor U26593 (N_26593,N_25275,N_25654);
xnor U26594 (N_26594,N_25960,N_25919);
nand U26595 (N_26595,N_25367,N_25031);
nand U26596 (N_26596,N_25162,N_25399);
nor U26597 (N_26597,N_25852,N_25190);
or U26598 (N_26598,N_25677,N_25835);
nand U26599 (N_26599,N_25869,N_25387);
and U26600 (N_26600,N_25409,N_25250);
or U26601 (N_26601,N_25243,N_25356);
nor U26602 (N_26602,N_25615,N_25535);
nand U26603 (N_26603,N_25610,N_25576);
nand U26604 (N_26604,N_25170,N_25479);
nor U26605 (N_26605,N_25329,N_25449);
nand U26606 (N_26606,N_25838,N_25311);
xor U26607 (N_26607,N_25883,N_25851);
xnor U26608 (N_26608,N_25066,N_25734);
nor U26609 (N_26609,N_25701,N_25592);
or U26610 (N_26610,N_25270,N_25496);
nand U26611 (N_26611,N_25756,N_25901);
or U26612 (N_26612,N_25135,N_25704);
nor U26613 (N_26613,N_25819,N_25743);
and U26614 (N_26614,N_25452,N_25506);
xor U26615 (N_26615,N_25492,N_25846);
nand U26616 (N_26616,N_25938,N_25232);
or U26617 (N_26617,N_25187,N_25758);
or U26618 (N_26618,N_25964,N_25976);
nand U26619 (N_26619,N_25909,N_25194);
or U26620 (N_26620,N_25459,N_25841);
or U26621 (N_26621,N_25721,N_25386);
or U26622 (N_26622,N_25636,N_25667);
xnor U26623 (N_26623,N_25286,N_25916);
nand U26624 (N_26624,N_25313,N_25099);
nand U26625 (N_26625,N_25478,N_25674);
or U26626 (N_26626,N_25986,N_25321);
xor U26627 (N_26627,N_25144,N_25357);
nor U26628 (N_26628,N_25165,N_25677);
and U26629 (N_26629,N_25778,N_25123);
or U26630 (N_26630,N_25145,N_25193);
nor U26631 (N_26631,N_25779,N_25721);
or U26632 (N_26632,N_25927,N_25392);
nand U26633 (N_26633,N_25609,N_25384);
and U26634 (N_26634,N_25629,N_25489);
nor U26635 (N_26635,N_25348,N_25564);
nand U26636 (N_26636,N_25036,N_25126);
or U26637 (N_26637,N_25566,N_25227);
and U26638 (N_26638,N_25239,N_25809);
and U26639 (N_26639,N_25039,N_25356);
nand U26640 (N_26640,N_25459,N_25523);
and U26641 (N_26641,N_25135,N_25359);
and U26642 (N_26642,N_25940,N_25455);
or U26643 (N_26643,N_25372,N_25200);
nor U26644 (N_26644,N_25204,N_25621);
or U26645 (N_26645,N_25561,N_25511);
xnor U26646 (N_26646,N_25562,N_25443);
and U26647 (N_26647,N_25651,N_25094);
nor U26648 (N_26648,N_25672,N_25559);
or U26649 (N_26649,N_25535,N_25381);
nand U26650 (N_26650,N_25081,N_25315);
or U26651 (N_26651,N_25596,N_25662);
nor U26652 (N_26652,N_25643,N_25284);
xor U26653 (N_26653,N_25245,N_25236);
nor U26654 (N_26654,N_25558,N_25315);
nor U26655 (N_26655,N_25975,N_25171);
and U26656 (N_26656,N_25111,N_25273);
and U26657 (N_26657,N_25124,N_25248);
and U26658 (N_26658,N_25281,N_25401);
or U26659 (N_26659,N_25032,N_25888);
nor U26660 (N_26660,N_25851,N_25828);
nor U26661 (N_26661,N_25224,N_25725);
nand U26662 (N_26662,N_25456,N_25665);
and U26663 (N_26663,N_25154,N_25574);
nand U26664 (N_26664,N_25286,N_25042);
xnor U26665 (N_26665,N_25628,N_25687);
nor U26666 (N_26666,N_25616,N_25885);
nor U26667 (N_26667,N_25646,N_25458);
or U26668 (N_26668,N_25039,N_25010);
and U26669 (N_26669,N_25639,N_25228);
nor U26670 (N_26670,N_25181,N_25073);
and U26671 (N_26671,N_25486,N_25827);
or U26672 (N_26672,N_25543,N_25472);
nor U26673 (N_26673,N_25172,N_25147);
and U26674 (N_26674,N_25734,N_25514);
and U26675 (N_26675,N_25667,N_25123);
xor U26676 (N_26676,N_25919,N_25567);
and U26677 (N_26677,N_25697,N_25103);
or U26678 (N_26678,N_25345,N_25795);
nor U26679 (N_26679,N_25065,N_25104);
or U26680 (N_26680,N_25494,N_25603);
nor U26681 (N_26681,N_25407,N_25314);
nor U26682 (N_26682,N_25371,N_25293);
nor U26683 (N_26683,N_25691,N_25537);
or U26684 (N_26684,N_25792,N_25908);
and U26685 (N_26685,N_25719,N_25214);
and U26686 (N_26686,N_25582,N_25297);
and U26687 (N_26687,N_25613,N_25564);
or U26688 (N_26688,N_25709,N_25109);
or U26689 (N_26689,N_25533,N_25871);
xor U26690 (N_26690,N_25454,N_25126);
xnor U26691 (N_26691,N_25639,N_25877);
or U26692 (N_26692,N_25834,N_25279);
xor U26693 (N_26693,N_25155,N_25864);
nand U26694 (N_26694,N_25506,N_25516);
nand U26695 (N_26695,N_25050,N_25859);
nor U26696 (N_26696,N_25064,N_25361);
and U26697 (N_26697,N_25702,N_25885);
or U26698 (N_26698,N_25812,N_25566);
and U26699 (N_26699,N_25175,N_25831);
nand U26700 (N_26700,N_25994,N_25007);
nand U26701 (N_26701,N_25530,N_25028);
nor U26702 (N_26702,N_25594,N_25985);
and U26703 (N_26703,N_25842,N_25871);
nor U26704 (N_26704,N_25963,N_25727);
nand U26705 (N_26705,N_25178,N_25176);
and U26706 (N_26706,N_25246,N_25806);
nand U26707 (N_26707,N_25556,N_25559);
and U26708 (N_26708,N_25466,N_25449);
or U26709 (N_26709,N_25587,N_25260);
xnor U26710 (N_26710,N_25103,N_25755);
nand U26711 (N_26711,N_25306,N_25343);
nor U26712 (N_26712,N_25059,N_25476);
xnor U26713 (N_26713,N_25610,N_25571);
and U26714 (N_26714,N_25126,N_25279);
and U26715 (N_26715,N_25822,N_25723);
nor U26716 (N_26716,N_25122,N_25872);
or U26717 (N_26717,N_25281,N_25061);
xor U26718 (N_26718,N_25827,N_25472);
and U26719 (N_26719,N_25624,N_25263);
or U26720 (N_26720,N_25612,N_25545);
and U26721 (N_26721,N_25382,N_25059);
and U26722 (N_26722,N_25374,N_25177);
nand U26723 (N_26723,N_25218,N_25626);
xnor U26724 (N_26724,N_25500,N_25124);
nor U26725 (N_26725,N_25374,N_25307);
nor U26726 (N_26726,N_25973,N_25663);
nor U26727 (N_26727,N_25897,N_25252);
nand U26728 (N_26728,N_25576,N_25967);
nor U26729 (N_26729,N_25873,N_25313);
or U26730 (N_26730,N_25520,N_25417);
and U26731 (N_26731,N_25651,N_25584);
nor U26732 (N_26732,N_25543,N_25838);
nand U26733 (N_26733,N_25186,N_25635);
nor U26734 (N_26734,N_25412,N_25312);
nand U26735 (N_26735,N_25536,N_25991);
and U26736 (N_26736,N_25632,N_25617);
or U26737 (N_26737,N_25745,N_25393);
nand U26738 (N_26738,N_25615,N_25008);
or U26739 (N_26739,N_25482,N_25433);
nor U26740 (N_26740,N_25211,N_25615);
xnor U26741 (N_26741,N_25095,N_25476);
nor U26742 (N_26742,N_25624,N_25303);
nor U26743 (N_26743,N_25720,N_25700);
or U26744 (N_26744,N_25603,N_25402);
nand U26745 (N_26745,N_25511,N_25111);
xnor U26746 (N_26746,N_25788,N_25432);
and U26747 (N_26747,N_25103,N_25739);
nor U26748 (N_26748,N_25371,N_25564);
nand U26749 (N_26749,N_25961,N_25430);
and U26750 (N_26750,N_25817,N_25748);
nor U26751 (N_26751,N_25356,N_25636);
nor U26752 (N_26752,N_25650,N_25460);
or U26753 (N_26753,N_25023,N_25345);
or U26754 (N_26754,N_25888,N_25574);
and U26755 (N_26755,N_25172,N_25759);
and U26756 (N_26756,N_25662,N_25176);
and U26757 (N_26757,N_25943,N_25716);
and U26758 (N_26758,N_25301,N_25553);
xnor U26759 (N_26759,N_25427,N_25466);
or U26760 (N_26760,N_25732,N_25916);
and U26761 (N_26761,N_25302,N_25755);
xnor U26762 (N_26762,N_25253,N_25098);
xor U26763 (N_26763,N_25770,N_25924);
nor U26764 (N_26764,N_25381,N_25407);
xor U26765 (N_26765,N_25901,N_25754);
xor U26766 (N_26766,N_25988,N_25075);
and U26767 (N_26767,N_25400,N_25774);
or U26768 (N_26768,N_25004,N_25078);
nand U26769 (N_26769,N_25790,N_25916);
and U26770 (N_26770,N_25554,N_25178);
nor U26771 (N_26771,N_25089,N_25428);
and U26772 (N_26772,N_25594,N_25158);
xnor U26773 (N_26773,N_25961,N_25626);
nand U26774 (N_26774,N_25609,N_25886);
nand U26775 (N_26775,N_25721,N_25830);
nor U26776 (N_26776,N_25950,N_25413);
or U26777 (N_26777,N_25847,N_25576);
or U26778 (N_26778,N_25656,N_25256);
and U26779 (N_26779,N_25678,N_25407);
nand U26780 (N_26780,N_25991,N_25437);
xor U26781 (N_26781,N_25739,N_25985);
and U26782 (N_26782,N_25584,N_25188);
or U26783 (N_26783,N_25392,N_25164);
and U26784 (N_26784,N_25548,N_25008);
or U26785 (N_26785,N_25451,N_25423);
nor U26786 (N_26786,N_25484,N_25543);
and U26787 (N_26787,N_25858,N_25717);
nand U26788 (N_26788,N_25408,N_25415);
or U26789 (N_26789,N_25944,N_25010);
and U26790 (N_26790,N_25666,N_25720);
xor U26791 (N_26791,N_25681,N_25639);
nor U26792 (N_26792,N_25816,N_25166);
nor U26793 (N_26793,N_25551,N_25710);
nor U26794 (N_26794,N_25126,N_25579);
or U26795 (N_26795,N_25682,N_25177);
nand U26796 (N_26796,N_25417,N_25864);
nor U26797 (N_26797,N_25278,N_25376);
nand U26798 (N_26798,N_25505,N_25773);
nand U26799 (N_26799,N_25764,N_25005);
and U26800 (N_26800,N_25143,N_25718);
nor U26801 (N_26801,N_25711,N_25006);
or U26802 (N_26802,N_25636,N_25672);
or U26803 (N_26803,N_25576,N_25461);
or U26804 (N_26804,N_25449,N_25042);
xnor U26805 (N_26805,N_25606,N_25738);
or U26806 (N_26806,N_25875,N_25794);
nor U26807 (N_26807,N_25555,N_25031);
nand U26808 (N_26808,N_25217,N_25510);
nor U26809 (N_26809,N_25029,N_25068);
xor U26810 (N_26810,N_25201,N_25714);
nand U26811 (N_26811,N_25772,N_25568);
and U26812 (N_26812,N_25907,N_25779);
and U26813 (N_26813,N_25476,N_25037);
xnor U26814 (N_26814,N_25037,N_25422);
xnor U26815 (N_26815,N_25532,N_25283);
xor U26816 (N_26816,N_25782,N_25124);
nor U26817 (N_26817,N_25614,N_25481);
or U26818 (N_26818,N_25403,N_25325);
or U26819 (N_26819,N_25496,N_25815);
and U26820 (N_26820,N_25630,N_25629);
and U26821 (N_26821,N_25563,N_25434);
nand U26822 (N_26822,N_25038,N_25727);
or U26823 (N_26823,N_25422,N_25618);
xnor U26824 (N_26824,N_25701,N_25627);
or U26825 (N_26825,N_25898,N_25921);
nand U26826 (N_26826,N_25740,N_25808);
nor U26827 (N_26827,N_25871,N_25811);
and U26828 (N_26828,N_25806,N_25449);
xor U26829 (N_26829,N_25843,N_25383);
and U26830 (N_26830,N_25022,N_25185);
xor U26831 (N_26831,N_25867,N_25579);
nand U26832 (N_26832,N_25235,N_25912);
xor U26833 (N_26833,N_25243,N_25106);
xnor U26834 (N_26834,N_25311,N_25603);
nor U26835 (N_26835,N_25139,N_25829);
xnor U26836 (N_26836,N_25363,N_25620);
and U26837 (N_26837,N_25951,N_25635);
and U26838 (N_26838,N_25642,N_25601);
nand U26839 (N_26839,N_25687,N_25088);
nand U26840 (N_26840,N_25249,N_25141);
and U26841 (N_26841,N_25543,N_25159);
nand U26842 (N_26842,N_25503,N_25315);
xnor U26843 (N_26843,N_25068,N_25475);
nor U26844 (N_26844,N_25087,N_25224);
and U26845 (N_26845,N_25522,N_25294);
and U26846 (N_26846,N_25946,N_25206);
nor U26847 (N_26847,N_25399,N_25595);
and U26848 (N_26848,N_25956,N_25871);
nand U26849 (N_26849,N_25321,N_25309);
nand U26850 (N_26850,N_25435,N_25766);
xor U26851 (N_26851,N_25315,N_25473);
xor U26852 (N_26852,N_25539,N_25548);
xor U26853 (N_26853,N_25907,N_25373);
or U26854 (N_26854,N_25091,N_25942);
or U26855 (N_26855,N_25283,N_25031);
xnor U26856 (N_26856,N_25141,N_25817);
nand U26857 (N_26857,N_25387,N_25558);
xor U26858 (N_26858,N_25873,N_25841);
xor U26859 (N_26859,N_25920,N_25149);
nor U26860 (N_26860,N_25590,N_25722);
nor U26861 (N_26861,N_25734,N_25220);
xor U26862 (N_26862,N_25440,N_25837);
or U26863 (N_26863,N_25112,N_25066);
nor U26864 (N_26864,N_25715,N_25912);
nor U26865 (N_26865,N_25755,N_25196);
nand U26866 (N_26866,N_25017,N_25369);
nor U26867 (N_26867,N_25420,N_25540);
xnor U26868 (N_26868,N_25862,N_25757);
xnor U26869 (N_26869,N_25946,N_25728);
or U26870 (N_26870,N_25474,N_25892);
and U26871 (N_26871,N_25235,N_25060);
nand U26872 (N_26872,N_25182,N_25320);
or U26873 (N_26873,N_25330,N_25314);
nor U26874 (N_26874,N_25078,N_25734);
nor U26875 (N_26875,N_25744,N_25639);
or U26876 (N_26876,N_25310,N_25704);
xnor U26877 (N_26877,N_25746,N_25266);
and U26878 (N_26878,N_25645,N_25540);
and U26879 (N_26879,N_25625,N_25472);
and U26880 (N_26880,N_25706,N_25055);
and U26881 (N_26881,N_25112,N_25284);
and U26882 (N_26882,N_25183,N_25524);
nor U26883 (N_26883,N_25454,N_25519);
nor U26884 (N_26884,N_25752,N_25261);
nand U26885 (N_26885,N_25709,N_25315);
xor U26886 (N_26886,N_25401,N_25566);
xnor U26887 (N_26887,N_25113,N_25075);
nor U26888 (N_26888,N_25829,N_25076);
and U26889 (N_26889,N_25058,N_25267);
and U26890 (N_26890,N_25587,N_25703);
nand U26891 (N_26891,N_25226,N_25945);
and U26892 (N_26892,N_25791,N_25016);
nand U26893 (N_26893,N_25615,N_25466);
nor U26894 (N_26894,N_25412,N_25772);
or U26895 (N_26895,N_25108,N_25716);
nand U26896 (N_26896,N_25122,N_25217);
nor U26897 (N_26897,N_25040,N_25104);
or U26898 (N_26898,N_25930,N_25239);
and U26899 (N_26899,N_25262,N_25721);
xnor U26900 (N_26900,N_25326,N_25917);
and U26901 (N_26901,N_25665,N_25340);
or U26902 (N_26902,N_25069,N_25850);
nor U26903 (N_26903,N_25662,N_25236);
or U26904 (N_26904,N_25645,N_25341);
nand U26905 (N_26905,N_25338,N_25575);
xor U26906 (N_26906,N_25190,N_25879);
xor U26907 (N_26907,N_25234,N_25101);
nand U26908 (N_26908,N_25274,N_25455);
or U26909 (N_26909,N_25771,N_25806);
xor U26910 (N_26910,N_25124,N_25677);
and U26911 (N_26911,N_25920,N_25650);
xor U26912 (N_26912,N_25671,N_25124);
or U26913 (N_26913,N_25409,N_25796);
xor U26914 (N_26914,N_25995,N_25053);
nor U26915 (N_26915,N_25000,N_25848);
xnor U26916 (N_26916,N_25872,N_25688);
and U26917 (N_26917,N_25099,N_25590);
and U26918 (N_26918,N_25539,N_25728);
and U26919 (N_26919,N_25884,N_25962);
and U26920 (N_26920,N_25372,N_25670);
nor U26921 (N_26921,N_25920,N_25895);
and U26922 (N_26922,N_25295,N_25335);
nand U26923 (N_26923,N_25169,N_25569);
xnor U26924 (N_26924,N_25211,N_25524);
xnor U26925 (N_26925,N_25937,N_25129);
xor U26926 (N_26926,N_25268,N_25056);
and U26927 (N_26927,N_25026,N_25778);
nand U26928 (N_26928,N_25626,N_25362);
and U26929 (N_26929,N_25280,N_25493);
and U26930 (N_26930,N_25751,N_25955);
nor U26931 (N_26931,N_25070,N_25091);
nor U26932 (N_26932,N_25861,N_25374);
nand U26933 (N_26933,N_25579,N_25835);
xor U26934 (N_26934,N_25599,N_25053);
nor U26935 (N_26935,N_25794,N_25714);
or U26936 (N_26936,N_25763,N_25708);
xnor U26937 (N_26937,N_25574,N_25467);
or U26938 (N_26938,N_25291,N_25901);
xnor U26939 (N_26939,N_25265,N_25554);
xor U26940 (N_26940,N_25016,N_25597);
and U26941 (N_26941,N_25314,N_25392);
xnor U26942 (N_26942,N_25474,N_25770);
and U26943 (N_26943,N_25540,N_25352);
nand U26944 (N_26944,N_25704,N_25814);
nand U26945 (N_26945,N_25743,N_25341);
xor U26946 (N_26946,N_25034,N_25367);
and U26947 (N_26947,N_25838,N_25570);
and U26948 (N_26948,N_25689,N_25323);
and U26949 (N_26949,N_25070,N_25786);
or U26950 (N_26950,N_25017,N_25305);
nor U26951 (N_26951,N_25082,N_25028);
xnor U26952 (N_26952,N_25185,N_25317);
xor U26953 (N_26953,N_25478,N_25281);
or U26954 (N_26954,N_25331,N_25992);
and U26955 (N_26955,N_25674,N_25659);
nand U26956 (N_26956,N_25064,N_25380);
or U26957 (N_26957,N_25052,N_25948);
or U26958 (N_26958,N_25468,N_25425);
nor U26959 (N_26959,N_25675,N_25429);
xor U26960 (N_26960,N_25410,N_25895);
nand U26961 (N_26961,N_25325,N_25836);
nand U26962 (N_26962,N_25374,N_25170);
nand U26963 (N_26963,N_25654,N_25312);
and U26964 (N_26964,N_25150,N_25256);
nor U26965 (N_26965,N_25996,N_25270);
and U26966 (N_26966,N_25184,N_25046);
nor U26967 (N_26967,N_25352,N_25367);
and U26968 (N_26968,N_25256,N_25350);
or U26969 (N_26969,N_25079,N_25324);
or U26970 (N_26970,N_25855,N_25320);
nor U26971 (N_26971,N_25400,N_25306);
and U26972 (N_26972,N_25273,N_25000);
and U26973 (N_26973,N_25584,N_25792);
xor U26974 (N_26974,N_25340,N_25319);
nand U26975 (N_26975,N_25921,N_25580);
nor U26976 (N_26976,N_25073,N_25922);
nor U26977 (N_26977,N_25915,N_25614);
or U26978 (N_26978,N_25352,N_25265);
and U26979 (N_26979,N_25971,N_25571);
nor U26980 (N_26980,N_25650,N_25169);
nand U26981 (N_26981,N_25465,N_25721);
and U26982 (N_26982,N_25608,N_25794);
nand U26983 (N_26983,N_25510,N_25105);
nor U26984 (N_26984,N_25125,N_25423);
nand U26985 (N_26985,N_25406,N_25557);
nor U26986 (N_26986,N_25679,N_25038);
or U26987 (N_26987,N_25931,N_25510);
xnor U26988 (N_26988,N_25463,N_25738);
nor U26989 (N_26989,N_25379,N_25314);
nor U26990 (N_26990,N_25722,N_25493);
nand U26991 (N_26991,N_25063,N_25442);
or U26992 (N_26992,N_25166,N_25449);
and U26993 (N_26993,N_25976,N_25042);
and U26994 (N_26994,N_25136,N_25329);
xor U26995 (N_26995,N_25641,N_25880);
and U26996 (N_26996,N_25855,N_25646);
nor U26997 (N_26997,N_25938,N_25919);
nand U26998 (N_26998,N_25060,N_25342);
or U26999 (N_26999,N_25006,N_25714);
and U27000 (N_27000,N_26261,N_26766);
nand U27001 (N_27001,N_26622,N_26494);
xor U27002 (N_27002,N_26938,N_26773);
nand U27003 (N_27003,N_26914,N_26923);
or U27004 (N_27004,N_26094,N_26597);
or U27005 (N_27005,N_26279,N_26987);
and U27006 (N_27006,N_26440,N_26876);
and U27007 (N_27007,N_26326,N_26423);
nor U27008 (N_27008,N_26752,N_26591);
xnor U27009 (N_27009,N_26366,N_26902);
nand U27010 (N_27010,N_26727,N_26436);
or U27011 (N_27011,N_26994,N_26697);
and U27012 (N_27012,N_26131,N_26439);
nor U27013 (N_27013,N_26571,N_26629);
xnor U27014 (N_27014,N_26883,N_26768);
xnor U27015 (N_27015,N_26174,N_26551);
or U27016 (N_27016,N_26189,N_26250);
or U27017 (N_27017,N_26302,N_26448);
xnor U27018 (N_27018,N_26529,N_26117);
nor U27019 (N_27019,N_26532,N_26788);
xnor U27020 (N_27020,N_26495,N_26054);
xor U27021 (N_27021,N_26413,N_26889);
nor U27022 (N_27022,N_26787,N_26866);
nand U27023 (N_27023,N_26760,N_26709);
nor U27024 (N_27024,N_26490,N_26926);
xor U27025 (N_27025,N_26941,N_26948);
and U27026 (N_27026,N_26352,N_26184);
xor U27027 (N_27027,N_26193,N_26148);
xor U27028 (N_27028,N_26801,N_26386);
and U27029 (N_27029,N_26980,N_26793);
and U27030 (N_27030,N_26166,N_26910);
nor U27031 (N_27031,N_26882,N_26238);
and U27032 (N_27032,N_26945,N_26735);
and U27033 (N_27033,N_26134,N_26310);
nor U27034 (N_27034,N_26606,N_26668);
and U27035 (N_27035,N_26065,N_26523);
nand U27036 (N_27036,N_26233,N_26008);
nand U27037 (N_27037,N_26960,N_26479);
xor U27038 (N_27038,N_26246,N_26718);
or U27039 (N_27039,N_26730,N_26103);
and U27040 (N_27040,N_26498,N_26916);
or U27041 (N_27041,N_26028,N_26073);
and U27042 (N_27042,N_26828,N_26677);
nand U27043 (N_27043,N_26299,N_26141);
and U27044 (N_27044,N_26743,N_26234);
nand U27045 (N_27045,N_26300,N_26930);
nand U27046 (N_27046,N_26698,N_26149);
nor U27047 (N_27047,N_26821,N_26625);
and U27048 (N_27048,N_26197,N_26936);
xor U27049 (N_27049,N_26818,N_26872);
nor U27050 (N_27050,N_26880,N_26268);
nand U27051 (N_27051,N_26464,N_26628);
xnor U27052 (N_27052,N_26408,N_26181);
nand U27053 (N_27053,N_26617,N_26297);
or U27054 (N_27054,N_26792,N_26833);
xor U27055 (N_27055,N_26483,N_26164);
and U27056 (N_27056,N_26858,N_26087);
xor U27057 (N_27057,N_26685,N_26072);
nor U27058 (N_27058,N_26430,N_26236);
nand U27059 (N_27059,N_26034,N_26319);
and U27060 (N_27060,N_26210,N_26771);
and U27061 (N_27061,N_26273,N_26040);
nand U27062 (N_27062,N_26074,N_26109);
nand U27063 (N_27063,N_26203,N_26558);
xor U27064 (N_27064,N_26586,N_26574);
xor U27065 (N_27065,N_26480,N_26069);
nor U27066 (N_27066,N_26006,N_26675);
and U27067 (N_27067,N_26982,N_26604);
nor U27068 (N_27068,N_26165,N_26043);
nor U27069 (N_27069,N_26294,N_26126);
nand U27070 (N_27070,N_26449,N_26021);
xor U27071 (N_27071,N_26831,N_26857);
nand U27072 (N_27072,N_26213,N_26224);
nor U27073 (N_27073,N_26135,N_26282);
nor U27074 (N_27074,N_26393,N_26318);
or U27075 (N_27075,N_26284,N_26999);
xor U27076 (N_27076,N_26847,N_26355);
and U27077 (N_27077,N_26075,N_26438);
xnor U27078 (N_27078,N_26239,N_26777);
nand U27079 (N_27079,N_26229,N_26437);
or U27080 (N_27080,N_26637,N_26200);
or U27081 (N_27081,N_26272,N_26425);
xnor U27082 (N_27082,N_26410,N_26487);
and U27083 (N_27083,N_26489,N_26886);
nand U27084 (N_27084,N_26461,N_26548);
and U27085 (N_27085,N_26559,N_26688);
nor U27086 (N_27086,N_26429,N_26491);
xnor U27087 (N_27087,N_26589,N_26156);
xnor U27088 (N_27088,N_26863,N_26391);
xnor U27089 (N_27089,N_26089,N_26255);
and U27090 (N_27090,N_26925,N_26751);
nor U27091 (N_27091,N_26368,N_26961);
nor U27092 (N_27092,N_26953,N_26879);
and U27093 (N_27093,N_26854,N_26515);
and U27094 (N_27094,N_26262,N_26747);
nand U27095 (N_27095,N_26292,N_26819);
and U27096 (N_27096,N_26922,N_26802);
xor U27097 (N_27097,N_26305,N_26765);
and U27098 (N_27098,N_26701,N_26612);
or U27099 (N_27099,N_26542,N_26965);
nand U27100 (N_27100,N_26599,N_26023);
and U27101 (N_27101,N_26215,N_26728);
nor U27102 (N_27102,N_26014,N_26151);
nand U27103 (N_27103,N_26419,N_26139);
or U27104 (N_27104,N_26125,N_26600);
nand U27105 (N_27105,N_26850,N_26578);
nand U27106 (N_27106,N_26387,N_26614);
and U27107 (N_27107,N_26372,N_26107);
nor U27108 (N_27108,N_26003,N_26144);
xor U27109 (N_27109,N_26052,N_26270);
xor U27110 (N_27110,N_26803,N_26679);
nand U27111 (N_27111,N_26114,N_26442);
nor U27112 (N_27112,N_26903,N_26807);
xnor U27113 (N_27113,N_26967,N_26281);
and U27114 (N_27114,N_26564,N_26348);
and U27115 (N_27115,N_26993,N_26186);
and U27116 (N_27116,N_26647,N_26266);
or U27117 (N_27117,N_26984,N_26301);
nor U27118 (N_27118,N_26457,N_26811);
or U27119 (N_27119,N_26650,N_26885);
and U27120 (N_27120,N_26039,N_26864);
nand U27121 (N_27121,N_26015,N_26211);
nand U27122 (N_27122,N_26737,N_26570);
nand U27123 (N_27123,N_26544,N_26526);
nand U27124 (N_27124,N_26700,N_26092);
or U27125 (N_27125,N_26509,N_26264);
or U27126 (N_27126,N_26082,N_26051);
xor U27127 (N_27127,N_26106,N_26928);
nand U27128 (N_27128,N_26329,N_26293);
or U27129 (N_27129,N_26682,N_26976);
and U27130 (N_27130,N_26549,N_26537);
xnor U27131 (N_27131,N_26363,N_26518);
nand U27132 (N_27132,N_26424,N_26340);
or U27133 (N_27133,N_26991,N_26814);
and U27134 (N_27134,N_26096,N_26249);
nor U27135 (N_27135,N_26108,N_26192);
xor U27136 (N_27136,N_26772,N_26669);
nor U27137 (N_27137,N_26603,N_26001);
xnor U27138 (N_27138,N_26050,N_26188);
nand U27139 (N_27139,N_26513,N_26016);
nor U27140 (N_27140,N_26180,N_26013);
nand U27141 (N_27141,N_26175,N_26163);
and U27142 (N_27142,N_26749,N_26426);
nor U27143 (N_27143,N_26733,N_26502);
and U27144 (N_27144,N_26855,N_26196);
nor U27145 (N_27145,N_26009,N_26214);
xnor U27146 (N_27146,N_26704,N_26547);
and U27147 (N_27147,N_26573,N_26970);
and U27148 (N_27148,N_26759,N_26332);
and U27149 (N_27149,N_26045,N_26198);
xnor U27150 (N_27150,N_26160,N_26243);
nor U27151 (N_27151,N_26252,N_26610);
nor U27152 (N_27152,N_26232,N_26240);
or U27153 (N_27153,N_26365,N_26929);
nand U27154 (N_27154,N_26983,N_26382);
nor U27155 (N_27155,N_26584,N_26183);
nor U27156 (N_27156,N_26639,N_26177);
and U27157 (N_27157,N_26271,N_26315);
xor U27158 (N_27158,N_26157,N_26690);
or U27159 (N_27159,N_26477,N_26694);
xnor U27160 (N_27160,N_26815,N_26036);
xnor U27161 (N_27161,N_26228,N_26744);
nand U27162 (N_27162,N_26101,N_26593);
or U27163 (N_27163,N_26364,N_26732);
and U27164 (N_27164,N_26714,N_26711);
or U27165 (N_27165,N_26935,N_26343);
and U27166 (N_27166,N_26746,N_26588);
and U27167 (N_27167,N_26396,N_26371);
nand U27168 (N_27168,N_26358,N_26167);
or U27169 (N_27169,N_26323,N_26949);
xnor U27170 (N_27170,N_26066,N_26415);
nand U27171 (N_27171,N_26624,N_26385);
nor U27172 (N_27172,N_26900,N_26607);
nand U27173 (N_27173,N_26826,N_26781);
nand U27174 (N_27174,N_26660,N_26404);
or U27175 (N_27175,N_26877,N_26245);
or U27176 (N_27176,N_26486,N_26680);
nand U27177 (N_27177,N_26140,N_26116);
nor U27178 (N_27178,N_26966,N_26105);
nand U27179 (N_27179,N_26247,N_26152);
or U27180 (N_27180,N_26875,N_26869);
nor U27181 (N_27181,N_26029,N_26241);
nor U27182 (N_27182,N_26905,N_26510);
nor U27183 (N_27183,N_26753,N_26538);
nand U27184 (N_27184,N_26920,N_26789);
and U27185 (N_27185,N_26652,N_26353);
nor U27186 (N_27186,N_26434,N_26964);
and U27187 (N_27187,N_26467,N_26068);
nand U27188 (N_27188,N_26049,N_26360);
and U27189 (N_27189,N_26286,N_26962);
or U27190 (N_27190,N_26018,N_26235);
nand U27191 (N_27191,N_26204,N_26002);
or U27192 (N_27192,N_26522,N_26626);
and U27193 (N_27193,N_26379,N_26859);
or U27194 (N_27194,N_26012,N_26492);
and U27195 (N_27195,N_26808,N_26825);
xnor U27196 (N_27196,N_26761,N_26525);
nor U27197 (N_27197,N_26102,N_26579);
nor U27198 (N_27198,N_26673,N_26779);
nor U27199 (N_27199,N_26635,N_26507);
xnor U27200 (N_27200,N_26758,N_26137);
nor U27201 (N_27201,N_26695,N_26242);
or U27202 (N_27202,N_26934,N_26552);
xor U27203 (N_27203,N_26696,N_26774);
or U27204 (N_27204,N_26767,N_26031);
nand U27205 (N_27205,N_26325,N_26474);
xnor U27206 (N_27206,N_26806,N_26741);
nor U27207 (N_27207,N_26170,N_26451);
nand U27208 (N_27208,N_26011,N_26540);
nor U27209 (N_27209,N_26832,N_26985);
xnor U27210 (N_27210,N_26959,N_26988);
xnor U27211 (N_27211,N_26873,N_26172);
nand U27212 (N_27212,N_26783,N_26511);
xnor U27213 (N_27213,N_26699,N_26534);
and U27214 (N_27214,N_26158,N_26121);
nor U27215 (N_27215,N_26208,N_26800);
xnor U27216 (N_27216,N_26336,N_26500);
nor U27217 (N_27217,N_26745,N_26084);
and U27218 (N_27218,N_26596,N_26621);
or U27219 (N_27219,N_26689,N_26503);
xnor U27220 (N_27220,N_26453,N_26473);
xor U27221 (N_27221,N_26226,N_26136);
and U27222 (N_27222,N_26852,N_26981);
or U27223 (N_27223,N_26078,N_26088);
nor U27224 (N_27224,N_26796,N_26918);
or U27225 (N_27225,N_26499,N_26356);
and U27226 (N_27226,N_26038,N_26159);
and U27227 (N_27227,N_26260,N_26362);
xor U27228 (N_27228,N_26100,N_26963);
and U27229 (N_27229,N_26007,N_26799);
and U27230 (N_27230,N_26894,N_26390);
nor U27231 (N_27231,N_26561,N_26230);
nor U27232 (N_27232,N_26638,N_26575);
and U27233 (N_27233,N_26402,N_26508);
xnor U27234 (N_27234,N_26354,N_26658);
nor U27235 (N_27235,N_26615,N_26025);
or U27236 (N_27236,N_26707,N_26587);
nand U27237 (N_27237,N_26345,N_26968);
and U27238 (N_27238,N_26418,N_26071);
or U27239 (N_27239,N_26032,N_26901);
and U27240 (N_27240,N_26915,N_26738);
and U27241 (N_27241,N_26291,N_26394);
nor U27242 (N_27242,N_26085,N_26651);
xor U27243 (N_27243,N_26784,N_26952);
nor U27244 (N_27244,N_26443,N_26304);
or U27245 (N_27245,N_26095,N_26602);
nor U27246 (N_27246,N_26601,N_26056);
xor U27247 (N_27247,N_26583,N_26342);
xnor U27248 (N_27248,N_26462,N_26795);
nand U27249 (N_27249,N_26311,N_26566);
and U27250 (N_27250,N_26339,N_26904);
xor U27251 (N_27251,N_26762,N_26205);
nor U27252 (N_27252,N_26545,N_26409);
nor U27253 (N_27253,N_26401,N_26667);
or U27254 (N_27254,N_26659,N_26527);
and U27255 (N_27255,N_26947,N_26620);
and U27256 (N_27256,N_26937,N_26162);
and U27257 (N_27257,N_26267,N_26729);
nor U27258 (N_27258,N_26455,N_26757);
nand U27259 (N_27259,N_26130,N_26791);
nand U27260 (N_27260,N_26562,N_26389);
nand U27261 (N_27261,N_26168,N_26324);
xnor U27262 (N_27262,N_26590,N_26259);
or U27263 (N_27263,N_26836,N_26520);
and U27264 (N_27264,N_26568,N_26878);
and U27265 (N_27265,N_26161,N_26307);
and U27266 (N_27266,N_26063,N_26898);
nor U27267 (N_27267,N_26496,N_26388);
nand U27268 (N_27268,N_26046,N_26576);
or U27269 (N_27269,N_26070,N_26227);
or U27270 (N_27270,N_26640,N_26906);
xnor U27271 (N_27271,N_26581,N_26124);
and U27272 (N_27272,N_26684,N_26219);
nor U27273 (N_27273,N_26506,N_26944);
and U27274 (N_27274,N_26222,N_26790);
and U27275 (N_27275,N_26153,N_26539);
or U27276 (N_27276,N_26725,N_26090);
and U27277 (N_27277,N_26335,N_26829);
nand U27278 (N_27278,N_26731,N_26104);
or U27279 (N_27279,N_26664,N_26411);
or U27280 (N_27280,N_26557,N_26816);
xnor U27281 (N_27281,N_26719,N_26482);
and U27282 (N_27282,N_26110,N_26739);
and U27283 (N_27283,N_26010,N_26027);
and U27284 (N_27284,N_26687,N_26917);
nor U27285 (N_27285,N_26907,N_26654);
and U27286 (N_27286,N_26672,N_26572);
and U27287 (N_27287,N_26649,N_26890);
nand U27288 (N_27288,N_26950,N_26810);
or U27289 (N_27289,N_26061,N_26838);
xnor U27290 (N_27290,N_26320,N_26035);
nand U27291 (N_27291,N_26077,N_26662);
xnor U27292 (N_27292,N_26887,N_26567);
xnor U27293 (N_27293,N_26417,N_26331);
nand U27294 (N_27294,N_26517,N_26083);
xnor U27295 (N_27295,N_26516,N_26710);
or U27296 (N_27296,N_26861,N_26721);
or U27297 (N_27297,N_26447,N_26111);
or U27298 (N_27298,N_26627,N_26399);
xor U27299 (N_27299,N_26406,N_26283);
nand U27300 (N_27300,N_26716,N_26726);
and U27301 (N_27301,N_26835,N_26550);
nor U27302 (N_27302,N_26862,N_26535);
nor U27303 (N_27303,N_26809,N_26099);
xor U27304 (N_27304,N_26265,N_26780);
nor U27305 (N_27305,N_26359,N_26909);
nor U27306 (N_27306,N_26512,N_26113);
nor U27307 (N_27307,N_26972,N_26805);
xnor U27308 (N_27308,N_26374,N_26059);
nand U27309 (N_27309,N_26846,N_26373);
or U27310 (N_27310,N_26642,N_26996);
or U27311 (N_27311,N_26093,N_26865);
nor U27312 (N_27312,N_26750,N_26998);
and U27313 (N_27313,N_26048,N_26251);
xnor U27314 (N_27314,N_26017,N_26956);
nor U27315 (N_27315,N_26755,N_26954);
and U27316 (N_27316,N_26403,N_26853);
xor U27317 (N_27317,N_26951,N_26543);
nand U27318 (N_27318,N_26913,N_26648);
xor U27319 (N_27319,N_26287,N_26715);
nor U27320 (N_27320,N_26636,N_26308);
xnor U27321 (N_27321,N_26127,N_26813);
xnor U27322 (N_27322,N_26632,N_26288);
or U27323 (N_27323,N_26475,N_26276);
and U27324 (N_27324,N_26678,N_26724);
or U27325 (N_27325,N_26185,N_26871);
or U27326 (N_27326,N_26493,N_26431);
or U27327 (N_27327,N_26908,N_26098);
nand U27328 (N_27328,N_26171,N_26663);
and U27329 (N_27329,N_26633,N_26874);
nand U27330 (N_27330,N_26969,N_26849);
and U27331 (N_27331,N_26129,N_26830);
and U27332 (N_27332,N_26646,N_26536);
nand U27333 (N_27333,N_26764,N_26702);
nand U27334 (N_27334,N_26361,N_26142);
or U27335 (N_27335,N_26081,N_26469);
xnor U27336 (N_27336,N_26316,N_26782);
nand U27337 (N_27337,N_26313,N_26921);
nand U27338 (N_27338,N_26786,N_26565);
nor U27339 (N_27339,N_26037,N_26296);
and U27340 (N_27340,N_26756,N_26618);
or U27341 (N_27341,N_26097,N_26258);
xor U27342 (N_27342,N_26497,N_26427);
and U27343 (N_27343,N_26519,N_26881);
nand U27344 (N_27344,N_26661,N_26720);
and U27345 (N_27345,N_26533,N_26312);
and U27346 (N_27346,N_26504,N_26369);
nor U27347 (N_27347,N_26754,N_26531);
xnor U27348 (N_27348,N_26563,N_26452);
xor U27349 (N_27349,N_26717,N_26884);
or U27350 (N_27350,N_26553,N_26178);
xor U27351 (N_27351,N_26692,N_26609);
xnor U27352 (N_27352,N_26804,N_26303);
nor U27353 (N_27353,N_26416,N_26631);
xor U27354 (N_27354,N_26693,N_26560);
nor U27355 (N_27355,N_26514,N_26785);
or U27356 (N_27356,N_26367,N_26770);
nand U27357 (N_27357,N_26263,N_26841);
nor U27358 (N_27358,N_26641,N_26115);
and U27359 (N_27359,N_26986,N_26444);
and U27360 (N_27360,N_26556,N_26932);
and U27361 (N_27361,N_26524,N_26798);
and U27362 (N_27362,N_26997,N_26407);
and U27363 (N_27363,N_26856,N_26120);
or U27364 (N_27364,N_26278,N_26223);
nor U27365 (N_27365,N_26338,N_26195);
xor U27366 (N_27366,N_26594,N_26657);
or U27367 (N_27367,N_26740,N_26280);
xnor U27368 (N_27368,N_26943,N_26895);
nand U27369 (N_27369,N_26187,N_26398);
and U27370 (N_27370,N_26257,N_26441);
nand U27371 (N_27371,N_26942,N_26484);
xor U27372 (N_27372,N_26817,N_26653);
or U27373 (N_27373,N_26346,N_26957);
nor U27374 (N_27374,N_26674,N_26256);
or U27375 (N_27375,N_26955,N_26843);
nand U27376 (N_27376,N_26445,N_26703);
nor U27377 (N_27377,N_26199,N_26191);
xnor U27378 (N_27378,N_26145,N_26979);
nor U27379 (N_27379,N_26897,N_26079);
and U27380 (N_27380,N_26220,N_26505);
nor U27381 (N_27381,N_26207,N_26611);
and U27382 (N_27382,N_26026,N_26501);
nand U27383 (N_27383,N_26309,N_26004);
xnor U27384 (N_27384,N_26824,N_26577);
and U27385 (N_27385,N_26582,N_26823);
nor U27386 (N_27386,N_26041,N_26488);
and U27387 (N_27387,N_26327,N_26975);
nand U27388 (N_27388,N_26289,N_26691);
nor U27389 (N_27389,N_26778,N_26169);
nand U27390 (N_27390,N_26958,N_26468);
or U27391 (N_27391,N_26734,N_26939);
xnor U27392 (N_27392,N_26794,N_26712);
nand U27393 (N_27393,N_26086,N_26554);
or U27394 (N_27394,N_26891,N_26713);
nand U27395 (N_27395,N_26446,N_26067);
or U27396 (N_27396,N_26030,N_26769);
and U27397 (N_27397,N_26397,N_26321);
nor U27398 (N_27398,N_26924,N_26822);
nor U27399 (N_27399,N_26400,N_26676);
or U27400 (N_27400,N_26655,N_26912);
and U27401 (N_27401,N_26645,N_26432);
nand U27402 (N_27402,N_26275,N_26990);
nor U27403 (N_27403,N_26112,N_26080);
and U27404 (N_27404,N_26834,N_26033);
and U27405 (N_27405,N_26351,N_26206);
or U27406 (N_27406,N_26024,N_26179);
xor U27407 (N_27407,N_26209,N_26347);
or U27408 (N_27408,N_26919,N_26459);
nand U27409 (N_27409,N_26306,N_26244);
and U27410 (N_27410,N_26630,N_26119);
nor U27411 (N_27411,N_26763,N_26330);
nand U27412 (N_27412,N_26465,N_26867);
nand U27413 (N_27413,N_26123,N_26995);
nand U27414 (N_27414,N_26370,N_26005);
nand U27415 (N_27415,N_26062,N_26665);
xor U27416 (N_27416,N_26060,N_26128);
nor U27417 (N_27417,N_26269,N_26435);
and U27418 (N_27418,N_26421,N_26019);
or U27419 (N_27419,N_26290,N_26931);
nor U27420 (N_27420,N_26454,N_26091);
and U27421 (N_27421,N_26405,N_26064);
and U27422 (N_27422,N_26349,N_26201);
nand U27423 (N_27423,N_26595,N_26940);
xnor U27424 (N_27424,N_26476,N_26053);
xnor U27425 (N_27425,N_26585,N_26322);
nor U27426 (N_27426,N_26253,N_26608);
nor U27427 (N_27427,N_26458,N_26118);
nor U27428 (N_27428,N_26182,N_26971);
nand U27429 (N_27429,N_26055,N_26428);
or U27430 (N_27430,N_26380,N_26892);
nor U27431 (N_27431,N_26317,N_26328);
or U27432 (N_27432,N_26216,N_26295);
xor U27433 (N_27433,N_26671,N_26237);
and U27434 (N_27434,N_26381,N_26973);
nor U27435 (N_27435,N_26616,N_26977);
nor U27436 (N_27436,N_26845,N_26057);
and U27437 (N_27437,N_26619,N_26470);
nor U27438 (N_27438,N_26058,N_26132);
nor U27439 (N_27439,N_26022,N_26978);
or U27440 (N_27440,N_26143,N_26974);
nor U27441 (N_27441,N_26357,N_26422);
and U27442 (N_27442,N_26530,N_26350);
nand U27443 (N_27443,N_26541,N_26569);
or U27444 (N_27444,N_26231,N_26314);
nor U27445 (N_27445,N_26274,N_26202);
or U27446 (N_27446,N_26133,N_26644);
or U27447 (N_27447,N_26384,N_26333);
nor U27448 (N_27448,N_26992,N_26686);
xnor U27449 (N_27449,N_26723,N_26217);
and U27450 (N_27450,N_26285,N_26375);
xnor U27451 (N_27451,N_26122,N_26592);
or U27452 (N_27452,N_26225,N_26154);
xor U27453 (N_27453,N_26989,N_26463);
nor U27454 (N_27454,N_26248,N_26748);
and U27455 (N_27455,N_26946,N_26471);
nor U27456 (N_27456,N_26546,N_26708);
and U27457 (N_27457,N_26146,N_26722);
and U27458 (N_27458,N_26000,N_26742);
nand U27459 (N_27459,N_26481,N_26776);
xnor U27460 (N_27460,N_26681,N_26298);
and U27461 (N_27461,N_26221,N_26666);
nand U27462 (N_27462,N_26190,N_26888);
nor U27463 (N_27463,N_26839,N_26848);
nor U27464 (N_27464,N_26218,N_26860);
xnor U27465 (N_27465,N_26334,N_26705);
or U27466 (N_27466,N_26383,N_26472);
nor U27467 (N_27467,N_26155,N_26842);
nor U27468 (N_27468,N_26683,N_26837);
or U27469 (N_27469,N_26377,N_26775);
nor U27470 (N_27470,N_26076,N_26605);
xnor U27471 (N_27471,N_26412,N_26706);
nor U27472 (N_27472,N_26844,N_26797);
xor U27473 (N_27473,N_26840,N_26414);
or U27474 (N_27474,N_26820,N_26042);
or U27475 (N_27475,N_26376,N_26392);
and U27476 (N_27476,N_26337,N_26868);
nor U27477 (N_27477,N_26047,N_26812);
nand U27478 (N_27478,N_26623,N_26044);
nor U27479 (N_27479,N_26521,N_26634);
xor U27480 (N_27480,N_26254,N_26147);
or U27481 (N_27481,N_26456,N_26194);
xnor U27482 (N_27482,N_26893,N_26643);
nor U27483 (N_27483,N_26670,N_26466);
or U27484 (N_27484,N_26378,N_26460);
nand U27485 (N_27485,N_26020,N_26420);
and U27486 (N_27486,N_26176,N_26613);
and U27487 (N_27487,N_26212,N_26555);
and U27488 (N_27488,N_26138,N_26870);
and U27489 (N_27489,N_26344,N_26736);
nand U27490 (N_27490,N_26341,N_26173);
nor U27491 (N_27491,N_26150,N_26933);
xor U27492 (N_27492,N_26656,N_26478);
or U27493 (N_27493,N_26450,N_26485);
nor U27494 (N_27494,N_26580,N_26598);
or U27495 (N_27495,N_26528,N_26851);
nand U27496 (N_27496,N_26433,N_26395);
nand U27497 (N_27497,N_26896,N_26899);
nand U27498 (N_27498,N_26911,N_26927);
nor U27499 (N_27499,N_26277,N_26827);
nor U27500 (N_27500,N_26755,N_26462);
nor U27501 (N_27501,N_26777,N_26487);
and U27502 (N_27502,N_26801,N_26305);
or U27503 (N_27503,N_26789,N_26928);
nand U27504 (N_27504,N_26921,N_26726);
and U27505 (N_27505,N_26331,N_26118);
and U27506 (N_27506,N_26107,N_26324);
or U27507 (N_27507,N_26098,N_26495);
nor U27508 (N_27508,N_26623,N_26587);
nor U27509 (N_27509,N_26516,N_26465);
or U27510 (N_27510,N_26764,N_26045);
xnor U27511 (N_27511,N_26596,N_26431);
nor U27512 (N_27512,N_26762,N_26258);
and U27513 (N_27513,N_26381,N_26885);
xnor U27514 (N_27514,N_26271,N_26639);
and U27515 (N_27515,N_26431,N_26011);
xnor U27516 (N_27516,N_26426,N_26587);
nor U27517 (N_27517,N_26283,N_26541);
or U27518 (N_27518,N_26125,N_26827);
nor U27519 (N_27519,N_26973,N_26465);
and U27520 (N_27520,N_26239,N_26415);
xor U27521 (N_27521,N_26667,N_26551);
and U27522 (N_27522,N_26010,N_26636);
and U27523 (N_27523,N_26555,N_26990);
nor U27524 (N_27524,N_26407,N_26851);
or U27525 (N_27525,N_26515,N_26013);
xnor U27526 (N_27526,N_26208,N_26343);
nand U27527 (N_27527,N_26141,N_26230);
xnor U27528 (N_27528,N_26742,N_26162);
and U27529 (N_27529,N_26422,N_26951);
xnor U27530 (N_27530,N_26171,N_26654);
and U27531 (N_27531,N_26085,N_26504);
and U27532 (N_27532,N_26538,N_26546);
or U27533 (N_27533,N_26773,N_26661);
nand U27534 (N_27534,N_26154,N_26594);
nor U27535 (N_27535,N_26504,N_26869);
or U27536 (N_27536,N_26923,N_26989);
nand U27537 (N_27537,N_26101,N_26438);
nand U27538 (N_27538,N_26171,N_26820);
and U27539 (N_27539,N_26342,N_26841);
or U27540 (N_27540,N_26629,N_26440);
and U27541 (N_27541,N_26487,N_26914);
or U27542 (N_27542,N_26895,N_26707);
nor U27543 (N_27543,N_26710,N_26730);
xnor U27544 (N_27544,N_26582,N_26576);
xnor U27545 (N_27545,N_26143,N_26372);
xor U27546 (N_27546,N_26207,N_26938);
nand U27547 (N_27547,N_26240,N_26740);
nor U27548 (N_27548,N_26631,N_26548);
and U27549 (N_27549,N_26796,N_26440);
or U27550 (N_27550,N_26107,N_26078);
xnor U27551 (N_27551,N_26748,N_26127);
nand U27552 (N_27552,N_26842,N_26374);
and U27553 (N_27553,N_26297,N_26605);
or U27554 (N_27554,N_26046,N_26018);
nand U27555 (N_27555,N_26228,N_26269);
or U27556 (N_27556,N_26227,N_26416);
xor U27557 (N_27557,N_26963,N_26096);
nor U27558 (N_27558,N_26317,N_26866);
and U27559 (N_27559,N_26202,N_26128);
and U27560 (N_27560,N_26889,N_26065);
nand U27561 (N_27561,N_26046,N_26026);
and U27562 (N_27562,N_26029,N_26987);
nor U27563 (N_27563,N_26500,N_26135);
xnor U27564 (N_27564,N_26143,N_26804);
xor U27565 (N_27565,N_26722,N_26608);
nor U27566 (N_27566,N_26520,N_26064);
or U27567 (N_27567,N_26859,N_26003);
xnor U27568 (N_27568,N_26878,N_26170);
and U27569 (N_27569,N_26901,N_26646);
and U27570 (N_27570,N_26218,N_26841);
and U27571 (N_27571,N_26282,N_26272);
nor U27572 (N_27572,N_26481,N_26129);
nor U27573 (N_27573,N_26166,N_26744);
or U27574 (N_27574,N_26939,N_26055);
nand U27575 (N_27575,N_26024,N_26188);
nand U27576 (N_27576,N_26475,N_26549);
and U27577 (N_27577,N_26460,N_26286);
or U27578 (N_27578,N_26708,N_26153);
or U27579 (N_27579,N_26563,N_26684);
or U27580 (N_27580,N_26089,N_26809);
nand U27581 (N_27581,N_26406,N_26553);
or U27582 (N_27582,N_26702,N_26673);
xor U27583 (N_27583,N_26017,N_26112);
xor U27584 (N_27584,N_26952,N_26465);
or U27585 (N_27585,N_26378,N_26953);
or U27586 (N_27586,N_26275,N_26485);
nor U27587 (N_27587,N_26572,N_26541);
or U27588 (N_27588,N_26410,N_26965);
xor U27589 (N_27589,N_26575,N_26480);
nor U27590 (N_27590,N_26185,N_26460);
and U27591 (N_27591,N_26703,N_26333);
nand U27592 (N_27592,N_26277,N_26455);
or U27593 (N_27593,N_26359,N_26301);
nor U27594 (N_27594,N_26128,N_26068);
nand U27595 (N_27595,N_26554,N_26886);
and U27596 (N_27596,N_26451,N_26014);
nor U27597 (N_27597,N_26037,N_26969);
nand U27598 (N_27598,N_26622,N_26315);
and U27599 (N_27599,N_26288,N_26830);
nor U27600 (N_27600,N_26352,N_26173);
nor U27601 (N_27601,N_26030,N_26454);
xnor U27602 (N_27602,N_26252,N_26449);
or U27603 (N_27603,N_26456,N_26633);
xor U27604 (N_27604,N_26203,N_26378);
or U27605 (N_27605,N_26942,N_26769);
and U27606 (N_27606,N_26128,N_26264);
nor U27607 (N_27607,N_26327,N_26889);
xnor U27608 (N_27608,N_26162,N_26459);
or U27609 (N_27609,N_26209,N_26879);
or U27610 (N_27610,N_26495,N_26449);
nand U27611 (N_27611,N_26390,N_26275);
xor U27612 (N_27612,N_26327,N_26750);
xor U27613 (N_27613,N_26360,N_26318);
nor U27614 (N_27614,N_26507,N_26295);
nand U27615 (N_27615,N_26393,N_26437);
xor U27616 (N_27616,N_26019,N_26830);
nor U27617 (N_27617,N_26621,N_26737);
xnor U27618 (N_27618,N_26551,N_26687);
nand U27619 (N_27619,N_26879,N_26732);
nand U27620 (N_27620,N_26643,N_26439);
xor U27621 (N_27621,N_26570,N_26251);
nor U27622 (N_27622,N_26791,N_26515);
or U27623 (N_27623,N_26368,N_26128);
nand U27624 (N_27624,N_26122,N_26423);
or U27625 (N_27625,N_26991,N_26543);
nand U27626 (N_27626,N_26221,N_26654);
or U27627 (N_27627,N_26113,N_26736);
nand U27628 (N_27628,N_26070,N_26023);
nor U27629 (N_27629,N_26030,N_26308);
or U27630 (N_27630,N_26608,N_26464);
xor U27631 (N_27631,N_26258,N_26998);
or U27632 (N_27632,N_26647,N_26091);
nand U27633 (N_27633,N_26053,N_26729);
nand U27634 (N_27634,N_26381,N_26021);
xor U27635 (N_27635,N_26785,N_26747);
nor U27636 (N_27636,N_26471,N_26151);
nand U27637 (N_27637,N_26785,N_26315);
nor U27638 (N_27638,N_26363,N_26690);
or U27639 (N_27639,N_26881,N_26385);
xnor U27640 (N_27640,N_26115,N_26434);
or U27641 (N_27641,N_26298,N_26474);
and U27642 (N_27642,N_26954,N_26669);
and U27643 (N_27643,N_26031,N_26204);
nor U27644 (N_27644,N_26991,N_26316);
and U27645 (N_27645,N_26561,N_26106);
and U27646 (N_27646,N_26032,N_26125);
or U27647 (N_27647,N_26818,N_26083);
nor U27648 (N_27648,N_26150,N_26788);
or U27649 (N_27649,N_26373,N_26614);
nand U27650 (N_27650,N_26197,N_26610);
and U27651 (N_27651,N_26271,N_26941);
xor U27652 (N_27652,N_26744,N_26116);
nor U27653 (N_27653,N_26309,N_26734);
nor U27654 (N_27654,N_26259,N_26886);
xor U27655 (N_27655,N_26175,N_26534);
and U27656 (N_27656,N_26857,N_26983);
nor U27657 (N_27657,N_26967,N_26346);
xnor U27658 (N_27658,N_26295,N_26509);
nand U27659 (N_27659,N_26088,N_26824);
xnor U27660 (N_27660,N_26423,N_26333);
nand U27661 (N_27661,N_26470,N_26581);
and U27662 (N_27662,N_26831,N_26488);
and U27663 (N_27663,N_26550,N_26140);
or U27664 (N_27664,N_26754,N_26396);
nor U27665 (N_27665,N_26368,N_26362);
and U27666 (N_27666,N_26068,N_26165);
nand U27667 (N_27667,N_26595,N_26093);
or U27668 (N_27668,N_26831,N_26588);
nand U27669 (N_27669,N_26376,N_26269);
nor U27670 (N_27670,N_26149,N_26749);
or U27671 (N_27671,N_26825,N_26112);
or U27672 (N_27672,N_26233,N_26147);
or U27673 (N_27673,N_26976,N_26326);
xnor U27674 (N_27674,N_26453,N_26909);
xnor U27675 (N_27675,N_26237,N_26778);
and U27676 (N_27676,N_26749,N_26575);
or U27677 (N_27677,N_26263,N_26634);
nand U27678 (N_27678,N_26445,N_26868);
and U27679 (N_27679,N_26081,N_26851);
nor U27680 (N_27680,N_26356,N_26781);
and U27681 (N_27681,N_26287,N_26366);
nand U27682 (N_27682,N_26651,N_26897);
and U27683 (N_27683,N_26552,N_26527);
nand U27684 (N_27684,N_26984,N_26573);
nand U27685 (N_27685,N_26255,N_26234);
or U27686 (N_27686,N_26439,N_26540);
and U27687 (N_27687,N_26876,N_26139);
or U27688 (N_27688,N_26504,N_26176);
and U27689 (N_27689,N_26545,N_26668);
nor U27690 (N_27690,N_26019,N_26471);
and U27691 (N_27691,N_26049,N_26013);
nor U27692 (N_27692,N_26654,N_26287);
xnor U27693 (N_27693,N_26134,N_26658);
nand U27694 (N_27694,N_26044,N_26145);
and U27695 (N_27695,N_26679,N_26267);
xor U27696 (N_27696,N_26785,N_26790);
xnor U27697 (N_27697,N_26244,N_26161);
and U27698 (N_27698,N_26226,N_26964);
nand U27699 (N_27699,N_26571,N_26895);
and U27700 (N_27700,N_26738,N_26637);
nand U27701 (N_27701,N_26468,N_26663);
nand U27702 (N_27702,N_26695,N_26588);
xor U27703 (N_27703,N_26154,N_26664);
nand U27704 (N_27704,N_26997,N_26512);
and U27705 (N_27705,N_26710,N_26991);
and U27706 (N_27706,N_26457,N_26001);
nand U27707 (N_27707,N_26186,N_26137);
nor U27708 (N_27708,N_26385,N_26791);
nor U27709 (N_27709,N_26291,N_26566);
or U27710 (N_27710,N_26531,N_26785);
nor U27711 (N_27711,N_26703,N_26878);
xnor U27712 (N_27712,N_26950,N_26804);
nand U27713 (N_27713,N_26936,N_26049);
and U27714 (N_27714,N_26958,N_26443);
or U27715 (N_27715,N_26180,N_26138);
and U27716 (N_27716,N_26825,N_26240);
xor U27717 (N_27717,N_26988,N_26162);
nand U27718 (N_27718,N_26102,N_26777);
nand U27719 (N_27719,N_26365,N_26278);
and U27720 (N_27720,N_26462,N_26275);
nand U27721 (N_27721,N_26800,N_26363);
or U27722 (N_27722,N_26655,N_26354);
nand U27723 (N_27723,N_26079,N_26668);
and U27724 (N_27724,N_26875,N_26052);
or U27725 (N_27725,N_26144,N_26321);
and U27726 (N_27726,N_26555,N_26970);
or U27727 (N_27727,N_26298,N_26048);
and U27728 (N_27728,N_26188,N_26643);
and U27729 (N_27729,N_26514,N_26265);
nor U27730 (N_27730,N_26630,N_26822);
nor U27731 (N_27731,N_26477,N_26961);
nor U27732 (N_27732,N_26964,N_26675);
nand U27733 (N_27733,N_26972,N_26920);
xnor U27734 (N_27734,N_26455,N_26181);
and U27735 (N_27735,N_26561,N_26772);
or U27736 (N_27736,N_26637,N_26547);
or U27737 (N_27737,N_26084,N_26252);
or U27738 (N_27738,N_26397,N_26178);
and U27739 (N_27739,N_26899,N_26222);
xor U27740 (N_27740,N_26289,N_26711);
or U27741 (N_27741,N_26576,N_26286);
or U27742 (N_27742,N_26372,N_26222);
nor U27743 (N_27743,N_26112,N_26674);
xnor U27744 (N_27744,N_26697,N_26082);
nor U27745 (N_27745,N_26994,N_26086);
and U27746 (N_27746,N_26870,N_26382);
xnor U27747 (N_27747,N_26503,N_26433);
nor U27748 (N_27748,N_26398,N_26518);
or U27749 (N_27749,N_26543,N_26184);
or U27750 (N_27750,N_26990,N_26463);
or U27751 (N_27751,N_26376,N_26665);
nand U27752 (N_27752,N_26347,N_26062);
nand U27753 (N_27753,N_26300,N_26859);
nand U27754 (N_27754,N_26520,N_26240);
nor U27755 (N_27755,N_26299,N_26282);
and U27756 (N_27756,N_26719,N_26398);
nand U27757 (N_27757,N_26768,N_26266);
nand U27758 (N_27758,N_26831,N_26216);
and U27759 (N_27759,N_26982,N_26726);
nand U27760 (N_27760,N_26534,N_26037);
nand U27761 (N_27761,N_26685,N_26268);
and U27762 (N_27762,N_26038,N_26415);
nand U27763 (N_27763,N_26680,N_26303);
xnor U27764 (N_27764,N_26233,N_26083);
xor U27765 (N_27765,N_26524,N_26516);
or U27766 (N_27766,N_26138,N_26991);
xor U27767 (N_27767,N_26343,N_26924);
nor U27768 (N_27768,N_26933,N_26501);
nand U27769 (N_27769,N_26557,N_26871);
or U27770 (N_27770,N_26124,N_26495);
xor U27771 (N_27771,N_26729,N_26050);
and U27772 (N_27772,N_26172,N_26484);
and U27773 (N_27773,N_26850,N_26909);
nand U27774 (N_27774,N_26815,N_26112);
or U27775 (N_27775,N_26140,N_26494);
xor U27776 (N_27776,N_26821,N_26883);
nand U27777 (N_27777,N_26106,N_26915);
nor U27778 (N_27778,N_26099,N_26015);
and U27779 (N_27779,N_26330,N_26493);
nand U27780 (N_27780,N_26039,N_26216);
or U27781 (N_27781,N_26344,N_26639);
or U27782 (N_27782,N_26474,N_26624);
nor U27783 (N_27783,N_26184,N_26452);
nand U27784 (N_27784,N_26870,N_26959);
and U27785 (N_27785,N_26747,N_26321);
nand U27786 (N_27786,N_26204,N_26179);
or U27787 (N_27787,N_26391,N_26670);
and U27788 (N_27788,N_26075,N_26053);
nand U27789 (N_27789,N_26440,N_26704);
nor U27790 (N_27790,N_26015,N_26764);
nor U27791 (N_27791,N_26995,N_26433);
or U27792 (N_27792,N_26063,N_26526);
or U27793 (N_27793,N_26395,N_26481);
xor U27794 (N_27794,N_26965,N_26746);
nor U27795 (N_27795,N_26043,N_26146);
and U27796 (N_27796,N_26751,N_26392);
xnor U27797 (N_27797,N_26709,N_26160);
xor U27798 (N_27798,N_26497,N_26140);
xor U27799 (N_27799,N_26010,N_26122);
nand U27800 (N_27800,N_26038,N_26615);
nor U27801 (N_27801,N_26312,N_26549);
and U27802 (N_27802,N_26883,N_26843);
and U27803 (N_27803,N_26192,N_26261);
nand U27804 (N_27804,N_26575,N_26173);
nor U27805 (N_27805,N_26937,N_26687);
and U27806 (N_27806,N_26431,N_26686);
nand U27807 (N_27807,N_26649,N_26762);
nor U27808 (N_27808,N_26724,N_26753);
or U27809 (N_27809,N_26019,N_26160);
nand U27810 (N_27810,N_26523,N_26435);
nor U27811 (N_27811,N_26181,N_26920);
nor U27812 (N_27812,N_26732,N_26060);
and U27813 (N_27813,N_26099,N_26213);
and U27814 (N_27814,N_26901,N_26270);
xor U27815 (N_27815,N_26144,N_26642);
or U27816 (N_27816,N_26550,N_26466);
or U27817 (N_27817,N_26046,N_26211);
or U27818 (N_27818,N_26156,N_26709);
xor U27819 (N_27819,N_26430,N_26196);
and U27820 (N_27820,N_26512,N_26187);
and U27821 (N_27821,N_26587,N_26314);
and U27822 (N_27822,N_26494,N_26479);
xor U27823 (N_27823,N_26530,N_26602);
and U27824 (N_27824,N_26463,N_26635);
and U27825 (N_27825,N_26061,N_26406);
or U27826 (N_27826,N_26059,N_26076);
and U27827 (N_27827,N_26918,N_26188);
nand U27828 (N_27828,N_26329,N_26823);
nand U27829 (N_27829,N_26896,N_26048);
or U27830 (N_27830,N_26237,N_26398);
and U27831 (N_27831,N_26584,N_26623);
nor U27832 (N_27832,N_26753,N_26570);
nand U27833 (N_27833,N_26058,N_26331);
nor U27834 (N_27834,N_26821,N_26234);
nand U27835 (N_27835,N_26888,N_26020);
xnor U27836 (N_27836,N_26245,N_26987);
xnor U27837 (N_27837,N_26969,N_26411);
and U27838 (N_27838,N_26320,N_26512);
nand U27839 (N_27839,N_26470,N_26027);
or U27840 (N_27840,N_26916,N_26582);
and U27841 (N_27841,N_26467,N_26676);
nor U27842 (N_27842,N_26071,N_26370);
nand U27843 (N_27843,N_26382,N_26116);
or U27844 (N_27844,N_26011,N_26308);
nand U27845 (N_27845,N_26227,N_26260);
nor U27846 (N_27846,N_26571,N_26172);
or U27847 (N_27847,N_26424,N_26290);
xnor U27848 (N_27848,N_26944,N_26709);
nor U27849 (N_27849,N_26823,N_26119);
nor U27850 (N_27850,N_26379,N_26898);
and U27851 (N_27851,N_26557,N_26708);
nor U27852 (N_27852,N_26175,N_26056);
xor U27853 (N_27853,N_26512,N_26553);
xnor U27854 (N_27854,N_26920,N_26949);
or U27855 (N_27855,N_26455,N_26651);
xnor U27856 (N_27856,N_26545,N_26103);
nand U27857 (N_27857,N_26886,N_26326);
or U27858 (N_27858,N_26789,N_26180);
nor U27859 (N_27859,N_26482,N_26764);
and U27860 (N_27860,N_26192,N_26421);
and U27861 (N_27861,N_26555,N_26453);
and U27862 (N_27862,N_26279,N_26273);
and U27863 (N_27863,N_26559,N_26847);
nor U27864 (N_27864,N_26382,N_26472);
nor U27865 (N_27865,N_26926,N_26060);
nand U27866 (N_27866,N_26030,N_26494);
nor U27867 (N_27867,N_26709,N_26793);
xnor U27868 (N_27868,N_26055,N_26067);
nand U27869 (N_27869,N_26740,N_26823);
xor U27870 (N_27870,N_26279,N_26448);
nor U27871 (N_27871,N_26069,N_26547);
and U27872 (N_27872,N_26616,N_26020);
xor U27873 (N_27873,N_26446,N_26714);
nor U27874 (N_27874,N_26782,N_26416);
nand U27875 (N_27875,N_26873,N_26745);
or U27876 (N_27876,N_26974,N_26300);
nor U27877 (N_27877,N_26641,N_26342);
xor U27878 (N_27878,N_26714,N_26382);
nand U27879 (N_27879,N_26150,N_26245);
nor U27880 (N_27880,N_26683,N_26513);
xnor U27881 (N_27881,N_26350,N_26103);
xnor U27882 (N_27882,N_26816,N_26736);
and U27883 (N_27883,N_26164,N_26384);
xor U27884 (N_27884,N_26389,N_26337);
xnor U27885 (N_27885,N_26540,N_26851);
or U27886 (N_27886,N_26101,N_26645);
nor U27887 (N_27887,N_26949,N_26469);
and U27888 (N_27888,N_26363,N_26199);
or U27889 (N_27889,N_26610,N_26679);
nand U27890 (N_27890,N_26666,N_26331);
or U27891 (N_27891,N_26875,N_26222);
xor U27892 (N_27892,N_26862,N_26121);
nor U27893 (N_27893,N_26475,N_26368);
or U27894 (N_27894,N_26222,N_26030);
nand U27895 (N_27895,N_26914,N_26325);
and U27896 (N_27896,N_26710,N_26677);
nand U27897 (N_27897,N_26334,N_26426);
nor U27898 (N_27898,N_26143,N_26718);
nand U27899 (N_27899,N_26686,N_26538);
xor U27900 (N_27900,N_26731,N_26318);
nand U27901 (N_27901,N_26857,N_26490);
nor U27902 (N_27902,N_26005,N_26125);
and U27903 (N_27903,N_26065,N_26145);
or U27904 (N_27904,N_26230,N_26350);
nor U27905 (N_27905,N_26892,N_26392);
or U27906 (N_27906,N_26791,N_26877);
xor U27907 (N_27907,N_26297,N_26839);
or U27908 (N_27908,N_26081,N_26774);
nor U27909 (N_27909,N_26741,N_26176);
and U27910 (N_27910,N_26527,N_26413);
nor U27911 (N_27911,N_26140,N_26079);
xor U27912 (N_27912,N_26775,N_26653);
or U27913 (N_27913,N_26392,N_26571);
and U27914 (N_27914,N_26190,N_26503);
xor U27915 (N_27915,N_26827,N_26387);
nand U27916 (N_27916,N_26001,N_26232);
and U27917 (N_27917,N_26005,N_26317);
nand U27918 (N_27918,N_26546,N_26889);
xor U27919 (N_27919,N_26567,N_26193);
and U27920 (N_27920,N_26956,N_26387);
xor U27921 (N_27921,N_26883,N_26849);
or U27922 (N_27922,N_26616,N_26867);
or U27923 (N_27923,N_26420,N_26244);
nor U27924 (N_27924,N_26159,N_26121);
nand U27925 (N_27925,N_26217,N_26894);
xor U27926 (N_27926,N_26025,N_26406);
and U27927 (N_27927,N_26047,N_26936);
and U27928 (N_27928,N_26574,N_26885);
nor U27929 (N_27929,N_26206,N_26221);
or U27930 (N_27930,N_26513,N_26537);
nor U27931 (N_27931,N_26482,N_26142);
nor U27932 (N_27932,N_26289,N_26874);
nor U27933 (N_27933,N_26367,N_26120);
and U27934 (N_27934,N_26778,N_26535);
nand U27935 (N_27935,N_26772,N_26009);
nor U27936 (N_27936,N_26312,N_26366);
xnor U27937 (N_27937,N_26481,N_26192);
xor U27938 (N_27938,N_26175,N_26019);
nor U27939 (N_27939,N_26639,N_26965);
nor U27940 (N_27940,N_26421,N_26989);
and U27941 (N_27941,N_26451,N_26328);
nand U27942 (N_27942,N_26916,N_26170);
xor U27943 (N_27943,N_26613,N_26016);
nand U27944 (N_27944,N_26478,N_26649);
nor U27945 (N_27945,N_26339,N_26809);
nor U27946 (N_27946,N_26468,N_26987);
xor U27947 (N_27947,N_26418,N_26763);
nand U27948 (N_27948,N_26141,N_26985);
xor U27949 (N_27949,N_26824,N_26016);
or U27950 (N_27950,N_26656,N_26486);
and U27951 (N_27951,N_26012,N_26458);
nor U27952 (N_27952,N_26313,N_26103);
nand U27953 (N_27953,N_26290,N_26423);
nand U27954 (N_27954,N_26960,N_26072);
or U27955 (N_27955,N_26167,N_26872);
nor U27956 (N_27956,N_26234,N_26547);
xnor U27957 (N_27957,N_26452,N_26494);
or U27958 (N_27958,N_26802,N_26255);
nand U27959 (N_27959,N_26108,N_26951);
or U27960 (N_27960,N_26557,N_26191);
xor U27961 (N_27961,N_26399,N_26773);
or U27962 (N_27962,N_26445,N_26068);
and U27963 (N_27963,N_26215,N_26375);
nor U27964 (N_27964,N_26690,N_26678);
nand U27965 (N_27965,N_26534,N_26507);
xor U27966 (N_27966,N_26327,N_26752);
xor U27967 (N_27967,N_26181,N_26658);
nor U27968 (N_27968,N_26176,N_26861);
or U27969 (N_27969,N_26368,N_26343);
xnor U27970 (N_27970,N_26519,N_26491);
and U27971 (N_27971,N_26147,N_26505);
nor U27972 (N_27972,N_26987,N_26455);
and U27973 (N_27973,N_26785,N_26696);
nand U27974 (N_27974,N_26247,N_26372);
xor U27975 (N_27975,N_26189,N_26623);
xnor U27976 (N_27976,N_26228,N_26267);
and U27977 (N_27977,N_26521,N_26664);
and U27978 (N_27978,N_26152,N_26573);
or U27979 (N_27979,N_26073,N_26178);
nand U27980 (N_27980,N_26651,N_26152);
xor U27981 (N_27981,N_26475,N_26494);
or U27982 (N_27982,N_26258,N_26780);
or U27983 (N_27983,N_26027,N_26920);
nor U27984 (N_27984,N_26613,N_26511);
and U27985 (N_27985,N_26249,N_26717);
nand U27986 (N_27986,N_26682,N_26818);
nor U27987 (N_27987,N_26110,N_26406);
nand U27988 (N_27988,N_26862,N_26585);
xnor U27989 (N_27989,N_26748,N_26538);
and U27990 (N_27990,N_26005,N_26990);
and U27991 (N_27991,N_26106,N_26836);
xnor U27992 (N_27992,N_26704,N_26899);
nor U27993 (N_27993,N_26286,N_26361);
and U27994 (N_27994,N_26032,N_26076);
nor U27995 (N_27995,N_26489,N_26857);
nor U27996 (N_27996,N_26801,N_26349);
or U27997 (N_27997,N_26646,N_26814);
xor U27998 (N_27998,N_26545,N_26285);
xnor U27999 (N_27999,N_26655,N_26933);
nand U28000 (N_28000,N_27589,N_27458);
nor U28001 (N_28001,N_27764,N_27260);
xnor U28002 (N_28002,N_27138,N_27600);
nor U28003 (N_28003,N_27960,N_27920);
nand U28004 (N_28004,N_27951,N_27567);
xnor U28005 (N_28005,N_27505,N_27916);
and U28006 (N_28006,N_27998,N_27294);
nor U28007 (N_28007,N_27148,N_27161);
or U28008 (N_28008,N_27980,N_27799);
or U28009 (N_28009,N_27947,N_27500);
or U28010 (N_28010,N_27970,N_27773);
or U28011 (N_28011,N_27893,N_27251);
nor U28012 (N_28012,N_27852,N_27489);
xnor U28013 (N_28013,N_27042,N_27413);
or U28014 (N_28014,N_27918,N_27605);
or U28015 (N_28015,N_27724,N_27023);
nand U28016 (N_28016,N_27757,N_27243);
nand U28017 (N_28017,N_27551,N_27792);
and U28018 (N_28018,N_27134,N_27327);
nor U28019 (N_28019,N_27795,N_27174);
nand U28020 (N_28020,N_27924,N_27295);
nand U28021 (N_28021,N_27865,N_27173);
nor U28022 (N_28022,N_27300,N_27798);
nor U28023 (N_28023,N_27695,N_27412);
and U28024 (N_28024,N_27350,N_27742);
and U28025 (N_28025,N_27287,N_27190);
nand U28026 (N_28026,N_27302,N_27217);
nor U28027 (N_28027,N_27168,N_27126);
nor U28028 (N_28028,N_27741,N_27603);
and U28029 (N_28029,N_27650,N_27649);
xor U28030 (N_28030,N_27698,N_27209);
and U28031 (N_28031,N_27283,N_27663);
or U28032 (N_28032,N_27112,N_27717);
or U28033 (N_28033,N_27523,N_27891);
xor U28034 (N_28034,N_27405,N_27305);
or U28035 (N_28035,N_27364,N_27638);
nand U28036 (N_28036,N_27468,N_27047);
or U28037 (N_28037,N_27384,N_27766);
or U28038 (N_28038,N_27417,N_27936);
xor U28039 (N_28039,N_27729,N_27850);
or U28040 (N_28040,N_27493,N_27485);
and U28041 (N_28041,N_27457,N_27187);
and U28042 (N_28042,N_27012,N_27574);
xnor U28043 (N_28043,N_27533,N_27314);
nand U28044 (N_28044,N_27946,N_27169);
and U28045 (N_28045,N_27027,N_27402);
or U28046 (N_28046,N_27986,N_27699);
and U28047 (N_28047,N_27044,N_27312);
or U28048 (N_28048,N_27552,N_27255);
nand U28049 (N_28049,N_27398,N_27547);
xor U28050 (N_28050,N_27376,N_27703);
nand U28051 (N_28051,N_27064,N_27240);
nor U28052 (N_28052,N_27440,N_27181);
and U28053 (N_28053,N_27677,N_27661);
nand U28054 (N_28054,N_27572,N_27232);
and U28055 (N_28055,N_27108,N_27634);
or U28056 (N_28056,N_27281,N_27514);
nand U28057 (N_28057,N_27751,N_27336);
xnor U28058 (N_28058,N_27212,N_27874);
nand U28059 (N_28059,N_27392,N_27414);
xnor U28060 (N_28060,N_27411,N_27261);
and U28061 (N_28061,N_27151,N_27651);
and U28062 (N_28062,N_27944,N_27241);
nor U28063 (N_28063,N_27107,N_27637);
and U28064 (N_28064,N_27885,N_27901);
and U28065 (N_28065,N_27563,N_27501);
nand U28066 (N_28066,N_27859,N_27539);
or U28067 (N_28067,N_27301,N_27610);
nor U28068 (N_28068,N_27668,N_27396);
xnor U28069 (N_28069,N_27085,N_27284);
or U28070 (N_28070,N_27842,N_27180);
nand U28071 (N_28071,N_27525,N_27503);
and U28072 (N_28072,N_27915,N_27821);
or U28073 (N_28073,N_27824,N_27297);
and U28074 (N_28074,N_27498,N_27774);
nor U28075 (N_28075,N_27534,N_27571);
and U28076 (N_28076,N_27016,N_27565);
xor U28077 (N_28077,N_27092,N_27478);
nand U28078 (N_28078,N_27671,N_27646);
nand U28079 (N_28079,N_27471,N_27976);
or U28080 (N_28080,N_27438,N_27965);
or U28081 (N_28081,N_27387,N_27278);
nand U28082 (N_28082,N_27189,N_27611);
xnor U28083 (N_28083,N_27706,N_27822);
nand U28084 (N_28084,N_27954,N_27644);
nor U28085 (N_28085,N_27046,N_27755);
nor U28086 (N_28086,N_27199,N_27556);
or U28087 (N_28087,N_27608,N_27761);
xor U28088 (N_28088,N_27121,N_27455);
xnor U28089 (N_28089,N_27059,N_27338);
or U28090 (N_28090,N_27910,N_27216);
xnor U28091 (N_28091,N_27194,N_27829);
xor U28092 (N_28092,N_27914,N_27504);
and U28093 (N_28093,N_27242,N_27329);
or U28094 (N_28094,N_27862,N_27367);
nor U28095 (N_28095,N_27456,N_27246);
nand U28096 (N_28096,N_27612,N_27927);
xor U28097 (N_28097,N_27239,N_27790);
or U28098 (N_28098,N_27981,N_27334);
or U28099 (N_28099,N_27351,N_27801);
nor U28100 (N_28100,N_27102,N_27021);
nand U28101 (N_28101,N_27379,N_27667);
nand U28102 (N_28102,N_27632,N_27013);
nor U28103 (N_28103,N_27544,N_27035);
and U28104 (N_28104,N_27690,N_27073);
xnor U28105 (N_28105,N_27256,N_27921);
and U28106 (N_28106,N_27075,N_27687);
nand U28107 (N_28107,N_27160,N_27867);
nor U28108 (N_28108,N_27911,N_27834);
or U28109 (N_28109,N_27250,N_27111);
nand U28110 (N_28110,N_27718,N_27346);
xor U28111 (N_28111,N_27487,N_27306);
nand U28112 (N_28112,N_27847,N_27840);
or U28113 (N_28113,N_27835,N_27601);
and U28114 (N_28114,N_27065,N_27370);
nand U28115 (N_28115,N_27641,N_27648);
nor U28116 (N_28116,N_27783,N_27486);
nor U28117 (N_28117,N_27701,N_27923);
and U28118 (N_28118,N_27756,N_27165);
nand U28119 (N_28119,N_27584,N_27995);
nand U28120 (N_28120,N_27769,N_27454);
nor U28121 (N_28121,N_27557,N_27818);
nor U28122 (N_28122,N_27462,N_27139);
xor U28123 (N_28123,N_27709,N_27322);
or U28124 (N_28124,N_27545,N_27389);
nand U28125 (N_28125,N_27495,N_27538);
nor U28126 (N_28126,N_27985,N_27407);
nand U28127 (N_28127,N_27938,N_27259);
or U28128 (N_28128,N_27307,N_27749);
nand U28129 (N_28129,N_27873,N_27760);
or U28130 (N_28130,N_27437,N_27031);
nor U28131 (N_28131,N_27685,N_27594);
nand U28132 (N_28132,N_27056,N_27592);
and U28133 (N_28133,N_27647,N_27153);
xnor U28134 (N_28134,N_27721,N_27740);
and U28135 (N_28135,N_27465,N_27894);
xor U28136 (N_28136,N_27812,N_27087);
and U28137 (N_28137,N_27786,N_27427);
nor U28138 (N_28138,N_27908,N_27028);
nor U28139 (N_28139,N_27282,N_27103);
or U28140 (N_28140,N_27024,N_27096);
or U28141 (N_28141,N_27508,N_27142);
and U28142 (N_28142,N_27130,N_27953);
or U28143 (N_28143,N_27735,N_27811);
nand U28144 (N_28144,N_27521,N_27436);
nand U28145 (N_28145,N_27658,N_27040);
nor U28146 (N_28146,N_27733,N_27330);
and U28147 (N_28147,N_27030,N_27320);
nand U28148 (N_28148,N_27186,N_27763);
nand U28149 (N_28149,N_27967,N_27039);
xor U28150 (N_28150,N_27206,N_27091);
and U28151 (N_28151,N_27994,N_27155);
xor U28152 (N_28152,N_27432,N_27288);
or U28153 (N_28153,N_27404,N_27378);
nand U28154 (N_28154,N_27990,N_27123);
xor U28155 (N_28155,N_27555,N_27984);
xnor U28156 (N_28156,N_27079,N_27449);
xor U28157 (N_28157,N_27089,N_27313);
nand U28158 (N_28158,N_27484,N_27248);
or U28159 (N_28159,N_27453,N_27948);
nand U28160 (N_28160,N_27502,N_27715);
nor U28161 (N_28161,N_27009,N_27443);
xor U28162 (N_28162,N_27005,N_27060);
xnor U28163 (N_28163,N_27309,N_27977);
nand U28164 (N_28164,N_27779,N_27140);
nand U28165 (N_28165,N_27499,N_27808);
or U28166 (N_28166,N_27176,N_27268);
nand U28167 (N_28167,N_27827,N_27767);
nand U28168 (N_28168,N_27682,N_27115);
nand U28169 (N_28169,N_27746,N_27974);
nand U28170 (N_28170,N_27917,N_27395);
nand U28171 (N_28171,N_27418,N_27365);
or U28172 (N_28172,N_27939,N_27122);
nand U28173 (N_28173,N_27654,N_27444);
or U28174 (N_28174,N_27897,N_27930);
nand U28175 (N_28175,N_27050,N_27802);
xor U28176 (N_28176,N_27510,N_27270);
xor U28177 (N_28177,N_27913,N_27477);
and U28178 (N_28178,N_27684,N_27999);
and U28179 (N_28179,N_27895,N_27043);
nor U28180 (N_28180,N_27884,N_27762);
xnor U28181 (N_28181,N_27158,N_27269);
nor U28182 (N_28182,N_27464,N_27643);
nand U28183 (N_28183,N_27640,N_27736);
nor U28184 (N_28184,N_27357,N_27575);
or U28185 (N_28185,N_27394,N_27452);
nand U28186 (N_28186,N_27739,N_27907);
xor U28187 (N_28187,N_27360,N_27274);
nor U28188 (N_28188,N_27955,N_27204);
xnor U28189 (N_28189,N_27467,N_27585);
xnor U28190 (N_28190,N_27292,N_27730);
xor U28191 (N_28191,N_27899,N_27037);
and U28192 (N_28192,N_27445,N_27355);
and U28193 (N_28193,N_27034,N_27618);
xor U28194 (N_28194,N_27135,N_27768);
nand U28195 (N_28195,N_27422,N_27672);
or U28196 (N_28196,N_27120,N_27748);
xnor U28197 (N_28197,N_27258,N_27285);
or U28198 (N_28198,N_27342,N_27473);
and U28199 (N_28199,N_27731,N_27881);
nor U28200 (N_28200,N_27383,N_27590);
or U28201 (N_28201,N_27882,N_27548);
nor U28202 (N_28202,N_27813,N_27286);
nand U28203 (N_28203,N_27922,N_27184);
nor U28204 (N_28204,N_27609,N_27653);
nand U28205 (N_28205,N_27235,N_27293);
and U28206 (N_28206,N_27315,N_27747);
nand U28207 (N_28207,N_27221,N_27424);
nand U28208 (N_28208,N_27400,N_27689);
and U28209 (N_28209,N_27657,N_27639);
and U28210 (N_28210,N_27195,N_27368);
nor U28211 (N_28211,N_27019,N_27596);
nor U28212 (N_28212,N_27833,N_27815);
nand U28213 (N_28213,N_27805,N_27772);
or U28214 (N_28214,N_27220,N_27159);
xor U28215 (N_28215,N_27511,N_27806);
nand U28216 (N_28216,N_27925,N_27428);
nand U28217 (N_28217,N_27616,N_27568);
nor U28218 (N_28218,N_27254,N_27780);
xor U28219 (N_28219,N_27866,N_27226);
nand U28220 (N_28220,N_27849,N_27324);
nand U28221 (N_28221,N_27391,N_27002);
nand U28222 (N_28222,N_27777,N_27014);
or U28223 (N_28223,N_27483,N_27228);
and U28224 (N_28224,N_27045,N_27621);
nand U28225 (N_28225,N_27083,N_27714);
nor U28226 (N_28226,N_27708,N_27333);
nand U28227 (N_28227,N_27758,N_27143);
or U28228 (N_28228,N_27020,N_27519);
nor U28229 (N_28229,N_27996,N_27223);
xor U28230 (N_28230,N_27903,N_27470);
nand U28231 (N_28231,N_27566,N_27507);
xor U28232 (N_28232,N_27201,N_27900);
xor U28233 (N_28233,N_27804,N_27426);
or U28234 (N_28234,N_27406,N_27474);
nand U28235 (N_28235,N_27694,N_27325);
nand U28236 (N_28236,N_27851,N_27561);
nor U28237 (N_28237,N_27854,N_27442);
xor U28238 (N_28238,N_27704,N_27172);
xor U28239 (N_28239,N_27509,N_27666);
nand U28240 (N_28240,N_27431,N_27304);
xor U28241 (N_28241,N_27871,N_27202);
nand U28242 (N_28242,N_27185,N_27257);
or U28243 (N_28243,N_27518,N_27193);
and U28244 (N_28244,N_27993,N_27167);
xor U28245 (N_28245,N_27529,N_27720);
nand U28246 (N_28246,N_27244,N_27110);
nor U28247 (N_28247,N_27385,N_27291);
and U28248 (N_28248,N_27581,N_27318);
or U28249 (N_28249,N_27488,N_27163);
nand U28250 (N_28250,N_27934,N_27554);
nand U28251 (N_28251,N_27249,N_27952);
xnor U28252 (N_28252,N_27613,N_27113);
and U28253 (N_28253,N_27353,N_27224);
nand U28254 (N_28254,N_27247,N_27188);
nor U28255 (N_28255,N_27230,N_27719);
xor U28256 (N_28256,N_27593,N_27789);
nor U28257 (N_28257,N_27054,N_27578);
and U28258 (N_28258,N_27912,N_27415);
or U28259 (N_28259,N_27481,N_27633);
xnor U28260 (N_28260,N_27057,N_27707);
xor U28261 (N_28261,N_27909,N_27652);
nand U28262 (N_28262,N_27550,N_27870);
nand U28263 (N_28263,N_27828,N_27032);
or U28264 (N_28264,N_27067,N_27631);
or U28265 (N_28265,N_27208,N_27071);
or U28266 (N_28266,N_27001,N_27372);
nor U28267 (N_28267,N_27041,N_27506);
nand U28268 (N_28268,N_27328,N_27515);
nand U28269 (N_28269,N_27989,N_27086);
nor U28270 (N_28270,N_27826,N_27157);
or U28271 (N_28271,N_27238,N_27620);
and U28272 (N_28272,N_27095,N_27814);
and U28273 (N_28273,N_27528,N_27408);
or U28274 (N_28274,N_27356,N_27141);
nand U28275 (N_28275,N_27928,N_27145);
nand U28276 (N_28276,N_27683,N_27029);
or U28277 (N_28277,N_27341,N_27058);
xor U28278 (N_28278,N_27000,N_27712);
xor U28279 (N_28279,N_27615,N_27642);
and U28280 (N_28280,N_27662,N_27132);
or U28281 (N_28281,N_27425,N_27179);
nor U28282 (N_28282,N_27214,N_27344);
or U28283 (N_28283,N_27697,N_27627);
xor U28284 (N_28284,N_27373,N_27591);
nand U28285 (N_28285,N_27359,N_27210);
nand U28286 (N_28286,N_27080,N_27800);
nand U28287 (N_28287,N_27997,N_27540);
or U28288 (N_28288,N_27880,N_27599);
or U28289 (N_28289,N_27765,N_27461);
and U28290 (N_28290,N_27737,N_27987);
xnor U28291 (N_28291,N_27945,N_27949);
nor U28292 (N_28292,N_27573,N_27705);
nor U28293 (N_28293,N_27175,N_27101);
or U28294 (N_28294,N_27265,N_27883);
xnor U28295 (N_28295,N_27723,N_27038);
xor U28296 (N_28296,N_27119,N_27797);
and U28297 (N_28297,N_27010,N_27093);
and U28298 (N_28298,N_27429,N_27303);
xnor U28299 (N_28299,N_27482,N_27597);
nor U28300 (N_28300,N_27381,N_27553);
nor U28301 (N_28301,N_27491,N_27441);
and U28302 (N_28302,N_27595,N_27878);
nor U28303 (N_28303,N_27535,N_27656);
nand U28304 (N_28304,N_27154,N_27586);
xnor U28305 (N_28305,N_27962,N_27966);
nand U28306 (N_28306,N_27207,N_27886);
nand U28307 (N_28307,N_27319,N_27670);
and U28308 (N_28308,N_27331,N_27564);
and U28309 (N_28309,N_27033,N_27604);
nor U28310 (N_28310,N_27036,N_27524);
nand U28311 (N_28311,N_27371,N_27754);
and U28312 (N_28312,N_27879,N_27479);
nor U28313 (N_28313,N_27317,N_27968);
or U28314 (N_28314,N_27361,N_27655);
nor U28315 (N_28315,N_27109,N_27088);
nand U28316 (N_28316,N_27512,N_27008);
and U28317 (N_28317,N_27077,N_27401);
xor U28318 (N_28318,N_27469,N_27776);
xor U28319 (N_28319,N_27926,N_27337);
and U28320 (N_28320,N_27399,N_27843);
and U28321 (N_28321,N_27678,N_27419);
and U28322 (N_28322,N_27062,N_27669);
nand U28323 (N_28323,N_27097,N_27074);
or U28324 (N_28324,N_27963,N_27352);
nand U28325 (N_28325,N_27081,N_27375);
and U28326 (N_28326,N_27098,N_27864);
or U28327 (N_28327,N_27770,N_27832);
and U28328 (N_28328,N_27700,N_27298);
nor U28329 (N_28329,N_27078,N_27788);
nand U28330 (N_28330,N_27076,N_27680);
xnor U28331 (N_28331,N_27796,N_27973);
nand U28332 (N_28332,N_27090,N_27558);
and U28333 (N_28333,N_27343,N_27490);
or U28334 (N_28334,N_27841,N_27084);
or U28335 (N_28335,N_27131,N_27825);
nor U28336 (N_28336,N_27875,N_27562);
or U28337 (N_28337,N_27816,N_27860);
or U28338 (N_28338,N_27846,N_27940);
nor U28339 (N_28339,N_27340,N_27803);
and U28340 (N_28340,N_27716,N_27136);
nor U28341 (N_28341,N_27403,N_27252);
or U28342 (N_28342,N_27211,N_27171);
nor U28343 (N_28343,N_27710,N_27681);
or U28344 (N_28344,N_27626,N_27975);
xor U28345 (N_28345,N_27602,N_27645);
nor U28346 (N_28346,N_27527,N_27686);
nor U28347 (N_28347,N_27466,N_27117);
or U28348 (N_28348,N_27991,N_27299);
or U28349 (N_28349,N_27791,N_27820);
or U28350 (N_28350,N_27614,N_27289);
and U28351 (N_28351,N_27377,N_27728);
nand U28352 (N_28352,N_27137,N_27225);
nor U28353 (N_28353,N_27711,N_27051);
nor U28354 (N_28354,N_27146,N_27410);
nand U28355 (N_28355,N_27857,N_27280);
nand U28356 (N_28356,N_27517,N_27713);
nor U28357 (N_28357,N_27362,N_27177);
nand U28358 (N_28358,N_27856,N_27972);
or U28359 (N_28359,N_27837,N_27950);
nor U28360 (N_28360,N_27889,N_27676);
nand U28361 (N_28361,N_27162,N_27659);
or U28362 (N_28362,N_27197,N_27892);
nor U28363 (N_28363,N_27339,N_27941);
and U28364 (N_28364,N_27476,N_27771);
nor U28365 (N_28365,N_27018,N_27082);
and U28366 (N_28366,N_27480,N_27855);
nor U28367 (N_28367,N_27127,N_27099);
nor U28368 (N_28368,N_27198,N_27752);
and U28369 (N_28369,N_27863,N_27560);
xnor U28370 (N_28370,N_27026,N_27022);
nor U28371 (N_28371,N_27205,N_27118);
or U28372 (N_28372,N_27147,N_27277);
xor U28373 (N_28373,N_27872,N_27233);
nand U28374 (N_28374,N_27133,N_27861);
and U28375 (N_28375,N_27170,N_27290);
or U28376 (N_28376,N_27830,N_27906);
and U28377 (N_28377,N_27055,N_27494);
and U28378 (N_28378,N_27348,N_27725);
and U28379 (N_28379,N_27619,N_27932);
nand U28380 (N_28380,N_27902,N_27231);
xor U28381 (N_28381,N_27049,N_27702);
or U28382 (N_28382,N_27809,N_27957);
nor U28383 (N_28383,N_27192,N_27459);
xnor U28384 (N_28384,N_27964,N_27434);
nor U28385 (N_28385,N_27156,N_27530);
nand U28386 (N_28386,N_27382,N_27890);
xor U28387 (N_28387,N_27347,N_27810);
and U28388 (N_28388,N_27450,N_27848);
nor U28389 (N_28389,N_27166,N_27366);
and U28390 (N_28390,N_27905,N_27775);
xnor U28391 (N_28391,N_27386,N_27679);
nor U28392 (N_28392,N_27688,N_27660);
nand U28393 (N_28393,N_27858,N_27817);
or U28394 (N_28394,N_27665,N_27275);
and U28395 (N_28395,N_27549,N_27520);
and U28396 (N_28396,N_27983,N_27296);
or U28397 (N_28397,N_27262,N_27513);
nand U28398 (N_28398,N_27496,N_27420);
and U28399 (N_28399,N_27937,N_27237);
nand U28400 (N_28400,N_27349,N_27526);
and U28401 (N_28401,N_27635,N_27577);
and U28402 (N_28402,N_27838,N_27622);
xnor U28403 (N_28403,N_27819,N_27006);
and U28404 (N_28404,N_27069,N_27272);
and U28405 (N_28405,N_27354,N_27380);
or U28406 (N_28406,N_27446,N_27178);
or U28407 (N_28407,N_27053,N_27007);
nor U28408 (N_28408,N_27839,N_27439);
or U28409 (N_28409,N_27421,N_27273);
nand U28410 (N_28410,N_27017,N_27793);
nor U28411 (N_28411,N_27784,N_27219);
or U28412 (N_28412,N_27100,N_27070);
or U28413 (N_28413,N_27978,N_27061);
nand U28414 (N_28414,N_27311,N_27222);
nor U28415 (N_28415,N_27321,N_27266);
nand U28416 (N_28416,N_27738,N_27323);
or U28417 (N_28417,N_27435,N_27781);
nand U28418 (N_28418,N_27674,N_27807);
nor U28419 (N_28419,N_27904,N_27125);
nor U28420 (N_28420,N_27196,N_27877);
and U28421 (N_28421,N_27416,N_27271);
nor U28422 (N_28422,N_27782,N_27072);
nand U28423 (N_28423,N_27588,N_27750);
nand U28424 (N_28424,N_27451,N_27543);
or U28425 (N_28425,N_27433,N_27144);
and U28426 (N_28426,N_27869,N_27263);
nor U28427 (N_28427,N_27958,N_27183);
nand U28428 (N_28428,N_27245,N_27388);
nor U28429 (N_28429,N_27492,N_27692);
nand U28430 (N_28430,N_27310,N_27823);
or U28431 (N_28431,N_27625,N_27358);
and U28432 (N_28432,N_27460,N_27004);
xnor U28433 (N_28433,N_27606,N_27229);
nor U28434 (N_28434,N_27743,N_27393);
nor U28435 (N_28435,N_27345,N_27582);
xor U28436 (N_28436,N_27559,N_27536);
nand U28437 (N_28437,N_27576,N_27979);
nand U28438 (N_28438,N_27264,N_27066);
nor U28439 (N_28439,N_27011,N_27215);
nand U28440 (N_28440,N_27935,N_27068);
and U28441 (N_28441,N_27150,N_27898);
xnor U28442 (N_28442,N_27579,N_27583);
or U28443 (N_28443,N_27693,N_27623);
nand U28444 (N_28444,N_27475,N_27629);
and U28445 (N_28445,N_27607,N_27931);
xor U28446 (N_28446,N_27374,N_27844);
and U28447 (N_28447,N_27956,N_27390);
nand U28448 (N_28448,N_27048,N_27203);
or U28449 (N_28449,N_27363,N_27279);
xnor U28450 (N_28450,N_27580,N_27430);
nand U28451 (N_28451,N_27876,N_27015);
or U28452 (N_28452,N_27003,N_27624);
nand U28453 (N_28453,N_27691,N_27369);
xor U28454 (N_28454,N_27942,N_27152);
and U28455 (N_28455,N_27753,N_27542);
nor U28456 (N_28456,N_27149,N_27182);
xnor U28457 (N_28457,N_27308,N_27778);
nor U28458 (N_28458,N_27234,N_27546);
nand U28459 (N_28459,N_27933,N_27845);
and U28460 (N_28460,N_27025,N_27887);
and U28461 (N_28461,N_27531,N_27675);
and U28462 (N_28462,N_27497,N_27191);
nand U28463 (N_28463,N_27094,N_27969);
and U28464 (N_28464,N_27063,N_27116);
xor U28465 (N_28465,N_27734,N_27276);
nand U28466 (N_28466,N_27732,N_27052);
nor U28467 (N_28467,N_27569,N_27124);
xnor U28468 (N_28468,N_27253,N_27617);
or U28469 (N_28469,N_27868,N_27472);
nor U28470 (N_28470,N_27522,N_27745);
and U28471 (N_28471,N_27129,N_27447);
nand U28472 (N_28472,N_27516,N_27722);
and U28473 (N_28473,N_27598,N_27236);
or U28474 (N_28474,N_27896,N_27673);
nand U28475 (N_28475,N_27164,N_27961);
or U28476 (N_28476,N_27988,N_27853);
xor U28477 (N_28477,N_27537,N_27726);
nand U28478 (N_28478,N_27696,N_27335);
nand U28479 (N_28479,N_27943,N_27794);
and U28480 (N_28480,N_27759,N_27929);
or U28481 (N_28481,N_27332,N_27200);
xnor U28482 (N_28482,N_27836,N_27727);
or U28483 (N_28483,N_27664,N_27831);
nor U28484 (N_28484,N_27213,N_27218);
and U28485 (N_28485,N_27463,N_27971);
nand U28486 (N_28486,N_27628,N_27744);
or U28487 (N_28487,N_27541,N_27397);
or U28488 (N_28488,N_27423,N_27636);
or U28489 (N_28489,N_27787,N_27992);
nor U28490 (N_28490,N_27959,N_27114);
nand U28491 (N_28491,N_27982,N_27326);
nand U28492 (N_28492,N_27919,N_27267);
xor U28493 (N_28493,N_27532,N_27570);
and U28494 (N_28494,N_27785,N_27587);
xor U28495 (N_28495,N_27888,N_27105);
xnor U28496 (N_28496,N_27227,N_27104);
nand U28497 (N_28497,N_27448,N_27128);
and U28498 (N_28498,N_27316,N_27106);
nand U28499 (N_28499,N_27630,N_27409);
nor U28500 (N_28500,N_27942,N_27022);
and U28501 (N_28501,N_27153,N_27526);
and U28502 (N_28502,N_27644,N_27171);
nor U28503 (N_28503,N_27710,N_27984);
nand U28504 (N_28504,N_27903,N_27906);
and U28505 (N_28505,N_27637,N_27101);
nand U28506 (N_28506,N_27283,N_27622);
and U28507 (N_28507,N_27826,N_27851);
or U28508 (N_28508,N_27331,N_27279);
and U28509 (N_28509,N_27998,N_27584);
nand U28510 (N_28510,N_27216,N_27906);
and U28511 (N_28511,N_27926,N_27300);
xnor U28512 (N_28512,N_27129,N_27837);
nor U28513 (N_28513,N_27409,N_27294);
nand U28514 (N_28514,N_27809,N_27681);
xnor U28515 (N_28515,N_27390,N_27100);
and U28516 (N_28516,N_27582,N_27073);
and U28517 (N_28517,N_27052,N_27035);
and U28518 (N_28518,N_27232,N_27358);
xnor U28519 (N_28519,N_27406,N_27113);
and U28520 (N_28520,N_27199,N_27013);
nor U28521 (N_28521,N_27330,N_27841);
and U28522 (N_28522,N_27297,N_27027);
xnor U28523 (N_28523,N_27932,N_27046);
or U28524 (N_28524,N_27347,N_27157);
xnor U28525 (N_28525,N_27905,N_27754);
and U28526 (N_28526,N_27798,N_27651);
or U28527 (N_28527,N_27983,N_27066);
xor U28528 (N_28528,N_27722,N_27817);
or U28529 (N_28529,N_27878,N_27729);
nand U28530 (N_28530,N_27948,N_27024);
xnor U28531 (N_28531,N_27993,N_27761);
and U28532 (N_28532,N_27585,N_27160);
nand U28533 (N_28533,N_27051,N_27492);
or U28534 (N_28534,N_27623,N_27026);
and U28535 (N_28535,N_27585,N_27440);
nand U28536 (N_28536,N_27914,N_27848);
and U28537 (N_28537,N_27275,N_27246);
and U28538 (N_28538,N_27173,N_27819);
and U28539 (N_28539,N_27734,N_27967);
and U28540 (N_28540,N_27035,N_27582);
or U28541 (N_28541,N_27214,N_27167);
or U28542 (N_28542,N_27003,N_27282);
nor U28543 (N_28543,N_27850,N_27357);
or U28544 (N_28544,N_27184,N_27835);
nor U28545 (N_28545,N_27356,N_27393);
or U28546 (N_28546,N_27373,N_27997);
nand U28547 (N_28547,N_27990,N_27646);
nand U28548 (N_28548,N_27208,N_27716);
nand U28549 (N_28549,N_27520,N_27934);
and U28550 (N_28550,N_27031,N_27397);
xnor U28551 (N_28551,N_27472,N_27371);
nand U28552 (N_28552,N_27332,N_27775);
xnor U28553 (N_28553,N_27677,N_27729);
and U28554 (N_28554,N_27974,N_27783);
or U28555 (N_28555,N_27071,N_27556);
or U28556 (N_28556,N_27085,N_27871);
or U28557 (N_28557,N_27535,N_27631);
xor U28558 (N_28558,N_27230,N_27759);
and U28559 (N_28559,N_27661,N_27339);
xnor U28560 (N_28560,N_27155,N_27020);
xnor U28561 (N_28561,N_27544,N_27903);
nand U28562 (N_28562,N_27687,N_27847);
xnor U28563 (N_28563,N_27936,N_27270);
nor U28564 (N_28564,N_27317,N_27236);
and U28565 (N_28565,N_27854,N_27776);
xor U28566 (N_28566,N_27299,N_27629);
nand U28567 (N_28567,N_27658,N_27461);
nand U28568 (N_28568,N_27557,N_27286);
xor U28569 (N_28569,N_27834,N_27385);
or U28570 (N_28570,N_27476,N_27666);
nand U28571 (N_28571,N_27377,N_27168);
nand U28572 (N_28572,N_27210,N_27938);
nand U28573 (N_28573,N_27490,N_27143);
or U28574 (N_28574,N_27411,N_27980);
nand U28575 (N_28575,N_27342,N_27700);
and U28576 (N_28576,N_27310,N_27934);
and U28577 (N_28577,N_27276,N_27292);
and U28578 (N_28578,N_27399,N_27882);
nand U28579 (N_28579,N_27808,N_27874);
or U28580 (N_28580,N_27613,N_27389);
xor U28581 (N_28581,N_27499,N_27221);
nand U28582 (N_28582,N_27401,N_27187);
nor U28583 (N_28583,N_27265,N_27590);
and U28584 (N_28584,N_27297,N_27679);
xor U28585 (N_28585,N_27609,N_27315);
nor U28586 (N_28586,N_27491,N_27192);
or U28587 (N_28587,N_27839,N_27212);
xnor U28588 (N_28588,N_27158,N_27852);
nor U28589 (N_28589,N_27921,N_27169);
xnor U28590 (N_28590,N_27141,N_27361);
xor U28591 (N_28591,N_27566,N_27417);
nand U28592 (N_28592,N_27437,N_27036);
or U28593 (N_28593,N_27960,N_27705);
nor U28594 (N_28594,N_27095,N_27580);
and U28595 (N_28595,N_27217,N_27864);
nand U28596 (N_28596,N_27019,N_27273);
nor U28597 (N_28597,N_27366,N_27680);
nor U28598 (N_28598,N_27806,N_27528);
nor U28599 (N_28599,N_27974,N_27149);
xnor U28600 (N_28600,N_27175,N_27886);
nor U28601 (N_28601,N_27633,N_27771);
nand U28602 (N_28602,N_27927,N_27648);
and U28603 (N_28603,N_27506,N_27156);
xnor U28604 (N_28604,N_27956,N_27802);
nor U28605 (N_28605,N_27915,N_27400);
nand U28606 (N_28606,N_27637,N_27866);
nor U28607 (N_28607,N_27185,N_27357);
nor U28608 (N_28608,N_27787,N_27573);
and U28609 (N_28609,N_27900,N_27393);
or U28610 (N_28610,N_27318,N_27190);
nand U28611 (N_28611,N_27558,N_27218);
xnor U28612 (N_28612,N_27230,N_27677);
and U28613 (N_28613,N_27791,N_27018);
and U28614 (N_28614,N_27933,N_27355);
nand U28615 (N_28615,N_27393,N_27851);
nor U28616 (N_28616,N_27848,N_27650);
nand U28617 (N_28617,N_27696,N_27214);
or U28618 (N_28618,N_27685,N_27077);
xnor U28619 (N_28619,N_27338,N_27307);
xor U28620 (N_28620,N_27888,N_27566);
and U28621 (N_28621,N_27034,N_27954);
and U28622 (N_28622,N_27048,N_27085);
nor U28623 (N_28623,N_27003,N_27968);
and U28624 (N_28624,N_27602,N_27116);
or U28625 (N_28625,N_27903,N_27371);
nor U28626 (N_28626,N_27624,N_27316);
and U28627 (N_28627,N_27786,N_27352);
nand U28628 (N_28628,N_27120,N_27341);
nor U28629 (N_28629,N_27321,N_27588);
or U28630 (N_28630,N_27164,N_27146);
nor U28631 (N_28631,N_27691,N_27961);
xnor U28632 (N_28632,N_27417,N_27524);
and U28633 (N_28633,N_27410,N_27327);
nor U28634 (N_28634,N_27406,N_27567);
or U28635 (N_28635,N_27047,N_27237);
and U28636 (N_28636,N_27853,N_27888);
nor U28637 (N_28637,N_27621,N_27747);
or U28638 (N_28638,N_27218,N_27299);
or U28639 (N_28639,N_27770,N_27689);
and U28640 (N_28640,N_27459,N_27605);
or U28641 (N_28641,N_27625,N_27406);
nand U28642 (N_28642,N_27063,N_27963);
or U28643 (N_28643,N_27212,N_27748);
nor U28644 (N_28644,N_27045,N_27133);
and U28645 (N_28645,N_27389,N_27057);
nor U28646 (N_28646,N_27731,N_27707);
nand U28647 (N_28647,N_27261,N_27235);
nand U28648 (N_28648,N_27210,N_27218);
or U28649 (N_28649,N_27442,N_27758);
and U28650 (N_28650,N_27394,N_27303);
xnor U28651 (N_28651,N_27502,N_27961);
nor U28652 (N_28652,N_27715,N_27615);
xor U28653 (N_28653,N_27103,N_27584);
and U28654 (N_28654,N_27525,N_27394);
nor U28655 (N_28655,N_27059,N_27378);
xnor U28656 (N_28656,N_27505,N_27457);
nor U28657 (N_28657,N_27879,N_27252);
nor U28658 (N_28658,N_27034,N_27486);
xor U28659 (N_28659,N_27805,N_27705);
and U28660 (N_28660,N_27096,N_27962);
nor U28661 (N_28661,N_27944,N_27302);
or U28662 (N_28662,N_27929,N_27343);
and U28663 (N_28663,N_27337,N_27237);
and U28664 (N_28664,N_27128,N_27545);
xor U28665 (N_28665,N_27704,N_27504);
and U28666 (N_28666,N_27730,N_27087);
or U28667 (N_28667,N_27415,N_27899);
nand U28668 (N_28668,N_27622,N_27384);
and U28669 (N_28669,N_27985,N_27726);
and U28670 (N_28670,N_27981,N_27233);
nor U28671 (N_28671,N_27327,N_27827);
or U28672 (N_28672,N_27556,N_27190);
nor U28673 (N_28673,N_27797,N_27952);
nand U28674 (N_28674,N_27913,N_27581);
nor U28675 (N_28675,N_27945,N_27918);
nand U28676 (N_28676,N_27584,N_27094);
nor U28677 (N_28677,N_27192,N_27257);
nand U28678 (N_28678,N_27840,N_27647);
nor U28679 (N_28679,N_27459,N_27760);
xnor U28680 (N_28680,N_27414,N_27479);
or U28681 (N_28681,N_27867,N_27799);
or U28682 (N_28682,N_27455,N_27889);
nor U28683 (N_28683,N_27828,N_27536);
nand U28684 (N_28684,N_27313,N_27688);
and U28685 (N_28685,N_27570,N_27987);
nand U28686 (N_28686,N_27741,N_27116);
and U28687 (N_28687,N_27268,N_27802);
or U28688 (N_28688,N_27209,N_27334);
xnor U28689 (N_28689,N_27932,N_27668);
nor U28690 (N_28690,N_27023,N_27335);
nand U28691 (N_28691,N_27258,N_27549);
and U28692 (N_28692,N_27168,N_27988);
and U28693 (N_28693,N_27805,N_27096);
or U28694 (N_28694,N_27331,N_27434);
xor U28695 (N_28695,N_27899,N_27094);
nor U28696 (N_28696,N_27277,N_27440);
or U28697 (N_28697,N_27838,N_27030);
xor U28698 (N_28698,N_27300,N_27715);
or U28699 (N_28699,N_27347,N_27566);
nand U28700 (N_28700,N_27902,N_27330);
xor U28701 (N_28701,N_27365,N_27424);
xnor U28702 (N_28702,N_27668,N_27841);
or U28703 (N_28703,N_27172,N_27284);
or U28704 (N_28704,N_27125,N_27814);
nor U28705 (N_28705,N_27817,N_27025);
nor U28706 (N_28706,N_27817,N_27608);
nor U28707 (N_28707,N_27904,N_27794);
or U28708 (N_28708,N_27170,N_27273);
nor U28709 (N_28709,N_27401,N_27093);
nand U28710 (N_28710,N_27308,N_27415);
nand U28711 (N_28711,N_27892,N_27593);
xnor U28712 (N_28712,N_27473,N_27974);
nor U28713 (N_28713,N_27774,N_27064);
or U28714 (N_28714,N_27489,N_27586);
nor U28715 (N_28715,N_27586,N_27591);
or U28716 (N_28716,N_27201,N_27502);
xor U28717 (N_28717,N_27882,N_27073);
nand U28718 (N_28718,N_27458,N_27628);
nand U28719 (N_28719,N_27142,N_27358);
nor U28720 (N_28720,N_27342,N_27742);
or U28721 (N_28721,N_27189,N_27473);
nor U28722 (N_28722,N_27091,N_27199);
nor U28723 (N_28723,N_27162,N_27559);
nand U28724 (N_28724,N_27696,N_27435);
and U28725 (N_28725,N_27713,N_27881);
xor U28726 (N_28726,N_27254,N_27748);
nand U28727 (N_28727,N_27137,N_27016);
and U28728 (N_28728,N_27602,N_27661);
and U28729 (N_28729,N_27808,N_27961);
xnor U28730 (N_28730,N_27123,N_27565);
and U28731 (N_28731,N_27223,N_27288);
nor U28732 (N_28732,N_27145,N_27696);
nor U28733 (N_28733,N_27816,N_27946);
and U28734 (N_28734,N_27677,N_27464);
nor U28735 (N_28735,N_27389,N_27908);
nand U28736 (N_28736,N_27985,N_27740);
nand U28737 (N_28737,N_27875,N_27114);
xor U28738 (N_28738,N_27350,N_27009);
or U28739 (N_28739,N_27262,N_27200);
and U28740 (N_28740,N_27167,N_27953);
xor U28741 (N_28741,N_27473,N_27510);
or U28742 (N_28742,N_27460,N_27941);
and U28743 (N_28743,N_27295,N_27495);
xor U28744 (N_28744,N_27397,N_27927);
xnor U28745 (N_28745,N_27795,N_27376);
nand U28746 (N_28746,N_27876,N_27128);
and U28747 (N_28747,N_27510,N_27756);
or U28748 (N_28748,N_27434,N_27059);
xnor U28749 (N_28749,N_27178,N_27714);
and U28750 (N_28750,N_27841,N_27442);
nor U28751 (N_28751,N_27799,N_27469);
and U28752 (N_28752,N_27930,N_27427);
nand U28753 (N_28753,N_27679,N_27173);
nand U28754 (N_28754,N_27545,N_27080);
or U28755 (N_28755,N_27416,N_27258);
xnor U28756 (N_28756,N_27916,N_27529);
nand U28757 (N_28757,N_27818,N_27084);
and U28758 (N_28758,N_27569,N_27210);
nand U28759 (N_28759,N_27256,N_27167);
nand U28760 (N_28760,N_27253,N_27911);
xor U28761 (N_28761,N_27040,N_27922);
and U28762 (N_28762,N_27853,N_27582);
nand U28763 (N_28763,N_27073,N_27565);
nor U28764 (N_28764,N_27846,N_27612);
nand U28765 (N_28765,N_27846,N_27994);
nand U28766 (N_28766,N_27664,N_27282);
nand U28767 (N_28767,N_27447,N_27029);
nand U28768 (N_28768,N_27732,N_27480);
nand U28769 (N_28769,N_27895,N_27172);
or U28770 (N_28770,N_27328,N_27870);
nand U28771 (N_28771,N_27740,N_27812);
xnor U28772 (N_28772,N_27558,N_27654);
nor U28773 (N_28773,N_27813,N_27090);
nor U28774 (N_28774,N_27243,N_27928);
nand U28775 (N_28775,N_27447,N_27376);
or U28776 (N_28776,N_27312,N_27487);
and U28777 (N_28777,N_27795,N_27372);
xnor U28778 (N_28778,N_27045,N_27326);
and U28779 (N_28779,N_27789,N_27703);
and U28780 (N_28780,N_27235,N_27368);
or U28781 (N_28781,N_27440,N_27931);
or U28782 (N_28782,N_27384,N_27663);
nor U28783 (N_28783,N_27027,N_27884);
nor U28784 (N_28784,N_27818,N_27555);
nor U28785 (N_28785,N_27602,N_27394);
xor U28786 (N_28786,N_27755,N_27270);
nor U28787 (N_28787,N_27694,N_27974);
nand U28788 (N_28788,N_27398,N_27915);
or U28789 (N_28789,N_27909,N_27582);
or U28790 (N_28790,N_27915,N_27192);
and U28791 (N_28791,N_27897,N_27274);
or U28792 (N_28792,N_27295,N_27400);
xnor U28793 (N_28793,N_27565,N_27385);
and U28794 (N_28794,N_27783,N_27665);
nor U28795 (N_28795,N_27785,N_27649);
nor U28796 (N_28796,N_27748,N_27555);
xnor U28797 (N_28797,N_27335,N_27420);
nand U28798 (N_28798,N_27699,N_27680);
and U28799 (N_28799,N_27396,N_27493);
and U28800 (N_28800,N_27379,N_27406);
nand U28801 (N_28801,N_27040,N_27076);
nor U28802 (N_28802,N_27213,N_27380);
or U28803 (N_28803,N_27210,N_27288);
and U28804 (N_28804,N_27555,N_27954);
and U28805 (N_28805,N_27933,N_27299);
xor U28806 (N_28806,N_27767,N_27146);
and U28807 (N_28807,N_27684,N_27844);
and U28808 (N_28808,N_27628,N_27770);
xor U28809 (N_28809,N_27087,N_27927);
nand U28810 (N_28810,N_27290,N_27944);
nor U28811 (N_28811,N_27053,N_27392);
and U28812 (N_28812,N_27543,N_27547);
or U28813 (N_28813,N_27524,N_27968);
or U28814 (N_28814,N_27166,N_27151);
nor U28815 (N_28815,N_27631,N_27723);
and U28816 (N_28816,N_27774,N_27506);
and U28817 (N_28817,N_27372,N_27521);
and U28818 (N_28818,N_27213,N_27456);
xor U28819 (N_28819,N_27470,N_27510);
nor U28820 (N_28820,N_27559,N_27893);
xnor U28821 (N_28821,N_27772,N_27536);
nor U28822 (N_28822,N_27452,N_27959);
nand U28823 (N_28823,N_27167,N_27905);
or U28824 (N_28824,N_27792,N_27738);
nor U28825 (N_28825,N_27300,N_27269);
nor U28826 (N_28826,N_27534,N_27445);
nor U28827 (N_28827,N_27361,N_27400);
nor U28828 (N_28828,N_27704,N_27717);
xor U28829 (N_28829,N_27807,N_27125);
nor U28830 (N_28830,N_27645,N_27540);
nand U28831 (N_28831,N_27553,N_27826);
and U28832 (N_28832,N_27348,N_27840);
or U28833 (N_28833,N_27882,N_27878);
nor U28834 (N_28834,N_27739,N_27378);
xnor U28835 (N_28835,N_27765,N_27380);
or U28836 (N_28836,N_27993,N_27405);
or U28837 (N_28837,N_27477,N_27459);
nand U28838 (N_28838,N_27434,N_27007);
or U28839 (N_28839,N_27094,N_27523);
and U28840 (N_28840,N_27030,N_27871);
or U28841 (N_28841,N_27397,N_27445);
or U28842 (N_28842,N_27619,N_27770);
or U28843 (N_28843,N_27483,N_27209);
nand U28844 (N_28844,N_27014,N_27332);
nor U28845 (N_28845,N_27791,N_27525);
and U28846 (N_28846,N_27049,N_27762);
xnor U28847 (N_28847,N_27430,N_27891);
and U28848 (N_28848,N_27509,N_27400);
or U28849 (N_28849,N_27898,N_27798);
xnor U28850 (N_28850,N_27014,N_27547);
or U28851 (N_28851,N_27950,N_27937);
and U28852 (N_28852,N_27575,N_27449);
nor U28853 (N_28853,N_27114,N_27294);
or U28854 (N_28854,N_27544,N_27942);
and U28855 (N_28855,N_27881,N_27265);
and U28856 (N_28856,N_27688,N_27909);
xor U28857 (N_28857,N_27231,N_27951);
and U28858 (N_28858,N_27549,N_27246);
xor U28859 (N_28859,N_27354,N_27559);
xnor U28860 (N_28860,N_27275,N_27548);
xor U28861 (N_28861,N_27262,N_27476);
xor U28862 (N_28862,N_27782,N_27842);
nand U28863 (N_28863,N_27144,N_27366);
nor U28864 (N_28864,N_27895,N_27469);
or U28865 (N_28865,N_27870,N_27002);
and U28866 (N_28866,N_27675,N_27147);
nor U28867 (N_28867,N_27669,N_27561);
or U28868 (N_28868,N_27538,N_27966);
nand U28869 (N_28869,N_27774,N_27011);
nand U28870 (N_28870,N_27694,N_27351);
xor U28871 (N_28871,N_27909,N_27463);
and U28872 (N_28872,N_27029,N_27868);
and U28873 (N_28873,N_27364,N_27021);
xor U28874 (N_28874,N_27729,N_27517);
xnor U28875 (N_28875,N_27387,N_27346);
nor U28876 (N_28876,N_27964,N_27194);
nand U28877 (N_28877,N_27689,N_27361);
nand U28878 (N_28878,N_27643,N_27797);
xor U28879 (N_28879,N_27742,N_27564);
nor U28880 (N_28880,N_27602,N_27148);
nand U28881 (N_28881,N_27856,N_27723);
xor U28882 (N_28882,N_27172,N_27123);
and U28883 (N_28883,N_27610,N_27928);
or U28884 (N_28884,N_27146,N_27954);
xor U28885 (N_28885,N_27485,N_27194);
nor U28886 (N_28886,N_27476,N_27515);
and U28887 (N_28887,N_27119,N_27634);
xnor U28888 (N_28888,N_27478,N_27232);
or U28889 (N_28889,N_27322,N_27375);
and U28890 (N_28890,N_27597,N_27573);
and U28891 (N_28891,N_27711,N_27682);
and U28892 (N_28892,N_27076,N_27737);
and U28893 (N_28893,N_27850,N_27332);
nand U28894 (N_28894,N_27633,N_27588);
and U28895 (N_28895,N_27789,N_27718);
nor U28896 (N_28896,N_27147,N_27263);
or U28897 (N_28897,N_27882,N_27125);
nand U28898 (N_28898,N_27483,N_27144);
nand U28899 (N_28899,N_27960,N_27051);
or U28900 (N_28900,N_27802,N_27817);
and U28901 (N_28901,N_27938,N_27889);
xnor U28902 (N_28902,N_27504,N_27161);
nor U28903 (N_28903,N_27455,N_27982);
nand U28904 (N_28904,N_27621,N_27038);
nor U28905 (N_28905,N_27752,N_27231);
and U28906 (N_28906,N_27870,N_27150);
nor U28907 (N_28907,N_27493,N_27044);
nand U28908 (N_28908,N_27119,N_27442);
and U28909 (N_28909,N_27393,N_27113);
nand U28910 (N_28910,N_27523,N_27207);
xor U28911 (N_28911,N_27871,N_27915);
or U28912 (N_28912,N_27886,N_27613);
and U28913 (N_28913,N_27917,N_27693);
nand U28914 (N_28914,N_27401,N_27924);
and U28915 (N_28915,N_27361,N_27391);
and U28916 (N_28916,N_27946,N_27880);
or U28917 (N_28917,N_27634,N_27374);
xnor U28918 (N_28918,N_27023,N_27263);
or U28919 (N_28919,N_27049,N_27423);
and U28920 (N_28920,N_27675,N_27563);
nand U28921 (N_28921,N_27610,N_27875);
xor U28922 (N_28922,N_27101,N_27409);
nor U28923 (N_28923,N_27735,N_27680);
or U28924 (N_28924,N_27791,N_27303);
or U28925 (N_28925,N_27473,N_27908);
xor U28926 (N_28926,N_27953,N_27876);
nor U28927 (N_28927,N_27506,N_27329);
or U28928 (N_28928,N_27515,N_27223);
and U28929 (N_28929,N_27085,N_27600);
nor U28930 (N_28930,N_27700,N_27872);
nand U28931 (N_28931,N_27382,N_27435);
and U28932 (N_28932,N_27500,N_27634);
and U28933 (N_28933,N_27172,N_27777);
and U28934 (N_28934,N_27256,N_27801);
nand U28935 (N_28935,N_27345,N_27984);
xor U28936 (N_28936,N_27074,N_27353);
and U28937 (N_28937,N_27182,N_27054);
nor U28938 (N_28938,N_27107,N_27725);
and U28939 (N_28939,N_27334,N_27925);
xnor U28940 (N_28940,N_27510,N_27849);
or U28941 (N_28941,N_27568,N_27626);
nand U28942 (N_28942,N_27711,N_27874);
or U28943 (N_28943,N_27871,N_27276);
and U28944 (N_28944,N_27997,N_27259);
and U28945 (N_28945,N_27057,N_27072);
and U28946 (N_28946,N_27133,N_27676);
nand U28947 (N_28947,N_27149,N_27385);
or U28948 (N_28948,N_27633,N_27072);
or U28949 (N_28949,N_27160,N_27854);
and U28950 (N_28950,N_27452,N_27814);
and U28951 (N_28951,N_27525,N_27192);
and U28952 (N_28952,N_27900,N_27692);
xor U28953 (N_28953,N_27803,N_27531);
or U28954 (N_28954,N_27417,N_27004);
and U28955 (N_28955,N_27603,N_27218);
and U28956 (N_28956,N_27733,N_27143);
nand U28957 (N_28957,N_27418,N_27322);
xor U28958 (N_28958,N_27597,N_27247);
xnor U28959 (N_28959,N_27599,N_27738);
and U28960 (N_28960,N_27849,N_27454);
xnor U28961 (N_28961,N_27996,N_27874);
nor U28962 (N_28962,N_27372,N_27104);
nor U28963 (N_28963,N_27877,N_27697);
nand U28964 (N_28964,N_27611,N_27687);
xnor U28965 (N_28965,N_27303,N_27044);
nand U28966 (N_28966,N_27894,N_27737);
nand U28967 (N_28967,N_27897,N_27527);
and U28968 (N_28968,N_27636,N_27826);
xor U28969 (N_28969,N_27589,N_27029);
xor U28970 (N_28970,N_27275,N_27413);
and U28971 (N_28971,N_27937,N_27518);
nand U28972 (N_28972,N_27637,N_27099);
and U28973 (N_28973,N_27633,N_27897);
nor U28974 (N_28974,N_27621,N_27633);
nor U28975 (N_28975,N_27476,N_27750);
or U28976 (N_28976,N_27162,N_27707);
and U28977 (N_28977,N_27092,N_27091);
xor U28978 (N_28978,N_27453,N_27931);
or U28979 (N_28979,N_27546,N_27105);
and U28980 (N_28980,N_27120,N_27173);
or U28981 (N_28981,N_27110,N_27487);
nand U28982 (N_28982,N_27472,N_27156);
nand U28983 (N_28983,N_27273,N_27933);
nor U28984 (N_28984,N_27409,N_27978);
or U28985 (N_28985,N_27905,N_27137);
and U28986 (N_28986,N_27148,N_27531);
or U28987 (N_28987,N_27663,N_27572);
and U28988 (N_28988,N_27339,N_27309);
nand U28989 (N_28989,N_27925,N_27840);
nor U28990 (N_28990,N_27237,N_27905);
and U28991 (N_28991,N_27330,N_27761);
xor U28992 (N_28992,N_27165,N_27991);
xor U28993 (N_28993,N_27327,N_27389);
nand U28994 (N_28994,N_27081,N_27126);
nor U28995 (N_28995,N_27893,N_27500);
or U28996 (N_28996,N_27979,N_27024);
and U28997 (N_28997,N_27951,N_27586);
xnor U28998 (N_28998,N_27805,N_27809);
and U28999 (N_28999,N_27063,N_27019);
and U29000 (N_29000,N_28501,N_28456);
or U29001 (N_29001,N_28414,N_28248);
or U29002 (N_29002,N_28965,N_28484);
xor U29003 (N_29003,N_28706,N_28832);
and U29004 (N_29004,N_28698,N_28566);
and U29005 (N_29005,N_28780,N_28664);
or U29006 (N_29006,N_28038,N_28629);
and U29007 (N_29007,N_28081,N_28144);
xnor U29008 (N_29008,N_28554,N_28959);
nand U29009 (N_29009,N_28788,N_28328);
nand U29010 (N_29010,N_28684,N_28445);
and U29011 (N_29011,N_28278,N_28578);
and U29012 (N_29012,N_28107,N_28624);
and U29013 (N_29013,N_28340,N_28114);
or U29014 (N_29014,N_28517,N_28619);
nand U29015 (N_29015,N_28504,N_28295);
and U29016 (N_29016,N_28928,N_28031);
nand U29017 (N_29017,N_28329,N_28796);
or U29018 (N_29018,N_28332,N_28151);
or U29019 (N_29019,N_28049,N_28431);
nand U29020 (N_29020,N_28660,N_28129);
xnor U29021 (N_29021,N_28705,N_28604);
and U29022 (N_29022,N_28206,N_28806);
xnor U29023 (N_29023,N_28347,N_28690);
nand U29024 (N_29024,N_28557,N_28016);
or U29025 (N_29025,N_28040,N_28791);
and U29026 (N_29026,N_28070,N_28886);
nor U29027 (N_29027,N_28012,N_28869);
xnor U29028 (N_29028,N_28822,N_28785);
xor U29029 (N_29029,N_28131,N_28100);
nand U29030 (N_29030,N_28801,N_28051);
and U29031 (N_29031,N_28905,N_28355);
xor U29032 (N_29032,N_28180,N_28429);
xor U29033 (N_29033,N_28699,N_28942);
or U29034 (N_29034,N_28458,N_28290);
xnor U29035 (N_29035,N_28688,N_28149);
or U29036 (N_29036,N_28298,N_28462);
or U29037 (N_29037,N_28628,N_28286);
or U29038 (N_29038,N_28715,N_28064);
and U29039 (N_29039,N_28982,N_28769);
xnor U29040 (N_29040,N_28083,N_28020);
xor U29041 (N_29041,N_28167,N_28103);
and U29042 (N_29042,N_28175,N_28187);
xor U29043 (N_29043,N_28090,N_28283);
nor U29044 (N_29044,N_28923,N_28954);
xor U29045 (N_29045,N_28205,N_28743);
and U29046 (N_29046,N_28249,N_28618);
xor U29047 (N_29047,N_28343,N_28021);
xnor U29048 (N_29048,N_28387,N_28874);
or U29049 (N_29049,N_28995,N_28211);
or U29050 (N_29050,N_28838,N_28480);
or U29051 (N_29051,N_28846,N_28765);
nand U29052 (N_29052,N_28652,N_28555);
and U29053 (N_29053,N_28738,N_28243);
nor U29054 (N_29054,N_28645,N_28666);
nor U29055 (N_29055,N_28888,N_28845);
or U29056 (N_29056,N_28018,N_28756);
and U29057 (N_29057,N_28539,N_28717);
nor U29058 (N_29058,N_28198,N_28703);
and U29059 (N_29059,N_28316,N_28241);
nand U29060 (N_29060,N_28068,N_28852);
xnor U29061 (N_29061,N_28086,N_28659);
xnor U29062 (N_29062,N_28321,N_28774);
xor U29063 (N_29063,N_28382,N_28908);
xor U29064 (N_29064,N_28779,N_28981);
xor U29065 (N_29065,N_28830,N_28558);
or U29066 (N_29066,N_28394,N_28572);
xor U29067 (N_29067,N_28957,N_28448);
and U29068 (N_29068,N_28045,N_28194);
xor U29069 (N_29069,N_28719,N_28369);
nor U29070 (N_29070,N_28677,N_28877);
nand U29071 (N_29071,N_28541,N_28342);
nor U29072 (N_29072,N_28204,N_28617);
nor U29073 (N_29073,N_28483,N_28140);
or U29074 (N_29074,N_28271,N_28697);
and U29075 (N_29075,N_28071,N_28457);
and U29076 (N_29076,N_28777,N_28672);
xor U29077 (N_29077,N_28804,N_28514);
nor U29078 (N_29078,N_28902,N_28236);
and U29079 (N_29079,N_28136,N_28401);
xor U29080 (N_29080,N_28179,N_28609);
and U29081 (N_29081,N_28190,N_28653);
nand U29082 (N_29082,N_28146,N_28816);
and U29083 (N_29083,N_28543,N_28354);
and U29084 (N_29084,N_28282,N_28800);
xor U29085 (N_29085,N_28824,N_28306);
nand U29086 (N_29086,N_28858,N_28868);
nand U29087 (N_29087,N_28899,N_28217);
nand U29088 (N_29088,N_28912,N_28900);
nor U29089 (N_29089,N_28178,N_28058);
or U29090 (N_29090,N_28790,N_28663);
nor U29091 (N_29091,N_28885,N_28926);
nand U29092 (N_29092,N_28571,N_28671);
nand U29093 (N_29093,N_28132,N_28574);
nand U29094 (N_29094,N_28422,N_28833);
nand U29095 (N_29095,N_28255,N_28296);
nor U29096 (N_29096,N_28904,N_28635);
xnor U29097 (N_29097,N_28240,N_28693);
nand U29098 (N_29098,N_28017,N_28610);
xnor U29099 (N_29099,N_28958,N_28466);
or U29100 (N_29100,N_28261,N_28828);
or U29101 (N_29101,N_28889,N_28265);
xnor U29102 (N_29102,N_28390,N_28542);
xor U29103 (N_29103,N_28365,N_28915);
nor U29104 (N_29104,N_28569,N_28985);
nand U29105 (N_29105,N_28360,N_28423);
xnor U29106 (N_29106,N_28246,N_28642);
or U29107 (N_29107,N_28091,N_28977);
or U29108 (N_29108,N_28124,N_28587);
nor U29109 (N_29109,N_28405,N_28510);
xor U29110 (N_29110,N_28815,N_28605);
or U29111 (N_29111,N_28043,N_28583);
nand U29112 (N_29112,N_28075,N_28884);
nand U29113 (N_29113,N_28106,N_28437);
xnor U29114 (N_29114,N_28661,N_28063);
xor U29115 (N_29115,N_28399,N_28223);
nor U29116 (N_29116,N_28277,N_28023);
and U29117 (N_29117,N_28503,N_28444);
or U29118 (N_29118,N_28507,N_28960);
nand U29119 (N_29119,N_28259,N_28389);
xnor U29120 (N_29120,N_28632,N_28536);
nand U29121 (N_29121,N_28513,N_28381);
nor U29122 (N_29122,N_28914,N_28611);
nand U29123 (N_29123,N_28521,N_28334);
and U29124 (N_29124,N_28455,N_28089);
and U29125 (N_29125,N_28742,N_28913);
or U29126 (N_29126,N_28077,N_28579);
nor U29127 (N_29127,N_28158,N_28173);
and U29128 (N_29128,N_28430,N_28475);
xnor U29129 (N_29129,N_28254,N_28512);
xnor U29130 (N_29130,N_28907,N_28922);
nor U29131 (N_29131,N_28764,N_28979);
nand U29132 (N_29132,N_28966,N_28850);
nor U29133 (N_29133,N_28096,N_28119);
nand U29134 (N_29134,N_28741,N_28324);
and U29135 (N_29135,N_28820,N_28084);
xor U29136 (N_29136,N_28792,N_28760);
xor U29137 (N_29137,N_28188,N_28710);
nor U29138 (N_29138,N_28166,N_28668);
xnor U29139 (N_29139,N_28770,N_28729);
nor U29140 (N_29140,N_28944,N_28681);
and U29141 (N_29141,N_28807,N_28320);
xnor U29142 (N_29142,N_28039,N_28358);
nor U29143 (N_29143,N_28171,N_28505);
nand U29144 (N_29144,N_28950,N_28116);
xnor U29145 (N_29145,N_28991,N_28150);
or U29146 (N_29146,N_28910,N_28172);
nor U29147 (N_29147,N_28613,N_28776);
xor U29148 (N_29148,N_28451,N_28214);
or U29149 (N_29149,N_28585,N_28099);
xor U29150 (N_29150,N_28812,N_28500);
nand U29151 (N_29151,N_28622,N_28753);
nor U29152 (N_29152,N_28999,N_28208);
xnor U29153 (N_29153,N_28032,N_28485);
nand U29154 (N_29154,N_28728,N_28933);
nand U29155 (N_29155,N_28808,N_28191);
nor U29156 (N_29156,N_28597,N_28141);
nor U29157 (N_29157,N_28819,N_28487);
nand U29158 (N_29158,N_28007,N_28392);
or U29159 (N_29159,N_28949,N_28641);
nand U29160 (N_29160,N_28643,N_28549);
xnor U29161 (N_29161,N_28526,N_28582);
or U29162 (N_29162,N_28887,N_28297);
nand U29163 (N_29163,N_28030,N_28798);
and U29164 (N_29164,N_28708,N_28990);
nand U29165 (N_29165,N_28294,N_28493);
nor U29166 (N_29166,N_28312,N_28094);
nand U29167 (N_29167,N_28386,N_28013);
or U29168 (N_29168,N_28257,N_28101);
and U29169 (N_29169,N_28714,N_28176);
nand U29170 (N_29170,N_28916,N_28184);
nand U29171 (N_29171,N_28955,N_28074);
nand U29172 (N_29172,N_28772,N_28408);
or U29173 (N_29173,N_28936,N_28145);
xor U29174 (N_29174,N_28123,N_28130);
or U29175 (N_29175,N_28199,N_28875);
and U29176 (N_29176,N_28417,N_28871);
nand U29177 (N_29177,N_28670,N_28065);
or U29178 (N_29178,N_28309,N_28285);
xor U29179 (N_29179,N_28799,N_28771);
and U29180 (N_29180,N_28658,N_28351);
or U29181 (N_29181,N_28657,N_28404);
nand U29182 (N_29182,N_28055,N_28528);
nor U29183 (N_29183,N_28047,N_28687);
and U29184 (N_29184,N_28281,N_28305);
nand U29185 (N_29185,N_28683,N_28441);
or U29186 (N_29186,N_28362,N_28720);
and U29187 (N_29187,N_28689,N_28425);
nand U29188 (N_29188,N_28436,N_28567);
nor U29189 (N_29189,N_28247,N_28925);
nor U29190 (N_29190,N_28440,N_28435);
nand U29191 (N_29191,N_28128,N_28280);
nand U29192 (N_29192,N_28491,N_28758);
or U29193 (N_29193,N_28856,N_28341);
xnor U29194 (N_29194,N_28842,N_28473);
nor U29195 (N_29195,N_28143,N_28215);
nand U29196 (N_29196,N_28268,N_28700);
xor U29197 (N_29197,N_28073,N_28793);
nand U29198 (N_29198,N_28046,N_28336);
xnor U29199 (N_29199,N_28607,N_28373);
nand U29200 (N_29200,N_28468,N_28576);
xor U29201 (N_29201,N_28872,N_28695);
nor U29202 (N_29202,N_28980,N_28454);
or U29203 (N_29203,N_28834,N_28213);
nand U29204 (N_29204,N_28943,N_28606);
nor U29205 (N_29205,N_28725,N_28426);
nand U29206 (N_29206,N_28827,N_28581);
xor U29207 (N_29207,N_28079,N_28533);
xnor U29208 (N_29208,N_28733,N_28037);
nor U29209 (N_29209,N_28522,N_28863);
or U29210 (N_29210,N_28163,N_28739);
or U29211 (N_29211,N_28797,N_28972);
nand U29212 (N_29212,N_28552,N_28495);
xor U29213 (N_29213,N_28357,N_28849);
nor U29214 (N_29214,N_28072,N_28269);
and U29215 (N_29215,N_28153,N_28831);
nand U29216 (N_29216,N_28478,N_28011);
and U29217 (N_29217,N_28301,N_28929);
nand U29218 (N_29218,N_28197,N_28380);
nand U29219 (N_29219,N_28773,N_28319);
nor U29220 (N_29220,N_28344,N_28449);
nand U29221 (N_29221,N_28335,N_28443);
or U29222 (N_29222,N_28718,N_28402);
nor U29223 (N_29223,N_28640,N_28034);
or U29224 (N_29224,N_28447,N_28655);
and U29225 (N_29225,N_28631,N_28962);
xor U29226 (N_29226,N_28366,N_28564);
xnor U29227 (N_29227,N_28292,N_28302);
or U29228 (N_29228,N_28497,N_28156);
nand U29229 (N_29229,N_28472,N_28104);
xor U29230 (N_29230,N_28623,N_28711);
or U29231 (N_29231,N_28327,N_28044);
or U29232 (N_29232,N_28596,N_28069);
nand U29233 (N_29233,N_28529,N_28299);
nor U29234 (N_29234,N_28275,N_28767);
nand U29235 (N_29235,N_28740,N_28917);
or U29236 (N_29236,N_28397,N_28761);
and U29237 (N_29237,N_28288,N_28676);
xor U29238 (N_29238,N_28696,N_28234);
or U29239 (N_29239,N_28967,N_28396);
xor U29240 (N_29240,N_28311,N_28494);
or U29241 (N_29241,N_28378,N_28679);
xor U29242 (N_29242,N_28766,N_28182);
nand U29243 (N_29243,N_28352,N_28775);
nand U29244 (N_29244,N_28303,N_28946);
nor U29245 (N_29245,N_28704,N_28398);
nand U29246 (N_29246,N_28250,N_28379);
or U29247 (N_29247,N_28759,N_28372);
nor U29248 (N_29248,N_28519,N_28008);
and U29249 (N_29249,N_28580,N_28847);
xnor U29250 (N_29250,N_28598,N_28548);
nor U29251 (N_29251,N_28573,N_28975);
nor U29252 (N_29252,N_28854,N_28147);
or U29253 (N_29253,N_28515,N_28228);
or U29254 (N_29254,N_28446,N_28052);
xor U29255 (N_29255,N_28464,N_28345);
nor U29256 (N_29256,N_28750,N_28844);
nand U29257 (N_29257,N_28486,N_28749);
xnor U29258 (N_29258,N_28562,N_28803);
and U29259 (N_29259,N_28675,N_28867);
nor U29260 (N_29260,N_28004,N_28196);
nand U29261 (N_29261,N_28721,N_28022);
and U29262 (N_29262,N_28538,N_28941);
nor U29263 (N_29263,N_28627,N_28127);
xnor U29264 (N_29264,N_28864,N_28821);
and U29265 (N_29265,N_28841,N_28656);
xor U29266 (N_29266,N_28968,N_28594);
xnor U29267 (N_29267,N_28986,N_28731);
or U29268 (N_29268,N_28921,N_28633);
nor U29269 (N_29269,N_28621,N_28452);
or U29270 (N_29270,N_28474,N_28823);
nand U29271 (N_29271,N_28019,N_28424);
xnor U29272 (N_29272,N_28577,N_28253);
or U29273 (N_29273,N_28918,N_28691);
and U29274 (N_29274,N_28097,N_28192);
nor U29275 (N_29275,N_28644,N_28202);
nand U29276 (N_29276,N_28951,N_28251);
or U29277 (N_29277,N_28836,N_28570);
and U29278 (N_29278,N_28245,N_28680);
nand U29279 (N_29279,N_28947,N_28974);
xor U29280 (N_29280,N_28825,N_28420);
nor U29281 (N_29281,N_28005,N_28233);
and U29282 (N_29282,N_28783,N_28238);
nand U29283 (N_29283,N_28882,N_28556);
nand U29284 (N_29284,N_28476,N_28109);
or U29285 (N_29285,N_28789,N_28135);
xor U29286 (N_29286,N_28155,N_28665);
xor U29287 (N_29287,N_28873,N_28252);
nand U29288 (N_29288,N_28006,N_28203);
nand U29289 (N_29289,N_28053,N_28961);
and U29290 (N_29290,N_28160,N_28612);
xnor U29291 (N_29291,N_28561,N_28839);
and U29292 (N_29292,N_28210,N_28048);
xor U29293 (N_29293,N_28744,N_28673);
nand U29294 (N_29294,N_28218,N_28209);
xor U29295 (N_29295,N_28161,N_28811);
xnor U29296 (N_29296,N_28125,N_28620);
or U29297 (N_29297,N_28862,N_28971);
nor U29298 (N_29298,N_28427,N_28222);
nor U29299 (N_29299,N_28270,N_28370);
nor U29300 (N_29300,N_28989,N_28459);
nand U29301 (N_29301,N_28630,N_28757);
and U29302 (N_29302,N_28300,N_28752);
nand U29303 (N_29303,N_28168,N_28407);
xnor U29304 (N_29304,N_28263,N_28927);
and U29305 (N_29305,N_28952,N_28216);
nor U29306 (N_29306,N_28326,N_28367);
nor U29307 (N_29307,N_28080,N_28590);
xor U29308 (N_29308,N_28393,N_28723);
or U29309 (N_29309,N_28421,N_28148);
or U29310 (N_29310,N_28919,N_28139);
and U29311 (N_29311,N_28066,N_28726);
and U29312 (N_29312,N_28502,N_28242);
and U29313 (N_29313,N_28551,N_28932);
nand U29314 (N_29314,N_28550,N_28460);
and U29315 (N_29315,N_28453,N_28553);
and U29316 (N_29316,N_28442,N_28225);
and U29317 (N_29317,N_28880,N_28639);
xor U29318 (N_29318,N_28057,N_28122);
nand U29319 (N_29319,N_28289,N_28395);
xnor U29320 (N_29320,N_28374,N_28050);
xor U29321 (N_29321,N_28105,N_28559);
or U29322 (N_29322,N_28010,N_28111);
or U29323 (N_29323,N_28088,N_28356);
nand U29324 (N_29324,N_28601,N_28786);
nand U29325 (N_29325,N_28102,N_28787);
nor U29326 (N_29326,N_28963,N_28428);
nand U29327 (N_29327,N_28809,N_28207);
or U29328 (N_29328,N_28463,N_28523);
and U29329 (N_29329,N_28778,N_28901);
xnor U29330 (N_29330,N_28813,N_28488);
and U29331 (N_29331,N_28227,N_28230);
or U29332 (N_29332,N_28406,N_28937);
and U29333 (N_29333,N_28185,N_28909);
nand U29334 (N_29334,N_28348,N_28054);
nor U29335 (N_29335,N_28865,N_28121);
nand U29336 (N_29336,N_28751,N_28036);
and U29337 (N_29337,N_28992,N_28226);
nand U29338 (N_29338,N_28498,N_28595);
or U29339 (N_29339,N_28322,N_28924);
or U29340 (N_29340,N_28713,N_28647);
and U29341 (N_29341,N_28108,N_28120);
nor U29342 (N_29342,N_28650,N_28634);
xnor U29343 (N_29343,N_28368,N_28667);
and U29344 (N_29344,N_28814,N_28266);
or U29345 (N_29345,N_28026,N_28520);
or U29346 (N_29346,N_28898,N_28000);
nand U29347 (N_29347,N_28076,N_28857);
and U29348 (N_29348,N_28892,N_28973);
nor U29349 (N_29349,N_28860,N_28138);
or U29350 (N_29350,N_28730,N_28893);
and U29351 (N_29351,N_28648,N_28859);
xor U29352 (N_29352,N_28669,N_28938);
nor U29353 (N_29353,N_28279,N_28896);
and U29354 (N_29354,N_28716,N_28231);
xor U29355 (N_29355,N_28537,N_28535);
nand U29356 (N_29356,N_28056,N_28126);
xor U29357 (N_29357,N_28317,N_28685);
nor U29358 (N_29358,N_28042,N_28035);
or U29359 (N_29359,N_28997,N_28575);
and U29360 (N_29360,N_28993,N_28547);
nand U29361 (N_29361,N_28383,N_28707);
xor U29362 (N_29362,N_28433,N_28152);
or U29363 (N_29363,N_28939,N_28264);
nor U29364 (N_29364,N_28608,N_28654);
or U29365 (N_29365,N_28747,N_28724);
nor U29366 (N_29366,N_28244,N_28256);
and U29367 (N_29367,N_28385,N_28337);
nand U29368 (N_29368,N_28384,N_28878);
or U29369 (N_29369,N_28411,N_28310);
and U29370 (N_29370,N_28200,N_28735);
nand U29371 (N_29371,N_28028,N_28376);
nor U29372 (N_29372,N_28059,N_28001);
and U29373 (N_29373,N_28763,N_28157);
nor U29374 (N_29374,N_28881,N_28930);
nor U29375 (N_29375,N_28015,N_28674);
nor U29376 (N_29376,N_28637,N_28636);
xor U29377 (N_29377,N_28477,N_28061);
and U29378 (N_29378,N_28260,N_28614);
and U29379 (N_29379,N_28870,N_28489);
nand U29380 (N_29380,N_28482,N_28784);
xor U29381 (N_29381,N_28692,N_28067);
and U29382 (N_29382,N_28524,N_28181);
and U29383 (N_29383,N_28220,N_28615);
nor U29384 (N_29384,N_28987,N_28755);
and U29385 (N_29385,N_28291,N_28174);
nor U29386 (N_29386,N_28984,N_28115);
nor U29387 (N_29387,N_28781,N_28722);
xor U29388 (N_29388,N_28239,N_28235);
nand U29389 (N_29389,N_28432,N_28732);
nor U29390 (N_29390,N_28201,N_28626);
nor U29391 (N_29391,N_28994,N_28906);
and U29392 (N_29392,N_28748,N_28272);
xnor U29393 (N_29393,N_28829,N_28212);
or U29394 (N_29394,N_28826,N_28532);
and U29395 (N_29395,N_28304,N_28866);
nand U29396 (N_29396,N_28325,N_28403);
nor U29397 (N_29397,N_28313,N_28409);
nor U29398 (N_29398,N_28469,N_28848);
xnor U29399 (N_29399,N_28391,N_28646);
or U29400 (N_29400,N_28586,N_28195);
and U29401 (N_29401,N_28388,N_28229);
nor U29402 (N_29402,N_28082,N_28479);
nand U29403 (N_29403,N_28592,N_28085);
or U29404 (N_29404,N_28600,N_28940);
xnor U29405 (N_29405,N_28170,N_28258);
nor U29406 (N_29406,N_28307,N_28419);
or U29407 (N_29407,N_28333,N_28353);
and U29408 (N_29408,N_28177,N_28438);
xor U29409 (N_29409,N_28511,N_28754);
nand U29410 (N_29410,N_28817,N_28400);
or U29411 (N_29411,N_28883,N_28638);
and U29412 (N_29412,N_28346,N_28948);
nor U29413 (N_29413,N_28560,N_28712);
and U29414 (N_29414,N_28371,N_28467);
nor U29415 (N_29415,N_28359,N_28033);
and U29416 (N_29416,N_28599,N_28330);
nor U29417 (N_29417,N_28092,N_28189);
xnor U29418 (N_29418,N_28891,N_28186);
or U29419 (N_29419,N_28686,N_28516);
xnor U29420 (N_29420,N_28142,N_28274);
xnor U29421 (N_29421,N_28794,N_28110);
and U29422 (N_29422,N_28339,N_28481);
nand U29423 (N_29423,N_28025,N_28041);
xnor U29424 (N_29424,N_28616,N_28287);
nor U29425 (N_29425,N_28293,N_28087);
nor U29426 (N_29426,N_28024,N_28361);
or U29427 (N_29427,N_28262,N_28527);
and U29428 (N_29428,N_28450,N_28953);
and U29429 (N_29429,N_28133,N_28903);
nand U29430 (N_29430,N_28745,N_28591);
nor U29431 (N_29431,N_28805,N_28471);
and U29432 (N_29432,N_28563,N_28509);
nor U29433 (N_29433,N_28589,N_28531);
or U29434 (N_29434,N_28835,N_28095);
and U29435 (N_29435,N_28651,N_28273);
nor U29436 (N_29436,N_28988,N_28118);
or U29437 (N_29437,N_28945,N_28237);
and U29438 (N_29438,N_28678,N_28534);
or U29439 (N_29439,N_28183,N_28546);
nor U29440 (N_29440,N_28978,N_28415);
xnor U29441 (N_29441,N_28470,N_28169);
xnor U29442 (N_29442,N_28920,N_28843);
xor U29443 (N_29443,N_28802,N_28593);
nor U29444 (N_29444,N_28009,N_28314);
nand U29445 (N_29445,N_28465,N_28350);
nand U29446 (N_29446,N_28709,N_28461);
or U29447 (N_29447,N_28439,N_28490);
xor U29448 (N_29448,N_28364,N_28544);
nand U29449 (N_29449,N_28837,N_28956);
nand U29450 (N_29450,N_28694,N_28662);
xnor U29451 (N_29451,N_28029,N_28818);
nor U29452 (N_29452,N_28737,N_28970);
or U29453 (N_29453,N_28861,N_28412);
nor U29454 (N_29454,N_28879,N_28002);
and U29455 (N_29455,N_28284,N_28232);
or U29456 (N_29456,N_28701,N_28315);
xor U29457 (N_29457,N_28768,N_28377);
nand U29458 (N_29458,N_28588,N_28062);
nor U29459 (N_29459,N_28876,N_28894);
or U29460 (N_29460,N_28060,N_28702);
xnor U29461 (N_29461,N_28318,N_28782);
or U29462 (N_29462,N_28413,N_28518);
nor U29463 (N_29463,N_28331,N_28983);
xnor U29464 (N_29464,N_28602,N_28113);
nand U29465 (N_29465,N_28969,N_28996);
nor U29466 (N_29466,N_28349,N_28810);
nor U29467 (N_29467,N_28276,N_28625);
nor U29468 (N_29468,N_28727,N_28736);
nand U29469 (N_29469,N_28897,N_28911);
nand U29470 (N_29470,N_28410,N_28193);
nand U29471 (N_29471,N_28098,N_28525);
nand U29472 (N_29472,N_28308,N_28164);
and U29473 (N_29473,N_28682,N_28434);
nand U29474 (N_29474,N_28162,N_28112);
nand U29475 (N_29475,N_28649,N_28545);
nand U29476 (N_29476,N_28078,N_28221);
or U29477 (N_29477,N_28976,N_28134);
and U29478 (N_29478,N_28935,N_28323);
xnor U29479 (N_29479,N_28734,N_28746);
xnor U29480 (N_29480,N_28851,N_28499);
xnor U29481 (N_29481,N_28895,N_28224);
or U29482 (N_29482,N_28418,N_28506);
xnor U29483 (N_29483,N_28219,N_28338);
or U29484 (N_29484,N_28267,N_28165);
nor U29485 (N_29485,N_28416,N_28890);
and U29486 (N_29486,N_28530,N_28508);
xor U29487 (N_29487,N_28934,N_28855);
xnor U29488 (N_29488,N_28964,N_28931);
xor U29489 (N_29489,N_28027,N_28093);
or U29490 (N_29490,N_28998,N_28014);
nor U29491 (N_29491,N_28492,N_28603);
nand U29492 (N_29492,N_28363,N_28565);
or U29493 (N_29493,N_28540,N_28568);
xor U29494 (N_29494,N_28795,N_28853);
and U29495 (N_29495,N_28154,N_28375);
nand U29496 (N_29496,N_28003,N_28840);
and U29497 (N_29497,N_28496,N_28762);
and U29498 (N_29498,N_28584,N_28137);
or U29499 (N_29499,N_28117,N_28159);
nand U29500 (N_29500,N_28582,N_28440);
and U29501 (N_29501,N_28249,N_28406);
nor U29502 (N_29502,N_28666,N_28746);
or U29503 (N_29503,N_28315,N_28211);
and U29504 (N_29504,N_28647,N_28575);
or U29505 (N_29505,N_28744,N_28954);
xor U29506 (N_29506,N_28613,N_28163);
nor U29507 (N_29507,N_28312,N_28256);
nor U29508 (N_29508,N_28086,N_28283);
xor U29509 (N_29509,N_28703,N_28569);
and U29510 (N_29510,N_28220,N_28791);
nor U29511 (N_29511,N_28100,N_28346);
xor U29512 (N_29512,N_28957,N_28853);
and U29513 (N_29513,N_28042,N_28115);
or U29514 (N_29514,N_28598,N_28899);
and U29515 (N_29515,N_28452,N_28083);
nand U29516 (N_29516,N_28100,N_28438);
or U29517 (N_29517,N_28319,N_28219);
nand U29518 (N_29518,N_28239,N_28700);
nand U29519 (N_29519,N_28084,N_28542);
xor U29520 (N_29520,N_28777,N_28626);
and U29521 (N_29521,N_28841,N_28515);
and U29522 (N_29522,N_28783,N_28467);
nand U29523 (N_29523,N_28407,N_28866);
and U29524 (N_29524,N_28751,N_28618);
xor U29525 (N_29525,N_28510,N_28419);
or U29526 (N_29526,N_28649,N_28903);
nor U29527 (N_29527,N_28773,N_28440);
nor U29528 (N_29528,N_28310,N_28397);
nand U29529 (N_29529,N_28800,N_28268);
and U29530 (N_29530,N_28342,N_28134);
and U29531 (N_29531,N_28377,N_28600);
or U29532 (N_29532,N_28019,N_28934);
xor U29533 (N_29533,N_28110,N_28100);
xnor U29534 (N_29534,N_28422,N_28690);
nand U29535 (N_29535,N_28080,N_28846);
nor U29536 (N_29536,N_28027,N_28237);
xor U29537 (N_29537,N_28606,N_28927);
and U29538 (N_29538,N_28617,N_28051);
or U29539 (N_29539,N_28205,N_28310);
or U29540 (N_29540,N_28689,N_28272);
or U29541 (N_29541,N_28168,N_28756);
nand U29542 (N_29542,N_28076,N_28985);
and U29543 (N_29543,N_28623,N_28558);
nor U29544 (N_29544,N_28515,N_28801);
and U29545 (N_29545,N_28700,N_28364);
or U29546 (N_29546,N_28453,N_28892);
and U29547 (N_29547,N_28861,N_28644);
or U29548 (N_29548,N_28230,N_28581);
nand U29549 (N_29549,N_28519,N_28093);
nor U29550 (N_29550,N_28096,N_28106);
xor U29551 (N_29551,N_28910,N_28025);
nand U29552 (N_29552,N_28181,N_28109);
xnor U29553 (N_29553,N_28146,N_28971);
nor U29554 (N_29554,N_28534,N_28248);
or U29555 (N_29555,N_28839,N_28191);
xnor U29556 (N_29556,N_28382,N_28090);
nand U29557 (N_29557,N_28686,N_28773);
or U29558 (N_29558,N_28113,N_28673);
and U29559 (N_29559,N_28726,N_28481);
nand U29560 (N_29560,N_28608,N_28878);
or U29561 (N_29561,N_28173,N_28807);
xnor U29562 (N_29562,N_28438,N_28625);
or U29563 (N_29563,N_28545,N_28466);
and U29564 (N_29564,N_28492,N_28197);
xor U29565 (N_29565,N_28578,N_28136);
and U29566 (N_29566,N_28565,N_28594);
or U29567 (N_29567,N_28953,N_28972);
or U29568 (N_29568,N_28340,N_28305);
or U29569 (N_29569,N_28387,N_28651);
and U29570 (N_29570,N_28818,N_28395);
or U29571 (N_29571,N_28576,N_28670);
and U29572 (N_29572,N_28566,N_28697);
or U29573 (N_29573,N_28295,N_28370);
and U29574 (N_29574,N_28023,N_28650);
nor U29575 (N_29575,N_28825,N_28619);
or U29576 (N_29576,N_28922,N_28680);
or U29577 (N_29577,N_28443,N_28103);
xnor U29578 (N_29578,N_28819,N_28529);
nor U29579 (N_29579,N_28379,N_28125);
nand U29580 (N_29580,N_28461,N_28233);
nand U29581 (N_29581,N_28253,N_28085);
or U29582 (N_29582,N_28035,N_28218);
xor U29583 (N_29583,N_28157,N_28358);
nand U29584 (N_29584,N_28254,N_28799);
and U29585 (N_29585,N_28851,N_28403);
nand U29586 (N_29586,N_28050,N_28848);
nor U29587 (N_29587,N_28306,N_28799);
and U29588 (N_29588,N_28160,N_28776);
nor U29589 (N_29589,N_28222,N_28749);
nor U29590 (N_29590,N_28567,N_28793);
and U29591 (N_29591,N_28339,N_28003);
or U29592 (N_29592,N_28859,N_28479);
nand U29593 (N_29593,N_28616,N_28429);
nand U29594 (N_29594,N_28399,N_28554);
and U29595 (N_29595,N_28211,N_28895);
nand U29596 (N_29596,N_28941,N_28439);
nand U29597 (N_29597,N_28971,N_28601);
nor U29598 (N_29598,N_28229,N_28255);
and U29599 (N_29599,N_28687,N_28857);
nand U29600 (N_29600,N_28830,N_28325);
nor U29601 (N_29601,N_28872,N_28995);
nand U29602 (N_29602,N_28011,N_28052);
xor U29603 (N_29603,N_28052,N_28586);
nor U29604 (N_29604,N_28789,N_28902);
nand U29605 (N_29605,N_28662,N_28565);
xnor U29606 (N_29606,N_28349,N_28321);
and U29607 (N_29607,N_28278,N_28253);
xor U29608 (N_29608,N_28010,N_28047);
xnor U29609 (N_29609,N_28938,N_28831);
nand U29610 (N_29610,N_28165,N_28496);
and U29611 (N_29611,N_28347,N_28090);
and U29612 (N_29612,N_28079,N_28300);
xnor U29613 (N_29613,N_28613,N_28499);
and U29614 (N_29614,N_28280,N_28988);
nor U29615 (N_29615,N_28052,N_28654);
and U29616 (N_29616,N_28132,N_28694);
xnor U29617 (N_29617,N_28064,N_28453);
and U29618 (N_29618,N_28095,N_28895);
xor U29619 (N_29619,N_28950,N_28008);
nand U29620 (N_29620,N_28786,N_28054);
and U29621 (N_29621,N_28643,N_28834);
nor U29622 (N_29622,N_28585,N_28603);
and U29623 (N_29623,N_28937,N_28754);
xnor U29624 (N_29624,N_28236,N_28754);
nand U29625 (N_29625,N_28996,N_28824);
nor U29626 (N_29626,N_28851,N_28573);
xor U29627 (N_29627,N_28539,N_28735);
and U29628 (N_29628,N_28981,N_28330);
nand U29629 (N_29629,N_28373,N_28417);
nand U29630 (N_29630,N_28668,N_28874);
nand U29631 (N_29631,N_28571,N_28996);
and U29632 (N_29632,N_28596,N_28293);
or U29633 (N_29633,N_28482,N_28693);
or U29634 (N_29634,N_28218,N_28831);
nand U29635 (N_29635,N_28736,N_28111);
nand U29636 (N_29636,N_28068,N_28012);
nor U29637 (N_29637,N_28886,N_28160);
or U29638 (N_29638,N_28657,N_28364);
or U29639 (N_29639,N_28150,N_28167);
nand U29640 (N_29640,N_28285,N_28049);
nand U29641 (N_29641,N_28557,N_28239);
and U29642 (N_29642,N_28949,N_28688);
or U29643 (N_29643,N_28141,N_28112);
nor U29644 (N_29644,N_28582,N_28016);
nor U29645 (N_29645,N_28113,N_28405);
and U29646 (N_29646,N_28894,N_28654);
or U29647 (N_29647,N_28302,N_28006);
nor U29648 (N_29648,N_28443,N_28886);
nand U29649 (N_29649,N_28887,N_28469);
xor U29650 (N_29650,N_28440,N_28875);
or U29651 (N_29651,N_28675,N_28605);
nand U29652 (N_29652,N_28587,N_28273);
nand U29653 (N_29653,N_28526,N_28643);
nor U29654 (N_29654,N_28553,N_28253);
xor U29655 (N_29655,N_28327,N_28417);
and U29656 (N_29656,N_28074,N_28210);
or U29657 (N_29657,N_28708,N_28540);
nor U29658 (N_29658,N_28137,N_28425);
xor U29659 (N_29659,N_28022,N_28426);
or U29660 (N_29660,N_28312,N_28019);
or U29661 (N_29661,N_28151,N_28459);
nor U29662 (N_29662,N_28378,N_28528);
and U29663 (N_29663,N_28341,N_28845);
and U29664 (N_29664,N_28783,N_28644);
xnor U29665 (N_29665,N_28599,N_28656);
nand U29666 (N_29666,N_28155,N_28840);
and U29667 (N_29667,N_28875,N_28343);
nor U29668 (N_29668,N_28676,N_28402);
and U29669 (N_29669,N_28176,N_28105);
or U29670 (N_29670,N_28261,N_28979);
and U29671 (N_29671,N_28937,N_28469);
or U29672 (N_29672,N_28090,N_28409);
or U29673 (N_29673,N_28721,N_28979);
xnor U29674 (N_29674,N_28820,N_28712);
nor U29675 (N_29675,N_28479,N_28141);
nand U29676 (N_29676,N_28819,N_28882);
nand U29677 (N_29677,N_28039,N_28114);
xor U29678 (N_29678,N_28935,N_28495);
or U29679 (N_29679,N_28757,N_28607);
nand U29680 (N_29680,N_28957,N_28995);
or U29681 (N_29681,N_28384,N_28184);
or U29682 (N_29682,N_28308,N_28055);
xor U29683 (N_29683,N_28004,N_28461);
xnor U29684 (N_29684,N_28008,N_28728);
nand U29685 (N_29685,N_28653,N_28802);
or U29686 (N_29686,N_28526,N_28710);
nor U29687 (N_29687,N_28734,N_28249);
nor U29688 (N_29688,N_28944,N_28805);
and U29689 (N_29689,N_28007,N_28147);
nor U29690 (N_29690,N_28093,N_28405);
nor U29691 (N_29691,N_28738,N_28136);
xnor U29692 (N_29692,N_28238,N_28336);
nand U29693 (N_29693,N_28613,N_28188);
or U29694 (N_29694,N_28065,N_28410);
or U29695 (N_29695,N_28749,N_28629);
or U29696 (N_29696,N_28474,N_28305);
nand U29697 (N_29697,N_28572,N_28757);
nor U29698 (N_29698,N_28587,N_28833);
nor U29699 (N_29699,N_28382,N_28293);
nor U29700 (N_29700,N_28077,N_28985);
nand U29701 (N_29701,N_28695,N_28746);
and U29702 (N_29702,N_28360,N_28020);
and U29703 (N_29703,N_28214,N_28035);
or U29704 (N_29704,N_28452,N_28139);
or U29705 (N_29705,N_28847,N_28924);
nor U29706 (N_29706,N_28061,N_28831);
nand U29707 (N_29707,N_28511,N_28745);
nand U29708 (N_29708,N_28378,N_28909);
xor U29709 (N_29709,N_28771,N_28939);
nand U29710 (N_29710,N_28445,N_28544);
or U29711 (N_29711,N_28864,N_28786);
xnor U29712 (N_29712,N_28283,N_28284);
and U29713 (N_29713,N_28621,N_28138);
xnor U29714 (N_29714,N_28978,N_28559);
nor U29715 (N_29715,N_28338,N_28776);
xor U29716 (N_29716,N_28149,N_28628);
or U29717 (N_29717,N_28231,N_28037);
xnor U29718 (N_29718,N_28017,N_28716);
or U29719 (N_29719,N_28676,N_28781);
or U29720 (N_29720,N_28345,N_28757);
nand U29721 (N_29721,N_28626,N_28655);
nand U29722 (N_29722,N_28643,N_28061);
xor U29723 (N_29723,N_28298,N_28118);
nand U29724 (N_29724,N_28197,N_28353);
nor U29725 (N_29725,N_28361,N_28998);
and U29726 (N_29726,N_28958,N_28851);
and U29727 (N_29727,N_28437,N_28319);
nor U29728 (N_29728,N_28271,N_28189);
or U29729 (N_29729,N_28092,N_28726);
xor U29730 (N_29730,N_28203,N_28175);
xor U29731 (N_29731,N_28874,N_28865);
xnor U29732 (N_29732,N_28528,N_28649);
nand U29733 (N_29733,N_28929,N_28181);
nor U29734 (N_29734,N_28768,N_28268);
or U29735 (N_29735,N_28406,N_28298);
nand U29736 (N_29736,N_28229,N_28282);
nand U29737 (N_29737,N_28335,N_28710);
and U29738 (N_29738,N_28558,N_28779);
and U29739 (N_29739,N_28299,N_28872);
or U29740 (N_29740,N_28475,N_28187);
xnor U29741 (N_29741,N_28787,N_28237);
nand U29742 (N_29742,N_28046,N_28440);
nand U29743 (N_29743,N_28143,N_28864);
and U29744 (N_29744,N_28555,N_28812);
nor U29745 (N_29745,N_28905,N_28019);
and U29746 (N_29746,N_28347,N_28641);
xnor U29747 (N_29747,N_28360,N_28065);
or U29748 (N_29748,N_28328,N_28468);
or U29749 (N_29749,N_28310,N_28739);
nor U29750 (N_29750,N_28875,N_28132);
xor U29751 (N_29751,N_28804,N_28879);
nand U29752 (N_29752,N_28950,N_28096);
nor U29753 (N_29753,N_28484,N_28754);
or U29754 (N_29754,N_28854,N_28070);
or U29755 (N_29755,N_28821,N_28311);
or U29756 (N_29756,N_28049,N_28083);
and U29757 (N_29757,N_28747,N_28106);
xnor U29758 (N_29758,N_28326,N_28645);
nand U29759 (N_29759,N_28497,N_28845);
xor U29760 (N_29760,N_28893,N_28515);
or U29761 (N_29761,N_28542,N_28152);
nor U29762 (N_29762,N_28938,N_28425);
and U29763 (N_29763,N_28265,N_28936);
nor U29764 (N_29764,N_28495,N_28031);
nand U29765 (N_29765,N_28571,N_28316);
nand U29766 (N_29766,N_28849,N_28941);
or U29767 (N_29767,N_28303,N_28424);
xor U29768 (N_29768,N_28999,N_28661);
or U29769 (N_29769,N_28733,N_28028);
or U29770 (N_29770,N_28190,N_28975);
or U29771 (N_29771,N_28287,N_28946);
xor U29772 (N_29772,N_28372,N_28876);
and U29773 (N_29773,N_28719,N_28607);
and U29774 (N_29774,N_28830,N_28695);
nor U29775 (N_29775,N_28511,N_28248);
nand U29776 (N_29776,N_28305,N_28038);
xor U29777 (N_29777,N_28432,N_28419);
or U29778 (N_29778,N_28474,N_28108);
nor U29779 (N_29779,N_28720,N_28395);
nand U29780 (N_29780,N_28105,N_28899);
or U29781 (N_29781,N_28438,N_28984);
nand U29782 (N_29782,N_28909,N_28749);
and U29783 (N_29783,N_28907,N_28123);
xor U29784 (N_29784,N_28577,N_28219);
xor U29785 (N_29785,N_28824,N_28489);
xor U29786 (N_29786,N_28339,N_28768);
and U29787 (N_29787,N_28684,N_28382);
or U29788 (N_29788,N_28178,N_28832);
and U29789 (N_29789,N_28821,N_28338);
xnor U29790 (N_29790,N_28400,N_28741);
nand U29791 (N_29791,N_28349,N_28879);
nor U29792 (N_29792,N_28896,N_28495);
or U29793 (N_29793,N_28160,N_28391);
nand U29794 (N_29794,N_28331,N_28746);
xor U29795 (N_29795,N_28105,N_28984);
nor U29796 (N_29796,N_28922,N_28785);
nor U29797 (N_29797,N_28086,N_28601);
nand U29798 (N_29798,N_28111,N_28854);
nand U29799 (N_29799,N_28249,N_28857);
nor U29800 (N_29800,N_28614,N_28837);
nand U29801 (N_29801,N_28943,N_28847);
xnor U29802 (N_29802,N_28177,N_28411);
or U29803 (N_29803,N_28375,N_28616);
and U29804 (N_29804,N_28510,N_28249);
nand U29805 (N_29805,N_28636,N_28352);
xnor U29806 (N_29806,N_28938,N_28686);
nand U29807 (N_29807,N_28423,N_28892);
xor U29808 (N_29808,N_28482,N_28402);
or U29809 (N_29809,N_28938,N_28266);
xnor U29810 (N_29810,N_28299,N_28865);
and U29811 (N_29811,N_28540,N_28514);
or U29812 (N_29812,N_28351,N_28574);
or U29813 (N_29813,N_28946,N_28970);
nor U29814 (N_29814,N_28372,N_28138);
or U29815 (N_29815,N_28105,N_28868);
xor U29816 (N_29816,N_28387,N_28285);
and U29817 (N_29817,N_28590,N_28201);
or U29818 (N_29818,N_28855,N_28622);
nand U29819 (N_29819,N_28366,N_28126);
nand U29820 (N_29820,N_28652,N_28659);
xor U29821 (N_29821,N_28913,N_28498);
or U29822 (N_29822,N_28058,N_28300);
nor U29823 (N_29823,N_28964,N_28744);
xnor U29824 (N_29824,N_28544,N_28343);
and U29825 (N_29825,N_28759,N_28659);
or U29826 (N_29826,N_28576,N_28734);
and U29827 (N_29827,N_28434,N_28782);
or U29828 (N_29828,N_28822,N_28062);
nand U29829 (N_29829,N_28742,N_28915);
and U29830 (N_29830,N_28479,N_28044);
xor U29831 (N_29831,N_28599,N_28817);
or U29832 (N_29832,N_28935,N_28611);
xor U29833 (N_29833,N_28494,N_28653);
or U29834 (N_29834,N_28356,N_28522);
nand U29835 (N_29835,N_28701,N_28362);
and U29836 (N_29836,N_28331,N_28885);
nor U29837 (N_29837,N_28651,N_28004);
or U29838 (N_29838,N_28672,N_28890);
xor U29839 (N_29839,N_28901,N_28898);
and U29840 (N_29840,N_28561,N_28037);
or U29841 (N_29841,N_28746,N_28074);
nand U29842 (N_29842,N_28848,N_28608);
nor U29843 (N_29843,N_28858,N_28284);
nand U29844 (N_29844,N_28276,N_28971);
or U29845 (N_29845,N_28683,N_28183);
nand U29846 (N_29846,N_28785,N_28410);
nor U29847 (N_29847,N_28457,N_28061);
nor U29848 (N_29848,N_28478,N_28898);
xor U29849 (N_29849,N_28473,N_28831);
or U29850 (N_29850,N_28558,N_28928);
xor U29851 (N_29851,N_28366,N_28809);
nand U29852 (N_29852,N_28615,N_28381);
or U29853 (N_29853,N_28160,N_28413);
nor U29854 (N_29854,N_28793,N_28998);
nor U29855 (N_29855,N_28589,N_28412);
and U29856 (N_29856,N_28774,N_28046);
xor U29857 (N_29857,N_28207,N_28558);
xnor U29858 (N_29858,N_28411,N_28084);
or U29859 (N_29859,N_28482,N_28090);
xnor U29860 (N_29860,N_28753,N_28071);
nor U29861 (N_29861,N_28571,N_28345);
xor U29862 (N_29862,N_28380,N_28254);
or U29863 (N_29863,N_28801,N_28995);
nor U29864 (N_29864,N_28061,N_28435);
nand U29865 (N_29865,N_28838,N_28028);
nor U29866 (N_29866,N_28503,N_28376);
or U29867 (N_29867,N_28335,N_28752);
or U29868 (N_29868,N_28073,N_28498);
or U29869 (N_29869,N_28078,N_28794);
nor U29870 (N_29870,N_28762,N_28794);
xnor U29871 (N_29871,N_28244,N_28706);
nor U29872 (N_29872,N_28586,N_28134);
and U29873 (N_29873,N_28640,N_28013);
and U29874 (N_29874,N_28868,N_28000);
nand U29875 (N_29875,N_28247,N_28267);
xnor U29876 (N_29876,N_28158,N_28490);
nand U29877 (N_29877,N_28924,N_28097);
or U29878 (N_29878,N_28735,N_28595);
or U29879 (N_29879,N_28899,N_28686);
xnor U29880 (N_29880,N_28738,N_28085);
or U29881 (N_29881,N_28287,N_28976);
nand U29882 (N_29882,N_28541,N_28815);
nand U29883 (N_29883,N_28471,N_28850);
xnor U29884 (N_29884,N_28306,N_28330);
or U29885 (N_29885,N_28709,N_28246);
and U29886 (N_29886,N_28911,N_28245);
xor U29887 (N_29887,N_28680,N_28332);
nand U29888 (N_29888,N_28652,N_28239);
or U29889 (N_29889,N_28073,N_28015);
or U29890 (N_29890,N_28399,N_28255);
xor U29891 (N_29891,N_28746,N_28864);
and U29892 (N_29892,N_28743,N_28434);
nor U29893 (N_29893,N_28878,N_28998);
xor U29894 (N_29894,N_28162,N_28227);
nor U29895 (N_29895,N_28756,N_28164);
nor U29896 (N_29896,N_28897,N_28880);
and U29897 (N_29897,N_28183,N_28741);
nand U29898 (N_29898,N_28931,N_28648);
nor U29899 (N_29899,N_28346,N_28963);
xor U29900 (N_29900,N_28033,N_28444);
xor U29901 (N_29901,N_28919,N_28635);
nor U29902 (N_29902,N_28253,N_28692);
and U29903 (N_29903,N_28630,N_28039);
and U29904 (N_29904,N_28773,N_28692);
xnor U29905 (N_29905,N_28612,N_28844);
or U29906 (N_29906,N_28258,N_28586);
and U29907 (N_29907,N_28931,N_28659);
nand U29908 (N_29908,N_28271,N_28826);
or U29909 (N_29909,N_28985,N_28536);
or U29910 (N_29910,N_28091,N_28544);
nand U29911 (N_29911,N_28397,N_28540);
or U29912 (N_29912,N_28890,N_28712);
nand U29913 (N_29913,N_28992,N_28902);
and U29914 (N_29914,N_28685,N_28501);
xor U29915 (N_29915,N_28147,N_28645);
and U29916 (N_29916,N_28819,N_28990);
or U29917 (N_29917,N_28025,N_28086);
or U29918 (N_29918,N_28631,N_28509);
nand U29919 (N_29919,N_28832,N_28527);
and U29920 (N_29920,N_28762,N_28472);
xor U29921 (N_29921,N_28082,N_28205);
or U29922 (N_29922,N_28310,N_28443);
nand U29923 (N_29923,N_28343,N_28009);
and U29924 (N_29924,N_28509,N_28617);
nand U29925 (N_29925,N_28827,N_28662);
and U29926 (N_29926,N_28718,N_28663);
xnor U29927 (N_29927,N_28031,N_28443);
xor U29928 (N_29928,N_28135,N_28825);
or U29929 (N_29929,N_28661,N_28237);
nor U29930 (N_29930,N_28215,N_28277);
nor U29931 (N_29931,N_28498,N_28397);
or U29932 (N_29932,N_28643,N_28380);
xnor U29933 (N_29933,N_28100,N_28879);
and U29934 (N_29934,N_28427,N_28692);
nand U29935 (N_29935,N_28670,N_28957);
or U29936 (N_29936,N_28529,N_28004);
and U29937 (N_29937,N_28671,N_28108);
and U29938 (N_29938,N_28238,N_28712);
nor U29939 (N_29939,N_28653,N_28049);
nand U29940 (N_29940,N_28529,N_28907);
or U29941 (N_29941,N_28728,N_28249);
xor U29942 (N_29942,N_28469,N_28145);
nor U29943 (N_29943,N_28180,N_28621);
or U29944 (N_29944,N_28500,N_28165);
and U29945 (N_29945,N_28717,N_28535);
or U29946 (N_29946,N_28764,N_28458);
and U29947 (N_29947,N_28974,N_28580);
xnor U29948 (N_29948,N_28940,N_28697);
xor U29949 (N_29949,N_28356,N_28476);
nand U29950 (N_29950,N_28269,N_28930);
and U29951 (N_29951,N_28469,N_28518);
nand U29952 (N_29952,N_28708,N_28496);
and U29953 (N_29953,N_28420,N_28920);
nor U29954 (N_29954,N_28701,N_28500);
or U29955 (N_29955,N_28551,N_28335);
or U29956 (N_29956,N_28867,N_28214);
xor U29957 (N_29957,N_28161,N_28667);
nand U29958 (N_29958,N_28519,N_28163);
nor U29959 (N_29959,N_28285,N_28646);
xnor U29960 (N_29960,N_28370,N_28459);
nand U29961 (N_29961,N_28230,N_28150);
xor U29962 (N_29962,N_28302,N_28696);
and U29963 (N_29963,N_28699,N_28251);
or U29964 (N_29964,N_28005,N_28764);
nand U29965 (N_29965,N_28410,N_28366);
nor U29966 (N_29966,N_28647,N_28069);
nor U29967 (N_29967,N_28028,N_28334);
nand U29968 (N_29968,N_28767,N_28906);
and U29969 (N_29969,N_28265,N_28059);
or U29970 (N_29970,N_28188,N_28900);
or U29971 (N_29971,N_28832,N_28516);
or U29972 (N_29972,N_28927,N_28527);
nor U29973 (N_29973,N_28366,N_28872);
or U29974 (N_29974,N_28575,N_28615);
and U29975 (N_29975,N_28012,N_28496);
xor U29976 (N_29976,N_28495,N_28536);
or U29977 (N_29977,N_28381,N_28012);
and U29978 (N_29978,N_28233,N_28235);
and U29979 (N_29979,N_28962,N_28415);
or U29980 (N_29980,N_28423,N_28809);
xnor U29981 (N_29981,N_28324,N_28408);
nor U29982 (N_29982,N_28786,N_28086);
nand U29983 (N_29983,N_28954,N_28811);
or U29984 (N_29984,N_28016,N_28198);
and U29985 (N_29985,N_28288,N_28072);
nor U29986 (N_29986,N_28588,N_28572);
or U29987 (N_29987,N_28497,N_28839);
and U29988 (N_29988,N_28810,N_28072);
and U29989 (N_29989,N_28780,N_28525);
nor U29990 (N_29990,N_28405,N_28395);
xnor U29991 (N_29991,N_28457,N_28032);
or U29992 (N_29992,N_28726,N_28169);
xnor U29993 (N_29993,N_28743,N_28972);
or U29994 (N_29994,N_28099,N_28311);
or U29995 (N_29995,N_28318,N_28051);
and U29996 (N_29996,N_28927,N_28317);
nand U29997 (N_29997,N_28958,N_28039);
or U29998 (N_29998,N_28149,N_28758);
nor U29999 (N_29999,N_28489,N_28145);
nand UO_0 (O_0,N_29789,N_29585);
nand UO_1 (O_1,N_29519,N_29674);
nand UO_2 (O_2,N_29084,N_29402);
or UO_3 (O_3,N_29305,N_29625);
nand UO_4 (O_4,N_29110,N_29572);
xnor UO_5 (O_5,N_29273,N_29465);
nand UO_6 (O_6,N_29897,N_29083);
xnor UO_7 (O_7,N_29453,N_29765);
nor UO_8 (O_8,N_29867,N_29731);
and UO_9 (O_9,N_29844,N_29068);
nor UO_10 (O_10,N_29853,N_29104);
nor UO_11 (O_11,N_29445,N_29299);
and UO_12 (O_12,N_29499,N_29406);
or UO_13 (O_13,N_29180,N_29633);
xor UO_14 (O_14,N_29728,N_29944);
nor UO_15 (O_15,N_29065,N_29599);
nor UO_16 (O_16,N_29513,N_29687);
and UO_17 (O_17,N_29602,N_29716);
xnor UO_18 (O_18,N_29972,N_29958);
nor UO_19 (O_19,N_29590,N_29541);
nor UO_20 (O_20,N_29534,N_29912);
or UO_21 (O_21,N_29089,N_29514);
xor UO_22 (O_22,N_29983,N_29381);
xnor UO_23 (O_23,N_29366,N_29531);
and UO_24 (O_24,N_29827,N_29634);
and UO_25 (O_25,N_29031,N_29702);
nor UO_26 (O_26,N_29353,N_29437);
and UO_27 (O_27,N_29303,N_29182);
or UO_28 (O_28,N_29036,N_29883);
xnor UO_29 (O_29,N_29394,N_29492);
nor UO_30 (O_30,N_29521,N_29044);
nand UO_31 (O_31,N_29715,N_29767);
xor UO_32 (O_32,N_29826,N_29420);
and UO_33 (O_33,N_29396,N_29335);
or UO_34 (O_34,N_29977,N_29183);
nand UO_35 (O_35,N_29607,N_29074);
and UO_36 (O_36,N_29734,N_29146);
and UO_37 (O_37,N_29876,N_29236);
and UO_38 (O_38,N_29473,N_29830);
and UO_39 (O_39,N_29120,N_29512);
nor UO_40 (O_40,N_29745,N_29331);
nand UO_41 (O_41,N_29943,N_29309);
nor UO_42 (O_42,N_29247,N_29907);
or UO_43 (O_43,N_29295,N_29004);
xnor UO_44 (O_44,N_29891,N_29707);
nand UO_45 (O_45,N_29987,N_29566);
or UO_46 (O_46,N_29302,N_29153);
xor UO_47 (O_47,N_29352,N_29109);
nor UO_48 (O_48,N_29312,N_29112);
nand UO_49 (O_49,N_29598,N_29538);
xor UO_50 (O_50,N_29685,N_29117);
nor UO_51 (O_51,N_29866,N_29037);
and UO_52 (O_52,N_29306,N_29328);
xor UO_53 (O_53,N_29484,N_29511);
and UO_54 (O_54,N_29547,N_29903);
or UO_55 (O_55,N_29881,N_29025);
nor UO_56 (O_56,N_29859,N_29419);
nand UO_57 (O_57,N_29933,N_29256);
xnor UO_58 (O_58,N_29754,N_29914);
or UO_59 (O_59,N_29479,N_29848);
nand UO_60 (O_60,N_29142,N_29232);
nand UO_61 (O_61,N_29191,N_29285);
and UO_62 (O_62,N_29626,N_29378);
xor UO_63 (O_63,N_29909,N_29532);
nand UO_64 (O_64,N_29087,N_29663);
and UO_65 (O_65,N_29207,N_29748);
nor UO_66 (O_66,N_29758,N_29069);
nor UO_67 (O_67,N_29385,N_29874);
or UO_68 (O_68,N_29121,N_29166);
nand UO_69 (O_69,N_29843,N_29281);
or UO_70 (O_70,N_29054,N_29341);
or UO_71 (O_71,N_29568,N_29583);
nor UO_72 (O_72,N_29497,N_29761);
nor UO_73 (O_73,N_29440,N_29759);
and UO_74 (O_74,N_29934,N_29214);
nand UO_75 (O_75,N_29956,N_29476);
xnor UO_76 (O_76,N_29581,N_29254);
and UO_77 (O_77,N_29670,N_29155);
xnor UO_78 (O_78,N_29710,N_29178);
or UO_79 (O_79,N_29164,N_29321);
nor UO_80 (O_80,N_29355,N_29204);
nand UO_81 (O_81,N_29387,N_29563);
and UO_82 (O_82,N_29475,N_29165);
and UO_83 (O_83,N_29882,N_29560);
xor UO_84 (O_84,N_29092,N_29757);
or UO_85 (O_85,N_29008,N_29222);
nor UO_86 (O_86,N_29549,N_29712);
nor UO_87 (O_87,N_29429,N_29284);
xnor UO_88 (O_88,N_29543,N_29713);
xnor UO_89 (O_89,N_29231,N_29393);
nor UO_90 (O_90,N_29435,N_29949);
and UO_91 (O_91,N_29116,N_29500);
xnor UO_92 (O_92,N_29212,N_29374);
nor UO_93 (O_93,N_29227,N_29668);
nor UO_94 (O_94,N_29265,N_29739);
xor UO_95 (O_95,N_29496,N_29854);
or UO_96 (O_96,N_29550,N_29013);
nand UO_97 (O_97,N_29470,N_29058);
nor UO_98 (O_98,N_29689,N_29539);
or UO_99 (O_99,N_29901,N_29009);
or UO_100 (O_100,N_29007,N_29810);
nand UO_101 (O_101,N_29884,N_29315);
nor UO_102 (O_102,N_29316,N_29151);
xor UO_103 (O_103,N_29570,N_29966);
nor UO_104 (O_104,N_29762,N_29662);
xnor UO_105 (O_105,N_29252,N_29443);
and UO_106 (O_106,N_29965,N_29067);
or UO_107 (O_107,N_29483,N_29923);
or UO_108 (O_108,N_29398,N_29071);
xnor UO_109 (O_109,N_29705,N_29307);
xnor UO_110 (O_110,N_29066,N_29750);
xnor UO_111 (O_111,N_29459,N_29718);
xor UO_112 (O_112,N_29801,N_29082);
nor UO_113 (O_113,N_29509,N_29242);
xor UO_114 (O_114,N_29487,N_29657);
nand UO_115 (O_115,N_29330,N_29641);
xnor UO_116 (O_116,N_29049,N_29928);
or UO_117 (O_117,N_29708,N_29729);
or UO_118 (O_118,N_29384,N_29682);
and UO_119 (O_119,N_29970,N_29170);
nand UO_120 (O_120,N_29442,N_29807);
nand UO_121 (O_121,N_29571,N_29733);
and UO_122 (O_122,N_29535,N_29526);
nor UO_123 (O_123,N_29819,N_29656);
or UO_124 (O_124,N_29413,N_29593);
or UO_125 (O_125,N_29989,N_29565);
xor UO_126 (O_126,N_29371,N_29039);
or UO_127 (O_127,N_29940,N_29474);
or UO_128 (O_128,N_29617,N_29438);
xnor UO_129 (O_129,N_29197,N_29606);
nand UO_130 (O_130,N_29805,N_29720);
xnor UO_131 (O_131,N_29529,N_29399);
nor UO_132 (O_132,N_29177,N_29555);
xnor UO_133 (O_133,N_29169,N_29464);
and UO_134 (O_134,N_29098,N_29589);
xor UO_135 (O_135,N_29900,N_29834);
nand UO_136 (O_136,N_29127,N_29503);
and UO_137 (O_137,N_29119,N_29377);
xor UO_138 (O_138,N_29508,N_29388);
and UO_139 (O_139,N_29821,N_29862);
nor UO_140 (O_140,N_29892,N_29020);
or UO_141 (O_141,N_29246,N_29596);
nor UO_142 (O_142,N_29783,N_29122);
and UO_143 (O_143,N_29213,N_29361);
and UO_144 (O_144,N_29806,N_29404);
or UO_145 (O_145,N_29038,N_29781);
nand UO_146 (O_146,N_29605,N_29665);
nor UO_147 (O_147,N_29160,N_29967);
xnor UO_148 (O_148,N_29224,N_29939);
nand UO_149 (O_149,N_29778,N_29086);
xor UO_150 (O_150,N_29491,N_29623);
and UO_151 (O_151,N_29879,N_29631);
xnor UO_152 (O_152,N_29850,N_29645);
xnor UO_153 (O_153,N_29209,N_29727);
nand UO_154 (O_154,N_29026,N_29017);
nand UO_155 (O_155,N_29426,N_29271);
or UO_156 (O_156,N_29869,N_29988);
and UO_157 (O_157,N_29288,N_29920);
nand UO_158 (O_158,N_29791,N_29875);
nor UO_159 (O_159,N_29911,N_29679);
nand UO_160 (O_160,N_29198,N_29184);
and UO_161 (O_161,N_29863,N_29595);
xor UO_162 (O_162,N_29363,N_29637);
and UO_163 (O_163,N_29005,N_29357);
or UO_164 (O_164,N_29698,N_29370);
or UO_165 (O_165,N_29202,N_29878);
or UO_166 (O_166,N_29811,N_29986);
or UO_167 (O_167,N_29980,N_29975);
xor UO_168 (O_168,N_29671,N_29055);
and UO_169 (O_169,N_29154,N_29741);
or UO_170 (O_170,N_29677,N_29035);
nand UO_171 (O_171,N_29622,N_29090);
nand UO_172 (O_172,N_29383,N_29436);
nor UO_173 (O_173,N_29841,N_29889);
nor UO_174 (O_174,N_29280,N_29612);
nor UO_175 (O_175,N_29235,N_29002);
nand UO_176 (O_176,N_29959,N_29400);
xor UO_177 (O_177,N_29955,N_29592);
nand UO_178 (O_178,N_29651,N_29237);
nor UO_179 (O_179,N_29836,N_29751);
or UO_180 (O_180,N_29888,N_29458);
and UO_181 (O_181,N_29211,N_29486);
nand UO_182 (O_182,N_29382,N_29558);
xor UO_183 (O_183,N_29332,N_29320);
nor UO_184 (O_184,N_29297,N_29991);
nand UO_185 (O_185,N_29048,N_29097);
and UO_186 (O_186,N_29530,N_29032);
xnor UO_187 (O_187,N_29604,N_29011);
xnor UO_188 (O_188,N_29792,N_29769);
nand UO_189 (O_189,N_29998,N_29216);
and UO_190 (O_190,N_29837,N_29638);
xor UO_191 (O_191,N_29194,N_29427);
nand UO_192 (O_192,N_29203,N_29157);
nand UO_193 (O_193,N_29345,N_29618);
nand UO_194 (O_194,N_29014,N_29945);
or UO_195 (O_195,N_29290,N_29283);
or UO_196 (O_196,N_29350,N_29851);
nor UO_197 (O_197,N_29188,N_29027);
or UO_198 (O_198,N_29905,N_29785);
and UO_199 (O_199,N_29999,N_29450);
nand UO_200 (O_200,N_29744,N_29310);
and UO_201 (O_201,N_29372,N_29409);
nor UO_202 (O_202,N_29777,N_29347);
and UO_203 (O_203,N_29106,N_29505);
or UO_204 (O_204,N_29796,N_29922);
nand UO_205 (O_205,N_29343,N_29276);
or UO_206 (O_206,N_29386,N_29747);
or UO_207 (O_207,N_29927,N_29260);
xnor UO_208 (O_208,N_29724,N_29871);
nand UO_209 (O_209,N_29717,N_29646);
nand UO_210 (O_210,N_29910,N_29144);
or UO_211 (O_211,N_29351,N_29093);
nand UO_212 (O_212,N_29323,N_29226);
or UO_213 (O_213,N_29666,N_29775);
and UO_214 (O_214,N_29217,N_29159);
nand UO_215 (O_215,N_29096,N_29449);
or UO_216 (O_216,N_29782,N_29793);
nand UO_217 (O_217,N_29849,N_29610);
xor UO_218 (O_218,N_29737,N_29838);
and UO_219 (O_219,N_29921,N_29193);
and UO_220 (O_220,N_29199,N_29824);
and UO_221 (O_221,N_29076,N_29664);
xnor UO_222 (O_222,N_29858,N_29141);
or UO_223 (O_223,N_29693,N_29375);
or UO_224 (O_224,N_29579,N_29763);
and UO_225 (O_225,N_29825,N_29738);
and UO_226 (O_226,N_29973,N_29251);
nand UO_227 (O_227,N_29131,N_29272);
and UO_228 (O_228,N_29709,N_29932);
xnor UO_229 (O_229,N_29149,N_29636);
or UO_230 (O_230,N_29060,N_29395);
nand UO_231 (O_231,N_29051,N_29522);
nor UO_232 (O_232,N_29424,N_29771);
nand UO_233 (O_233,N_29640,N_29407);
xor UO_234 (O_234,N_29845,N_29723);
and UO_235 (O_235,N_29990,N_29052);
and UO_236 (O_236,N_29814,N_29130);
nand UO_237 (O_237,N_29263,N_29997);
and UO_238 (O_238,N_29033,N_29085);
or UO_239 (O_239,N_29621,N_29412);
nor UO_240 (O_240,N_29803,N_29336);
nand UO_241 (O_241,N_29070,N_29798);
or UO_242 (O_242,N_29174,N_29749);
xnor UO_243 (O_243,N_29576,N_29902);
nand UO_244 (O_244,N_29969,N_29041);
or UO_245 (O_245,N_29894,N_29168);
xnor UO_246 (O_246,N_29773,N_29423);
or UO_247 (O_247,N_29551,N_29012);
nand UO_248 (O_248,N_29971,N_29957);
nand UO_249 (O_249,N_29294,N_29688);
and UO_250 (O_250,N_29896,N_29463);
nor UO_251 (O_251,N_29692,N_29860);
nor UO_252 (O_252,N_29322,N_29886);
or UO_253 (O_253,N_29691,N_29468);
xnor UO_254 (O_254,N_29735,N_29301);
nor UO_255 (O_255,N_29984,N_29397);
nand UO_256 (O_256,N_29802,N_29286);
xor UO_257 (O_257,N_29416,N_29173);
or UO_258 (O_258,N_29003,N_29405);
and UO_259 (O_259,N_29313,N_29015);
and UO_260 (O_260,N_29839,N_29135);
nand UO_261 (O_261,N_29241,N_29954);
nand UO_262 (O_262,N_29552,N_29291);
nand UO_263 (O_263,N_29813,N_29893);
and UO_264 (O_264,N_29118,N_29342);
or UO_265 (O_265,N_29454,N_29078);
and UO_266 (O_266,N_29495,N_29156);
nand UO_267 (O_267,N_29580,N_29392);
or UO_268 (O_268,N_29577,N_29628);
nor UO_269 (O_269,N_29681,N_29644);
nand UO_270 (O_270,N_29061,N_29455);
nand UO_271 (O_271,N_29714,N_29730);
nand UO_272 (O_272,N_29648,N_29652);
nor UO_273 (O_273,N_29201,N_29292);
or UO_274 (O_274,N_29091,N_29196);
nand UO_275 (O_275,N_29578,N_29358);
or UO_276 (O_276,N_29359,N_29546);
nor UO_277 (O_277,N_29161,N_29000);
and UO_278 (O_278,N_29278,N_29139);
and UO_279 (O_279,N_29208,N_29129);
nor UO_280 (O_280,N_29620,N_29390);
nand UO_281 (O_281,N_29616,N_29536);
and UO_282 (O_282,N_29525,N_29334);
xnor UO_283 (O_283,N_29527,N_29123);
or UO_284 (O_284,N_29561,N_29653);
nand UO_285 (O_285,N_29742,N_29953);
nor UO_286 (O_286,N_29079,N_29433);
xnor UO_287 (O_287,N_29770,N_29736);
or UO_288 (O_288,N_29573,N_29456);
and UO_289 (O_289,N_29482,N_29772);
nand UO_290 (O_290,N_29132,N_29700);
nand UO_291 (O_291,N_29311,N_29963);
or UO_292 (O_292,N_29072,N_29138);
nor UO_293 (O_293,N_29057,N_29516);
nor UO_294 (O_294,N_29308,N_29143);
or UO_295 (O_295,N_29029,N_29947);
xor UO_296 (O_296,N_29215,N_29642);
and UO_297 (O_297,N_29829,N_29439);
nand UO_298 (O_298,N_29134,N_29812);
nor UO_299 (O_299,N_29873,N_29554);
xor UO_300 (O_300,N_29993,N_29533);
and UO_301 (O_301,N_29895,N_29441);
xnor UO_302 (O_302,N_29167,N_29187);
and UO_303 (O_303,N_29504,N_29995);
or UO_304 (O_304,N_29111,N_29600);
or UO_305 (O_305,N_29417,N_29979);
or UO_306 (O_306,N_29403,N_29948);
nor UO_307 (O_307,N_29520,N_29507);
nand UO_308 (O_308,N_29324,N_29186);
or UO_309 (O_309,N_29815,N_29823);
nand UO_310 (O_310,N_29447,N_29494);
nor UO_311 (O_311,N_29107,N_29658);
nor UO_312 (O_312,N_29243,N_29269);
nand UO_313 (O_313,N_29220,N_29150);
or UO_314 (O_314,N_29799,N_29746);
or UO_315 (O_315,N_29906,N_29899);
xnor UO_316 (O_316,N_29006,N_29282);
xnor UO_317 (O_317,N_29887,N_29696);
or UO_318 (O_318,N_29175,N_29063);
nand UO_319 (O_319,N_29654,N_29635);
nand UO_320 (O_320,N_29961,N_29101);
nand UO_321 (O_321,N_29128,N_29695);
and UO_322 (O_322,N_29794,N_29711);
or UO_323 (O_323,N_29189,N_29376);
or UO_324 (O_324,N_29152,N_29493);
or UO_325 (O_325,N_29472,N_29672);
nor UO_326 (O_326,N_29103,N_29304);
xor UO_327 (O_327,N_29701,N_29266);
or UO_328 (O_328,N_29978,N_29743);
xor UO_329 (O_329,N_29451,N_29205);
or UO_330 (O_330,N_29289,N_29756);
nand UO_331 (O_331,N_29591,N_29466);
nand UO_332 (O_332,N_29223,N_29938);
nor UO_333 (O_333,N_29753,N_29348);
and UO_334 (O_334,N_29619,N_29726);
nor UO_335 (O_335,N_29075,N_29239);
or UO_336 (O_336,N_29485,N_29327);
nor UO_337 (O_337,N_29904,N_29515);
nand UO_338 (O_338,N_29721,N_29820);
or UO_339 (O_339,N_29608,N_29976);
xor UO_340 (O_340,N_29210,N_29171);
or UO_341 (O_341,N_29982,N_29542);
nand UO_342 (O_342,N_29916,N_29809);
xnor UO_343 (O_343,N_29544,N_29462);
and UO_344 (O_344,N_29469,N_29680);
nand UO_345 (O_345,N_29800,N_29996);
or UO_346 (O_346,N_29234,N_29244);
xor UO_347 (O_347,N_29941,N_29125);
nor UO_348 (O_348,N_29339,N_29362);
or UO_349 (O_349,N_29857,N_29444);
and UO_350 (O_350,N_29597,N_29100);
nor UO_351 (O_351,N_29010,N_29760);
nor UO_352 (O_352,N_29267,N_29557);
nor UO_353 (O_353,N_29669,N_29457);
xnor UO_354 (O_354,N_29262,N_29019);
and UO_355 (O_355,N_29338,N_29414);
and UO_356 (O_356,N_29056,N_29408);
xnor UO_357 (O_357,N_29962,N_29569);
xor UO_358 (O_358,N_29936,N_29917);
nand UO_359 (O_359,N_29919,N_29163);
or UO_360 (O_360,N_29425,N_29890);
or UO_361 (O_361,N_29360,N_29258);
xor UO_362 (O_362,N_29981,N_29298);
xnor UO_363 (O_363,N_29248,N_29719);
nand UO_364 (O_364,N_29113,N_29176);
nor UO_365 (O_365,N_29471,N_29575);
nand UO_366 (O_366,N_29562,N_29181);
nor UO_367 (O_367,N_29985,N_29524);
nor UO_368 (O_368,N_29279,N_29864);
and UO_369 (O_369,N_29686,N_29856);
or UO_370 (O_370,N_29831,N_29219);
nor UO_371 (O_371,N_29461,N_29059);
nand UO_372 (O_372,N_29105,N_29564);
and UO_373 (O_373,N_29601,N_29460);
and UO_374 (O_374,N_29629,N_29992);
nand UO_375 (O_375,N_29832,N_29683);
or UO_376 (O_376,N_29942,N_29274);
xnor UO_377 (O_377,N_29929,N_29255);
nand UO_378 (O_378,N_29797,N_29047);
or UO_379 (O_379,N_29567,N_29639);
nor UO_380 (O_380,N_29808,N_29379);
xor UO_381 (O_381,N_29421,N_29314);
and UO_382 (O_382,N_29344,N_29603);
and UO_383 (O_383,N_29488,N_29268);
or UO_384 (O_384,N_29221,N_29935);
or UO_385 (O_385,N_29594,N_29667);
xor UO_386 (O_386,N_29245,N_29676);
or UO_387 (O_387,N_29467,N_29647);
or UO_388 (O_388,N_29369,N_29249);
nand UO_389 (O_389,N_29994,N_29478);
xnor UO_390 (O_390,N_29287,N_29477);
and UO_391 (O_391,N_29960,N_29296);
nand UO_392 (O_392,N_29852,N_29264);
nand UO_393 (O_393,N_29088,N_29365);
nand UO_394 (O_394,N_29452,N_29974);
xor UO_395 (O_395,N_29432,N_29545);
xnor UO_396 (O_396,N_29001,N_29489);
nor UO_397 (O_397,N_29584,N_29018);
nand UO_398 (O_398,N_29430,N_29043);
nor UO_399 (O_399,N_29816,N_29659);
and UO_400 (O_400,N_29835,N_29480);
xnor UO_401 (O_401,N_29023,N_29660);
xnor UO_402 (O_402,N_29077,N_29846);
or UO_403 (O_403,N_29586,N_29136);
or UO_404 (O_404,N_29418,N_29333);
or UO_405 (O_405,N_29225,N_29779);
nor UO_406 (O_406,N_29053,N_29588);
xor UO_407 (O_407,N_29776,N_29795);
nand UO_408 (O_408,N_29913,N_29349);
nand UO_409 (O_409,N_29162,N_29095);
nand UO_410 (O_410,N_29930,N_29238);
nor UO_411 (O_411,N_29021,N_29675);
xor UO_412 (O_412,N_29609,N_29300);
or UO_413 (O_413,N_29915,N_29102);
or UO_414 (O_414,N_29885,N_29764);
or UO_415 (O_415,N_29126,N_29732);
nor UO_416 (O_416,N_29655,N_29045);
or UO_417 (O_417,N_29788,N_29368);
nand UO_418 (O_418,N_29137,N_29818);
xnor UO_419 (O_419,N_29179,N_29034);
xor UO_420 (O_420,N_29627,N_29050);
xor UO_421 (O_421,N_29080,N_29148);
nand UO_422 (O_422,N_29926,N_29073);
or UO_423 (O_423,N_29704,N_29448);
nand UO_424 (O_424,N_29337,N_29250);
or UO_425 (O_425,N_29861,N_29556);
xor UO_426 (O_426,N_29523,N_29356);
nand UO_427 (O_427,N_29952,N_29872);
xor UO_428 (O_428,N_29540,N_29725);
nand UO_429 (O_429,N_29918,N_29703);
xnor UO_430 (O_430,N_29946,N_29632);
nor UO_431 (O_431,N_29804,N_29253);
or UO_432 (O_432,N_29615,N_29172);
nand UO_433 (O_433,N_29855,N_29042);
or UO_434 (O_434,N_29510,N_29833);
nor UO_435 (O_435,N_29822,N_29030);
xnor UO_436 (O_436,N_29229,N_29261);
xnor UO_437 (O_437,N_29446,N_29099);
nand UO_438 (O_438,N_29190,N_29147);
nand UO_439 (O_439,N_29022,N_29094);
nor UO_440 (O_440,N_29502,N_29329);
xnor UO_441 (O_441,N_29192,N_29373);
xnor UO_442 (O_442,N_29115,N_29548);
nand UO_443 (O_443,N_29145,N_29401);
nor UO_444 (O_444,N_29828,N_29880);
nand UO_445 (O_445,N_29790,N_29650);
nand UO_446 (O_446,N_29694,N_29755);
xnor UO_447 (O_447,N_29140,N_29410);
xor UO_448 (O_448,N_29752,N_29870);
or UO_449 (O_449,N_29699,N_29490);
nand UO_450 (O_450,N_29517,N_29501);
nand UO_451 (O_451,N_29422,N_29740);
nor UO_452 (O_452,N_29865,N_29951);
and UO_453 (O_453,N_29518,N_29124);
nand UO_454 (O_454,N_29624,N_29766);
nor UO_455 (O_455,N_29431,N_29200);
or UO_456 (O_456,N_29706,N_29908);
and UO_457 (O_457,N_29206,N_29481);
xor UO_458 (O_458,N_29937,N_29380);
xnor UO_459 (O_459,N_29024,N_29228);
xor UO_460 (O_460,N_29649,N_29319);
nand UO_461 (O_461,N_29780,N_29768);
xor UO_462 (O_462,N_29233,N_29678);
nor UO_463 (O_463,N_29877,N_29925);
xor UO_464 (O_464,N_29411,N_29690);
nor UO_465 (O_465,N_29195,N_29697);
xnor UO_466 (O_466,N_29354,N_29259);
nand UO_467 (O_467,N_29661,N_29275);
nor UO_468 (O_468,N_29218,N_29062);
xor UO_469 (O_469,N_29964,N_29787);
nand UO_470 (O_470,N_29643,N_29326);
or UO_471 (O_471,N_29270,N_29046);
nand UO_472 (O_472,N_29114,N_29931);
xnor UO_473 (O_473,N_29230,N_29293);
nor UO_474 (O_474,N_29817,N_29574);
nor UO_475 (O_475,N_29684,N_29968);
and UO_476 (O_476,N_29614,N_29277);
xor UO_477 (O_477,N_29318,N_29924);
or UO_478 (O_478,N_29840,N_29847);
nor UO_479 (O_479,N_29391,N_29364);
nand UO_480 (O_480,N_29950,N_29537);
xnor UO_481 (O_481,N_29784,N_29028);
xor UO_482 (O_482,N_29587,N_29428);
xor UO_483 (O_483,N_29498,N_29040);
xnor UO_484 (O_484,N_29389,N_29774);
or UO_485 (O_485,N_29064,N_29325);
nand UO_486 (O_486,N_29158,N_29367);
nand UO_487 (O_487,N_29611,N_29613);
nand UO_488 (O_488,N_29553,N_29346);
xnor UO_489 (O_489,N_29868,N_29133);
or UO_490 (O_490,N_29108,N_29630);
nor UO_491 (O_491,N_29016,N_29722);
or UO_492 (O_492,N_29240,N_29434);
or UO_493 (O_493,N_29415,N_29559);
nor UO_494 (O_494,N_29081,N_29898);
xor UO_495 (O_495,N_29582,N_29317);
or UO_496 (O_496,N_29673,N_29340);
and UO_497 (O_497,N_29842,N_29257);
nor UO_498 (O_498,N_29185,N_29506);
or UO_499 (O_499,N_29528,N_29786);
nand UO_500 (O_500,N_29634,N_29904);
or UO_501 (O_501,N_29277,N_29280);
nand UO_502 (O_502,N_29200,N_29104);
nand UO_503 (O_503,N_29520,N_29353);
and UO_504 (O_504,N_29523,N_29453);
or UO_505 (O_505,N_29881,N_29238);
nand UO_506 (O_506,N_29745,N_29044);
or UO_507 (O_507,N_29995,N_29241);
nor UO_508 (O_508,N_29627,N_29169);
or UO_509 (O_509,N_29610,N_29277);
nand UO_510 (O_510,N_29062,N_29265);
or UO_511 (O_511,N_29535,N_29474);
and UO_512 (O_512,N_29305,N_29136);
or UO_513 (O_513,N_29315,N_29576);
nor UO_514 (O_514,N_29159,N_29376);
and UO_515 (O_515,N_29237,N_29677);
xnor UO_516 (O_516,N_29742,N_29299);
nor UO_517 (O_517,N_29228,N_29031);
or UO_518 (O_518,N_29022,N_29473);
and UO_519 (O_519,N_29848,N_29624);
xor UO_520 (O_520,N_29361,N_29864);
xor UO_521 (O_521,N_29976,N_29578);
xor UO_522 (O_522,N_29850,N_29567);
xor UO_523 (O_523,N_29658,N_29063);
nor UO_524 (O_524,N_29267,N_29134);
nand UO_525 (O_525,N_29925,N_29884);
nor UO_526 (O_526,N_29353,N_29938);
nor UO_527 (O_527,N_29620,N_29124);
nand UO_528 (O_528,N_29134,N_29120);
xnor UO_529 (O_529,N_29477,N_29693);
nand UO_530 (O_530,N_29384,N_29309);
nor UO_531 (O_531,N_29646,N_29600);
nor UO_532 (O_532,N_29384,N_29104);
xor UO_533 (O_533,N_29018,N_29113);
and UO_534 (O_534,N_29487,N_29049);
and UO_535 (O_535,N_29219,N_29088);
nor UO_536 (O_536,N_29087,N_29507);
xor UO_537 (O_537,N_29718,N_29661);
xor UO_538 (O_538,N_29035,N_29186);
or UO_539 (O_539,N_29561,N_29684);
nor UO_540 (O_540,N_29739,N_29573);
nand UO_541 (O_541,N_29257,N_29426);
or UO_542 (O_542,N_29111,N_29209);
nor UO_543 (O_543,N_29011,N_29284);
nor UO_544 (O_544,N_29061,N_29877);
nand UO_545 (O_545,N_29342,N_29156);
nand UO_546 (O_546,N_29844,N_29632);
and UO_547 (O_547,N_29801,N_29755);
nand UO_548 (O_548,N_29366,N_29865);
xnor UO_549 (O_549,N_29348,N_29556);
or UO_550 (O_550,N_29730,N_29435);
or UO_551 (O_551,N_29925,N_29411);
or UO_552 (O_552,N_29772,N_29348);
and UO_553 (O_553,N_29946,N_29151);
nand UO_554 (O_554,N_29886,N_29015);
and UO_555 (O_555,N_29828,N_29401);
nor UO_556 (O_556,N_29680,N_29983);
xor UO_557 (O_557,N_29708,N_29744);
nand UO_558 (O_558,N_29288,N_29489);
and UO_559 (O_559,N_29858,N_29114);
xor UO_560 (O_560,N_29515,N_29832);
and UO_561 (O_561,N_29948,N_29270);
nor UO_562 (O_562,N_29459,N_29982);
nand UO_563 (O_563,N_29476,N_29880);
or UO_564 (O_564,N_29146,N_29160);
or UO_565 (O_565,N_29323,N_29481);
or UO_566 (O_566,N_29172,N_29492);
and UO_567 (O_567,N_29111,N_29751);
nor UO_568 (O_568,N_29989,N_29003);
and UO_569 (O_569,N_29577,N_29065);
nor UO_570 (O_570,N_29771,N_29248);
nor UO_571 (O_571,N_29120,N_29687);
or UO_572 (O_572,N_29550,N_29797);
nor UO_573 (O_573,N_29597,N_29587);
xnor UO_574 (O_574,N_29355,N_29734);
or UO_575 (O_575,N_29761,N_29830);
nand UO_576 (O_576,N_29175,N_29458);
nor UO_577 (O_577,N_29291,N_29405);
and UO_578 (O_578,N_29823,N_29461);
xor UO_579 (O_579,N_29290,N_29225);
nor UO_580 (O_580,N_29511,N_29017);
xor UO_581 (O_581,N_29657,N_29200);
nand UO_582 (O_582,N_29449,N_29454);
and UO_583 (O_583,N_29105,N_29882);
xnor UO_584 (O_584,N_29131,N_29207);
xnor UO_585 (O_585,N_29916,N_29709);
and UO_586 (O_586,N_29003,N_29314);
xor UO_587 (O_587,N_29115,N_29784);
and UO_588 (O_588,N_29856,N_29143);
xnor UO_589 (O_589,N_29705,N_29814);
and UO_590 (O_590,N_29983,N_29027);
nor UO_591 (O_591,N_29676,N_29435);
xnor UO_592 (O_592,N_29101,N_29319);
and UO_593 (O_593,N_29898,N_29235);
xnor UO_594 (O_594,N_29822,N_29518);
nand UO_595 (O_595,N_29388,N_29046);
nor UO_596 (O_596,N_29252,N_29354);
xnor UO_597 (O_597,N_29109,N_29960);
nand UO_598 (O_598,N_29318,N_29166);
or UO_599 (O_599,N_29596,N_29426);
nand UO_600 (O_600,N_29877,N_29689);
nor UO_601 (O_601,N_29402,N_29401);
or UO_602 (O_602,N_29745,N_29386);
or UO_603 (O_603,N_29611,N_29903);
or UO_604 (O_604,N_29659,N_29152);
nand UO_605 (O_605,N_29884,N_29352);
xor UO_606 (O_606,N_29194,N_29449);
or UO_607 (O_607,N_29875,N_29785);
and UO_608 (O_608,N_29731,N_29953);
nor UO_609 (O_609,N_29542,N_29819);
nor UO_610 (O_610,N_29753,N_29266);
xnor UO_611 (O_611,N_29255,N_29868);
and UO_612 (O_612,N_29503,N_29638);
and UO_613 (O_613,N_29157,N_29403);
and UO_614 (O_614,N_29842,N_29779);
nor UO_615 (O_615,N_29439,N_29065);
xnor UO_616 (O_616,N_29282,N_29113);
nor UO_617 (O_617,N_29243,N_29873);
and UO_618 (O_618,N_29957,N_29191);
xnor UO_619 (O_619,N_29881,N_29964);
nor UO_620 (O_620,N_29506,N_29422);
and UO_621 (O_621,N_29363,N_29400);
and UO_622 (O_622,N_29804,N_29839);
or UO_623 (O_623,N_29061,N_29030);
and UO_624 (O_624,N_29011,N_29287);
or UO_625 (O_625,N_29878,N_29915);
xnor UO_626 (O_626,N_29613,N_29944);
and UO_627 (O_627,N_29967,N_29753);
and UO_628 (O_628,N_29775,N_29296);
or UO_629 (O_629,N_29633,N_29292);
nand UO_630 (O_630,N_29436,N_29565);
xnor UO_631 (O_631,N_29152,N_29298);
and UO_632 (O_632,N_29098,N_29669);
or UO_633 (O_633,N_29871,N_29920);
nand UO_634 (O_634,N_29426,N_29059);
xnor UO_635 (O_635,N_29223,N_29585);
xnor UO_636 (O_636,N_29198,N_29285);
xnor UO_637 (O_637,N_29261,N_29314);
nor UO_638 (O_638,N_29617,N_29718);
or UO_639 (O_639,N_29318,N_29937);
or UO_640 (O_640,N_29803,N_29136);
or UO_641 (O_641,N_29201,N_29734);
or UO_642 (O_642,N_29542,N_29334);
nand UO_643 (O_643,N_29915,N_29236);
and UO_644 (O_644,N_29021,N_29620);
nor UO_645 (O_645,N_29481,N_29809);
and UO_646 (O_646,N_29930,N_29741);
nand UO_647 (O_647,N_29751,N_29367);
nand UO_648 (O_648,N_29639,N_29354);
and UO_649 (O_649,N_29837,N_29319);
nor UO_650 (O_650,N_29133,N_29813);
and UO_651 (O_651,N_29274,N_29037);
nand UO_652 (O_652,N_29016,N_29100);
and UO_653 (O_653,N_29496,N_29442);
nand UO_654 (O_654,N_29540,N_29802);
nand UO_655 (O_655,N_29409,N_29696);
nor UO_656 (O_656,N_29828,N_29556);
xor UO_657 (O_657,N_29390,N_29988);
and UO_658 (O_658,N_29596,N_29677);
xnor UO_659 (O_659,N_29810,N_29831);
nand UO_660 (O_660,N_29542,N_29806);
and UO_661 (O_661,N_29808,N_29775);
xnor UO_662 (O_662,N_29445,N_29230);
or UO_663 (O_663,N_29999,N_29098);
and UO_664 (O_664,N_29655,N_29168);
or UO_665 (O_665,N_29852,N_29390);
or UO_666 (O_666,N_29361,N_29420);
nor UO_667 (O_667,N_29348,N_29380);
and UO_668 (O_668,N_29318,N_29981);
nor UO_669 (O_669,N_29747,N_29014);
nand UO_670 (O_670,N_29017,N_29122);
or UO_671 (O_671,N_29009,N_29376);
and UO_672 (O_672,N_29662,N_29191);
nor UO_673 (O_673,N_29071,N_29819);
nand UO_674 (O_674,N_29702,N_29937);
or UO_675 (O_675,N_29979,N_29717);
nor UO_676 (O_676,N_29479,N_29576);
xnor UO_677 (O_677,N_29697,N_29242);
xor UO_678 (O_678,N_29428,N_29638);
or UO_679 (O_679,N_29368,N_29870);
nor UO_680 (O_680,N_29014,N_29831);
nand UO_681 (O_681,N_29155,N_29952);
and UO_682 (O_682,N_29349,N_29464);
and UO_683 (O_683,N_29343,N_29718);
nor UO_684 (O_684,N_29706,N_29933);
nor UO_685 (O_685,N_29348,N_29211);
nand UO_686 (O_686,N_29192,N_29388);
xor UO_687 (O_687,N_29331,N_29269);
nor UO_688 (O_688,N_29531,N_29338);
nor UO_689 (O_689,N_29028,N_29983);
nor UO_690 (O_690,N_29719,N_29198);
nor UO_691 (O_691,N_29239,N_29579);
or UO_692 (O_692,N_29218,N_29068);
nand UO_693 (O_693,N_29965,N_29708);
or UO_694 (O_694,N_29076,N_29079);
and UO_695 (O_695,N_29088,N_29948);
xnor UO_696 (O_696,N_29258,N_29954);
nand UO_697 (O_697,N_29870,N_29332);
or UO_698 (O_698,N_29919,N_29807);
nor UO_699 (O_699,N_29256,N_29257);
xor UO_700 (O_700,N_29116,N_29563);
or UO_701 (O_701,N_29924,N_29095);
xnor UO_702 (O_702,N_29023,N_29830);
nand UO_703 (O_703,N_29408,N_29261);
and UO_704 (O_704,N_29609,N_29477);
nand UO_705 (O_705,N_29527,N_29734);
nor UO_706 (O_706,N_29865,N_29301);
nor UO_707 (O_707,N_29489,N_29271);
and UO_708 (O_708,N_29091,N_29620);
and UO_709 (O_709,N_29104,N_29325);
nand UO_710 (O_710,N_29900,N_29820);
xnor UO_711 (O_711,N_29896,N_29255);
xnor UO_712 (O_712,N_29316,N_29147);
nor UO_713 (O_713,N_29579,N_29609);
nand UO_714 (O_714,N_29594,N_29234);
nand UO_715 (O_715,N_29683,N_29569);
and UO_716 (O_716,N_29251,N_29731);
xnor UO_717 (O_717,N_29666,N_29929);
xor UO_718 (O_718,N_29506,N_29181);
nand UO_719 (O_719,N_29399,N_29266);
nor UO_720 (O_720,N_29603,N_29130);
nand UO_721 (O_721,N_29514,N_29596);
and UO_722 (O_722,N_29252,N_29535);
nand UO_723 (O_723,N_29468,N_29996);
xor UO_724 (O_724,N_29944,N_29810);
nor UO_725 (O_725,N_29261,N_29558);
and UO_726 (O_726,N_29451,N_29024);
xor UO_727 (O_727,N_29944,N_29174);
and UO_728 (O_728,N_29190,N_29647);
xor UO_729 (O_729,N_29826,N_29281);
or UO_730 (O_730,N_29647,N_29479);
xor UO_731 (O_731,N_29404,N_29637);
nor UO_732 (O_732,N_29312,N_29763);
or UO_733 (O_733,N_29927,N_29954);
xnor UO_734 (O_734,N_29493,N_29032);
xnor UO_735 (O_735,N_29543,N_29604);
xnor UO_736 (O_736,N_29448,N_29558);
or UO_737 (O_737,N_29743,N_29165);
and UO_738 (O_738,N_29978,N_29515);
xor UO_739 (O_739,N_29875,N_29171);
xor UO_740 (O_740,N_29883,N_29831);
xor UO_741 (O_741,N_29654,N_29389);
nor UO_742 (O_742,N_29417,N_29192);
and UO_743 (O_743,N_29361,N_29437);
or UO_744 (O_744,N_29532,N_29343);
nor UO_745 (O_745,N_29400,N_29756);
and UO_746 (O_746,N_29128,N_29079);
nor UO_747 (O_747,N_29859,N_29588);
nor UO_748 (O_748,N_29795,N_29240);
xor UO_749 (O_749,N_29948,N_29210);
nor UO_750 (O_750,N_29361,N_29742);
nor UO_751 (O_751,N_29350,N_29305);
and UO_752 (O_752,N_29506,N_29709);
or UO_753 (O_753,N_29460,N_29689);
nand UO_754 (O_754,N_29640,N_29670);
and UO_755 (O_755,N_29499,N_29655);
nand UO_756 (O_756,N_29674,N_29599);
or UO_757 (O_757,N_29586,N_29403);
xnor UO_758 (O_758,N_29842,N_29272);
and UO_759 (O_759,N_29071,N_29499);
xnor UO_760 (O_760,N_29542,N_29673);
nand UO_761 (O_761,N_29583,N_29532);
xnor UO_762 (O_762,N_29393,N_29987);
or UO_763 (O_763,N_29938,N_29345);
nand UO_764 (O_764,N_29196,N_29199);
and UO_765 (O_765,N_29684,N_29667);
xnor UO_766 (O_766,N_29244,N_29083);
or UO_767 (O_767,N_29852,N_29452);
xor UO_768 (O_768,N_29812,N_29567);
nand UO_769 (O_769,N_29284,N_29881);
and UO_770 (O_770,N_29018,N_29217);
nor UO_771 (O_771,N_29061,N_29344);
nand UO_772 (O_772,N_29164,N_29378);
and UO_773 (O_773,N_29068,N_29119);
xor UO_774 (O_774,N_29435,N_29116);
and UO_775 (O_775,N_29907,N_29354);
xor UO_776 (O_776,N_29039,N_29140);
nand UO_777 (O_777,N_29995,N_29623);
xnor UO_778 (O_778,N_29313,N_29954);
nor UO_779 (O_779,N_29910,N_29555);
and UO_780 (O_780,N_29469,N_29299);
nor UO_781 (O_781,N_29534,N_29339);
or UO_782 (O_782,N_29355,N_29152);
and UO_783 (O_783,N_29895,N_29610);
and UO_784 (O_784,N_29557,N_29449);
xnor UO_785 (O_785,N_29325,N_29624);
and UO_786 (O_786,N_29679,N_29152);
nor UO_787 (O_787,N_29984,N_29761);
or UO_788 (O_788,N_29952,N_29227);
xnor UO_789 (O_789,N_29730,N_29657);
or UO_790 (O_790,N_29064,N_29246);
nor UO_791 (O_791,N_29667,N_29374);
nor UO_792 (O_792,N_29465,N_29565);
and UO_793 (O_793,N_29058,N_29708);
and UO_794 (O_794,N_29849,N_29395);
or UO_795 (O_795,N_29217,N_29135);
xnor UO_796 (O_796,N_29786,N_29516);
or UO_797 (O_797,N_29085,N_29776);
xor UO_798 (O_798,N_29306,N_29848);
xnor UO_799 (O_799,N_29982,N_29174);
nor UO_800 (O_800,N_29339,N_29463);
nor UO_801 (O_801,N_29788,N_29093);
xnor UO_802 (O_802,N_29627,N_29494);
xnor UO_803 (O_803,N_29863,N_29626);
xor UO_804 (O_804,N_29663,N_29668);
nor UO_805 (O_805,N_29625,N_29500);
xnor UO_806 (O_806,N_29057,N_29931);
nand UO_807 (O_807,N_29794,N_29073);
xnor UO_808 (O_808,N_29763,N_29957);
xnor UO_809 (O_809,N_29343,N_29595);
nor UO_810 (O_810,N_29277,N_29312);
nand UO_811 (O_811,N_29073,N_29642);
and UO_812 (O_812,N_29841,N_29850);
nand UO_813 (O_813,N_29632,N_29798);
nor UO_814 (O_814,N_29822,N_29493);
and UO_815 (O_815,N_29403,N_29915);
or UO_816 (O_816,N_29466,N_29659);
nand UO_817 (O_817,N_29484,N_29084);
xnor UO_818 (O_818,N_29404,N_29318);
or UO_819 (O_819,N_29769,N_29788);
or UO_820 (O_820,N_29946,N_29741);
nand UO_821 (O_821,N_29894,N_29186);
nand UO_822 (O_822,N_29320,N_29419);
nor UO_823 (O_823,N_29632,N_29198);
xor UO_824 (O_824,N_29270,N_29478);
nor UO_825 (O_825,N_29361,N_29243);
nor UO_826 (O_826,N_29721,N_29578);
xnor UO_827 (O_827,N_29110,N_29353);
and UO_828 (O_828,N_29800,N_29164);
or UO_829 (O_829,N_29805,N_29897);
nor UO_830 (O_830,N_29332,N_29063);
nand UO_831 (O_831,N_29961,N_29924);
or UO_832 (O_832,N_29420,N_29440);
or UO_833 (O_833,N_29309,N_29320);
or UO_834 (O_834,N_29367,N_29283);
xnor UO_835 (O_835,N_29415,N_29450);
nor UO_836 (O_836,N_29843,N_29339);
nor UO_837 (O_837,N_29812,N_29915);
xor UO_838 (O_838,N_29013,N_29245);
or UO_839 (O_839,N_29721,N_29380);
or UO_840 (O_840,N_29004,N_29555);
xnor UO_841 (O_841,N_29267,N_29123);
nand UO_842 (O_842,N_29039,N_29127);
and UO_843 (O_843,N_29037,N_29298);
and UO_844 (O_844,N_29667,N_29784);
or UO_845 (O_845,N_29044,N_29055);
nand UO_846 (O_846,N_29434,N_29371);
xor UO_847 (O_847,N_29118,N_29602);
xnor UO_848 (O_848,N_29026,N_29883);
nand UO_849 (O_849,N_29939,N_29341);
and UO_850 (O_850,N_29985,N_29328);
nor UO_851 (O_851,N_29940,N_29418);
and UO_852 (O_852,N_29794,N_29441);
or UO_853 (O_853,N_29110,N_29655);
nand UO_854 (O_854,N_29658,N_29770);
xor UO_855 (O_855,N_29952,N_29056);
xnor UO_856 (O_856,N_29935,N_29275);
or UO_857 (O_857,N_29413,N_29058);
or UO_858 (O_858,N_29900,N_29396);
nor UO_859 (O_859,N_29119,N_29945);
nor UO_860 (O_860,N_29005,N_29838);
or UO_861 (O_861,N_29820,N_29234);
and UO_862 (O_862,N_29536,N_29412);
xor UO_863 (O_863,N_29879,N_29947);
xor UO_864 (O_864,N_29161,N_29536);
nor UO_865 (O_865,N_29565,N_29844);
nand UO_866 (O_866,N_29665,N_29236);
nor UO_867 (O_867,N_29961,N_29219);
nand UO_868 (O_868,N_29875,N_29573);
or UO_869 (O_869,N_29284,N_29327);
nand UO_870 (O_870,N_29073,N_29617);
xnor UO_871 (O_871,N_29347,N_29120);
xor UO_872 (O_872,N_29428,N_29516);
xor UO_873 (O_873,N_29238,N_29602);
or UO_874 (O_874,N_29699,N_29483);
and UO_875 (O_875,N_29234,N_29419);
nor UO_876 (O_876,N_29038,N_29941);
and UO_877 (O_877,N_29410,N_29186);
and UO_878 (O_878,N_29438,N_29337);
xor UO_879 (O_879,N_29410,N_29001);
nor UO_880 (O_880,N_29004,N_29566);
nand UO_881 (O_881,N_29655,N_29299);
xnor UO_882 (O_882,N_29402,N_29589);
nand UO_883 (O_883,N_29432,N_29142);
and UO_884 (O_884,N_29129,N_29901);
xnor UO_885 (O_885,N_29508,N_29972);
xnor UO_886 (O_886,N_29546,N_29454);
nor UO_887 (O_887,N_29343,N_29407);
nor UO_888 (O_888,N_29693,N_29202);
xnor UO_889 (O_889,N_29761,N_29221);
and UO_890 (O_890,N_29493,N_29855);
or UO_891 (O_891,N_29186,N_29141);
nand UO_892 (O_892,N_29058,N_29232);
and UO_893 (O_893,N_29581,N_29399);
xor UO_894 (O_894,N_29567,N_29809);
or UO_895 (O_895,N_29145,N_29330);
or UO_896 (O_896,N_29345,N_29547);
or UO_897 (O_897,N_29763,N_29693);
and UO_898 (O_898,N_29890,N_29519);
and UO_899 (O_899,N_29008,N_29036);
nand UO_900 (O_900,N_29012,N_29426);
or UO_901 (O_901,N_29597,N_29636);
nand UO_902 (O_902,N_29938,N_29434);
and UO_903 (O_903,N_29180,N_29910);
nand UO_904 (O_904,N_29747,N_29820);
nor UO_905 (O_905,N_29180,N_29611);
nor UO_906 (O_906,N_29856,N_29352);
and UO_907 (O_907,N_29786,N_29343);
or UO_908 (O_908,N_29700,N_29872);
xor UO_909 (O_909,N_29347,N_29707);
nor UO_910 (O_910,N_29112,N_29918);
xnor UO_911 (O_911,N_29106,N_29275);
nor UO_912 (O_912,N_29214,N_29381);
nor UO_913 (O_913,N_29401,N_29323);
nor UO_914 (O_914,N_29759,N_29730);
and UO_915 (O_915,N_29783,N_29833);
nand UO_916 (O_916,N_29835,N_29610);
nor UO_917 (O_917,N_29197,N_29069);
nor UO_918 (O_918,N_29714,N_29811);
and UO_919 (O_919,N_29935,N_29126);
and UO_920 (O_920,N_29385,N_29497);
or UO_921 (O_921,N_29111,N_29161);
or UO_922 (O_922,N_29784,N_29942);
and UO_923 (O_923,N_29354,N_29353);
or UO_924 (O_924,N_29613,N_29469);
nor UO_925 (O_925,N_29330,N_29081);
xor UO_926 (O_926,N_29819,N_29111);
nand UO_927 (O_927,N_29766,N_29075);
and UO_928 (O_928,N_29971,N_29189);
nand UO_929 (O_929,N_29053,N_29883);
xor UO_930 (O_930,N_29408,N_29102);
and UO_931 (O_931,N_29341,N_29533);
nand UO_932 (O_932,N_29003,N_29925);
xnor UO_933 (O_933,N_29230,N_29338);
or UO_934 (O_934,N_29614,N_29039);
or UO_935 (O_935,N_29461,N_29245);
nor UO_936 (O_936,N_29898,N_29442);
xnor UO_937 (O_937,N_29271,N_29239);
xnor UO_938 (O_938,N_29329,N_29382);
xnor UO_939 (O_939,N_29206,N_29283);
xor UO_940 (O_940,N_29740,N_29228);
and UO_941 (O_941,N_29490,N_29833);
or UO_942 (O_942,N_29624,N_29754);
nor UO_943 (O_943,N_29450,N_29306);
nand UO_944 (O_944,N_29348,N_29056);
and UO_945 (O_945,N_29935,N_29233);
nand UO_946 (O_946,N_29801,N_29462);
xnor UO_947 (O_947,N_29784,N_29907);
or UO_948 (O_948,N_29169,N_29591);
nand UO_949 (O_949,N_29689,N_29152);
xnor UO_950 (O_950,N_29462,N_29413);
nor UO_951 (O_951,N_29383,N_29492);
or UO_952 (O_952,N_29987,N_29688);
or UO_953 (O_953,N_29187,N_29419);
nand UO_954 (O_954,N_29674,N_29377);
or UO_955 (O_955,N_29664,N_29338);
nand UO_956 (O_956,N_29010,N_29726);
or UO_957 (O_957,N_29787,N_29376);
and UO_958 (O_958,N_29800,N_29047);
nor UO_959 (O_959,N_29977,N_29205);
and UO_960 (O_960,N_29115,N_29862);
xnor UO_961 (O_961,N_29099,N_29157);
xor UO_962 (O_962,N_29037,N_29547);
nand UO_963 (O_963,N_29683,N_29821);
and UO_964 (O_964,N_29046,N_29312);
xnor UO_965 (O_965,N_29522,N_29833);
and UO_966 (O_966,N_29800,N_29254);
nand UO_967 (O_967,N_29369,N_29418);
and UO_968 (O_968,N_29841,N_29219);
or UO_969 (O_969,N_29975,N_29521);
xnor UO_970 (O_970,N_29939,N_29465);
or UO_971 (O_971,N_29539,N_29799);
xor UO_972 (O_972,N_29960,N_29511);
and UO_973 (O_973,N_29065,N_29507);
and UO_974 (O_974,N_29697,N_29379);
or UO_975 (O_975,N_29652,N_29808);
or UO_976 (O_976,N_29388,N_29845);
and UO_977 (O_977,N_29174,N_29616);
nand UO_978 (O_978,N_29632,N_29838);
and UO_979 (O_979,N_29990,N_29661);
nand UO_980 (O_980,N_29310,N_29732);
and UO_981 (O_981,N_29933,N_29671);
or UO_982 (O_982,N_29474,N_29274);
and UO_983 (O_983,N_29834,N_29650);
nand UO_984 (O_984,N_29334,N_29024);
nand UO_985 (O_985,N_29930,N_29088);
or UO_986 (O_986,N_29873,N_29691);
or UO_987 (O_987,N_29189,N_29062);
xor UO_988 (O_988,N_29813,N_29035);
xnor UO_989 (O_989,N_29172,N_29362);
nand UO_990 (O_990,N_29159,N_29872);
nor UO_991 (O_991,N_29071,N_29452);
nand UO_992 (O_992,N_29962,N_29200);
or UO_993 (O_993,N_29193,N_29715);
nand UO_994 (O_994,N_29239,N_29084);
and UO_995 (O_995,N_29268,N_29658);
nand UO_996 (O_996,N_29578,N_29608);
nor UO_997 (O_997,N_29238,N_29860);
and UO_998 (O_998,N_29186,N_29875);
and UO_999 (O_999,N_29376,N_29213);
nand UO_1000 (O_1000,N_29875,N_29997);
and UO_1001 (O_1001,N_29036,N_29255);
nor UO_1002 (O_1002,N_29367,N_29123);
xnor UO_1003 (O_1003,N_29035,N_29079);
nand UO_1004 (O_1004,N_29622,N_29125);
or UO_1005 (O_1005,N_29315,N_29304);
xnor UO_1006 (O_1006,N_29820,N_29334);
nand UO_1007 (O_1007,N_29144,N_29816);
and UO_1008 (O_1008,N_29692,N_29431);
or UO_1009 (O_1009,N_29206,N_29942);
and UO_1010 (O_1010,N_29495,N_29732);
nor UO_1011 (O_1011,N_29661,N_29204);
nand UO_1012 (O_1012,N_29021,N_29924);
xor UO_1013 (O_1013,N_29238,N_29417);
and UO_1014 (O_1014,N_29986,N_29989);
nand UO_1015 (O_1015,N_29839,N_29765);
and UO_1016 (O_1016,N_29374,N_29491);
xnor UO_1017 (O_1017,N_29516,N_29040);
nor UO_1018 (O_1018,N_29691,N_29665);
and UO_1019 (O_1019,N_29689,N_29203);
nor UO_1020 (O_1020,N_29903,N_29019);
or UO_1021 (O_1021,N_29937,N_29060);
nor UO_1022 (O_1022,N_29039,N_29286);
xor UO_1023 (O_1023,N_29415,N_29743);
nor UO_1024 (O_1024,N_29686,N_29134);
nand UO_1025 (O_1025,N_29508,N_29349);
nand UO_1026 (O_1026,N_29715,N_29249);
nand UO_1027 (O_1027,N_29537,N_29611);
or UO_1028 (O_1028,N_29904,N_29313);
xnor UO_1029 (O_1029,N_29364,N_29337);
and UO_1030 (O_1030,N_29389,N_29328);
nand UO_1031 (O_1031,N_29268,N_29864);
and UO_1032 (O_1032,N_29478,N_29697);
nand UO_1033 (O_1033,N_29441,N_29651);
and UO_1034 (O_1034,N_29583,N_29323);
or UO_1035 (O_1035,N_29753,N_29423);
nor UO_1036 (O_1036,N_29263,N_29274);
and UO_1037 (O_1037,N_29794,N_29388);
nand UO_1038 (O_1038,N_29428,N_29364);
or UO_1039 (O_1039,N_29657,N_29459);
or UO_1040 (O_1040,N_29002,N_29987);
or UO_1041 (O_1041,N_29992,N_29256);
or UO_1042 (O_1042,N_29168,N_29689);
or UO_1043 (O_1043,N_29958,N_29837);
xor UO_1044 (O_1044,N_29342,N_29462);
xnor UO_1045 (O_1045,N_29781,N_29255);
or UO_1046 (O_1046,N_29433,N_29454);
xor UO_1047 (O_1047,N_29579,N_29253);
and UO_1048 (O_1048,N_29560,N_29476);
and UO_1049 (O_1049,N_29984,N_29634);
nor UO_1050 (O_1050,N_29025,N_29928);
or UO_1051 (O_1051,N_29984,N_29033);
nand UO_1052 (O_1052,N_29385,N_29550);
xnor UO_1053 (O_1053,N_29042,N_29447);
nand UO_1054 (O_1054,N_29202,N_29688);
nor UO_1055 (O_1055,N_29413,N_29053);
or UO_1056 (O_1056,N_29656,N_29006);
xor UO_1057 (O_1057,N_29467,N_29434);
nor UO_1058 (O_1058,N_29967,N_29646);
nor UO_1059 (O_1059,N_29651,N_29678);
xnor UO_1060 (O_1060,N_29288,N_29974);
xor UO_1061 (O_1061,N_29972,N_29007);
or UO_1062 (O_1062,N_29525,N_29400);
xnor UO_1063 (O_1063,N_29182,N_29810);
nor UO_1064 (O_1064,N_29681,N_29465);
nor UO_1065 (O_1065,N_29451,N_29905);
nand UO_1066 (O_1066,N_29445,N_29219);
nor UO_1067 (O_1067,N_29461,N_29704);
xnor UO_1068 (O_1068,N_29335,N_29765);
or UO_1069 (O_1069,N_29257,N_29776);
nand UO_1070 (O_1070,N_29915,N_29950);
nor UO_1071 (O_1071,N_29039,N_29009);
nor UO_1072 (O_1072,N_29042,N_29129);
nand UO_1073 (O_1073,N_29473,N_29497);
or UO_1074 (O_1074,N_29257,N_29677);
nand UO_1075 (O_1075,N_29351,N_29079);
or UO_1076 (O_1076,N_29625,N_29866);
nand UO_1077 (O_1077,N_29629,N_29862);
nand UO_1078 (O_1078,N_29440,N_29136);
nor UO_1079 (O_1079,N_29213,N_29828);
xnor UO_1080 (O_1080,N_29235,N_29062);
nor UO_1081 (O_1081,N_29078,N_29842);
and UO_1082 (O_1082,N_29898,N_29954);
and UO_1083 (O_1083,N_29089,N_29840);
xnor UO_1084 (O_1084,N_29131,N_29625);
or UO_1085 (O_1085,N_29265,N_29699);
nor UO_1086 (O_1086,N_29681,N_29560);
and UO_1087 (O_1087,N_29821,N_29534);
nor UO_1088 (O_1088,N_29920,N_29893);
xnor UO_1089 (O_1089,N_29771,N_29551);
nor UO_1090 (O_1090,N_29077,N_29124);
xor UO_1091 (O_1091,N_29927,N_29268);
xnor UO_1092 (O_1092,N_29325,N_29352);
or UO_1093 (O_1093,N_29182,N_29683);
nand UO_1094 (O_1094,N_29282,N_29031);
or UO_1095 (O_1095,N_29638,N_29045);
or UO_1096 (O_1096,N_29920,N_29472);
xor UO_1097 (O_1097,N_29402,N_29791);
nand UO_1098 (O_1098,N_29577,N_29760);
nand UO_1099 (O_1099,N_29773,N_29718);
or UO_1100 (O_1100,N_29148,N_29942);
nand UO_1101 (O_1101,N_29389,N_29354);
nor UO_1102 (O_1102,N_29053,N_29052);
and UO_1103 (O_1103,N_29858,N_29393);
xnor UO_1104 (O_1104,N_29937,N_29487);
nand UO_1105 (O_1105,N_29233,N_29317);
xor UO_1106 (O_1106,N_29505,N_29170);
xnor UO_1107 (O_1107,N_29191,N_29559);
nor UO_1108 (O_1108,N_29724,N_29461);
or UO_1109 (O_1109,N_29720,N_29662);
or UO_1110 (O_1110,N_29079,N_29409);
and UO_1111 (O_1111,N_29858,N_29555);
nor UO_1112 (O_1112,N_29408,N_29665);
nand UO_1113 (O_1113,N_29824,N_29032);
nor UO_1114 (O_1114,N_29716,N_29019);
nor UO_1115 (O_1115,N_29409,N_29535);
xor UO_1116 (O_1116,N_29119,N_29872);
or UO_1117 (O_1117,N_29222,N_29385);
xnor UO_1118 (O_1118,N_29885,N_29748);
and UO_1119 (O_1119,N_29726,N_29417);
and UO_1120 (O_1120,N_29161,N_29879);
or UO_1121 (O_1121,N_29393,N_29590);
nand UO_1122 (O_1122,N_29170,N_29423);
nor UO_1123 (O_1123,N_29157,N_29670);
and UO_1124 (O_1124,N_29444,N_29288);
nand UO_1125 (O_1125,N_29383,N_29182);
or UO_1126 (O_1126,N_29058,N_29469);
nor UO_1127 (O_1127,N_29686,N_29377);
nand UO_1128 (O_1128,N_29722,N_29977);
nand UO_1129 (O_1129,N_29036,N_29616);
nor UO_1130 (O_1130,N_29005,N_29576);
or UO_1131 (O_1131,N_29239,N_29308);
and UO_1132 (O_1132,N_29070,N_29956);
nor UO_1133 (O_1133,N_29795,N_29942);
xor UO_1134 (O_1134,N_29220,N_29688);
nor UO_1135 (O_1135,N_29430,N_29945);
or UO_1136 (O_1136,N_29453,N_29121);
and UO_1137 (O_1137,N_29717,N_29234);
xor UO_1138 (O_1138,N_29958,N_29626);
xnor UO_1139 (O_1139,N_29794,N_29442);
or UO_1140 (O_1140,N_29942,N_29782);
xor UO_1141 (O_1141,N_29711,N_29422);
or UO_1142 (O_1142,N_29628,N_29205);
nand UO_1143 (O_1143,N_29450,N_29661);
or UO_1144 (O_1144,N_29218,N_29883);
and UO_1145 (O_1145,N_29654,N_29644);
and UO_1146 (O_1146,N_29355,N_29260);
and UO_1147 (O_1147,N_29608,N_29633);
nor UO_1148 (O_1148,N_29929,N_29687);
nor UO_1149 (O_1149,N_29743,N_29766);
nor UO_1150 (O_1150,N_29436,N_29147);
xor UO_1151 (O_1151,N_29773,N_29398);
or UO_1152 (O_1152,N_29590,N_29549);
nor UO_1153 (O_1153,N_29569,N_29552);
xnor UO_1154 (O_1154,N_29750,N_29970);
nor UO_1155 (O_1155,N_29959,N_29639);
nand UO_1156 (O_1156,N_29515,N_29754);
or UO_1157 (O_1157,N_29148,N_29116);
and UO_1158 (O_1158,N_29045,N_29348);
or UO_1159 (O_1159,N_29159,N_29890);
xnor UO_1160 (O_1160,N_29167,N_29782);
and UO_1161 (O_1161,N_29078,N_29991);
nand UO_1162 (O_1162,N_29680,N_29711);
or UO_1163 (O_1163,N_29421,N_29495);
nand UO_1164 (O_1164,N_29601,N_29716);
xor UO_1165 (O_1165,N_29857,N_29436);
xor UO_1166 (O_1166,N_29341,N_29020);
xor UO_1167 (O_1167,N_29074,N_29137);
xor UO_1168 (O_1168,N_29792,N_29984);
xnor UO_1169 (O_1169,N_29931,N_29157);
and UO_1170 (O_1170,N_29547,N_29535);
or UO_1171 (O_1171,N_29718,N_29378);
xor UO_1172 (O_1172,N_29603,N_29655);
xnor UO_1173 (O_1173,N_29137,N_29804);
or UO_1174 (O_1174,N_29903,N_29237);
nand UO_1175 (O_1175,N_29379,N_29085);
or UO_1176 (O_1176,N_29470,N_29646);
nand UO_1177 (O_1177,N_29015,N_29392);
nand UO_1178 (O_1178,N_29104,N_29570);
and UO_1179 (O_1179,N_29443,N_29851);
or UO_1180 (O_1180,N_29009,N_29962);
xor UO_1181 (O_1181,N_29376,N_29304);
xor UO_1182 (O_1182,N_29900,N_29328);
nor UO_1183 (O_1183,N_29871,N_29405);
nand UO_1184 (O_1184,N_29628,N_29648);
and UO_1185 (O_1185,N_29360,N_29497);
xnor UO_1186 (O_1186,N_29484,N_29622);
and UO_1187 (O_1187,N_29337,N_29802);
or UO_1188 (O_1188,N_29117,N_29369);
nor UO_1189 (O_1189,N_29239,N_29585);
nor UO_1190 (O_1190,N_29210,N_29563);
nand UO_1191 (O_1191,N_29025,N_29996);
and UO_1192 (O_1192,N_29329,N_29916);
xor UO_1193 (O_1193,N_29435,N_29652);
and UO_1194 (O_1194,N_29364,N_29380);
nor UO_1195 (O_1195,N_29608,N_29999);
xor UO_1196 (O_1196,N_29374,N_29222);
xor UO_1197 (O_1197,N_29275,N_29905);
nand UO_1198 (O_1198,N_29347,N_29108);
and UO_1199 (O_1199,N_29357,N_29058);
or UO_1200 (O_1200,N_29796,N_29437);
xor UO_1201 (O_1201,N_29579,N_29278);
nor UO_1202 (O_1202,N_29957,N_29759);
nor UO_1203 (O_1203,N_29330,N_29039);
nor UO_1204 (O_1204,N_29422,N_29350);
nor UO_1205 (O_1205,N_29040,N_29120);
or UO_1206 (O_1206,N_29943,N_29353);
nand UO_1207 (O_1207,N_29844,N_29418);
and UO_1208 (O_1208,N_29860,N_29967);
xor UO_1209 (O_1209,N_29555,N_29500);
nand UO_1210 (O_1210,N_29481,N_29782);
and UO_1211 (O_1211,N_29056,N_29827);
nor UO_1212 (O_1212,N_29809,N_29202);
nor UO_1213 (O_1213,N_29833,N_29850);
xor UO_1214 (O_1214,N_29810,N_29816);
nand UO_1215 (O_1215,N_29401,N_29896);
and UO_1216 (O_1216,N_29542,N_29989);
and UO_1217 (O_1217,N_29270,N_29365);
nor UO_1218 (O_1218,N_29567,N_29289);
nor UO_1219 (O_1219,N_29470,N_29462);
and UO_1220 (O_1220,N_29103,N_29444);
xnor UO_1221 (O_1221,N_29215,N_29265);
xor UO_1222 (O_1222,N_29786,N_29739);
nand UO_1223 (O_1223,N_29416,N_29283);
xor UO_1224 (O_1224,N_29864,N_29053);
nand UO_1225 (O_1225,N_29163,N_29622);
nor UO_1226 (O_1226,N_29268,N_29072);
and UO_1227 (O_1227,N_29601,N_29274);
and UO_1228 (O_1228,N_29344,N_29266);
nand UO_1229 (O_1229,N_29992,N_29895);
or UO_1230 (O_1230,N_29695,N_29971);
and UO_1231 (O_1231,N_29348,N_29510);
xor UO_1232 (O_1232,N_29104,N_29957);
nand UO_1233 (O_1233,N_29169,N_29748);
nand UO_1234 (O_1234,N_29519,N_29773);
or UO_1235 (O_1235,N_29932,N_29012);
xnor UO_1236 (O_1236,N_29389,N_29293);
or UO_1237 (O_1237,N_29575,N_29236);
or UO_1238 (O_1238,N_29662,N_29017);
nand UO_1239 (O_1239,N_29400,N_29589);
nand UO_1240 (O_1240,N_29180,N_29338);
nand UO_1241 (O_1241,N_29607,N_29365);
or UO_1242 (O_1242,N_29396,N_29110);
nand UO_1243 (O_1243,N_29184,N_29107);
nand UO_1244 (O_1244,N_29520,N_29259);
and UO_1245 (O_1245,N_29123,N_29906);
nor UO_1246 (O_1246,N_29777,N_29198);
nor UO_1247 (O_1247,N_29390,N_29292);
nor UO_1248 (O_1248,N_29326,N_29190);
xor UO_1249 (O_1249,N_29387,N_29867);
nand UO_1250 (O_1250,N_29539,N_29557);
nor UO_1251 (O_1251,N_29307,N_29868);
nor UO_1252 (O_1252,N_29274,N_29066);
nor UO_1253 (O_1253,N_29162,N_29125);
or UO_1254 (O_1254,N_29024,N_29747);
xor UO_1255 (O_1255,N_29392,N_29672);
or UO_1256 (O_1256,N_29031,N_29730);
and UO_1257 (O_1257,N_29882,N_29265);
and UO_1258 (O_1258,N_29617,N_29101);
or UO_1259 (O_1259,N_29907,N_29971);
nor UO_1260 (O_1260,N_29127,N_29652);
nand UO_1261 (O_1261,N_29231,N_29015);
nand UO_1262 (O_1262,N_29086,N_29702);
nand UO_1263 (O_1263,N_29082,N_29059);
xor UO_1264 (O_1264,N_29199,N_29647);
or UO_1265 (O_1265,N_29244,N_29922);
and UO_1266 (O_1266,N_29810,N_29017);
nand UO_1267 (O_1267,N_29462,N_29490);
nand UO_1268 (O_1268,N_29894,N_29613);
and UO_1269 (O_1269,N_29118,N_29206);
and UO_1270 (O_1270,N_29654,N_29396);
xor UO_1271 (O_1271,N_29046,N_29529);
nor UO_1272 (O_1272,N_29494,N_29625);
xnor UO_1273 (O_1273,N_29851,N_29206);
xnor UO_1274 (O_1274,N_29143,N_29623);
and UO_1275 (O_1275,N_29885,N_29753);
and UO_1276 (O_1276,N_29563,N_29957);
and UO_1277 (O_1277,N_29659,N_29465);
and UO_1278 (O_1278,N_29563,N_29660);
nor UO_1279 (O_1279,N_29730,N_29612);
nand UO_1280 (O_1280,N_29253,N_29715);
nor UO_1281 (O_1281,N_29081,N_29262);
and UO_1282 (O_1282,N_29385,N_29153);
nor UO_1283 (O_1283,N_29808,N_29871);
and UO_1284 (O_1284,N_29347,N_29215);
and UO_1285 (O_1285,N_29623,N_29475);
and UO_1286 (O_1286,N_29774,N_29996);
nor UO_1287 (O_1287,N_29786,N_29085);
and UO_1288 (O_1288,N_29053,N_29127);
nand UO_1289 (O_1289,N_29068,N_29637);
nand UO_1290 (O_1290,N_29585,N_29978);
nor UO_1291 (O_1291,N_29272,N_29782);
and UO_1292 (O_1292,N_29304,N_29431);
nand UO_1293 (O_1293,N_29217,N_29759);
or UO_1294 (O_1294,N_29053,N_29503);
or UO_1295 (O_1295,N_29433,N_29322);
and UO_1296 (O_1296,N_29909,N_29914);
or UO_1297 (O_1297,N_29602,N_29272);
nand UO_1298 (O_1298,N_29891,N_29887);
xor UO_1299 (O_1299,N_29143,N_29174);
and UO_1300 (O_1300,N_29172,N_29612);
nand UO_1301 (O_1301,N_29952,N_29980);
and UO_1302 (O_1302,N_29899,N_29534);
or UO_1303 (O_1303,N_29462,N_29689);
and UO_1304 (O_1304,N_29631,N_29370);
or UO_1305 (O_1305,N_29703,N_29510);
or UO_1306 (O_1306,N_29871,N_29296);
nand UO_1307 (O_1307,N_29801,N_29151);
and UO_1308 (O_1308,N_29146,N_29054);
nor UO_1309 (O_1309,N_29255,N_29981);
nor UO_1310 (O_1310,N_29243,N_29893);
nand UO_1311 (O_1311,N_29268,N_29535);
nor UO_1312 (O_1312,N_29988,N_29811);
xor UO_1313 (O_1313,N_29874,N_29403);
and UO_1314 (O_1314,N_29414,N_29172);
and UO_1315 (O_1315,N_29051,N_29290);
or UO_1316 (O_1316,N_29163,N_29021);
and UO_1317 (O_1317,N_29611,N_29547);
nand UO_1318 (O_1318,N_29695,N_29179);
and UO_1319 (O_1319,N_29196,N_29991);
nand UO_1320 (O_1320,N_29923,N_29153);
and UO_1321 (O_1321,N_29486,N_29051);
or UO_1322 (O_1322,N_29547,N_29118);
nand UO_1323 (O_1323,N_29459,N_29210);
nand UO_1324 (O_1324,N_29459,N_29819);
and UO_1325 (O_1325,N_29881,N_29113);
nor UO_1326 (O_1326,N_29416,N_29313);
nand UO_1327 (O_1327,N_29491,N_29031);
and UO_1328 (O_1328,N_29551,N_29903);
and UO_1329 (O_1329,N_29951,N_29584);
or UO_1330 (O_1330,N_29600,N_29862);
or UO_1331 (O_1331,N_29667,N_29816);
xor UO_1332 (O_1332,N_29257,N_29290);
nand UO_1333 (O_1333,N_29002,N_29869);
nor UO_1334 (O_1334,N_29366,N_29257);
nor UO_1335 (O_1335,N_29136,N_29173);
nand UO_1336 (O_1336,N_29378,N_29268);
nand UO_1337 (O_1337,N_29568,N_29725);
xor UO_1338 (O_1338,N_29404,N_29278);
nor UO_1339 (O_1339,N_29597,N_29631);
nor UO_1340 (O_1340,N_29565,N_29238);
xor UO_1341 (O_1341,N_29768,N_29182);
or UO_1342 (O_1342,N_29112,N_29256);
xor UO_1343 (O_1343,N_29325,N_29771);
nor UO_1344 (O_1344,N_29061,N_29555);
xor UO_1345 (O_1345,N_29211,N_29245);
or UO_1346 (O_1346,N_29504,N_29636);
nor UO_1347 (O_1347,N_29233,N_29048);
xnor UO_1348 (O_1348,N_29893,N_29621);
nor UO_1349 (O_1349,N_29320,N_29274);
xnor UO_1350 (O_1350,N_29562,N_29141);
or UO_1351 (O_1351,N_29333,N_29364);
nand UO_1352 (O_1352,N_29277,N_29518);
nand UO_1353 (O_1353,N_29395,N_29442);
nand UO_1354 (O_1354,N_29470,N_29236);
xnor UO_1355 (O_1355,N_29011,N_29374);
nor UO_1356 (O_1356,N_29584,N_29723);
xor UO_1357 (O_1357,N_29534,N_29920);
nand UO_1358 (O_1358,N_29722,N_29042);
and UO_1359 (O_1359,N_29681,N_29263);
or UO_1360 (O_1360,N_29243,N_29270);
or UO_1361 (O_1361,N_29517,N_29956);
nor UO_1362 (O_1362,N_29687,N_29090);
and UO_1363 (O_1363,N_29337,N_29040);
nor UO_1364 (O_1364,N_29954,N_29968);
and UO_1365 (O_1365,N_29188,N_29050);
xor UO_1366 (O_1366,N_29151,N_29855);
xor UO_1367 (O_1367,N_29067,N_29455);
or UO_1368 (O_1368,N_29695,N_29456);
xnor UO_1369 (O_1369,N_29408,N_29896);
or UO_1370 (O_1370,N_29740,N_29702);
xnor UO_1371 (O_1371,N_29245,N_29728);
and UO_1372 (O_1372,N_29587,N_29956);
nor UO_1373 (O_1373,N_29564,N_29352);
or UO_1374 (O_1374,N_29352,N_29992);
nor UO_1375 (O_1375,N_29948,N_29292);
nand UO_1376 (O_1376,N_29191,N_29343);
xor UO_1377 (O_1377,N_29569,N_29440);
nor UO_1378 (O_1378,N_29711,N_29036);
nor UO_1379 (O_1379,N_29150,N_29133);
nand UO_1380 (O_1380,N_29497,N_29080);
and UO_1381 (O_1381,N_29771,N_29313);
xor UO_1382 (O_1382,N_29974,N_29183);
nor UO_1383 (O_1383,N_29405,N_29357);
and UO_1384 (O_1384,N_29089,N_29301);
and UO_1385 (O_1385,N_29829,N_29924);
nand UO_1386 (O_1386,N_29331,N_29008);
nand UO_1387 (O_1387,N_29994,N_29697);
nand UO_1388 (O_1388,N_29208,N_29744);
and UO_1389 (O_1389,N_29436,N_29146);
and UO_1390 (O_1390,N_29520,N_29979);
or UO_1391 (O_1391,N_29477,N_29150);
and UO_1392 (O_1392,N_29803,N_29145);
xor UO_1393 (O_1393,N_29161,N_29572);
and UO_1394 (O_1394,N_29472,N_29565);
nand UO_1395 (O_1395,N_29262,N_29412);
xnor UO_1396 (O_1396,N_29468,N_29982);
nand UO_1397 (O_1397,N_29819,N_29788);
and UO_1398 (O_1398,N_29117,N_29881);
xor UO_1399 (O_1399,N_29919,N_29151);
nand UO_1400 (O_1400,N_29787,N_29900);
xnor UO_1401 (O_1401,N_29101,N_29766);
or UO_1402 (O_1402,N_29569,N_29816);
nand UO_1403 (O_1403,N_29509,N_29347);
and UO_1404 (O_1404,N_29692,N_29774);
and UO_1405 (O_1405,N_29827,N_29657);
nand UO_1406 (O_1406,N_29479,N_29456);
and UO_1407 (O_1407,N_29017,N_29571);
or UO_1408 (O_1408,N_29278,N_29623);
nor UO_1409 (O_1409,N_29801,N_29236);
and UO_1410 (O_1410,N_29509,N_29253);
xnor UO_1411 (O_1411,N_29543,N_29644);
or UO_1412 (O_1412,N_29164,N_29185);
or UO_1413 (O_1413,N_29286,N_29057);
nand UO_1414 (O_1414,N_29088,N_29060);
nor UO_1415 (O_1415,N_29198,N_29084);
xnor UO_1416 (O_1416,N_29846,N_29799);
nand UO_1417 (O_1417,N_29433,N_29757);
xor UO_1418 (O_1418,N_29519,N_29181);
nor UO_1419 (O_1419,N_29163,N_29090);
nor UO_1420 (O_1420,N_29893,N_29887);
xnor UO_1421 (O_1421,N_29180,N_29883);
nand UO_1422 (O_1422,N_29585,N_29092);
nor UO_1423 (O_1423,N_29026,N_29581);
xor UO_1424 (O_1424,N_29340,N_29770);
nand UO_1425 (O_1425,N_29443,N_29871);
nor UO_1426 (O_1426,N_29916,N_29109);
and UO_1427 (O_1427,N_29388,N_29237);
and UO_1428 (O_1428,N_29318,N_29825);
xor UO_1429 (O_1429,N_29049,N_29110);
xor UO_1430 (O_1430,N_29307,N_29946);
nor UO_1431 (O_1431,N_29439,N_29434);
or UO_1432 (O_1432,N_29529,N_29759);
and UO_1433 (O_1433,N_29895,N_29689);
or UO_1434 (O_1434,N_29558,N_29938);
xor UO_1435 (O_1435,N_29647,N_29972);
or UO_1436 (O_1436,N_29009,N_29893);
and UO_1437 (O_1437,N_29702,N_29980);
and UO_1438 (O_1438,N_29634,N_29166);
xor UO_1439 (O_1439,N_29305,N_29587);
nor UO_1440 (O_1440,N_29717,N_29769);
xnor UO_1441 (O_1441,N_29355,N_29923);
nand UO_1442 (O_1442,N_29693,N_29158);
xnor UO_1443 (O_1443,N_29773,N_29301);
and UO_1444 (O_1444,N_29890,N_29493);
xnor UO_1445 (O_1445,N_29523,N_29148);
xnor UO_1446 (O_1446,N_29181,N_29105);
or UO_1447 (O_1447,N_29217,N_29670);
nand UO_1448 (O_1448,N_29457,N_29681);
nand UO_1449 (O_1449,N_29279,N_29599);
nand UO_1450 (O_1450,N_29585,N_29888);
nand UO_1451 (O_1451,N_29953,N_29461);
xor UO_1452 (O_1452,N_29483,N_29080);
and UO_1453 (O_1453,N_29552,N_29838);
nand UO_1454 (O_1454,N_29662,N_29393);
or UO_1455 (O_1455,N_29607,N_29541);
nand UO_1456 (O_1456,N_29878,N_29067);
nor UO_1457 (O_1457,N_29042,N_29734);
or UO_1458 (O_1458,N_29267,N_29509);
nand UO_1459 (O_1459,N_29720,N_29620);
nand UO_1460 (O_1460,N_29468,N_29815);
nor UO_1461 (O_1461,N_29746,N_29787);
nand UO_1462 (O_1462,N_29055,N_29246);
nand UO_1463 (O_1463,N_29962,N_29715);
nand UO_1464 (O_1464,N_29773,N_29563);
or UO_1465 (O_1465,N_29146,N_29434);
xor UO_1466 (O_1466,N_29714,N_29307);
and UO_1467 (O_1467,N_29823,N_29157);
nand UO_1468 (O_1468,N_29716,N_29012);
or UO_1469 (O_1469,N_29675,N_29873);
xnor UO_1470 (O_1470,N_29270,N_29239);
and UO_1471 (O_1471,N_29922,N_29093);
nand UO_1472 (O_1472,N_29261,N_29707);
or UO_1473 (O_1473,N_29159,N_29189);
nand UO_1474 (O_1474,N_29366,N_29801);
xor UO_1475 (O_1475,N_29517,N_29816);
nor UO_1476 (O_1476,N_29331,N_29489);
or UO_1477 (O_1477,N_29179,N_29108);
nor UO_1478 (O_1478,N_29807,N_29251);
and UO_1479 (O_1479,N_29591,N_29146);
nor UO_1480 (O_1480,N_29881,N_29833);
xnor UO_1481 (O_1481,N_29419,N_29571);
nand UO_1482 (O_1482,N_29086,N_29472);
nand UO_1483 (O_1483,N_29267,N_29737);
nor UO_1484 (O_1484,N_29484,N_29951);
nor UO_1485 (O_1485,N_29715,N_29204);
nor UO_1486 (O_1486,N_29348,N_29578);
xor UO_1487 (O_1487,N_29353,N_29430);
xor UO_1488 (O_1488,N_29321,N_29036);
and UO_1489 (O_1489,N_29464,N_29355);
xor UO_1490 (O_1490,N_29360,N_29095);
nor UO_1491 (O_1491,N_29670,N_29551);
nor UO_1492 (O_1492,N_29119,N_29435);
nor UO_1493 (O_1493,N_29069,N_29199);
or UO_1494 (O_1494,N_29927,N_29361);
and UO_1495 (O_1495,N_29787,N_29190);
nand UO_1496 (O_1496,N_29306,N_29771);
or UO_1497 (O_1497,N_29962,N_29660);
and UO_1498 (O_1498,N_29794,N_29619);
and UO_1499 (O_1499,N_29068,N_29489);
nor UO_1500 (O_1500,N_29252,N_29046);
and UO_1501 (O_1501,N_29145,N_29268);
xor UO_1502 (O_1502,N_29890,N_29582);
and UO_1503 (O_1503,N_29788,N_29686);
xor UO_1504 (O_1504,N_29886,N_29983);
and UO_1505 (O_1505,N_29426,N_29696);
or UO_1506 (O_1506,N_29020,N_29860);
or UO_1507 (O_1507,N_29778,N_29947);
or UO_1508 (O_1508,N_29690,N_29840);
nand UO_1509 (O_1509,N_29858,N_29337);
and UO_1510 (O_1510,N_29571,N_29584);
nor UO_1511 (O_1511,N_29829,N_29671);
xnor UO_1512 (O_1512,N_29685,N_29440);
and UO_1513 (O_1513,N_29261,N_29099);
and UO_1514 (O_1514,N_29086,N_29695);
nand UO_1515 (O_1515,N_29976,N_29134);
nor UO_1516 (O_1516,N_29475,N_29759);
nand UO_1517 (O_1517,N_29098,N_29947);
xor UO_1518 (O_1518,N_29633,N_29171);
nand UO_1519 (O_1519,N_29100,N_29359);
nor UO_1520 (O_1520,N_29076,N_29802);
nor UO_1521 (O_1521,N_29866,N_29925);
or UO_1522 (O_1522,N_29603,N_29142);
and UO_1523 (O_1523,N_29519,N_29453);
nand UO_1524 (O_1524,N_29289,N_29022);
nor UO_1525 (O_1525,N_29197,N_29299);
and UO_1526 (O_1526,N_29418,N_29534);
or UO_1527 (O_1527,N_29743,N_29332);
nand UO_1528 (O_1528,N_29596,N_29355);
or UO_1529 (O_1529,N_29560,N_29970);
xnor UO_1530 (O_1530,N_29429,N_29718);
xor UO_1531 (O_1531,N_29801,N_29640);
nand UO_1532 (O_1532,N_29275,N_29775);
nor UO_1533 (O_1533,N_29428,N_29585);
nand UO_1534 (O_1534,N_29111,N_29870);
nor UO_1535 (O_1535,N_29925,N_29764);
or UO_1536 (O_1536,N_29796,N_29489);
or UO_1537 (O_1537,N_29736,N_29376);
nor UO_1538 (O_1538,N_29920,N_29667);
nor UO_1539 (O_1539,N_29234,N_29749);
and UO_1540 (O_1540,N_29313,N_29384);
or UO_1541 (O_1541,N_29840,N_29209);
xor UO_1542 (O_1542,N_29960,N_29146);
and UO_1543 (O_1543,N_29467,N_29678);
nand UO_1544 (O_1544,N_29482,N_29243);
or UO_1545 (O_1545,N_29370,N_29818);
and UO_1546 (O_1546,N_29988,N_29821);
nor UO_1547 (O_1547,N_29853,N_29582);
xor UO_1548 (O_1548,N_29432,N_29650);
or UO_1549 (O_1549,N_29521,N_29743);
xnor UO_1550 (O_1550,N_29832,N_29248);
xor UO_1551 (O_1551,N_29582,N_29021);
xor UO_1552 (O_1552,N_29564,N_29533);
xor UO_1553 (O_1553,N_29766,N_29082);
nand UO_1554 (O_1554,N_29892,N_29974);
and UO_1555 (O_1555,N_29114,N_29515);
xnor UO_1556 (O_1556,N_29487,N_29666);
xor UO_1557 (O_1557,N_29539,N_29936);
xnor UO_1558 (O_1558,N_29844,N_29944);
nand UO_1559 (O_1559,N_29300,N_29782);
or UO_1560 (O_1560,N_29887,N_29349);
xor UO_1561 (O_1561,N_29967,N_29484);
xor UO_1562 (O_1562,N_29837,N_29238);
or UO_1563 (O_1563,N_29156,N_29628);
or UO_1564 (O_1564,N_29810,N_29893);
nand UO_1565 (O_1565,N_29417,N_29494);
or UO_1566 (O_1566,N_29219,N_29500);
or UO_1567 (O_1567,N_29708,N_29892);
xnor UO_1568 (O_1568,N_29157,N_29492);
xnor UO_1569 (O_1569,N_29621,N_29749);
xnor UO_1570 (O_1570,N_29462,N_29353);
nor UO_1571 (O_1571,N_29056,N_29958);
nor UO_1572 (O_1572,N_29414,N_29948);
nand UO_1573 (O_1573,N_29797,N_29091);
xnor UO_1574 (O_1574,N_29704,N_29209);
and UO_1575 (O_1575,N_29808,N_29281);
nand UO_1576 (O_1576,N_29626,N_29581);
nor UO_1577 (O_1577,N_29017,N_29690);
nand UO_1578 (O_1578,N_29907,N_29674);
nor UO_1579 (O_1579,N_29584,N_29156);
nor UO_1580 (O_1580,N_29349,N_29578);
or UO_1581 (O_1581,N_29053,N_29535);
and UO_1582 (O_1582,N_29416,N_29371);
nand UO_1583 (O_1583,N_29413,N_29230);
or UO_1584 (O_1584,N_29420,N_29476);
nand UO_1585 (O_1585,N_29561,N_29523);
and UO_1586 (O_1586,N_29125,N_29240);
nor UO_1587 (O_1587,N_29694,N_29172);
nor UO_1588 (O_1588,N_29942,N_29649);
xor UO_1589 (O_1589,N_29534,N_29410);
nor UO_1590 (O_1590,N_29229,N_29888);
and UO_1591 (O_1591,N_29415,N_29686);
nand UO_1592 (O_1592,N_29356,N_29948);
xnor UO_1593 (O_1593,N_29798,N_29354);
nor UO_1594 (O_1594,N_29714,N_29906);
or UO_1595 (O_1595,N_29572,N_29645);
xor UO_1596 (O_1596,N_29887,N_29657);
and UO_1597 (O_1597,N_29920,N_29998);
xnor UO_1598 (O_1598,N_29779,N_29628);
or UO_1599 (O_1599,N_29020,N_29895);
and UO_1600 (O_1600,N_29556,N_29815);
and UO_1601 (O_1601,N_29344,N_29208);
xor UO_1602 (O_1602,N_29691,N_29082);
or UO_1603 (O_1603,N_29201,N_29400);
and UO_1604 (O_1604,N_29274,N_29132);
nor UO_1605 (O_1605,N_29245,N_29598);
or UO_1606 (O_1606,N_29196,N_29184);
or UO_1607 (O_1607,N_29862,N_29931);
or UO_1608 (O_1608,N_29928,N_29614);
nor UO_1609 (O_1609,N_29747,N_29367);
nand UO_1610 (O_1610,N_29671,N_29891);
xnor UO_1611 (O_1611,N_29210,N_29392);
nand UO_1612 (O_1612,N_29115,N_29786);
and UO_1613 (O_1613,N_29535,N_29010);
and UO_1614 (O_1614,N_29658,N_29363);
or UO_1615 (O_1615,N_29843,N_29507);
xor UO_1616 (O_1616,N_29423,N_29965);
nand UO_1617 (O_1617,N_29814,N_29054);
xnor UO_1618 (O_1618,N_29499,N_29611);
and UO_1619 (O_1619,N_29556,N_29877);
nor UO_1620 (O_1620,N_29310,N_29259);
xor UO_1621 (O_1621,N_29787,N_29199);
or UO_1622 (O_1622,N_29295,N_29438);
nand UO_1623 (O_1623,N_29836,N_29581);
xnor UO_1624 (O_1624,N_29576,N_29696);
nand UO_1625 (O_1625,N_29795,N_29558);
and UO_1626 (O_1626,N_29508,N_29091);
and UO_1627 (O_1627,N_29800,N_29642);
nand UO_1628 (O_1628,N_29729,N_29404);
or UO_1629 (O_1629,N_29037,N_29530);
nand UO_1630 (O_1630,N_29060,N_29268);
xor UO_1631 (O_1631,N_29337,N_29251);
xnor UO_1632 (O_1632,N_29506,N_29332);
nand UO_1633 (O_1633,N_29169,N_29231);
nor UO_1634 (O_1634,N_29924,N_29231);
nand UO_1635 (O_1635,N_29131,N_29642);
nand UO_1636 (O_1636,N_29575,N_29802);
or UO_1637 (O_1637,N_29734,N_29207);
or UO_1638 (O_1638,N_29327,N_29696);
or UO_1639 (O_1639,N_29856,N_29130);
and UO_1640 (O_1640,N_29522,N_29191);
or UO_1641 (O_1641,N_29322,N_29226);
xor UO_1642 (O_1642,N_29768,N_29335);
and UO_1643 (O_1643,N_29066,N_29130);
nor UO_1644 (O_1644,N_29831,N_29413);
and UO_1645 (O_1645,N_29712,N_29770);
or UO_1646 (O_1646,N_29798,N_29694);
and UO_1647 (O_1647,N_29515,N_29320);
nand UO_1648 (O_1648,N_29408,N_29389);
or UO_1649 (O_1649,N_29771,N_29385);
nand UO_1650 (O_1650,N_29511,N_29528);
xnor UO_1651 (O_1651,N_29740,N_29320);
nand UO_1652 (O_1652,N_29713,N_29809);
xor UO_1653 (O_1653,N_29525,N_29122);
xnor UO_1654 (O_1654,N_29420,N_29916);
or UO_1655 (O_1655,N_29112,N_29222);
xnor UO_1656 (O_1656,N_29193,N_29367);
nand UO_1657 (O_1657,N_29820,N_29181);
nand UO_1658 (O_1658,N_29395,N_29665);
or UO_1659 (O_1659,N_29943,N_29572);
xnor UO_1660 (O_1660,N_29701,N_29461);
and UO_1661 (O_1661,N_29376,N_29779);
nor UO_1662 (O_1662,N_29123,N_29323);
nor UO_1663 (O_1663,N_29266,N_29450);
or UO_1664 (O_1664,N_29195,N_29451);
or UO_1665 (O_1665,N_29904,N_29754);
or UO_1666 (O_1666,N_29975,N_29224);
or UO_1667 (O_1667,N_29156,N_29130);
nor UO_1668 (O_1668,N_29602,N_29730);
nor UO_1669 (O_1669,N_29724,N_29622);
or UO_1670 (O_1670,N_29260,N_29248);
and UO_1671 (O_1671,N_29192,N_29983);
nand UO_1672 (O_1672,N_29720,N_29084);
or UO_1673 (O_1673,N_29057,N_29647);
nor UO_1674 (O_1674,N_29239,N_29857);
nor UO_1675 (O_1675,N_29529,N_29752);
and UO_1676 (O_1676,N_29955,N_29187);
and UO_1677 (O_1677,N_29640,N_29539);
and UO_1678 (O_1678,N_29994,N_29935);
xor UO_1679 (O_1679,N_29456,N_29148);
or UO_1680 (O_1680,N_29428,N_29748);
and UO_1681 (O_1681,N_29714,N_29682);
or UO_1682 (O_1682,N_29928,N_29974);
or UO_1683 (O_1683,N_29201,N_29246);
xnor UO_1684 (O_1684,N_29482,N_29797);
or UO_1685 (O_1685,N_29899,N_29520);
or UO_1686 (O_1686,N_29032,N_29300);
nand UO_1687 (O_1687,N_29887,N_29318);
and UO_1688 (O_1688,N_29886,N_29901);
and UO_1689 (O_1689,N_29693,N_29308);
or UO_1690 (O_1690,N_29012,N_29037);
and UO_1691 (O_1691,N_29246,N_29131);
xor UO_1692 (O_1692,N_29805,N_29953);
nor UO_1693 (O_1693,N_29920,N_29193);
and UO_1694 (O_1694,N_29256,N_29510);
and UO_1695 (O_1695,N_29998,N_29404);
and UO_1696 (O_1696,N_29251,N_29550);
and UO_1697 (O_1697,N_29996,N_29249);
nand UO_1698 (O_1698,N_29529,N_29817);
nand UO_1699 (O_1699,N_29898,N_29384);
nor UO_1700 (O_1700,N_29258,N_29610);
nand UO_1701 (O_1701,N_29620,N_29844);
nand UO_1702 (O_1702,N_29829,N_29040);
or UO_1703 (O_1703,N_29417,N_29380);
nand UO_1704 (O_1704,N_29968,N_29405);
or UO_1705 (O_1705,N_29035,N_29117);
or UO_1706 (O_1706,N_29298,N_29511);
and UO_1707 (O_1707,N_29870,N_29967);
nor UO_1708 (O_1708,N_29079,N_29441);
nand UO_1709 (O_1709,N_29408,N_29431);
xor UO_1710 (O_1710,N_29338,N_29481);
or UO_1711 (O_1711,N_29861,N_29762);
and UO_1712 (O_1712,N_29185,N_29895);
nand UO_1713 (O_1713,N_29208,N_29742);
nor UO_1714 (O_1714,N_29707,N_29812);
or UO_1715 (O_1715,N_29289,N_29013);
nor UO_1716 (O_1716,N_29897,N_29196);
nor UO_1717 (O_1717,N_29326,N_29261);
or UO_1718 (O_1718,N_29772,N_29863);
and UO_1719 (O_1719,N_29889,N_29178);
and UO_1720 (O_1720,N_29015,N_29480);
or UO_1721 (O_1721,N_29287,N_29851);
nor UO_1722 (O_1722,N_29572,N_29637);
nor UO_1723 (O_1723,N_29261,N_29630);
nor UO_1724 (O_1724,N_29062,N_29304);
xor UO_1725 (O_1725,N_29391,N_29451);
nor UO_1726 (O_1726,N_29915,N_29269);
and UO_1727 (O_1727,N_29478,N_29756);
nand UO_1728 (O_1728,N_29415,N_29672);
nand UO_1729 (O_1729,N_29097,N_29644);
or UO_1730 (O_1730,N_29445,N_29177);
xnor UO_1731 (O_1731,N_29745,N_29207);
and UO_1732 (O_1732,N_29351,N_29115);
nand UO_1733 (O_1733,N_29452,N_29613);
nor UO_1734 (O_1734,N_29788,N_29590);
nand UO_1735 (O_1735,N_29182,N_29626);
or UO_1736 (O_1736,N_29181,N_29130);
nor UO_1737 (O_1737,N_29296,N_29667);
nor UO_1738 (O_1738,N_29176,N_29877);
nand UO_1739 (O_1739,N_29845,N_29680);
nand UO_1740 (O_1740,N_29426,N_29607);
nand UO_1741 (O_1741,N_29945,N_29829);
nor UO_1742 (O_1742,N_29812,N_29670);
and UO_1743 (O_1743,N_29574,N_29662);
or UO_1744 (O_1744,N_29991,N_29276);
and UO_1745 (O_1745,N_29689,N_29466);
xor UO_1746 (O_1746,N_29233,N_29930);
or UO_1747 (O_1747,N_29036,N_29315);
and UO_1748 (O_1748,N_29511,N_29130);
or UO_1749 (O_1749,N_29282,N_29572);
and UO_1750 (O_1750,N_29123,N_29859);
nor UO_1751 (O_1751,N_29857,N_29120);
and UO_1752 (O_1752,N_29310,N_29706);
xor UO_1753 (O_1753,N_29884,N_29979);
nor UO_1754 (O_1754,N_29397,N_29347);
xor UO_1755 (O_1755,N_29223,N_29759);
or UO_1756 (O_1756,N_29646,N_29093);
and UO_1757 (O_1757,N_29466,N_29264);
and UO_1758 (O_1758,N_29718,N_29638);
xor UO_1759 (O_1759,N_29137,N_29869);
or UO_1760 (O_1760,N_29852,N_29439);
nand UO_1761 (O_1761,N_29671,N_29265);
xnor UO_1762 (O_1762,N_29043,N_29437);
xor UO_1763 (O_1763,N_29377,N_29510);
or UO_1764 (O_1764,N_29359,N_29016);
xor UO_1765 (O_1765,N_29636,N_29801);
and UO_1766 (O_1766,N_29786,N_29253);
and UO_1767 (O_1767,N_29279,N_29715);
and UO_1768 (O_1768,N_29839,N_29673);
or UO_1769 (O_1769,N_29026,N_29928);
nand UO_1770 (O_1770,N_29178,N_29396);
nor UO_1771 (O_1771,N_29184,N_29323);
or UO_1772 (O_1772,N_29378,N_29138);
nand UO_1773 (O_1773,N_29315,N_29027);
nor UO_1774 (O_1774,N_29637,N_29264);
xnor UO_1775 (O_1775,N_29384,N_29798);
xnor UO_1776 (O_1776,N_29576,N_29639);
nor UO_1777 (O_1777,N_29334,N_29928);
and UO_1778 (O_1778,N_29990,N_29212);
or UO_1779 (O_1779,N_29590,N_29028);
xnor UO_1780 (O_1780,N_29013,N_29700);
and UO_1781 (O_1781,N_29459,N_29222);
or UO_1782 (O_1782,N_29945,N_29605);
and UO_1783 (O_1783,N_29864,N_29680);
xor UO_1784 (O_1784,N_29428,N_29465);
and UO_1785 (O_1785,N_29336,N_29826);
nor UO_1786 (O_1786,N_29452,N_29901);
xor UO_1787 (O_1787,N_29269,N_29271);
and UO_1788 (O_1788,N_29227,N_29767);
nand UO_1789 (O_1789,N_29708,N_29648);
xor UO_1790 (O_1790,N_29270,N_29521);
or UO_1791 (O_1791,N_29166,N_29151);
nand UO_1792 (O_1792,N_29620,N_29128);
nor UO_1793 (O_1793,N_29044,N_29559);
nor UO_1794 (O_1794,N_29498,N_29041);
nand UO_1795 (O_1795,N_29591,N_29792);
nand UO_1796 (O_1796,N_29467,N_29376);
nand UO_1797 (O_1797,N_29731,N_29813);
nor UO_1798 (O_1798,N_29264,N_29770);
or UO_1799 (O_1799,N_29909,N_29959);
xor UO_1800 (O_1800,N_29561,N_29496);
nor UO_1801 (O_1801,N_29675,N_29788);
or UO_1802 (O_1802,N_29398,N_29821);
nor UO_1803 (O_1803,N_29306,N_29345);
nor UO_1804 (O_1804,N_29312,N_29243);
xnor UO_1805 (O_1805,N_29214,N_29680);
xnor UO_1806 (O_1806,N_29748,N_29980);
or UO_1807 (O_1807,N_29236,N_29109);
or UO_1808 (O_1808,N_29979,N_29108);
and UO_1809 (O_1809,N_29734,N_29962);
nor UO_1810 (O_1810,N_29278,N_29938);
or UO_1811 (O_1811,N_29183,N_29564);
and UO_1812 (O_1812,N_29710,N_29404);
xor UO_1813 (O_1813,N_29644,N_29673);
or UO_1814 (O_1814,N_29682,N_29748);
or UO_1815 (O_1815,N_29280,N_29168);
xnor UO_1816 (O_1816,N_29148,N_29634);
and UO_1817 (O_1817,N_29644,N_29757);
xor UO_1818 (O_1818,N_29019,N_29194);
and UO_1819 (O_1819,N_29257,N_29292);
nor UO_1820 (O_1820,N_29248,N_29636);
or UO_1821 (O_1821,N_29454,N_29180);
nand UO_1822 (O_1822,N_29864,N_29467);
or UO_1823 (O_1823,N_29483,N_29354);
or UO_1824 (O_1824,N_29474,N_29134);
or UO_1825 (O_1825,N_29502,N_29821);
nand UO_1826 (O_1826,N_29026,N_29991);
nor UO_1827 (O_1827,N_29570,N_29089);
xnor UO_1828 (O_1828,N_29036,N_29825);
xor UO_1829 (O_1829,N_29854,N_29865);
xnor UO_1830 (O_1830,N_29475,N_29393);
xor UO_1831 (O_1831,N_29151,N_29023);
nand UO_1832 (O_1832,N_29511,N_29727);
and UO_1833 (O_1833,N_29953,N_29637);
xnor UO_1834 (O_1834,N_29687,N_29047);
and UO_1835 (O_1835,N_29036,N_29786);
and UO_1836 (O_1836,N_29269,N_29650);
and UO_1837 (O_1837,N_29226,N_29220);
nor UO_1838 (O_1838,N_29858,N_29297);
or UO_1839 (O_1839,N_29114,N_29989);
and UO_1840 (O_1840,N_29356,N_29541);
nor UO_1841 (O_1841,N_29406,N_29072);
or UO_1842 (O_1842,N_29972,N_29702);
xor UO_1843 (O_1843,N_29053,N_29225);
nor UO_1844 (O_1844,N_29655,N_29025);
or UO_1845 (O_1845,N_29109,N_29592);
or UO_1846 (O_1846,N_29670,N_29556);
nor UO_1847 (O_1847,N_29806,N_29430);
or UO_1848 (O_1848,N_29745,N_29417);
or UO_1849 (O_1849,N_29509,N_29489);
nor UO_1850 (O_1850,N_29143,N_29734);
and UO_1851 (O_1851,N_29167,N_29952);
nor UO_1852 (O_1852,N_29753,N_29940);
xor UO_1853 (O_1853,N_29576,N_29194);
nand UO_1854 (O_1854,N_29773,N_29324);
nand UO_1855 (O_1855,N_29386,N_29205);
nor UO_1856 (O_1856,N_29180,N_29112);
or UO_1857 (O_1857,N_29227,N_29384);
and UO_1858 (O_1858,N_29079,N_29590);
nand UO_1859 (O_1859,N_29249,N_29412);
and UO_1860 (O_1860,N_29936,N_29295);
and UO_1861 (O_1861,N_29727,N_29018);
nand UO_1862 (O_1862,N_29535,N_29712);
and UO_1863 (O_1863,N_29324,N_29997);
and UO_1864 (O_1864,N_29709,N_29106);
nand UO_1865 (O_1865,N_29763,N_29268);
nor UO_1866 (O_1866,N_29693,N_29595);
xor UO_1867 (O_1867,N_29012,N_29211);
and UO_1868 (O_1868,N_29183,N_29450);
xnor UO_1869 (O_1869,N_29010,N_29470);
or UO_1870 (O_1870,N_29821,N_29692);
xor UO_1871 (O_1871,N_29582,N_29164);
xor UO_1872 (O_1872,N_29507,N_29754);
and UO_1873 (O_1873,N_29108,N_29456);
nor UO_1874 (O_1874,N_29964,N_29446);
nand UO_1875 (O_1875,N_29843,N_29363);
nor UO_1876 (O_1876,N_29088,N_29050);
or UO_1877 (O_1877,N_29276,N_29865);
nor UO_1878 (O_1878,N_29548,N_29746);
and UO_1879 (O_1879,N_29396,N_29065);
xnor UO_1880 (O_1880,N_29428,N_29636);
nor UO_1881 (O_1881,N_29523,N_29554);
xor UO_1882 (O_1882,N_29054,N_29190);
and UO_1883 (O_1883,N_29022,N_29705);
or UO_1884 (O_1884,N_29335,N_29821);
nand UO_1885 (O_1885,N_29800,N_29847);
nand UO_1886 (O_1886,N_29169,N_29640);
nor UO_1887 (O_1887,N_29306,N_29073);
xor UO_1888 (O_1888,N_29102,N_29219);
or UO_1889 (O_1889,N_29265,N_29755);
xnor UO_1890 (O_1890,N_29036,N_29840);
or UO_1891 (O_1891,N_29833,N_29702);
and UO_1892 (O_1892,N_29354,N_29789);
and UO_1893 (O_1893,N_29343,N_29190);
nand UO_1894 (O_1894,N_29649,N_29203);
nand UO_1895 (O_1895,N_29776,N_29637);
nor UO_1896 (O_1896,N_29681,N_29631);
xnor UO_1897 (O_1897,N_29367,N_29388);
nor UO_1898 (O_1898,N_29518,N_29593);
and UO_1899 (O_1899,N_29534,N_29576);
nor UO_1900 (O_1900,N_29388,N_29523);
nor UO_1901 (O_1901,N_29859,N_29769);
xnor UO_1902 (O_1902,N_29579,N_29264);
or UO_1903 (O_1903,N_29742,N_29611);
xnor UO_1904 (O_1904,N_29710,N_29220);
nand UO_1905 (O_1905,N_29200,N_29698);
or UO_1906 (O_1906,N_29819,N_29011);
nor UO_1907 (O_1907,N_29543,N_29247);
xnor UO_1908 (O_1908,N_29517,N_29923);
or UO_1909 (O_1909,N_29663,N_29737);
nor UO_1910 (O_1910,N_29352,N_29354);
or UO_1911 (O_1911,N_29585,N_29896);
and UO_1912 (O_1912,N_29685,N_29075);
xor UO_1913 (O_1913,N_29682,N_29552);
xor UO_1914 (O_1914,N_29708,N_29093);
nand UO_1915 (O_1915,N_29283,N_29103);
nand UO_1916 (O_1916,N_29033,N_29102);
or UO_1917 (O_1917,N_29897,N_29659);
or UO_1918 (O_1918,N_29854,N_29583);
xor UO_1919 (O_1919,N_29576,N_29267);
nand UO_1920 (O_1920,N_29484,N_29616);
xnor UO_1921 (O_1921,N_29840,N_29830);
xor UO_1922 (O_1922,N_29377,N_29348);
nand UO_1923 (O_1923,N_29655,N_29839);
xor UO_1924 (O_1924,N_29899,N_29040);
and UO_1925 (O_1925,N_29486,N_29950);
or UO_1926 (O_1926,N_29819,N_29322);
nand UO_1927 (O_1927,N_29145,N_29569);
nand UO_1928 (O_1928,N_29696,N_29228);
or UO_1929 (O_1929,N_29082,N_29056);
and UO_1930 (O_1930,N_29709,N_29918);
nand UO_1931 (O_1931,N_29494,N_29492);
nor UO_1932 (O_1932,N_29500,N_29251);
and UO_1933 (O_1933,N_29665,N_29506);
xnor UO_1934 (O_1934,N_29551,N_29474);
xnor UO_1935 (O_1935,N_29771,N_29361);
xnor UO_1936 (O_1936,N_29846,N_29392);
and UO_1937 (O_1937,N_29073,N_29757);
or UO_1938 (O_1938,N_29395,N_29528);
nand UO_1939 (O_1939,N_29781,N_29252);
xor UO_1940 (O_1940,N_29992,N_29588);
and UO_1941 (O_1941,N_29286,N_29889);
nor UO_1942 (O_1942,N_29024,N_29428);
nor UO_1943 (O_1943,N_29591,N_29685);
nor UO_1944 (O_1944,N_29526,N_29252);
xor UO_1945 (O_1945,N_29071,N_29921);
and UO_1946 (O_1946,N_29147,N_29381);
or UO_1947 (O_1947,N_29741,N_29402);
nand UO_1948 (O_1948,N_29868,N_29367);
nor UO_1949 (O_1949,N_29831,N_29164);
and UO_1950 (O_1950,N_29985,N_29923);
nand UO_1951 (O_1951,N_29148,N_29466);
nand UO_1952 (O_1952,N_29760,N_29171);
and UO_1953 (O_1953,N_29318,N_29261);
or UO_1954 (O_1954,N_29659,N_29310);
and UO_1955 (O_1955,N_29602,N_29114);
xnor UO_1956 (O_1956,N_29909,N_29786);
nor UO_1957 (O_1957,N_29583,N_29462);
nand UO_1958 (O_1958,N_29424,N_29226);
xor UO_1959 (O_1959,N_29609,N_29820);
and UO_1960 (O_1960,N_29772,N_29907);
and UO_1961 (O_1961,N_29390,N_29880);
or UO_1962 (O_1962,N_29262,N_29050);
nand UO_1963 (O_1963,N_29915,N_29796);
and UO_1964 (O_1964,N_29384,N_29177);
and UO_1965 (O_1965,N_29061,N_29648);
nor UO_1966 (O_1966,N_29178,N_29502);
and UO_1967 (O_1967,N_29567,N_29131);
or UO_1968 (O_1968,N_29807,N_29899);
or UO_1969 (O_1969,N_29941,N_29579);
nand UO_1970 (O_1970,N_29496,N_29086);
or UO_1971 (O_1971,N_29467,N_29146);
nand UO_1972 (O_1972,N_29348,N_29938);
nor UO_1973 (O_1973,N_29125,N_29607);
nor UO_1974 (O_1974,N_29960,N_29749);
and UO_1975 (O_1975,N_29411,N_29792);
nand UO_1976 (O_1976,N_29668,N_29194);
nor UO_1977 (O_1977,N_29516,N_29945);
and UO_1978 (O_1978,N_29870,N_29343);
nand UO_1979 (O_1979,N_29957,N_29472);
nor UO_1980 (O_1980,N_29436,N_29235);
xnor UO_1981 (O_1981,N_29257,N_29672);
nand UO_1982 (O_1982,N_29161,N_29992);
nor UO_1983 (O_1983,N_29262,N_29871);
or UO_1984 (O_1984,N_29788,N_29717);
nand UO_1985 (O_1985,N_29973,N_29839);
or UO_1986 (O_1986,N_29210,N_29441);
and UO_1987 (O_1987,N_29897,N_29972);
nor UO_1988 (O_1988,N_29740,N_29162);
nor UO_1989 (O_1989,N_29599,N_29368);
nor UO_1990 (O_1990,N_29292,N_29808);
or UO_1991 (O_1991,N_29800,N_29218);
and UO_1992 (O_1992,N_29530,N_29268);
nor UO_1993 (O_1993,N_29636,N_29281);
or UO_1994 (O_1994,N_29576,N_29498);
nand UO_1995 (O_1995,N_29022,N_29419);
xnor UO_1996 (O_1996,N_29059,N_29519);
nor UO_1997 (O_1997,N_29318,N_29722);
xor UO_1998 (O_1998,N_29958,N_29826);
or UO_1999 (O_1999,N_29621,N_29778);
xnor UO_2000 (O_2000,N_29419,N_29295);
nor UO_2001 (O_2001,N_29606,N_29101);
nand UO_2002 (O_2002,N_29191,N_29926);
nor UO_2003 (O_2003,N_29582,N_29811);
nand UO_2004 (O_2004,N_29495,N_29192);
nor UO_2005 (O_2005,N_29066,N_29042);
nand UO_2006 (O_2006,N_29788,N_29591);
xor UO_2007 (O_2007,N_29815,N_29548);
xor UO_2008 (O_2008,N_29962,N_29985);
xor UO_2009 (O_2009,N_29686,N_29863);
nor UO_2010 (O_2010,N_29642,N_29999);
nor UO_2011 (O_2011,N_29718,N_29428);
or UO_2012 (O_2012,N_29600,N_29723);
or UO_2013 (O_2013,N_29981,N_29734);
nand UO_2014 (O_2014,N_29950,N_29738);
and UO_2015 (O_2015,N_29656,N_29868);
and UO_2016 (O_2016,N_29391,N_29190);
xor UO_2017 (O_2017,N_29779,N_29409);
xnor UO_2018 (O_2018,N_29307,N_29064);
and UO_2019 (O_2019,N_29810,N_29199);
nand UO_2020 (O_2020,N_29052,N_29004);
nand UO_2021 (O_2021,N_29996,N_29905);
or UO_2022 (O_2022,N_29433,N_29231);
nand UO_2023 (O_2023,N_29101,N_29905);
or UO_2024 (O_2024,N_29078,N_29268);
and UO_2025 (O_2025,N_29254,N_29822);
nor UO_2026 (O_2026,N_29234,N_29192);
xnor UO_2027 (O_2027,N_29946,N_29234);
or UO_2028 (O_2028,N_29799,N_29118);
and UO_2029 (O_2029,N_29972,N_29245);
nand UO_2030 (O_2030,N_29355,N_29089);
and UO_2031 (O_2031,N_29225,N_29433);
xnor UO_2032 (O_2032,N_29259,N_29101);
nor UO_2033 (O_2033,N_29516,N_29884);
or UO_2034 (O_2034,N_29875,N_29746);
and UO_2035 (O_2035,N_29669,N_29358);
xnor UO_2036 (O_2036,N_29538,N_29402);
nand UO_2037 (O_2037,N_29034,N_29602);
or UO_2038 (O_2038,N_29868,N_29607);
and UO_2039 (O_2039,N_29156,N_29896);
or UO_2040 (O_2040,N_29409,N_29955);
xor UO_2041 (O_2041,N_29063,N_29874);
or UO_2042 (O_2042,N_29412,N_29828);
xnor UO_2043 (O_2043,N_29450,N_29247);
and UO_2044 (O_2044,N_29026,N_29694);
and UO_2045 (O_2045,N_29936,N_29293);
nor UO_2046 (O_2046,N_29209,N_29278);
nand UO_2047 (O_2047,N_29189,N_29640);
nor UO_2048 (O_2048,N_29377,N_29899);
nor UO_2049 (O_2049,N_29777,N_29478);
or UO_2050 (O_2050,N_29425,N_29644);
or UO_2051 (O_2051,N_29897,N_29118);
or UO_2052 (O_2052,N_29555,N_29042);
or UO_2053 (O_2053,N_29596,N_29302);
nor UO_2054 (O_2054,N_29570,N_29386);
or UO_2055 (O_2055,N_29305,N_29100);
and UO_2056 (O_2056,N_29708,N_29317);
xnor UO_2057 (O_2057,N_29329,N_29761);
nand UO_2058 (O_2058,N_29841,N_29367);
xor UO_2059 (O_2059,N_29426,N_29829);
xnor UO_2060 (O_2060,N_29876,N_29302);
nand UO_2061 (O_2061,N_29762,N_29597);
or UO_2062 (O_2062,N_29370,N_29486);
or UO_2063 (O_2063,N_29925,N_29652);
or UO_2064 (O_2064,N_29051,N_29031);
xor UO_2065 (O_2065,N_29722,N_29656);
nor UO_2066 (O_2066,N_29011,N_29237);
xnor UO_2067 (O_2067,N_29259,N_29016);
nor UO_2068 (O_2068,N_29041,N_29833);
nand UO_2069 (O_2069,N_29758,N_29060);
nand UO_2070 (O_2070,N_29502,N_29501);
nor UO_2071 (O_2071,N_29124,N_29631);
nand UO_2072 (O_2072,N_29738,N_29146);
nor UO_2073 (O_2073,N_29380,N_29011);
xnor UO_2074 (O_2074,N_29217,N_29565);
or UO_2075 (O_2075,N_29598,N_29175);
nor UO_2076 (O_2076,N_29437,N_29945);
nand UO_2077 (O_2077,N_29605,N_29540);
xnor UO_2078 (O_2078,N_29005,N_29465);
nor UO_2079 (O_2079,N_29520,N_29959);
nor UO_2080 (O_2080,N_29879,N_29862);
or UO_2081 (O_2081,N_29874,N_29236);
xor UO_2082 (O_2082,N_29437,N_29334);
nor UO_2083 (O_2083,N_29592,N_29631);
xnor UO_2084 (O_2084,N_29284,N_29894);
nand UO_2085 (O_2085,N_29889,N_29649);
xor UO_2086 (O_2086,N_29039,N_29356);
xnor UO_2087 (O_2087,N_29678,N_29438);
nand UO_2088 (O_2088,N_29273,N_29784);
nand UO_2089 (O_2089,N_29890,N_29485);
xnor UO_2090 (O_2090,N_29069,N_29498);
nand UO_2091 (O_2091,N_29069,N_29281);
nor UO_2092 (O_2092,N_29160,N_29193);
nand UO_2093 (O_2093,N_29054,N_29186);
nand UO_2094 (O_2094,N_29883,N_29774);
nor UO_2095 (O_2095,N_29342,N_29783);
xnor UO_2096 (O_2096,N_29569,N_29862);
and UO_2097 (O_2097,N_29335,N_29404);
or UO_2098 (O_2098,N_29106,N_29186);
and UO_2099 (O_2099,N_29796,N_29893);
xor UO_2100 (O_2100,N_29959,N_29460);
nor UO_2101 (O_2101,N_29107,N_29178);
xnor UO_2102 (O_2102,N_29408,N_29830);
xnor UO_2103 (O_2103,N_29199,N_29026);
or UO_2104 (O_2104,N_29606,N_29763);
nor UO_2105 (O_2105,N_29084,N_29167);
nor UO_2106 (O_2106,N_29444,N_29230);
nor UO_2107 (O_2107,N_29635,N_29607);
xnor UO_2108 (O_2108,N_29762,N_29554);
and UO_2109 (O_2109,N_29613,N_29598);
nand UO_2110 (O_2110,N_29548,N_29050);
or UO_2111 (O_2111,N_29914,N_29188);
and UO_2112 (O_2112,N_29262,N_29995);
or UO_2113 (O_2113,N_29929,N_29949);
xnor UO_2114 (O_2114,N_29179,N_29400);
xnor UO_2115 (O_2115,N_29110,N_29311);
nand UO_2116 (O_2116,N_29824,N_29537);
or UO_2117 (O_2117,N_29539,N_29123);
nand UO_2118 (O_2118,N_29611,N_29367);
xor UO_2119 (O_2119,N_29075,N_29510);
nor UO_2120 (O_2120,N_29456,N_29458);
or UO_2121 (O_2121,N_29849,N_29310);
or UO_2122 (O_2122,N_29389,N_29197);
nand UO_2123 (O_2123,N_29937,N_29800);
nor UO_2124 (O_2124,N_29421,N_29061);
nand UO_2125 (O_2125,N_29314,N_29764);
xnor UO_2126 (O_2126,N_29395,N_29451);
xnor UO_2127 (O_2127,N_29458,N_29067);
xnor UO_2128 (O_2128,N_29794,N_29340);
nor UO_2129 (O_2129,N_29732,N_29779);
and UO_2130 (O_2130,N_29640,N_29152);
or UO_2131 (O_2131,N_29649,N_29742);
xnor UO_2132 (O_2132,N_29008,N_29532);
nand UO_2133 (O_2133,N_29645,N_29747);
nor UO_2134 (O_2134,N_29176,N_29848);
nand UO_2135 (O_2135,N_29636,N_29800);
and UO_2136 (O_2136,N_29536,N_29426);
and UO_2137 (O_2137,N_29580,N_29053);
or UO_2138 (O_2138,N_29432,N_29166);
and UO_2139 (O_2139,N_29314,N_29196);
xor UO_2140 (O_2140,N_29673,N_29608);
nand UO_2141 (O_2141,N_29134,N_29981);
and UO_2142 (O_2142,N_29399,N_29297);
or UO_2143 (O_2143,N_29240,N_29626);
nand UO_2144 (O_2144,N_29107,N_29157);
and UO_2145 (O_2145,N_29776,N_29292);
and UO_2146 (O_2146,N_29032,N_29767);
or UO_2147 (O_2147,N_29252,N_29989);
xor UO_2148 (O_2148,N_29101,N_29549);
or UO_2149 (O_2149,N_29458,N_29798);
nor UO_2150 (O_2150,N_29118,N_29574);
and UO_2151 (O_2151,N_29418,N_29122);
and UO_2152 (O_2152,N_29559,N_29869);
or UO_2153 (O_2153,N_29428,N_29786);
nor UO_2154 (O_2154,N_29869,N_29684);
or UO_2155 (O_2155,N_29263,N_29661);
or UO_2156 (O_2156,N_29778,N_29156);
xor UO_2157 (O_2157,N_29268,N_29397);
nor UO_2158 (O_2158,N_29468,N_29706);
and UO_2159 (O_2159,N_29518,N_29002);
nand UO_2160 (O_2160,N_29892,N_29258);
nand UO_2161 (O_2161,N_29062,N_29664);
xor UO_2162 (O_2162,N_29420,N_29173);
nand UO_2163 (O_2163,N_29698,N_29469);
or UO_2164 (O_2164,N_29492,N_29421);
and UO_2165 (O_2165,N_29550,N_29716);
nand UO_2166 (O_2166,N_29438,N_29951);
or UO_2167 (O_2167,N_29297,N_29265);
and UO_2168 (O_2168,N_29410,N_29849);
nand UO_2169 (O_2169,N_29443,N_29744);
xnor UO_2170 (O_2170,N_29265,N_29236);
and UO_2171 (O_2171,N_29263,N_29877);
xor UO_2172 (O_2172,N_29812,N_29228);
and UO_2173 (O_2173,N_29504,N_29552);
or UO_2174 (O_2174,N_29231,N_29154);
and UO_2175 (O_2175,N_29763,N_29843);
xnor UO_2176 (O_2176,N_29398,N_29008);
nor UO_2177 (O_2177,N_29221,N_29783);
and UO_2178 (O_2178,N_29232,N_29783);
and UO_2179 (O_2179,N_29933,N_29558);
xor UO_2180 (O_2180,N_29026,N_29966);
or UO_2181 (O_2181,N_29051,N_29577);
nor UO_2182 (O_2182,N_29883,N_29646);
and UO_2183 (O_2183,N_29518,N_29835);
nand UO_2184 (O_2184,N_29946,N_29698);
xnor UO_2185 (O_2185,N_29016,N_29012);
nand UO_2186 (O_2186,N_29135,N_29456);
and UO_2187 (O_2187,N_29511,N_29750);
nor UO_2188 (O_2188,N_29312,N_29441);
xnor UO_2189 (O_2189,N_29576,N_29243);
nor UO_2190 (O_2190,N_29164,N_29120);
nand UO_2191 (O_2191,N_29398,N_29084);
or UO_2192 (O_2192,N_29391,N_29487);
nand UO_2193 (O_2193,N_29326,N_29614);
xor UO_2194 (O_2194,N_29710,N_29532);
nand UO_2195 (O_2195,N_29703,N_29668);
xor UO_2196 (O_2196,N_29426,N_29666);
or UO_2197 (O_2197,N_29068,N_29472);
and UO_2198 (O_2198,N_29570,N_29535);
nor UO_2199 (O_2199,N_29974,N_29906);
nand UO_2200 (O_2200,N_29632,N_29060);
or UO_2201 (O_2201,N_29629,N_29777);
xor UO_2202 (O_2202,N_29540,N_29747);
or UO_2203 (O_2203,N_29818,N_29696);
or UO_2204 (O_2204,N_29121,N_29997);
nor UO_2205 (O_2205,N_29247,N_29990);
nor UO_2206 (O_2206,N_29730,N_29317);
xnor UO_2207 (O_2207,N_29108,N_29957);
nor UO_2208 (O_2208,N_29460,N_29007);
nor UO_2209 (O_2209,N_29103,N_29852);
or UO_2210 (O_2210,N_29112,N_29121);
or UO_2211 (O_2211,N_29357,N_29363);
or UO_2212 (O_2212,N_29048,N_29808);
nor UO_2213 (O_2213,N_29637,N_29215);
and UO_2214 (O_2214,N_29623,N_29116);
nand UO_2215 (O_2215,N_29214,N_29207);
or UO_2216 (O_2216,N_29835,N_29062);
nand UO_2217 (O_2217,N_29683,N_29625);
nand UO_2218 (O_2218,N_29446,N_29748);
xnor UO_2219 (O_2219,N_29744,N_29025);
nor UO_2220 (O_2220,N_29010,N_29768);
nor UO_2221 (O_2221,N_29284,N_29972);
or UO_2222 (O_2222,N_29367,N_29632);
nor UO_2223 (O_2223,N_29802,N_29753);
or UO_2224 (O_2224,N_29928,N_29281);
and UO_2225 (O_2225,N_29790,N_29786);
xnor UO_2226 (O_2226,N_29323,N_29785);
or UO_2227 (O_2227,N_29232,N_29418);
nand UO_2228 (O_2228,N_29837,N_29380);
and UO_2229 (O_2229,N_29082,N_29246);
and UO_2230 (O_2230,N_29842,N_29846);
nand UO_2231 (O_2231,N_29708,N_29021);
nor UO_2232 (O_2232,N_29880,N_29268);
nand UO_2233 (O_2233,N_29180,N_29940);
and UO_2234 (O_2234,N_29980,N_29507);
or UO_2235 (O_2235,N_29317,N_29841);
or UO_2236 (O_2236,N_29605,N_29753);
nor UO_2237 (O_2237,N_29768,N_29842);
xor UO_2238 (O_2238,N_29620,N_29884);
xnor UO_2239 (O_2239,N_29697,N_29021);
nor UO_2240 (O_2240,N_29075,N_29594);
and UO_2241 (O_2241,N_29430,N_29246);
and UO_2242 (O_2242,N_29484,N_29801);
nor UO_2243 (O_2243,N_29046,N_29231);
and UO_2244 (O_2244,N_29247,N_29329);
and UO_2245 (O_2245,N_29720,N_29659);
and UO_2246 (O_2246,N_29111,N_29250);
nor UO_2247 (O_2247,N_29646,N_29285);
xor UO_2248 (O_2248,N_29145,N_29933);
xnor UO_2249 (O_2249,N_29496,N_29049);
nand UO_2250 (O_2250,N_29690,N_29009);
xor UO_2251 (O_2251,N_29277,N_29249);
nor UO_2252 (O_2252,N_29297,N_29691);
and UO_2253 (O_2253,N_29636,N_29595);
nand UO_2254 (O_2254,N_29630,N_29448);
nor UO_2255 (O_2255,N_29153,N_29214);
or UO_2256 (O_2256,N_29671,N_29298);
xnor UO_2257 (O_2257,N_29046,N_29207);
nand UO_2258 (O_2258,N_29020,N_29473);
xnor UO_2259 (O_2259,N_29213,N_29894);
xnor UO_2260 (O_2260,N_29421,N_29764);
xor UO_2261 (O_2261,N_29526,N_29749);
and UO_2262 (O_2262,N_29664,N_29978);
nand UO_2263 (O_2263,N_29466,N_29037);
nor UO_2264 (O_2264,N_29564,N_29423);
nor UO_2265 (O_2265,N_29758,N_29386);
or UO_2266 (O_2266,N_29014,N_29785);
nor UO_2267 (O_2267,N_29202,N_29253);
xor UO_2268 (O_2268,N_29577,N_29594);
or UO_2269 (O_2269,N_29371,N_29278);
or UO_2270 (O_2270,N_29070,N_29968);
nand UO_2271 (O_2271,N_29513,N_29957);
and UO_2272 (O_2272,N_29976,N_29988);
nand UO_2273 (O_2273,N_29628,N_29050);
nor UO_2274 (O_2274,N_29241,N_29200);
nand UO_2275 (O_2275,N_29477,N_29415);
nand UO_2276 (O_2276,N_29740,N_29171);
xnor UO_2277 (O_2277,N_29508,N_29981);
nand UO_2278 (O_2278,N_29038,N_29118);
nor UO_2279 (O_2279,N_29366,N_29148);
nand UO_2280 (O_2280,N_29393,N_29584);
xnor UO_2281 (O_2281,N_29814,N_29962);
and UO_2282 (O_2282,N_29179,N_29096);
and UO_2283 (O_2283,N_29877,N_29733);
xor UO_2284 (O_2284,N_29576,N_29107);
xnor UO_2285 (O_2285,N_29726,N_29355);
xnor UO_2286 (O_2286,N_29643,N_29094);
nand UO_2287 (O_2287,N_29579,N_29269);
or UO_2288 (O_2288,N_29613,N_29564);
nand UO_2289 (O_2289,N_29958,N_29504);
xor UO_2290 (O_2290,N_29221,N_29234);
nand UO_2291 (O_2291,N_29319,N_29321);
nand UO_2292 (O_2292,N_29152,N_29147);
nand UO_2293 (O_2293,N_29299,N_29024);
xor UO_2294 (O_2294,N_29721,N_29033);
xor UO_2295 (O_2295,N_29232,N_29689);
and UO_2296 (O_2296,N_29713,N_29619);
nand UO_2297 (O_2297,N_29717,N_29252);
and UO_2298 (O_2298,N_29278,N_29497);
nand UO_2299 (O_2299,N_29405,N_29298);
nand UO_2300 (O_2300,N_29408,N_29860);
and UO_2301 (O_2301,N_29390,N_29008);
nand UO_2302 (O_2302,N_29601,N_29609);
and UO_2303 (O_2303,N_29572,N_29781);
or UO_2304 (O_2304,N_29484,N_29904);
nor UO_2305 (O_2305,N_29832,N_29804);
and UO_2306 (O_2306,N_29781,N_29652);
nor UO_2307 (O_2307,N_29263,N_29828);
nand UO_2308 (O_2308,N_29701,N_29832);
and UO_2309 (O_2309,N_29873,N_29489);
xnor UO_2310 (O_2310,N_29391,N_29070);
and UO_2311 (O_2311,N_29059,N_29681);
or UO_2312 (O_2312,N_29501,N_29524);
nand UO_2313 (O_2313,N_29212,N_29923);
nor UO_2314 (O_2314,N_29040,N_29068);
xor UO_2315 (O_2315,N_29145,N_29063);
and UO_2316 (O_2316,N_29650,N_29291);
nand UO_2317 (O_2317,N_29037,N_29894);
and UO_2318 (O_2318,N_29537,N_29943);
or UO_2319 (O_2319,N_29374,N_29373);
xnor UO_2320 (O_2320,N_29647,N_29401);
xnor UO_2321 (O_2321,N_29569,N_29117);
or UO_2322 (O_2322,N_29114,N_29269);
and UO_2323 (O_2323,N_29440,N_29095);
xor UO_2324 (O_2324,N_29864,N_29961);
xor UO_2325 (O_2325,N_29583,N_29981);
and UO_2326 (O_2326,N_29650,N_29379);
nor UO_2327 (O_2327,N_29942,N_29797);
or UO_2328 (O_2328,N_29671,N_29777);
or UO_2329 (O_2329,N_29067,N_29120);
xnor UO_2330 (O_2330,N_29595,N_29253);
and UO_2331 (O_2331,N_29492,N_29769);
xor UO_2332 (O_2332,N_29622,N_29524);
nand UO_2333 (O_2333,N_29771,N_29673);
nand UO_2334 (O_2334,N_29581,N_29651);
nand UO_2335 (O_2335,N_29745,N_29448);
xnor UO_2336 (O_2336,N_29858,N_29760);
xnor UO_2337 (O_2337,N_29872,N_29214);
or UO_2338 (O_2338,N_29878,N_29161);
nand UO_2339 (O_2339,N_29255,N_29416);
nand UO_2340 (O_2340,N_29107,N_29332);
xor UO_2341 (O_2341,N_29386,N_29465);
and UO_2342 (O_2342,N_29197,N_29720);
and UO_2343 (O_2343,N_29182,N_29743);
and UO_2344 (O_2344,N_29038,N_29293);
and UO_2345 (O_2345,N_29727,N_29105);
xor UO_2346 (O_2346,N_29831,N_29018);
or UO_2347 (O_2347,N_29685,N_29111);
nand UO_2348 (O_2348,N_29267,N_29842);
nand UO_2349 (O_2349,N_29818,N_29794);
nand UO_2350 (O_2350,N_29186,N_29325);
xnor UO_2351 (O_2351,N_29140,N_29183);
nor UO_2352 (O_2352,N_29309,N_29571);
nand UO_2353 (O_2353,N_29186,N_29252);
nand UO_2354 (O_2354,N_29635,N_29347);
and UO_2355 (O_2355,N_29090,N_29563);
nor UO_2356 (O_2356,N_29373,N_29871);
nor UO_2357 (O_2357,N_29486,N_29217);
nor UO_2358 (O_2358,N_29995,N_29178);
xor UO_2359 (O_2359,N_29743,N_29970);
and UO_2360 (O_2360,N_29047,N_29702);
nand UO_2361 (O_2361,N_29286,N_29203);
xor UO_2362 (O_2362,N_29056,N_29281);
or UO_2363 (O_2363,N_29505,N_29622);
or UO_2364 (O_2364,N_29169,N_29974);
nor UO_2365 (O_2365,N_29517,N_29338);
nand UO_2366 (O_2366,N_29252,N_29550);
and UO_2367 (O_2367,N_29272,N_29090);
nor UO_2368 (O_2368,N_29782,N_29103);
nor UO_2369 (O_2369,N_29898,N_29246);
xnor UO_2370 (O_2370,N_29454,N_29084);
or UO_2371 (O_2371,N_29800,N_29900);
xor UO_2372 (O_2372,N_29347,N_29432);
or UO_2373 (O_2373,N_29776,N_29787);
xor UO_2374 (O_2374,N_29097,N_29769);
and UO_2375 (O_2375,N_29130,N_29446);
and UO_2376 (O_2376,N_29240,N_29163);
or UO_2377 (O_2377,N_29263,N_29397);
nand UO_2378 (O_2378,N_29832,N_29186);
nor UO_2379 (O_2379,N_29924,N_29779);
or UO_2380 (O_2380,N_29839,N_29054);
nor UO_2381 (O_2381,N_29262,N_29326);
nor UO_2382 (O_2382,N_29291,N_29868);
or UO_2383 (O_2383,N_29732,N_29400);
and UO_2384 (O_2384,N_29659,N_29841);
xnor UO_2385 (O_2385,N_29487,N_29360);
or UO_2386 (O_2386,N_29481,N_29154);
xnor UO_2387 (O_2387,N_29365,N_29917);
xor UO_2388 (O_2388,N_29483,N_29885);
nand UO_2389 (O_2389,N_29056,N_29845);
xnor UO_2390 (O_2390,N_29601,N_29951);
or UO_2391 (O_2391,N_29338,N_29048);
xnor UO_2392 (O_2392,N_29418,N_29329);
nand UO_2393 (O_2393,N_29724,N_29472);
nand UO_2394 (O_2394,N_29762,N_29154);
nor UO_2395 (O_2395,N_29746,N_29684);
nor UO_2396 (O_2396,N_29536,N_29642);
xnor UO_2397 (O_2397,N_29383,N_29698);
xnor UO_2398 (O_2398,N_29484,N_29539);
nor UO_2399 (O_2399,N_29646,N_29918);
nand UO_2400 (O_2400,N_29411,N_29464);
and UO_2401 (O_2401,N_29143,N_29461);
nor UO_2402 (O_2402,N_29296,N_29791);
or UO_2403 (O_2403,N_29408,N_29347);
or UO_2404 (O_2404,N_29303,N_29815);
and UO_2405 (O_2405,N_29017,N_29098);
nor UO_2406 (O_2406,N_29906,N_29169);
xor UO_2407 (O_2407,N_29711,N_29211);
and UO_2408 (O_2408,N_29956,N_29255);
nand UO_2409 (O_2409,N_29752,N_29662);
and UO_2410 (O_2410,N_29880,N_29258);
and UO_2411 (O_2411,N_29904,N_29844);
xnor UO_2412 (O_2412,N_29662,N_29944);
nand UO_2413 (O_2413,N_29715,N_29228);
nand UO_2414 (O_2414,N_29759,N_29819);
nand UO_2415 (O_2415,N_29277,N_29235);
or UO_2416 (O_2416,N_29224,N_29782);
and UO_2417 (O_2417,N_29791,N_29913);
and UO_2418 (O_2418,N_29248,N_29059);
nand UO_2419 (O_2419,N_29122,N_29930);
and UO_2420 (O_2420,N_29619,N_29506);
xnor UO_2421 (O_2421,N_29545,N_29490);
or UO_2422 (O_2422,N_29861,N_29386);
xor UO_2423 (O_2423,N_29604,N_29280);
xnor UO_2424 (O_2424,N_29160,N_29026);
nand UO_2425 (O_2425,N_29825,N_29329);
nor UO_2426 (O_2426,N_29642,N_29089);
and UO_2427 (O_2427,N_29379,N_29895);
nor UO_2428 (O_2428,N_29950,N_29633);
xor UO_2429 (O_2429,N_29687,N_29223);
xnor UO_2430 (O_2430,N_29687,N_29366);
nand UO_2431 (O_2431,N_29208,N_29018);
nand UO_2432 (O_2432,N_29945,N_29401);
nor UO_2433 (O_2433,N_29601,N_29731);
nor UO_2434 (O_2434,N_29782,N_29986);
nand UO_2435 (O_2435,N_29465,N_29814);
nand UO_2436 (O_2436,N_29265,N_29696);
and UO_2437 (O_2437,N_29121,N_29760);
and UO_2438 (O_2438,N_29960,N_29563);
nand UO_2439 (O_2439,N_29796,N_29409);
xor UO_2440 (O_2440,N_29373,N_29854);
or UO_2441 (O_2441,N_29577,N_29268);
and UO_2442 (O_2442,N_29915,N_29021);
xnor UO_2443 (O_2443,N_29254,N_29665);
or UO_2444 (O_2444,N_29015,N_29399);
or UO_2445 (O_2445,N_29247,N_29365);
and UO_2446 (O_2446,N_29481,N_29475);
nor UO_2447 (O_2447,N_29035,N_29454);
nor UO_2448 (O_2448,N_29034,N_29432);
nand UO_2449 (O_2449,N_29328,N_29999);
and UO_2450 (O_2450,N_29340,N_29781);
and UO_2451 (O_2451,N_29783,N_29927);
nor UO_2452 (O_2452,N_29651,N_29573);
xnor UO_2453 (O_2453,N_29042,N_29848);
or UO_2454 (O_2454,N_29564,N_29242);
and UO_2455 (O_2455,N_29984,N_29964);
xor UO_2456 (O_2456,N_29988,N_29955);
xor UO_2457 (O_2457,N_29587,N_29071);
nand UO_2458 (O_2458,N_29295,N_29721);
and UO_2459 (O_2459,N_29765,N_29585);
nand UO_2460 (O_2460,N_29058,N_29512);
or UO_2461 (O_2461,N_29342,N_29703);
and UO_2462 (O_2462,N_29376,N_29717);
or UO_2463 (O_2463,N_29743,N_29750);
or UO_2464 (O_2464,N_29273,N_29247);
or UO_2465 (O_2465,N_29351,N_29069);
or UO_2466 (O_2466,N_29313,N_29187);
and UO_2467 (O_2467,N_29280,N_29818);
or UO_2468 (O_2468,N_29347,N_29479);
or UO_2469 (O_2469,N_29433,N_29410);
and UO_2470 (O_2470,N_29728,N_29233);
nor UO_2471 (O_2471,N_29029,N_29598);
xnor UO_2472 (O_2472,N_29506,N_29871);
or UO_2473 (O_2473,N_29119,N_29467);
and UO_2474 (O_2474,N_29377,N_29680);
or UO_2475 (O_2475,N_29276,N_29202);
nand UO_2476 (O_2476,N_29080,N_29196);
or UO_2477 (O_2477,N_29943,N_29079);
or UO_2478 (O_2478,N_29885,N_29677);
or UO_2479 (O_2479,N_29267,N_29760);
or UO_2480 (O_2480,N_29633,N_29928);
nand UO_2481 (O_2481,N_29777,N_29743);
xnor UO_2482 (O_2482,N_29196,N_29005);
and UO_2483 (O_2483,N_29509,N_29613);
nand UO_2484 (O_2484,N_29090,N_29138);
xor UO_2485 (O_2485,N_29832,N_29924);
nor UO_2486 (O_2486,N_29804,N_29239);
nand UO_2487 (O_2487,N_29771,N_29702);
xnor UO_2488 (O_2488,N_29250,N_29560);
xor UO_2489 (O_2489,N_29490,N_29213);
or UO_2490 (O_2490,N_29791,N_29777);
and UO_2491 (O_2491,N_29704,N_29037);
and UO_2492 (O_2492,N_29140,N_29677);
and UO_2493 (O_2493,N_29413,N_29914);
xor UO_2494 (O_2494,N_29738,N_29845);
or UO_2495 (O_2495,N_29915,N_29405);
and UO_2496 (O_2496,N_29180,N_29377);
or UO_2497 (O_2497,N_29239,N_29703);
nor UO_2498 (O_2498,N_29536,N_29777);
nor UO_2499 (O_2499,N_29029,N_29020);
and UO_2500 (O_2500,N_29726,N_29777);
and UO_2501 (O_2501,N_29697,N_29313);
or UO_2502 (O_2502,N_29799,N_29217);
nor UO_2503 (O_2503,N_29333,N_29989);
nor UO_2504 (O_2504,N_29542,N_29233);
or UO_2505 (O_2505,N_29285,N_29593);
nand UO_2506 (O_2506,N_29160,N_29960);
nor UO_2507 (O_2507,N_29695,N_29222);
and UO_2508 (O_2508,N_29383,N_29226);
nor UO_2509 (O_2509,N_29051,N_29925);
and UO_2510 (O_2510,N_29225,N_29956);
and UO_2511 (O_2511,N_29631,N_29817);
nor UO_2512 (O_2512,N_29010,N_29327);
xnor UO_2513 (O_2513,N_29799,N_29002);
and UO_2514 (O_2514,N_29107,N_29162);
xnor UO_2515 (O_2515,N_29269,N_29112);
xnor UO_2516 (O_2516,N_29752,N_29673);
and UO_2517 (O_2517,N_29854,N_29213);
nor UO_2518 (O_2518,N_29152,N_29168);
nor UO_2519 (O_2519,N_29890,N_29072);
xor UO_2520 (O_2520,N_29439,N_29818);
xor UO_2521 (O_2521,N_29124,N_29126);
nor UO_2522 (O_2522,N_29214,N_29287);
and UO_2523 (O_2523,N_29139,N_29487);
xor UO_2524 (O_2524,N_29978,N_29129);
and UO_2525 (O_2525,N_29099,N_29906);
nand UO_2526 (O_2526,N_29941,N_29225);
nor UO_2527 (O_2527,N_29515,N_29816);
and UO_2528 (O_2528,N_29597,N_29947);
and UO_2529 (O_2529,N_29504,N_29387);
nor UO_2530 (O_2530,N_29087,N_29153);
or UO_2531 (O_2531,N_29493,N_29522);
and UO_2532 (O_2532,N_29421,N_29453);
nand UO_2533 (O_2533,N_29548,N_29414);
or UO_2534 (O_2534,N_29353,N_29254);
or UO_2535 (O_2535,N_29114,N_29584);
nor UO_2536 (O_2536,N_29571,N_29020);
and UO_2537 (O_2537,N_29185,N_29893);
and UO_2538 (O_2538,N_29520,N_29365);
xor UO_2539 (O_2539,N_29416,N_29647);
or UO_2540 (O_2540,N_29146,N_29089);
and UO_2541 (O_2541,N_29952,N_29508);
xnor UO_2542 (O_2542,N_29444,N_29178);
and UO_2543 (O_2543,N_29770,N_29814);
and UO_2544 (O_2544,N_29927,N_29760);
and UO_2545 (O_2545,N_29234,N_29831);
and UO_2546 (O_2546,N_29224,N_29018);
xnor UO_2547 (O_2547,N_29937,N_29050);
xor UO_2548 (O_2548,N_29688,N_29915);
nand UO_2549 (O_2549,N_29106,N_29498);
xor UO_2550 (O_2550,N_29902,N_29245);
nand UO_2551 (O_2551,N_29899,N_29942);
xnor UO_2552 (O_2552,N_29729,N_29741);
nand UO_2553 (O_2553,N_29824,N_29574);
nor UO_2554 (O_2554,N_29432,N_29089);
and UO_2555 (O_2555,N_29451,N_29680);
and UO_2556 (O_2556,N_29441,N_29806);
or UO_2557 (O_2557,N_29538,N_29026);
and UO_2558 (O_2558,N_29566,N_29735);
xor UO_2559 (O_2559,N_29316,N_29878);
xor UO_2560 (O_2560,N_29302,N_29740);
nand UO_2561 (O_2561,N_29134,N_29596);
nand UO_2562 (O_2562,N_29573,N_29122);
and UO_2563 (O_2563,N_29857,N_29069);
nand UO_2564 (O_2564,N_29688,N_29098);
nand UO_2565 (O_2565,N_29165,N_29239);
xor UO_2566 (O_2566,N_29895,N_29423);
or UO_2567 (O_2567,N_29714,N_29270);
xnor UO_2568 (O_2568,N_29041,N_29171);
xnor UO_2569 (O_2569,N_29467,N_29233);
nor UO_2570 (O_2570,N_29400,N_29344);
nand UO_2571 (O_2571,N_29516,N_29407);
or UO_2572 (O_2572,N_29013,N_29240);
xor UO_2573 (O_2573,N_29489,N_29321);
or UO_2574 (O_2574,N_29396,N_29972);
nand UO_2575 (O_2575,N_29743,N_29820);
nand UO_2576 (O_2576,N_29521,N_29166);
nand UO_2577 (O_2577,N_29785,N_29984);
and UO_2578 (O_2578,N_29011,N_29302);
or UO_2579 (O_2579,N_29850,N_29785);
xnor UO_2580 (O_2580,N_29850,N_29852);
nor UO_2581 (O_2581,N_29924,N_29117);
nor UO_2582 (O_2582,N_29994,N_29206);
and UO_2583 (O_2583,N_29064,N_29642);
nor UO_2584 (O_2584,N_29441,N_29655);
nor UO_2585 (O_2585,N_29513,N_29870);
and UO_2586 (O_2586,N_29994,N_29212);
and UO_2587 (O_2587,N_29380,N_29522);
xnor UO_2588 (O_2588,N_29038,N_29499);
or UO_2589 (O_2589,N_29017,N_29025);
xor UO_2590 (O_2590,N_29624,N_29781);
nor UO_2591 (O_2591,N_29962,N_29107);
nand UO_2592 (O_2592,N_29749,N_29425);
or UO_2593 (O_2593,N_29249,N_29282);
xnor UO_2594 (O_2594,N_29736,N_29966);
and UO_2595 (O_2595,N_29432,N_29452);
or UO_2596 (O_2596,N_29663,N_29287);
xor UO_2597 (O_2597,N_29916,N_29944);
nor UO_2598 (O_2598,N_29826,N_29228);
nand UO_2599 (O_2599,N_29569,N_29339);
nand UO_2600 (O_2600,N_29869,N_29108);
and UO_2601 (O_2601,N_29168,N_29533);
nor UO_2602 (O_2602,N_29380,N_29121);
and UO_2603 (O_2603,N_29670,N_29292);
nand UO_2604 (O_2604,N_29985,N_29783);
nand UO_2605 (O_2605,N_29195,N_29105);
and UO_2606 (O_2606,N_29743,N_29836);
or UO_2607 (O_2607,N_29369,N_29266);
xor UO_2608 (O_2608,N_29246,N_29027);
nand UO_2609 (O_2609,N_29127,N_29634);
xor UO_2610 (O_2610,N_29000,N_29540);
xor UO_2611 (O_2611,N_29761,N_29612);
nand UO_2612 (O_2612,N_29469,N_29176);
nand UO_2613 (O_2613,N_29112,N_29114);
or UO_2614 (O_2614,N_29856,N_29181);
or UO_2615 (O_2615,N_29228,N_29717);
and UO_2616 (O_2616,N_29743,N_29335);
or UO_2617 (O_2617,N_29053,N_29316);
nor UO_2618 (O_2618,N_29059,N_29969);
nand UO_2619 (O_2619,N_29871,N_29102);
and UO_2620 (O_2620,N_29827,N_29733);
and UO_2621 (O_2621,N_29804,N_29465);
nand UO_2622 (O_2622,N_29873,N_29070);
xnor UO_2623 (O_2623,N_29050,N_29199);
nand UO_2624 (O_2624,N_29451,N_29427);
nand UO_2625 (O_2625,N_29310,N_29743);
and UO_2626 (O_2626,N_29219,N_29534);
nand UO_2627 (O_2627,N_29709,N_29858);
and UO_2628 (O_2628,N_29968,N_29912);
and UO_2629 (O_2629,N_29229,N_29455);
nor UO_2630 (O_2630,N_29222,N_29114);
xor UO_2631 (O_2631,N_29690,N_29752);
nor UO_2632 (O_2632,N_29931,N_29228);
nor UO_2633 (O_2633,N_29763,N_29346);
nand UO_2634 (O_2634,N_29518,N_29795);
xor UO_2635 (O_2635,N_29760,N_29098);
xnor UO_2636 (O_2636,N_29739,N_29915);
xor UO_2637 (O_2637,N_29129,N_29701);
xor UO_2638 (O_2638,N_29010,N_29647);
xnor UO_2639 (O_2639,N_29454,N_29575);
nor UO_2640 (O_2640,N_29155,N_29882);
nand UO_2641 (O_2641,N_29592,N_29872);
or UO_2642 (O_2642,N_29339,N_29220);
nor UO_2643 (O_2643,N_29218,N_29865);
and UO_2644 (O_2644,N_29361,N_29900);
xor UO_2645 (O_2645,N_29164,N_29222);
xnor UO_2646 (O_2646,N_29691,N_29398);
xnor UO_2647 (O_2647,N_29117,N_29528);
xnor UO_2648 (O_2648,N_29609,N_29854);
xnor UO_2649 (O_2649,N_29247,N_29376);
and UO_2650 (O_2650,N_29112,N_29638);
nand UO_2651 (O_2651,N_29478,N_29127);
and UO_2652 (O_2652,N_29785,N_29274);
and UO_2653 (O_2653,N_29425,N_29682);
nand UO_2654 (O_2654,N_29140,N_29685);
nor UO_2655 (O_2655,N_29120,N_29545);
xnor UO_2656 (O_2656,N_29486,N_29759);
nand UO_2657 (O_2657,N_29533,N_29181);
xor UO_2658 (O_2658,N_29464,N_29768);
and UO_2659 (O_2659,N_29943,N_29308);
nand UO_2660 (O_2660,N_29233,N_29434);
and UO_2661 (O_2661,N_29156,N_29390);
xor UO_2662 (O_2662,N_29488,N_29986);
nor UO_2663 (O_2663,N_29473,N_29863);
or UO_2664 (O_2664,N_29201,N_29300);
nand UO_2665 (O_2665,N_29169,N_29294);
nor UO_2666 (O_2666,N_29935,N_29819);
nor UO_2667 (O_2667,N_29550,N_29486);
nand UO_2668 (O_2668,N_29200,N_29474);
or UO_2669 (O_2669,N_29614,N_29322);
xor UO_2670 (O_2670,N_29217,N_29584);
and UO_2671 (O_2671,N_29845,N_29698);
nor UO_2672 (O_2672,N_29855,N_29964);
and UO_2673 (O_2673,N_29474,N_29949);
nor UO_2674 (O_2674,N_29957,N_29919);
and UO_2675 (O_2675,N_29975,N_29216);
xnor UO_2676 (O_2676,N_29139,N_29257);
nor UO_2677 (O_2677,N_29307,N_29460);
and UO_2678 (O_2678,N_29675,N_29854);
and UO_2679 (O_2679,N_29818,N_29566);
xnor UO_2680 (O_2680,N_29868,N_29041);
nand UO_2681 (O_2681,N_29401,N_29890);
xor UO_2682 (O_2682,N_29112,N_29274);
nand UO_2683 (O_2683,N_29770,N_29877);
xnor UO_2684 (O_2684,N_29757,N_29947);
or UO_2685 (O_2685,N_29677,N_29850);
or UO_2686 (O_2686,N_29668,N_29604);
or UO_2687 (O_2687,N_29936,N_29985);
xor UO_2688 (O_2688,N_29983,N_29078);
nand UO_2689 (O_2689,N_29592,N_29460);
and UO_2690 (O_2690,N_29150,N_29221);
or UO_2691 (O_2691,N_29187,N_29032);
nor UO_2692 (O_2692,N_29899,N_29188);
xnor UO_2693 (O_2693,N_29358,N_29719);
and UO_2694 (O_2694,N_29987,N_29363);
or UO_2695 (O_2695,N_29530,N_29644);
or UO_2696 (O_2696,N_29646,N_29695);
nor UO_2697 (O_2697,N_29805,N_29588);
nor UO_2698 (O_2698,N_29284,N_29962);
xnor UO_2699 (O_2699,N_29154,N_29921);
nor UO_2700 (O_2700,N_29847,N_29819);
nor UO_2701 (O_2701,N_29542,N_29763);
and UO_2702 (O_2702,N_29923,N_29555);
and UO_2703 (O_2703,N_29576,N_29110);
nor UO_2704 (O_2704,N_29383,N_29316);
xor UO_2705 (O_2705,N_29147,N_29722);
nor UO_2706 (O_2706,N_29046,N_29285);
xor UO_2707 (O_2707,N_29879,N_29527);
nor UO_2708 (O_2708,N_29324,N_29502);
xnor UO_2709 (O_2709,N_29496,N_29979);
xor UO_2710 (O_2710,N_29029,N_29032);
and UO_2711 (O_2711,N_29291,N_29141);
xnor UO_2712 (O_2712,N_29455,N_29636);
nor UO_2713 (O_2713,N_29084,N_29792);
or UO_2714 (O_2714,N_29124,N_29037);
or UO_2715 (O_2715,N_29075,N_29718);
and UO_2716 (O_2716,N_29904,N_29214);
or UO_2717 (O_2717,N_29152,N_29015);
and UO_2718 (O_2718,N_29819,N_29967);
nor UO_2719 (O_2719,N_29817,N_29394);
and UO_2720 (O_2720,N_29800,N_29313);
or UO_2721 (O_2721,N_29016,N_29285);
nor UO_2722 (O_2722,N_29686,N_29772);
nand UO_2723 (O_2723,N_29801,N_29444);
nand UO_2724 (O_2724,N_29313,N_29687);
xnor UO_2725 (O_2725,N_29172,N_29840);
or UO_2726 (O_2726,N_29132,N_29099);
nand UO_2727 (O_2727,N_29563,N_29801);
or UO_2728 (O_2728,N_29706,N_29623);
xor UO_2729 (O_2729,N_29283,N_29293);
nor UO_2730 (O_2730,N_29276,N_29923);
or UO_2731 (O_2731,N_29146,N_29044);
and UO_2732 (O_2732,N_29628,N_29928);
nor UO_2733 (O_2733,N_29735,N_29048);
nand UO_2734 (O_2734,N_29910,N_29126);
xnor UO_2735 (O_2735,N_29100,N_29916);
or UO_2736 (O_2736,N_29397,N_29595);
nor UO_2737 (O_2737,N_29415,N_29201);
or UO_2738 (O_2738,N_29788,N_29287);
nand UO_2739 (O_2739,N_29603,N_29366);
and UO_2740 (O_2740,N_29871,N_29603);
xor UO_2741 (O_2741,N_29801,N_29234);
xor UO_2742 (O_2742,N_29025,N_29528);
nor UO_2743 (O_2743,N_29178,N_29985);
and UO_2744 (O_2744,N_29933,N_29662);
nor UO_2745 (O_2745,N_29491,N_29034);
nand UO_2746 (O_2746,N_29530,N_29475);
xnor UO_2747 (O_2747,N_29626,N_29294);
xor UO_2748 (O_2748,N_29001,N_29851);
xor UO_2749 (O_2749,N_29452,N_29644);
and UO_2750 (O_2750,N_29573,N_29523);
or UO_2751 (O_2751,N_29625,N_29657);
nor UO_2752 (O_2752,N_29910,N_29953);
nor UO_2753 (O_2753,N_29605,N_29053);
nor UO_2754 (O_2754,N_29554,N_29854);
nor UO_2755 (O_2755,N_29216,N_29526);
nor UO_2756 (O_2756,N_29768,N_29496);
nor UO_2757 (O_2757,N_29850,N_29755);
or UO_2758 (O_2758,N_29093,N_29213);
and UO_2759 (O_2759,N_29376,N_29796);
nor UO_2760 (O_2760,N_29211,N_29885);
nand UO_2761 (O_2761,N_29698,N_29665);
xnor UO_2762 (O_2762,N_29080,N_29210);
and UO_2763 (O_2763,N_29095,N_29533);
and UO_2764 (O_2764,N_29977,N_29282);
nand UO_2765 (O_2765,N_29753,N_29028);
or UO_2766 (O_2766,N_29828,N_29735);
and UO_2767 (O_2767,N_29066,N_29692);
or UO_2768 (O_2768,N_29544,N_29026);
nand UO_2769 (O_2769,N_29181,N_29707);
nand UO_2770 (O_2770,N_29536,N_29971);
xor UO_2771 (O_2771,N_29567,N_29383);
nor UO_2772 (O_2772,N_29355,N_29034);
or UO_2773 (O_2773,N_29095,N_29747);
nor UO_2774 (O_2774,N_29331,N_29059);
xor UO_2775 (O_2775,N_29447,N_29173);
or UO_2776 (O_2776,N_29317,N_29728);
nand UO_2777 (O_2777,N_29601,N_29581);
xnor UO_2778 (O_2778,N_29055,N_29584);
or UO_2779 (O_2779,N_29226,N_29536);
and UO_2780 (O_2780,N_29040,N_29597);
nand UO_2781 (O_2781,N_29517,N_29385);
or UO_2782 (O_2782,N_29181,N_29718);
or UO_2783 (O_2783,N_29311,N_29945);
xnor UO_2784 (O_2784,N_29210,N_29607);
or UO_2785 (O_2785,N_29440,N_29648);
nand UO_2786 (O_2786,N_29893,N_29177);
nand UO_2787 (O_2787,N_29457,N_29528);
xor UO_2788 (O_2788,N_29310,N_29409);
nand UO_2789 (O_2789,N_29935,N_29363);
nor UO_2790 (O_2790,N_29116,N_29471);
and UO_2791 (O_2791,N_29882,N_29426);
and UO_2792 (O_2792,N_29718,N_29601);
nand UO_2793 (O_2793,N_29164,N_29538);
nand UO_2794 (O_2794,N_29775,N_29261);
xor UO_2795 (O_2795,N_29574,N_29235);
xor UO_2796 (O_2796,N_29849,N_29174);
nand UO_2797 (O_2797,N_29219,N_29485);
xnor UO_2798 (O_2798,N_29687,N_29070);
and UO_2799 (O_2799,N_29829,N_29773);
and UO_2800 (O_2800,N_29362,N_29752);
nand UO_2801 (O_2801,N_29652,N_29687);
or UO_2802 (O_2802,N_29592,N_29531);
or UO_2803 (O_2803,N_29259,N_29723);
or UO_2804 (O_2804,N_29606,N_29859);
or UO_2805 (O_2805,N_29843,N_29030);
xor UO_2806 (O_2806,N_29074,N_29543);
nor UO_2807 (O_2807,N_29618,N_29723);
xor UO_2808 (O_2808,N_29946,N_29726);
xor UO_2809 (O_2809,N_29421,N_29906);
xor UO_2810 (O_2810,N_29609,N_29547);
or UO_2811 (O_2811,N_29232,N_29667);
xnor UO_2812 (O_2812,N_29169,N_29527);
nand UO_2813 (O_2813,N_29569,N_29548);
nand UO_2814 (O_2814,N_29320,N_29402);
or UO_2815 (O_2815,N_29227,N_29707);
or UO_2816 (O_2816,N_29500,N_29361);
and UO_2817 (O_2817,N_29166,N_29329);
nand UO_2818 (O_2818,N_29877,N_29998);
nor UO_2819 (O_2819,N_29995,N_29883);
or UO_2820 (O_2820,N_29057,N_29554);
and UO_2821 (O_2821,N_29267,N_29624);
and UO_2822 (O_2822,N_29595,N_29360);
xor UO_2823 (O_2823,N_29560,N_29906);
nor UO_2824 (O_2824,N_29263,N_29291);
nor UO_2825 (O_2825,N_29487,N_29066);
xor UO_2826 (O_2826,N_29207,N_29874);
and UO_2827 (O_2827,N_29999,N_29434);
nor UO_2828 (O_2828,N_29081,N_29774);
xor UO_2829 (O_2829,N_29856,N_29667);
nor UO_2830 (O_2830,N_29463,N_29070);
nor UO_2831 (O_2831,N_29306,N_29342);
or UO_2832 (O_2832,N_29238,N_29056);
nor UO_2833 (O_2833,N_29626,N_29335);
and UO_2834 (O_2834,N_29336,N_29623);
xnor UO_2835 (O_2835,N_29827,N_29927);
xor UO_2836 (O_2836,N_29995,N_29037);
and UO_2837 (O_2837,N_29165,N_29489);
nor UO_2838 (O_2838,N_29127,N_29601);
nor UO_2839 (O_2839,N_29614,N_29179);
xor UO_2840 (O_2840,N_29496,N_29173);
and UO_2841 (O_2841,N_29009,N_29041);
or UO_2842 (O_2842,N_29822,N_29509);
nand UO_2843 (O_2843,N_29788,N_29806);
xor UO_2844 (O_2844,N_29318,N_29122);
nand UO_2845 (O_2845,N_29763,N_29080);
xnor UO_2846 (O_2846,N_29297,N_29710);
xnor UO_2847 (O_2847,N_29373,N_29210);
nor UO_2848 (O_2848,N_29631,N_29148);
nor UO_2849 (O_2849,N_29872,N_29419);
nor UO_2850 (O_2850,N_29994,N_29900);
nor UO_2851 (O_2851,N_29250,N_29156);
nor UO_2852 (O_2852,N_29180,N_29619);
nand UO_2853 (O_2853,N_29310,N_29042);
nor UO_2854 (O_2854,N_29603,N_29825);
nand UO_2855 (O_2855,N_29609,N_29603);
and UO_2856 (O_2856,N_29544,N_29250);
nand UO_2857 (O_2857,N_29232,N_29525);
and UO_2858 (O_2858,N_29523,N_29866);
or UO_2859 (O_2859,N_29591,N_29120);
xnor UO_2860 (O_2860,N_29622,N_29536);
nor UO_2861 (O_2861,N_29065,N_29261);
xor UO_2862 (O_2862,N_29630,N_29605);
and UO_2863 (O_2863,N_29433,N_29554);
or UO_2864 (O_2864,N_29729,N_29051);
nor UO_2865 (O_2865,N_29264,N_29072);
xnor UO_2866 (O_2866,N_29314,N_29919);
nor UO_2867 (O_2867,N_29695,N_29813);
nand UO_2868 (O_2868,N_29252,N_29326);
nor UO_2869 (O_2869,N_29663,N_29869);
nand UO_2870 (O_2870,N_29860,N_29937);
or UO_2871 (O_2871,N_29488,N_29806);
and UO_2872 (O_2872,N_29153,N_29752);
or UO_2873 (O_2873,N_29547,N_29333);
or UO_2874 (O_2874,N_29141,N_29893);
and UO_2875 (O_2875,N_29168,N_29861);
nand UO_2876 (O_2876,N_29287,N_29444);
and UO_2877 (O_2877,N_29967,N_29920);
or UO_2878 (O_2878,N_29440,N_29611);
and UO_2879 (O_2879,N_29577,N_29215);
nor UO_2880 (O_2880,N_29438,N_29005);
nand UO_2881 (O_2881,N_29863,N_29076);
xor UO_2882 (O_2882,N_29374,N_29737);
or UO_2883 (O_2883,N_29101,N_29895);
xnor UO_2884 (O_2884,N_29661,N_29919);
and UO_2885 (O_2885,N_29156,N_29976);
xor UO_2886 (O_2886,N_29236,N_29093);
xor UO_2887 (O_2887,N_29572,N_29075);
or UO_2888 (O_2888,N_29221,N_29157);
or UO_2889 (O_2889,N_29341,N_29068);
or UO_2890 (O_2890,N_29519,N_29123);
and UO_2891 (O_2891,N_29634,N_29173);
or UO_2892 (O_2892,N_29463,N_29180);
xor UO_2893 (O_2893,N_29420,N_29739);
xnor UO_2894 (O_2894,N_29469,N_29579);
or UO_2895 (O_2895,N_29989,N_29582);
or UO_2896 (O_2896,N_29174,N_29514);
nor UO_2897 (O_2897,N_29553,N_29201);
and UO_2898 (O_2898,N_29000,N_29907);
nand UO_2899 (O_2899,N_29424,N_29406);
nor UO_2900 (O_2900,N_29645,N_29107);
or UO_2901 (O_2901,N_29165,N_29047);
or UO_2902 (O_2902,N_29601,N_29847);
nor UO_2903 (O_2903,N_29891,N_29896);
and UO_2904 (O_2904,N_29532,N_29131);
nor UO_2905 (O_2905,N_29606,N_29900);
or UO_2906 (O_2906,N_29910,N_29824);
nor UO_2907 (O_2907,N_29012,N_29446);
xnor UO_2908 (O_2908,N_29121,N_29795);
nor UO_2909 (O_2909,N_29733,N_29189);
nor UO_2910 (O_2910,N_29766,N_29912);
and UO_2911 (O_2911,N_29636,N_29909);
or UO_2912 (O_2912,N_29794,N_29788);
nor UO_2913 (O_2913,N_29645,N_29479);
nor UO_2914 (O_2914,N_29194,N_29282);
and UO_2915 (O_2915,N_29053,N_29954);
nand UO_2916 (O_2916,N_29074,N_29300);
xnor UO_2917 (O_2917,N_29467,N_29136);
or UO_2918 (O_2918,N_29402,N_29959);
nand UO_2919 (O_2919,N_29578,N_29999);
or UO_2920 (O_2920,N_29568,N_29961);
nor UO_2921 (O_2921,N_29203,N_29562);
and UO_2922 (O_2922,N_29303,N_29860);
nand UO_2923 (O_2923,N_29760,N_29081);
nor UO_2924 (O_2924,N_29841,N_29364);
nor UO_2925 (O_2925,N_29156,N_29060);
or UO_2926 (O_2926,N_29373,N_29527);
or UO_2927 (O_2927,N_29888,N_29564);
xnor UO_2928 (O_2928,N_29618,N_29516);
nor UO_2929 (O_2929,N_29736,N_29375);
or UO_2930 (O_2930,N_29875,N_29627);
or UO_2931 (O_2931,N_29255,N_29756);
xor UO_2932 (O_2932,N_29658,N_29808);
xnor UO_2933 (O_2933,N_29956,N_29708);
xor UO_2934 (O_2934,N_29514,N_29270);
nor UO_2935 (O_2935,N_29788,N_29381);
nor UO_2936 (O_2936,N_29124,N_29103);
nand UO_2937 (O_2937,N_29485,N_29590);
xor UO_2938 (O_2938,N_29880,N_29821);
nor UO_2939 (O_2939,N_29026,N_29475);
xor UO_2940 (O_2940,N_29244,N_29502);
and UO_2941 (O_2941,N_29577,N_29936);
nand UO_2942 (O_2942,N_29567,N_29732);
and UO_2943 (O_2943,N_29002,N_29561);
nor UO_2944 (O_2944,N_29644,N_29705);
nand UO_2945 (O_2945,N_29596,N_29925);
and UO_2946 (O_2946,N_29131,N_29742);
or UO_2947 (O_2947,N_29795,N_29295);
and UO_2948 (O_2948,N_29070,N_29239);
and UO_2949 (O_2949,N_29045,N_29245);
nor UO_2950 (O_2950,N_29482,N_29557);
nand UO_2951 (O_2951,N_29639,N_29606);
and UO_2952 (O_2952,N_29277,N_29480);
or UO_2953 (O_2953,N_29435,N_29078);
nor UO_2954 (O_2954,N_29733,N_29130);
and UO_2955 (O_2955,N_29735,N_29948);
or UO_2956 (O_2956,N_29351,N_29645);
or UO_2957 (O_2957,N_29156,N_29216);
xor UO_2958 (O_2958,N_29929,N_29707);
xnor UO_2959 (O_2959,N_29510,N_29747);
nand UO_2960 (O_2960,N_29526,N_29791);
nor UO_2961 (O_2961,N_29849,N_29657);
nand UO_2962 (O_2962,N_29830,N_29333);
nor UO_2963 (O_2963,N_29092,N_29660);
or UO_2964 (O_2964,N_29429,N_29496);
and UO_2965 (O_2965,N_29691,N_29200);
and UO_2966 (O_2966,N_29771,N_29156);
nor UO_2967 (O_2967,N_29551,N_29314);
xor UO_2968 (O_2968,N_29084,N_29733);
and UO_2969 (O_2969,N_29910,N_29931);
xnor UO_2970 (O_2970,N_29753,N_29852);
or UO_2971 (O_2971,N_29387,N_29195);
and UO_2972 (O_2972,N_29066,N_29155);
nand UO_2973 (O_2973,N_29176,N_29633);
nor UO_2974 (O_2974,N_29746,N_29123);
nor UO_2975 (O_2975,N_29306,N_29335);
xnor UO_2976 (O_2976,N_29996,N_29537);
nand UO_2977 (O_2977,N_29478,N_29114);
and UO_2978 (O_2978,N_29414,N_29174);
nand UO_2979 (O_2979,N_29635,N_29408);
nand UO_2980 (O_2980,N_29360,N_29587);
and UO_2981 (O_2981,N_29140,N_29956);
and UO_2982 (O_2982,N_29498,N_29771);
xnor UO_2983 (O_2983,N_29680,N_29885);
nor UO_2984 (O_2984,N_29597,N_29344);
nor UO_2985 (O_2985,N_29129,N_29094);
or UO_2986 (O_2986,N_29316,N_29476);
xor UO_2987 (O_2987,N_29377,N_29315);
nand UO_2988 (O_2988,N_29173,N_29226);
nand UO_2989 (O_2989,N_29767,N_29505);
and UO_2990 (O_2990,N_29014,N_29416);
or UO_2991 (O_2991,N_29739,N_29814);
and UO_2992 (O_2992,N_29067,N_29579);
xor UO_2993 (O_2993,N_29241,N_29262);
or UO_2994 (O_2994,N_29947,N_29558);
or UO_2995 (O_2995,N_29849,N_29049);
nand UO_2996 (O_2996,N_29385,N_29302);
or UO_2997 (O_2997,N_29906,N_29480);
nor UO_2998 (O_2998,N_29101,N_29335);
xnor UO_2999 (O_2999,N_29912,N_29404);
and UO_3000 (O_3000,N_29118,N_29980);
nand UO_3001 (O_3001,N_29413,N_29908);
nand UO_3002 (O_3002,N_29896,N_29034);
nor UO_3003 (O_3003,N_29950,N_29232);
xor UO_3004 (O_3004,N_29918,N_29038);
or UO_3005 (O_3005,N_29759,N_29021);
nor UO_3006 (O_3006,N_29904,N_29026);
xor UO_3007 (O_3007,N_29794,N_29757);
xor UO_3008 (O_3008,N_29502,N_29522);
and UO_3009 (O_3009,N_29337,N_29958);
nand UO_3010 (O_3010,N_29972,N_29757);
nand UO_3011 (O_3011,N_29784,N_29587);
and UO_3012 (O_3012,N_29508,N_29712);
and UO_3013 (O_3013,N_29476,N_29408);
nand UO_3014 (O_3014,N_29895,N_29968);
xor UO_3015 (O_3015,N_29055,N_29250);
xnor UO_3016 (O_3016,N_29998,N_29978);
and UO_3017 (O_3017,N_29518,N_29463);
and UO_3018 (O_3018,N_29985,N_29068);
nor UO_3019 (O_3019,N_29654,N_29702);
and UO_3020 (O_3020,N_29463,N_29992);
nor UO_3021 (O_3021,N_29141,N_29404);
nand UO_3022 (O_3022,N_29723,N_29934);
xnor UO_3023 (O_3023,N_29220,N_29279);
or UO_3024 (O_3024,N_29669,N_29767);
and UO_3025 (O_3025,N_29341,N_29222);
nor UO_3026 (O_3026,N_29284,N_29582);
or UO_3027 (O_3027,N_29303,N_29773);
and UO_3028 (O_3028,N_29237,N_29576);
xnor UO_3029 (O_3029,N_29104,N_29598);
and UO_3030 (O_3030,N_29797,N_29287);
nor UO_3031 (O_3031,N_29751,N_29256);
and UO_3032 (O_3032,N_29802,N_29003);
nor UO_3033 (O_3033,N_29199,N_29371);
and UO_3034 (O_3034,N_29277,N_29787);
nor UO_3035 (O_3035,N_29943,N_29306);
nand UO_3036 (O_3036,N_29420,N_29042);
nor UO_3037 (O_3037,N_29357,N_29501);
nand UO_3038 (O_3038,N_29569,N_29403);
or UO_3039 (O_3039,N_29959,N_29312);
or UO_3040 (O_3040,N_29104,N_29459);
nand UO_3041 (O_3041,N_29212,N_29320);
xor UO_3042 (O_3042,N_29032,N_29778);
or UO_3043 (O_3043,N_29029,N_29492);
xnor UO_3044 (O_3044,N_29956,N_29482);
or UO_3045 (O_3045,N_29494,N_29872);
nor UO_3046 (O_3046,N_29796,N_29646);
nand UO_3047 (O_3047,N_29129,N_29051);
nor UO_3048 (O_3048,N_29709,N_29000);
and UO_3049 (O_3049,N_29800,N_29611);
nor UO_3050 (O_3050,N_29415,N_29385);
or UO_3051 (O_3051,N_29834,N_29892);
and UO_3052 (O_3052,N_29144,N_29540);
and UO_3053 (O_3053,N_29662,N_29660);
xnor UO_3054 (O_3054,N_29757,N_29850);
xnor UO_3055 (O_3055,N_29044,N_29996);
nand UO_3056 (O_3056,N_29949,N_29779);
or UO_3057 (O_3057,N_29586,N_29878);
or UO_3058 (O_3058,N_29178,N_29518);
and UO_3059 (O_3059,N_29084,N_29542);
and UO_3060 (O_3060,N_29201,N_29242);
nor UO_3061 (O_3061,N_29998,N_29774);
nand UO_3062 (O_3062,N_29028,N_29283);
xnor UO_3063 (O_3063,N_29445,N_29237);
nand UO_3064 (O_3064,N_29645,N_29113);
xor UO_3065 (O_3065,N_29368,N_29969);
or UO_3066 (O_3066,N_29101,N_29334);
nand UO_3067 (O_3067,N_29165,N_29811);
nor UO_3068 (O_3068,N_29826,N_29717);
xnor UO_3069 (O_3069,N_29550,N_29580);
nor UO_3070 (O_3070,N_29388,N_29326);
nor UO_3071 (O_3071,N_29791,N_29275);
or UO_3072 (O_3072,N_29596,N_29185);
or UO_3073 (O_3073,N_29214,N_29885);
xor UO_3074 (O_3074,N_29281,N_29116);
and UO_3075 (O_3075,N_29596,N_29824);
nand UO_3076 (O_3076,N_29615,N_29583);
nand UO_3077 (O_3077,N_29720,N_29921);
xnor UO_3078 (O_3078,N_29772,N_29688);
nor UO_3079 (O_3079,N_29711,N_29370);
nor UO_3080 (O_3080,N_29408,N_29562);
or UO_3081 (O_3081,N_29674,N_29815);
nor UO_3082 (O_3082,N_29292,N_29786);
and UO_3083 (O_3083,N_29985,N_29565);
nand UO_3084 (O_3084,N_29480,N_29201);
xor UO_3085 (O_3085,N_29621,N_29864);
nor UO_3086 (O_3086,N_29377,N_29768);
nand UO_3087 (O_3087,N_29855,N_29062);
or UO_3088 (O_3088,N_29380,N_29411);
nor UO_3089 (O_3089,N_29748,N_29586);
and UO_3090 (O_3090,N_29566,N_29583);
xor UO_3091 (O_3091,N_29352,N_29373);
and UO_3092 (O_3092,N_29865,N_29381);
nor UO_3093 (O_3093,N_29444,N_29785);
nor UO_3094 (O_3094,N_29268,N_29810);
and UO_3095 (O_3095,N_29196,N_29495);
nand UO_3096 (O_3096,N_29344,N_29195);
xnor UO_3097 (O_3097,N_29429,N_29582);
xor UO_3098 (O_3098,N_29810,N_29497);
nor UO_3099 (O_3099,N_29973,N_29862);
xnor UO_3100 (O_3100,N_29687,N_29179);
or UO_3101 (O_3101,N_29373,N_29552);
and UO_3102 (O_3102,N_29056,N_29917);
nand UO_3103 (O_3103,N_29598,N_29297);
nor UO_3104 (O_3104,N_29071,N_29268);
xor UO_3105 (O_3105,N_29103,N_29996);
nand UO_3106 (O_3106,N_29403,N_29473);
nor UO_3107 (O_3107,N_29247,N_29797);
xnor UO_3108 (O_3108,N_29077,N_29682);
nor UO_3109 (O_3109,N_29625,N_29122);
nand UO_3110 (O_3110,N_29983,N_29699);
or UO_3111 (O_3111,N_29490,N_29889);
nor UO_3112 (O_3112,N_29461,N_29560);
and UO_3113 (O_3113,N_29956,N_29083);
xnor UO_3114 (O_3114,N_29450,N_29271);
nor UO_3115 (O_3115,N_29981,N_29606);
nor UO_3116 (O_3116,N_29643,N_29033);
and UO_3117 (O_3117,N_29506,N_29559);
and UO_3118 (O_3118,N_29963,N_29886);
or UO_3119 (O_3119,N_29123,N_29271);
or UO_3120 (O_3120,N_29775,N_29450);
nand UO_3121 (O_3121,N_29345,N_29346);
nor UO_3122 (O_3122,N_29621,N_29559);
nand UO_3123 (O_3123,N_29607,N_29118);
or UO_3124 (O_3124,N_29097,N_29192);
or UO_3125 (O_3125,N_29692,N_29997);
and UO_3126 (O_3126,N_29833,N_29003);
or UO_3127 (O_3127,N_29006,N_29065);
nor UO_3128 (O_3128,N_29739,N_29112);
nand UO_3129 (O_3129,N_29963,N_29377);
and UO_3130 (O_3130,N_29985,N_29485);
and UO_3131 (O_3131,N_29521,N_29273);
nand UO_3132 (O_3132,N_29581,N_29889);
and UO_3133 (O_3133,N_29492,N_29644);
and UO_3134 (O_3134,N_29349,N_29788);
or UO_3135 (O_3135,N_29969,N_29437);
and UO_3136 (O_3136,N_29351,N_29901);
or UO_3137 (O_3137,N_29726,N_29821);
xnor UO_3138 (O_3138,N_29194,N_29355);
and UO_3139 (O_3139,N_29054,N_29098);
or UO_3140 (O_3140,N_29378,N_29786);
and UO_3141 (O_3141,N_29003,N_29474);
or UO_3142 (O_3142,N_29601,N_29273);
nand UO_3143 (O_3143,N_29791,N_29696);
and UO_3144 (O_3144,N_29214,N_29481);
nand UO_3145 (O_3145,N_29025,N_29768);
or UO_3146 (O_3146,N_29967,N_29245);
xor UO_3147 (O_3147,N_29784,N_29573);
or UO_3148 (O_3148,N_29218,N_29157);
and UO_3149 (O_3149,N_29835,N_29279);
nor UO_3150 (O_3150,N_29223,N_29919);
nand UO_3151 (O_3151,N_29658,N_29463);
and UO_3152 (O_3152,N_29409,N_29129);
xor UO_3153 (O_3153,N_29926,N_29514);
nor UO_3154 (O_3154,N_29492,N_29071);
nand UO_3155 (O_3155,N_29286,N_29862);
xnor UO_3156 (O_3156,N_29902,N_29701);
or UO_3157 (O_3157,N_29524,N_29118);
nor UO_3158 (O_3158,N_29619,N_29935);
xnor UO_3159 (O_3159,N_29634,N_29224);
nand UO_3160 (O_3160,N_29063,N_29318);
and UO_3161 (O_3161,N_29803,N_29876);
xnor UO_3162 (O_3162,N_29405,N_29229);
xnor UO_3163 (O_3163,N_29153,N_29150);
nor UO_3164 (O_3164,N_29073,N_29870);
xnor UO_3165 (O_3165,N_29130,N_29707);
or UO_3166 (O_3166,N_29197,N_29380);
or UO_3167 (O_3167,N_29911,N_29917);
or UO_3168 (O_3168,N_29278,N_29470);
or UO_3169 (O_3169,N_29550,N_29041);
or UO_3170 (O_3170,N_29964,N_29110);
xnor UO_3171 (O_3171,N_29640,N_29288);
nand UO_3172 (O_3172,N_29917,N_29198);
or UO_3173 (O_3173,N_29218,N_29567);
nand UO_3174 (O_3174,N_29345,N_29936);
and UO_3175 (O_3175,N_29869,N_29363);
and UO_3176 (O_3176,N_29869,N_29463);
xnor UO_3177 (O_3177,N_29602,N_29481);
xor UO_3178 (O_3178,N_29580,N_29907);
xnor UO_3179 (O_3179,N_29151,N_29888);
or UO_3180 (O_3180,N_29893,N_29146);
nand UO_3181 (O_3181,N_29194,N_29306);
nor UO_3182 (O_3182,N_29757,N_29187);
or UO_3183 (O_3183,N_29482,N_29384);
xnor UO_3184 (O_3184,N_29310,N_29836);
xor UO_3185 (O_3185,N_29070,N_29471);
nand UO_3186 (O_3186,N_29451,N_29679);
and UO_3187 (O_3187,N_29613,N_29479);
nand UO_3188 (O_3188,N_29042,N_29175);
and UO_3189 (O_3189,N_29811,N_29297);
xnor UO_3190 (O_3190,N_29958,N_29215);
nand UO_3191 (O_3191,N_29998,N_29821);
and UO_3192 (O_3192,N_29185,N_29844);
nor UO_3193 (O_3193,N_29387,N_29663);
nor UO_3194 (O_3194,N_29120,N_29292);
xnor UO_3195 (O_3195,N_29276,N_29954);
nor UO_3196 (O_3196,N_29199,N_29667);
and UO_3197 (O_3197,N_29759,N_29936);
or UO_3198 (O_3198,N_29267,N_29452);
nor UO_3199 (O_3199,N_29991,N_29545);
nand UO_3200 (O_3200,N_29384,N_29984);
nand UO_3201 (O_3201,N_29075,N_29873);
and UO_3202 (O_3202,N_29029,N_29447);
nand UO_3203 (O_3203,N_29658,N_29849);
nor UO_3204 (O_3204,N_29749,N_29432);
nand UO_3205 (O_3205,N_29068,N_29374);
nand UO_3206 (O_3206,N_29471,N_29606);
nor UO_3207 (O_3207,N_29498,N_29416);
xnor UO_3208 (O_3208,N_29885,N_29002);
xor UO_3209 (O_3209,N_29345,N_29435);
nor UO_3210 (O_3210,N_29527,N_29331);
or UO_3211 (O_3211,N_29639,N_29134);
nand UO_3212 (O_3212,N_29755,N_29315);
xor UO_3213 (O_3213,N_29205,N_29279);
nand UO_3214 (O_3214,N_29081,N_29160);
and UO_3215 (O_3215,N_29328,N_29654);
nand UO_3216 (O_3216,N_29197,N_29462);
and UO_3217 (O_3217,N_29533,N_29354);
nor UO_3218 (O_3218,N_29576,N_29503);
nor UO_3219 (O_3219,N_29206,N_29584);
or UO_3220 (O_3220,N_29712,N_29877);
xnor UO_3221 (O_3221,N_29531,N_29857);
xor UO_3222 (O_3222,N_29608,N_29277);
or UO_3223 (O_3223,N_29938,N_29095);
nor UO_3224 (O_3224,N_29953,N_29066);
nor UO_3225 (O_3225,N_29310,N_29115);
and UO_3226 (O_3226,N_29997,N_29821);
and UO_3227 (O_3227,N_29638,N_29351);
xnor UO_3228 (O_3228,N_29748,N_29909);
and UO_3229 (O_3229,N_29613,N_29783);
nand UO_3230 (O_3230,N_29732,N_29638);
or UO_3231 (O_3231,N_29798,N_29829);
and UO_3232 (O_3232,N_29650,N_29669);
xnor UO_3233 (O_3233,N_29965,N_29226);
xnor UO_3234 (O_3234,N_29082,N_29985);
xnor UO_3235 (O_3235,N_29345,N_29434);
and UO_3236 (O_3236,N_29565,N_29935);
or UO_3237 (O_3237,N_29374,N_29079);
nor UO_3238 (O_3238,N_29331,N_29921);
xnor UO_3239 (O_3239,N_29024,N_29746);
nor UO_3240 (O_3240,N_29222,N_29898);
nand UO_3241 (O_3241,N_29881,N_29734);
or UO_3242 (O_3242,N_29959,N_29233);
and UO_3243 (O_3243,N_29961,N_29679);
xnor UO_3244 (O_3244,N_29703,N_29677);
nor UO_3245 (O_3245,N_29855,N_29602);
nand UO_3246 (O_3246,N_29316,N_29911);
and UO_3247 (O_3247,N_29291,N_29853);
or UO_3248 (O_3248,N_29074,N_29934);
nand UO_3249 (O_3249,N_29315,N_29838);
nand UO_3250 (O_3250,N_29399,N_29087);
nor UO_3251 (O_3251,N_29678,N_29484);
xnor UO_3252 (O_3252,N_29334,N_29511);
nor UO_3253 (O_3253,N_29553,N_29760);
xor UO_3254 (O_3254,N_29073,N_29783);
or UO_3255 (O_3255,N_29257,N_29782);
or UO_3256 (O_3256,N_29863,N_29337);
nor UO_3257 (O_3257,N_29509,N_29959);
xnor UO_3258 (O_3258,N_29037,N_29865);
nor UO_3259 (O_3259,N_29190,N_29252);
nand UO_3260 (O_3260,N_29058,N_29207);
or UO_3261 (O_3261,N_29246,N_29209);
nand UO_3262 (O_3262,N_29134,N_29943);
or UO_3263 (O_3263,N_29304,N_29242);
or UO_3264 (O_3264,N_29473,N_29924);
xnor UO_3265 (O_3265,N_29180,N_29140);
and UO_3266 (O_3266,N_29020,N_29296);
and UO_3267 (O_3267,N_29334,N_29915);
or UO_3268 (O_3268,N_29281,N_29119);
nand UO_3269 (O_3269,N_29450,N_29065);
and UO_3270 (O_3270,N_29785,N_29494);
nor UO_3271 (O_3271,N_29663,N_29348);
xnor UO_3272 (O_3272,N_29185,N_29290);
nand UO_3273 (O_3273,N_29507,N_29274);
or UO_3274 (O_3274,N_29280,N_29578);
and UO_3275 (O_3275,N_29331,N_29309);
nand UO_3276 (O_3276,N_29040,N_29543);
or UO_3277 (O_3277,N_29620,N_29041);
and UO_3278 (O_3278,N_29139,N_29081);
and UO_3279 (O_3279,N_29044,N_29861);
and UO_3280 (O_3280,N_29086,N_29332);
nor UO_3281 (O_3281,N_29468,N_29711);
nand UO_3282 (O_3282,N_29758,N_29189);
or UO_3283 (O_3283,N_29991,N_29113);
and UO_3284 (O_3284,N_29998,N_29198);
and UO_3285 (O_3285,N_29859,N_29982);
or UO_3286 (O_3286,N_29285,N_29392);
or UO_3287 (O_3287,N_29088,N_29926);
xnor UO_3288 (O_3288,N_29509,N_29807);
nor UO_3289 (O_3289,N_29310,N_29578);
or UO_3290 (O_3290,N_29376,N_29748);
nor UO_3291 (O_3291,N_29942,N_29757);
and UO_3292 (O_3292,N_29901,N_29631);
nand UO_3293 (O_3293,N_29313,N_29097);
and UO_3294 (O_3294,N_29571,N_29767);
or UO_3295 (O_3295,N_29203,N_29434);
nand UO_3296 (O_3296,N_29417,N_29746);
and UO_3297 (O_3297,N_29962,N_29230);
nand UO_3298 (O_3298,N_29184,N_29951);
or UO_3299 (O_3299,N_29452,N_29473);
or UO_3300 (O_3300,N_29299,N_29582);
nand UO_3301 (O_3301,N_29469,N_29495);
or UO_3302 (O_3302,N_29924,N_29198);
nand UO_3303 (O_3303,N_29242,N_29516);
nor UO_3304 (O_3304,N_29400,N_29289);
xor UO_3305 (O_3305,N_29794,N_29990);
nand UO_3306 (O_3306,N_29911,N_29175);
nor UO_3307 (O_3307,N_29582,N_29641);
or UO_3308 (O_3308,N_29242,N_29848);
nor UO_3309 (O_3309,N_29249,N_29488);
nor UO_3310 (O_3310,N_29146,N_29015);
or UO_3311 (O_3311,N_29884,N_29890);
nor UO_3312 (O_3312,N_29550,N_29965);
nor UO_3313 (O_3313,N_29529,N_29376);
nand UO_3314 (O_3314,N_29387,N_29266);
nor UO_3315 (O_3315,N_29035,N_29473);
nand UO_3316 (O_3316,N_29624,N_29774);
or UO_3317 (O_3317,N_29125,N_29521);
and UO_3318 (O_3318,N_29518,N_29023);
nand UO_3319 (O_3319,N_29299,N_29952);
xnor UO_3320 (O_3320,N_29272,N_29174);
nor UO_3321 (O_3321,N_29488,N_29571);
or UO_3322 (O_3322,N_29458,N_29684);
or UO_3323 (O_3323,N_29077,N_29982);
or UO_3324 (O_3324,N_29967,N_29490);
nand UO_3325 (O_3325,N_29041,N_29573);
or UO_3326 (O_3326,N_29944,N_29189);
nor UO_3327 (O_3327,N_29126,N_29385);
nor UO_3328 (O_3328,N_29133,N_29725);
nand UO_3329 (O_3329,N_29794,N_29013);
or UO_3330 (O_3330,N_29334,N_29796);
xor UO_3331 (O_3331,N_29548,N_29488);
nor UO_3332 (O_3332,N_29071,N_29486);
and UO_3333 (O_3333,N_29232,N_29578);
nand UO_3334 (O_3334,N_29434,N_29248);
xor UO_3335 (O_3335,N_29502,N_29878);
or UO_3336 (O_3336,N_29757,N_29891);
nor UO_3337 (O_3337,N_29648,N_29495);
or UO_3338 (O_3338,N_29838,N_29282);
and UO_3339 (O_3339,N_29097,N_29243);
and UO_3340 (O_3340,N_29186,N_29150);
and UO_3341 (O_3341,N_29627,N_29002);
nand UO_3342 (O_3342,N_29685,N_29259);
nor UO_3343 (O_3343,N_29275,N_29773);
nand UO_3344 (O_3344,N_29579,N_29283);
or UO_3345 (O_3345,N_29358,N_29766);
and UO_3346 (O_3346,N_29975,N_29012);
or UO_3347 (O_3347,N_29156,N_29963);
nor UO_3348 (O_3348,N_29465,N_29133);
nand UO_3349 (O_3349,N_29639,N_29346);
nand UO_3350 (O_3350,N_29288,N_29754);
xnor UO_3351 (O_3351,N_29921,N_29396);
nand UO_3352 (O_3352,N_29617,N_29429);
nand UO_3353 (O_3353,N_29630,N_29941);
nor UO_3354 (O_3354,N_29997,N_29177);
or UO_3355 (O_3355,N_29597,N_29584);
and UO_3356 (O_3356,N_29688,N_29218);
and UO_3357 (O_3357,N_29855,N_29698);
nor UO_3358 (O_3358,N_29357,N_29230);
nor UO_3359 (O_3359,N_29031,N_29469);
or UO_3360 (O_3360,N_29007,N_29413);
and UO_3361 (O_3361,N_29873,N_29360);
nand UO_3362 (O_3362,N_29300,N_29119);
nor UO_3363 (O_3363,N_29787,N_29792);
or UO_3364 (O_3364,N_29861,N_29772);
xnor UO_3365 (O_3365,N_29901,N_29110);
nand UO_3366 (O_3366,N_29964,N_29031);
xnor UO_3367 (O_3367,N_29229,N_29677);
xor UO_3368 (O_3368,N_29596,N_29770);
or UO_3369 (O_3369,N_29490,N_29917);
nor UO_3370 (O_3370,N_29846,N_29322);
xnor UO_3371 (O_3371,N_29516,N_29721);
and UO_3372 (O_3372,N_29388,N_29542);
or UO_3373 (O_3373,N_29380,N_29112);
nor UO_3374 (O_3374,N_29294,N_29222);
nand UO_3375 (O_3375,N_29588,N_29820);
and UO_3376 (O_3376,N_29928,N_29521);
nor UO_3377 (O_3377,N_29915,N_29802);
or UO_3378 (O_3378,N_29514,N_29066);
nand UO_3379 (O_3379,N_29465,N_29490);
and UO_3380 (O_3380,N_29299,N_29610);
nand UO_3381 (O_3381,N_29348,N_29681);
nor UO_3382 (O_3382,N_29801,N_29799);
xnor UO_3383 (O_3383,N_29292,N_29783);
nor UO_3384 (O_3384,N_29236,N_29695);
nor UO_3385 (O_3385,N_29875,N_29341);
xor UO_3386 (O_3386,N_29397,N_29189);
or UO_3387 (O_3387,N_29661,N_29526);
or UO_3388 (O_3388,N_29999,N_29539);
xor UO_3389 (O_3389,N_29108,N_29448);
nand UO_3390 (O_3390,N_29520,N_29764);
xor UO_3391 (O_3391,N_29296,N_29694);
and UO_3392 (O_3392,N_29173,N_29975);
xnor UO_3393 (O_3393,N_29259,N_29370);
xor UO_3394 (O_3394,N_29033,N_29274);
and UO_3395 (O_3395,N_29651,N_29404);
nand UO_3396 (O_3396,N_29824,N_29276);
and UO_3397 (O_3397,N_29845,N_29811);
or UO_3398 (O_3398,N_29133,N_29780);
and UO_3399 (O_3399,N_29388,N_29306);
or UO_3400 (O_3400,N_29356,N_29321);
nand UO_3401 (O_3401,N_29993,N_29370);
nor UO_3402 (O_3402,N_29863,N_29208);
and UO_3403 (O_3403,N_29548,N_29604);
nand UO_3404 (O_3404,N_29177,N_29337);
or UO_3405 (O_3405,N_29499,N_29833);
and UO_3406 (O_3406,N_29255,N_29284);
nand UO_3407 (O_3407,N_29940,N_29258);
or UO_3408 (O_3408,N_29947,N_29787);
nand UO_3409 (O_3409,N_29524,N_29044);
xor UO_3410 (O_3410,N_29918,N_29297);
nor UO_3411 (O_3411,N_29005,N_29437);
nor UO_3412 (O_3412,N_29848,N_29765);
nand UO_3413 (O_3413,N_29139,N_29718);
and UO_3414 (O_3414,N_29744,N_29224);
xnor UO_3415 (O_3415,N_29809,N_29129);
nor UO_3416 (O_3416,N_29718,N_29502);
xor UO_3417 (O_3417,N_29027,N_29817);
or UO_3418 (O_3418,N_29990,N_29113);
nand UO_3419 (O_3419,N_29802,N_29747);
xor UO_3420 (O_3420,N_29976,N_29543);
and UO_3421 (O_3421,N_29580,N_29299);
xor UO_3422 (O_3422,N_29523,N_29994);
xnor UO_3423 (O_3423,N_29625,N_29110);
and UO_3424 (O_3424,N_29703,N_29901);
or UO_3425 (O_3425,N_29342,N_29043);
xor UO_3426 (O_3426,N_29211,N_29042);
and UO_3427 (O_3427,N_29695,N_29454);
and UO_3428 (O_3428,N_29155,N_29465);
nor UO_3429 (O_3429,N_29499,N_29915);
and UO_3430 (O_3430,N_29926,N_29325);
and UO_3431 (O_3431,N_29238,N_29374);
nor UO_3432 (O_3432,N_29120,N_29329);
or UO_3433 (O_3433,N_29014,N_29435);
nand UO_3434 (O_3434,N_29092,N_29831);
nand UO_3435 (O_3435,N_29662,N_29072);
or UO_3436 (O_3436,N_29598,N_29925);
xnor UO_3437 (O_3437,N_29622,N_29581);
xor UO_3438 (O_3438,N_29535,N_29265);
nor UO_3439 (O_3439,N_29552,N_29689);
nand UO_3440 (O_3440,N_29075,N_29507);
nor UO_3441 (O_3441,N_29316,N_29587);
and UO_3442 (O_3442,N_29415,N_29226);
xnor UO_3443 (O_3443,N_29734,N_29700);
and UO_3444 (O_3444,N_29411,N_29528);
and UO_3445 (O_3445,N_29960,N_29864);
and UO_3446 (O_3446,N_29393,N_29986);
or UO_3447 (O_3447,N_29607,N_29483);
nor UO_3448 (O_3448,N_29969,N_29030);
nor UO_3449 (O_3449,N_29554,N_29501);
nor UO_3450 (O_3450,N_29192,N_29499);
nand UO_3451 (O_3451,N_29803,N_29139);
nor UO_3452 (O_3452,N_29980,N_29570);
xnor UO_3453 (O_3453,N_29496,N_29117);
nand UO_3454 (O_3454,N_29948,N_29491);
nand UO_3455 (O_3455,N_29521,N_29890);
and UO_3456 (O_3456,N_29488,N_29894);
and UO_3457 (O_3457,N_29842,N_29393);
or UO_3458 (O_3458,N_29121,N_29036);
nor UO_3459 (O_3459,N_29710,N_29840);
nor UO_3460 (O_3460,N_29750,N_29084);
xnor UO_3461 (O_3461,N_29940,N_29005);
and UO_3462 (O_3462,N_29167,N_29594);
xnor UO_3463 (O_3463,N_29715,N_29759);
or UO_3464 (O_3464,N_29461,N_29968);
nand UO_3465 (O_3465,N_29200,N_29024);
nor UO_3466 (O_3466,N_29185,N_29538);
nand UO_3467 (O_3467,N_29335,N_29323);
and UO_3468 (O_3468,N_29748,N_29972);
or UO_3469 (O_3469,N_29051,N_29891);
nor UO_3470 (O_3470,N_29786,N_29271);
nand UO_3471 (O_3471,N_29689,N_29283);
or UO_3472 (O_3472,N_29515,N_29882);
xor UO_3473 (O_3473,N_29990,N_29485);
xor UO_3474 (O_3474,N_29774,N_29181);
nor UO_3475 (O_3475,N_29212,N_29512);
or UO_3476 (O_3476,N_29958,N_29789);
xnor UO_3477 (O_3477,N_29124,N_29358);
nor UO_3478 (O_3478,N_29636,N_29526);
nand UO_3479 (O_3479,N_29791,N_29360);
or UO_3480 (O_3480,N_29960,N_29614);
xnor UO_3481 (O_3481,N_29344,N_29166);
nor UO_3482 (O_3482,N_29755,N_29370);
nand UO_3483 (O_3483,N_29111,N_29960);
and UO_3484 (O_3484,N_29883,N_29018);
nand UO_3485 (O_3485,N_29436,N_29279);
or UO_3486 (O_3486,N_29601,N_29344);
and UO_3487 (O_3487,N_29553,N_29722);
nor UO_3488 (O_3488,N_29730,N_29377);
or UO_3489 (O_3489,N_29503,N_29801);
xnor UO_3490 (O_3490,N_29073,N_29651);
and UO_3491 (O_3491,N_29801,N_29972);
xor UO_3492 (O_3492,N_29665,N_29405);
nor UO_3493 (O_3493,N_29725,N_29766);
nand UO_3494 (O_3494,N_29437,N_29044);
xor UO_3495 (O_3495,N_29339,N_29373);
and UO_3496 (O_3496,N_29738,N_29535);
nand UO_3497 (O_3497,N_29112,N_29788);
nand UO_3498 (O_3498,N_29614,N_29680);
or UO_3499 (O_3499,N_29834,N_29430);
endmodule