module basic_1500_15000_2000_5_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_532,In_571);
xor U1 (N_1,In_1378,In_262);
nand U2 (N_2,In_104,In_126);
xor U3 (N_3,In_1397,In_1411);
nor U4 (N_4,In_263,In_1228);
nor U5 (N_5,In_279,In_201);
and U6 (N_6,In_1143,In_401);
and U7 (N_7,In_925,In_620);
nand U8 (N_8,In_528,In_525);
xor U9 (N_9,In_276,In_41);
or U10 (N_10,In_1457,In_1480);
nand U11 (N_11,In_1085,In_834);
and U12 (N_12,In_1366,In_754);
and U13 (N_13,In_940,In_779);
and U14 (N_14,In_1118,In_495);
and U15 (N_15,In_1120,In_357);
and U16 (N_16,In_911,In_893);
and U17 (N_17,In_36,In_151);
nor U18 (N_18,In_773,In_709);
nand U19 (N_19,In_924,In_683);
nand U20 (N_20,In_1356,In_469);
nand U21 (N_21,In_243,In_206);
or U22 (N_22,In_1313,In_188);
xor U23 (N_23,In_857,In_213);
nor U24 (N_24,In_252,In_13);
or U25 (N_25,In_706,In_162);
nor U26 (N_26,In_778,In_83);
and U27 (N_27,In_1316,In_556);
nor U28 (N_28,In_1109,In_403);
nor U29 (N_29,In_356,In_1271);
or U30 (N_30,In_1408,In_740);
nand U31 (N_31,In_300,In_536);
nor U32 (N_32,In_1182,In_247);
nor U33 (N_33,In_1089,In_1068);
nand U34 (N_34,In_1107,In_96);
and U35 (N_35,In_202,In_886);
and U36 (N_36,In_1393,In_1070);
or U37 (N_37,In_759,In_1202);
xnor U38 (N_38,In_49,In_286);
nor U39 (N_39,In_54,In_1223);
nor U40 (N_40,In_1336,In_119);
nor U41 (N_41,In_242,In_394);
nand U42 (N_42,In_187,In_877);
and U43 (N_43,In_1350,In_458);
xor U44 (N_44,In_359,In_261);
nand U45 (N_45,In_170,In_310);
xnor U46 (N_46,In_1155,In_309);
and U47 (N_47,In_806,In_1023);
and U48 (N_48,In_1440,In_579);
nor U49 (N_49,In_1424,In_22);
or U50 (N_50,In_636,In_1133);
nor U51 (N_51,In_1475,In_1226);
or U52 (N_52,In_230,In_1205);
and U53 (N_53,In_623,In_1498);
and U54 (N_54,In_1353,In_913);
nand U55 (N_55,In_685,In_402);
nor U56 (N_56,In_526,In_687);
and U57 (N_57,In_57,In_1465);
or U58 (N_58,In_1087,In_838);
or U59 (N_59,In_796,In_116);
nor U60 (N_60,In_437,In_1293);
nor U61 (N_61,In_1381,In_1317);
nor U62 (N_62,In_374,In_781);
nor U63 (N_63,In_1191,In_208);
or U64 (N_64,In_430,In_541);
or U65 (N_65,In_248,In_757);
and U66 (N_66,In_756,In_210);
or U67 (N_67,In_282,In_1490);
nand U68 (N_68,In_1010,In_852);
and U69 (N_69,In_1362,In_415);
or U70 (N_70,In_1468,In_502);
nand U71 (N_71,In_738,In_179);
or U72 (N_72,In_1448,In_922);
or U73 (N_73,In_652,In_1102);
and U74 (N_74,In_1207,In_292);
xnor U75 (N_75,In_74,In_1215);
or U76 (N_76,In_815,In_86);
or U77 (N_77,In_1281,In_1332);
and U78 (N_78,In_1328,In_963);
xnor U79 (N_79,In_375,In_166);
nor U80 (N_80,In_1265,In_810);
nor U81 (N_81,In_61,In_584);
nor U82 (N_82,In_379,In_828);
nand U83 (N_83,In_1084,In_939);
nor U84 (N_84,In_204,In_1487);
or U85 (N_85,In_1279,In_735);
nor U86 (N_86,In_559,In_100);
nand U87 (N_87,In_1050,In_351);
nor U88 (N_88,In_1462,In_1301);
and U89 (N_89,In_360,In_10);
xnor U90 (N_90,In_81,In_4);
nand U91 (N_91,In_751,In_1288);
nand U92 (N_92,In_589,In_580);
and U93 (N_93,In_1098,In_1277);
nor U94 (N_94,In_1134,In_325);
nand U95 (N_95,In_1062,In_448);
nor U96 (N_96,In_1478,In_544);
nor U97 (N_97,In_957,In_1493);
nand U98 (N_98,In_987,In_1347);
or U99 (N_99,In_1456,In_986);
or U100 (N_100,In_227,In_745);
or U101 (N_101,In_1030,In_499);
nor U102 (N_102,In_741,In_943);
or U103 (N_103,In_395,In_1259);
nor U104 (N_104,In_1167,In_820);
xor U105 (N_105,In_1237,In_1321);
nand U106 (N_106,In_1451,In_529);
or U107 (N_107,In_829,In_1095);
and U108 (N_108,In_144,In_915);
or U109 (N_109,In_624,In_1203);
or U110 (N_110,In_366,In_1492);
nand U111 (N_111,In_1260,In_297);
and U112 (N_112,In_1004,In_138);
xnor U113 (N_113,In_868,In_181);
nand U114 (N_114,In_1398,In_481);
nand U115 (N_115,In_514,In_389);
nor U116 (N_116,In_871,In_207);
nor U117 (N_117,In_148,In_1150);
or U118 (N_118,In_225,In_258);
or U119 (N_119,In_1358,In_960);
or U120 (N_120,In_919,In_1414);
and U121 (N_121,In_1444,In_762);
nor U122 (N_122,In_1446,In_605);
and U123 (N_123,In_1242,In_1272);
nor U124 (N_124,In_555,In_878);
or U125 (N_125,In_324,In_369);
nand U126 (N_126,In_472,In_1142);
or U127 (N_127,In_447,In_197);
xor U128 (N_128,In_133,In_720);
or U129 (N_129,In_90,In_1461);
and U130 (N_130,In_1053,In_327);
or U131 (N_131,In_409,In_1043);
nand U132 (N_132,In_152,In_1429);
or U133 (N_133,In_1141,In_135);
or U134 (N_134,In_221,In_164);
xnor U135 (N_135,In_2,In_681);
nor U136 (N_136,In_1357,In_819);
or U137 (N_137,In_404,In_1015);
and U138 (N_138,In_15,In_643);
nand U139 (N_139,In_1125,In_700);
xnor U140 (N_140,In_274,In_1379);
nor U141 (N_141,In_1229,In_542);
nor U142 (N_142,In_543,In_1322);
or U143 (N_143,In_927,In_546);
nand U144 (N_144,In_937,In_933);
nor U145 (N_145,In_1274,In_51);
and U146 (N_146,In_280,In_855);
and U147 (N_147,In_1076,In_43);
xor U148 (N_148,In_1391,In_1477);
nor U149 (N_149,In_947,In_1310);
nor U150 (N_150,In_1374,In_640);
nor U151 (N_151,In_220,In_244);
xnor U152 (N_152,In_1264,In_1403);
nor U153 (N_153,In_34,In_1359);
xor U154 (N_154,In_1390,In_518);
xor U155 (N_155,In_102,In_1476);
nand U156 (N_156,In_811,In_607);
and U157 (N_157,In_131,In_537);
and U158 (N_158,In_1018,In_20);
nor U159 (N_159,In_35,In_438);
nor U160 (N_160,In_147,In_1427);
nor U161 (N_161,In_265,In_1042);
nand U162 (N_162,In_572,In_482);
xnor U163 (N_163,In_1021,In_634);
or U164 (N_164,In_1256,In_1270);
nor U165 (N_165,In_88,In_731);
and U166 (N_166,In_862,In_1294);
or U167 (N_167,In_1209,In_121);
nor U168 (N_168,In_733,In_1485);
nor U169 (N_169,In_1022,In_1466);
nor U170 (N_170,In_1307,In_386);
nand U171 (N_171,In_991,In_1075);
xnor U172 (N_172,In_920,In_747);
xnor U173 (N_173,In_334,In_1335);
or U174 (N_174,In_874,In_647);
or U175 (N_175,In_229,In_744);
nor U176 (N_176,In_906,In_663);
nor U177 (N_177,In_818,In_507);
nand U178 (N_178,In_1063,In_696);
and U179 (N_179,In_538,In_501);
nand U180 (N_180,In_677,In_979);
or U181 (N_181,In_40,In_672);
nand U182 (N_182,In_949,In_770);
or U183 (N_183,In_1188,In_355);
and U184 (N_184,In_842,In_1096);
or U185 (N_185,In_902,In_1405);
nor U186 (N_186,In_1262,In_446);
nand U187 (N_187,In_965,In_996);
nand U188 (N_188,In_1333,In_308);
nor U189 (N_189,In_1238,In_112);
and U190 (N_190,In_1101,In_851);
nor U191 (N_191,In_1329,In_461);
and U192 (N_192,In_353,In_191);
or U193 (N_193,In_154,In_1304);
or U194 (N_194,In_753,In_273);
nor U195 (N_195,In_1421,In_803);
nand U196 (N_196,In_184,In_644);
and U197 (N_197,In_460,In_1211);
nand U198 (N_198,In_406,In_1069);
xor U199 (N_199,In_711,In_805);
nand U200 (N_200,In_0,In_1132);
nor U201 (N_201,In_516,In_408);
or U202 (N_202,In_1146,In_413);
nand U203 (N_203,In_1020,In_39);
and U204 (N_204,In_392,In_880);
nand U205 (N_205,In_328,In_716);
or U206 (N_206,In_304,In_52);
or U207 (N_207,In_646,In_732);
nor U208 (N_208,In_68,In_178);
nand U209 (N_209,In_824,In_1412);
and U210 (N_210,In_75,In_349);
or U211 (N_211,In_1241,In_1417);
nand U212 (N_212,In_581,In_1436);
or U213 (N_213,In_586,In_671);
nand U214 (N_214,In_944,In_1073);
nand U215 (N_215,In_1305,In_1292);
nor U216 (N_216,In_926,In_434);
or U217 (N_217,In_218,In_952);
xor U218 (N_218,In_1368,In_508);
and U219 (N_219,In_400,In_942);
nor U220 (N_220,In_1311,In_466);
nor U221 (N_221,In_776,In_1257);
nor U222 (N_222,In_710,In_266);
or U223 (N_223,In_938,In_573);
or U224 (N_224,In_109,In_1131);
and U225 (N_225,In_480,In_1437);
xor U226 (N_226,In_1162,In_1151);
nor U227 (N_227,In_698,In_728);
and U228 (N_228,In_895,In_270);
nor U229 (N_229,In_76,In_969);
and U230 (N_230,In_808,In_1136);
xnor U231 (N_231,In_569,In_1140);
and U232 (N_232,In_335,In_908);
nand U233 (N_233,In_761,In_718);
xor U234 (N_234,In_748,In_1097);
and U235 (N_235,In_1326,In_802);
nor U236 (N_236,In_1029,In_330);
or U237 (N_237,In_989,In_124);
and U238 (N_238,In_1005,In_24);
nand U239 (N_239,In_648,In_1110);
nor U240 (N_240,In_739,In_1275);
nand U241 (N_241,In_105,In_697);
or U242 (N_242,In_1036,In_85);
and U243 (N_243,In_990,In_1365);
or U244 (N_244,In_346,In_574);
and U245 (N_245,In_365,In_1467);
nand U246 (N_246,In_1181,In_867);
and U247 (N_247,In_695,In_1320);
nand U248 (N_248,In_250,In_1334);
or U249 (N_249,In_470,In_115);
or U250 (N_250,In_1312,In_433);
and U251 (N_251,In_1491,In_175);
and U252 (N_252,In_752,In_132);
nand U253 (N_253,In_1037,In_494);
or U254 (N_254,In_84,In_419);
nor U255 (N_255,In_553,In_1454);
xnor U256 (N_256,In_577,In_1006);
and U257 (N_257,In_1337,In_1208);
and U258 (N_258,In_576,In_338);
and U259 (N_259,In_1026,In_251);
or U260 (N_260,In_373,In_682);
nor U261 (N_261,In_876,In_606);
nor U262 (N_262,In_339,In_680);
and U263 (N_263,In_897,In_44);
nor U264 (N_264,In_72,In_656);
xnor U265 (N_265,In_301,In_55);
nor U266 (N_266,In_540,In_113);
or U267 (N_267,In_928,In_63);
nand U268 (N_268,In_859,In_1090);
or U269 (N_269,In_734,In_14);
and U270 (N_270,In_176,In_964);
xor U271 (N_271,In_194,In_608);
nand U272 (N_272,In_1173,In_1175);
nor U273 (N_273,In_669,In_567);
nand U274 (N_274,In_699,In_595);
and U275 (N_275,In_332,In_436);
nand U276 (N_276,In_93,In_490);
or U277 (N_277,In_1471,In_984);
and U278 (N_278,In_1168,In_527);
and U279 (N_279,In_1054,In_725);
and U280 (N_280,In_1342,In_625);
nor U281 (N_281,In_423,In_1296);
and U282 (N_282,In_385,In_658);
nor U283 (N_283,In_1106,In_73);
or U284 (N_284,In_1013,In_896);
xor U285 (N_285,In_846,In_281);
and U286 (N_286,In_1383,In_1180);
and U287 (N_287,In_1283,In_420);
nor U288 (N_288,In_167,In_412);
nor U289 (N_289,In_492,In_869);
and U290 (N_290,In_767,In_195);
or U291 (N_291,In_1302,In_600);
and U292 (N_292,In_723,In_1375);
nor U293 (N_293,In_1367,In_1447);
and U294 (N_294,In_1240,In_180);
xnor U295 (N_295,In_789,In_111);
nor U296 (N_296,In_78,In_1082);
nand U297 (N_297,In_1179,In_106);
or U298 (N_298,In_390,In_724);
nor U299 (N_299,In_594,In_117);
or U300 (N_300,In_936,In_995);
nand U301 (N_301,In_228,In_1452);
and U302 (N_302,In_186,In_814);
or U303 (N_303,In_649,In_107);
and U304 (N_304,In_833,In_916);
nor U305 (N_305,In_563,In_189);
and U306 (N_306,In_533,In_323);
and U307 (N_307,In_630,In_1413);
and U308 (N_308,In_1000,In_1276);
nor U309 (N_309,In_58,In_233);
nand U310 (N_310,In_861,In_642);
nor U311 (N_311,In_903,In_294);
and U312 (N_312,In_530,In_712);
or U313 (N_313,In_539,In_1079);
xor U314 (N_314,In_303,In_200);
or U315 (N_315,In_664,In_1399);
nor U316 (N_316,In_1269,In_1244);
and U317 (N_317,In_1033,In_1388);
nor U318 (N_318,In_435,In_427);
or U319 (N_319,In_1348,In_890);
and U320 (N_320,In_449,In_632);
nand U321 (N_321,In_616,In_1172);
and U322 (N_322,In_475,In_491);
nand U323 (N_323,In_451,In_340);
xnor U324 (N_324,In_666,In_585);
xor U325 (N_325,In_976,In_848);
nor U326 (N_326,In_614,In_593);
or U327 (N_327,In_344,In_800);
and U328 (N_328,In_1287,In_1119);
nor U329 (N_329,In_804,In_825);
nand U330 (N_330,In_1138,In_1174);
and U331 (N_331,In_67,In_1177);
nand U332 (N_332,In_1345,In_1031);
xnor U333 (N_333,In_923,In_1420);
or U334 (N_334,In_160,In_1423);
nor U335 (N_335,In_1415,In_760);
nor U336 (N_336,In_882,In_1387);
and U337 (N_337,In_1318,In_56);
and U338 (N_338,In_1161,In_1327);
and U339 (N_339,In_799,In_3);
nand U340 (N_340,In_1112,In_1434);
nand U341 (N_341,In_823,In_343);
or U342 (N_342,In_654,In_1113);
xnor U343 (N_343,In_235,In_1135);
or U344 (N_344,In_153,In_467);
nor U345 (N_345,In_1486,In_764);
nor U346 (N_346,In_97,In_974);
nand U347 (N_347,In_565,In_1443);
or U348 (N_348,In_224,In_1124);
nand U349 (N_349,In_1245,In_239);
or U350 (N_350,In_1396,In_1071);
nor U351 (N_351,In_1212,In_534);
or U352 (N_352,In_1234,In_231);
nand U353 (N_353,In_904,In_524);
and U354 (N_354,In_719,In_418);
or U355 (N_355,In_1370,In_50);
nor U356 (N_356,In_1116,In_477);
or U357 (N_357,In_1494,In_80);
or U358 (N_358,In_245,In_452);
and U359 (N_359,In_1278,In_602);
nor U360 (N_360,In_517,In_892);
nor U361 (N_361,In_1267,In_839);
and U362 (N_362,In_238,In_156);
or U363 (N_363,In_889,In_1230);
or U364 (N_364,In_1239,In_885);
or U365 (N_365,In_463,In_705);
and U366 (N_366,In_1066,In_879);
and U367 (N_367,In_165,In_1011);
nor U368 (N_368,In_171,In_442);
or U369 (N_369,In_1057,In_1380);
and U370 (N_370,In_407,In_707);
nor U371 (N_371,In_199,In_651);
nor U372 (N_372,In_1210,In_758);
and U373 (N_373,In_485,In_959);
or U374 (N_374,In_1016,In_1221);
nor U375 (N_375,In_278,In_429);
nand U376 (N_376,In_256,In_590);
or U377 (N_377,In_535,In_547);
or U378 (N_378,In_1371,In_1341);
nor U379 (N_379,In_1213,In_305);
nor U380 (N_380,In_1419,In_561);
and U381 (N_381,In_450,In_440);
nor U382 (N_382,In_489,In_1499);
or U383 (N_383,In_259,In_1198);
xor U384 (N_384,In_635,In_500);
nor U385 (N_385,In_617,In_16);
nor U386 (N_386,In_1183,In_1196);
nand U387 (N_387,In_275,In_322);
nor U388 (N_388,In_1377,In_424);
nand U389 (N_389,In_341,In_1450);
and U390 (N_390,In_1472,In_907);
nand U391 (N_391,In_854,In_1236);
and U392 (N_392,In_807,In_844);
and U393 (N_393,In_772,In_793);
xnor U394 (N_394,In_691,In_596);
nor U395 (N_395,In_1280,In_1343);
or U396 (N_396,In_1045,In_240);
and U397 (N_397,In_578,In_136);
or U398 (N_398,In_841,In_255);
and U399 (N_399,In_388,In_860);
nor U400 (N_400,In_1268,In_18);
or U401 (N_401,In_1459,In_1048);
nor U402 (N_402,In_174,In_587);
or U403 (N_403,In_32,In_30);
nand U404 (N_404,In_702,In_765);
nand U405 (N_405,In_575,In_704);
or U406 (N_406,In_597,In_1035);
and U407 (N_407,In_750,In_237);
or U408 (N_408,In_284,In_271);
nor U409 (N_409,In_383,In_1159);
nor U410 (N_410,In_592,In_1483);
nand U411 (N_411,In_746,In_708);
xor U412 (N_412,In_150,In_1139);
nor U413 (N_413,In_1441,In_791);
or U414 (N_414,In_619,In_158);
or U415 (N_415,In_1064,In_417);
and U416 (N_416,In_82,In_333);
and U417 (N_417,In_1204,In_1);
nor U418 (N_418,In_1438,In_684);
and U419 (N_419,In_342,In_1289);
nand U420 (N_420,In_474,In_254);
nor U421 (N_421,In_1290,In_633);
xor U422 (N_422,In_1263,In_319);
and U423 (N_423,In_866,In_405);
and U424 (N_424,In_1189,In_899);
xnor U425 (N_425,In_1418,In_326);
and U426 (N_426,In_826,In_1014);
and U427 (N_427,In_384,In_444);
nand U428 (N_428,In_1349,In_693);
or U429 (N_429,In_1319,In_1474);
or U430 (N_430,In_931,In_831);
or U431 (N_431,In_506,In_1364);
nand U432 (N_432,In_1086,In_566);
nand U433 (N_433,In_416,In_531);
nand U434 (N_434,In_1148,In_42);
nand U435 (N_435,In_935,In_142);
and U436 (N_436,In_679,In_473);
xnor U437 (N_437,In_288,In_604);
nor U438 (N_438,In_1430,In_1416);
xnor U439 (N_439,In_881,In_123);
and U440 (N_440,In_223,In_843);
or U441 (N_441,In_582,In_603);
nor U442 (N_442,In_557,In_670);
nand U443 (N_443,In_1130,In_146);
nor U444 (N_444,In_1017,In_715);
or U445 (N_445,In_1484,In_1195);
nand U446 (N_446,In_1315,In_1147);
or U447 (N_447,In_1473,In_613);
nand U448 (N_448,In_914,In_521);
or U449 (N_449,In_362,In_512);
or U450 (N_450,In_377,In_1410);
nand U451 (N_451,In_982,In_1382);
or U452 (N_452,In_290,In_497);
and U453 (N_453,In_1426,In_350);
or U454 (N_454,In_1369,In_95);
nor U455 (N_455,In_638,In_1104);
nand U456 (N_456,In_1115,In_289);
and U457 (N_457,In_909,In_769);
and U458 (N_458,In_850,In_662);
nand U459 (N_459,In_1093,In_1051);
or U460 (N_460,In_1024,In_380);
and U461 (N_461,In_1308,In_898);
or U462 (N_462,In_376,In_1220);
or U463 (N_463,In_992,In_971);
and U464 (N_464,In_214,In_37);
or U465 (N_465,In_967,In_794);
and U466 (N_466,In_311,In_1144);
and U467 (N_467,In_883,In_1009);
xnor U468 (N_468,In_441,In_505);
nand U469 (N_469,In_1072,In_1291);
and U470 (N_470,In_1165,In_1249);
nor U471 (N_471,In_1060,In_583);
nor U472 (N_472,In_62,In_1394);
and U473 (N_473,In_94,In_714);
xor U474 (N_474,In_1100,In_849);
nand U475 (N_475,In_777,In_961);
or U476 (N_476,In_1061,In_945);
or U477 (N_477,In_168,In_622);
or U478 (N_478,In_872,In_29);
nor U479 (N_479,In_432,In_127);
and U480 (N_480,In_414,In_551);
or U481 (N_481,In_1186,In_1284);
and U482 (N_482,In_894,In_721);
xor U483 (N_483,In_1355,In_6);
xnor U484 (N_484,In_337,In_47);
nor U485 (N_485,In_125,In_382);
nor U486 (N_486,In_293,In_856);
nor U487 (N_487,In_372,In_550);
nor U488 (N_488,In_1235,In_1481);
nor U489 (N_489,In_1433,In_410);
and U490 (N_490,In_285,In_1128);
and U491 (N_491,In_978,In_422);
nand U492 (N_492,In_599,In_9);
nor U493 (N_493,In_1149,In_503);
and U494 (N_494,In_784,In_345);
nor U495 (N_495,In_26,In_69);
nor U496 (N_496,In_722,In_785);
nand U497 (N_497,In_790,In_498);
xor U498 (N_498,In_997,In_510);
and U499 (N_499,In_198,In_1246);
nand U500 (N_500,In_177,In_190);
nand U501 (N_501,In_1250,In_295);
nand U502 (N_502,In_1435,In_31);
nand U503 (N_503,In_713,In_1121);
nor U504 (N_504,In_610,In_591);
nor U505 (N_505,In_1254,In_941);
nor U506 (N_506,In_968,In_1298);
or U507 (N_507,In_774,In_1297);
and U508 (N_508,In_101,In_668);
xnor U509 (N_509,In_12,In_291);
nor U510 (N_510,In_1145,In_493);
nand U511 (N_511,In_970,In_378);
and U512 (N_512,In_520,In_99);
or U513 (N_513,In_901,In_1360);
nand U514 (N_514,In_439,In_108);
nand U515 (N_515,In_1152,In_797);
nor U516 (N_516,In_1123,In_917);
and U517 (N_517,In_1495,In_686);
and U518 (N_518,In_149,In_1432);
nand U519 (N_519,In_1058,In_455);
nor U520 (N_520,In_1187,In_1224);
xor U521 (N_521,In_1386,In_798);
nand U522 (N_522,In_1199,In_1400);
and U523 (N_523,In_766,In_511);
nor U524 (N_524,In_873,In_1083);
xnor U525 (N_525,In_1169,In_1346);
nor U526 (N_526,In_361,In_912);
or U527 (N_527,In_562,In_320);
nand U528 (N_528,In_23,In_1339);
xnor U529 (N_529,In_523,In_316);
and U530 (N_530,In_130,In_1171);
and U531 (N_531,In_958,In_19);
or U532 (N_532,In_212,In_1081);
nand U533 (N_533,In_269,In_118);
nor U534 (N_534,In_471,In_155);
and U535 (N_535,In_476,In_205);
and U536 (N_536,In_1194,In_5);
xor U537 (N_537,In_317,In_203);
nor U538 (N_538,In_185,In_1439);
nand U539 (N_539,In_788,In_628);
nor U540 (N_540,In_1074,In_629);
or U541 (N_541,In_318,In_657);
nor U542 (N_542,In_1217,In_813);
and U543 (N_543,In_929,In_426);
xnor U544 (N_544,In_977,In_1025);
nand U545 (N_545,In_688,In_64);
and U546 (N_546,In_358,In_1201);
or U547 (N_547,In_1306,In_79);
nor U548 (N_548,In_627,In_570);
or U549 (N_549,In_268,In_1185);
or U550 (N_550,In_817,In_232);
nand U551 (N_551,In_771,In_1049);
nor U552 (N_552,In_216,In_425);
xnor U553 (N_553,In_1266,In_980);
nand U554 (N_554,In_283,In_1314);
or U555 (N_555,In_953,In_1225);
nand U556 (N_556,In_639,In_809);
or U557 (N_557,In_1323,In_910);
nor U558 (N_558,In_730,In_1137);
or U559 (N_559,In_1114,In_645);
and U560 (N_560,In_1157,In_621);
and U561 (N_561,In_727,In_1406);
and U562 (N_562,In_701,In_479);
nand U563 (N_563,In_1046,In_717);
nor U564 (N_564,In_38,In_956);
nand U565 (N_565,In_1038,In_196);
nand U566 (N_566,In_736,In_1056);
and U567 (N_567,In_1309,In_694);
nand U568 (N_568,In_1232,In_1092);
or U569 (N_569,In_1041,In_558);
nand U570 (N_570,In_1324,In_1219);
nor U571 (N_571,In_1482,In_486);
and U572 (N_572,In_918,In_674);
and U573 (N_573,In_1453,In_1285);
nor U574 (N_574,In_1344,In_267);
nand U575 (N_575,In_1040,In_1197);
xor U576 (N_576,In_1166,In_1354);
or U577 (N_577,In_1214,In_21);
and U578 (N_578,In_655,In_128);
xnor U579 (N_579,In_302,In_993);
and U580 (N_580,In_1300,In_329);
nand U581 (N_581,In_832,In_1080);
and U582 (N_582,In_858,In_1184);
and U583 (N_583,In_89,In_891);
nor U584 (N_584,In_122,In_137);
or U585 (N_585,In_161,In_665);
nand U586 (N_586,In_487,In_1352);
and U587 (N_587,In_1361,In_336);
and U588 (N_588,In_98,In_1401);
xnor U589 (N_589,In_1470,In_1178);
nand U590 (N_590,In_1248,In_1055);
nand U591 (N_591,In_863,In_552);
nand U592 (N_592,In_737,In_1044);
nor U593 (N_593,In_519,In_900);
nor U594 (N_594,In_192,In_1258);
nor U595 (N_595,In_1460,In_835);
or U596 (N_596,In_659,In_249);
and U597 (N_597,In_1442,In_1028);
xor U598 (N_598,In_70,In_1282);
nor U599 (N_599,In_830,In_387);
and U600 (N_600,In_981,In_763);
nor U601 (N_601,In_1002,In_884);
and U602 (N_602,In_1216,In_431);
or U603 (N_603,In_1088,In_241);
xnor U604 (N_604,In_1153,In_615);
xnor U605 (N_605,In_887,In_1407);
xnor U606 (N_606,In_465,In_364);
and U607 (N_607,In_222,In_837);
nor U608 (N_608,In_816,In_66);
and U609 (N_609,In_609,In_87);
nor U610 (N_610,In_370,In_236);
nor U611 (N_611,In_549,In_331);
nand U612 (N_612,In_234,In_1170);
nor U613 (N_613,In_445,In_313);
nand U614 (N_614,In_845,In_139);
or U615 (N_615,In_77,In_1469);
nor U616 (N_616,In_246,In_397);
nand U617 (N_617,In_675,In_1261);
nor U618 (N_618,In_676,In_637);
nor U619 (N_619,In_368,In_65);
or U620 (N_620,In_1372,In_1019);
nor U621 (N_621,In_60,In_1247);
and U622 (N_622,In_847,In_453);
and U623 (N_623,In_611,In_1340);
or U624 (N_624,In_1385,In_661);
nand U625 (N_625,In_786,In_618);
nor U626 (N_626,In_354,In_143);
and U627 (N_627,In_399,In_783);
nor U628 (N_628,In_1331,In_1154);
nand U629 (N_629,In_780,In_755);
or U630 (N_630,In_729,In_1445);
or U631 (N_631,In_1330,In_114);
or U632 (N_632,In_159,In_264);
nor U633 (N_633,In_836,In_307);
and U634 (N_634,In_1078,In_129);
xnor U635 (N_635,In_875,In_253);
nand U636 (N_636,In_1376,In_457);
nor U637 (N_637,In_398,In_504);
xor U638 (N_638,In_1039,In_905);
or U639 (N_639,In_1122,In_1488);
nand U640 (N_640,In_1422,In_1067);
nand U641 (N_641,In_272,In_1449);
nand U642 (N_642,In_775,In_948);
or U643 (N_643,In_921,In_973);
or U644 (N_644,In_1163,In_496);
xor U645 (N_645,In_994,In_1392);
or U646 (N_646,In_33,In_934);
nor U647 (N_647,In_1243,In_955);
or U648 (N_648,In_193,In_812);
nor U649 (N_649,In_673,In_1363);
nand U650 (N_650,In_1425,In_314);
and U651 (N_651,In_975,In_25);
and U652 (N_652,In_371,In_1001);
or U653 (N_653,In_1091,In_888);
and U654 (N_654,In_1111,In_689);
and U655 (N_655,In_985,In_1489);
or U656 (N_656,In_827,In_478);
nor U657 (N_657,In_703,In_998);
or U658 (N_658,In_141,In_792);
xor U659 (N_659,In_367,In_554);
and U660 (N_660,In_443,In_183);
or U661 (N_661,In_140,In_690);
nand U662 (N_662,In_27,In_588);
and U663 (N_663,In_1034,In_1252);
xnor U664 (N_664,In_983,In_110);
and U665 (N_665,In_795,In_954);
nand U666 (N_666,In_1032,In_1227);
nand U667 (N_667,In_1402,In_1108);
and U668 (N_668,In_7,In_1325);
or U669 (N_669,In_459,In_363);
and U670 (N_670,In_483,In_145);
or U671 (N_671,In_568,In_17);
and U672 (N_672,In_513,In_1027);
or U673 (N_673,In_660,In_1160);
nor U674 (N_674,In_1464,In_1007);
nand U675 (N_675,In_801,In_840);
nor U676 (N_676,In_853,In_1384);
nand U677 (N_677,In_53,In_1338);
nand U678 (N_678,In_1233,In_598);
and U679 (N_679,In_1463,In_1105);
or U680 (N_680,In_1431,In_1373);
nand U681 (N_681,In_522,In_601);
or U682 (N_682,In_91,In_1156);
xor U683 (N_683,In_103,In_428);
and U684 (N_684,In_612,In_157);
nor U685 (N_685,In_1126,In_1251);
nor U686 (N_686,In_999,In_468);
or U687 (N_687,In_1286,In_211);
or U688 (N_688,In_631,In_1455);
nor U689 (N_689,In_1129,In_1351);
or U690 (N_690,In_951,In_641);
nand U691 (N_691,In_219,In_287);
nand U692 (N_692,In_456,In_421);
or U693 (N_693,In_726,In_209);
nand U694 (N_694,In_352,In_321);
xnor U695 (N_695,In_870,In_1497);
xnor U696 (N_696,In_299,In_1395);
nand U697 (N_697,In_217,In_1052);
or U698 (N_698,In_1158,In_1255);
nor U699 (N_699,In_822,In_11);
nand U700 (N_700,In_650,In_515);
nand U701 (N_701,In_391,In_1479);
nand U702 (N_702,In_787,In_28);
and U703 (N_703,In_742,In_260);
or U704 (N_704,In_1103,In_1099);
nor U705 (N_705,In_315,In_1176);
nand U706 (N_706,In_932,In_678);
nand U707 (N_707,In_454,In_1299);
and U708 (N_708,In_411,In_59);
and U709 (N_709,In_396,In_1409);
nand U710 (N_710,In_173,In_1065);
nand U711 (N_711,In_1117,In_312);
nand U712 (N_712,In_1496,In_743);
nand U713 (N_713,In_865,In_930);
nand U714 (N_714,In_163,In_1389);
and U715 (N_715,In_626,In_1012);
nor U716 (N_716,In_1458,In_45);
and U717 (N_717,In_1222,In_46);
nand U718 (N_718,In_92,In_1206);
nand U719 (N_719,In_488,In_768);
nand U720 (N_720,In_464,In_1200);
nor U721 (N_721,In_548,In_1127);
and U722 (N_722,In_48,In_1193);
nand U723 (N_723,In_257,In_692);
and U724 (N_724,In_950,In_1218);
and U725 (N_725,In_1047,In_946);
or U726 (N_726,In_484,In_1190);
and U727 (N_727,In_215,In_1295);
nand U728 (N_728,In_962,In_393);
or U729 (N_729,In_988,In_306);
nor U730 (N_730,In_1164,In_182);
nand U731 (N_731,In_667,In_972);
xor U732 (N_732,In_381,In_509);
nor U733 (N_733,In_1253,In_226);
and U734 (N_734,In_1273,In_120);
nand U735 (N_735,In_277,In_8);
xor U736 (N_736,In_1008,In_821);
nor U737 (N_737,In_1077,In_1059);
and U738 (N_738,In_749,In_1404);
nor U739 (N_739,In_462,In_560);
or U740 (N_740,In_1003,In_134);
nor U741 (N_741,In_1428,In_1192);
nor U742 (N_742,In_172,In_864);
nand U743 (N_743,In_298,In_169);
and U744 (N_744,In_1094,In_1303);
nand U745 (N_745,In_1231,In_296);
or U746 (N_746,In_564,In_966);
or U747 (N_747,In_545,In_348);
nor U748 (N_748,In_782,In_653);
or U749 (N_749,In_71,In_347);
nand U750 (N_750,In_282,In_992);
or U751 (N_751,In_1316,In_478);
nand U752 (N_752,In_1213,In_407);
nor U753 (N_753,In_1124,In_265);
or U754 (N_754,In_1338,In_4);
and U755 (N_755,In_1467,In_1302);
and U756 (N_756,In_76,In_691);
and U757 (N_757,In_992,In_980);
nand U758 (N_758,In_1239,In_665);
and U759 (N_759,In_1245,In_1497);
and U760 (N_760,In_1323,In_142);
nor U761 (N_761,In_767,In_1370);
nand U762 (N_762,In_851,In_1095);
nor U763 (N_763,In_609,In_1366);
nor U764 (N_764,In_1466,In_641);
nor U765 (N_765,In_335,In_198);
xnor U766 (N_766,In_1438,In_244);
or U767 (N_767,In_629,In_809);
nand U768 (N_768,In_201,In_1232);
or U769 (N_769,In_267,In_338);
and U770 (N_770,In_1169,In_1284);
and U771 (N_771,In_356,In_1432);
nand U772 (N_772,In_1498,In_1235);
nor U773 (N_773,In_478,In_110);
or U774 (N_774,In_494,In_151);
nor U775 (N_775,In_1368,In_360);
or U776 (N_776,In_864,In_191);
nor U777 (N_777,In_61,In_409);
and U778 (N_778,In_1436,In_512);
nor U779 (N_779,In_1416,In_1201);
and U780 (N_780,In_364,In_1305);
nor U781 (N_781,In_337,In_856);
nor U782 (N_782,In_1302,In_342);
nand U783 (N_783,In_1130,In_575);
and U784 (N_784,In_41,In_918);
nand U785 (N_785,In_768,In_827);
or U786 (N_786,In_1376,In_1232);
or U787 (N_787,In_254,In_268);
and U788 (N_788,In_1128,In_1496);
nand U789 (N_789,In_1267,In_513);
nand U790 (N_790,In_961,In_570);
and U791 (N_791,In_139,In_1434);
nand U792 (N_792,In_49,In_1247);
or U793 (N_793,In_852,In_251);
nor U794 (N_794,In_156,In_1248);
and U795 (N_795,In_977,In_547);
xnor U796 (N_796,In_964,In_1494);
nor U797 (N_797,In_758,In_227);
nor U798 (N_798,In_346,In_669);
nand U799 (N_799,In_1144,In_188);
or U800 (N_800,In_783,In_574);
nor U801 (N_801,In_593,In_689);
or U802 (N_802,In_698,In_1033);
or U803 (N_803,In_957,In_741);
nand U804 (N_804,In_1078,In_484);
nand U805 (N_805,In_1275,In_645);
or U806 (N_806,In_1217,In_381);
nand U807 (N_807,In_58,In_241);
and U808 (N_808,In_948,In_719);
nor U809 (N_809,In_451,In_913);
nor U810 (N_810,In_65,In_1300);
nand U811 (N_811,In_52,In_799);
nand U812 (N_812,In_1422,In_386);
nand U813 (N_813,In_1236,In_1282);
or U814 (N_814,In_1084,In_83);
nor U815 (N_815,In_648,In_686);
and U816 (N_816,In_1350,In_913);
nand U817 (N_817,In_1481,In_282);
nand U818 (N_818,In_1217,In_635);
nor U819 (N_819,In_1203,In_1490);
nand U820 (N_820,In_1443,In_56);
nor U821 (N_821,In_823,In_105);
and U822 (N_822,In_1467,In_45);
nand U823 (N_823,In_954,In_546);
or U824 (N_824,In_3,In_1452);
nor U825 (N_825,In_568,In_1134);
and U826 (N_826,In_69,In_201);
and U827 (N_827,In_154,In_217);
and U828 (N_828,In_705,In_983);
or U829 (N_829,In_766,In_1320);
and U830 (N_830,In_604,In_1423);
and U831 (N_831,In_1083,In_987);
nand U832 (N_832,In_286,In_695);
nand U833 (N_833,In_385,In_977);
or U834 (N_834,In_162,In_278);
xnor U835 (N_835,In_1090,In_879);
or U836 (N_836,In_113,In_276);
nor U837 (N_837,In_1162,In_431);
or U838 (N_838,In_846,In_1408);
and U839 (N_839,In_1407,In_1477);
nand U840 (N_840,In_581,In_54);
nand U841 (N_841,In_645,In_9);
and U842 (N_842,In_913,In_9);
or U843 (N_843,In_1462,In_1210);
or U844 (N_844,In_889,In_955);
or U845 (N_845,In_518,In_861);
and U846 (N_846,In_1086,In_50);
and U847 (N_847,In_936,In_57);
or U848 (N_848,In_566,In_1310);
nand U849 (N_849,In_516,In_1141);
or U850 (N_850,In_277,In_303);
or U851 (N_851,In_333,In_801);
nor U852 (N_852,In_491,In_894);
or U853 (N_853,In_1236,In_398);
or U854 (N_854,In_616,In_435);
nand U855 (N_855,In_565,In_473);
and U856 (N_856,In_397,In_897);
nor U857 (N_857,In_316,In_1485);
nor U858 (N_858,In_98,In_1024);
and U859 (N_859,In_335,In_1288);
nand U860 (N_860,In_1096,In_235);
nand U861 (N_861,In_1497,In_666);
nand U862 (N_862,In_470,In_1400);
nor U863 (N_863,In_121,In_393);
and U864 (N_864,In_537,In_282);
nor U865 (N_865,In_370,In_1471);
and U866 (N_866,In_1252,In_1227);
and U867 (N_867,In_147,In_669);
nor U868 (N_868,In_1323,In_199);
xor U869 (N_869,In_33,In_1058);
and U870 (N_870,In_188,In_1374);
nor U871 (N_871,In_1142,In_76);
and U872 (N_872,In_1298,In_13);
and U873 (N_873,In_740,In_595);
and U874 (N_874,In_9,In_135);
nand U875 (N_875,In_1208,In_1205);
and U876 (N_876,In_507,In_1459);
nor U877 (N_877,In_805,In_761);
xnor U878 (N_878,In_175,In_314);
nand U879 (N_879,In_864,In_897);
xnor U880 (N_880,In_380,In_1233);
or U881 (N_881,In_486,In_442);
nand U882 (N_882,In_1040,In_1260);
or U883 (N_883,In_320,In_433);
and U884 (N_884,In_1039,In_752);
xnor U885 (N_885,In_935,In_355);
or U886 (N_886,In_1122,In_180);
nor U887 (N_887,In_9,In_368);
nand U888 (N_888,In_900,In_361);
and U889 (N_889,In_605,In_1275);
nor U890 (N_890,In_1106,In_1212);
nand U891 (N_891,In_206,In_700);
nand U892 (N_892,In_1448,In_819);
nor U893 (N_893,In_1398,In_298);
nor U894 (N_894,In_508,In_325);
xnor U895 (N_895,In_352,In_24);
or U896 (N_896,In_1296,In_1441);
nor U897 (N_897,In_12,In_1408);
xor U898 (N_898,In_1237,In_604);
nand U899 (N_899,In_785,In_610);
nand U900 (N_900,In_404,In_990);
nand U901 (N_901,In_364,In_1066);
nor U902 (N_902,In_1249,In_1255);
or U903 (N_903,In_290,In_633);
nor U904 (N_904,In_611,In_153);
or U905 (N_905,In_543,In_451);
and U906 (N_906,In_447,In_810);
nor U907 (N_907,In_1206,In_41);
or U908 (N_908,In_477,In_1143);
and U909 (N_909,In_1364,In_232);
and U910 (N_910,In_501,In_828);
nand U911 (N_911,In_820,In_841);
or U912 (N_912,In_990,In_570);
nand U913 (N_913,In_305,In_304);
nor U914 (N_914,In_802,In_212);
or U915 (N_915,In_533,In_293);
nor U916 (N_916,In_338,In_1092);
and U917 (N_917,In_155,In_738);
xor U918 (N_918,In_541,In_1139);
nor U919 (N_919,In_1186,In_739);
nand U920 (N_920,In_332,In_806);
or U921 (N_921,In_1464,In_1203);
xor U922 (N_922,In_875,In_700);
and U923 (N_923,In_552,In_868);
xor U924 (N_924,In_801,In_1002);
nand U925 (N_925,In_166,In_1323);
or U926 (N_926,In_1366,In_424);
or U927 (N_927,In_884,In_849);
nor U928 (N_928,In_81,In_458);
and U929 (N_929,In_1076,In_524);
nand U930 (N_930,In_1335,In_1448);
or U931 (N_931,In_955,In_486);
nor U932 (N_932,In_1182,In_48);
or U933 (N_933,In_530,In_766);
nor U934 (N_934,In_865,In_1242);
nand U935 (N_935,In_23,In_1326);
or U936 (N_936,In_1011,In_532);
nand U937 (N_937,In_1048,In_25);
and U938 (N_938,In_426,In_269);
and U939 (N_939,In_925,In_221);
nor U940 (N_940,In_378,In_241);
nand U941 (N_941,In_1396,In_1068);
nor U942 (N_942,In_135,In_1401);
and U943 (N_943,In_1446,In_653);
and U944 (N_944,In_1225,In_458);
and U945 (N_945,In_653,In_776);
nand U946 (N_946,In_1484,In_251);
or U947 (N_947,In_377,In_128);
nand U948 (N_948,In_891,In_824);
and U949 (N_949,In_1365,In_396);
and U950 (N_950,In_3,In_360);
and U951 (N_951,In_971,In_1398);
xnor U952 (N_952,In_788,In_114);
or U953 (N_953,In_1486,In_1196);
and U954 (N_954,In_980,In_381);
xnor U955 (N_955,In_598,In_468);
nor U956 (N_956,In_812,In_1420);
nor U957 (N_957,In_333,In_934);
or U958 (N_958,In_274,In_1385);
or U959 (N_959,In_54,In_519);
and U960 (N_960,In_757,In_574);
or U961 (N_961,In_917,In_1385);
xnor U962 (N_962,In_836,In_831);
nand U963 (N_963,In_975,In_261);
or U964 (N_964,In_1128,In_507);
or U965 (N_965,In_678,In_580);
or U966 (N_966,In_91,In_823);
or U967 (N_967,In_1075,In_89);
xor U968 (N_968,In_807,In_587);
and U969 (N_969,In_643,In_1285);
nand U970 (N_970,In_198,In_1207);
or U971 (N_971,In_131,In_1471);
or U972 (N_972,In_1089,In_133);
and U973 (N_973,In_904,In_185);
or U974 (N_974,In_1125,In_803);
nor U975 (N_975,In_1457,In_480);
nor U976 (N_976,In_410,In_687);
and U977 (N_977,In_585,In_968);
or U978 (N_978,In_483,In_578);
nand U979 (N_979,In_703,In_1145);
nand U980 (N_980,In_1060,In_804);
xor U981 (N_981,In_711,In_1203);
or U982 (N_982,In_1254,In_215);
and U983 (N_983,In_1248,In_1120);
nand U984 (N_984,In_666,In_1125);
nor U985 (N_985,In_196,In_377);
and U986 (N_986,In_572,In_574);
nand U987 (N_987,In_241,In_201);
xor U988 (N_988,In_1412,In_1406);
and U989 (N_989,In_1122,In_224);
nor U990 (N_990,In_1278,In_1005);
nand U991 (N_991,In_3,In_550);
nor U992 (N_992,In_1243,In_1067);
or U993 (N_993,In_69,In_753);
nand U994 (N_994,In_123,In_1427);
nand U995 (N_995,In_377,In_799);
nor U996 (N_996,In_19,In_839);
nor U997 (N_997,In_180,In_570);
or U998 (N_998,In_832,In_846);
or U999 (N_999,In_288,In_601);
or U1000 (N_1000,In_458,In_827);
nand U1001 (N_1001,In_599,In_465);
or U1002 (N_1002,In_814,In_1469);
or U1003 (N_1003,In_1476,In_270);
nand U1004 (N_1004,In_1376,In_168);
and U1005 (N_1005,In_72,In_741);
and U1006 (N_1006,In_293,In_1112);
nor U1007 (N_1007,In_681,In_806);
nor U1008 (N_1008,In_1254,In_1459);
nand U1009 (N_1009,In_169,In_695);
nor U1010 (N_1010,In_269,In_1306);
and U1011 (N_1011,In_790,In_1127);
nor U1012 (N_1012,In_344,In_1129);
nand U1013 (N_1013,In_25,In_981);
or U1014 (N_1014,In_720,In_440);
nand U1015 (N_1015,In_277,In_187);
nand U1016 (N_1016,In_193,In_1003);
xor U1017 (N_1017,In_179,In_832);
and U1018 (N_1018,In_965,In_382);
and U1019 (N_1019,In_484,In_319);
or U1020 (N_1020,In_298,In_325);
xnor U1021 (N_1021,In_443,In_104);
or U1022 (N_1022,In_1438,In_450);
nand U1023 (N_1023,In_864,In_462);
or U1024 (N_1024,In_1301,In_448);
xnor U1025 (N_1025,In_746,In_894);
nand U1026 (N_1026,In_110,In_1394);
nor U1027 (N_1027,In_84,In_735);
or U1028 (N_1028,In_1026,In_781);
nor U1029 (N_1029,In_1445,In_1394);
and U1030 (N_1030,In_1224,In_684);
nand U1031 (N_1031,In_888,In_940);
and U1032 (N_1032,In_429,In_181);
and U1033 (N_1033,In_81,In_1376);
and U1034 (N_1034,In_1273,In_130);
or U1035 (N_1035,In_857,In_616);
xnor U1036 (N_1036,In_901,In_1234);
or U1037 (N_1037,In_1063,In_70);
or U1038 (N_1038,In_590,In_870);
nand U1039 (N_1039,In_523,In_606);
and U1040 (N_1040,In_1465,In_211);
nor U1041 (N_1041,In_467,In_417);
nand U1042 (N_1042,In_395,In_921);
nand U1043 (N_1043,In_1171,In_1090);
nand U1044 (N_1044,In_1078,In_1212);
and U1045 (N_1045,In_385,In_688);
nand U1046 (N_1046,In_705,In_35);
and U1047 (N_1047,In_303,In_610);
nand U1048 (N_1048,In_425,In_1112);
and U1049 (N_1049,In_653,In_1104);
or U1050 (N_1050,In_1166,In_848);
and U1051 (N_1051,In_312,In_253);
xnor U1052 (N_1052,In_907,In_1251);
xor U1053 (N_1053,In_667,In_370);
and U1054 (N_1054,In_1499,In_1081);
nand U1055 (N_1055,In_1493,In_422);
or U1056 (N_1056,In_703,In_484);
and U1057 (N_1057,In_1404,In_71);
or U1058 (N_1058,In_1486,In_211);
and U1059 (N_1059,In_1450,In_1226);
nor U1060 (N_1060,In_940,In_629);
and U1061 (N_1061,In_1395,In_1048);
and U1062 (N_1062,In_1176,In_61);
nor U1063 (N_1063,In_553,In_169);
nor U1064 (N_1064,In_61,In_469);
nand U1065 (N_1065,In_403,In_851);
nor U1066 (N_1066,In_635,In_1053);
and U1067 (N_1067,In_33,In_674);
xnor U1068 (N_1068,In_970,In_314);
nand U1069 (N_1069,In_1160,In_1290);
and U1070 (N_1070,In_416,In_1211);
or U1071 (N_1071,In_134,In_1335);
xnor U1072 (N_1072,In_190,In_925);
or U1073 (N_1073,In_158,In_140);
nor U1074 (N_1074,In_251,In_462);
or U1075 (N_1075,In_214,In_299);
nand U1076 (N_1076,In_1114,In_261);
and U1077 (N_1077,In_553,In_829);
or U1078 (N_1078,In_1075,In_253);
or U1079 (N_1079,In_153,In_1157);
and U1080 (N_1080,In_189,In_1233);
nor U1081 (N_1081,In_601,In_142);
and U1082 (N_1082,In_328,In_1380);
nand U1083 (N_1083,In_426,In_129);
nor U1084 (N_1084,In_908,In_1204);
and U1085 (N_1085,In_996,In_1033);
or U1086 (N_1086,In_724,In_62);
and U1087 (N_1087,In_1306,In_964);
or U1088 (N_1088,In_1355,In_1421);
nand U1089 (N_1089,In_408,In_1071);
or U1090 (N_1090,In_849,In_1027);
or U1091 (N_1091,In_1433,In_721);
xnor U1092 (N_1092,In_697,In_835);
nor U1093 (N_1093,In_270,In_1111);
xor U1094 (N_1094,In_307,In_306);
nand U1095 (N_1095,In_704,In_307);
nand U1096 (N_1096,In_495,In_1290);
nor U1097 (N_1097,In_433,In_733);
or U1098 (N_1098,In_591,In_104);
nor U1099 (N_1099,In_512,In_91);
nand U1100 (N_1100,In_675,In_25);
and U1101 (N_1101,In_1234,In_1426);
or U1102 (N_1102,In_938,In_232);
nor U1103 (N_1103,In_144,In_1088);
and U1104 (N_1104,In_573,In_1263);
or U1105 (N_1105,In_443,In_520);
and U1106 (N_1106,In_143,In_1116);
nand U1107 (N_1107,In_311,In_1244);
or U1108 (N_1108,In_591,In_362);
or U1109 (N_1109,In_945,In_619);
and U1110 (N_1110,In_1199,In_1067);
and U1111 (N_1111,In_776,In_968);
and U1112 (N_1112,In_223,In_325);
and U1113 (N_1113,In_1376,In_607);
and U1114 (N_1114,In_989,In_453);
or U1115 (N_1115,In_283,In_124);
and U1116 (N_1116,In_1200,In_407);
nor U1117 (N_1117,In_1105,In_515);
and U1118 (N_1118,In_392,In_271);
nor U1119 (N_1119,In_129,In_1317);
nor U1120 (N_1120,In_1038,In_111);
xor U1121 (N_1121,In_1109,In_1431);
or U1122 (N_1122,In_646,In_1072);
and U1123 (N_1123,In_1084,In_587);
nand U1124 (N_1124,In_1161,In_762);
and U1125 (N_1125,In_41,In_420);
xnor U1126 (N_1126,In_914,In_565);
xor U1127 (N_1127,In_356,In_1279);
and U1128 (N_1128,In_640,In_1197);
or U1129 (N_1129,In_970,In_808);
nor U1130 (N_1130,In_721,In_1441);
or U1131 (N_1131,In_911,In_1413);
nor U1132 (N_1132,In_6,In_848);
or U1133 (N_1133,In_424,In_88);
nor U1134 (N_1134,In_304,In_352);
nor U1135 (N_1135,In_173,In_571);
or U1136 (N_1136,In_1047,In_1212);
or U1137 (N_1137,In_468,In_785);
and U1138 (N_1138,In_1395,In_308);
nand U1139 (N_1139,In_1462,In_1419);
and U1140 (N_1140,In_425,In_1336);
nor U1141 (N_1141,In_1348,In_1006);
or U1142 (N_1142,In_671,In_430);
nand U1143 (N_1143,In_430,In_502);
and U1144 (N_1144,In_353,In_911);
xor U1145 (N_1145,In_1013,In_199);
nor U1146 (N_1146,In_428,In_545);
nor U1147 (N_1147,In_1495,In_1476);
nand U1148 (N_1148,In_943,In_1359);
or U1149 (N_1149,In_830,In_116);
and U1150 (N_1150,In_143,In_1384);
nand U1151 (N_1151,In_539,In_970);
nor U1152 (N_1152,In_661,In_827);
nor U1153 (N_1153,In_34,In_896);
nand U1154 (N_1154,In_1089,In_1380);
nor U1155 (N_1155,In_658,In_169);
nor U1156 (N_1156,In_1003,In_598);
nand U1157 (N_1157,In_934,In_664);
or U1158 (N_1158,In_69,In_1260);
or U1159 (N_1159,In_989,In_1071);
nand U1160 (N_1160,In_1059,In_187);
nor U1161 (N_1161,In_1424,In_180);
nor U1162 (N_1162,In_1166,In_364);
and U1163 (N_1163,In_268,In_231);
and U1164 (N_1164,In_1247,In_122);
nand U1165 (N_1165,In_554,In_587);
nor U1166 (N_1166,In_227,In_91);
nor U1167 (N_1167,In_1343,In_465);
xnor U1168 (N_1168,In_1251,In_1402);
or U1169 (N_1169,In_807,In_241);
and U1170 (N_1170,In_244,In_467);
and U1171 (N_1171,In_658,In_940);
nor U1172 (N_1172,In_1419,In_768);
and U1173 (N_1173,In_472,In_1023);
or U1174 (N_1174,In_207,In_615);
or U1175 (N_1175,In_1167,In_256);
nor U1176 (N_1176,In_1084,In_1402);
nand U1177 (N_1177,In_757,In_1382);
or U1178 (N_1178,In_885,In_911);
and U1179 (N_1179,In_843,In_432);
or U1180 (N_1180,In_673,In_109);
and U1181 (N_1181,In_1188,In_610);
or U1182 (N_1182,In_1489,In_780);
nand U1183 (N_1183,In_11,In_943);
and U1184 (N_1184,In_763,In_713);
nor U1185 (N_1185,In_1323,In_1225);
xnor U1186 (N_1186,In_367,In_1406);
or U1187 (N_1187,In_998,In_1405);
or U1188 (N_1188,In_1497,In_1326);
nor U1189 (N_1189,In_1287,In_1101);
nand U1190 (N_1190,In_763,In_95);
nand U1191 (N_1191,In_288,In_800);
nor U1192 (N_1192,In_1305,In_451);
or U1193 (N_1193,In_101,In_435);
nor U1194 (N_1194,In_1112,In_418);
and U1195 (N_1195,In_1202,In_1357);
nor U1196 (N_1196,In_365,In_799);
or U1197 (N_1197,In_411,In_1489);
nor U1198 (N_1198,In_135,In_581);
nor U1199 (N_1199,In_1101,In_469);
and U1200 (N_1200,In_184,In_364);
and U1201 (N_1201,In_1070,In_1485);
and U1202 (N_1202,In_1115,In_911);
and U1203 (N_1203,In_856,In_821);
or U1204 (N_1204,In_643,In_562);
xor U1205 (N_1205,In_1328,In_428);
or U1206 (N_1206,In_472,In_864);
or U1207 (N_1207,In_301,In_932);
nor U1208 (N_1208,In_877,In_278);
nor U1209 (N_1209,In_649,In_1497);
nor U1210 (N_1210,In_144,In_638);
or U1211 (N_1211,In_168,In_724);
and U1212 (N_1212,In_990,In_574);
and U1213 (N_1213,In_803,In_768);
nand U1214 (N_1214,In_1069,In_806);
nand U1215 (N_1215,In_917,In_678);
or U1216 (N_1216,In_393,In_1259);
and U1217 (N_1217,In_353,In_1391);
nand U1218 (N_1218,In_648,In_548);
and U1219 (N_1219,In_489,In_1155);
or U1220 (N_1220,In_671,In_553);
and U1221 (N_1221,In_698,In_1387);
nor U1222 (N_1222,In_299,In_1266);
nand U1223 (N_1223,In_1483,In_349);
or U1224 (N_1224,In_1146,In_604);
nand U1225 (N_1225,In_1210,In_790);
or U1226 (N_1226,In_122,In_830);
xor U1227 (N_1227,In_1289,In_633);
or U1228 (N_1228,In_788,In_424);
and U1229 (N_1229,In_43,In_318);
and U1230 (N_1230,In_51,In_89);
and U1231 (N_1231,In_205,In_571);
nand U1232 (N_1232,In_883,In_916);
and U1233 (N_1233,In_872,In_835);
nor U1234 (N_1234,In_923,In_134);
xnor U1235 (N_1235,In_27,In_650);
nor U1236 (N_1236,In_1131,In_13);
and U1237 (N_1237,In_735,In_1187);
nand U1238 (N_1238,In_313,In_378);
nor U1239 (N_1239,In_103,In_650);
and U1240 (N_1240,In_384,In_454);
nor U1241 (N_1241,In_566,In_625);
nand U1242 (N_1242,In_1,In_1312);
nor U1243 (N_1243,In_407,In_725);
and U1244 (N_1244,In_893,In_62);
nor U1245 (N_1245,In_279,In_1474);
or U1246 (N_1246,In_1069,In_1416);
and U1247 (N_1247,In_1021,In_814);
and U1248 (N_1248,In_554,In_1325);
and U1249 (N_1249,In_13,In_1150);
nor U1250 (N_1250,In_611,In_524);
and U1251 (N_1251,In_18,In_1258);
nand U1252 (N_1252,In_1047,In_1474);
nor U1253 (N_1253,In_584,In_503);
nand U1254 (N_1254,In_41,In_921);
nor U1255 (N_1255,In_116,In_1138);
or U1256 (N_1256,In_1147,In_354);
or U1257 (N_1257,In_1003,In_35);
or U1258 (N_1258,In_1396,In_580);
nand U1259 (N_1259,In_466,In_1491);
nor U1260 (N_1260,In_343,In_75);
and U1261 (N_1261,In_1404,In_1368);
or U1262 (N_1262,In_1023,In_1254);
or U1263 (N_1263,In_395,In_358);
xor U1264 (N_1264,In_28,In_898);
nand U1265 (N_1265,In_708,In_958);
and U1266 (N_1266,In_1271,In_89);
nand U1267 (N_1267,In_280,In_36);
nand U1268 (N_1268,In_1465,In_897);
or U1269 (N_1269,In_765,In_1206);
nand U1270 (N_1270,In_1257,In_529);
nor U1271 (N_1271,In_711,In_1358);
and U1272 (N_1272,In_245,In_958);
xor U1273 (N_1273,In_1271,In_503);
nand U1274 (N_1274,In_1408,In_1443);
nand U1275 (N_1275,In_645,In_1384);
or U1276 (N_1276,In_239,In_1294);
nor U1277 (N_1277,In_1410,In_1205);
and U1278 (N_1278,In_1000,In_955);
and U1279 (N_1279,In_702,In_951);
or U1280 (N_1280,In_920,In_211);
nand U1281 (N_1281,In_991,In_40);
nand U1282 (N_1282,In_917,In_769);
and U1283 (N_1283,In_1060,In_500);
and U1284 (N_1284,In_1304,In_702);
nand U1285 (N_1285,In_19,In_197);
nor U1286 (N_1286,In_1294,In_289);
or U1287 (N_1287,In_571,In_29);
nor U1288 (N_1288,In_630,In_919);
nor U1289 (N_1289,In_1036,In_282);
nor U1290 (N_1290,In_1404,In_682);
nor U1291 (N_1291,In_1269,In_1209);
nor U1292 (N_1292,In_1467,In_1434);
nand U1293 (N_1293,In_1405,In_1315);
or U1294 (N_1294,In_192,In_438);
or U1295 (N_1295,In_990,In_854);
xor U1296 (N_1296,In_708,In_1125);
nand U1297 (N_1297,In_819,In_841);
and U1298 (N_1298,In_234,In_169);
nor U1299 (N_1299,In_992,In_923);
nor U1300 (N_1300,In_15,In_373);
nand U1301 (N_1301,In_606,In_786);
nor U1302 (N_1302,In_1326,In_1263);
nand U1303 (N_1303,In_823,In_216);
or U1304 (N_1304,In_450,In_808);
nand U1305 (N_1305,In_591,In_961);
or U1306 (N_1306,In_1072,In_496);
xor U1307 (N_1307,In_1206,In_1431);
nor U1308 (N_1308,In_523,In_147);
nor U1309 (N_1309,In_1117,In_883);
xor U1310 (N_1310,In_1000,In_18);
or U1311 (N_1311,In_570,In_469);
nor U1312 (N_1312,In_370,In_241);
and U1313 (N_1313,In_207,In_861);
or U1314 (N_1314,In_664,In_866);
nor U1315 (N_1315,In_1271,In_857);
nand U1316 (N_1316,In_541,In_756);
and U1317 (N_1317,In_229,In_1308);
or U1318 (N_1318,In_825,In_1169);
or U1319 (N_1319,In_178,In_964);
or U1320 (N_1320,In_589,In_390);
and U1321 (N_1321,In_156,In_584);
and U1322 (N_1322,In_1150,In_831);
xnor U1323 (N_1323,In_1283,In_1408);
and U1324 (N_1324,In_386,In_1411);
nand U1325 (N_1325,In_120,In_931);
nor U1326 (N_1326,In_857,In_1359);
nor U1327 (N_1327,In_593,In_624);
nand U1328 (N_1328,In_100,In_525);
nor U1329 (N_1329,In_668,In_962);
nand U1330 (N_1330,In_557,In_162);
nor U1331 (N_1331,In_96,In_737);
and U1332 (N_1332,In_193,In_989);
nand U1333 (N_1333,In_1306,In_1139);
xnor U1334 (N_1334,In_1242,In_841);
or U1335 (N_1335,In_196,In_616);
xor U1336 (N_1336,In_1007,In_533);
and U1337 (N_1337,In_1352,In_490);
and U1338 (N_1338,In_551,In_806);
nand U1339 (N_1339,In_1301,In_706);
and U1340 (N_1340,In_10,In_405);
nand U1341 (N_1341,In_184,In_292);
and U1342 (N_1342,In_307,In_240);
and U1343 (N_1343,In_606,In_495);
and U1344 (N_1344,In_644,In_1086);
nor U1345 (N_1345,In_840,In_681);
and U1346 (N_1346,In_608,In_264);
nor U1347 (N_1347,In_574,In_1427);
nand U1348 (N_1348,In_1316,In_293);
and U1349 (N_1349,In_919,In_1234);
nand U1350 (N_1350,In_858,In_1488);
nor U1351 (N_1351,In_1363,In_1181);
nor U1352 (N_1352,In_240,In_120);
xnor U1353 (N_1353,In_1181,In_1293);
or U1354 (N_1354,In_1310,In_502);
or U1355 (N_1355,In_1329,In_834);
or U1356 (N_1356,In_574,In_229);
xnor U1357 (N_1357,In_1009,In_988);
xnor U1358 (N_1358,In_228,In_355);
nand U1359 (N_1359,In_171,In_1357);
nor U1360 (N_1360,In_421,In_842);
nand U1361 (N_1361,In_1156,In_1373);
and U1362 (N_1362,In_1251,In_678);
or U1363 (N_1363,In_1423,In_1035);
and U1364 (N_1364,In_157,In_647);
and U1365 (N_1365,In_929,In_1181);
and U1366 (N_1366,In_810,In_722);
nand U1367 (N_1367,In_899,In_686);
nor U1368 (N_1368,In_662,In_1131);
and U1369 (N_1369,In_1277,In_362);
nor U1370 (N_1370,In_164,In_1493);
and U1371 (N_1371,In_1186,In_629);
nand U1372 (N_1372,In_954,In_927);
nor U1373 (N_1373,In_346,In_84);
and U1374 (N_1374,In_247,In_192);
nor U1375 (N_1375,In_1017,In_1057);
or U1376 (N_1376,In_1058,In_522);
nor U1377 (N_1377,In_1158,In_238);
or U1378 (N_1378,In_434,In_1441);
nor U1379 (N_1379,In_720,In_790);
or U1380 (N_1380,In_802,In_93);
xor U1381 (N_1381,In_108,In_632);
nand U1382 (N_1382,In_1261,In_1089);
xor U1383 (N_1383,In_480,In_357);
nor U1384 (N_1384,In_830,In_1435);
nor U1385 (N_1385,In_650,In_724);
and U1386 (N_1386,In_510,In_323);
and U1387 (N_1387,In_63,In_357);
nor U1388 (N_1388,In_1093,In_194);
nand U1389 (N_1389,In_1332,In_663);
nand U1390 (N_1390,In_457,In_283);
nor U1391 (N_1391,In_276,In_773);
or U1392 (N_1392,In_835,In_192);
xnor U1393 (N_1393,In_1037,In_1384);
nand U1394 (N_1394,In_1255,In_1200);
nor U1395 (N_1395,In_874,In_1026);
nor U1396 (N_1396,In_812,In_289);
nand U1397 (N_1397,In_925,In_861);
and U1398 (N_1398,In_40,In_1261);
and U1399 (N_1399,In_109,In_1461);
or U1400 (N_1400,In_607,In_1441);
xor U1401 (N_1401,In_1221,In_698);
xnor U1402 (N_1402,In_466,In_243);
nor U1403 (N_1403,In_1303,In_175);
and U1404 (N_1404,In_1055,In_1410);
nand U1405 (N_1405,In_936,In_444);
nand U1406 (N_1406,In_145,In_383);
or U1407 (N_1407,In_1150,In_305);
nand U1408 (N_1408,In_127,In_1113);
and U1409 (N_1409,In_425,In_512);
nand U1410 (N_1410,In_700,In_1174);
or U1411 (N_1411,In_191,In_226);
xnor U1412 (N_1412,In_925,In_689);
or U1413 (N_1413,In_1039,In_969);
or U1414 (N_1414,In_949,In_415);
nand U1415 (N_1415,In_194,In_1433);
nor U1416 (N_1416,In_1165,In_1071);
and U1417 (N_1417,In_1301,In_769);
nor U1418 (N_1418,In_506,In_278);
nand U1419 (N_1419,In_889,In_1070);
nor U1420 (N_1420,In_591,In_235);
and U1421 (N_1421,In_889,In_847);
and U1422 (N_1422,In_980,In_1349);
xnor U1423 (N_1423,In_527,In_967);
or U1424 (N_1424,In_99,In_1299);
or U1425 (N_1425,In_602,In_1472);
and U1426 (N_1426,In_313,In_1470);
or U1427 (N_1427,In_699,In_814);
xnor U1428 (N_1428,In_244,In_419);
nor U1429 (N_1429,In_676,In_529);
or U1430 (N_1430,In_579,In_527);
xor U1431 (N_1431,In_1203,In_379);
and U1432 (N_1432,In_1265,In_713);
and U1433 (N_1433,In_67,In_302);
and U1434 (N_1434,In_1073,In_1474);
and U1435 (N_1435,In_901,In_1);
nor U1436 (N_1436,In_157,In_1232);
nor U1437 (N_1437,In_283,In_705);
nor U1438 (N_1438,In_235,In_539);
or U1439 (N_1439,In_112,In_201);
xnor U1440 (N_1440,In_998,In_660);
nand U1441 (N_1441,In_1488,In_135);
nor U1442 (N_1442,In_1405,In_914);
nor U1443 (N_1443,In_556,In_1227);
or U1444 (N_1444,In_186,In_1315);
nand U1445 (N_1445,In_95,In_293);
and U1446 (N_1446,In_232,In_1481);
nor U1447 (N_1447,In_1459,In_802);
and U1448 (N_1448,In_605,In_1445);
and U1449 (N_1449,In_262,In_172);
nand U1450 (N_1450,In_290,In_2);
nand U1451 (N_1451,In_354,In_942);
nor U1452 (N_1452,In_133,In_1148);
nor U1453 (N_1453,In_1115,In_653);
nand U1454 (N_1454,In_1456,In_965);
xnor U1455 (N_1455,In_675,In_91);
or U1456 (N_1456,In_378,In_288);
and U1457 (N_1457,In_567,In_1363);
nor U1458 (N_1458,In_952,In_1118);
nor U1459 (N_1459,In_704,In_247);
and U1460 (N_1460,In_911,In_1312);
nand U1461 (N_1461,In_567,In_419);
nand U1462 (N_1462,In_480,In_1392);
and U1463 (N_1463,In_1071,In_694);
and U1464 (N_1464,In_446,In_1220);
nor U1465 (N_1465,In_94,In_391);
nand U1466 (N_1466,In_1036,In_804);
nand U1467 (N_1467,In_1480,In_681);
and U1468 (N_1468,In_130,In_1055);
nor U1469 (N_1469,In_6,In_408);
xor U1470 (N_1470,In_235,In_841);
and U1471 (N_1471,In_1182,In_344);
and U1472 (N_1472,In_763,In_416);
nor U1473 (N_1473,In_547,In_351);
and U1474 (N_1474,In_959,In_834);
or U1475 (N_1475,In_646,In_1120);
and U1476 (N_1476,In_652,In_877);
xor U1477 (N_1477,In_428,In_135);
and U1478 (N_1478,In_475,In_436);
or U1479 (N_1479,In_112,In_1131);
or U1480 (N_1480,In_283,In_1289);
nor U1481 (N_1481,In_248,In_872);
or U1482 (N_1482,In_718,In_549);
and U1483 (N_1483,In_1182,In_1386);
xor U1484 (N_1484,In_1286,In_1350);
nor U1485 (N_1485,In_900,In_1255);
nor U1486 (N_1486,In_134,In_808);
or U1487 (N_1487,In_1179,In_8);
or U1488 (N_1488,In_137,In_427);
and U1489 (N_1489,In_60,In_91);
or U1490 (N_1490,In_37,In_1008);
xnor U1491 (N_1491,In_55,In_1099);
and U1492 (N_1492,In_528,In_603);
and U1493 (N_1493,In_1347,In_1381);
nand U1494 (N_1494,In_854,In_1314);
xnor U1495 (N_1495,In_1353,In_766);
nor U1496 (N_1496,In_974,In_1397);
nand U1497 (N_1497,In_801,In_940);
nand U1498 (N_1498,In_1008,In_85);
nand U1499 (N_1499,In_44,In_800);
nor U1500 (N_1500,In_1369,In_1471);
or U1501 (N_1501,In_1281,In_1470);
and U1502 (N_1502,In_875,In_394);
nor U1503 (N_1503,In_302,In_1361);
xor U1504 (N_1504,In_488,In_1468);
xnor U1505 (N_1505,In_1362,In_260);
or U1506 (N_1506,In_532,In_1064);
nand U1507 (N_1507,In_662,In_894);
nor U1508 (N_1508,In_699,In_1096);
and U1509 (N_1509,In_537,In_104);
nand U1510 (N_1510,In_1001,In_1200);
nand U1511 (N_1511,In_557,In_1240);
xnor U1512 (N_1512,In_823,In_715);
nand U1513 (N_1513,In_1346,In_599);
and U1514 (N_1514,In_931,In_1100);
xnor U1515 (N_1515,In_1259,In_1308);
nor U1516 (N_1516,In_1223,In_144);
or U1517 (N_1517,In_343,In_189);
nand U1518 (N_1518,In_483,In_1435);
nor U1519 (N_1519,In_989,In_347);
nand U1520 (N_1520,In_457,In_901);
and U1521 (N_1521,In_242,In_675);
nor U1522 (N_1522,In_626,In_907);
nor U1523 (N_1523,In_461,In_415);
nand U1524 (N_1524,In_452,In_1303);
and U1525 (N_1525,In_1264,In_386);
nand U1526 (N_1526,In_1151,In_240);
nand U1527 (N_1527,In_33,In_631);
xor U1528 (N_1528,In_88,In_423);
or U1529 (N_1529,In_19,In_1240);
xnor U1530 (N_1530,In_1203,In_1242);
nor U1531 (N_1531,In_142,In_776);
nand U1532 (N_1532,In_462,In_1448);
nand U1533 (N_1533,In_414,In_758);
and U1534 (N_1534,In_1216,In_1084);
nand U1535 (N_1535,In_1372,In_921);
nor U1536 (N_1536,In_512,In_1068);
or U1537 (N_1537,In_1177,In_1331);
or U1538 (N_1538,In_525,In_366);
and U1539 (N_1539,In_891,In_476);
nand U1540 (N_1540,In_478,In_760);
or U1541 (N_1541,In_294,In_1113);
nand U1542 (N_1542,In_9,In_1413);
and U1543 (N_1543,In_1301,In_837);
and U1544 (N_1544,In_969,In_1230);
and U1545 (N_1545,In_1405,In_343);
nand U1546 (N_1546,In_1025,In_1170);
and U1547 (N_1547,In_763,In_787);
and U1548 (N_1548,In_822,In_1435);
nor U1549 (N_1549,In_1405,In_53);
nor U1550 (N_1550,In_750,In_669);
and U1551 (N_1551,In_1323,In_1001);
nor U1552 (N_1552,In_1087,In_1448);
nand U1553 (N_1553,In_1082,In_184);
xnor U1554 (N_1554,In_803,In_1207);
nand U1555 (N_1555,In_256,In_568);
xor U1556 (N_1556,In_1073,In_654);
or U1557 (N_1557,In_232,In_900);
or U1558 (N_1558,In_1314,In_634);
nand U1559 (N_1559,In_415,In_387);
nand U1560 (N_1560,In_240,In_338);
or U1561 (N_1561,In_587,In_1133);
and U1562 (N_1562,In_1095,In_136);
nor U1563 (N_1563,In_844,In_700);
or U1564 (N_1564,In_1097,In_1077);
and U1565 (N_1565,In_951,In_836);
and U1566 (N_1566,In_251,In_711);
nand U1567 (N_1567,In_208,In_875);
xor U1568 (N_1568,In_1208,In_678);
or U1569 (N_1569,In_202,In_531);
and U1570 (N_1570,In_1294,In_516);
nand U1571 (N_1571,In_830,In_516);
or U1572 (N_1572,In_855,In_787);
and U1573 (N_1573,In_737,In_1443);
and U1574 (N_1574,In_282,In_1416);
and U1575 (N_1575,In_559,In_323);
nor U1576 (N_1576,In_848,In_106);
nor U1577 (N_1577,In_670,In_96);
and U1578 (N_1578,In_1125,In_176);
nand U1579 (N_1579,In_5,In_24);
and U1580 (N_1580,In_696,In_317);
or U1581 (N_1581,In_295,In_674);
nand U1582 (N_1582,In_28,In_225);
nand U1583 (N_1583,In_441,In_39);
nor U1584 (N_1584,In_1029,In_690);
nand U1585 (N_1585,In_849,In_644);
nor U1586 (N_1586,In_1436,In_837);
nor U1587 (N_1587,In_150,In_1122);
nand U1588 (N_1588,In_694,In_963);
and U1589 (N_1589,In_368,In_1175);
nand U1590 (N_1590,In_1364,In_116);
and U1591 (N_1591,In_597,In_1165);
nor U1592 (N_1592,In_608,In_804);
and U1593 (N_1593,In_1132,In_132);
nand U1594 (N_1594,In_658,In_390);
and U1595 (N_1595,In_676,In_642);
and U1596 (N_1596,In_837,In_570);
or U1597 (N_1597,In_1172,In_1395);
nand U1598 (N_1598,In_266,In_1255);
nand U1599 (N_1599,In_1315,In_541);
and U1600 (N_1600,In_657,In_677);
nand U1601 (N_1601,In_884,In_613);
nand U1602 (N_1602,In_706,In_1224);
or U1603 (N_1603,In_1338,In_228);
nor U1604 (N_1604,In_1184,In_1497);
and U1605 (N_1605,In_1447,In_535);
and U1606 (N_1606,In_393,In_344);
or U1607 (N_1607,In_863,In_888);
or U1608 (N_1608,In_277,In_879);
nor U1609 (N_1609,In_65,In_995);
nor U1610 (N_1610,In_901,In_1110);
nand U1611 (N_1611,In_305,In_1178);
nand U1612 (N_1612,In_968,In_929);
xnor U1613 (N_1613,In_795,In_457);
or U1614 (N_1614,In_1384,In_1280);
nor U1615 (N_1615,In_444,In_1007);
xnor U1616 (N_1616,In_1212,In_704);
nor U1617 (N_1617,In_732,In_1459);
or U1618 (N_1618,In_779,In_505);
nand U1619 (N_1619,In_808,In_1457);
nand U1620 (N_1620,In_17,In_159);
nor U1621 (N_1621,In_1132,In_512);
xor U1622 (N_1622,In_1326,In_1020);
and U1623 (N_1623,In_323,In_65);
xor U1624 (N_1624,In_755,In_945);
nand U1625 (N_1625,In_204,In_167);
nand U1626 (N_1626,In_193,In_796);
or U1627 (N_1627,In_1082,In_1191);
or U1628 (N_1628,In_496,In_214);
and U1629 (N_1629,In_1317,In_50);
and U1630 (N_1630,In_1260,In_790);
and U1631 (N_1631,In_1119,In_160);
nand U1632 (N_1632,In_959,In_1221);
or U1633 (N_1633,In_858,In_1214);
and U1634 (N_1634,In_999,In_60);
or U1635 (N_1635,In_639,In_1470);
and U1636 (N_1636,In_1059,In_1066);
and U1637 (N_1637,In_136,In_1225);
nor U1638 (N_1638,In_1,In_304);
nand U1639 (N_1639,In_1173,In_723);
or U1640 (N_1640,In_830,In_52);
nor U1641 (N_1641,In_180,In_519);
nor U1642 (N_1642,In_417,In_446);
nor U1643 (N_1643,In_1018,In_730);
nand U1644 (N_1644,In_684,In_1337);
nand U1645 (N_1645,In_86,In_773);
nand U1646 (N_1646,In_507,In_435);
nand U1647 (N_1647,In_547,In_1366);
or U1648 (N_1648,In_970,In_525);
or U1649 (N_1649,In_1240,In_1363);
nor U1650 (N_1650,In_599,In_27);
or U1651 (N_1651,In_231,In_940);
nand U1652 (N_1652,In_858,In_957);
or U1653 (N_1653,In_494,In_290);
or U1654 (N_1654,In_140,In_359);
or U1655 (N_1655,In_1314,In_1103);
or U1656 (N_1656,In_40,In_1428);
or U1657 (N_1657,In_547,In_882);
and U1658 (N_1658,In_1140,In_685);
and U1659 (N_1659,In_212,In_873);
xor U1660 (N_1660,In_890,In_112);
nor U1661 (N_1661,In_436,In_121);
xnor U1662 (N_1662,In_1343,In_165);
nand U1663 (N_1663,In_701,In_328);
xor U1664 (N_1664,In_478,In_494);
and U1665 (N_1665,In_1496,In_262);
xor U1666 (N_1666,In_603,In_1193);
nor U1667 (N_1667,In_930,In_1439);
or U1668 (N_1668,In_953,In_1202);
and U1669 (N_1669,In_1285,In_945);
nand U1670 (N_1670,In_763,In_996);
nand U1671 (N_1671,In_392,In_582);
or U1672 (N_1672,In_937,In_1085);
or U1673 (N_1673,In_1350,In_492);
and U1674 (N_1674,In_1047,In_895);
or U1675 (N_1675,In_1130,In_299);
or U1676 (N_1676,In_241,In_1104);
xor U1677 (N_1677,In_243,In_570);
nand U1678 (N_1678,In_1303,In_1166);
nand U1679 (N_1679,In_103,In_1164);
nand U1680 (N_1680,In_881,In_962);
or U1681 (N_1681,In_1469,In_1357);
or U1682 (N_1682,In_354,In_570);
nand U1683 (N_1683,In_645,In_819);
nor U1684 (N_1684,In_883,In_302);
and U1685 (N_1685,In_215,In_612);
nand U1686 (N_1686,In_1396,In_1357);
nor U1687 (N_1687,In_560,In_524);
or U1688 (N_1688,In_858,In_232);
and U1689 (N_1689,In_1447,In_418);
nor U1690 (N_1690,In_927,In_1208);
nor U1691 (N_1691,In_675,In_769);
and U1692 (N_1692,In_368,In_896);
or U1693 (N_1693,In_1246,In_852);
xnor U1694 (N_1694,In_772,In_902);
nand U1695 (N_1695,In_490,In_868);
nand U1696 (N_1696,In_28,In_808);
and U1697 (N_1697,In_1049,In_996);
xor U1698 (N_1698,In_935,In_377);
or U1699 (N_1699,In_657,In_1297);
nor U1700 (N_1700,In_707,In_1129);
or U1701 (N_1701,In_1213,In_1237);
and U1702 (N_1702,In_1435,In_1144);
or U1703 (N_1703,In_859,In_354);
nand U1704 (N_1704,In_189,In_219);
or U1705 (N_1705,In_113,In_1398);
and U1706 (N_1706,In_938,In_196);
or U1707 (N_1707,In_477,In_1347);
or U1708 (N_1708,In_844,In_488);
nor U1709 (N_1709,In_1060,In_1334);
or U1710 (N_1710,In_1420,In_1378);
xnor U1711 (N_1711,In_898,In_1029);
nor U1712 (N_1712,In_198,In_220);
and U1713 (N_1713,In_1095,In_1177);
nand U1714 (N_1714,In_643,In_230);
or U1715 (N_1715,In_1306,In_1454);
and U1716 (N_1716,In_868,In_533);
or U1717 (N_1717,In_1459,In_327);
nor U1718 (N_1718,In_368,In_950);
nor U1719 (N_1719,In_1479,In_723);
nand U1720 (N_1720,In_96,In_198);
nor U1721 (N_1721,In_84,In_92);
nand U1722 (N_1722,In_1109,In_70);
or U1723 (N_1723,In_88,In_235);
nand U1724 (N_1724,In_1336,In_857);
nand U1725 (N_1725,In_1375,In_371);
or U1726 (N_1726,In_950,In_1006);
and U1727 (N_1727,In_257,In_976);
nor U1728 (N_1728,In_673,In_203);
and U1729 (N_1729,In_39,In_262);
and U1730 (N_1730,In_227,In_1108);
nand U1731 (N_1731,In_159,In_1154);
nand U1732 (N_1732,In_1219,In_1175);
nand U1733 (N_1733,In_301,In_227);
and U1734 (N_1734,In_768,In_1405);
nand U1735 (N_1735,In_1219,In_517);
nor U1736 (N_1736,In_1104,In_731);
nand U1737 (N_1737,In_1432,In_188);
nand U1738 (N_1738,In_757,In_1215);
xor U1739 (N_1739,In_687,In_411);
nor U1740 (N_1740,In_121,In_885);
and U1741 (N_1741,In_301,In_356);
xor U1742 (N_1742,In_23,In_297);
or U1743 (N_1743,In_1154,In_221);
and U1744 (N_1744,In_935,In_232);
xnor U1745 (N_1745,In_19,In_66);
and U1746 (N_1746,In_1139,In_1182);
nand U1747 (N_1747,In_826,In_971);
or U1748 (N_1748,In_726,In_1137);
nor U1749 (N_1749,In_585,In_725);
nand U1750 (N_1750,In_843,In_827);
nand U1751 (N_1751,In_1187,In_989);
xor U1752 (N_1752,In_559,In_416);
and U1753 (N_1753,In_929,In_148);
nor U1754 (N_1754,In_911,In_1151);
or U1755 (N_1755,In_569,In_1046);
nand U1756 (N_1756,In_1074,In_522);
and U1757 (N_1757,In_239,In_1053);
or U1758 (N_1758,In_765,In_1496);
or U1759 (N_1759,In_773,In_1461);
and U1760 (N_1760,In_629,In_290);
nand U1761 (N_1761,In_138,In_1138);
or U1762 (N_1762,In_530,In_1313);
xnor U1763 (N_1763,In_209,In_485);
nand U1764 (N_1764,In_18,In_211);
nand U1765 (N_1765,In_180,In_1360);
and U1766 (N_1766,In_277,In_1080);
nor U1767 (N_1767,In_318,In_461);
nand U1768 (N_1768,In_1419,In_1055);
nand U1769 (N_1769,In_191,In_1445);
or U1770 (N_1770,In_971,In_1098);
or U1771 (N_1771,In_1162,In_921);
and U1772 (N_1772,In_388,In_1317);
nor U1773 (N_1773,In_631,In_381);
nor U1774 (N_1774,In_1173,In_1230);
and U1775 (N_1775,In_1463,In_174);
xor U1776 (N_1776,In_1196,In_301);
nand U1777 (N_1777,In_779,In_127);
xnor U1778 (N_1778,In_57,In_1391);
xor U1779 (N_1779,In_536,In_1254);
or U1780 (N_1780,In_344,In_1142);
or U1781 (N_1781,In_1057,In_750);
nor U1782 (N_1782,In_509,In_1454);
and U1783 (N_1783,In_566,In_1276);
or U1784 (N_1784,In_733,In_1486);
or U1785 (N_1785,In_919,In_1337);
nand U1786 (N_1786,In_1040,In_653);
nor U1787 (N_1787,In_387,In_1018);
nand U1788 (N_1788,In_1155,In_61);
and U1789 (N_1789,In_78,In_1477);
and U1790 (N_1790,In_1044,In_948);
and U1791 (N_1791,In_1243,In_1432);
or U1792 (N_1792,In_1326,In_1289);
or U1793 (N_1793,In_95,In_234);
xnor U1794 (N_1794,In_22,In_654);
and U1795 (N_1795,In_967,In_1352);
or U1796 (N_1796,In_1223,In_671);
nor U1797 (N_1797,In_126,In_748);
nor U1798 (N_1798,In_13,In_612);
nand U1799 (N_1799,In_1216,In_480);
nand U1800 (N_1800,In_1297,In_1481);
nand U1801 (N_1801,In_1111,In_1361);
and U1802 (N_1802,In_931,In_412);
or U1803 (N_1803,In_1036,In_1142);
or U1804 (N_1804,In_1440,In_374);
nor U1805 (N_1805,In_328,In_877);
and U1806 (N_1806,In_424,In_372);
nand U1807 (N_1807,In_1081,In_1018);
and U1808 (N_1808,In_970,In_67);
or U1809 (N_1809,In_1395,In_1265);
and U1810 (N_1810,In_673,In_1320);
nand U1811 (N_1811,In_1159,In_7);
nand U1812 (N_1812,In_1388,In_549);
xor U1813 (N_1813,In_32,In_1013);
and U1814 (N_1814,In_555,In_725);
nand U1815 (N_1815,In_1004,In_662);
nand U1816 (N_1816,In_482,In_3);
nor U1817 (N_1817,In_459,In_862);
and U1818 (N_1818,In_310,In_1088);
nor U1819 (N_1819,In_513,In_826);
and U1820 (N_1820,In_387,In_1211);
nor U1821 (N_1821,In_656,In_1193);
and U1822 (N_1822,In_601,In_458);
and U1823 (N_1823,In_537,In_1485);
nor U1824 (N_1824,In_171,In_1214);
or U1825 (N_1825,In_6,In_885);
xor U1826 (N_1826,In_721,In_1132);
or U1827 (N_1827,In_17,In_1368);
or U1828 (N_1828,In_484,In_1119);
nor U1829 (N_1829,In_1241,In_1264);
nand U1830 (N_1830,In_401,In_11);
xnor U1831 (N_1831,In_605,In_1217);
nor U1832 (N_1832,In_674,In_682);
and U1833 (N_1833,In_469,In_1410);
nand U1834 (N_1834,In_713,In_813);
nor U1835 (N_1835,In_434,In_578);
nor U1836 (N_1836,In_539,In_297);
nand U1837 (N_1837,In_668,In_48);
or U1838 (N_1838,In_328,In_1386);
or U1839 (N_1839,In_453,In_1152);
nor U1840 (N_1840,In_1088,In_1147);
and U1841 (N_1841,In_1126,In_1318);
nand U1842 (N_1842,In_1427,In_1380);
nor U1843 (N_1843,In_1172,In_1239);
nand U1844 (N_1844,In_150,In_1106);
or U1845 (N_1845,In_747,In_29);
nor U1846 (N_1846,In_872,In_1068);
or U1847 (N_1847,In_1304,In_810);
nand U1848 (N_1848,In_108,In_501);
and U1849 (N_1849,In_102,In_654);
or U1850 (N_1850,In_1072,In_1046);
or U1851 (N_1851,In_384,In_504);
and U1852 (N_1852,In_1267,In_1072);
nor U1853 (N_1853,In_478,In_170);
nand U1854 (N_1854,In_243,In_971);
and U1855 (N_1855,In_733,In_1379);
xor U1856 (N_1856,In_214,In_1262);
nor U1857 (N_1857,In_903,In_1067);
nor U1858 (N_1858,In_1180,In_1261);
or U1859 (N_1859,In_1171,In_756);
nor U1860 (N_1860,In_779,In_53);
nor U1861 (N_1861,In_586,In_919);
nand U1862 (N_1862,In_725,In_96);
nor U1863 (N_1863,In_1040,In_964);
and U1864 (N_1864,In_927,In_518);
and U1865 (N_1865,In_1284,In_1297);
nand U1866 (N_1866,In_764,In_1268);
nand U1867 (N_1867,In_1046,In_1134);
nor U1868 (N_1868,In_1018,In_153);
nand U1869 (N_1869,In_1440,In_959);
or U1870 (N_1870,In_298,In_559);
nand U1871 (N_1871,In_706,In_365);
xnor U1872 (N_1872,In_1148,In_802);
or U1873 (N_1873,In_353,In_599);
nand U1874 (N_1874,In_959,In_1495);
or U1875 (N_1875,In_1387,In_269);
nor U1876 (N_1876,In_411,In_138);
and U1877 (N_1877,In_821,In_83);
or U1878 (N_1878,In_1004,In_1099);
nor U1879 (N_1879,In_1412,In_270);
xor U1880 (N_1880,In_699,In_615);
and U1881 (N_1881,In_900,In_550);
nor U1882 (N_1882,In_913,In_520);
or U1883 (N_1883,In_651,In_57);
and U1884 (N_1884,In_258,In_689);
xor U1885 (N_1885,In_538,In_217);
nor U1886 (N_1886,In_81,In_706);
or U1887 (N_1887,In_798,In_636);
and U1888 (N_1888,In_1368,In_1093);
nand U1889 (N_1889,In_672,In_1196);
and U1890 (N_1890,In_382,In_378);
and U1891 (N_1891,In_259,In_1278);
xor U1892 (N_1892,In_1296,In_143);
nand U1893 (N_1893,In_167,In_1079);
or U1894 (N_1894,In_290,In_246);
and U1895 (N_1895,In_442,In_240);
or U1896 (N_1896,In_1405,In_702);
or U1897 (N_1897,In_1131,In_464);
or U1898 (N_1898,In_643,In_182);
nor U1899 (N_1899,In_51,In_1385);
xor U1900 (N_1900,In_1111,In_526);
or U1901 (N_1901,In_1494,In_670);
nor U1902 (N_1902,In_1462,In_558);
or U1903 (N_1903,In_1299,In_553);
nand U1904 (N_1904,In_160,In_859);
and U1905 (N_1905,In_733,In_1037);
xnor U1906 (N_1906,In_284,In_156);
xnor U1907 (N_1907,In_732,In_50);
nand U1908 (N_1908,In_1157,In_717);
or U1909 (N_1909,In_861,In_435);
nor U1910 (N_1910,In_261,In_477);
or U1911 (N_1911,In_1483,In_1242);
and U1912 (N_1912,In_1320,In_1477);
nor U1913 (N_1913,In_803,In_1100);
and U1914 (N_1914,In_1465,In_143);
nand U1915 (N_1915,In_852,In_836);
or U1916 (N_1916,In_1201,In_456);
nor U1917 (N_1917,In_15,In_26);
or U1918 (N_1918,In_1308,In_342);
and U1919 (N_1919,In_1041,In_1114);
or U1920 (N_1920,In_603,In_1408);
nor U1921 (N_1921,In_422,In_447);
or U1922 (N_1922,In_977,In_602);
and U1923 (N_1923,In_381,In_915);
and U1924 (N_1924,In_929,In_481);
xnor U1925 (N_1925,In_52,In_38);
and U1926 (N_1926,In_1132,In_112);
xor U1927 (N_1927,In_1493,In_824);
nand U1928 (N_1928,In_1057,In_19);
nor U1929 (N_1929,In_53,In_1003);
nor U1930 (N_1930,In_502,In_1408);
nor U1931 (N_1931,In_658,In_1308);
xor U1932 (N_1932,In_1461,In_294);
nor U1933 (N_1933,In_1051,In_1487);
or U1934 (N_1934,In_1327,In_1453);
xor U1935 (N_1935,In_667,In_103);
nor U1936 (N_1936,In_1181,In_1281);
and U1937 (N_1937,In_654,In_428);
or U1938 (N_1938,In_1281,In_289);
nor U1939 (N_1939,In_203,In_648);
nand U1940 (N_1940,In_1127,In_1039);
nand U1941 (N_1941,In_1169,In_329);
nor U1942 (N_1942,In_1310,In_898);
and U1943 (N_1943,In_591,In_1226);
nand U1944 (N_1944,In_526,In_409);
or U1945 (N_1945,In_150,In_825);
nand U1946 (N_1946,In_893,In_408);
or U1947 (N_1947,In_793,In_891);
or U1948 (N_1948,In_100,In_222);
nor U1949 (N_1949,In_1202,In_1407);
or U1950 (N_1950,In_754,In_238);
nor U1951 (N_1951,In_28,In_99);
xor U1952 (N_1952,In_1475,In_782);
nand U1953 (N_1953,In_912,In_738);
nor U1954 (N_1954,In_380,In_801);
or U1955 (N_1955,In_898,In_236);
nand U1956 (N_1956,In_1042,In_1122);
and U1957 (N_1957,In_453,In_500);
and U1958 (N_1958,In_1333,In_821);
nor U1959 (N_1959,In_621,In_1406);
and U1960 (N_1960,In_143,In_1469);
or U1961 (N_1961,In_124,In_428);
nor U1962 (N_1962,In_206,In_90);
nand U1963 (N_1963,In_118,In_404);
nor U1964 (N_1964,In_1202,In_399);
nand U1965 (N_1965,In_157,In_266);
or U1966 (N_1966,In_267,In_278);
or U1967 (N_1967,In_1364,In_594);
nor U1968 (N_1968,In_903,In_655);
nand U1969 (N_1969,In_426,In_863);
or U1970 (N_1970,In_520,In_181);
and U1971 (N_1971,In_1443,In_437);
nor U1972 (N_1972,In_1174,In_592);
or U1973 (N_1973,In_1307,In_1301);
nor U1974 (N_1974,In_935,In_879);
and U1975 (N_1975,In_601,In_646);
and U1976 (N_1976,In_869,In_468);
nor U1977 (N_1977,In_1008,In_1231);
and U1978 (N_1978,In_457,In_1468);
nor U1979 (N_1979,In_64,In_753);
nand U1980 (N_1980,In_1374,In_885);
nor U1981 (N_1981,In_411,In_521);
and U1982 (N_1982,In_721,In_1084);
and U1983 (N_1983,In_155,In_1346);
nand U1984 (N_1984,In_393,In_252);
nor U1985 (N_1985,In_680,In_47);
or U1986 (N_1986,In_654,In_762);
and U1987 (N_1987,In_855,In_525);
or U1988 (N_1988,In_883,In_1059);
nand U1989 (N_1989,In_1430,In_356);
xnor U1990 (N_1990,In_313,In_32);
nor U1991 (N_1991,In_1299,In_157);
nand U1992 (N_1992,In_1015,In_326);
xnor U1993 (N_1993,In_85,In_598);
xor U1994 (N_1994,In_20,In_763);
xor U1995 (N_1995,In_95,In_1007);
and U1996 (N_1996,In_813,In_54);
or U1997 (N_1997,In_1236,In_298);
nand U1998 (N_1998,In_577,In_795);
and U1999 (N_1999,In_730,In_498);
or U2000 (N_2000,In_204,In_554);
and U2001 (N_2001,In_203,In_793);
and U2002 (N_2002,In_333,In_63);
and U2003 (N_2003,In_1417,In_1257);
or U2004 (N_2004,In_1357,In_977);
nor U2005 (N_2005,In_266,In_904);
and U2006 (N_2006,In_1332,In_234);
and U2007 (N_2007,In_1467,In_1052);
or U2008 (N_2008,In_1235,In_1068);
or U2009 (N_2009,In_1044,In_787);
or U2010 (N_2010,In_1278,In_895);
nand U2011 (N_2011,In_259,In_403);
xor U2012 (N_2012,In_1260,In_178);
nor U2013 (N_2013,In_949,In_1445);
or U2014 (N_2014,In_737,In_1113);
or U2015 (N_2015,In_1432,In_573);
nor U2016 (N_2016,In_195,In_796);
nand U2017 (N_2017,In_1074,In_667);
nor U2018 (N_2018,In_1386,In_1333);
or U2019 (N_2019,In_1357,In_609);
or U2020 (N_2020,In_851,In_385);
or U2021 (N_2021,In_212,In_357);
or U2022 (N_2022,In_720,In_1029);
nor U2023 (N_2023,In_416,In_1498);
and U2024 (N_2024,In_503,In_309);
nor U2025 (N_2025,In_677,In_186);
nand U2026 (N_2026,In_1032,In_986);
or U2027 (N_2027,In_687,In_913);
xnor U2028 (N_2028,In_995,In_361);
and U2029 (N_2029,In_1139,In_608);
nand U2030 (N_2030,In_1294,In_545);
nor U2031 (N_2031,In_592,In_824);
xor U2032 (N_2032,In_500,In_84);
nor U2033 (N_2033,In_1285,In_95);
and U2034 (N_2034,In_1366,In_457);
nor U2035 (N_2035,In_571,In_306);
nor U2036 (N_2036,In_1424,In_111);
and U2037 (N_2037,In_1431,In_934);
nor U2038 (N_2038,In_369,In_821);
nor U2039 (N_2039,In_1477,In_622);
nor U2040 (N_2040,In_31,In_644);
or U2041 (N_2041,In_1355,In_617);
and U2042 (N_2042,In_444,In_641);
and U2043 (N_2043,In_527,In_1022);
and U2044 (N_2044,In_502,In_636);
and U2045 (N_2045,In_909,In_900);
or U2046 (N_2046,In_1107,In_992);
nand U2047 (N_2047,In_1444,In_1319);
nor U2048 (N_2048,In_1340,In_889);
or U2049 (N_2049,In_515,In_1482);
xnor U2050 (N_2050,In_37,In_244);
and U2051 (N_2051,In_451,In_374);
and U2052 (N_2052,In_894,In_871);
and U2053 (N_2053,In_377,In_431);
or U2054 (N_2054,In_1226,In_568);
nor U2055 (N_2055,In_979,In_1163);
nor U2056 (N_2056,In_901,In_954);
xor U2057 (N_2057,In_1296,In_730);
nor U2058 (N_2058,In_841,In_1063);
or U2059 (N_2059,In_826,In_330);
and U2060 (N_2060,In_266,In_1009);
and U2061 (N_2061,In_908,In_857);
or U2062 (N_2062,In_1391,In_621);
xor U2063 (N_2063,In_1169,In_1301);
nor U2064 (N_2064,In_1482,In_1004);
nand U2065 (N_2065,In_384,In_271);
and U2066 (N_2066,In_472,In_1479);
or U2067 (N_2067,In_382,In_354);
nor U2068 (N_2068,In_1373,In_1099);
and U2069 (N_2069,In_163,In_1281);
or U2070 (N_2070,In_1438,In_40);
nand U2071 (N_2071,In_863,In_559);
nor U2072 (N_2072,In_332,In_309);
or U2073 (N_2073,In_745,In_302);
nor U2074 (N_2074,In_527,In_142);
or U2075 (N_2075,In_1386,In_593);
xnor U2076 (N_2076,In_585,In_1457);
and U2077 (N_2077,In_940,In_6);
or U2078 (N_2078,In_548,In_1328);
or U2079 (N_2079,In_423,In_1334);
nor U2080 (N_2080,In_1323,In_1037);
xor U2081 (N_2081,In_107,In_739);
nor U2082 (N_2082,In_854,In_818);
nor U2083 (N_2083,In_969,In_92);
and U2084 (N_2084,In_1263,In_460);
nand U2085 (N_2085,In_190,In_55);
or U2086 (N_2086,In_950,In_1162);
and U2087 (N_2087,In_1296,In_457);
nor U2088 (N_2088,In_234,In_547);
or U2089 (N_2089,In_1307,In_749);
or U2090 (N_2090,In_1304,In_265);
xnor U2091 (N_2091,In_1464,In_970);
and U2092 (N_2092,In_1219,In_179);
nor U2093 (N_2093,In_985,In_439);
nor U2094 (N_2094,In_972,In_168);
nor U2095 (N_2095,In_185,In_52);
or U2096 (N_2096,In_927,In_403);
or U2097 (N_2097,In_1109,In_913);
nor U2098 (N_2098,In_1089,In_1012);
nand U2099 (N_2099,In_221,In_1126);
nand U2100 (N_2100,In_810,In_634);
or U2101 (N_2101,In_1010,In_700);
nor U2102 (N_2102,In_1315,In_1422);
or U2103 (N_2103,In_131,In_1333);
or U2104 (N_2104,In_1334,In_687);
nand U2105 (N_2105,In_665,In_105);
and U2106 (N_2106,In_844,In_349);
and U2107 (N_2107,In_794,In_1246);
and U2108 (N_2108,In_112,In_34);
and U2109 (N_2109,In_1414,In_179);
or U2110 (N_2110,In_715,In_99);
nand U2111 (N_2111,In_116,In_426);
nand U2112 (N_2112,In_40,In_1408);
and U2113 (N_2113,In_823,In_881);
and U2114 (N_2114,In_1474,In_1255);
nand U2115 (N_2115,In_1421,In_80);
xor U2116 (N_2116,In_1397,In_616);
or U2117 (N_2117,In_1232,In_250);
nand U2118 (N_2118,In_1331,In_1414);
nor U2119 (N_2119,In_616,In_1050);
or U2120 (N_2120,In_1381,In_56);
and U2121 (N_2121,In_806,In_87);
nor U2122 (N_2122,In_1377,In_1100);
nor U2123 (N_2123,In_587,In_913);
and U2124 (N_2124,In_838,In_701);
nand U2125 (N_2125,In_795,In_468);
nand U2126 (N_2126,In_1057,In_491);
nand U2127 (N_2127,In_309,In_123);
nor U2128 (N_2128,In_932,In_1174);
or U2129 (N_2129,In_886,In_286);
or U2130 (N_2130,In_1045,In_1459);
xnor U2131 (N_2131,In_1411,In_1468);
or U2132 (N_2132,In_1283,In_83);
nand U2133 (N_2133,In_118,In_1140);
or U2134 (N_2134,In_995,In_705);
and U2135 (N_2135,In_839,In_244);
or U2136 (N_2136,In_1039,In_748);
nor U2137 (N_2137,In_912,In_455);
or U2138 (N_2138,In_179,In_204);
and U2139 (N_2139,In_110,In_873);
nor U2140 (N_2140,In_686,In_1236);
and U2141 (N_2141,In_998,In_1419);
nor U2142 (N_2142,In_596,In_256);
xnor U2143 (N_2143,In_733,In_81);
nor U2144 (N_2144,In_1415,In_394);
and U2145 (N_2145,In_1259,In_381);
and U2146 (N_2146,In_307,In_71);
nor U2147 (N_2147,In_1214,In_1222);
nand U2148 (N_2148,In_1166,In_94);
nand U2149 (N_2149,In_713,In_668);
xor U2150 (N_2150,In_186,In_1132);
or U2151 (N_2151,In_191,In_1130);
nand U2152 (N_2152,In_1384,In_561);
nor U2153 (N_2153,In_1471,In_882);
and U2154 (N_2154,In_128,In_465);
xnor U2155 (N_2155,In_1211,In_728);
nand U2156 (N_2156,In_1424,In_1254);
or U2157 (N_2157,In_1230,In_895);
and U2158 (N_2158,In_923,In_395);
and U2159 (N_2159,In_769,In_386);
nand U2160 (N_2160,In_13,In_1014);
or U2161 (N_2161,In_330,In_184);
or U2162 (N_2162,In_1497,In_804);
nor U2163 (N_2163,In_524,In_1349);
nor U2164 (N_2164,In_334,In_923);
and U2165 (N_2165,In_1125,In_1448);
nor U2166 (N_2166,In_345,In_264);
xor U2167 (N_2167,In_872,In_22);
xor U2168 (N_2168,In_1202,In_826);
and U2169 (N_2169,In_141,In_1100);
nor U2170 (N_2170,In_420,In_1208);
nor U2171 (N_2171,In_581,In_1145);
nor U2172 (N_2172,In_1279,In_1157);
or U2173 (N_2173,In_1449,In_226);
or U2174 (N_2174,In_215,In_1114);
or U2175 (N_2175,In_601,In_5);
nor U2176 (N_2176,In_749,In_740);
and U2177 (N_2177,In_368,In_599);
nor U2178 (N_2178,In_1268,In_1360);
nand U2179 (N_2179,In_1404,In_1234);
or U2180 (N_2180,In_1368,In_146);
or U2181 (N_2181,In_124,In_1434);
nand U2182 (N_2182,In_400,In_1013);
nand U2183 (N_2183,In_874,In_1397);
and U2184 (N_2184,In_437,In_1128);
nand U2185 (N_2185,In_286,In_39);
or U2186 (N_2186,In_397,In_151);
or U2187 (N_2187,In_1465,In_1372);
or U2188 (N_2188,In_1184,In_749);
nor U2189 (N_2189,In_224,In_175);
nand U2190 (N_2190,In_888,In_885);
nor U2191 (N_2191,In_538,In_768);
nand U2192 (N_2192,In_462,In_457);
nand U2193 (N_2193,In_643,In_1218);
nand U2194 (N_2194,In_1014,In_1096);
xnor U2195 (N_2195,In_604,In_1057);
nand U2196 (N_2196,In_1463,In_960);
or U2197 (N_2197,In_1144,In_501);
or U2198 (N_2198,In_721,In_682);
or U2199 (N_2199,In_699,In_192);
nor U2200 (N_2200,In_1130,In_790);
or U2201 (N_2201,In_346,In_215);
nand U2202 (N_2202,In_1043,In_991);
and U2203 (N_2203,In_1253,In_792);
nor U2204 (N_2204,In_1171,In_1263);
nor U2205 (N_2205,In_453,In_1122);
nand U2206 (N_2206,In_1256,In_1381);
or U2207 (N_2207,In_416,In_784);
nor U2208 (N_2208,In_538,In_712);
nor U2209 (N_2209,In_182,In_682);
and U2210 (N_2210,In_413,In_79);
xnor U2211 (N_2211,In_258,In_704);
nand U2212 (N_2212,In_254,In_479);
nor U2213 (N_2213,In_1359,In_311);
nor U2214 (N_2214,In_259,In_242);
nor U2215 (N_2215,In_294,In_390);
and U2216 (N_2216,In_403,In_522);
and U2217 (N_2217,In_816,In_815);
nand U2218 (N_2218,In_636,In_674);
nor U2219 (N_2219,In_413,In_401);
nand U2220 (N_2220,In_246,In_1332);
and U2221 (N_2221,In_1147,In_548);
nand U2222 (N_2222,In_1279,In_894);
or U2223 (N_2223,In_264,In_1114);
and U2224 (N_2224,In_1322,In_1408);
and U2225 (N_2225,In_1310,In_749);
nor U2226 (N_2226,In_507,In_234);
and U2227 (N_2227,In_185,In_187);
or U2228 (N_2228,In_104,In_786);
and U2229 (N_2229,In_599,In_161);
nor U2230 (N_2230,In_350,In_40);
or U2231 (N_2231,In_1359,In_1265);
or U2232 (N_2232,In_381,In_52);
xor U2233 (N_2233,In_334,In_170);
or U2234 (N_2234,In_736,In_243);
nand U2235 (N_2235,In_553,In_1494);
and U2236 (N_2236,In_747,In_895);
nor U2237 (N_2237,In_1329,In_289);
xnor U2238 (N_2238,In_1288,In_514);
and U2239 (N_2239,In_474,In_506);
or U2240 (N_2240,In_1120,In_992);
and U2241 (N_2241,In_173,In_121);
nand U2242 (N_2242,In_1436,In_624);
and U2243 (N_2243,In_1419,In_884);
or U2244 (N_2244,In_1022,In_1362);
nor U2245 (N_2245,In_852,In_435);
and U2246 (N_2246,In_1188,In_625);
xor U2247 (N_2247,In_1325,In_339);
or U2248 (N_2248,In_1166,In_898);
nand U2249 (N_2249,In_496,In_1233);
nand U2250 (N_2250,In_708,In_1317);
nor U2251 (N_2251,In_293,In_993);
nand U2252 (N_2252,In_216,In_1174);
or U2253 (N_2253,In_1315,In_1444);
nor U2254 (N_2254,In_294,In_753);
and U2255 (N_2255,In_976,In_401);
xnor U2256 (N_2256,In_509,In_716);
or U2257 (N_2257,In_795,In_870);
and U2258 (N_2258,In_1,In_362);
xor U2259 (N_2259,In_481,In_474);
or U2260 (N_2260,In_985,In_59);
nand U2261 (N_2261,In_870,In_876);
or U2262 (N_2262,In_337,In_896);
xnor U2263 (N_2263,In_164,In_831);
nor U2264 (N_2264,In_736,In_1079);
nor U2265 (N_2265,In_636,In_1208);
xor U2266 (N_2266,In_443,In_1323);
nand U2267 (N_2267,In_560,In_478);
nand U2268 (N_2268,In_703,In_982);
nor U2269 (N_2269,In_494,In_1047);
and U2270 (N_2270,In_498,In_60);
nand U2271 (N_2271,In_597,In_804);
nor U2272 (N_2272,In_5,In_195);
nand U2273 (N_2273,In_610,In_1408);
nand U2274 (N_2274,In_1353,In_956);
or U2275 (N_2275,In_73,In_844);
nand U2276 (N_2276,In_1147,In_907);
nand U2277 (N_2277,In_1088,In_967);
and U2278 (N_2278,In_704,In_130);
nor U2279 (N_2279,In_245,In_11);
nand U2280 (N_2280,In_1376,In_1204);
xnor U2281 (N_2281,In_1206,In_525);
and U2282 (N_2282,In_1252,In_424);
or U2283 (N_2283,In_422,In_557);
and U2284 (N_2284,In_717,In_1053);
nor U2285 (N_2285,In_347,In_1399);
nand U2286 (N_2286,In_1421,In_1121);
or U2287 (N_2287,In_1463,In_59);
xnor U2288 (N_2288,In_1042,In_148);
nand U2289 (N_2289,In_250,In_288);
or U2290 (N_2290,In_1316,In_41);
xnor U2291 (N_2291,In_1055,In_707);
and U2292 (N_2292,In_399,In_213);
and U2293 (N_2293,In_1139,In_793);
nand U2294 (N_2294,In_149,In_122);
or U2295 (N_2295,In_1290,In_961);
or U2296 (N_2296,In_838,In_1439);
nand U2297 (N_2297,In_34,In_270);
or U2298 (N_2298,In_498,In_864);
nand U2299 (N_2299,In_858,In_352);
and U2300 (N_2300,In_151,In_19);
and U2301 (N_2301,In_1096,In_774);
nand U2302 (N_2302,In_534,In_218);
nor U2303 (N_2303,In_152,In_1150);
and U2304 (N_2304,In_366,In_828);
nor U2305 (N_2305,In_1064,In_328);
nand U2306 (N_2306,In_769,In_723);
xor U2307 (N_2307,In_1024,In_884);
nor U2308 (N_2308,In_122,In_1185);
nor U2309 (N_2309,In_1040,In_1294);
nor U2310 (N_2310,In_747,In_387);
nand U2311 (N_2311,In_1247,In_134);
and U2312 (N_2312,In_700,In_34);
nor U2313 (N_2313,In_869,In_1214);
and U2314 (N_2314,In_1038,In_1307);
and U2315 (N_2315,In_1194,In_1208);
or U2316 (N_2316,In_663,In_203);
nor U2317 (N_2317,In_1466,In_775);
xor U2318 (N_2318,In_5,In_1285);
and U2319 (N_2319,In_1336,In_1199);
nand U2320 (N_2320,In_582,In_600);
and U2321 (N_2321,In_442,In_1465);
or U2322 (N_2322,In_263,In_1265);
nand U2323 (N_2323,In_855,In_1208);
or U2324 (N_2324,In_1082,In_1038);
and U2325 (N_2325,In_1137,In_667);
nor U2326 (N_2326,In_1068,In_703);
nor U2327 (N_2327,In_166,In_1023);
nand U2328 (N_2328,In_145,In_991);
nor U2329 (N_2329,In_267,In_12);
and U2330 (N_2330,In_1005,In_1177);
and U2331 (N_2331,In_801,In_87);
xnor U2332 (N_2332,In_1205,In_1267);
nor U2333 (N_2333,In_607,In_212);
or U2334 (N_2334,In_1050,In_197);
nand U2335 (N_2335,In_32,In_1484);
or U2336 (N_2336,In_1064,In_450);
nand U2337 (N_2337,In_208,In_1472);
nor U2338 (N_2338,In_399,In_415);
or U2339 (N_2339,In_840,In_1205);
or U2340 (N_2340,In_64,In_555);
and U2341 (N_2341,In_1223,In_1413);
nor U2342 (N_2342,In_341,In_300);
or U2343 (N_2343,In_261,In_348);
nand U2344 (N_2344,In_600,In_520);
xnor U2345 (N_2345,In_1424,In_1067);
and U2346 (N_2346,In_1239,In_142);
nand U2347 (N_2347,In_1438,In_1352);
xor U2348 (N_2348,In_823,In_680);
or U2349 (N_2349,In_901,In_624);
xor U2350 (N_2350,In_187,In_1100);
xnor U2351 (N_2351,In_1332,In_569);
and U2352 (N_2352,In_1495,In_962);
nor U2353 (N_2353,In_1229,In_1139);
and U2354 (N_2354,In_502,In_1177);
or U2355 (N_2355,In_652,In_205);
nor U2356 (N_2356,In_1416,In_15);
nor U2357 (N_2357,In_128,In_988);
and U2358 (N_2358,In_400,In_1125);
nor U2359 (N_2359,In_363,In_315);
nor U2360 (N_2360,In_871,In_742);
nand U2361 (N_2361,In_991,In_1325);
nor U2362 (N_2362,In_641,In_564);
or U2363 (N_2363,In_500,In_1143);
or U2364 (N_2364,In_493,In_871);
and U2365 (N_2365,In_370,In_1105);
xnor U2366 (N_2366,In_1380,In_81);
nand U2367 (N_2367,In_381,In_76);
xor U2368 (N_2368,In_565,In_1284);
or U2369 (N_2369,In_1266,In_82);
nand U2370 (N_2370,In_860,In_351);
or U2371 (N_2371,In_1103,In_56);
nand U2372 (N_2372,In_114,In_905);
and U2373 (N_2373,In_853,In_792);
nor U2374 (N_2374,In_540,In_659);
and U2375 (N_2375,In_675,In_509);
nand U2376 (N_2376,In_508,In_1319);
nand U2377 (N_2377,In_751,In_1070);
xnor U2378 (N_2378,In_195,In_302);
and U2379 (N_2379,In_1287,In_1058);
nor U2380 (N_2380,In_927,In_59);
or U2381 (N_2381,In_1277,In_391);
nand U2382 (N_2382,In_926,In_458);
or U2383 (N_2383,In_1425,In_1060);
and U2384 (N_2384,In_913,In_202);
nand U2385 (N_2385,In_871,In_575);
and U2386 (N_2386,In_1090,In_476);
and U2387 (N_2387,In_496,In_410);
and U2388 (N_2388,In_658,In_1330);
and U2389 (N_2389,In_985,In_1496);
nor U2390 (N_2390,In_1283,In_103);
nor U2391 (N_2391,In_733,In_536);
and U2392 (N_2392,In_525,In_636);
nor U2393 (N_2393,In_711,In_1353);
nor U2394 (N_2394,In_32,In_697);
and U2395 (N_2395,In_1158,In_138);
or U2396 (N_2396,In_1254,In_362);
nor U2397 (N_2397,In_930,In_759);
nand U2398 (N_2398,In_1481,In_588);
or U2399 (N_2399,In_272,In_985);
nor U2400 (N_2400,In_325,In_1488);
nor U2401 (N_2401,In_990,In_885);
or U2402 (N_2402,In_996,In_3);
nand U2403 (N_2403,In_246,In_362);
or U2404 (N_2404,In_33,In_793);
xnor U2405 (N_2405,In_493,In_793);
nor U2406 (N_2406,In_400,In_220);
nor U2407 (N_2407,In_635,In_751);
xnor U2408 (N_2408,In_1021,In_978);
nor U2409 (N_2409,In_341,In_1125);
nor U2410 (N_2410,In_893,In_21);
or U2411 (N_2411,In_89,In_704);
or U2412 (N_2412,In_1484,In_948);
nand U2413 (N_2413,In_217,In_563);
and U2414 (N_2414,In_735,In_539);
nor U2415 (N_2415,In_1136,In_191);
nand U2416 (N_2416,In_300,In_416);
or U2417 (N_2417,In_836,In_168);
or U2418 (N_2418,In_1470,In_549);
nor U2419 (N_2419,In_281,In_1413);
and U2420 (N_2420,In_266,In_716);
nor U2421 (N_2421,In_748,In_513);
or U2422 (N_2422,In_396,In_1335);
and U2423 (N_2423,In_381,In_903);
nor U2424 (N_2424,In_969,In_1460);
or U2425 (N_2425,In_958,In_1001);
nand U2426 (N_2426,In_648,In_567);
or U2427 (N_2427,In_1399,In_692);
and U2428 (N_2428,In_969,In_1278);
nor U2429 (N_2429,In_1498,In_568);
nand U2430 (N_2430,In_181,In_1056);
nor U2431 (N_2431,In_52,In_1371);
and U2432 (N_2432,In_33,In_352);
nor U2433 (N_2433,In_684,In_803);
nor U2434 (N_2434,In_781,In_54);
nand U2435 (N_2435,In_135,In_902);
and U2436 (N_2436,In_364,In_889);
nand U2437 (N_2437,In_604,In_251);
xor U2438 (N_2438,In_502,In_891);
nor U2439 (N_2439,In_263,In_1461);
and U2440 (N_2440,In_1383,In_1021);
xor U2441 (N_2441,In_639,In_233);
or U2442 (N_2442,In_830,In_732);
and U2443 (N_2443,In_1181,In_24);
xnor U2444 (N_2444,In_996,In_697);
and U2445 (N_2445,In_1318,In_133);
nor U2446 (N_2446,In_315,In_695);
and U2447 (N_2447,In_652,In_52);
nor U2448 (N_2448,In_1349,In_240);
or U2449 (N_2449,In_322,In_200);
or U2450 (N_2450,In_1302,In_1477);
or U2451 (N_2451,In_1465,In_943);
nor U2452 (N_2452,In_1449,In_1006);
and U2453 (N_2453,In_88,In_1005);
nand U2454 (N_2454,In_730,In_1352);
nor U2455 (N_2455,In_688,In_947);
nor U2456 (N_2456,In_317,In_949);
xor U2457 (N_2457,In_338,In_379);
nand U2458 (N_2458,In_305,In_906);
or U2459 (N_2459,In_1296,In_864);
nand U2460 (N_2460,In_72,In_145);
nand U2461 (N_2461,In_646,In_948);
nand U2462 (N_2462,In_1209,In_148);
nand U2463 (N_2463,In_893,In_153);
and U2464 (N_2464,In_1377,In_1013);
or U2465 (N_2465,In_312,In_1289);
nand U2466 (N_2466,In_1130,In_623);
nor U2467 (N_2467,In_355,In_113);
xor U2468 (N_2468,In_1050,In_593);
and U2469 (N_2469,In_772,In_1197);
nor U2470 (N_2470,In_1385,In_851);
or U2471 (N_2471,In_1425,In_642);
and U2472 (N_2472,In_1208,In_848);
nor U2473 (N_2473,In_1152,In_618);
or U2474 (N_2474,In_111,In_619);
or U2475 (N_2475,In_1400,In_168);
nor U2476 (N_2476,In_12,In_220);
nand U2477 (N_2477,In_360,In_380);
nand U2478 (N_2478,In_1194,In_1301);
nand U2479 (N_2479,In_4,In_771);
and U2480 (N_2480,In_863,In_879);
nor U2481 (N_2481,In_1467,In_386);
xor U2482 (N_2482,In_306,In_341);
and U2483 (N_2483,In_50,In_1205);
and U2484 (N_2484,In_1446,In_16);
nor U2485 (N_2485,In_1406,In_1293);
nand U2486 (N_2486,In_462,In_724);
or U2487 (N_2487,In_1490,In_152);
or U2488 (N_2488,In_777,In_700);
nor U2489 (N_2489,In_662,In_1373);
and U2490 (N_2490,In_1495,In_79);
nand U2491 (N_2491,In_1435,In_347);
xor U2492 (N_2492,In_1293,In_1374);
and U2493 (N_2493,In_34,In_797);
and U2494 (N_2494,In_3,In_510);
xor U2495 (N_2495,In_260,In_1011);
nand U2496 (N_2496,In_44,In_1271);
nor U2497 (N_2497,In_306,In_1384);
nand U2498 (N_2498,In_303,In_442);
and U2499 (N_2499,In_280,In_636);
and U2500 (N_2500,In_758,In_537);
nand U2501 (N_2501,In_40,In_479);
nand U2502 (N_2502,In_383,In_1363);
nand U2503 (N_2503,In_363,In_652);
and U2504 (N_2504,In_553,In_330);
xor U2505 (N_2505,In_218,In_148);
nand U2506 (N_2506,In_381,In_1344);
nor U2507 (N_2507,In_1333,In_1035);
nor U2508 (N_2508,In_711,In_619);
and U2509 (N_2509,In_472,In_76);
xor U2510 (N_2510,In_567,In_1177);
and U2511 (N_2511,In_1182,In_107);
or U2512 (N_2512,In_1443,In_822);
nor U2513 (N_2513,In_1188,In_1107);
nor U2514 (N_2514,In_1014,In_645);
nor U2515 (N_2515,In_1090,In_34);
xor U2516 (N_2516,In_315,In_1464);
nand U2517 (N_2517,In_614,In_201);
or U2518 (N_2518,In_1378,In_729);
and U2519 (N_2519,In_463,In_167);
nand U2520 (N_2520,In_982,In_481);
xnor U2521 (N_2521,In_1028,In_723);
nor U2522 (N_2522,In_494,In_622);
nor U2523 (N_2523,In_280,In_609);
and U2524 (N_2524,In_658,In_1051);
xor U2525 (N_2525,In_764,In_808);
nand U2526 (N_2526,In_82,In_769);
and U2527 (N_2527,In_1180,In_1183);
or U2528 (N_2528,In_237,In_780);
or U2529 (N_2529,In_1212,In_295);
nor U2530 (N_2530,In_518,In_586);
or U2531 (N_2531,In_351,In_872);
or U2532 (N_2532,In_378,In_393);
or U2533 (N_2533,In_1134,In_929);
and U2534 (N_2534,In_379,In_198);
and U2535 (N_2535,In_504,In_1417);
nand U2536 (N_2536,In_220,In_343);
xnor U2537 (N_2537,In_1034,In_156);
nand U2538 (N_2538,In_990,In_949);
and U2539 (N_2539,In_721,In_1014);
nand U2540 (N_2540,In_1321,In_362);
xnor U2541 (N_2541,In_558,In_326);
nand U2542 (N_2542,In_1080,In_303);
or U2543 (N_2543,In_188,In_19);
or U2544 (N_2544,In_42,In_241);
and U2545 (N_2545,In_292,In_364);
nor U2546 (N_2546,In_1286,In_1077);
nand U2547 (N_2547,In_366,In_407);
and U2548 (N_2548,In_763,In_645);
xnor U2549 (N_2549,In_253,In_1236);
xnor U2550 (N_2550,In_701,In_706);
nand U2551 (N_2551,In_1197,In_1090);
or U2552 (N_2552,In_949,In_1199);
or U2553 (N_2553,In_491,In_411);
or U2554 (N_2554,In_645,In_585);
nand U2555 (N_2555,In_1266,In_698);
nor U2556 (N_2556,In_161,In_281);
nor U2557 (N_2557,In_1043,In_60);
nor U2558 (N_2558,In_434,In_685);
nor U2559 (N_2559,In_1203,In_94);
nor U2560 (N_2560,In_100,In_660);
nand U2561 (N_2561,In_1152,In_365);
or U2562 (N_2562,In_129,In_18);
or U2563 (N_2563,In_662,In_540);
and U2564 (N_2564,In_1484,In_710);
xnor U2565 (N_2565,In_321,In_193);
nand U2566 (N_2566,In_146,In_320);
xnor U2567 (N_2567,In_969,In_1018);
xor U2568 (N_2568,In_150,In_870);
or U2569 (N_2569,In_581,In_601);
and U2570 (N_2570,In_1089,In_79);
or U2571 (N_2571,In_1423,In_1313);
xor U2572 (N_2572,In_1459,In_646);
nand U2573 (N_2573,In_326,In_1336);
nand U2574 (N_2574,In_423,In_366);
xnor U2575 (N_2575,In_559,In_24);
or U2576 (N_2576,In_595,In_174);
nor U2577 (N_2577,In_917,In_884);
or U2578 (N_2578,In_1284,In_1413);
nand U2579 (N_2579,In_753,In_969);
xor U2580 (N_2580,In_606,In_1477);
and U2581 (N_2581,In_159,In_1493);
nand U2582 (N_2582,In_424,In_776);
or U2583 (N_2583,In_1377,In_348);
nand U2584 (N_2584,In_472,In_480);
nor U2585 (N_2585,In_415,In_1139);
nor U2586 (N_2586,In_911,In_71);
nand U2587 (N_2587,In_1423,In_415);
and U2588 (N_2588,In_544,In_788);
nand U2589 (N_2589,In_593,In_682);
xor U2590 (N_2590,In_686,In_371);
nand U2591 (N_2591,In_959,In_1140);
and U2592 (N_2592,In_944,In_1052);
and U2593 (N_2593,In_1034,In_545);
nand U2594 (N_2594,In_310,In_630);
and U2595 (N_2595,In_751,In_539);
and U2596 (N_2596,In_527,In_1252);
nand U2597 (N_2597,In_317,In_591);
nand U2598 (N_2598,In_0,In_510);
xnor U2599 (N_2599,In_1387,In_700);
and U2600 (N_2600,In_694,In_428);
or U2601 (N_2601,In_831,In_580);
or U2602 (N_2602,In_669,In_697);
and U2603 (N_2603,In_821,In_410);
nand U2604 (N_2604,In_182,In_961);
nor U2605 (N_2605,In_435,In_774);
nor U2606 (N_2606,In_726,In_1275);
or U2607 (N_2607,In_331,In_813);
and U2608 (N_2608,In_806,In_618);
and U2609 (N_2609,In_1352,In_784);
nor U2610 (N_2610,In_711,In_283);
and U2611 (N_2611,In_99,In_1426);
nor U2612 (N_2612,In_496,In_879);
or U2613 (N_2613,In_960,In_609);
and U2614 (N_2614,In_1478,In_930);
nand U2615 (N_2615,In_1362,In_1238);
nand U2616 (N_2616,In_1355,In_1006);
nand U2617 (N_2617,In_1313,In_634);
or U2618 (N_2618,In_916,In_531);
and U2619 (N_2619,In_1282,In_1230);
nand U2620 (N_2620,In_782,In_571);
and U2621 (N_2621,In_595,In_520);
or U2622 (N_2622,In_349,In_289);
nor U2623 (N_2623,In_1196,In_37);
and U2624 (N_2624,In_680,In_464);
nor U2625 (N_2625,In_809,In_515);
or U2626 (N_2626,In_1219,In_987);
nand U2627 (N_2627,In_1348,In_425);
or U2628 (N_2628,In_950,In_1259);
or U2629 (N_2629,In_840,In_281);
and U2630 (N_2630,In_921,In_1477);
and U2631 (N_2631,In_1362,In_780);
nor U2632 (N_2632,In_346,In_973);
and U2633 (N_2633,In_1158,In_881);
xnor U2634 (N_2634,In_1263,In_875);
nor U2635 (N_2635,In_903,In_598);
nor U2636 (N_2636,In_724,In_307);
or U2637 (N_2637,In_737,In_973);
or U2638 (N_2638,In_137,In_842);
nor U2639 (N_2639,In_1460,In_1463);
nor U2640 (N_2640,In_61,In_691);
and U2641 (N_2641,In_82,In_908);
and U2642 (N_2642,In_1199,In_608);
xor U2643 (N_2643,In_505,In_1109);
or U2644 (N_2644,In_1461,In_225);
and U2645 (N_2645,In_5,In_630);
nor U2646 (N_2646,In_181,In_1042);
nor U2647 (N_2647,In_859,In_393);
or U2648 (N_2648,In_819,In_804);
or U2649 (N_2649,In_248,In_1346);
nor U2650 (N_2650,In_508,In_1417);
nand U2651 (N_2651,In_810,In_270);
xnor U2652 (N_2652,In_365,In_73);
nor U2653 (N_2653,In_6,In_172);
and U2654 (N_2654,In_836,In_1232);
nor U2655 (N_2655,In_434,In_806);
nor U2656 (N_2656,In_1419,In_625);
xor U2657 (N_2657,In_357,In_457);
or U2658 (N_2658,In_1262,In_525);
and U2659 (N_2659,In_547,In_788);
nand U2660 (N_2660,In_867,In_1268);
or U2661 (N_2661,In_1326,In_213);
nand U2662 (N_2662,In_288,In_642);
nand U2663 (N_2663,In_624,In_441);
or U2664 (N_2664,In_1496,In_1216);
or U2665 (N_2665,In_113,In_270);
or U2666 (N_2666,In_1261,In_133);
nand U2667 (N_2667,In_1341,In_1123);
and U2668 (N_2668,In_1150,In_1353);
or U2669 (N_2669,In_1350,In_1047);
and U2670 (N_2670,In_1048,In_975);
or U2671 (N_2671,In_1162,In_21);
and U2672 (N_2672,In_1154,In_703);
or U2673 (N_2673,In_748,In_20);
or U2674 (N_2674,In_836,In_1071);
nor U2675 (N_2675,In_842,In_460);
and U2676 (N_2676,In_56,In_889);
nor U2677 (N_2677,In_694,In_988);
nand U2678 (N_2678,In_1067,In_42);
or U2679 (N_2679,In_423,In_1432);
xor U2680 (N_2680,In_1285,In_226);
or U2681 (N_2681,In_334,In_1062);
nand U2682 (N_2682,In_642,In_703);
nand U2683 (N_2683,In_144,In_793);
xnor U2684 (N_2684,In_1174,In_1236);
nand U2685 (N_2685,In_295,In_1243);
nor U2686 (N_2686,In_43,In_288);
nor U2687 (N_2687,In_20,In_305);
nand U2688 (N_2688,In_295,In_598);
nand U2689 (N_2689,In_751,In_1345);
nand U2690 (N_2690,In_422,In_1409);
and U2691 (N_2691,In_99,In_1064);
or U2692 (N_2692,In_1370,In_741);
and U2693 (N_2693,In_1412,In_89);
nor U2694 (N_2694,In_434,In_945);
or U2695 (N_2695,In_1164,In_459);
nand U2696 (N_2696,In_645,In_292);
or U2697 (N_2697,In_283,In_1154);
or U2698 (N_2698,In_350,In_10);
and U2699 (N_2699,In_867,In_814);
xnor U2700 (N_2700,In_1349,In_1327);
or U2701 (N_2701,In_664,In_1);
xor U2702 (N_2702,In_94,In_718);
or U2703 (N_2703,In_947,In_448);
nor U2704 (N_2704,In_696,In_441);
nand U2705 (N_2705,In_319,In_780);
or U2706 (N_2706,In_678,In_460);
xnor U2707 (N_2707,In_1165,In_242);
or U2708 (N_2708,In_338,In_77);
nand U2709 (N_2709,In_1268,In_914);
nor U2710 (N_2710,In_78,In_355);
and U2711 (N_2711,In_1016,In_175);
xor U2712 (N_2712,In_357,In_870);
nand U2713 (N_2713,In_23,In_796);
nand U2714 (N_2714,In_1061,In_375);
nand U2715 (N_2715,In_813,In_13);
nor U2716 (N_2716,In_975,In_318);
xor U2717 (N_2717,In_1174,In_1261);
or U2718 (N_2718,In_372,In_1192);
and U2719 (N_2719,In_844,In_160);
xnor U2720 (N_2720,In_1280,In_74);
nor U2721 (N_2721,In_1180,In_181);
or U2722 (N_2722,In_1324,In_1189);
and U2723 (N_2723,In_1486,In_227);
nor U2724 (N_2724,In_1275,In_772);
nand U2725 (N_2725,In_1105,In_825);
nor U2726 (N_2726,In_174,In_1106);
and U2727 (N_2727,In_1073,In_814);
nor U2728 (N_2728,In_949,In_400);
or U2729 (N_2729,In_1485,In_149);
nand U2730 (N_2730,In_940,In_1449);
and U2731 (N_2731,In_193,In_345);
xnor U2732 (N_2732,In_221,In_340);
nor U2733 (N_2733,In_667,In_359);
nand U2734 (N_2734,In_1327,In_726);
or U2735 (N_2735,In_1468,In_366);
and U2736 (N_2736,In_981,In_1054);
and U2737 (N_2737,In_109,In_1173);
xnor U2738 (N_2738,In_1470,In_201);
and U2739 (N_2739,In_738,In_469);
or U2740 (N_2740,In_1129,In_952);
nor U2741 (N_2741,In_442,In_188);
or U2742 (N_2742,In_155,In_83);
xor U2743 (N_2743,In_1379,In_954);
nor U2744 (N_2744,In_750,In_255);
nand U2745 (N_2745,In_1300,In_1059);
nor U2746 (N_2746,In_1279,In_1363);
nor U2747 (N_2747,In_1200,In_163);
xor U2748 (N_2748,In_157,In_5);
or U2749 (N_2749,In_912,In_925);
and U2750 (N_2750,In_248,In_1249);
nand U2751 (N_2751,In_636,In_566);
nand U2752 (N_2752,In_1022,In_618);
nor U2753 (N_2753,In_862,In_550);
nand U2754 (N_2754,In_936,In_505);
nor U2755 (N_2755,In_524,In_1139);
nor U2756 (N_2756,In_1031,In_739);
nand U2757 (N_2757,In_1186,In_1313);
xnor U2758 (N_2758,In_1391,In_740);
nor U2759 (N_2759,In_303,In_640);
nand U2760 (N_2760,In_621,In_475);
and U2761 (N_2761,In_610,In_499);
and U2762 (N_2762,In_575,In_1019);
nand U2763 (N_2763,In_574,In_483);
nand U2764 (N_2764,In_8,In_310);
nand U2765 (N_2765,In_121,In_711);
and U2766 (N_2766,In_1381,In_450);
and U2767 (N_2767,In_48,In_1302);
nor U2768 (N_2768,In_198,In_395);
nor U2769 (N_2769,In_632,In_15);
and U2770 (N_2770,In_1058,In_726);
and U2771 (N_2771,In_369,In_954);
nand U2772 (N_2772,In_991,In_142);
nor U2773 (N_2773,In_902,In_675);
and U2774 (N_2774,In_325,In_110);
or U2775 (N_2775,In_1304,In_68);
nor U2776 (N_2776,In_64,In_684);
xnor U2777 (N_2777,In_1488,In_144);
nand U2778 (N_2778,In_1142,In_798);
nand U2779 (N_2779,In_996,In_1488);
and U2780 (N_2780,In_302,In_295);
or U2781 (N_2781,In_332,In_1494);
or U2782 (N_2782,In_420,In_293);
and U2783 (N_2783,In_62,In_612);
nand U2784 (N_2784,In_1228,In_1304);
nor U2785 (N_2785,In_145,In_1179);
nor U2786 (N_2786,In_1358,In_90);
nor U2787 (N_2787,In_1065,In_1449);
and U2788 (N_2788,In_581,In_1100);
or U2789 (N_2789,In_877,In_1090);
nor U2790 (N_2790,In_14,In_497);
nor U2791 (N_2791,In_102,In_969);
and U2792 (N_2792,In_1446,In_78);
nand U2793 (N_2793,In_607,In_1412);
and U2794 (N_2794,In_1241,In_824);
and U2795 (N_2795,In_1033,In_788);
or U2796 (N_2796,In_1033,In_1298);
nand U2797 (N_2797,In_1468,In_433);
xnor U2798 (N_2798,In_288,In_1035);
nand U2799 (N_2799,In_1479,In_433);
xor U2800 (N_2800,In_1295,In_717);
nor U2801 (N_2801,In_971,In_601);
or U2802 (N_2802,In_1263,In_317);
and U2803 (N_2803,In_847,In_153);
nand U2804 (N_2804,In_680,In_1368);
nand U2805 (N_2805,In_1122,In_692);
nor U2806 (N_2806,In_953,In_390);
and U2807 (N_2807,In_449,In_89);
nor U2808 (N_2808,In_1033,In_1237);
or U2809 (N_2809,In_1306,In_49);
xor U2810 (N_2810,In_317,In_106);
nand U2811 (N_2811,In_312,In_1186);
and U2812 (N_2812,In_1448,In_583);
nor U2813 (N_2813,In_1150,In_118);
and U2814 (N_2814,In_114,In_1333);
nand U2815 (N_2815,In_707,In_431);
and U2816 (N_2816,In_598,In_341);
nand U2817 (N_2817,In_946,In_976);
or U2818 (N_2818,In_687,In_1442);
nand U2819 (N_2819,In_372,In_169);
or U2820 (N_2820,In_758,In_266);
and U2821 (N_2821,In_864,In_771);
nand U2822 (N_2822,In_357,In_776);
nor U2823 (N_2823,In_1461,In_27);
nor U2824 (N_2824,In_1454,In_538);
or U2825 (N_2825,In_849,In_221);
xor U2826 (N_2826,In_743,In_290);
nor U2827 (N_2827,In_810,In_577);
or U2828 (N_2828,In_1048,In_602);
and U2829 (N_2829,In_354,In_1116);
xnor U2830 (N_2830,In_537,In_216);
nor U2831 (N_2831,In_875,In_730);
xnor U2832 (N_2832,In_156,In_185);
nand U2833 (N_2833,In_1406,In_1346);
and U2834 (N_2834,In_710,In_124);
and U2835 (N_2835,In_489,In_670);
nand U2836 (N_2836,In_1469,In_114);
nor U2837 (N_2837,In_919,In_1293);
and U2838 (N_2838,In_1408,In_698);
and U2839 (N_2839,In_393,In_893);
nand U2840 (N_2840,In_1057,In_323);
nor U2841 (N_2841,In_633,In_660);
nor U2842 (N_2842,In_461,In_43);
nand U2843 (N_2843,In_774,In_325);
nand U2844 (N_2844,In_226,In_814);
nand U2845 (N_2845,In_657,In_1408);
nor U2846 (N_2846,In_514,In_993);
and U2847 (N_2847,In_256,In_671);
nand U2848 (N_2848,In_1263,In_458);
nor U2849 (N_2849,In_728,In_540);
nor U2850 (N_2850,In_1414,In_1307);
or U2851 (N_2851,In_838,In_1114);
or U2852 (N_2852,In_603,In_565);
nand U2853 (N_2853,In_866,In_583);
or U2854 (N_2854,In_1214,In_762);
nor U2855 (N_2855,In_362,In_781);
xnor U2856 (N_2856,In_1242,In_642);
xnor U2857 (N_2857,In_3,In_774);
nand U2858 (N_2858,In_657,In_496);
xnor U2859 (N_2859,In_1169,In_951);
xnor U2860 (N_2860,In_1029,In_857);
nor U2861 (N_2861,In_161,In_326);
nand U2862 (N_2862,In_1054,In_172);
nand U2863 (N_2863,In_437,In_577);
or U2864 (N_2864,In_445,In_480);
nor U2865 (N_2865,In_743,In_117);
nand U2866 (N_2866,In_1443,In_346);
or U2867 (N_2867,In_1346,In_356);
or U2868 (N_2868,In_1093,In_408);
xor U2869 (N_2869,In_84,In_1223);
xnor U2870 (N_2870,In_954,In_610);
and U2871 (N_2871,In_1008,In_946);
nand U2872 (N_2872,In_845,In_463);
xnor U2873 (N_2873,In_30,In_1498);
nand U2874 (N_2874,In_460,In_199);
nor U2875 (N_2875,In_654,In_605);
xnor U2876 (N_2876,In_1165,In_1246);
or U2877 (N_2877,In_448,In_958);
xnor U2878 (N_2878,In_1065,In_573);
and U2879 (N_2879,In_1442,In_70);
nor U2880 (N_2880,In_1297,In_1282);
or U2881 (N_2881,In_466,In_902);
nor U2882 (N_2882,In_149,In_678);
or U2883 (N_2883,In_743,In_918);
nand U2884 (N_2884,In_366,In_626);
nand U2885 (N_2885,In_1322,In_632);
nor U2886 (N_2886,In_410,In_28);
nor U2887 (N_2887,In_604,In_231);
and U2888 (N_2888,In_1292,In_1287);
nand U2889 (N_2889,In_1024,In_530);
nand U2890 (N_2890,In_1174,In_381);
or U2891 (N_2891,In_1472,In_855);
or U2892 (N_2892,In_1373,In_1379);
or U2893 (N_2893,In_684,In_812);
nor U2894 (N_2894,In_1256,In_986);
or U2895 (N_2895,In_605,In_955);
nor U2896 (N_2896,In_1376,In_1144);
nand U2897 (N_2897,In_177,In_180);
and U2898 (N_2898,In_1478,In_778);
nand U2899 (N_2899,In_141,In_1270);
or U2900 (N_2900,In_160,In_1354);
or U2901 (N_2901,In_159,In_899);
and U2902 (N_2902,In_286,In_374);
nor U2903 (N_2903,In_700,In_1326);
nand U2904 (N_2904,In_782,In_438);
nor U2905 (N_2905,In_1181,In_884);
nand U2906 (N_2906,In_439,In_332);
nor U2907 (N_2907,In_573,In_978);
and U2908 (N_2908,In_1303,In_700);
and U2909 (N_2909,In_724,In_1383);
and U2910 (N_2910,In_440,In_710);
or U2911 (N_2911,In_253,In_1279);
nand U2912 (N_2912,In_1499,In_1186);
and U2913 (N_2913,In_807,In_392);
or U2914 (N_2914,In_935,In_890);
nor U2915 (N_2915,In_1091,In_603);
or U2916 (N_2916,In_561,In_1234);
xor U2917 (N_2917,In_1243,In_1463);
or U2918 (N_2918,In_464,In_721);
nor U2919 (N_2919,In_532,In_597);
and U2920 (N_2920,In_514,In_967);
or U2921 (N_2921,In_1298,In_160);
nand U2922 (N_2922,In_1142,In_973);
nor U2923 (N_2923,In_210,In_537);
or U2924 (N_2924,In_585,In_1303);
nor U2925 (N_2925,In_1411,In_217);
and U2926 (N_2926,In_1051,In_747);
nand U2927 (N_2927,In_1343,In_1394);
or U2928 (N_2928,In_1213,In_583);
nor U2929 (N_2929,In_190,In_1188);
nand U2930 (N_2930,In_901,In_1178);
nor U2931 (N_2931,In_653,In_1400);
nor U2932 (N_2932,In_744,In_1143);
or U2933 (N_2933,In_798,In_1069);
nand U2934 (N_2934,In_332,In_1499);
xor U2935 (N_2935,In_714,In_1278);
xnor U2936 (N_2936,In_1042,In_411);
nor U2937 (N_2937,In_589,In_1073);
nor U2938 (N_2938,In_143,In_997);
nand U2939 (N_2939,In_1461,In_1142);
nor U2940 (N_2940,In_588,In_885);
nor U2941 (N_2941,In_1238,In_880);
and U2942 (N_2942,In_799,In_307);
nor U2943 (N_2943,In_621,In_255);
and U2944 (N_2944,In_1299,In_336);
nand U2945 (N_2945,In_855,In_282);
nor U2946 (N_2946,In_1317,In_464);
nor U2947 (N_2947,In_255,In_440);
nand U2948 (N_2948,In_1222,In_411);
nand U2949 (N_2949,In_293,In_918);
nand U2950 (N_2950,In_213,In_367);
nand U2951 (N_2951,In_738,In_514);
and U2952 (N_2952,In_987,In_1415);
nand U2953 (N_2953,In_63,In_91);
and U2954 (N_2954,In_322,In_590);
xor U2955 (N_2955,In_711,In_229);
nor U2956 (N_2956,In_1364,In_1005);
nor U2957 (N_2957,In_1272,In_253);
and U2958 (N_2958,In_867,In_714);
or U2959 (N_2959,In_174,In_204);
and U2960 (N_2960,In_1469,In_1156);
xnor U2961 (N_2961,In_37,In_1240);
or U2962 (N_2962,In_714,In_653);
nand U2963 (N_2963,In_279,In_1219);
nand U2964 (N_2964,In_119,In_1091);
nor U2965 (N_2965,In_641,In_787);
and U2966 (N_2966,In_216,In_1488);
and U2967 (N_2967,In_1349,In_1437);
and U2968 (N_2968,In_1062,In_324);
nor U2969 (N_2969,In_1498,In_921);
xnor U2970 (N_2970,In_1116,In_38);
or U2971 (N_2971,In_1424,In_253);
xor U2972 (N_2972,In_48,In_1154);
and U2973 (N_2973,In_1249,In_903);
and U2974 (N_2974,In_808,In_317);
nand U2975 (N_2975,In_542,In_1056);
nor U2976 (N_2976,In_492,In_1330);
nor U2977 (N_2977,In_665,In_124);
nand U2978 (N_2978,In_1151,In_523);
nand U2979 (N_2979,In_961,In_314);
or U2980 (N_2980,In_815,In_105);
and U2981 (N_2981,In_1342,In_659);
and U2982 (N_2982,In_412,In_1091);
nor U2983 (N_2983,In_1245,In_1136);
and U2984 (N_2984,In_77,In_142);
or U2985 (N_2985,In_309,In_1130);
nand U2986 (N_2986,In_726,In_215);
nor U2987 (N_2987,In_212,In_233);
nand U2988 (N_2988,In_1378,In_1146);
xnor U2989 (N_2989,In_193,In_1310);
and U2990 (N_2990,In_1163,In_248);
nand U2991 (N_2991,In_1233,In_1404);
or U2992 (N_2992,In_615,In_1147);
nor U2993 (N_2993,In_475,In_257);
nor U2994 (N_2994,In_1150,In_1442);
nor U2995 (N_2995,In_250,In_639);
nor U2996 (N_2996,In_717,In_897);
nor U2997 (N_2997,In_455,In_1185);
or U2998 (N_2998,In_559,In_246);
or U2999 (N_2999,In_203,In_561);
nand U3000 (N_3000,N_1175,N_1345);
or U3001 (N_3001,N_6,N_589);
and U3002 (N_3002,N_2290,N_395);
xor U3003 (N_3003,N_2042,N_1853);
or U3004 (N_3004,N_543,N_1543);
and U3005 (N_3005,N_2185,N_1442);
nor U3006 (N_3006,N_91,N_448);
and U3007 (N_3007,N_2194,N_2075);
and U3008 (N_3008,N_979,N_1876);
and U3009 (N_3009,N_2444,N_1036);
nand U3010 (N_3010,N_116,N_1745);
nand U3011 (N_3011,N_1051,N_2678);
and U3012 (N_3012,N_2221,N_936);
or U3013 (N_3013,N_970,N_1172);
nand U3014 (N_3014,N_1819,N_1576);
or U3015 (N_3015,N_859,N_2993);
and U3016 (N_3016,N_2601,N_481);
or U3017 (N_3017,N_1326,N_1188);
and U3018 (N_3018,N_1417,N_2328);
nor U3019 (N_3019,N_2521,N_1547);
or U3020 (N_3020,N_2284,N_2522);
and U3021 (N_3021,N_2548,N_178);
and U3022 (N_3022,N_1756,N_2100);
or U3023 (N_3023,N_2389,N_1041);
nor U3024 (N_3024,N_851,N_260);
and U3025 (N_3025,N_469,N_1696);
or U3026 (N_3026,N_510,N_682);
xnor U3027 (N_3027,N_2200,N_611);
or U3028 (N_3028,N_313,N_2062);
nand U3029 (N_3029,N_1142,N_276);
nor U3030 (N_3030,N_2241,N_858);
nand U3031 (N_3031,N_376,N_79);
or U3032 (N_3032,N_645,N_226);
or U3033 (N_3033,N_1080,N_660);
and U3034 (N_3034,N_1094,N_2168);
or U3035 (N_3035,N_2503,N_2554);
and U3036 (N_3036,N_1771,N_1362);
and U3037 (N_3037,N_2416,N_121);
xor U3038 (N_3038,N_2064,N_2225);
nor U3039 (N_3039,N_1789,N_1243);
or U3040 (N_3040,N_2442,N_2486);
or U3041 (N_3041,N_2836,N_102);
nor U3042 (N_3042,N_72,N_1602);
nor U3043 (N_3043,N_2512,N_2545);
nor U3044 (N_3044,N_967,N_1831);
or U3045 (N_3045,N_1770,N_2080);
nand U3046 (N_3046,N_1485,N_1758);
nand U3047 (N_3047,N_278,N_2806);
nor U3048 (N_3048,N_1753,N_2923);
xnor U3049 (N_3049,N_406,N_8);
or U3050 (N_3050,N_1062,N_497);
or U3051 (N_3051,N_777,N_542);
xnor U3052 (N_3052,N_2296,N_1426);
nor U3053 (N_3053,N_2203,N_2038);
nor U3054 (N_3054,N_2013,N_961);
nor U3055 (N_3055,N_257,N_1215);
or U3056 (N_3056,N_45,N_2291);
xnor U3057 (N_3057,N_1286,N_1290);
nor U3058 (N_3058,N_1500,N_2795);
or U3059 (N_3059,N_1261,N_929);
nor U3060 (N_3060,N_427,N_1450);
xor U3061 (N_3061,N_1058,N_2541);
or U3062 (N_3062,N_2857,N_1922);
nor U3063 (N_3063,N_838,N_2798);
and U3064 (N_3064,N_2269,N_1887);
nand U3065 (N_3065,N_648,N_1757);
nor U3066 (N_3066,N_2010,N_1901);
and U3067 (N_3067,N_1519,N_1454);
nor U3068 (N_3068,N_1119,N_1480);
or U3069 (N_3069,N_1681,N_799);
nor U3070 (N_3070,N_1407,N_2621);
nand U3071 (N_3071,N_797,N_2178);
and U3072 (N_3072,N_2292,N_356);
or U3073 (N_3073,N_1586,N_605);
xnor U3074 (N_3074,N_1455,N_2353);
nand U3075 (N_3075,N_2327,N_2563);
and U3076 (N_3076,N_2189,N_2330);
and U3077 (N_3077,N_2305,N_1106);
nand U3078 (N_3078,N_656,N_179);
and U3079 (N_3079,N_839,N_2591);
nand U3080 (N_3080,N_2282,N_2137);
or U3081 (N_3081,N_1779,N_1039);
nand U3082 (N_3082,N_1137,N_142);
and U3083 (N_3083,N_517,N_1239);
nor U3084 (N_3084,N_1538,N_1697);
and U3085 (N_3085,N_2164,N_1025);
and U3086 (N_3086,N_1312,N_775);
and U3087 (N_3087,N_2415,N_138);
and U3088 (N_3088,N_124,N_2248);
xor U3089 (N_3089,N_2264,N_1109);
nor U3090 (N_3090,N_1662,N_1324);
nand U3091 (N_3091,N_1231,N_2147);
or U3092 (N_3092,N_1105,N_2287);
nor U3093 (N_3093,N_2577,N_506);
or U3094 (N_3094,N_403,N_1221);
nor U3095 (N_3095,N_1459,N_240);
nand U3096 (N_3096,N_1552,N_1280);
or U3097 (N_3097,N_1823,N_1673);
or U3098 (N_3098,N_2125,N_2155);
or U3099 (N_3099,N_225,N_2050);
nand U3100 (N_3100,N_1120,N_1490);
nand U3101 (N_3101,N_399,N_2602);
and U3102 (N_3102,N_1600,N_466);
or U3103 (N_3103,N_2868,N_1037);
and U3104 (N_3104,N_1850,N_445);
nand U3105 (N_3105,N_744,N_2054);
nand U3106 (N_3106,N_2238,N_2344);
and U3107 (N_3107,N_2253,N_455);
nor U3108 (N_3108,N_1319,N_2371);
and U3109 (N_3109,N_2373,N_1002);
nand U3110 (N_3110,N_2136,N_2703);
nand U3111 (N_3111,N_2640,N_1619);
or U3112 (N_3112,N_2524,N_1683);
or U3113 (N_3113,N_1100,N_2025);
and U3114 (N_3114,N_1020,N_1699);
and U3115 (N_3115,N_2994,N_493);
or U3116 (N_3116,N_562,N_1323);
and U3117 (N_3117,N_103,N_2874);
or U3118 (N_3118,N_702,N_1361);
or U3119 (N_3119,N_2466,N_378);
or U3120 (N_3120,N_1179,N_2504);
xnor U3121 (N_3121,N_675,N_783);
nor U3122 (N_3122,N_2097,N_1655);
nand U3123 (N_3123,N_640,N_2308);
nand U3124 (N_3124,N_1688,N_1408);
nor U3125 (N_3125,N_1936,N_2793);
or U3126 (N_3126,N_2193,N_2707);
nor U3127 (N_3127,N_773,N_734);
nand U3128 (N_3128,N_1928,N_2052);
or U3129 (N_3129,N_1768,N_2905);
and U3130 (N_3130,N_1759,N_1372);
or U3131 (N_3131,N_1629,N_2260);
nor U3132 (N_3132,N_342,N_2511);
nand U3133 (N_3133,N_1028,N_1401);
and U3134 (N_3134,N_76,N_1820);
or U3135 (N_3135,N_853,N_26);
nand U3136 (N_3136,N_243,N_172);
or U3137 (N_3137,N_1703,N_1065);
and U3138 (N_3138,N_1659,N_2576);
nor U3139 (N_3139,N_1118,N_355);
or U3140 (N_3140,N_1712,N_1856);
nor U3141 (N_3141,N_41,N_1382);
and U3142 (N_3142,N_1515,N_1103);
and U3143 (N_3143,N_426,N_2870);
or U3144 (N_3144,N_423,N_1321);
nor U3145 (N_3145,N_89,N_1405);
nand U3146 (N_3146,N_2679,N_279);
xor U3147 (N_3147,N_2632,N_495);
nand U3148 (N_3148,N_2370,N_610);
or U3149 (N_3149,N_2564,N_1066);
nor U3150 (N_3150,N_1872,N_2907);
nor U3151 (N_3151,N_2711,N_860);
nor U3152 (N_3152,N_2633,N_126);
or U3153 (N_3153,N_255,N_2885);
nor U3154 (N_3154,N_889,N_2560);
or U3155 (N_3155,N_900,N_1915);
nand U3156 (N_3156,N_221,N_1102);
and U3157 (N_3157,N_1945,N_2830);
xnor U3158 (N_3158,N_1909,N_2172);
or U3159 (N_3159,N_244,N_1236);
nand U3160 (N_3160,N_987,N_1007);
nand U3161 (N_3161,N_614,N_33);
xnor U3162 (N_3162,N_380,N_2005);
nor U3163 (N_3163,N_2598,N_2951);
nand U3164 (N_3164,N_837,N_812);
or U3165 (N_3165,N_2761,N_2778);
and U3166 (N_3166,N_2686,N_1775);
or U3167 (N_3167,N_252,N_2334);
nand U3168 (N_3168,N_820,N_2614);
nor U3169 (N_3169,N_271,N_291);
nand U3170 (N_3170,N_104,N_1948);
nand U3171 (N_3171,N_2805,N_105);
xnor U3172 (N_3172,N_1839,N_934);
or U3173 (N_3173,N_2099,N_16);
nand U3174 (N_3174,N_1706,N_1514);
or U3175 (N_3175,N_2413,N_1391);
nor U3176 (N_3176,N_1938,N_277);
nand U3177 (N_3177,N_396,N_2822);
or U3178 (N_3178,N_364,N_2255);
xnor U3179 (N_3179,N_208,N_1388);
or U3180 (N_3180,N_2692,N_2086);
nor U3181 (N_3181,N_603,N_1708);
and U3182 (N_3182,N_75,N_2457);
and U3183 (N_3183,N_841,N_1487);
and U3184 (N_3184,N_1709,N_1446);
nand U3185 (N_3185,N_1539,N_262);
nand U3186 (N_3186,N_2072,N_1976);
and U3187 (N_3187,N_397,N_2683);
xnor U3188 (N_3188,N_317,N_2908);
nor U3189 (N_3189,N_459,N_281);
nor U3190 (N_3190,N_84,N_1496);
and U3191 (N_3191,N_654,N_2842);
nor U3192 (N_3192,N_2694,N_2324);
and U3193 (N_3193,N_2398,N_548);
or U3194 (N_3194,N_1344,N_2397);
nor U3195 (N_3195,N_2517,N_1615);
and U3196 (N_3196,N_1184,N_2910);
and U3197 (N_3197,N_1988,N_2819);
or U3198 (N_3198,N_625,N_2505);
or U3199 (N_3199,N_1849,N_1468);
or U3200 (N_3200,N_2906,N_253);
nand U3201 (N_3201,N_442,N_995);
or U3202 (N_3202,N_1420,N_2572);
nor U3203 (N_3203,N_350,N_2379);
xnor U3204 (N_3204,N_2783,N_1916);
nand U3205 (N_3205,N_204,N_192);
and U3206 (N_3206,N_98,N_1773);
nor U3207 (N_3207,N_646,N_2500);
and U3208 (N_3208,N_1129,N_2360);
and U3209 (N_3209,N_1717,N_2687);
nor U3210 (N_3210,N_701,N_1999);
xnor U3211 (N_3211,N_2975,N_974);
or U3212 (N_3212,N_2258,N_2232);
nand U3213 (N_3213,N_2816,N_490);
or U3214 (N_3214,N_218,N_2044);
nand U3215 (N_3215,N_852,N_2135);
xnor U3216 (N_3216,N_1516,N_986);
xnor U3217 (N_3217,N_1626,N_1840);
xor U3218 (N_3218,N_1322,N_312);
nand U3219 (N_3219,N_1350,N_2917);
and U3220 (N_3220,N_691,N_508);
and U3221 (N_3221,N_861,N_1349);
nand U3222 (N_3222,N_112,N_2838);
or U3223 (N_3223,N_752,N_1306);
or U3224 (N_3224,N_306,N_1605);
nand U3225 (N_3225,N_1656,N_2104);
or U3226 (N_3226,N_2408,N_712);
or U3227 (N_3227,N_2095,N_1674);
or U3228 (N_3228,N_764,N_2740);
or U3229 (N_3229,N_266,N_1110);
and U3230 (N_3230,N_1633,N_896);
and U3231 (N_3231,N_2508,N_2863);
nor U3232 (N_3232,N_2514,N_2930);
or U3233 (N_3233,N_818,N_1074);
and U3234 (N_3234,N_1273,N_2573);
or U3235 (N_3235,N_227,N_2578);
nor U3236 (N_3236,N_2856,N_612);
and U3237 (N_3237,N_2755,N_1896);
nand U3238 (N_3238,N_1206,N_1743);
nand U3239 (N_3239,N_2550,N_1776);
xor U3240 (N_3240,N_897,N_2719);
and U3241 (N_3241,N_2841,N_2592);
and U3242 (N_3242,N_1634,N_1059);
nor U3243 (N_3243,N_420,N_2642);
nand U3244 (N_3244,N_1282,N_1472);
and U3245 (N_3245,N_2471,N_1499);
or U3246 (N_3246,N_2832,N_703);
nor U3247 (N_3247,N_487,N_1648);
nor U3248 (N_3248,N_383,N_1264);
xnor U3249 (N_3249,N_713,N_1995);
nand U3250 (N_3250,N_1439,N_2134);
nor U3251 (N_3251,N_584,N_1877);
nor U3252 (N_3252,N_267,N_2748);
or U3253 (N_3253,N_882,N_2478);
and U3254 (N_3254,N_553,N_2892);
nand U3255 (N_3255,N_2432,N_601);
and U3256 (N_3256,N_846,N_2593);
or U3257 (N_3257,N_789,N_351);
nand U3258 (N_3258,N_2276,N_2720);
nor U3259 (N_3259,N_2585,N_693);
nor U3260 (N_3260,N_2810,N_1380);
and U3261 (N_3261,N_1297,N_2094);
or U3262 (N_3262,N_1809,N_44);
or U3263 (N_3263,N_419,N_1377);
or U3264 (N_3264,N_1241,N_1004);
or U3265 (N_3265,N_1238,N_2428);
and U3266 (N_3266,N_2055,N_1192);
or U3267 (N_3267,N_2551,N_1890);
nor U3268 (N_3268,N_2228,N_1604);
nand U3269 (N_3269,N_1707,N_2317);
nand U3270 (N_3270,N_1777,N_140);
nor U3271 (N_3271,N_1957,N_369);
nand U3272 (N_3272,N_2977,N_1894);
xor U3273 (N_3273,N_1974,N_2767);
nand U3274 (N_3274,N_739,N_1695);
nand U3275 (N_3275,N_1630,N_2441);
or U3276 (N_3276,N_1166,N_763);
nand U3277 (N_3277,N_794,N_2881);
nand U3278 (N_3278,N_2823,N_2244);
nor U3279 (N_3279,N_298,N_432);
nor U3280 (N_3280,N_2162,N_2350);
or U3281 (N_3281,N_1222,N_1846);
or U3282 (N_3282,N_1276,N_1603);
or U3283 (N_3283,N_2927,N_1885);
xor U3284 (N_3284,N_2026,N_792);
or U3285 (N_3285,N_1389,N_738);
or U3286 (N_3286,N_107,N_2698);
or U3287 (N_3287,N_1851,N_66);
nand U3288 (N_3288,N_880,N_2009);
or U3289 (N_3289,N_2668,N_136);
nor U3290 (N_3290,N_217,N_700);
xor U3291 (N_3291,N_629,N_1645);
nand U3292 (N_3292,N_2312,N_2973);
nor U3293 (N_3293,N_2760,N_1577);
nor U3294 (N_3294,N_2959,N_926);
nand U3295 (N_3295,N_1738,N_1888);
or U3296 (N_3296,N_2467,N_1003);
and U3297 (N_3297,N_2877,N_1671);
or U3298 (N_3298,N_2583,N_343);
nor U3299 (N_3299,N_169,N_2159);
or U3300 (N_3300,N_2995,N_165);
nor U3301 (N_3301,N_2865,N_2498);
and U3302 (N_3302,N_1933,N_1608);
nand U3303 (N_3303,N_1223,N_2230);
nand U3304 (N_3304,N_771,N_2958);
nand U3305 (N_3305,N_22,N_1943);
nand U3306 (N_3306,N_2676,N_2293);
and U3307 (N_3307,N_514,N_2542);
or U3308 (N_3308,N_65,N_1649);
nand U3309 (N_3309,N_195,N_2695);
or U3310 (N_3310,N_719,N_2682);
nor U3311 (N_3311,N_326,N_1298);
or U3312 (N_3312,N_491,N_2000);
nor U3313 (N_3313,N_647,N_709);
and U3314 (N_3314,N_2462,N_2181);
xor U3315 (N_3315,N_1652,N_55);
or U3316 (N_3316,N_139,N_1798);
and U3317 (N_3317,N_536,N_1169);
or U3318 (N_3318,N_173,N_202);
xor U3319 (N_3319,N_207,N_1997);
and U3320 (N_3320,N_945,N_231);
nand U3321 (N_3321,N_602,N_292);
nand U3322 (N_3322,N_1765,N_154);
nor U3323 (N_3323,N_2937,N_616);
nor U3324 (N_3324,N_2997,N_831);
xnor U3325 (N_3325,N_1469,N_2739);
nor U3326 (N_3326,N_2021,N_440);
nor U3327 (N_3327,N_1536,N_31);
and U3328 (N_3328,N_594,N_2051);
or U3329 (N_3329,N_120,N_391);
nor U3330 (N_3330,N_489,N_1225);
nand U3331 (N_3331,N_916,N_101);
and U3332 (N_3332,N_1396,N_2488);
nor U3333 (N_3333,N_2928,N_515);
and U3334 (N_3334,N_1842,N_371);
or U3335 (N_3335,N_2252,N_1657);
or U3336 (N_3336,N_714,N_2947);
nand U3337 (N_3337,N_1736,N_521);
nand U3338 (N_3338,N_2700,N_907);
nand U3339 (N_3339,N_2979,N_1330);
and U3340 (N_3340,N_1787,N_309);
xnor U3341 (N_3341,N_1267,N_1219);
nor U3342 (N_3342,N_1752,N_441);
and U3343 (N_3343,N_505,N_1095);
or U3344 (N_3344,N_2153,N_1445);
or U3345 (N_3345,N_2089,N_507);
xor U3346 (N_3346,N_776,N_1087);
or U3347 (N_3347,N_1249,N_152);
nor U3348 (N_3348,N_2510,N_2056);
nand U3349 (N_3349,N_1589,N_2801);
nor U3350 (N_3350,N_573,N_1715);
nor U3351 (N_3351,N_1475,N_147);
nor U3352 (N_3352,N_2812,N_2029);
nor U3353 (N_3353,N_2256,N_149);
or U3354 (N_3354,N_1363,N_421);
or U3355 (N_3355,N_994,N_1);
nor U3356 (N_3356,N_1425,N_598);
nor U3357 (N_3357,N_206,N_2869);
nand U3358 (N_3358,N_2229,N_1931);
and U3359 (N_3359,N_2983,N_1555);
nand U3360 (N_3360,N_981,N_1484);
nor U3361 (N_3361,N_1399,N_2078);
or U3362 (N_3362,N_539,N_942);
and U3363 (N_3363,N_2424,N_2169);
nand U3364 (N_3364,N_595,N_2886);
and U3365 (N_3365,N_1669,N_1376);
and U3366 (N_3366,N_809,N_2582);
nor U3367 (N_3367,N_731,N_1618);
and U3368 (N_3368,N_318,N_1963);
nand U3369 (N_3369,N_2407,N_2362);
nor U3370 (N_3370,N_46,N_1268);
xor U3371 (N_3371,N_1146,N_2743);
nor U3372 (N_3372,N_1226,N_1573);
nand U3373 (N_3373,N_2161,N_470);
nand U3374 (N_3374,N_2821,N_1014);
or U3375 (N_3375,N_2012,N_879);
and U3376 (N_3376,N_1742,N_2297);
or U3377 (N_3377,N_2913,N_1415);
or U3378 (N_3378,N_1892,N_2775);
and U3379 (N_3379,N_1968,N_802);
and U3380 (N_3380,N_1390,N_2532);
and U3381 (N_3381,N_1788,N_1320);
or U3382 (N_3382,N_597,N_2537);
nand U3383 (N_3383,N_1262,N_1187);
nor U3384 (N_3384,N_1947,N_791);
nand U3385 (N_3385,N_30,N_137);
and U3386 (N_3386,N_1147,N_1005);
and U3387 (N_3387,N_1111,N_2879);
or U3388 (N_3388,N_134,N_1461);
and U3389 (N_3389,N_1127,N_1598);
nor U3390 (N_3390,N_1006,N_2348);
or U3391 (N_3391,N_2262,N_162);
and U3392 (N_3392,N_1675,N_2620);
nor U3393 (N_3393,N_2789,N_828);
or U3394 (N_3394,N_1139,N_411);
nand U3395 (N_3395,N_624,N_2434);
nor U3396 (N_3396,N_2184,N_1857);
nand U3397 (N_3397,N_428,N_1878);
and U3398 (N_3398,N_2076,N_424);
nand U3399 (N_3399,N_17,N_1635);
nor U3400 (N_3400,N_1911,N_2289);
or U3401 (N_3401,N_511,N_2672);
and U3402 (N_3402,N_917,N_1451);
nor U3403 (N_3403,N_2603,N_912);
nand U3404 (N_3404,N_962,N_867);
and U3405 (N_3405,N_429,N_2002);
nor U3406 (N_3406,N_759,N_1607);
xor U3407 (N_3407,N_1220,N_1647);
xnor U3408 (N_3408,N_2705,N_1534);
or U3409 (N_3409,N_15,N_1981);
nor U3410 (N_3410,N_2448,N_1755);
xnor U3411 (N_3411,N_1413,N_2961);
or U3412 (N_3412,N_478,N_2986);
and U3413 (N_3413,N_2939,N_2876);
nand U3414 (N_3414,N_2242,N_870);
nor U3415 (N_3415,N_2309,N_1265);
and U3416 (N_3416,N_1452,N_732);
nand U3417 (N_3417,N_1984,N_1960);
or U3418 (N_3418,N_1895,N_1200);
and U3419 (N_3419,N_2302,N_581);
nor U3420 (N_3420,N_444,N_405);
xor U3421 (N_3421,N_2300,N_1875);
and U3422 (N_3422,N_944,N_2851);
nand U3423 (N_3423,N_1724,N_2069);
and U3424 (N_3424,N_678,N_2479);
and U3425 (N_3425,N_2105,N_2644);
and U3426 (N_3426,N_2962,N_2691);
or U3427 (N_3427,N_70,N_1279);
or U3428 (N_3428,N_1889,N_1148);
and U3429 (N_3429,N_1786,N_456);
xor U3430 (N_3430,N_2048,N_78);
and U3431 (N_3431,N_1342,N_891);
or U3432 (N_3432,N_2059,N_1258);
nor U3433 (N_3433,N_1898,N_2343);
and U3434 (N_3434,N_2087,N_368);
xnor U3435 (N_3435,N_1692,N_1728);
nor U3436 (N_3436,N_2113,N_1791);
and U3437 (N_3437,N_2492,N_1131);
and U3438 (N_3438,N_1357,N_118);
and U3439 (N_3439,N_567,N_2319);
nor U3440 (N_3440,N_2182,N_2880);
nor U3441 (N_3441,N_849,N_2716);
and U3442 (N_3442,N_1274,N_1956);
xor U3443 (N_3443,N_2867,N_1572);
nand U3444 (N_3444,N_1606,N_407);
xor U3445 (N_3445,N_2304,N_2447);
nor U3446 (N_3446,N_1821,N_997);
and U3447 (N_3447,N_817,N_928);
xor U3448 (N_3448,N_1880,N_117);
nand U3449 (N_3449,N_2747,N_943);
nand U3450 (N_3450,N_2144,N_830);
nor U3451 (N_3451,N_360,N_2364);
xor U3452 (N_3452,N_574,N_1218);
or U3453 (N_3453,N_303,N_1244);
nor U3454 (N_3454,N_1660,N_2756);
nand U3455 (N_3455,N_108,N_1245);
and U3456 (N_3456,N_2233,N_300);
or U3457 (N_3457,N_642,N_1073);
nand U3458 (N_3458,N_2998,N_422);
or U3459 (N_3459,N_684,N_2173);
xnor U3460 (N_3460,N_668,N_433);
nand U3461 (N_3461,N_999,N_2049);
nor U3462 (N_3462,N_845,N_2384);
nand U3463 (N_3463,N_617,N_2629);
and U3464 (N_3464,N_1559,N_1881);
or U3465 (N_3465,N_1723,N_1827);
nor U3466 (N_3466,N_1848,N_463);
or U3467 (N_3467,N_2534,N_2045);
and U3468 (N_3468,N_2223,N_180);
and U3469 (N_3469,N_615,N_1162);
xnor U3470 (N_3470,N_2320,N_2465);
or U3471 (N_3471,N_546,N_1061);
or U3472 (N_3472,N_2753,N_2143);
or U3473 (N_3473,N_1012,N_2664);
nor U3474 (N_3474,N_164,N_881);
and U3475 (N_3475,N_1368,N_1702);
or U3476 (N_3476,N_2699,N_414);
or U3477 (N_3477,N_1101,N_2502);
nor U3478 (N_3478,N_1374,N_1526);
and U3479 (N_3479,N_756,N_753);
nor U3480 (N_3480,N_49,N_1959);
and U3481 (N_3481,N_1124,N_110);
and U3482 (N_3482,N_2938,N_1980);
nand U3483 (N_3483,N_924,N_2745);
nand U3484 (N_3484,N_248,N_2204);
xor U3485 (N_3485,N_969,N_1735);
nor U3486 (N_3486,N_733,N_1115);
and U3487 (N_3487,N_1233,N_2952);
xnor U3488 (N_3488,N_1203,N_2476);
nand U3489 (N_3489,N_2531,N_2065);
nor U3490 (N_3490,N_43,N_1570);
or U3491 (N_3491,N_2061,N_2209);
nand U3492 (N_3492,N_235,N_2646);
xnor U3493 (N_3493,N_710,N_2561);
or U3494 (N_3494,N_125,N_1492);
or U3495 (N_3495,N_2540,N_834);
or U3496 (N_3496,N_2526,N_2390);
nand U3497 (N_3497,N_280,N_1479);
or U3498 (N_3498,N_1055,N_779);
and U3499 (N_3499,N_2190,N_932);
and U3500 (N_3500,N_596,N_2539);
nand U3501 (N_3501,N_1161,N_2310);
xor U3502 (N_3502,N_2299,N_1199);
xnor U3503 (N_3503,N_2452,N_2265);
and U3504 (N_3504,N_282,N_1811);
xnor U3505 (N_3505,N_209,N_1034);
and U3506 (N_3506,N_2982,N_2053);
nor U3507 (N_3507,N_1949,N_840);
and U3508 (N_3508,N_2831,N_1581);
and U3509 (N_3509,N_1272,N_274);
or U3510 (N_3510,N_2904,N_1309);
and U3511 (N_3511,N_1954,N_1072);
and U3512 (N_3512,N_755,N_664);
xnor U3513 (N_3513,N_1339,N_2475);
nor U3514 (N_3514,N_2595,N_1263);
or U3515 (N_3515,N_2762,N_718);
nand U3516 (N_3516,N_57,N_532);
and U3517 (N_3517,N_1457,N_450);
or U3518 (N_3518,N_2079,N_922);
nand U3519 (N_3519,N_1822,N_1293);
nor U3520 (N_3520,N_2346,N_461);
nor U3521 (N_3521,N_2387,N_2318);
nand U3522 (N_3522,N_1625,N_452);
nor U3523 (N_3523,N_189,N_529);
and U3524 (N_3524,N_2422,N_1315);
nor U3525 (N_3525,N_1270,N_400);
or U3526 (N_3526,N_2198,N_872);
or U3527 (N_3527,N_1523,N_447);
xnor U3528 (N_3528,N_2931,N_665);
nand U3529 (N_3529,N_2118,N_1590);
or U3530 (N_3530,N_135,N_2688);
and U3531 (N_3531,N_2547,N_2520);
nor U3532 (N_3532,N_1833,N_769);
xnor U3533 (N_3533,N_1818,N_2680);
nor U3534 (N_3534,N_2410,N_446);
or U3535 (N_3535,N_2849,N_144);
nand U3536 (N_3536,N_1428,N_2623);
and U3537 (N_3537,N_2170,N_2734);
or U3538 (N_3538,N_1790,N_1566);
or U3539 (N_3539,N_1303,N_2213);
nor U3540 (N_3540,N_373,N_498);
nor U3541 (N_3541,N_14,N_1501);
and U3542 (N_3542,N_2925,N_1171);
or U3543 (N_3543,N_2670,N_2280);
or U3544 (N_3544,N_2468,N_249);
nand U3545 (N_3545,N_1504,N_1722);
or U3546 (N_3546,N_468,N_613);
or U3547 (N_3547,N_2174,N_2976);
nor U3548 (N_3548,N_1117,N_1521);
nand U3549 (N_3549,N_1568,N_2945);
nor U3550 (N_3550,N_2336,N_2709);
nand U3551 (N_3551,N_2536,N_1392);
or U3552 (N_3552,N_2096,N_197);
nand U3553 (N_3553,N_1835,N_1527);
and U3554 (N_3554,N_1214,N_793);
or U3555 (N_3555,N_2638,N_389);
and U3556 (N_3556,N_1955,N_1906);
nand U3557 (N_3557,N_1204,N_1278);
nor U3558 (N_3558,N_132,N_2140);
xnor U3559 (N_3559,N_971,N_2889);
nor U3560 (N_3560,N_1337,N_485);
nand U3561 (N_3561,N_2896,N_367);
or U3562 (N_3562,N_1921,N_650);
nand U3563 (N_3563,N_711,N_1793);
nor U3564 (N_3564,N_2660,N_296);
and U3565 (N_3565,N_641,N_1522);
nor U3566 (N_3566,N_254,N_375);
xor U3567 (N_3567,N_653,N_1000);
nor U3568 (N_3568,N_854,N_2655);
and U3569 (N_3569,N_2314,N_1760);
nand U3570 (N_3570,N_337,N_86);
nor U3571 (N_3571,N_2763,N_2989);
nor U3572 (N_3572,N_705,N_2247);
nand U3573 (N_3573,N_2912,N_263);
nand U3574 (N_3574,N_2843,N_9);
or U3575 (N_3575,N_2110,N_460);
and U3576 (N_3576,N_2967,N_2586);
nand U3577 (N_3577,N_1930,N_1832);
nand U3578 (N_3578,N_1801,N_2964);
nor U3579 (N_3579,N_1186,N_785);
nor U3580 (N_3580,N_1664,N_2388);
nor U3581 (N_3581,N_811,N_2406);
nand U3582 (N_3582,N_352,N_2667);
and U3583 (N_3583,N_2298,N_346);
and U3584 (N_3584,N_2957,N_503);
nor U3585 (N_3585,N_216,N_374);
nand U3586 (N_3586,N_2007,N_947);
nand U3587 (N_3587,N_1386,N_946);
xnor U3588 (N_3588,N_2111,N_1477);
xnor U3589 (N_3589,N_2610,N_2018);
nand U3590 (N_3590,N_1700,N_1740);
or U3591 (N_3591,N_2575,N_569);
and U3592 (N_3592,N_2329,N_2893);
or U3593 (N_3593,N_2914,N_925);
or U3594 (N_3594,N_471,N_1182);
nor U3595 (N_3595,N_1749,N_1797);
xor U3596 (N_3596,N_2392,N_307);
and U3597 (N_3597,N_1116,N_1067);
or U3598 (N_3598,N_2259,N_2933);
or U3599 (N_3599,N_1173,N_1287);
nand U3600 (N_3600,N_2588,N_1541);
or U3601 (N_3601,N_826,N_2685);
nor U3602 (N_3602,N_741,N_1412);
and U3603 (N_3603,N_2919,N_554);
xor U3604 (N_3604,N_620,N_913);
or U3605 (N_3605,N_1558,N_10);
or U3606 (N_3606,N_2850,N_1926);
nand U3607 (N_3607,N_1296,N_1017);
xnor U3608 (N_3608,N_2126,N_1518);
nor U3609 (N_3609,N_2160,N_275);
nand U3610 (N_3610,N_600,N_1077);
and U3611 (N_3611,N_1462,N_2953);
nor U3612 (N_3612,N_361,N_1311);
nand U3613 (N_3613,N_1348,N_2356);
and U3614 (N_3614,N_32,N_1294);
nor U3615 (N_3615,N_2712,N_2523);
or U3616 (N_3616,N_2773,N_2477);
nand U3617 (N_3617,N_513,N_1178);
nand U3618 (N_3618,N_500,N_2439);
or U3619 (N_3619,N_582,N_1237);
nor U3620 (N_3620,N_2799,N_1579);
nor U3621 (N_3621,N_1197,N_1737);
xnor U3622 (N_3622,N_2808,N_1524);
nand U3623 (N_3623,N_2663,N_295);
or U3624 (N_3624,N_1359,N_2794);
or U3625 (N_3625,N_2139,N_1562);
or U3626 (N_3626,N_2758,N_2058);
xnor U3627 (N_3627,N_2559,N_2435);
or U3628 (N_3628,N_607,N_176);
and U3629 (N_3629,N_2417,N_1048);
nand U3630 (N_3630,N_2257,N_220);
and U3631 (N_3631,N_1181,N_2622);
nand U3632 (N_3632,N_836,N_2219);
or U3633 (N_3633,N_2385,N_1043);
nand U3634 (N_3634,N_1435,N_2458);
nor U3635 (N_3635,N_2771,N_708);
and U3636 (N_3636,N_2496,N_1411);
and U3637 (N_3637,N_146,N_2423);
and U3638 (N_3638,N_2440,N_1213);
or U3639 (N_3639,N_1158,N_1358);
and U3640 (N_3640,N_2809,N_438);
nor U3641 (N_3641,N_2436,N_2777);
and U3642 (N_3642,N_1403,N_1686);
nor U3643 (N_3643,N_2131,N_2834);
nor U3644 (N_3644,N_344,N_931);
and U3645 (N_3645,N_1597,N_1714);
or U3646 (N_3646,N_2764,N_1919);
or U3647 (N_3647,N_2567,N_1644);
nor U3648 (N_3648,N_2196,N_1112);
and U3649 (N_3649,N_2226,N_69);
nand U3650 (N_3650,N_1886,N_2571);
xor U3651 (N_3651,N_1718,N_1130);
or U3652 (N_3652,N_2286,N_1525);
nor U3653 (N_3653,N_814,N_224);
xnor U3654 (N_3654,N_2449,N_1196);
nor U3655 (N_3655,N_475,N_80);
or U3656 (N_3656,N_676,N_630);
nand U3657 (N_3657,N_1308,N_504);
and U3658 (N_3658,N_2565,N_1395);
or U3659 (N_3659,N_2991,N_1334);
or U3660 (N_3660,N_305,N_545);
and U3661 (N_3661,N_2884,N_1295);
nand U3662 (N_3662,N_38,N_123);
nand U3663 (N_3663,N_2191,N_1642);
nand U3664 (N_3664,N_1862,N_2032);
and U3665 (N_3665,N_2323,N_2083);
nor U3666 (N_3666,N_2331,N_914);
and U3667 (N_3667,N_2224,N_2941);
nand U3668 (N_3668,N_2948,N_2250);
and U3669 (N_3669,N_1332,N_1436);
nor U3670 (N_3670,N_1551,N_1805);
nor U3671 (N_3671,N_512,N_1601);
and U3672 (N_3672,N_394,N_1438);
xor U3673 (N_3673,N_1104,N_766);
and U3674 (N_3674,N_24,N_1064);
nor U3675 (N_3675,N_2120,N_90);
xnor U3676 (N_3676,N_716,N_2367);
and U3677 (N_3677,N_1232,N_2311);
nand U3678 (N_3678,N_2600,N_2090);
and U3679 (N_3679,N_2992,N_2121);
and U3680 (N_3680,N_2954,N_1316);
and U3681 (N_3681,N_1331,N_319);
nand U3682 (N_3682,N_435,N_1165);
and U3683 (N_3683,N_2845,N_832);
nand U3684 (N_3684,N_1964,N_2461);
nand U3685 (N_3685,N_320,N_1946);
nand U3686 (N_3686,N_1335,N_1082);
nor U3687 (N_3687,N_1935,N_1168);
and U3688 (N_3688,N_2063,N_2708);
nor U3689 (N_3689,N_1378,N_1253);
nand U3690 (N_3690,N_434,N_1027);
nor U3691 (N_3691,N_2335,N_2231);
or U3692 (N_3692,N_2741,N_643);
nor U3693 (N_3693,N_1932,N_1661);
nand U3694 (N_3694,N_2107,N_1108);
nand U3695 (N_3695,N_663,N_467);
xor U3696 (N_3696,N_2815,N_1704);
xor U3697 (N_3697,N_2506,N_2754);
and U3698 (N_3698,N_2141,N_2491);
and U3699 (N_3699,N_704,N_1247);
xor U3700 (N_3700,N_2996,N_1090);
or U3701 (N_3701,N_1754,N_2180);
nand U3702 (N_3702,N_2751,N_1563);
nand U3703 (N_3703,N_599,N_1585);
nand U3704 (N_3704,N_906,N_2909);
nand U3705 (N_3705,N_590,N_790);
nor U3706 (N_3706,N_2490,N_679);
nand U3707 (N_3707,N_2955,N_1125);
xnor U3708 (N_3708,N_1410,N_2464);
and U3709 (N_3709,N_1744,N_815);
nor U3710 (N_3710,N_39,N_2272);
nor U3711 (N_3711,N_649,N_1815);
and U3712 (N_3712,N_2339,N_449);
and U3713 (N_3713,N_1140,N_2530);
nor U3714 (N_3714,N_160,N_801);
or U3715 (N_3715,N_1986,N_1680);
or U3716 (N_3716,N_439,N_2188);
nor U3717 (N_3717,N_2192,N_2891);
or U3718 (N_3718,N_1670,N_476);
nor U3719 (N_3719,N_1154,N_2899);
nor U3720 (N_3720,N_1235,N_1632);
nor U3721 (N_3721,N_1817,N_2085);
nand U3722 (N_3722,N_2966,N_2022);
and U3723 (N_3723,N_2119,N_1716);
nor U3724 (N_3724,N_1400,N_2101);
nand U3725 (N_3725,N_321,N_2802);
or U3726 (N_3726,N_729,N_2214);
or U3727 (N_3727,N_155,N_2750);
nand U3728 (N_3728,N_2400,N_2940);
and U3729 (N_3729,N_1698,N_247);
xor U3730 (N_3730,N_1347,N_453);
and U3731 (N_3731,N_901,N_2395);
nor U3732 (N_3732,N_1741,N_2728);
nor U3733 (N_3733,N_2112,N_417);
nor U3734 (N_3734,N_1246,N_1640);
nor U3735 (N_3735,N_2718,N_2267);
nor U3736 (N_3736,N_855,N_1992);
nand U3737 (N_3737,N_1612,N_2372);
and U3738 (N_3738,N_2507,N_509);
nand U3739 (N_3739,N_1828,N_109);
nor U3740 (N_3740,N_148,N_1070);
nand U3741 (N_3741,N_1592,N_1611);
or U3742 (N_3742,N_2661,N_457);
or U3743 (N_3743,N_2731,N_1825);
or U3744 (N_3744,N_2669,N_2199);
and U3745 (N_3745,N_2270,N_12);
and U3746 (N_3746,N_258,N_2227);
and U3747 (N_3747,N_1532,N_242);
and U3748 (N_3748,N_2974,N_530);
xnor U3749 (N_3749,N_696,N_1925);
nor U3750 (N_3750,N_1912,N_1701);
nand U3751 (N_3751,N_1370,N_1201);
nor U3752 (N_3752,N_2594,N_83);
nor U3753 (N_3753,N_2606,N_1934);
and U3754 (N_3754,N_2445,N_805);
and U3755 (N_3755,N_551,N_2084);
xnor U3756 (N_3756,N_1429,N_2662);
nor U3757 (N_3757,N_2800,N_2853);
and U3758 (N_3758,N_2456,N_1160);
or U3759 (N_3759,N_2901,N_1792);
or U3760 (N_3760,N_2942,N_56);
or U3761 (N_3761,N_2584,N_2030);
or U3762 (N_3762,N_2929,N_387);
or U3763 (N_3763,N_869,N_1685);
and U3764 (N_3764,N_1750,N_2612);
or U3765 (N_3765,N_877,N_1993);
nor U3766 (N_3766,N_2737,N_1202);
nand U3767 (N_3767,N_1989,N_1520);
and U3768 (N_3768,N_1802,N_2721);
nand U3769 (N_3769,N_634,N_883);
or U3770 (N_3770,N_99,N_2151);
nor U3771 (N_3771,N_1679,N_2553);
nand U3772 (N_3772,N_1766,N_798);
and U3773 (N_3773,N_2046,N_246);
nand U3774 (N_3774,N_1317,N_1234);
and U3775 (N_3775,N_674,N_578);
nor U3776 (N_3776,N_547,N_717);
nand U3777 (N_3777,N_133,N_1387);
and U3778 (N_3778,N_2627,N_1624);
or U3779 (N_3779,N_823,N_502);
xnor U3780 (N_3780,N_53,N_1511);
and U3781 (N_3781,N_1505,N_2790);
nor U3782 (N_3782,N_2186,N_2443);
nor U3783 (N_3783,N_570,N_158);
and U3784 (N_3784,N_730,N_2971);
and U3785 (N_3785,N_1891,N_892);
or U3786 (N_3786,N_2527,N_1157);
or U3787 (N_3787,N_1421,N_1052);
nor U3788 (N_3788,N_2035,N_2597);
nand U3789 (N_3789,N_561,N_1859);
xnor U3790 (N_3790,N_363,N_2128);
nand U3791 (N_3791,N_130,N_2365);
nand U3792 (N_3792,N_672,N_2855);
or U3793 (N_3793,N_2787,N_1024);
nor U3794 (N_3794,N_833,N_2166);
and U3795 (N_3795,N_658,N_2780);
nor U3796 (N_3796,N_1217,N_2001);
and U3797 (N_3797,N_2854,N_2568);
nand U3798 (N_3798,N_745,N_1453);
or U3799 (N_3799,N_1732,N_384);
nor U3800 (N_3800,N_2779,N_984);
nand U3801 (N_3801,N_284,N_1560);
and U3802 (N_3802,N_2383,N_2766);
nor U3803 (N_3803,N_1803,N_1965);
or U3804 (N_3804,N_2117,N_1939);
nand U3805 (N_3805,N_1561,N_951);
nand U3806 (N_3806,N_354,N_1506);
and U3807 (N_3807,N_2016,N_878);
nor U3808 (N_3808,N_483,N_2828);
or U3809 (N_3809,N_304,N_1096);
nand U3810 (N_3810,N_163,N_2481);
and U3811 (N_3811,N_200,N_2338);
nand U3812 (N_3812,N_2431,N_1571);
and U3813 (N_3813,N_810,N_2202);
nor U3814 (N_3814,N_287,N_237);
nand U3815 (N_3815,N_2357,N_1883);
and U3816 (N_3816,N_1733,N_2653);
nor U3817 (N_3817,N_1069,N_2846);
nand U3818 (N_3818,N_401,N_1304);
or U3819 (N_3819,N_329,N_2999);
nor U3820 (N_3820,N_1567,N_297);
nand U3821 (N_3821,N_1667,N_1998);
or U3822 (N_3822,N_681,N_1150);
nand U3823 (N_3823,N_156,N_2489);
nor U3824 (N_3824,N_842,N_1650);
and U3825 (N_3825,N_1975,N_106);
xor U3826 (N_3826,N_1152,N_153);
and U3827 (N_3827,N_265,N_903);
nor U3828 (N_3828,N_2848,N_1734);
nand U3829 (N_3829,N_2480,N_1427);
nor U3830 (N_3830,N_2482,N_2702);
or U3831 (N_3831,N_166,N_1300);
and U3832 (N_3832,N_2207,N_2017);
and U3833 (N_3833,N_2878,N_2450);
nand U3834 (N_3834,N_182,N_965);
and U3835 (N_3835,N_638,N_2710);
or U3836 (N_3836,N_119,N_1546);
and U3837 (N_3837,N_1078,N_2386);
nor U3838 (N_3838,N_2414,N_1900);
nand U3839 (N_3839,N_1195,N_2538);
and U3840 (N_3840,N_2618,N_492);
or U3841 (N_3841,N_2091,N_1163);
nor U3842 (N_3842,N_2611,N_1318);
nand U3843 (N_3843,N_2533,N_2237);
nor U3844 (N_3844,N_2645,N_1483);
xnor U3845 (N_3845,N_1464,N_2949);
nor U3846 (N_3846,N_621,N_2014);
and U3847 (N_3847,N_2261,N_930);
xor U3848 (N_3848,N_1210,N_2249);
or U3849 (N_3849,N_2935,N_129);
nand U3850 (N_3850,N_1351,N_819);
and U3851 (N_3851,N_2254,N_2742);
nand U3852 (N_3852,N_1971,N_1010);
or U3853 (N_3853,N_362,N_2375);
nand U3854 (N_3854,N_1489,N_963);
or U3855 (N_3855,N_2150,N_534);
or U3856 (N_3856,N_2677,N_1016);
or U3857 (N_3857,N_74,N_632);
nand U3858 (N_3858,N_1402,N_150);
nor U3859 (N_3859,N_2405,N_1441);
nor U3860 (N_3860,N_1207,N_2326);
xnor U3861 (N_3861,N_1996,N_2429);
or U3862 (N_3862,N_1385,N_1812);
nor U3863 (N_3863,N_1193,N_1177);
nor U3864 (N_3864,N_2403,N_637);
and U3865 (N_3865,N_323,N_1599);
xor U3866 (N_3866,N_604,N_2549);
and U3867 (N_3867,N_2201,N_480);
xor U3868 (N_3868,N_559,N_2156);
and U3869 (N_3869,N_1967,N_1151);
and U3870 (N_3870,N_302,N_87);
nor U3871 (N_3871,N_1449,N_692);
or U3872 (N_3872,N_1431,N_1973);
nor U3873 (N_3873,N_2082,N_1868);
and U3874 (N_3874,N_157,N_1432);
nand U3875 (N_3875,N_213,N_290);
nand U3876 (N_3876,N_2943,N_2988);
nand U3877 (N_3877,N_856,N_816);
nand U3878 (N_3878,N_193,N_365);
nor U3879 (N_3879,N_1283,N_938);
xor U3880 (N_3880,N_2460,N_1837);
nand U3881 (N_3881,N_754,N_2011);
nor U3882 (N_3882,N_2455,N_1228);
or U3883 (N_3883,N_765,N_538);
nand U3884 (N_3884,N_1011,N_1613);
nor U3885 (N_3885,N_2033,N_315);
nand U3886 (N_3886,N_586,N_2145);
nor U3887 (N_3887,N_425,N_474);
nor U3888 (N_3888,N_2132,N_2725);
or U3889 (N_3889,N_1212,N_2179);
and U3890 (N_3890,N_948,N_1194);
xor U3891 (N_3891,N_1705,N_2840);
nand U3892 (N_3892,N_1682,N_2722);
and U3893 (N_3893,N_2495,N_1216);
nand U3894 (N_3894,N_2418,N_168);
nand U3895 (N_3895,N_2903,N_2835);
or U3896 (N_3896,N_141,N_1902);
or U3897 (N_3897,N_1711,N_1870);
and U3898 (N_3898,N_1953,N_2784);
or U3899 (N_3899,N_772,N_2825);
nand U3900 (N_3900,N_1040,N_550);
nor U3901 (N_3901,N_2003,N_2738);
nand U3902 (N_3902,N_2351,N_706);
or U3903 (N_3903,N_813,N_957);
and U3904 (N_3904,N_1867,N_2637);
and U3905 (N_3905,N_2274,N_1155);
nand U3906 (N_3906,N_2844,N_273);
and U3907 (N_3907,N_2788,N_2454);
or U3908 (N_3908,N_743,N_2352);
xnor U3909 (N_3909,N_579,N_1135);
and U3910 (N_3910,N_2736,N_2278);
and U3911 (N_3911,N_572,N_2656);
nand U3912 (N_3912,N_1582,N_2);
or U3913 (N_3913,N_1575,N_2864);
or U3914 (N_3914,N_698,N_338);
or U3915 (N_3915,N_808,N_2349);
and U3916 (N_3916,N_2081,N_953);
xnor U3917 (N_3917,N_1463,N_1373);
nor U3918 (N_3918,N_21,N_1257);
nor U3919 (N_3919,N_1136,N_1513);
or U3920 (N_3920,N_524,N_2872);
nor U3921 (N_3921,N_2281,N_223);
nor U3922 (N_3922,N_2666,N_336);
and U3923 (N_3923,N_1369,N_1394);
nor U3924 (N_3924,N_410,N_2366);
nor U3925 (N_3925,N_2715,N_464);
xnor U3926 (N_3926,N_2401,N_1627);
xnor U3927 (N_3927,N_2067,N_1126);
nand U3928 (N_3928,N_2036,N_2006);
nor U3929 (N_3929,N_2074,N_633);
nand U3930 (N_3930,N_2696,N_2240);
and U3931 (N_3931,N_1259,N_885);
or U3932 (N_3932,N_1031,N_2757);
and U3933 (N_3933,N_1772,N_1548);
and U3934 (N_3934,N_2501,N_835);
nor U3935 (N_3935,N_960,N_50);
nor U3936 (N_3936,N_1448,N_1987);
nor U3937 (N_3937,N_1029,N_848);
nor U3938 (N_3938,N_1379,N_1356);
or U3939 (N_3939,N_2970,N_1580);
or U3940 (N_3940,N_2723,N_657);
or U3941 (N_3941,N_1950,N_1198);
nor U3942 (N_3942,N_2525,N_1540);
or U3943 (N_3943,N_2474,N_727);
nor U3944 (N_3944,N_1528,N_2420);
or U3945 (N_3945,N_1255,N_1569);
and U3946 (N_3946,N_2427,N_1583);
nor U3947 (N_3947,N_1084,N_2382);
nor U3948 (N_3948,N_325,N_1076);
nand U3949 (N_3949,N_2187,N_1191);
and U3950 (N_3950,N_2774,N_1493);
nand U3951 (N_3951,N_1153,N_1869);
and U3952 (N_3952,N_2918,N_742);
and U3953 (N_3953,N_23,N_270);
nand U3954 (N_3954,N_259,N_786);
nor U3955 (N_3955,N_2149,N_377);
nand U3956 (N_3956,N_2246,N_1008);
nor U3957 (N_3957,N_1512,N_680);
xnor U3958 (N_3958,N_341,N_796);
and U3959 (N_3959,N_1676,N_973);
or U3960 (N_3960,N_1689,N_2608);
nor U3961 (N_3961,N_1434,N_111);
nor U3962 (N_3962,N_537,N_2965);
nand U3963 (N_3963,N_494,N_1970);
and U3964 (N_3964,N_1444,N_122);
or U3965 (N_3965,N_1229,N_71);
and U3966 (N_3966,N_2732,N_1144);
or U3967 (N_3967,N_1423,N_688);
nor U3968 (N_3968,N_1871,N_2639);
and U3969 (N_3969,N_2605,N_1763);
nand U3970 (N_3970,N_728,N_238);
or U3971 (N_3971,N_847,N_264);
nor U3972 (N_3972,N_1574,N_1897);
nor U3973 (N_3973,N_1054,N_1677);
or U3974 (N_3974,N_2972,N_366);
xor U3975 (N_3975,N_1355,N_746);
nand U3976 (N_3976,N_1333,N_18);
or U3977 (N_3977,N_2714,N_940);
nand U3978 (N_3978,N_662,N_781);
and U3979 (N_3979,N_1476,N_1731);
xor U3980 (N_3980,N_51,N_2544);
and U3981 (N_3981,N_1961,N_2271);
nor U3982 (N_3982,N_2411,N_2277);
nor U3983 (N_3983,N_697,N_1784);
nor U3984 (N_3984,N_2167,N_2027);
xor U3985 (N_3985,N_2581,N_418);
and U3986 (N_3986,N_409,N_293);
or U3987 (N_3987,N_2681,N_2345);
or U3988 (N_3988,N_1774,N_2306);
or U3989 (N_3989,N_528,N_1292);
nand U3990 (N_3990,N_723,N_628);
or U3991 (N_3991,N_2613,N_2624);
or U3992 (N_3992,N_2516,N_322);
nor U3993 (N_3993,N_593,N_2861);
xor U3994 (N_3994,N_1256,N_430);
or U3995 (N_3995,N_585,N_2628);
nand U3996 (N_3996,N_58,N_1929);
nor U3997 (N_3997,N_2673,N_484);
or U3998 (N_3998,N_1328,N_2981);
nand U3999 (N_3999,N_1185,N_1800);
or U4000 (N_4000,N_372,N_1834);
nor U4001 (N_4001,N_2785,N_1621);
and U4002 (N_4002,N_686,N_876);
nor U4003 (N_4003,N_52,N_721);
nand U4004 (N_4004,N_64,N_1651);
nand U4005 (N_4005,N_1098,N_736);
xor U4006 (N_4006,N_62,N_1488);
and U4007 (N_4007,N_707,N_2275);
nor U4008 (N_4008,N_952,N_1937);
nor U4009 (N_4009,N_241,N_2404);
nand U4010 (N_4010,N_950,N_1719);
or U4011 (N_4011,N_331,N_2615);
nand U4012 (N_4012,N_2235,N_1170);
or U4013 (N_4013,N_115,N_2619);
nand U4014 (N_4014,N_2782,N_1440);
or U4015 (N_4015,N_1991,N_88);
and U4016 (N_4016,N_308,N_2217);
or U4017 (N_4017,N_1071,N_2944);
and U4018 (N_4018,N_735,N_1952);
nor U4019 (N_4019,N_2797,N_555);
nand U4020 (N_4020,N_1138,N_1486);
and U4021 (N_4021,N_299,N_236);
nor U4022 (N_4022,N_2648,N_1353);
or U4023 (N_4023,N_330,N_2759);
nor U4024 (N_4024,N_2900,N_61);
nand U4025 (N_4025,N_767,N_622);
or U4026 (N_4026,N_2735,N_2657);
or U4027 (N_4027,N_2123,N_1962);
nor U4028 (N_4028,N_1254,N_268);
and U4029 (N_4029,N_1639,N_1720);
nor U4030 (N_4030,N_1271,N_884);
nor U4031 (N_4031,N_2358,N_966);
or U4032 (N_4032,N_2115,N_690);
or U4033 (N_4033,N_982,N_2043);
nand U4034 (N_4034,N_2347,N_2987);
and U4035 (N_4035,N_2251,N_412);
and U4036 (N_4036,N_2066,N_1183);
nand U4037 (N_4037,N_54,N_488);
nand U4038 (N_4038,N_904,N_170);
and U4039 (N_4039,N_1535,N_2426);
nor U4040 (N_4040,N_968,N_996);
nor U4041 (N_4041,N_1658,N_923);
xor U4042 (N_4042,N_1979,N_2894);
nor U4043 (N_4043,N_2499,N_990);
nand U4044 (N_4044,N_1508,N_677);
or U4045 (N_4045,N_927,N_131);
nor U4046 (N_4046,N_1769,N_1047);
or U4047 (N_4047,N_2412,N_873);
and U4048 (N_4048,N_1466,N_1710);
nand U4049 (N_4049,N_2652,N_2871);
nand U4050 (N_4050,N_1553,N_803);
and U4051 (N_4051,N_2781,N_587);
nor U4052 (N_4052,N_921,N_1035);
nand U4053 (N_4053,N_715,N_1281);
or U4054 (N_4054,N_564,N_2285);
nor U4055 (N_4055,N_525,N_2376);
nand U4056 (N_4056,N_482,N_286);
nor U4057 (N_4057,N_2634,N_2430);
and U4058 (N_4058,N_1128,N_1556);
or U4059 (N_4059,N_2453,N_27);
nor U4060 (N_4060,N_1565,N_2263);
or U4061 (N_4061,N_100,N_1277);
nor U4062 (N_4062,N_48,N_1227);
or U4063 (N_4063,N_2333,N_2354);
nor U4064 (N_4064,N_2103,N_2515);
nand U4065 (N_4065,N_2911,N_1329);
and U4066 (N_4066,N_251,N_2866);
and U4067 (N_4067,N_1668,N_1113);
xnor U4068 (N_4068,N_1414,N_2206);
xnor U4069 (N_4069,N_2222,N_239);
nor U4070 (N_4070,N_1978,N_770);
nand U4071 (N_4071,N_549,N_1905);
or U4072 (N_4072,N_96,N_1056);
and U4073 (N_4073,N_1748,N_2963);
xnor U4074 (N_4074,N_1982,N_1636);
or U4075 (N_4075,N_627,N_1721);
and U4076 (N_4076,N_2433,N_1517);
nand U4077 (N_4077,N_1424,N_761);
nand U4078 (N_4078,N_2266,N_1913);
nor U4079 (N_4079,N_843,N_2827);
and U4080 (N_4080,N_324,N_1852);
nor U4081 (N_4081,N_975,N_1785);
or U4082 (N_4082,N_1063,N_47);
or U4083 (N_4083,N_310,N_1564);
nand U4084 (N_4084,N_128,N_1549);
or U4085 (N_4085,N_2729,N_393);
and U4086 (N_4086,N_1285,N_2243);
or U4087 (N_4087,N_1609,N_1507);
and U4088 (N_4088,N_431,N_1149);
nor U4089 (N_4089,N_1032,N_1904);
nor U4090 (N_4090,N_1908,N_2770);
nand U4091 (N_4091,N_2215,N_1917);
or U4092 (N_4092,N_1097,N_2047);
and U4093 (N_4093,N_1884,N_2690);
nor U4094 (N_4094,N_937,N_683);
nor U4095 (N_4095,N_1914,N_1141);
xnor U4096 (N_4096,N_2706,N_77);
and U4097 (N_4097,N_1305,N_2746);
xor U4098 (N_4098,N_2359,N_473);
or U4099 (N_4099,N_250,N_1537);
and U4100 (N_4100,N_1086,N_2487);
and U4101 (N_4101,N_2152,N_720);
and U4102 (N_4102,N_1189,N_2890);
or U4103 (N_4103,N_245,N_256);
or U4104 (N_4104,N_1284,N_2008);
or U4105 (N_4105,N_1384,N_890);
and U4106 (N_4106,N_2968,N_2211);
nand U4107 (N_4107,N_2163,N_2071);
or U4108 (N_4108,N_2607,N_918);
or U4109 (N_4109,N_1019,N_2391);
nor U4110 (N_4110,N_1068,N_2915);
nand U4111 (N_4111,N_902,N_2234);
nor U4112 (N_4112,N_327,N_964);
nor U4113 (N_4113,N_800,N_2093);
nor U4114 (N_4114,N_2106,N_1958);
nand U4115 (N_4115,N_2028,N_222);
nor U4116 (N_4116,N_2847,N_501);
xnor U4117 (N_4117,N_1364,N_1751);
and U4118 (N_4118,N_2826,N_939);
nor U4119 (N_4119,N_636,N_1481);
and U4120 (N_4120,N_991,N_747);
nor U4121 (N_4121,N_1465,N_13);
and U4122 (N_4122,N_1690,N_2658);
nor U4123 (N_4123,N_40,N_97);
nand U4124 (N_4124,N_1727,N_451);
or U4125 (N_4125,N_2596,N_2804);
xor U4126 (N_4126,N_609,N_340);
and U4127 (N_4127,N_626,N_232);
nor U4128 (N_4128,N_188,N_1352);
nand U4129 (N_4129,N_857,N_2769);
or U4130 (N_4130,N_1879,N_386);
nor U4131 (N_4131,N_1495,N_201);
or U4132 (N_4132,N_2220,N_2922);
xnor U4133 (N_4133,N_2616,N_1240);
and U4134 (N_4134,N_2684,N_316);
nand U4135 (N_4135,N_436,N_1795);
or U4136 (N_4136,N_151,N_1046);
nand U4137 (N_4137,N_2446,N_2674);
and U4138 (N_4138,N_1122,N_531);
or U4139 (N_4139,N_1550,N_2315);
nand U4140 (N_4140,N_988,N_2837);
nor U4141 (N_4141,N_1013,N_1808);
nor U4142 (N_4142,N_1088,N_1620);
and U4143 (N_4143,N_1340,N_1180);
nor U4144 (N_4144,N_2814,N_1972);
and U4145 (N_4145,N_1346,N_272);
or U4146 (N_4146,N_886,N_1250);
nor U4147 (N_4147,N_2273,N_1893);
or U4148 (N_4148,N_2717,N_1778);
nor U4149 (N_4149,N_2088,N_1864);
nor U4150 (N_4150,N_1672,N_577);
and U4151 (N_4151,N_724,N_28);
nand U4152 (N_4152,N_1288,N_2556);
and U4153 (N_4153,N_1291,N_289);
or U4154 (N_4154,N_333,N_1530);
and U4155 (N_4155,N_1075,N_1176);
nor U4156 (N_4156,N_454,N_1474);
nor U4157 (N_4157,N_194,N_822);
and U4158 (N_4158,N_2294,N_212);
nand U4159 (N_4159,N_143,N_1794);
or U4160 (N_4160,N_1343,N_1341);
and U4161 (N_4161,N_1616,N_2895);
nor U4162 (N_4162,N_673,N_1354);
nand U4163 (N_4163,N_1060,N_2860);
nor U4164 (N_4164,N_2665,N_844);
nor U4165 (N_4165,N_1994,N_888);
or U4166 (N_4166,N_1447,N_127);
and U4167 (N_4167,N_2636,N_2368);
or U4168 (N_4168,N_496,N_145);
or U4169 (N_4169,N_2378,N_1023);
nor U4170 (N_4170,N_1807,N_1663);
nand U4171 (N_4171,N_2040,N_1242);
nand U4172 (N_4172,N_2631,N_2473);
nand U4173 (N_4173,N_2157,N_2381);
and U4174 (N_4174,N_1910,N_2421);
nor U4175 (N_4175,N_1977,N_398);
nor U4176 (N_4176,N_219,N_25);
or U4177 (N_4177,N_392,N_1847);
and U4178 (N_4178,N_748,N_1829);
or U4179 (N_4179,N_1205,N_2609);
or U4180 (N_4180,N_580,N_760);
or U4181 (N_4181,N_2659,N_522);
nand U4182 (N_4182,N_575,N_2154);
or U4183 (N_4183,N_1826,N_1594);
or U4184 (N_4184,N_527,N_1783);
nor U4185 (N_4185,N_978,N_2956);
or U4186 (N_4186,N_1209,N_1646);
and U4187 (N_4187,N_2023,N_1762);
nor U4188 (N_4188,N_2859,N_2902);
or U4189 (N_4189,N_2803,N_985);
and U4190 (N_4190,N_1057,N_2807);
nor U4191 (N_4191,N_2142,N_2817);
nor U4192 (N_4192,N_2590,N_2239);
nor U4193 (N_4193,N_1780,N_2990);
nor U4194 (N_4194,N_1367,N_1091);
nor U4195 (N_4195,N_1966,N_874);
nor U4196 (N_4196,N_1907,N_1614);
and U4197 (N_4197,N_518,N_1855);
xnor U4198 (N_4198,N_1799,N_535);
or U4199 (N_4199,N_2037,N_941);
nand U4200 (N_4200,N_381,N_2102);
and U4201 (N_4201,N_385,N_94);
or U4202 (N_4202,N_1089,N_1918);
nand U4203 (N_4203,N_1327,N_2689);
or U4204 (N_4204,N_7,N_1143);
and U4205 (N_4205,N_353,N_229);
nor U4206 (N_4206,N_740,N_1478);
and U4207 (N_4207,N_408,N_479);
or U4208 (N_4208,N_2960,N_552);
or U4209 (N_4209,N_2796,N_2342);
xnor U4210 (N_4210,N_2833,N_2579);
nand U4211 (N_4211,N_2288,N_1208);
xnor U4212 (N_4212,N_2887,N_2697);
and U4213 (N_4213,N_2650,N_2158);
and U4214 (N_4214,N_2070,N_576);
and U4215 (N_4215,N_2587,N_2518);
and U4216 (N_4216,N_2399,N_269);
and U4217 (N_4217,N_114,N_1289);
or U4218 (N_4218,N_35,N_184);
nor U4219 (N_4219,N_2325,N_1764);
and U4220 (N_4220,N_560,N_1310);
nand U4221 (N_4221,N_1637,N_1018);
and U4222 (N_4222,N_2898,N_345);
nor U4223 (N_4223,N_695,N_196);
nor U4224 (N_4224,N_2396,N_1882);
nor U4225 (N_4225,N_2630,N_1079);
and U4226 (N_4226,N_669,N_2862);
nand U4227 (N_4227,N_1730,N_2485);
nor U4228 (N_4228,N_1083,N_1015);
or U4229 (N_4229,N_1224,N_685);
or U4230 (N_4230,N_2114,N_1266);
nand U4231 (N_4231,N_1617,N_827);
or U4232 (N_4232,N_1085,N_1533);
or U4233 (N_4233,N_804,N_1022);
and U4234 (N_4234,N_63,N_214);
nor U4235 (N_4235,N_1049,N_1596);
and U4236 (N_4236,N_566,N_458);
or U4237 (N_4237,N_768,N_1030);
nor U4238 (N_4238,N_821,N_1371);
and U4239 (N_4239,N_95,N_1767);
or U4240 (N_4240,N_285,N_59);
nor U4241 (N_4241,N_1366,N_185);
nor U4242 (N_4242,N_1739,N_1836);
or U4243 (N_4243,N_1509,N_2195);
nand U4244 (N_4244,N_2535,N_1746);
and U4245 (N_4245,N_2176,N_2558);
nand U4246 (N_4246,N_2236,N_2546);
nand U4247 (N_4247,N_899,N_1033);
or U4248 (N_4248,N_34,N_1211);
nand U4249 (N_4249,N_866,N_920);
or U4250 (N_4250,N_2924,N_2041);
nor U4251 (N_4251,N_725,N_205);
and U4252 (N_4252,N_1491,N_955);
nor U4253 (N_4253,N_2459,N_864);
and U4254 (N_4254,N_462,N_1813);
and U4255 (N_4255,N_203,N_499);
nor U4256 (N_4256,N_2409,N_2340);
nor U4257 (N_4257,N_1529,N_1393);
and U4258 (N_4258,N_2704,N_2216);
nor U4259 (N_4259,N_1114,N_1494);
or U4260 (N_4260,N_2092,N_1665);
nand U4261 (N_4261,N_2978,N_1299);
and U4262 (N_4262,N_1398,N_2566);
nor U4263 (N_4263,N_787,N_93);
nor U4264 (N_4264,N_1623,N_762);
nand U4265 (N_4265,N_175,N_1409);
or U4266 (N_4266,N_388,N_347);
or U4267 (N_4267,N_465,N_2574);
xnor U4268 (N_4268,N_2604,N_2752);
and U4269 (N_4269,N_92,N_357);
and U4270 (N_4270,N_895,N_2177);
or U4271 (N_4271,N_1416,N_2004);
nor U4272 (N_4272,N_233,N_1302);
nand U4273 (N_4273,N_159,N_1458);
nor U4274 (N_4274,N_2897,N_1591);
nand U4275 (N_4275,N_863,N_1482);
and U4276 (N_4276,N_1638,N_1858);
and U4277 (N_4277,N_1026,N_1383);
nand U4278 (N_4278,N_477,N_2130);
and U4279 (N_4279,N_2820,N_2148);
nand U4280 (N_4280,N_2245,N_687);
or U4281 (N_4281,N_36,N_2649);
or U4282 (N_4282,N_2980,N_2675);
and U4283 (N_4283,N_1782,N_29);
nor U4284 (N_4284,N_588,N_2519);
xnor U4285 (N_4285,N_1190,N_2133);
nor U4286 (N_4286,N_2934,N_2932);
or U4287 (N_4287,N_1336,N_4);
nor U4288 (N_4288,N_2321,N_933);
nand U4289 (N_4289,N_1816,N_1678);
nor U4290 (N_4290,N_358,N_2916);
and U4291 (N_4291,N_1471,N_1927);
nor U4292 (N_4292,N_1021,N_1422);
and U4293 (N_4293,N_228,N_1042);
nor U4294 (N_4294,N_824,N_404);
nand U4295 (N_4295,N_671,N_1873);
nand U4296 (N_4296,N_670,N_949);
or U4297 (N_4297,N_1806,N_1164);
or U4298 (N_4298,N_2208,N_2279);
or U4299 (N_4299,N_2713,N_1260);
or U4300 (N_4300,N_1641,N_187);
xor U4301 (N_4301,N_2969,N_67);
nor U4302 (N_4302,N_1814,N_2493);
or U4303 (N_4303,N_1301,N_2873);
nand U4304 (N_4304,N_2730,N_472);
nand U4305 (N_4305,N_2552,N_782);
and U4306 (N_4306,N_989,N_174);
xnor U4307 (N_4307,N_1841,N_905);
and U4308 (N_4308,N_348,N_2369);
and U4309 (N_4309,N_606,N_1693);
nor U4310 (N_4310,N_2791,N_0);
nor U4311 (N_4311,N_520,N_1406);
nor U4312 (N_4312,N_910,N_2926);
and U4313 (N_4313,N_1622,N_1081);
or U4314 (N_4314,N_1761,N_413);
or U4315 (N_4315,N_2701,N_2393);
nor U4316 (N_4316,N_42,N_694);
nor U4317 (N_4317,N_1252,N_608);
and U4318 (N_4318,N_1654,N_2589);
or U4319 (N_4319,N_1726,N_167);
nor U4320 (N_4320,N_332,N_1174);
xor U4321 (N_4321,N_2744,N_2402);
xor U4322 (N_4322,N_2205,N_544);
or U4323 (N_4323,N_2380,N_2374);
xor U4324 (N_4324,N_519,N_1940);
xor U4325 (N_4325,N_2765,N_1473);
or U4326 (N_4326,N_486,N_2883);
or U4327 (N_4327,N_2175,N_1643);
and U4328 (N_4328,N_689,N_2122);
nand U4329 (N_4329,N_2268,N_1865);
and U4330 (N_4330,N_402,N_2562);
nand U4331 (N_4331,N_370,N_2332);
nor U4332 (N_4332,N_2034,N_958);
and U4333 (N_4333,N_1923,N_1531);
or U4334 (N_4334,N_2555,N_437);
xor U4335 (N_4335,N_2569,N_1156);
nand U4336 (N_4336,N_339,N_2946);
and U4337 (N_4337,N_1099,N_2419);
nand U4338 (N_4338,N_868,N_1687);
and U4339 (N_4339,N_60,N_2654);
nor U4340 (N_4340,N_563,N_2543);
nor U4341 (N_4341,N_2057,N_655);
nand U4342 (N_4342,N_2015,N_887);
or U4343 (N_4343,N_893,N_2472);
nand U4344 (N_4344,N_652,N_2394);
nand U4345 (N_4345,N_2210,N_591);
nand U4346 (N_4346,N_1460,N_2852);
or U4347 (N_4347,N_230,N_644);
or U4348 (N_4348,N_758,N_2580);
and U4349 (N_4349,N_862,N_751);
nor U4350 (N_4350,N_1796,N_1230);
or U4351 (N_4351,N_2875,N_2361);
and U4352 (N_4352,N_2073,N_2355);
nor U4353 (N_4353,N_73,N_1666);
nor U4354 (N_4354,N_2341,N_1470);
and U4355 (N_4355,N_2813,N_2858);
nor U4356 (N_4356,N_807,N_1653);
nand U4357 (N_4357,N_1804,N_1584);
or U4358 (N_4358,N_1418,N_1924);
nor U4359 (N_4359,N_161,N_774);
xor U4360 (N_4360,N_1044,N_1430);
and U4361 (N_4361,N_749,N_2733);
and U4362 (N_4362,N_571,N_2109);
nor U4363 (N_4363,N_2772,N_1433);
or U4364 (N_4364,N_2138,N_2483);
xnor U4365 (N_4365,N_618,N_314);
nand U4366 (N_4366,N_2724,N_2171);
and U4367 (N_4367,N_2020,N_1133);
or U4368 (N_4368,N_993,N_2212);
nor U4369 (N_4369,N_540,N_2484);
nand U4370 (N_4370,N_2437,N_1503);
xor U4371 (N_4371,N_443,N_113);
nand U4372 (N_4372,N_568,N_1944);
and U4373 (N_4373,N_1838,N_20);
nor U4374 (N_4374,N_1951,N_2882);
and U4375 (N_4375,N_2625,N_778);
or U4376 (N_4376,N_359,N_1313);
nor U4377 (N_4377,N_177,N_183);
xnor U4378 (N_4378,N_85,N_2451);
and U4379 (N_4379,N_1045,N_210);
nor U4380 (N_4380,N_2693,N_1325);
nor U4381 (N_4381,N_19,N_1542);
or U4382 (N_4382,N_1381,N_541);
and U4383 (N_4383,N_635,N_198);
xnor U4384 (N_4384,N_757,N_1510);
and U4385 (N_4385,N_1588,N_1338);
nand U4386 (N_4386,N_1467,N_2124);
nand U4387 (N_4387,N_959,N_908);
nor U4388 (N_4388,N_788,N_565);
xor U4389 (N_4389,N_11,N_186);
and U4390 (N_4390,N_1781,N_2146);
nor U4391 (N_4391,N_1691,N_2322);
xor U4392 (N_4392,N_2651,N_2108);
nand U4393 (N_4393,N_2818,N_3);
nor U4394 (N_4394,N_1360,N_2749);
nor U4395 (N_4395,N_619,N_1404);
and U4396 (N_4396,N_379,N_2776);
and U4397 (N_4397,N_722,N_1844);
nand U4398 (N_4398,N_2824,N_283);
nand U4399 (N_4399,N_2626,N_1969);
or U4400 (N_4400,N_850,N_37);
nor U4401 (N_4401,N_1093,N_972);
xor U4402 (N_4402,N_1053,N_2197);
xnor U4403 (N_4403,N_2129,N_1845);
nor U4404 (N_4404,N_2019,N_871);
and U4405 (N_4405,N_1545,N_2313);
nand U4406 (N_4406,N_1397,N_1725);
nand U4407 (N_4407,N_349,N_2529);
nor U4408 (N_4408,N_1983,N_2635);
nor U4409 (N_4409,N_983,N_2307);
or U4410 (N_4410,N_935,N_1437);
or U4411 (N_4411,N_2494,N_829);
or U4412 (N_4412,N_556,N_1365);
or U4413 (N_4413,N_1861,N_2303);
nand U4414 (N_4414,N_557,N_2469);
and U4415 (N_4415,N_865,N_1684);
nand U4416 (N_4416,N_1899,N_1498);
and U4417 (N_4417,N_1121,N_1275);
or U4418 (N_4418,N_2165,N_2295);
and U4419 (N_4419,N_190,N_2377);
or U4420 (N_4420,N_2068,N_2183);
and U4421 (N_4421,N_784,N_261);
nor U4422 (N_4422,N_1269,N_2316);
nand U4423 (N_4423,N_335,N_81);
nand U4424 (N_4424,N_2985,N_2218);
nor U4425 (N_4425,N_1107,N_2283);
nor U4426 (N_4426,N_1009,N_1610);
or U4427 (N_4427,N_2363,N_1314);
or U4428 (N_4428,N_2936,N_1747);
and U4429 (N_4429,N_2570,N_825);
nand U4430 (N_4430,N_1866,N_2425);
or U4431 (N_4431,N_2024,N_2792);
and U4432 (N_4432,N_1587,N_2888);
nand U4433 (N_4433,N_558,N_181);
xnor U4434 (N_4434,N_334,N_171);
nor U4435 (N_4435,N_1628,N_992);
xnor U4436 (N_4436,N_623,N_1419);
or U4437 (N_4437,N_301,N_1874);
nand U4438 (N_4438,N_1544,N_1159);
nand U4439 (N_4439,N_2829,N_894);
xor U4440 (N_4440,N_592,N_1123);
nand U4441 (N_4441,N_2839,N_1843);
and U4442 (N_4442,N_2077,N_415);
xor U4443 (N_4443,N_5,N_328);
and U4444 (N_4444,N_1038,N_2726);
nand U4445 (N_4445,N_1860,N_699);
nor U4446 (N_4446,N_651,N_659);
and U4447 (N_4447,N_2643,N_1942);
xor U4448 (N_4448,N_2463,N_211);
xnor U4449 (N_4449,N_1375,N_1863);
nor U4450 (N_4450,N_795,N_516);
or U4451 (N_4451,N_915,N_909);
nand U4452 (N_4452,N_526,N_2768);
nor U4453 (N_4453,N_898,N_1578);
nand U4454 (N_4454,N_2116,N_1920);
nand U4455 (N_4455,N_2031,N_533);
or U4456 (N_4456,N_956,N_311);
nand U4457 (N_4457,N_1941,N_191);
nor U4458 (N_4458,N_1854,N_382);
xnor U4459 (N_4459,N_2039,N_911);
and U4460 (N_4460,N_1595,N_2438);
nand U4461 (N_4461,N_1729,N_583);
nor U4462 (N_4462,N_2617,N_288);
and U4463 (N_4463,N_1990,N_1554);
nand U4464 (N_4464,N_416,N_2921);
or U4465 (N_4465,N_215,N_639);
nor U4466 (N_4466,N_1443,N_294);
nor U4467 (N_4467,N_2127,N_1593);
nand U4468 (N_4468,N_1985,N_2301);
nor U4469 (N_4469,N_2557,N_2098);
nor U4470 (N_4470,N_1248,N_2528);
nor U4471 (N_4471,N_2509,N_1050);
or U4472 (N_4472,N_2337,N_2727);
nand U4473 (N_4473,N_875,N_2786);
nand U4474 (N_4474,N_631,N_2984);
xnor U4475 (N_4475,N_68,N_2060);
or U4476 (N_4476,N_82,N_1167);
nor U4477 (N_4477,N_1713,N_1903);
or U4478 (N_4478,N_2599,N_919);
or U4479 (N_4479,N_1092,N_661);
nor U4480 (N_4480,N_2950,N_1557);
or U4481 (N_4481,N_523,N_1456);
or U4482 (N_4482,N_780,N_1145);
or U4483 (N_4483,N_390,N_1307);
and U4484 (N_4484,N_976,N_726);
or U4485 (N_4485,N_2641,N_1694);
and U4486 (N_4486,N_666,N_1132);
xor U4487 (N_4487,N_806,N_1251);
or U4488 (N_4488,N_1134,N_2497);
xor U4489 (N_4489,N_1824,N_667);
nor U4490 (N_4490,N_1631,N_980);
and U4491 (N_4491,N_234,N_1830);
and U4492 (N_4492,N_1810,N_2647);
and U4493 (N_4493,N_2513,N_998);
nand U4494 (N_4494,N_1502,N_737);
or U4495 (N_4495,N_2671,N_1001);
or U4496 (N_4496,N_2811,N_954);
nand U4497 (N_4497,N_2470,N_199);
and U4498 (N_4498,N_2920,N_1497);
nor U4499 (N_4499,N_750,N_977);
and U4500 (N_4500,N_1319,N_1666);
nand U4501 (N_4501,N_595,N_901);
nor U4502 (N_4502,N_407,N_2354);
nor U4503 (N_4503,N_559,N_1884);
and U4504 (N_4504,N_2030,N_2946);
nand U4505 (N_4505,N_510,N_689);
nand U4506 (N_4506,N_2972,N_1986);
nor U4507 (N_4507,N_1502,N_710);
and U4508 (N_4508,N_2462,N_1850);
and U4509 (N_4509,N_1113,N_369);
and U4510 (N_4510,N_2803,N_1839);
or U4511 (N_4511,N_74,N_966);
and U4512 (N_4512,N_2902,N_824);
or U4513 (N_4513,N_2318,N_470);
and U4514 (N_4514,N_704,N_1506);
nor U4515 (N_4515,N_759,N_2121);
or U4516 (N_4516,N_1763,N_831);
or U4517 (N_4517,N_1220,N_2726);
nor U4518 (N_4518,N_2381,N_1488);
nor U4519 (N_4519,N_1361,N_334);
and U4520 (N_4520,N_1701,N_1104);
or U4521 (N_4521,N_788,N_1179);
nand U4522 (N_4522,N_1970,N_2868);
or U4523 (N_4523,N_1011,N_2780);
and U4524 (N_4524,N_1399,N_948);
xnor U4525 (N_4525,N_1970,N_802);
nor U4526 (N_4526,N_140,N_58);
nor U4527 (N_4527,N_1248,N_727);
nor U4528 (N_4528,N_260,N_2083);
or U4529 (N_4529,N_970,N_1218);
and U4530 (N_4530,N_299,N_1726);
or U4531 (N_4531,N_357,N_428);
nor U4532 (N_4532,N_182,N_2650);
xor U4533 (N_4533,N_696,N_519);
nand U4534 (N_4534,N_1647,N_1372);
and U4535 (N_4535,N_2580,N_2715);
and U4536 (N_4536,N_2132,N_2809);
nor U4537 (N_4537,N_2928,N_155);
or U4538 (N_4538,N_2311,N_2797);
nand U4539 (N_4539,N_592,N_1338);
or U4540 (N_4540,N_2802,N_394);
xnor U4541 (N_4541,N_2674,N_399);
and U4542 (N_4542,N_2448,N_1831);
nor U4543 (N_4543,N_2065,N_2854);
or U4544 (N_4544,N_92,N_2848);
or U4545 (N_4545,N_2356,N_957);
xnor U4546 (N_4546,N_1996,N_486);
nand U4547 (N_4547,N_904,N_775);
and U4548 (N_4548,N_1560,N_1925);
nor U4549 (N_4549,N_341,N_1285);
nand U4550 (N_4550,N_2957,N_1860);
nand U4551 (N_4551,N_418,N_2770);
nor U4552 (N_4552,N_288,N_486);
nand U4553 (N_4553,N_531,N_1346);
nand U4554 (N_4554,N_275,N_2212);
xnor U4555 (N_4555,N_1565,N_2678);
or U4556 (N_4556,N_450,N_123);
nor U4557 (N_4557,N_2546,N_277);
nor U4558 (N_4558,N_1013,N_2808);
nand U4559 (N_4559,N_1906,N_2482);
and U4560 (N_4560,N_1186,N_317);
nand U4561 (N_4561,N_846,N_564);
nand U4562 (N_4562,N_2080,N_156);
or U4563 (N_4563,N_2022,N_222);
and U4564 (N_4564,N_2305,N_1916);
and U4565 (N_4565,N_2636,N_2668);
and U4566 (N_4566,N_2502,N_1065);
xor U4567 (N_4567,N_2900,N_2203);
nand U4568 (N_4568,N_2650,N_1181);
or U4569 (N_4569,N_615,N_970);
nor U4570 (N_4570,N_633,N_2040);
nor U4571 (N_4571,N_514,N_1811);
and U4572 (N_4572,N_1826,N_2382);
nor U4573 (N_4573,N_1123,N_1923);
and U4574 (N_4574,N_1320,N_2546);
xor U4575 (N_4575,N_1004,N_2279);
or U4576 (N_4576,N_146,N_961);
or U4577 (N_4577,N_1174,N_1828);
or U4578 (N_4578,N_557,N_46);
and U4579 (N_4579,N_1751,N_1685);
and U4580 (N_4580,N_123,N_308);
and U4581 (N_4581,N_1417,N_2408);
nand U4582 (N_4582,N_339,N_1915);
xor U4583 (N_4583,N_1908,N_1466);
nand U4584 (N_4584,N_1364,N_1439);
or U4585 (N_4585,N_387,N_2926);
nor U4586 (N_4586,N_2589,N_651);
and U4587 (N_4587,N_1741,N_2359);
nand U4588 (N_4588,N_1550,N_1566);
nor U4589 (N_4589,N_87,N_432);
nor U4590 (N_4590,N_1597,N_2960);
nand U4591 (N_4591,N_2884,N_1197);
nand U4592 (N_4592,N_1208,N_544);
and U4593 (N_4593,N_1968,N_886);
or U4594 (N_4594,N_795,N_660);
nand U4595 (N_4595,N_942,N_1716);
nor U4596 (N_4596,N_204,N_1607);
or U4597 (N_4597,N_522,N_2878);
nor U4598 (N_4598,N_2494,N_1234);
or U4599 (N_4599,N_1334,N_1445);
nor U4600 (N_4600,N_724,N_2997);
or U4601 (N_4601,N_1351,N_2462);
and U4602 (N_4602,N_1499,N_706);
nand U4603 (N_4603,N_2984,N_1451);
or U4604 (N_4604,N_2536,N_1384);
nand U4605 (N_4605,N_2390,N_914);
and U4606 (N_4606,N_2372,N_1991);
or U4607 (N_4607,N_1590,N_2550);
or U4608 (N_4608,N_578,N_2313);
nand U4609 (N_4609,N_1266,N_390);
nor U4610 (N_4610,N_192,N_369);
or U4611 (N_4611,N_2856,N_1896);
nor U4612 (N_4612,N_1374,N_2075);
or U4613 (N_4613,N_1656,N_2526);
and U4614 (N_4614,N_2690,N_2759);
or U4615 (N_4615,N_1209,N_2986);
and U4616 (N_4616,N_1601,N_2318);
or U4617 (N_4617,N_1531,N_1613);
and U4618 (N_4618,N_1002,N_2055);
and U4619 (N_4619,N_248,N_236);
nand U4620 (N_4620,N_998,N_1489);
and U4621 (N_4621,N_1229,N_1214);
or U4622 (N_4622,N_1948,N_1886);
nor U4623 (N_4623,N_1381,N_2831);
or U4624 (N_4624,N_781,N_696);
or U4625 (N_4625,N_967,N_18);
nand U4626 (N_4626,N_2333,N_1323);
and U4627 (N_4627,N_2846,N_1786);
and U4628 (N_4628,N_1497,N_2244);
and U4629 (N_4629,N_2881,N_1674);
nor U4630 (N_4630,N_443,N_1617);
nor U4631 (N_4631,N_2510,N_1989);
or U4632 (N_4632,N_1412,N_706);
nor U4633 (N_4633,N_400,N_1998);
and U4634 (N_4634,N_1994,N_2441);
xor U4635 (N_4635,N_1815,N_94);
nor U4636 (N_4636,N_978,N_1780);
nor U4637 (N_4637,N_2052,N_657);
and U4638 (N_4638,N_986,N_555);
nor U4639 (N_4639,N_1011,N_1885);
or U4640 (N_4640,N_1856,N_1457);
nor U4641 (N_4641,N_2893,N_2914);
xnor U4642 (N_4642,N_1277,N_1438);
nand U4643 (N_4643,N_2686,N_1528);
nor U4644 (N_4644,N_2507,N_2163);
and U4645 (N_4645,N_29,N_2301);
nand U4646 (N_4646,N_2545,N_1256);
or U4647 (N_4647,N_2975,N_661);
nand U4648 (N_4648,N_2957,N_2790);
nand U4649 (N_4649,N_2894,N_1955);
nor U4650 (N_4650,N_1705,N_1673);
and U4651 (N_4651,N_2603,N_2520);
nor U4652 (N_4652,N_635,N_974);
and U4653 (N_4653,N_707,N_2486);
and U4654 (N_4654,N_2433,N_2889);
or U4655 (N_4655,N_7,N_1189);
nand U4656 (N_4656,N_1279,N_2132);
or U4657 (N_4657,N_1295,N_2067);
and U4658 (N_4658,N_1102,N_1319);
and U4659 (N_4659,N_73,N_76);
nand U4660 (N_4660,N_1753,N_1421);
and U4661 (N_4661,N_985,N_350);
nor U4662 (N_4662,N_784,N_2993);
nor U4663 (N_4663,N_932,N_636);
and U4664 (N_4664,N_2799,N_1051);
or U4665 (N_4665,N_317,N_1461);
and U4666 (N_4666,N_2323,N_2508);
nand U4667 (N_4667,N_2206,N_2746);
and U4668 (N_4668,N_149,N_1223);
and U4669 (N_4669,N_2076,N_2611);
nand U4670 (N_4670,N_2179,N_1353);
xnor U4671 (N_4671,N_1443,N_2884);
xnor U4672 (N_4672,N_1693,N_130);
nor U4673 (N_4673,N_411,N_76);
nand U4674 (N_4674,N_1755,N_2356);
and U4675 (N_4675,N_2715,N_1674);
nand U4676 (N_4676,N_1273,N_2360);
and U4677 (N_4677,N_2522,N_2718);
xnor U4678 (N_4678,N_971,N_2545);
or U4679 (N_4679,N_203,N_702);
nor U4680 (N_4680,N_57,N_899);
and U4681 (N_4681,N_711,N_1325);
and U4682 (N_4682,N_1980,N_638);
xnor U4683 (N_4683,N_707,N_2644);
nor U4684 (N_4684,N_2262,N_1379);
and U4685 (N_4685,N_2411,N_2501);
or U4686 (N_4686,N_1256,N_363);
and U4687 (N_4687,N_273,N_539);
nor U4688 (N_4688,N_936,N_908);
nor U4689 (N_4689,N_2950,N_2092);
nand U4690 (N_4690,N_12,N_1094);
nand U4691 (N_4691,N_741,N_706);
nand U4692 (N_4692,N_536,N_1222);
nand U4693 (N_4693,N_1947,N_2843);
and U4694 (N_4694,N_2239,N_1995);
nor U4695 (N_4695,N_99,N_2150);
xor U4696 (N_4696,N_2449,N_1735);
or U4697 (N_4697,N_1215,N_1238);
nand U4698 (N_4698,N_1168,N_977);
and U4699 (N_4699,N_2597,N_2054);
nand U4700 (N_4700,N_2197,N_1304);
nor U4701 (N_4701,N_2442,N_492);
nand U4702 (N_4702,N_131,N_374);
xnor U4703 (N_4703,N_2986,N_566);
and U4704 (N_4704,N_630,N_2313);
nor U4705 (N_4705,N_1752,N_1082);
nor U4706 (N_4706,N_776,N_1121);
nor U4707 (N_4707,N_1005,N_1629);
xnor U4708 (N_4708,N_1477,N_2436);
and U4709 (N_4709,N_1437,N_1012);
nand U4710 (N_4710,N_2770,N_1069);
nor U4711 (N_4711,N_1642,N_875);
nor U4712 (N_4712,N_2368,N_1643);
or U4713 (N_4713,N_2726,N_311);
nor U4714 (N_4714,N_2999,N_2309);
nor U4715 (N_4715,N_1382,N_2732);
and U4716 (N_4716,N_1657,N_2265);
nor U4717 (N_4717,N_162,N_2851);
nor U4718 (N_4718,N_2496,N_2302);
nor U4719 (N_4719,N_2394,N_1346);
nor U4720 (N_4720,N_2908,N_29);
nand U4721 (N_4721,N_537,N_2942);
nor U4722 (N_4722,N_2629,N_2771);
and U4723 (N_4723,N_1542,N_2968);
nor U4724 (N_4724,N_1700,N_2819);
nand U4725 (N_4725,N_2851,N_1859);
and U4726 (N_4726,N_1614,N_2176);
nand U4727 (N_4727,N_1237,N_2597);
nand U4728 (N_4728,N_1658,N_273);
and U4729 (N_4729,N_1891,N_1621);
nand U4730 (N_4730,N_860,N_1432);
and U4731 (N_4731,N_2686,N_1662);
and U4732 (N_4732,N_1250,N_192);
and U4733 (N_4733,N_2902,N_981);
and U4734 (N_4734,N_2417,N_741);
nor U4735 (N_4735,N_1026,N_2151);
nor U4736 (N_4736,N_866,N_2565);
or U4737 (N_4737,N_1964,N_580);
nand U4738 (N_4738,N_1617,N_807);
and U4739 (N_4739,N_1665,N_222);
nand U4740 (N_4740,N_2662,N_689);
or U4741 (N_4741,N_2441,N_2768);
and U4742 (N_4742,N_2779,N_917);
nor U4743 (N_4743,N_733,N_1090);
nor U4744 (N_4744,N_2952,N_157);
xor U4745 (N_4745,N_58,N_264);
or U4746 (N_4746,N_1766,N_1020);
nor U4747 (N_4747,N_1837,N_2506);
nand U4748 (N_4748,N_940,N_2965);
or U4749 (N_4749,N_2155,N_1985);
or U4750 (N_4750,N_1890,N_2036);
nor U4751 (N_4751,N_2532,N_2776);
or U4752 (N_4752,N_1294,N_2111);
nand U4753 (N_4753,N_1173,N_1543);
nand U4754 (N_4754,N_323,N_207);
or U4755 (N_4755,N_176,N_14);
nor U4756 (N_4756,N_1045,N_2927);
xor U4757 (N_4757,N_57,N_2984);
xor U4758 (N_4758,N_2976,N_846);
xnor U4759 (N_4759,N_887,N_730);
or U4760 (N_4760,N_1575,N_1548);
nor U4761 (N_4761,N_498,N_18);
nor U4762 (N_4762,N_1383,N_1975);
and U4763 (N_4763,N_1936,N_2222);
xnor U4764 (N_4764,N_1062,N_66);
nand U4765 (N_4765,N_711,N_2608);
or U4766 (N_4766,N_1069,N_2044);
nor U4767 (N_4767,N_1018,N_8);
nand U4768 (N_4768,N_821,N_871);
nor U4769 (N_4769,N_1742,N_2984);
nand U4770 (N_4770,N_1247,N_525);
and U4771 (N_4771,N_2386,N_1377);
nand U4772 (N_4772,N_1112,N_1653);
nor U4773 (N_4773,N_2091,N_1670);
nor U4774 (N_4774,N_1271,N_124);
and U4775 (N_4775,N_804,N_334);
nor U4776 (N_4776,N_1760,N_1863);
and U4777 (N_4777,N_121,N_754);
nor U4778 (N_4778,N_52,N_756);
and U4779 (N_4779,N_2675,N_983);
nand U4780 (N_4780,N_899,N_2845);
and U4781 (N_4781,N_742,N_1528);
nand U4782 (N_4782,N_2395,N_1363);
and U4783 (N_4783,N_1706,N_1374);
or U4784 (N_4784,N_2194,N_1300);
or U4785 (N_4785,N_1531,N_181);
nand U4786 (N_4786,N_1386,N_2411);
and U4787 (N_4787,N_1635,N_2756);
nand U4788 (N_4788,N_215,N_107);
or U4789 (N_4789,N_959,N_18);
nor U4790 (N_4790,N_2976,N_2402);
or U4791 (N_4791,N_2435,N_1632);
nor U4792 (N_4792,N_136,N_2592);
and U4793 (N_4793,N_1669,N_1508);
nand U4794 (N_4794,N_826,N_723);
or U4795 (N_4795,N_657,N_1560);
xnor U4796 (N_4796,N_2441,N_2925);
nor U4797 (N_4797,N_2839,N_2851);
and U4798 (N_4798,N_2117,N_989);
or U4799 (N_4799,N_2118,N_882);
and U4800 (N_4800,N_404,N_487);
xnor U4801 (N_4801,N_1691,N_505);
and U4802 (N_4802,N_2934,N_2335);
nand U4803 (N_4803,N_177,N_2897);
xnor U4804 (N_4804,N_1178,N_140);
nand U4805 (N_4805,N_2246,N_789);
and U4806 (N_4806,N_617,N_733);
or U4807 (N_4807,N_759,N_2935);
xor U4808 (N_4808,N_705,N_1768);
xor U4809 (N_4809,N_834,N_1521);
nand U4810 (N_4810,N_1145,N_2258);
nand U4811 (N_4811,N_1802,N_501);
or U4812 (N_4812,N_278,N_2612);
xor U4813 (N_4813,N_2948,N_2015);
or U4814 (N_4814,N_2778,N_2048);
nor U4815 (N_4815,N_1542,N_1224);
nor U4816 (N_4816,N_726,N_1587);
or U4817 (N_4817,N_1168,N_1651);
nand U4818 (N_4818,N_2561,N_448);
or U4819 (N_4819,N_2524,N_244);
xnor U4820 (N_4820,N_1404,N_1524);
or U4821 (N_4821,N_1216,N_1843);
or U4822 (N_4822,N_1952,N_517);
or U4823 (N_4823,N_223,N_2580);
and U4824 (N_4824,N_700,N_1508);
or U4825 (N_4825,N_2415,N_37);
xnor U4826 (N_4826,N_280,N_158);
or U4827 (N_4827,N_1779,N_2793);
or U4828 (N_4828,N_2157,N_578);
or U4829 (N_4829,N_817,N_1518);
xnor U4830 (N_4830,N_1355,N_17);
nand U4831 (N_4831,N_2363,N_1981);
nand U4832 (N_4832,N_2452,N_464);
nor U4833 (N_4833,N_689,N_1229);
xnor U4834 (N_4834,N_813,N_2274);
nand U4835 (N_4835,N_2078,N_1935);
nor U4836 (N_4836,N_1322,N_2683);
nor U4837 (N_4837,N_1705,N_2608);
xnor U4838 (N_4838,N_2528,N_987);
and U4839 (N_4839,N_1497,N_1479);
and U4840 (N_4840,N_1378,N_476);
nor U4841 (N_4841,N_2035,N_2339);
or U4842 (N_4842,N_985,N_2893);
and U4843 (N_4843,N_2603,N_2185);
nand U4844 (N_4844,N_1532,N_1947);
and U4845 (N_4845,N_1926,N_1958);
nor U4846 (N_4846,N_172,N_235);
or U4847 (N_4847,N_1645,N_2836);
or U4848 (N_4848,N_389,N_1126);
nor U4849 (N_4849,N_2976,N_1598);
xnor U4850 (N_4850,N_1278,N_2483);
or U4851 (N_4851,N_2749,N_1384);
or U4852 (N_4852,N_1797,N_1914);
xnor U4853 (N_4853,N_1077,N_2259);
nor U4854 (N_4854,N_1620,N_692);
and U4855 (N_4855,N_1052,N_2431);
xnor U4856 (N_4856,N_1831,N_2204);
and U4857 (N_4857,N_1286,N_2105);
nor U4858 (N_4858,N_2266,N_2766);
nor U4859 (N_4859,N_2046,N_2466);
nand U4860 (N_4860,N_1176,N_737);
or U4861 (N_4861,N_379,N_579);
or U4862 (N_4862,N_434,N_1261);
and U4863 (N_4863,N_241,N_2963);
and U4864 (N_4864,N_1037,N_1076);
and U4865 (N_4865,N_1646,N_2075);
nor U4866 (N_4866,N_1995,N_280);
nor U4867 (N_4867,N_2956,N_193);
or U4868 (N_4868,N_852,N_301);
nand U4869 (N_4869,N_1081,N_1528);
nand U4870 (N_4870,N_2280,N_517);
or U4871 (N_4871,N_2321,N_278);
or U4872 (N_4872,N_1618,N_2632);
xor U4873 (N_4873,N_2575,N_714);
xor U4874 (N_4874,N_775,N_2884);
nor U4875 (N_4875,N_1660,N_311);
or U4876 (N_4876,N_1624,N_406);
xnor U4877 (N_4877,N_2220,N_969);
and U4878 (N_4878,N_2410,N_1570);
nor U4879 (N_4879,N_2698,N_1474);
nor U4880 (N_4880,N_2753,N_224);
or U4881 (N_4881,N_2559,N_1531);
or U4882 (N_4882,N_2691,N_1098);
nand U4883 (N_4883,N_418,N_2051);
nand U4884 (N_4884,N_2632,N_2745);
and U4885 (N_4885,N_703,N_539);
xor U4886 (N_4886,N_2485,N_1041);
or U4887 (N_4887,N_602,N_2318);
nand U4888 (N_4888,N_962,N_263);
or U4889 (N_4889,N_1106,N_579);
and U4890 (N_4890,N_2444,N_1122);
nor U4891 (N_4891,N_2421,N_2372);
or U4892 (N_4892,N_1341,N_1521);
and U4893 (N_4893,N_1562,N_963);
nand U4894 (N_4894,N_2838,N_325);
and U4895 (N_4895,N_1223,N_194);
nor U4896 (N_4896,N_409,N_133);
nor U4897 (N_4897,N_2708,N_2426);
nand U4898 (N_4898,N_1787,N_2997);
nor U4899 (N_4899,N_1914,N_2036);
and U4900 (N_4900,N_1934,N_1529);
nor U4901 (N_4901,N_1708,N_26);
nor U4902 (N_4902,N_2416,N_2961);
xor U4903 (N_4903,N_2815,N_812);
or U4904 (N_4904,N_28,N_835);
xor U4905 (N_4905,N_380,N_2025);
or U4906 (N_4906,N_1478,N_1543);
or U4907 (N_4907,N_2277,N_1152);
or U4908 (N_4908,N_1634,N_958);
xor U4909 (N_4909,N_1091,N_1189);
and U4910 (N_4910,N_1448,N_2199);
nand U4911 (N_4911,N_2586,N_1343);
nor U4912 (N_4912,N_866,N_582);
nor U4913 (N_4913,N_285,N_2586);
nand U4914 (N_4914,N_2696,N_360);
or U4915 (N_4915,N_423,N_65);
nand U4916 (N_4916,N_1894,N_693);
nand U4917 (N_4917,N_1147,N_2227);
or U4918 (N_4918,N_2371,N_1212);
nand U4919 (N_4919,N_2813,N_1026);
nor U4920 (N_4920,N_2677,N_1377);
and U4921 (N_4921,N_534,N_2596);
or U4922 (N_4922,N_1839,N_2402);
and U4923 (N_4923,N_346,N_42);
nand U4924 (N_4924,N_440,N_2574);
nor U4925 (N_4925,N_514,N_1046);
nor U4926 (N_4926,N_1065,N_1003);
nor U4927 (N_4927,N_339,N_2973);
or U4928 (N_4928,N_880,N_2389);
or U4929 (N_4929,N_1249,N_2100);
or U4930 (N_4930,N_2639,N_984);
and U4931 (N_4931,N_710,N_456);
nor U4932 (N_4932,N_945,N_2988);
nand U4933 (N_4933,N_1702,N_1099);
or U4934 (N_4934,N_2591,N_520);
or U4935 (N_4935,N_2364,N_393);
nor U4936 (N_4936,N_2573,N_1158);
xnor U4937 (N_4937,N_860,N_2103);
or U4938 (N_4938,N_1587,N_229);
nor U4939 (N_4939,N_2388,N_782);
nor U4940 (N_4940,N_21,N_1779);
nor U4941 (N_4941,N_1306,N_2316);
xor U4942 (N_4942,N_30,N_2526);
and U4943 (N_4943,N_1497,N_942);
and U4944 (N_4944,N_147,N_530);
nand U4945 (N_4945,N_1498,N_2252);
nor U4946 (N_4946,N_224,N_2633);
nand U4947 (N_4947,N_472,N_1916);
nand U4948 (N_4948,N_631,N_1305);
xnor U4949 (N_4949,N_1229,N_1082);
xor U4950 (N_4950,N_2098,N_1618);
and U4951 (N_4951,N_1658,N_2352);
and U4952 (N_4952,N_2173,N_2293);
or U4953 (N_4953,N_1551,N_2981);
nor U4954 (N_4954,N_882,N_2319);
nand U4955 (N_4955,N_2886,N_1110);
or U4956 (N_4956,N_161,N_2771);
xor U4957 (N_4957,N_789,N_296);
nor U4958 (N_4958,N_125,N_1362);
or U4959 (N_4959,N_2396,N_1102);
nand U4960 (N_4960,N_223,N_1152);
or U4961 (N_4961,N_2741,N_2599);
and U4962 (N_4962,N_2297,N_795);
nor U4963 (N_4963,N_2579,N_2164);
nand U4964 (N_4964,N_2646,N_2603);
nor U4965 (N_4965,N_1076,N_2416);
or U4966 (N_4966,N_1460,N_2665);
nor U4967 (N_4967,N_421,N_2613);
nor U4968 (N_4968,N_2792,N_62);
and U4969 (N_4969,N_752,N_1179);
or U4970 (N_4970,N_2299,N_678);
xnor U4971 (N_4971,N_506,N_492);
or U4972 (N_4972,N_2587,N_396);
or U4973 (N_4973,N_960,N_2326);
and U4974 (N_4974,N_631,N_1520);
nor U4975 (N_4975,N_1648,N_865);
or U4976 (N_4976,N_26,N_2122);
nand U4977 (N_4977,N_1289,N_246);
nand U4978 (N_4978,N_716,N_1741);
and U4979 (N_4979,N_2782,N_579);
nand U4980 (N_4980,N_2547,N_2219);
or U4981 (N_4981,N_665,N_791);
xor U4982 (N_4982,N_2639,N_654);
and U4983 (N_4983,N_1667,N_2490);
and U4984 (N_4984,N_906,N_431);
xor U4985 (N_4985,N_451,N_2509);
or U4986 (N_4986,N_601,N_2102);
nand U4987 (N_4987,N_980,N_489);
or U4988 (N_4988,N_2399,N_1359);
nor U4989 (N_4989,N_75,N_2263);
nor U4990 (N_4990,N_2701,N_1244);
and U4991 (N_4991,N_368,N_2241);
nor U4992 (N_4992,N_296,N_907);
or U4993 (N_4993,N_1292,N_1499);
xor U4994 (N_4994,N_788,N_2545);
and U4995 (N_4995,N_2392,N_1710);
nor U4996 (N_4996,N_135,N_867);
and U4997 (N_4997,N_133,N_83);
or U4998 (N_4998,N_2493,N_1939);
and U4999 (N_4999,N_2799,N_2052);
or U5000 (N_5000,N_252,N_2443);
nand U5001 (N_5001,N_181,N_2977);
or U5002 (N_5002,N_808,N_1296);
or U5003 (N_5003,N_760,N_706);
nand U5004 (N_5004,N_2115,N_1358);
nor U5005 (N_5005,N_1464,N_174);
nand U5006 (N_5006,N_2085,N_1156);
nand U5007 (N_5007,N_2865,N_2107);
nor U5008 (N_5008,N_412,N_622);
nand U5009 (N_5009,N_184,N_1473);
nor U5010 (N_5010,N_1605,N_2627);
xor U5011 (N_5011,N_2605,N_2435);
nand U5012 (N_5012,N_642,N_1671);
and U5013 (N_5013,N_2348,N_1192);
xor U5014 (N_5014,N_732,N_725);
and U5015 (N_5015,N_2903,N_398);
nor U5016 (N_5016,N_135,N_1469);
nand U5017 (N_5017,N_953,N_1798);
xor U5018 (N_5018,N_1335,N_856);
or U5019 (N_5019,N_937,N_1685);
or U5020 (N_5020,N_2417,N_2779);
nand U5021 (N_5021,N_693,N_2940);
xnor U5022 (N_5022,N_2660,N_471);
and U5023 (N_5023,N_2435,N_2232);
or U5024 (N_5024,N_855,N_2109);
nor U5025 (N_5025,N_2519,N_2732);
and U5026 (N_5026,N_2272,N_63);
nor U5027 (N_5027,N_100,N_1484);
nand U5028 (N_5028,N_1337,N_1413);
nand U5029 (N_5029,N_530,N_1287);
xor U5030 (N_5030,N_2396,N_2825);
nor U5031 (N_5031,N_1762,N_2549);
nand U5032 (N_5032,N_2644,N_2226);
nor U5033 (N_5033,N_2997,N_1412);
or U5034 (N_5034,N_494,N_1565);
nor U5035 (N_5035,N_1524,N_2286);
and U5036 (N_5036,N_1386,N_2443);
or U5037 (N_5037,N_902,N_191);
or U5038 (N_5038,N_1966,N_50);
and U5039 (N_5039,N_906,N_2217);
nand U5040 (N_5040,N_589,N_1525);
or U5041 (N_5041,N_1121,N_2940);
nand U5042 (N_5042,N_263,N_1953);
and U5043 (N_5043,N_1389,N_570);
nor U5044 (N_5044,N_2818,N_2480);
nor U5045 (N_5045,N_2829,N_1667);
nand U5046 (N_5046,N_1503,N_900);
or U5047 (N_5047,N_1420,N_2646);
xor U5048 (N_5048,N_2391,N_592);
or U5049 (N_5049,N_980,N_1756);
and U5050 (N_5050,N_1758,N_1735);
nand U5051 (N_5051,N_2701,N_2366);
nand U5052 (N_5052,N_564,N_1516);
nand U5053 (N_5053,N_1231,N_2268);
nand U5054 (N_5054,N_2940,N_1512);
nand U5055 (N_5055,N_1284,N_2818);
and U5056 (N_5056,N_731,N_1486);
nand U5057 (N_5057,N_2665,N_210);
or U5058 (N_5058,N_2074,N_1819);
nor U5059 (N_5059,N_1477,N_1942);
nand U5060 (N_5060,N_2006,N_648);
or U5061 (N_5061,N_2133,N_2585);
and U5062 (N_5062,N_783,N_62);
nand U5063 (N_5063,N_1427,N_2253);
and U5064 (N_5064,N_1449,N_2438);
or U5065 (N_5065,N_956,N_2418);
nand U5066 (N_5066,N_242,N_1125);
or U5067 (N_5067,N_62,N_1466);
and U5068 (N_5068,N_2495,N_1277);
nor U5069 (N_5069,N_2691,N_2240);
and U5070 (N_5070,N_656,N_2773);
and U5071 (N_5071,N_1623,N_768);
nor U5072 (N_5072,N_1991,N_2706);
and U5073 (N_5073,N_2426,N_1049);
nor U5074 (N_5074,N_2942,N_670);
and U5075 (N_5075,N_502,N_2013);
and U5076 (N_5076,N_2534,N_1082);
nand U5077 (N_5077,N_1182,N_1618);
and U5078 (N_5078,N_1741,N_1914);
nand U5079 (N_5079,N_1126,N_2358);
nor U5080 (N_5080,N_271,N_2215);
and U5081 (N_5081,N_1825,N_180);
nand U5082 (N_5082,N_1052,N_1567);
or U5083 (N_5083,N_780,N_1352);
or U5084 (N_5084,N_2112,N_1658);
nand U5085 (N_5085,N_464,N_1644);
and U5086 (N_5086,N_1653,N_1482);
and U5087 (N_5087,N_2236,N_1881);
or U5088 (N_5088,N_1527,N_181);
nor U5089 (N_5089,N_334,N_2919);
xor U5090 (N_5090,N_1723,N_1390);
xor U5091 (N_5091,N_1746,N_2414);
and U5092 (N_5092,N_2255,N_2548);
or U5093 (N_5093,N_233,N_505);
nand U5094 (N_5094,N_709,N_1821);
and U5095 (N_5095,N_144,N_1415);
or U5096 (N_5096,N_2322,N_763);
or U5097 (N_5097,N_1006,N_495);
nand U5098 (N_5098,N_677,N_2594);
nand U5099 (N_5099,N_1868,N_772);
nor U5100 (N_5100,N_2471,N_659);
and U5101 (N_5101,N_1852,N_2209);
nand U5102 (N_5102,N_2175,N_2930);
or U5103 (N_5103,N_1648,N_191);
nor U5104 (N_5104,N_1417,N_907);
nand U5105 (N_5105,N_1520,N_376);
and U5106 (N_5106,N_1384,N_707);
nor U5107 (N_5107,N_1709,N_1229);
nand U5108 (N_5108,N_1549,N_471);
nand U5109 (N_5109,N_1419,N_1199);
or U5110 (N_5110,N_1074,N_1980);
and U5111 (N_5111,N_823,N_1053);
nand U5112 (N_5112,N_2324,N_594);
and U5113 (N_5113,N_2970,N_1583);
or U5114 (N_5114,N_1567,N_497);
or U5115 (N_5115,N_1009,N_2431);
and U5116 (N_5116,N_915,N_1796);
xor U5117 (N_5117,N_1098,N_1335);
or U5118 (N_5118,N_2920,N_18);
nand U5119 (N_5119,N_2437,N_2143);
nor U5120 (N_5120,N_1398,N_1658);
nand U5121 (N_5121,N_253,N_2837);
nor U5122 (N_5122,N_84,N_2386);
or U5123 (N_5123,N_2591,N_1720);
nor U5124 (N_5124,N_2721,N_1414);
or U5125 (N_5125,N_1790,N_2823);
xor U5126 (N_5126,N_1564,N_1619);
or U5127 (N_5127,N_1657,N_2160);
xnor U5128 (N_5128,N_933,N_1743);
nor U5129 (N_5129,N_1520,N_2597);
nor U5130 (N_5130,N_344,N_2593);
nor U5131 (N_5131,N_313,N_836);
nor U5132 (N_5132,N_1342,N_687);
nand U5133 (N_5133,N_2144,N_502);
and U5134 (N_5134,N_1359,N_1200);
xor U5135 (N_5135,N_1538,N_156);
nor U5136 (N_5136,N_950,N_370);
nor U5137 (N_5137,N_990,N_1951);
or U5138 (N_5138,N_703,N_2914);
or U5139 (N_5139,N_2558,N_1102);
nor U5140 (N_5140,N_2839,N_530);
and U5141 (N_5141,N_2168,N_778);
nand U5142 (N_5142,N_1127,N_1636);
nor U5143 (N_5143,N_1586,N_959);
nor U5144 (N_5144,N_1478,N_2589);
or U5145 (N_5145,N_2853,N_1816);
and U5146 (N_5146,N_1333,N_621);
or U5147 (N_5147,N_2676,N_1220);
nor U5148 (N_5148,N_1040,N_2214);
or U5149 (N_5149,N_2789,N_1516);
xnor U5150 (N_5150,N_856,N_2231);
nand U5151 (N_5151,N_2499,N_1919);
nand U5152 (N_5152,N_2700,N_480);
and U5153 (N_5153,N_1363,N_2196);
or U5154 (N_5154,N_1937,N_2067);
or U5155 (N_5155,N_443,N_1794);
and U5156 (N_5156,N_584,N_1501);
or U5157 (N_5157,N_556,N_2216);
xor U5158 (N_5158,N_1583,N_384);
nand U5159 (N_5159,N_580,N_642);
xnor U5160 (N_5160,N_960,N_1340);
nand U5161 (N_5161,N_2313,N_887);
nor U5162 (N_5162,N_1346,N_926);
nand U5163 (N_5163,N_567,N_1645);
and U5164 (N_5164,N_263,N_204);
and U5165 (N_5165,N_334,N_234);
or U5166 (N_5166,N_721,N_672);
and U5167 (N_5167,N_323,N_2137);
nor U5168 (N_5168,N_2973,N_1609);
nor U5169 (N_5169,N_1023,N_2000);
nand U5170 (N_5170,N_2319,N_985);
and U5171 (N_5171,N_2567,N_1768);
nand U5172 (N_5172,N_351,N_2415);
or U5173 (N_5173,N_446,N_610);
or U5174 (N_5174,N_152,N_2563);
or U5175 (N_5175,N_1007,N_1077);
and U5176 (N_5176,N_737,N_1410);
nand U5177 (N_5177,N_2416,N_2290);
and U5178 (N_5178,N_306,N_1938);
xor U5179 (N_5179,N_1913,N_1544);
nand U5180 (N_5180,N_2802,N_950);
nor U5181 (N_5181,N_846,N_893);
nand U5182 (N_5182,N_759,N_2838);
nand U5183 (N_5183,N_1092,N_604);
nand U5184 (N_5184,N_367,N_30);
or U5185 (N_5185,N_1327,N_218);
nor U5186 (N_5186,N_689,N_984);
nor U5187 (N_5187,N_2654,N_2514);
nor U5188 (N_5188,N_1226,N_2620);
or U5189 (N_5189,N_949,N_1658);
or U5190 (N_5190,N_463,N_417);
and U5191 (N_5191,N_646,N_256);
or U5192 (N_5192,N_2259,N_1421);
or U5193 (N_5193,N_966,N_223);
nor U5194 (N_5194,N_2580,N_269);
nand U5195 (N_5195,N_2984,N_1593);
or U5196 (N_5196,N_1441,N_2303);
nand U5197 (N_5197,N_1294,N_954);
or U5198 (N_5198,N_1713,N_471);
or U5199 (N_5199,N_692,N_1696);
nand U5200 (N_5200,N_523,N_1667);
nand U5201 (N_5201,N_2950,N_293);
or U5202 (N_5202,N_546,N_2376);
xor U5203 (N_5203,N_296,N_1295);
xor U5204 (N_5204,N_1416,N_1849);
xor U5205 (N_5205,N_970,N_444);
nor U5206 (N_5206,N_1685,N_7);
nor U5207 (N_5207,N_665,N_1969);
nor U5208 (N_5208,N_545,N_673);
nand U5209 (N_5209,N_180,N_234);
and U5210 (N_5210,N_2534,N_2925);
or U5211 (N_5211,N_78,N_607);
or U5212 (N_5212,N_2533,N_467);
nand U5213 (N_5213,N_0,N_605);
or U5214 (N_5214,N_1087,N_281);
or U5215 (N_5215,N_398,N_1915);
nor U5216 (N_5216,N_873,N_744);
and U5217 (N_5217,N_2638,N_2586);
nor U5218 (N_5218,N_2287,N_2092);
xor U5219 (N_5219,N_1230,N_1491);
or U5220 (N_5220,N_1891,N_1939);
nor U5221 (N_5221,N_1016,N_2545);
or U5222 (N_5222,N_2740,N_2294);
xnor U5223 (N_5223,N_1386,N_2925);
nand U5224 (N_5224,N_261,N_2229);
and U5225 (N_5225,N_2303,N_1549);
and U5226 (N_5226,N_1690,N_2462);
nor U5227 (N_5227,N_1748,N_673);
and U5228 (N_5228,N_2217,N_1220);
and U5229 (N_5229,N_1623,N_2781);
xnor U5230 (N_5230,N_1851,N_1822);
or U5231 (N_5231,N_264,N_222);
xnor U5232 (N_5232,N_1771,N_144);
xnor U5233 (N_5233,N_715,N_10);
or U5234 (N_5234,N_790,N_2887);
or U5235 (N_5235,N_2512,N_624);
xnor U5236 (N_5236,N_1792,N_1289);
nand U5237 (N_5237,N_521,N_2204);
nand U5238 (N_5238,N_753,N_36);
or U5239 (N_5239,N_1419,N_2637);
nand U5240 (N_5240,N_2561,N_2383);
nand U5241 (N_5241,N_720,N_112);
nor U5242 (N_5242,N_328,N_1977);
and U5243 (N_5243,N_978,N_2369);
nor U5244 (N_5244,N_827,N_1067);
nand U5245 (N_5245,N_941,N_1027);
or U5246 (N_5246,N_1539,N_2528);
and U5247 (N_5247,N_971,N_1401);
nor U5248 (N_5248,N_423,N_2195);
nand U5249 (N_5249,N_2876,N_2013);
or U5250 (N_5250,N_1621,N_1364);
nor U5251 (N_5251,N_2473,N_412);
or U5252 (N_5252,N_2809,N_2741);
nor U5253 (N_5253,N_2547,N_837);
nand U5254 (N_5254,N_2228,N_164);
or U5255 (N_5255,N_637,N_721);
and U5256 (N_5256,N_2204,N_1971);
xnor U5257 (N_5257,N_1099,N_2641);
and U5258 (N_5258,N_2839,N_2625);
xnor U5259 (N_5259,N_1098,N_1698);
or U5260 (N_5260,N_1742,N_1513);
xnor U5261 (N_5261,N_745,N_394);
nor U5262 (N_5262,N_381,N_1060);
or U5263 (N_5263,N_1522,N_2113);
or U5264 (N_5264,N_490,N_2605);
nor U5265 (N_5265,N_885,N_341);
or U5266 (N_5266,N_393,N_2658);
nand U5267 (N_5267,N_1706,N_2397);
and U5268 (N_5268,N_2190,N_2520);
nand U5269 (N_5269,N_556,N_2993);
xor U5270 (N_5270,N_1392,N_117);
and U5271 (N_5271,N_2690,N_2346);
or U5272 (N_5272,N_651,N_1533);
or U5273 (N_5273,N_2030,N_1392);
nand U5274 (N_5274,N_2291,N_1744);
or U5275 (N_5275,N_2323,N_508);
or U5276 (N_5276,N_90,N_303);
or U5277 (N_5277,N_1106,N_2942);
nor U5278 (N_5278,N_547,N_1625);
and U5279 (N_5279,N_802,N_2783);
and U5280 (N_5280,N_1788,N_1851);
nand U5281 (N_5281,N_1603,N_1279);
nor U5282 (N_5282,N_1011,N_122);
nor U5283 (N_5283,N_1869,N_1079);
and U5284 (N_5284,N_2480,N_1342);
xnor U5285 (N_5285,N_1742,N_505);
or U5286 (N_5286,N_1241,N_1355);
and U5287 (N_5287,N_1785,N_2330);
xnor U5288 (N_5288,N_1049,N_2329);
or U5289 (N_5289,N_212,N_383);
and U5290 (N_5290,N_1777,N_2427);
and U5291 (N_5291,N_1303,N_1447);
and U5292 (N_5292,N_879,N_164);
and U5293 (N_5293,N_2200,N_479);
nor U5294 (N_5294,N_2008,N_750);
and U5295 (N_5295,N_2260,N_2728);
and U5296 (N_5296,N_2003,N_2135);
nor U5297 (N_5297,N_1943,N_2235);
nand U5298 (N_5298,N_989,N_2725);
or U5299 (N_5299,N_927,N_2473);
or U5300 (N_5300,N_2099,N_973);
nand U5301 (N_5301,N_2789,N_1152);
and U5302 (N_5302,N_1410,N_1572);
nor U5303 (N_5303,N_2508,N_2884);
and U5304 (N_5304,N_595,N_2709);
nand U5305 (N_5305,N_298,N_164);
nor U5306 (N_5306,N_700,N_306);
nand U5307 (N_5307,N_2629,N_1229);
and U5308 (N_5308,N_1423,N_504);
nor U5309 (N_5309,N_691,N_966);
nor U5310 (N_5310,N_1557,N_37);
nand U5311 (N_5311,N_2194,N_105);
nor U5312 (N_5312,N_2629,N_2141);
or U5313 (N_5313,N_546,N_2470);
and U5314 (N_5314,N_2935,N_2298);
xnor U5315 (N_5315,N_633,N_2856);
and U5316 (N_5316,N_1087,N_214);
nor U5317 (N_5317,N_1435,N_317);
or U5318 (N_5318,N_1791,N_669);
nand U5319 (N_5319,N_1354,N_281);
nand U5320 (N_5320,N_2680,N_684);
and U5321 (N_5321,N_2552,N_1737);
xor U5322 (N_5322,N_2245,N_2658);
or U5323 (N_5323,N_236,N_169);
nor U5324 (N_5324,N_1164,N_937);
nor U5325 (N_5325,N_2844,N_986);
or U5326 (N_5326,N_2433,N_602);
and U5327 (N_5327,N_649,N_1352);
or U5328 (N_5328,N_2864,N_2168);
nand U5329 (N_5329,N_2766,N_2865);
nor U5330 (N_5330,N_1622,N_1795);
and U5331 (N_5331,N_1122,N_1537);
nand U5332 (N_5332,N_1513,N_186);
and U5333 (N_5333,N_1422,N_131);
nor U5334 (N_5334,N_25,N_2282);
or U5335 (N_5335,N_496,N_2604);
nor U5336 (N_5336,N_498,N_2901);
xor U5337 (N_5337,N_1081,N_2151);
and U5338 (N_5338,N_1525,N_856);
nand U5339 (N_5339,N_2536,N_759);
nor U5340 (N_5340,N_2771,N_323);
nand U5341 (N_5341,N_1862,N_2602);
or U5342 (N_5342,N_1926,N_453);
nor U5343 (N_5343,N_906,N_741);
and U5344 (N_5344,N_2100,N_931);
and U5345 (N_5345,N_2833,N_1934);
nor U5346 (N_5346,N_1347,N_1089);
nand U5347 (N_5347,N_1850,N_1437);
or U5348 (N_5348,N_2977,N_52);
xnor U5349 (N_5349,N_2365,N_109);
and U5350 (N_5350,N_1478,N_1085);
or U5351 (N_5351,N_1425,N_2966);
xnor U5352 (N_5352,N_2421,N_1227);
xnor U5353 (N_5353,N_99,N_1467);
or U5354 (N_5354,N_1022,N_1548);
nor U5355 (N_5355,N_1854,N_20);
or U5356 (N_5356,N_114,N_1481);
xor U5357 (N_5357,N_1513,N_2853);
and U5358 (N_5358,N_1125,N_2032);
xnor U5359 (N_5359,N_422,N_624);
nand U5360 (N_5360,N_484,N_2547);
nor U5361 (N_5361,N_2379,N_2403);
nand U5362 (N_5362,N_1413,N_577);
and U5363 (N_5363,N_2616,N_1580);
or U5364 (N_5364,N_2185,N_1630);
or U5365 (N_5365,N_257,N_1896);
nor U5366 (N_5366,N_1381,N_264);
and U5367 (N_5367,N_2108,N_2797);
nand U5368 (N_5368,N_1966,N_1535);
nor U5369 (N_5369,N_2433,N_1171);
nand U5370 (N_5370,N_1347,N_2183);
or U5371 (N_5371,N_1014,N_2663);
nand U5372 (N_5372,N_430,N_1752);
nand U5373 (N_5373,N_1801,N_907);
nand U5374 (N_5374,N_2256,N_327);
and U5375 (N_5375,N_1375,N_330);
or U5376 (N_5376,N_287,N_2470);
nand U5377 (N_5377,N_1063,N_1076);
or U5378 (N_5378,N_732,N_75);
nor U5379 (N_5379,N_2309,N_2207);
and U5380 (N_5380,N_1149,N_1831);
or U5381 (N_5381,N_499,N_2765);
and U5382 (N_5382,N_1228,N_205);
nand U5383 (N_5383,N_438,N_1396);
and U5384 (N_5384,N_2538,N_2142);
nand U5385 (N_5385,N_2850,N_1556);
nand U5386 (N_5386,N_2284,N_808);
and U5387 (N_5387,N_727,N_2463);
or U5388 (N_5388,N_636,N_2940);
xor U5389 (N_5389,N_398,N_2257);
or U5390 (N_5390,N_715,N_535);
and U5391 (N_5391,N_897,N_2527);
nor U5392 (N_5392,N_1127,N_625);
nor U5393 (N_5393,N_551,N_580);
nor U5394 (N_5394,N_2862,N_30);
nand U5395 (N_5395,N_2268,N_925);
nor U5396 (N_5396,N_662,N_273);
nor U5397 (N_5397,N_1592,N_738);
nor U5398 (N_5398,N_1922,N_668);
xor U5399 (N_5399,N_1932,N_1504);
nor U5400 (N_5400,N_1205,N_2006);
nor U5401 (N_5401,N_1653,N_939);
xor U5402 (N_5402,N_915,N_2778);
or U5403 (N_5403,N_1078,N_1796);
nor U5404 (N_5404,N_1777,N_487);
or U5405 (N_5405,N_2820,N_658);
or U5406 (N_5406,N_751,N_600);
nand U5407 (N_5407,N_388,N_2197);
or U5408 (N_5408,N_2637,N_1631);
or U5409 (N_5409,N_2900,N_1977);
nand U5410 (N_5410,N_606,N_166);
nand U5411 (N_5411,N_1389,N_2395);
and U5412 (N_5412,N_1193,N_2129);
and U5413 (N_5413,N_608,N_870);
nand U5414 (N_5414,N_1650,N_1381);
nor U5415 (N_5415,N_1502,N_2992);
or U5416 (N_5416,N_187,N_1283);
and U5417 (N_5417,N_2551,N_2045);
and U5418 (N_5418,N_2279,N_2746);
xnor U5419 (N_5419,N_1618,N_106);
nand U5420 (N_5420,N_1356,N_1253);
nor U5421 (N_5421,N_825,N_1278);
or U5422 (N_5422,N_2232,N_338);
nand U5423 (N_5423,N_547,N_376);
xor U5424 (N_5424,N_2224,N_2179);
nand U5425 (N_5425,N_2772,N_2312);
or U5426 (N_5426,N_1129,N_290);
nand U5427 (N_5427,N_213,N_1773);
or U5428 (N_5428,N_2973,N_2411);
nor U5429 (N_5429,N_2997,N_1442);
and U5430 (N_5430,N_1616,N_2749);
and U5431 (N_5431,N_289,N_1334);
nor U5432 (N_5432,N_1235,N_2144);
and U5433 (N_5433,N_1010,N_14);
and U5434 (N_5434,N_2088,N_914);
nor U5435 (N_5435,N_1897,N_917);
nor U5436 (N_5436,N_901,N_2822);
or U5437 (N_5437,N_1909,N_1654);
nor U5438 (N_5438,N_144,N_472);
nor U5439 (N_5439,N_434,N_2537);
nor U5440 (N_5440,N_63,N_1195);
nor U5441 (N_5441,N_2307,N_1768);
and U5442 (N_5442,N_2264,N_2996);
nand U5443 (N_5443,N_160,N_2014);
or U5444 (N_5444,N_1229,N_695);
or U5445 (N_5445,N_2205,N_2221);
and U5446 (N_5446,N_1474,N_995);
or U5447 (N_5447,N_916,N_2921);
nand U5448 (N_5448,N_807,N_2201);
nor U5449 (N_5449,N_2798,N_1016);
nor U5450 (N_5450,N_1536,N_1936);
or U5451 (N_5451,N_980,N_2204);
nor U5452 (N_5452,N_850,N_155);
nor U5453 (N_5453,N_1617,N_2146);
nor U5454 (N_5454,N_2177,N_2894);
nand U5455 (N_5455,N_60,N_408);
nand U5456 (N_5456,N_2971,N_1840);
xor U5457 (N_5457,N_1950,N_2732);
nand U5458 (N_5458,N_254,N_1247);
and U5459 (N_5459,N_47,N_1261);
nor U5460 (N_5460,N_950,N_415);
nor U5461 (N_5461,N_1629,N_2437);
or U5462 (N_5462,N_0,N_1994);
xor U5463 (N_5463,N_2854,N_1926);
nor U5464 (N_5464,N_2626,N_1873);
and U5465 (N_5465,N_682,N_2319);
nand U5466 (N_5466,N_702,N_2318);
or U5467 (N_5467,N_1623,N_1226);
or U5468 (N_5468,N_1727,N_1666);
nor U5469 (N_5469,N_926,N_348);
nor U5470 (N_5470,N_1936,N_1609);
and U5471 (N_5471,N_897,N_2370);
and U5472 (N_5472,N_388,N_1795);
nand U5473 (N_5473,N_13,N_489);
and U5474 (N_5474,N_2224,N_429);
nor U5475 (N_5475,N_2645,N_1705);
nand U5476 (N_5476,N_1439,N_1401);
or U5477 (N_5477,N_809,N_457);
xnor U5478 (N_5478,N_650,N_2227);
xor U5479 (N_5479,N_2685,N_1117);
nand U5480 (N_5480,N_94,N_2423);
nor U5481 (N_5481,N_693,N_1223);
nor U5482 (N_5482,N_2097,N_1707);
nand U5483 (N_5483,N_2561,N_1771);
and U5484 (N_5484,N_1370,N_2367);
and U5485 (N_5485,N_151,N_1224);
and U5486 (N_5486,N_2758,N_1828);
nand U5487 (N_5487,N_1549,N_1957);
nor U5488 (N_5488,N_2259,N_1333);
xor U5489 (N_5489,N_739,N_2247);
or U5490 (N_5490,N_724,N_1164);
or U5491 (N_5491,N_723,N_2866);
nor U5492 (N_5492,N_2985,N_960);
and U5493 (N_5493,N_2197,N_1735);
nand U5494 (N_5494,N_67,N_185);
and U5495 (N_5495,N_2038,N_2976);
nand U5496 (N_5496,N_826,N_2773);
or U5497 (N_5497,N_612,N_981);
or U5498 (N_5498,N_724,N_974);
and U5499 (N_5499,N_806,N_1900);
nand U5500 (N_5500,N_546,N_2889);
nand U5501 (N_5501,N_1975,N_916);
and U5502 (N_5502,N_757,N_690);
or U5503 (N_5503,N_2952,N_2345);
or U5504 (N_5504,N_2453,N_1193);
and U5505 (N_5505,N_1570,N_2809);
or U5506 (N_5506,N_177,N_2727);
or U5507 (N_5507,N_1971,N_593);
and U5508 (N_5508,N_915,N_2031);
nand U5509 (N_5509,N_745,N_2094);
nand U5510 (N_5510,N_1993,N_516);
nand U5511 (N_5511,N_1297,N_2521);
and U5512 (N_5512,N_2498,N_785);
nor U5513 (N_5513,N_350,N_1672);
and U5514 (N_5514,N_2614,N_659);
nand U5515 (N_5515,N_363,N_103);
nor U5516 (N_5516,N_2494,N_770);
and U5517 (N_5517,N_559,N_2220);
nand U5518 (N_5518,N_1210,N_969);
and U5519 (N_5519,N_2151,N_160);
or U5520 (N_5520,N_1494,N_286);
and U5521 (N_5521,N_1209,N_1038);
or U5522 (N_5522,N_1681,N_1805);
nand U5523 (N_5523,N_2990,N_2);
or U5524 (N_5524,N_2190,N_606);
or U5525 (N_5525,N_1538,N_2810);
or U5526 (N_5526,N_2005,N_1062);
nor U5527 (N_5527,N_840,N_2573);
nand U5528 (N_5528,N_2663,N_2436);
or U5529 (N_5529,N_1022,N_227);
nor U5530 (N_5530,N_1673,N_1248);
and U5531 (N_5531,N_1760,N_1665);
nor U5532 (N_5532,N_814,N_2837);
or U5533 (N_5533,N_2649,N_2372);
and U5534 (N_5534,N_1766,N_2268);
xnor U5535 (N_5535,N_468,N_2752);
nor U5536 (N_5536,N_1328,N_331);
nor U5537 (N_5537,N_2442,N_2669);
and U5538 (N_5538,N_2864,N_526);
and U5539 (N_5539,N_877,N_430);
nor U5540 (N_5540,N_2342,N_850);
and U5541 (N_5541,N_2825,N_1392);
nor U5542 (N_5542,N_2742,N_180);
nor U5543 (N_5543,N_177,N_2988);
nor U5544 (N_5544,N_863,N_718);
nand U5545 (N_5545,N_1778,N_286);
nand U5546 (N_5546,N_2289,N_1211);
nand U5547 (N_5547,N_2231,N_1415);
and U5548 (N_5548,N_403,N_1946);
xor U5549 (N_5549,N_923,N_2958);
nand U5550 (N_5550,N_1364,N_1935);
or U5551 (N_5551,N_647,N_1589);
or U5552 (N_5552,N_926,N_1139);
or U5553 (N_5553,N_235,N_2250);
and U5554 (N_5554,N_987,N_2486);
or U5555 (N_5555,N_1297,N_886);
xnor U5556 (N_5556,N_371,N_667);
or U5557 (N_5557,N_963,N_1052);
or U5558 (N_5558,N_1343,N_1179);
nor U5559 (N_5559,N_397,N_1378);
and U5560 (N_5560,N_2555,N_1842);
and U5561 (N_5561,N_2540,N_996);
nand U5562 (N_5562,N_1011,N_2125);
and U5563 (N_5563,N_1709,N_2230);
and U5564 (N_5564,N_2377,N_1151);
nor U5565 (N_5565,N_622,N_1368);
or U5566 (N_5566,N_2286,N_2900);
nor U5567 (N_5567,N_1847,N_2524);
or U5568 (N_5568,N_1110,N_246);
xnor U5569 (N_5569,N_1288,N_2726);
and U5570 (N_5570,N_2157,N_710);
or U5571 (N_5571,N_708,N_1247);
and U5572 (N_5572,N_2594,N_858);
or U5573 (N_5573,N_1610,N_439);
and U5574 (N_5574,N_2201,N_1413);
or U5575 (N_5575,N_776,N_438);
and U5576 (N_5576,N_1374,N_2463);
xnor U5577 (N_5577,N_1024,N_1467);
nor U5578 (N_5578,N_1670,N_2452);
nor U5579 (N_5579,N_1460,N_703);
nor U5580 (N_5580,N_852,N_2544);
nor U5581 (N_5581,N_2569,N_1974);
and U5582 (N_5582,N_1552,N_1513);
or U5583 (N_5583,N_1725,N_1974);
nand U5584 (N_5584,N_1388,N_483);
nor U5585 (N_5585,N_2831,N_1928);
or U5586 (N_5586,N_1084,N_29);
nor U5587 (N_5587,N_242,N_924);
nand U5588 (N_5588,N_2699,N_340);
and U5589 (N_5589,N_1157,N_120);
or U5590 (N_5590,N_207,N_2420);
and U5591 (N_5591,N_1248,N_1175);
or U5592 (N_5592,N_1476,N_2818);
nor U5593 (N_5593,N_2459,N_1788);
nand U5594 (N_5594,N_1719,N_1072);
xor U5595 (N_5595,N_2661,N_2079);
nand U5596 (N_5596,N_100,N_2309);
nor U5597 (N_5597,N_1377,N_1240);
nor U5598 (N_5598,N_2858,N_889);
nor U5599 (N_5599,N_391,N_2504);
or U5600 (N_5600,N_2966,N_1662);
nor U5601 (N_5601,N_2393,N_158);
xor U5602 (N_5602,N_487,N_1392);
nor U5603 (N_5603,N_1455,N_2002);
or U5604 (N_5604,N_126,N_2156);
nand U5605 (N_5605,N_1866,N_544);
or U5606 (N_5606,N_1431,N_536);
and U5607 (N_5607,N_958,N_350);
and U5608 (N_5608,N_1915,N_1648);
or U5609 (N_5609,N_1008,N_532);
and U5610 (N_5610,N_785,N_2513);
nor U5611 (N_5611,N_2504,N_1214);
nor U5612 (N_5612,N_2824,N_1684);
or U5613 (N_5613,N_1511,N_851);
nor U5614 (N_5614,N_606,N_532);
or U5615 (N_5615,N_739,N_281);
or U5616 (N_5616,N_1993,N_2120);
or U5617 (N_5617,N_821,N_841);
and U5618 (N_5618,N_1396,N_1043);
nand U5619 (N_5619,N_2621,N_1875);
or U5620 (N_5620,N_1339,N_1784);
nor U5621 (N_5621,N_1402,N_2758);
or U5622 (N_5622,N_659,N_2035);
or U5623 (N_5623,N_2679,N_1743);
and U5624 (N_5624,N_923,N_1609);
nor U5625 (N_5625,N_1373,N_719);
nor U5626 (N_5626,N_416,N_1098);
nor U5627 (N_5627,N_1598,N_796);
or U5628 (N_5628,N_1011,N_2121);
and U5629 (N_5629,N_297,N_2700);
or U5630 (N_5630,N_2953,N_801);
or U5631 (N_5631,N_133,N_2685);
nand U5632 (N_5632,N_1203,N_1807);
and U5633 (N_5633,N_2897,N_2109);
nand U5634 (N_5634,N_2165,N_2354);
nor U5635 (N_5635,N_2505,N_1999);
nand U5636 (N_5636,N_1298,N_1587);
nand U5637 (N_5637,N_1786,N_400);
xnor U5638 (N_5638,N_2765,N_2435);
and U5639 (N_5639,N_1704,N_2945);
xnor U5640 (N_5640,N_1443,N_1183);
or U5641 (N_5641,N_950,N_2838);
nor U5642 (N_5642,N_2732,N_912);
or U5643 (N_5643,N_2785,N_599);
nand U5644 (N_5644,N_2990,N_2125);
or U5645 (N_5645,N_1158,N_1164);
xnor U5646 (N_5646,N_1284,N_2771);
or U5647 (N_5647,N_2741,N_640);
or U5648 (N_5648,N_282,N_294);
nor U5649 (N_5649,N_814,N_1289);
or U5650 (N_5650,N_766,N_2384);
or U5651 (N_5651,N_2345,N_1658);
nor U5652 (N_5652,N_1872,N_44);
nor U5653 (N_5653,N_1845,N_1561);
nor U5654 (N_5654,N_2237,N_2555);
and U5655 (N_5655,N_1506,N_208);
nor U5656 (N_5656,N_2523,N_421);
nand U5657 (N_5657,N_1177,N_356);
nor U5658 (N_5658,N_2449,N_2975);
nor U5659 (N_5659,N_885,N_2664);
nor U5660 (N_5660,N_2000,N_358);
and U5661 (N_5661,N_2853,N_434);
nor U5662 (N_5662,N_1427,N_1738);
nor U5663 (N_5663,N_1236,N_183);
nand U5664 (N_5664,N_963,N_830);
nand U5665 (N_5665,N_794,N_83);
nor U5666 (N_5666,N_399,N_123);
nand U5667 (N_5667,N_2878,N_2679);
and U5668 (N_5668,N_1384,N_1485);
or U5669 (N_5669,N_1895,N_158);
or U5670 (N_5670,N_1762,N_1462);
xnor U5671 (N_5671,N_535,N_34);
xnor U5672 (N_5672,N_2446,N_2074);
or U5673 (N_5673,N_1550,N_2187);
and U5674 (N_5674,N_1590,N_2137);
xnor U5675 (N_5675,N_368,N_2835);
xor U5676 (N_5676,N_1865,N_534);
nand U5677 (N_5677,N_619,N_2340);
xnor U5678 (N_5678,N_1877,N_2725);
and U5679 (N_5679,N_2050,N_433);
nor U5680 (N_5680,N_2031,N_376);
or U5681 (N_5681,N_2320,N_282);
nand U5682 (N_5682,N_1004,N_1763);
nor U5683 (N_5683,N_2253,N_2908);
and U5684 (N_5684,N_1822,N_2300);
xor U5685 (N_5685,N_2480,N_890);
nor U5686 (N_5686,N_2982,N_1411);
and U5687 (N_5687,N_841,N_1042);
nor U5688 (N_5688,N_2669,N_105);
or U5689 (N_5689,N_1845,N_524);
nor U5690 (N_5690,N_1969,N_2360);
nor U5691 (N_5691,N_2860,N_1051);
or U5692 (N_5692,N_1567,N_652);
nor U5693 (N_5693,N_2797,N_597);
and U5694 (N_5694,N_2059,N_161);
and U5695 (N_5695,N_447,N_2926);
nand U5696 (N_5696,N_2648,N_1125);
or U5697 (N_5697,N_1623,N_2176);
and U5698 (N_5698,N_2786,N_1913);
xor U5699 (N_5699,N_771,N_2432);
nor U5700 (N_5700,N_661,N_1329);
and U5701 (N_5701,N_832,N_481);
nor U5702 (N_5702,N_1808,N_2145);
or U5703 (N_5703,N_2629,N_2857);
or U5704 (N_5704,N_1499,N_791);
and U5705 (N_5705,N_2615,N_250);
nand U5706 (N_5706,N_405,N_1328);
xnor U5707 (N_5707,N_290,N_1734);
nor U5708 (N_5708,N_2351,N_125);
and U5709 (N_5709,N_463,N_1412);
or U5710 (N_5710,N_204,N_1066);
and U5711 (N_5711,N_191,N_1408);
and U5712 (N_5712,N_1871,N_2221);
and U5713 (N_5713,N_885,N_751);
nor U5714 (N_5714,N_1483,N_2572);
nand U5715 (N_5715,N_2478,N_124);
nor U5716 (N_5716,N_2759,N_1349);
or U5717 (N_5717,N_1455,N_241);
nand U5718 (N_5718,N_2621,N_2006);
xor U5719 (N_5719,N_1167,N_2770);
nor U5720 (N_5720,N_93,N_2893);
nand U5721 (N_5721,N_363,N_2624);
and U5722 (N_5722,N_1172,N_2257);
or U5723 (N_5723,N_2252,N_1521);
nand U5724 (N_5724,N_2243,N_1212);
nand U5725 (N_5725,N_2108,N_2509);
and U5726 (N_5726,N_233,N_1943);
nand U5727 (N_5727,N_1043,N_1682);
and U5728 (N_5728,N_1718,N_2793);
nor U5729 (N_5729,N_2490,N_1484);
nand U5730 (N_5730,N_1034,N_2714);
xor U5731 (N_5731,N_2285,N_858);
or U5732 (N_5732,N_2905,N_2266);
or U5733 (N_5733,N_2855,N_687);
nor U5734 (N_5734,N_2880,N_673);
and U5735 (N_5735,N_2828,N_146);
or U5736 (N_5736,N_2515,N_2784);
and U5737 (N_5737,N_2339,N_661);
xor U5738 (N_5738,N_1352,N_1688);
and U5739 (N_5739,N_1455,N_1641);
xnor U5740 (N_5740,N_925,N_558);
or U5741 (N_5741,N_412,N_137);
xnor U5742 (N_5742,N_377,N_2824);
or U5743 (N_5743,N_1584,N_809);
xor U5744 (N_5744,N_1920,N_658);
and U5745 (N_5745,N_2981,N_118);
and U5746 (N_5746,N_1318,N_138);
nand U5747 (N_5747,N_1953,N_294);
and U5748 (N_5748,N_1256,N_2454);
nor U5749 (N_5749,N_657,N_1808);
nor U5750 (N_5750,N_60,N_1209);
and U5751 (N_5751,N_1167,N_2587);
and U5752 (N_5752,N_1188,N_1727);
or U5753 (N_5753,N_396,N_871);
and U5754 (N_5754,N_2370,N_2773);
and U5755 (N_5755,N_2768,N_447);
nand U5756 (N_5756,N_1913,N_1298);
or U5757 (N_5757,N_2482,N_94);
nor U5758 (N_5758,N_1771,N_2132);
xnor U5759 (N_5759,N_1557,N_2873);
nor U5760 (N_5760,N_1531,N_2802);
and U5761 (N_5761,N_2706,N_245);
and U5762 (N_5762,N_1730,N_1516);
and U5763 (N_5763,N_1736,N_443);
and U5764 (N_5764,N_493,N_2527);
nand U5765 (N_5765,N_1662,N_149);
nand U5766 (N_5766,N_1253,N_2005);
nor U5767 (N_5767,N_2369,N_2705);
or U5768 (N_5768,N_172,N_888);
xnor U5769 (N_5769,N_1638,N_2996);
nand U5770 (N_5770,N_2270,N_1299);
and U5771 (N_5771,N_24,N_1603);
nand U5772 (N_5772,N_1927,N_1571);
xnor U5773 (N_5773,N_786,N_1264);
nand U5774 (N_5774,N_719,N_1096);
nand U5775 (N_5775,N_1182,N_1172);
or U5776 (N_5776,N_2951,N_1710);
or U5777 (N_5777,N_1404,N_622);
nor U5778 (N_5778,N_2479,N_650);
nand U5779 (N_5779,N_917,N_2577);
or U5780 (N_5780,N_2026,N_2431);
xor U5781 (N_5781,N_533,N_2353);
nand U5782 (N_5782,N_1770,N_2317);
xor U5783 (N_5783,N_2301,N_2942);
nor U5784 (N_5784,N_2772,N_2276);
nand U5785 (N_5785,N_830,N_1725);
or U5786 (N_5786,N_2191,N_2639);
or U5787 (N_5787,N_2590,N_12);
and U5788 (N_5788,N_2532,N_770);
xnor U5789 (N_5789,N_2172,N_1773);
or U5790 (N_5790,N_979,N_2834);
nor U5791 (N_5791,N_2657,N_2517);
or U5792 (N_5792,N_413,N_190);
nand U5793 (N_5793,N_552,N_1466);
nand U5794 (N_5794,N_747,N_945);
and U5795 (N_5795,N_2636,N_2886);
xor U5796 (N_5796,N_17,N_2460);
and U5797 (N_5797,N_1150,N_1008);
nand U5798 (N_5798,N_2819,N_2847);
nor U5799 (N_5799,N_970,N_805);
nand U5800 (N_5800,N_2375,N_2518);
xor U5801 (N_5801,N_583,N_135);
nor U5802 (N_5802,N_979,N_205);
or U5803 (N_5803,N_368,N_2877);
xor U5804 (N_5804,N_1673,N_1954);
nand U5805 (N_5805,N_28,N_617);
and U5806 (N_5806,N_2316,N_272);
and U5807 (N_5807,N_2834,N_2633);
nor U5808 (N_5808,N_110,N_2393);
nor U5809 (N_5809,N_1331,N_333);
nand U5810 (N_5810,N_190,N_2744);
and U5811 (N_5811,N_1176,N_528);
and U5812 (N_5812,N_1223,N_2356);
and U5813 (N_5813,N_2353,N_1015);
or U5814 (N_5814,N_2790,N_920);
or U5815 (N_5815,N_2137,N_2860);
nand U5816 (N_5816,N_2467,N_2663);
or U5817 (N_5817,N_1477,N_2301);
or U5818 (N_5818,N_1121,N_1927);
nand U5819 (N_5819,N_2287,N_673);
nor U5820 (N_5820,N_1346,N_1500);
and U5821 (N_5821,N_2926,N_345);
nor U5822 (N_5822,N_1435,N_640);
nor U5823 (N_5823,N_1876,N_1096);
nand U5824 (N_5824,N_2198,N_325);
xnor U5825 (N_5825,N_641,N_658);
nand U5826 (N_5826,N_2048,N_2719);
nor U5827 (N_5827,N_1709,N_1633);
and U5828 (N_5828,N_1558,N_22);
and U5829 (N_5829,N_1072,N_572);
xnor U5830 (N_5830,N_1959,N_2757);
and U5831 (N_5831,N_963,N_1589);
or U5832 (N_5832,N_2875,N_2507);
nor U5833 (N_5833,N_1806,N_796);
or U5834 (N_5834,N_2370,N_2097);
nor U5835 (N_5835,N_2348,N_2044);
and U5836 (N_5836,N_2965,N_1583);
and U5837 (N_5837,N_2425,N_1009);
or U5838 (N_5838,N_1568,N_2147);
and U5839 (N_5839,N_538,N_1534);
nand U5840 (N_5840,N_1961,N_1551);
or U5841 (N_5841,N_56,N_2760);
nand U5842 (N_5842,N_2620,N_1208);
nand U5843 (N_5843,N_1945,N_1975);
nor U5844 (N_5844,N_1303,N_2544);
and U5845 (N_5845,N_672,N_231);
and U5846 (N_5846,N_336,N_641);
nand U5847 (N_5847,N_1900,N_1973);
xor U5848 (N_5848,N_1612,N_2579);
nor U5849 (N_5849,N_1823,N_561);
nand U5850 (N_5850,N_2077,N_2508);
xnor U5851 (N_5851,N_1695,N_1258);
nor U5852 (N_5852,N_245,N_1750);
and U5853 (N_5853,N_1350,N_1951);
nor U5854 (N_5854,N_2993,N_1527);
and U5855 (N_5855,N_781,N_2006);
and U5856 (N_5856,N_43,N_2963);
nand U5857 (N_5857,N_1131,N_1502);
and U5858 (N_5858,N_145,N_2238);
nand U5859 (N_5859,N_2964,N_1475);
and U5860 (N_5860,N_2686,N_1215);
nand U5861 (N_5861,N_757,N_598);
or U5862 (N_5862,N_1018,N_2510);
and U5863 (N_5863,N_2597,N_872);
and U5864 (N_5864,N_2956,N_1678);
xnor U5865 (N_5865,N_2338,N_1286);
and U5866 (N_5866,N_282,N_1261);
and U5867 (N_5867,N_2666,N_2472);
xnor U5868 (N_5868,N_2481,N_384);
or U5869 (N_5869,N_1546,N_810);
or U5870 (N_5870,N_785,N_703);
nand U5871 (N_5871,N_1778,N_2373);
xor U5872 (N_5872,N_236,N_1740);
and U5873 (N_5873,N_1831,N_1229);
and U5874 (N_5874,N_1555,N_892);
and U5875 (N_5875,N_2655,N_2874);
nor U5876 (N_5876,N_756,N_2871);
nor U5877 (N_5877,N_2172,N_2952);
nand U5878 (N_5878,N_2466,N_2917);
and U5879 (N_5879,N_1595,N_2205);
nand U5880 (N_5880,N_1285,N_42);
nand U5881 (N_5881,N_1041,N_2015);
xor U5882 (N_5882,N_2984,N_897);
and U5883 (N_5883,N_1266,N_2800);
nand U5884 (N_5884,N_948,N_2847);
or U5885 (N_5885,N_1253,N_446);
and U5886 (N_5886,N_2375,N_2629);
and U5887 (N_5887,N_302,N_1314);
xor U5888 (N_5888,N_1557,N_92);
and U5889 (N_5889,N_2260,N_1710);
xor U5890 (N_5890,N_1932,N_316);
nand U5891 (N_5891,N_1830,N_1054);
and U5892 (N_5892,N_446,N_762);
nand U5893 (N_5893,N_775,N_1463);
nor U5894 (N_5894,N_2382,N_582);
or U5895 (N_5895,N_1502,N_2442);
or U5896 (N_5896,N_492,N_973);
nor U5897 (N_5897,N_36,N_1784);
or U5898 (N_5898,N_2824,N_1657);
nor U5899 (N_5899,N_2091,N_2583);
nand U5900 (N_5900,N_533,N_144);
nand U5901 (N_5901,N_19,N_759);
nor U5902 (N_5902,N_318,N_2213);
or U5903 (N_5903,N_673,N_516);
nor U5904 (N_5904,N_1906,N_1108);
xnor U5905 (N_5905,N_2813,N_2862);
nor U5906 (N_5906,N_1980,N_2335);
nor U5907 (N_5907,N_583,N_1103);
and U5908 (N_5908,N_1727,N_745);
nor U5909 (N_5909,N_684,N_2036);
nand U5910 (N_5910,N_1403,N_1309);
xor U5911 (N_5911,N_1034,N_2509);
nand U5912 (N_5912,N_2096,N_748);
or U5913 (N_5913,N_36,N_1142);
nand U5914 (N_5914,N_2524,N_729);
and U5915 (N_5915,N_1081,N_819);
or U5916 (N_5916,N_1318,N_2232);
nor U5917 (N_5917,N_738,N_2032);
nor U5918 (N_5918,N_568,N_66);
nand U5919 (N_5919,N_1718,N_1560);
and U5920 (N_5920,N_2915,N_208);
nand U5921 (N_5921,N_1359,N_1994);
xnor U5922 (N_5922,N_218,N_1669);
nor U5923 (N_5923,N_2158,N_2858);
nand U5924 (N_5924,N_2536,N_957);
nor U5925 (N_5925,N_1971,N_2860);
or U5926 (N_5926,N_1752,N_808);
and U5927 (N_5927,N_1806,N_1497);
nand U5928 (N_5928,N_45,N_162);
and U5929 (N_5929,N_131,N_2152);
nand U5930 (N_5930,N_2358,N_932);
nor U5931 (N_5931,N_2467,N_367);
or U5932 (N_5932,N_1732,N_850);
nand U5933 (N_5933,N_2131,N_393);
nand U5934 (N_5934,N_629,N_2230);
or U5935 (N_5935,N_1765,N_2507);
or U5936 (N_5936,N_2296,N_2390);
and U5937 (N_5937,N_1251,N_1059);
xor U5938 (N_5938,N_2715,N_709);
and U5939 (N_5939,N_1553,N_2836);
nand U5940 (N_5940,N_1622,N_254);
nor U5941 (N_5941,N_466,N_860);
and U5942 (N_5942,N_385,N_984);
nand U5943 (N_5943,N_2034,N_2961);
and U5944 (N_5944,N_270,N_2436);
or U5945 (N_5945,N_1083,N_2727);
or U5946 (N_5946,N_702,N_476);
nand U5947 (N_5947,N_373,N_639);
or U5948 (N_5948,N_1991,N_2167);
and U5949 (N_5949,N_2990,N_676);
nor U5950 (N_5950,N_418,N_510);
nor U5951 (N_5951,N_1104,N_2122);
and U5952 (N_5952,N_965,N_2602);
and U5953 (N_5953,N_2133,N_310);
xor U5954 (N_5954,N_2282,N_2687);
and U5955 (N_5955,N_1768,N_620);
or U5956 (N_5956,N_2327,N_1618);
nand U5957 (N_5957,N_590,N_805);
or U5958 (N_5958,N_2781,N_1425);
or U5959 (N_5959,N_2014,N_418);
nor U5960 (N_5960,N_2048,N_2586);
and U5961 (N_5961,N_2123,N_1003);
nand U5962 (N_5962,N_1018,N_2169);
nor U5963 (N_5963,N_1691,N_618);
and U5964 (N_5964,N_1064,N_792);
or U5965 (N_5965,N_1338,N_2143);
or U5966 (N_5966,N_779,N_201);
nor U5967 (N_5967,N_2622,N_672);
nand U5968 (N_5968,N_1586,N_2041);
and U5969 (N_5969,N_2260,N_478);
and U5970 (N_5970,N_2203,N_517);
nand U5971 (N_5971,N_2936,N_2719);
nand U5972 (N_5972,N_1635,N_1226);
and U5973 (N_5973,N_206,N_1059);
xnor U5974 (N_5974,N_2476,N_2861);
nor U5975 (N_5975,N_1533,N_831);
or U5976 (N_5976,N_2505,N_2583);
and U5977 (N_5977,N_873,N_28);
nand U5978 (N_5978,N_385,N_957);
nor U5979 (N_5979,N_1247,N_1443);
or U5980 (N_5980,N_2502,N_1207);
nand U5981 (N_5981,N_1526,N_2306);
or U5982 (N_5982,N_456,N_1915);
nand U5983 (N_5983,N_540,N_1718);
nand U5984 (N_5984,N_644,N_1276);
xnor U5985 (N_5985,N_1553,N_1630);
nand U5986 (N_5986,N_1187,N_743);
nand U5987 (N_5987,N_294,N_2208);
and U5988 (N_5988,N_994,N_417);
xnor U5989 (N_5989,N_2380,N_2640);
nand U5990 (N_5990,N_359,N_1256);
nor U5991 (N_5991,N_464,N_1007);
and U5992 (N_5992,N_1405,N_2855);
nand U5993 (N_5993,N_1966,N_970);
nor U5994 (N_5994,N_313,N_1908);
or U5995 (N_5995,N_2143,N_102);
and U5996 (N_5996,N_1071,N_1163);
or U5997 (N_5997,N_2924,N_2540);
nand U5998 (N_5998,N_604,N_716);
nor U5999 (N_5999,N_1760,N_204);
and U6000 (N_6000,N_3326,N_3637);
xor U6001 (N_6001,N_4679,N_3478);
nor U6002 (N_6002,N_3633,N_3571);
or U6003 (N_6003,N_4578,N_5162);
nor U6004 (N_6004,N_4155,N_3759);
nand U6005 (N_6005,N_3573,N_5665);
nor U6006 (N_6006,N_4579,N_5553);
and U6007 (N_6007,N_5249,N_3232);
and U6008 (N_6008,N_3661,N_3163);
and U6009 (N_6009,N_3275,N_5779);
xor U6010 (N_6010,N_4939,N_3320);
and U6011 (N_6011,N_5936,N_3386);
nor U6012 (N_6012,N_5886,N_3952);
xor U6013 (N_6013,N_4322,N_5172);
and U6014 (N_6014,N_4933,N_4045);
and U6015 (N_6015,N_5550,N_4123);
or U6016 (N_6016,N_4079,N_4686);
and U6017 (N_6017,N_3156,N_4633);
nand U6018 (N_6018,N_5065,N_4273);
nand U6019 (N_6019,N_3070,N_5207);
nor U6020 (N_6020,N_3942,N_4543);
nand U6021 (N_6021,N_3984,N_5239);
nor U6022 (N_6022,N_4417,N_5658);
nand U6023 (N_6023,N_3592,N_5827);
nand U6024 (N_6024,N_3263,N_5090);
xnor U6025 (N_6025,N_5456,N_3498);
and U6026 (N_6026,N_4501,N_5606);
and U6027 (N_6027,N_5136,N_3417);
and U6028 (N_6028,N_3769,N_3814);
nor U6029 (N_6029,N_5119,N_3047);
nor U6030 (N_6030,N_4702,N_4326);
nand U6031 (N_6031,N_4335,N_3024);
nand U6032 (N_6032,N_5433,N_3338);
or U6033 (N_6033,N_3919,N_3424);
nand U6034 (N_6034,N_5714,N_3569);
and U6035 (N_6035,N_4877,N_3535);
nand U6036 (N_6036,N_3043,N_3651);
nand U6037 (N_6037,N_5648,N_5262);
nor U6038 (N_6038,N_5414,N_5156);
nor U6039 (N_6039,N_4650,N_3312);
nor U6040 (N_6040,N_4558,N_3574);
and U6041 (N_6041,N_3492,N_3887);
nor U6042 (N_6042,N_3961,N_3395);
xnor U6043 (N_6043,N_5727,N_3739);
nor U6044 (N_6044,N_5989,N_4762);
nand U6045 (N_6045,N_5890,N_4177);
or U6046 (N_6046,N_3844,N_5051);
or U6047 (N_6047,N_5612,N_5687);
and U6048 (N_6048,N_4860,N_5095);
nand U6049 (N_6049,N_4592,N_4420);
or U6050 (N_6050,N_4264,N_4638);
nand U6051 (N_6051,N_5318,N_5694);
and U6052 (N_6052,N_5463,N_5724);
nor U6053 (N_6053,N_3467,N_3257);
and U6054 (N_6054,N_4824,N_4365);
xor U6055 (N_6055,N_3223,N_5723);
nor U6056 (N_6056,N_3144,N_4913);
nor U6057 (N_6057,N_3458,N_3079);
and U6058 (N_6058,N_3974,N_3044);
or U6059 (N_6059,N_4173,N_5331);
and U6060 (N_6060,N_5880,N_3175);
nand U6061 (N_6061,N_5669,N_3512);
nor U6062 (N_6062,N_5001,N_5222);
and U6063 (N_6063,N_4338,N_4000);
or U6064 (N_6064,N_5767,N_5511);
nor U6065 (N_6065,N_5971,N_3048);
nor U6066 (N_6066,N_4904,N_5871);
nor U6067 (N_6067,N_5264,N_4965);
nand U6068 (N_6068,N_3322,N_5442);
nor U6069 (N_6069,N_3114,N_3815);
and U6070 (N_6070,N_4018,N_3051);
or U6071 (N_6071,N_3189,N_3210);
or U6072 (N_6072,N_5475,N_3034);
and U6073 (N_6073,N_3450,N_5309);
or U6074 (N_6074,N_5600,N_5234);
or U6075 (N_6075,N_3117,N_3828);
nor U6076 (N_6076,N_5226,N_4526);
nand U6077 (N_6077,N_5556,N_4493);
nand U6078 (N_6078,N_4059,N_5942);
xor U6079 (N_6079,N_3783,N_4183);
or U6080 (N_6080,N_3292,N_3726);
nand U6081 (N_6081,N_5028,N_3860);
or U6082 (N_6082,N_5684,N_3122);
nor U6083 (N_6083,N_3861,N_4185);
and U6084 (N_6084,N_5151,N_3001);
or U6085 (N_6085,N_3052,N_5220);
nor U6086 (N_6086,N_5899,N_3606);
nand U6087 (N_6087,N_4768,N_3266);
and U6088 (N_6088,N_5039,N_5465);
nand U6089 (N_6089,N_3853,N_3094);
nand U6090 (N_6090,N_5398,N_3293);
nand U6091 (N_6091,N_4828,N_5773);
nand U6092 (N_6092,N_3221,N_4424);
and U6093 (N_6093,N_3724,N_5063);
and U6094 (N_6094,N_3028,N_5733);
nor U6095 (N_6095,N_4942,N_5011);
nand U6096 (N_6096,N_4569,N_5225);
nand U6097 (N_6097,N_4363,N_5452);
or U6098 (N_6098,N_5980,N_5032);
nand U6099 (N_6099,N_5285,N_3566);
and U6100 (N_6100,N_4978,N_3323);
nor U6101 (N_6101,N_3626,N_4687);
and U6102 (N_6102,N_5029,N_5596);
or U6103 (N_6103,N_4149,N_5181);
or U6104 (N_6104,N_5924,N_3743);
and U6105 (N_6105,N_5143,N_5699);
nor U6106 (N_6106,N_5616,N_3063);
and U6107 (N_6107,N_5895,N_4980);
or U6108 (N_6108,N_4022,N_3826);
nand U6109 (N_6109,N_3180,N_4977);
nand U6110 (N_6110,N_3895,N_3434);
or U6111 (N_6111,N_4647,N_4253);
and U6112 (N_6112,N_4533,N_5732);
nor U6113 (N_6113,N_3238,N_3894);
or U6114 (N_6114,N_3858,N_4790);
or U6115 (N_6115,N_3857,N_5708);
or U6116 (N_6116,N_5251,N_5254);
nor U6117 (N_6117,N_4673,N_4994);
xor U6118 (N_6118,N_5988,N_3406);
xor U6119 (N_6119,N_4707,N_3225);
or U6120 (N_6120,N_3982,N_5903);
and U6121 (N_6121,N_3041,N_5843);
nand U6122 (N_6122,N_3521,N_4622);
nor U6123 (N_6123,N_4370,N_3937);
and U6124 (N_6124,N_4812,N_4236);
nand U6125 (N_6125,N_3009,N_4274);
nand U6126 (N_6126,N_3443,N_3883);
and U6127 (N_6127,N_4716,N_3598);
nor U6128 (N_6128,N_3357,N_5490);
and U6129 (N_6129,N_5084,N_5918);
nand U6130 (N_6130,N_3012,N_5628);
xor U6131 (N_6131,N_3704,N_4029);
or U6132 (N_6132,N_5337,N_4730);
and U6133 (N_6133,N_5009,N_3800);
nor U6134 (N_6134,N_4349,N_5963);
nor U6135 (N_6135,N_3004,N_3440);
and U6136 (N_6136,N_4785,N_5154);
or U6137 (N_6137,N_4864,N_4728);
nand U6138 (N_6138,N_4343,N_3855);
nor U6139 (N_6139,N_3825,N_4636);
nand U6140 (N_6140,N_3329,N_4637);
nor U6141 (N_6141,N_3442,N_3420);
or U6142 (N_6142,N_5752,N_4474);
xnor U6143 (N_6143,N_5757,N_3080);
nand U6144 (N_6144,N_5476,N_4040);
and U6145 (N_6145,N_3113,N_3614);
and U6146 (N_6146,N_5979,N_3816);
xnor U6147 (N_6147,N_5747,N_3946);
xor U6148 (N_6148,N_4844,N_3646);
nor U6149 (N_6149,N_3480,N_4139);
nor U6150 (N_6150,N_4550,N_3732);
nor U6151 (N_6151,N_4103,N_4934);
or U6152 (N_6152,N_5073,N_3132);
and U6153 (N_6153,N_4186,N_4714);
xor U6154 (N_6154,N_3709,N_5951);
or U6155 (N_6155,N_5253,N_3397);
and U6156 (N_6156,N_3025,N_5021);
or U6157 (N_6157,N_4778,N_5521);
or U6158 (N_6158,N_4083,N_3227);
and U6159 (N_6159,N_4729,N_5698);
nor U6160 (N_6160,N_4591,N_5623);
nor U6161 (N_6161,N_4846,N_3603);
nor U6162 (N_6162,N_5962,N_3030);
nand U6163 (N_6163,N_4331,N_5939);
nand U6164 (N_6164,N_5881,N_4685);
nor U6165 (N_6165,N_4376,N_3073);
or U6166 (N_6166,N_5587,N_5347);
and U6167 (N_6167,N_4415,N_5124);
and U6168 (N_6168,N_5026,N_5920);
or U6169 (N_6169,N_5816,N_3243);
nand U6170 (N_6170,N_5422,N_5639);
xnor U6171 (N_6171,N_4397,N_5873);
and U6172 (N_6172,N_4110,N_5281);
nor U6173 (N_6173,N_5471,N_4195);
or U6174 (N_6174,N_5604,N_3682);
nor U6175 (N_6175,N_4053,N_5683);
or U6176 (N_6176,N_4069,N_5646);
nand U6177 (N_6177,N_5245,N_3920);
or U6178 (N_6178,N_4175,N_5589);
nor U6179 (N_6179,N_4404,N_3040);
nand U6180 (N_6180,N_3668,N_5856);
and U6181 (N_6181,N_4789,N_5275);
nor U6182 (N_6182,N_5466,N_4922);
xnor U6183 (N_6183,N_3115,N_3679);
xor U6184 (N_6184,N_4241,N_3700);
and U6185 (N_6185,N_4263,N_4613);
or U6186 (N_6186,N_3445,N_4483);
nand U6187 (N_6187,N_4771,N_3170);
nor U6188 (N_6188,N_4085,N_3631);
nor U6189 (N_6189,N_5328,N_4138);
xnor U6190 (N_6190,N_5975,N_3546);
or U6191 (N_6191,N_4239,N_5908);
nand U6192 (N_6192,N_4567,N_4586);
or U6193 (N_6193,N_4403,N_3552);
or U6194 (N_6194,N_3347,N_5450);
or U6195 (N_6195,N_3559,N_5799);
nand U6196 (N_6196,N_3688,N_5591);
nor U6197 (N_6197,N_4750,N_3253);
and U6198 (N_6198,N_3037,N_5440);
and U6199 (N_6199,N_3091,N_3587);
or U6200 (N_6200,N_3068,N_3452);
nor U6201 (N_6201,N_5375,N_5602);
or U6202 (N_6202,N_3274,N_5389);
and U6203 (N_6203,N_5932,N_3354);
nand U6204 (N_6204,N_5355,N_4899);
or U6205 (N_6205,N_4160,N_4879);
nand U6206 (N_6206,N_5570,N_4845);
xor U6207 (N_6207,N_4512,N_3314);
and U6208 (N_6208,N_3813,N_5755);
or U6209 (N_6209,N_3110,N_5108);
xnor U6210 (N_6210,N_3186,N_4436);
or U6211 (N_6211,N_3918,N_3568);
nor U6212 (N_6212,N_3062,N_4670);
or U6213 (N_6213,N_3555,N_3950);
nor U6214 (N_6214,N_5758,N_5560);
and U6215 (N_6215,N_3794,N_5887);
xnor U6216 (N_6216,N_3584,N_5297);
xor U6217 (N_6217,N_3746,N_5541);
or U6218 (N_6218,N_3702,N_5301);
nand U6219 (N_6219,N_3871,N_3538);
nand U6220 (N_6220,N_3508,N_5786);
nand U6221 (N_6221,N_4639,N_4725);
or U6222 (N_6222,N_5661,N_4475);
or U6223 (N_6223,N_4166,N_3738);
and U6224 (N_6224,N_5449,N_4168);
nor U6225 (N_6225,N_3328,N_3909);
nor U6226 (N_6226,N_4495,N_5125);
nand U6227 (N_6227,N_5282,N_3967);
nand U6228 (N_6228,N_3716,N_3582);
and U6229 (N_6229,N_4025,N_4389);
or U6230 (N_6230,N_5734,N_4581);
xnor U6231 (N_6231,N_4060,N_5808);
or U6232 (N_6232,N_3847,N_4499);
or U6233 (N_6233,N_5842,N_5536);
and U6234 (N_6234,N_3151,N_3665);
or U6235 (N_6235,N_5884,N_5362);
or U6236 (N_6236,N_5031,N_5605);
nand U6237 (N_6237,N_3510,N_3152);
xor U6238 (N_6238,N_5346,N_3933);
and U6239 (N_6239,N_3388,N_3905);
xnor U6240 (N_6240,N_5014,N_4458);
and U6241 (N_6241,N_4602,N_3910);
and U6242 (N_6242,N_5292,N_4169);
nor U6243 (N_6243,N_4156,N_5807);
or U6244 (N_6244,N_3447,N_3359);
and U6245 (N_6245,N_5915,N_4858);
nor U6246 (N_6246,N_3987,N_5429);
nor U6247 (N_6247,N_3495,N_4076);
xor U6248 (N_6248,N_3053,N_3237);
nand U6249 (N_6249,N_5603,N_5242);
or U6250 (N_6250,N_4615,N_5561);
and U6251 (N_6251,N_3519,N_5861);
or U6252 (N_6252,N_5682,N_5000);
and U6253 (N_6253,N_4523,N_3008);
or U6254 (N_6254,N_4838,N_3294);
and U6255 (N_6255,N_4668,N_4692);
nand U6256 (N_6256,N_3288,N_4813);
xor U6257 (N_6257,N_5488,N_4940);
nor U6258 (N_6258,N_3766,N_4950);
or U6259 (N_6259,N_3057,N_4963);
nor U6260 (N_6260,N_4293,N_5634);
and U6261 (N_6261,N_4215,N_3764);
nor U6262 (N_6262,N_3513,N_3026);
xnor U6263 (N_6263,N_4881,N_3055);
nand U6264 (N_6264,N_4769,N_5965);
or U6265 (N_6265,N_5625,N_3457);
or U6266 (N_6266,N_5211,N_3362);
and U6267 (N_6267,N_5320,N_5569);
nand U6268 (N_6268,N_4607,N_3818);
or U6269 (N_6269,N_5329,N_5846);
and U6270 (N_6270,N_3319,N_3205);
nor U6271 (N_6271,N_4416,N_5037);
nor U6272 (N_6272,N_3986,N_4981);
nor U6273 (N_6273,N_4063,N_3140);
nor U6274 (N_6274,N_5759,N_4793);
nor U6275 (N_6275,N_3579,N_4278);
nand U6276 (N_6276,N_5159,N_4600);
nand U6277 (N_6277,N_3046,N_4114);
nand U6278 (N_6278,N_4362,N_4822);
or U6279 (N_6279,N_5956,N_5060);
nor U6280 (N_6280,N_4430,N_3064);
or U6281 (N_6281,N_4211,N_4459);
and U6282 (N_6282,N_3361,N_3585);
nor U6283 (N_6283,N_4905,N_3981);
or U6284 (N_6284,N_3074,N_5715);
or U6285 (N_6285,N_3250,N_3496);
and U6286 (N_6286,N_5268,N_5957);
xnor U6287 (N_6287,N_5023,N_5680);
and U6288 (N_6288,N_4540,N_3756);
and U6289 (N_6289,N_5812,N_4301);
nand U6290 (N_6290,N_4583,N_5312);
nand U6291 (N_6291,N_4991,N_5215);
nor U6292 (N_6292,N_5121,N_3696);
and U6293 (N_6293,N_4494,N_5325);
and U6294 (N_6294,N_4918,N_3042);
nand U6295 (N_6295,N_4504,N_4228);
nand U6296 (N_6296,N_5614,N_3324);
nand U6297 (N_6297,N_5183,N_5735);
or U6298 (N_6298,N_3681,N_5504);
nor U6299 (N_6299,N_5558,N_4820);
xnor U6300 (N_6300,N_3137,N_3075);
and U6301 (N_6301,N_5319,N_5016);
nor U6302 (N_6302,N_4425,N_4438);
nand U6303 (N_6303,N_4594,N_3565);
or U6304 (N_6304,N_5195,N_5232);
and U6305 (N_6305,N_4706,N_5845);
and U6306 (N_6306,N_4989,N_3462);
nor U6307 (N_6307,N_3972,N_3259);
or U6308 (N_6308,N_4212,N_3372);
or U6309 (N_6309,N_5955,N_4008);
and U6310 (N_6310,N_3256,N_3570);
nand U6311 (N_6311,N_3414,N_4791);
nand U6312 (N_6312,N_4926,N_3805);
and U6313 (N_6313,N_5677,N_5455);
and U6314 (N_6314,N_3964,N_5091);
nand U6315 (N_6315,N_4485,N_4170);
or U6316 (N_6316,N_3581,N_3544);
nand U6317 (N_6317,N_3504,N_5306);
or U6318 (N_6318,N_5323,N_3547);
or U6319 (N_6319,N_5228,N_3841);
or U6320 (N_6320,N_4121,N_4737);
nor U6321 (N_6321,N_4953,N_5404);
and U6322 (N_6322,N_4122,N_3628);
or U6323 (N_6323,N_5917,N_4055);
and U6324 (N_6324,N_3712,N_4068);
xnor U6325 (N_6325,N_4258,N_4551);
and U6326 (N_6326,N_4286,N_3315);
nand U6327 (N_6327,N_3873,N_5788);
nand U6328 (N_6328,N_3387,N_4782);
and U6329 (N_6329,N_3929,N_5659);
xnor U6330 (N_6330,N_4112,N_5233);
or U6331 (N_6331,N_4518,N_5529);
nand U6332 (N_6332,N_4145,N_3620);
and U6333 (N_6333,N_3799,N_3490);
or U6334 (N_6334,N_3820,N_5823);
xnor U6335 (N_6335,N_3890,N_3460);
nand U6336 (N_6336,N_5847,N_3369);
nand U6337 (N_6337,N_4111,N_4159);
nand U6338 (N_6338,N_4695,N_3583);
nor U6339 (N_6339,N_5720,N_5274);
xor U6340 (N_6340,N_4410,N_5789);
nor U6341 (N_6341,N_4826,N_4298);
and U6342 (N_6342,N_4198,N_3242);
or U6343 (N_6343,N_4976,N_3914);
nand U6344 (N_6344,N_5040,N_4208);
and U6345 (N_6345,N_4004,N_4683);
and U6346 (N_6346,N_3105,N_3863);
xnor U6347 (N_6347,N_4344,N_3394);
or U6348 (N_6348,N_3777,N_5302);
nand U6349 (N_6349,N_5822,N_3334);
nand U6350 (N_6350,N_5510,N_4931);
nor U6351 (N_6351,N_4509,N_3965);
nand U6352 (N_6352,N_3744,N_3059);
nor U6353 (N_6353,N_5022,N_3134);
or U6354 (N_6354,N_4229,N_4130);
nand U6355 (N_6355,N_5701,N_3683);
and U6356 (N_6356,N_4271,N_3183);
nor U6357 (N_6357,N_4947,N_5227);
nand U6358 (N_6358,N_4300,N_3507);
xnor U6359 (N_6359,N_4927,N_4369);
or U6360 (N_6360,N_4759,N_3228);
nand U6361 (N_6361,N_4697,N_3203);
or U6362 (N_6362,N_4154,N_3882);
xnor U6363 (N_6363,N_4391,N_4314);
xor U6364 (N_6364,N_4988,N_4192);
and U6365 (N_6365,N_3071,N_4887);
xnor U6366 (N_6366,N_5574,N_3821);
nor U6367 (N_6367,N_4761,N_5041);
or U6368 (N_6368,N_5202,N_3705);
nor U6369 (N_6369,N_4658,N_4890);
xor U6370 (N_6370,N_5821,N_4892);
or U6371 (N_6371,N_4783,N_4405);
nand U6372 (N_6372,N_3669,N_5826);
nor U6373 (N_6373,N_5985,N_4066);
xnor U6374 (N_6374,N_4776,N_3456);
nand U6375 (N_6375,N_5984,N_4672);
xor U6376 (N_6376,N_4411,N_4912);
nor U6377 (N_6377,N_5030,N_3648);
nor U6378 (N_6378,N_4447,N_4560);
or U6379 (N_6379,N_4452,N_3590);
nor U6380 (N_6380,N_3100,N_4061);
nand U6381 (N_6381,N_4099,N_5563);
nor U6382 (N_6382,N_3917,N_3304);
nor U6383 (N_6383,N_5394,N_5870);
and U6384 (N_6384,N_3234,N_3831);
or U6385 (N_6385,N_4595,N_5185);
nor U6386 (N_6386,N_3021,N_5384);
or U6387 (N_6387,N_5425,N_4830);
or U6388 (N_6388,N_3903,N_3806);
and U6389 (N_6389,N_4364,N_4460);
nand U6390 (N_6390,N_3306,N_4146);
nand U6391 (N_6391,N_4664,N_5969);
nor U6392 (N_6392,N_3823,N_5891);
nand U6393 (N_6393,N_3488,N_5730);
and U6394 (N_6394,N_5096,N_5224);
nand U6395 (N_6395,N_4648,N_4665);
and U6396 (N_6396,N_5961,N_4187);
and U6397 (N_6397,N_5130,N_4559);
or U6398 (N_6398,N_4641,N_3339);
or U6399 (N_6399,N_3613,N_5753);
or U6400 (N_6400,N_3138,N_4189);
and U6401 (N_6401,N_5298,N_4954);
and U6402 (N_6402,N_4557,N_5927);
and U6403 (N_6403,N_3567,N_5689);
nor U6404 (N_6404,N_4479,N_5695);
nor U6405 (N_6405,N_5717,N_4466);
and U6406 (N_6406,N_3978,N_5796);
xor U6407 (N_6407,N_3997,N_5746);
and U6408 (N_6408,N_5348,N_4958);
nor U6409 (N_6409,N_5248,N_4006);
nor U6410 (N_6410,N_4002,N_4463);
and U6411 (N_6411,N_5514,N_4917);
nand U6412 (N_6412,N_4484,N_4279);
nor U6413 (N_6413,N_4593,N_4107);
nor U6414 (N_6414,N_3086,N_3482);
xor U6415 (N_6415,N_4440,N_3699);
xor U6416 (N_6416,N_3425,N_5489);
and U6417 (N_6417,N_5244,N_4281);
nand U6418 (N_6418,N_4084,N_5586);
nand U6419 (N_6419,N_5164,N_4357);
or U6420 (N_6420,N_5152,N_3220);
or U6421 (N_6421,N_4895,N_5357);
or U6422 (N_6422,N_5377,N_5685);
nor U6423 (N_6423,N_5356,N_4347);
or U6424 (N_6424,N_3290,N_4445);
nor U6425 (N_6425,N_5054,N_5163);
and U6426 (N_6426,N_4589,N_3718);
and U6427 (N_6427,N_4719,N_4677);
xor U6428 (N_6428,N_3177,N_4428);
nand U6429 (N_6429,N_3139,N_4903);
nor U6430 (N_6430,N_5792,N_4294);
and U6431 (N_6431,N_3532,N_4657);
and U6432 (N_6432,N_3382,N_5700);
and U6433 (N_6433,N_3448,N_4880);
nor U6434 (N_6434,N_5548,N_4603);
nand U6435 (N_6435,N_4318,N_3674);
and U6436 (N_6436,N_4840,N_4694);
nand U6437 (N_6437,N_5378,N_4078);
and U6438 (N_6438,N_3380,N_5327);
nor U6439 (N_6439,N_4444,N_4222);
xor U6440 (N_6440,N_3755,N_4091);
or U6441 (N_6441,N_5006,N_3418);
xnor U6442 (N_6442,N_5933,N_5388);
nor U6443 (N_6443,N_4851,N_3384);
and U6444 (N_6444,N_5116,N_4072);
and U6445 (N_6445,N_5019,N_5068);
or U6446 (N_6446,N_3723,N_4983);
nand U6447 (N_6447,N_4167,N_4616);
nor U6448 (N_6448,N_3287,N_4036);
or U6449 (N_6449,N_3449,N_5609);
nor U6450 (N_6450,N_4381,N_4773);
nand U6451 (N_6451,N_4515,N_5173);
nand U6452 (N_6452,N_5597,N_5142);
and U6453 (N_6453,N_4896,N_3506);
xnor U6454 (N_6454,N_4237,N_5247);
nor U6455 (N_6455,N_4042,N_3940);
or U6456 (N_6456,N_3888,N_5112);
or U6457 (N_6457,N_5213,N_3497);
nand U6458 (N_6458,N_3983,N_3770);
nor U6459 (N_6459,N_4467,N_3522);
or U6460 (N_6460,N_3992,N_5057);
or U6461 (N_6461,N_3686,N_4815);
and U6462 (N_6462,N_5279,N_3849);
nor U6463 (N_6463,N_5813,N_5836);
xor U6464 (N_6464,N_3654,N_5007);
or U6465 (N_6465,N_3084,N_3531);
or U6466 (N_6466,N_5139,N_3647);
nor U6467 (N_6467,N_4221,N_5518);
or U6468 (N_6468,N_5210,N_3352);
nor U6469 (N_6469,N_4207,N_3902);
or U6470 (N_6470,N_4774,N_3801);
nand U6471 (N_6471,N_5869,N_5435);
nand U6472 (N_6472,N_3518,N_4179);
or U6473 (N_6473,N_3989,N_3353);
and U6474 (N_6474,N_3615,N_3426);
xnor U6475 (N_6475,N_3106,N_4486);
nand U6476 (N_6476,N_5825,N_5771);
and U6477 (N_6477,N_3515,N_5966);
nor U6478 (N_6478,N_4623,N_5524);
nor U6479 (N_6479,N_5766,N_3416);
and U6480 (N_6480,N_4629,N_5187);
nor U6481 (N_6481,N_5371,N_5793);
and U6482 (N_6482,N_4872,N_3365);
or U6483 (N_6483,N_4847,N_4441);
nor U6484 (N_6484,N_4334,N_5652);
and U6485 (N_6485,N_3350,N_4755);
nand U6486 (N_6486,N_4539,N_4032);
nand U6487 (N_6487,N_5086,N_3408);
and U6488 (N_6488,N_4088,N_3586);
or U6489 (N_6489,N_5800,N_5740);
nor U6490 (N_6490,N_3872,N_5495);
or U6491 (N_6491,N_3087,N_4724);
nor U6492 (N_6492,N_4684,N_3778);
nand U6493 (N_6493,N_4307,N_5517);
or U6494 (N_6494,N_5676,N_5145);
and U6495 (N_6495,N_5970,N_5650);
nor U6496 (N_6496,N_5053,N_3127);
or U6497 (N_6497,N_4998,N_4224);
nand U6498 (N_6498,N_5397,N_3431);
nor U6499 (N_6499,N_3897,N_4137);
and U6500 (N_6500,N_5351,N_4407);
xnor U6501 (N_6501,N_4104,N_4193);
nor U6502 (N_6502,N_5905,N_5167);
or U6503 (N_6503,N_3649,N_4775);
nand U6504 (N_6504,N_3485,N_5479);
or U6505 (N_6505,N_5539,N_5993);
nor U6506 (N_6506,N_4124,N_5911);
nor U6507 (N_6507,N_4049,N_3795);
xor U6508 (N_6508,N_5947,N_5523);
or U6509 (N_6509,N_4262,N_5778);
or U6510 (N_6510,N_3944,N_5256);
nor U6511 (N_6511,N_3934,N_3370);
nor U6512 (N_6512,N_3404,N_3331);
nand U6513 (N_6513,N_4544,N_4070);
and U6514 (N_6514,N_5543,N_5153);
or U6515 (N_6515,N_3302,N_4507);
and U6516 (N_6516,N_3733,N_3092);
nand U6517 (N_6517,N_4891,N_4039);
nor U6518 (N_6518,N_5745,N_3019);
nor U6519 (N_6519,N_4333,N_5408);
nand U6520 (N_6520,N_3533,N_4327);
nor U6521 (N_6521,N_5333,N_4865);
nor U6522 (N_6522,N_4946,N_4627);
nor U6523 (N_6523,N_4948,N_5967);
and U6524 (N_6524,N_3793,N_5585);
and U6525 (N_6525,N_4556,N_3121);
nand U6526 (N_6526,N_3135,N_4951);
and U6527 (N_6527,N_5423,N_3099);
or U6528 (N_6528,N_5624,N_3687);
or U6529 (N_6529,N_3411,N_5428);
nor U6530 (N_6530,N_4355,N_5340);
and U6531 (N_6531,N_3659,N_3768);
nor U6532 (N_6532,N_5937,N_3734);
nor U6533 (N_6533,N_5396,N_4752);
or U6534 (N_6534,N_4478,N_4564);
nand U6535 (N_6535,N_5446,N_5810);
or U6536 (N_6536,N_5830,N_5568);
xnor U6537 (N_6537,N_5322,N_4973);
nor U6538 (N_6538,N_5629,N_3802);
nor U6539 (N_6539,N_3787,N_5672);
nand U6540 (N_6540,N_3049,N_5102);
nor U6541 (N_6541,N_5573,N_3599);
xnor U6542 (N_6542,N_3672,N_3842);
xor U6543 (N_6543,N_4654,N_3713);
nor U6544 (N_6544,N_5854,N_3854);
or U6545 (N_6545,N_3627,N_4713);
nand U6546 (N_6546,N_5611,N_5252);
or U6547 (N_6547,N_3742,N_3542);
nor U6548 (N_6548,N_5742,N_4141);
nand U6549 (N_6549,N_4580,N_4243);
and U6550 (N_6550,N_5223,N_4213);
nand U6551 (N_6551,N_3167,N_3172);
nor U6552 (N_6552,N_5255,N_4412);
or U6553 (N_6553,N_4194,N_5904);
nand U6554 (N_6554,N_5157,N_5772);
nor U6555 (N_6555,N_3195,N_4832);
and U6556 (N_6556,N_3824,N_5697);
nor U6557 (N_6557,N_3162,N_4450);
and U6558 (N_6558,N_3430,N_5462);
or U6559 (N_6559,N_5642,N_3465);
or U6560 (N_6560,N_4854,N_5660);
xnor U6561 (N_6561,N_3325,N_4026);
and U6562 (N_6562,N_3727,N_3520);
and U6563 (N_6563,N_4659,N_3564);
and U6564 (N_6564,N_3428,N_3159);
or U6565 (N_6565,N_5549,N_3891);
and U6566 (N_6566,N_4311,N_4628);
and U6567 (N_6567,N_4267,N_5286);
xnor U6568 (N_6568,N_3796,N_3261);
or U6569 (N_6569,N_5712,N_5820);
nand U6570 (N_6570,N_5653,N_5829);
and U6571 (N_6571,N_4470,N_3703);
nor U6572 (N_6572,N_5718,N_4715);
and U6573 (N_6573,N_3407,N_3150);
and U6574 (N_6574,N_5101,N_3469);
nor U6575 (N_6575,N_3859,N_5170);
nand U6576 (N_6576,N_4739,N_5284);
xor U6577 (N_6577,N_3212,N_4599);
and U6578 (N_6578,N_4968,N_3893);
nand U6579 (N_6579,N_3481,N_3255);
and U6580 (N_6580,N_3245,N_5209);
xor U6581 (N_6581,N_4214,N_4608);
or U6582 (N_6582,N_4784,N_5707);
or U6583 (N_6583,N_5851,N_4218);
nand U6584 (N_6584,N_4604,N_4868);
and U6585 (N_6585,N_5582,N_5017);
and U6586 (N_6586,N_5696,N_4516);
and U6587 (N_6587,N_3278,N_5907);
nand U6588 (N_6588,N_3503,N_5482);
and U6589 (N_6589,N_4909,N_5872);
nand U6590 (N_6590,N_3077,N_5841);
nor U6591 (N_6591,N_5212,N_5678);
nor U6592 (N_6592,N_4626,N_4320);
nor U6593 (N_6593,N_4077,N_5693);
nand U6594 (N_6594,N_3721,N_3345);
nand U6595 (N_6595,N_3398,N_3307);
nand U6596 (N_6596,N_3541,N_4624);
xnor U6597 (N_6597,N_3487,N_3422);
and U6598 (N_6598,N_5277,N_5246);
and U6599 (N_6599,N_3179,N_5118);
xnor U6600 (N_6600,N_3123,N_5754);
and U6601 (N_6601,N_4244,N_4709);
nor U6602 (N_6602,N_3808,N_4688);
and U6603 (N_6603,N_5567,N_3671);
nor U6604 (N_6604,N_4161,N_4573);
nor U6605 (N_6605,N_3358,N_5487);
and U6606 (N_6606,N_3701,N_3185);
nor U6607 (N_6607,N_5580,N_3736);
xnor U6608 (N_6608,N_4582,N_3757);
nor U6609 (N_6609,N_3168,N_4699);
or U6610 (N_6610,N_5149,N_5166);
nor U6611 (N_6611,N_3088,N_5618);
nand U6612 (N_6612,N_4990,N_3090);
and U6613 (N_6613,N_5995,N_5241);
nor U6614 (N_6614,N_4517,N_3509);
nor U6615 (N_6615,N_4422,N_5361);
and U6616 (N_6616,N_3036,N_4502);
and U6617 (N_6617,N_4044,N_4995);
and U6618 (N_6618,N_5443,N_3340);
nor U6619 (N_6619,N_4013,N_5990);
nor U6620 (N_6620,N_4984,N_5819);
and U6621 (N_6621,N_4992,N_4093);
nor U6622 (N_6622,N_4794,N_3349);
or U6623 (N_6623,N_3685,N_5801);
xnor U6624 (N_6624,N_3093,N_4574);
or U6625 (N_6625,N_4238,N_3775);
and U6626 (N_6626,N_5928,N_5010);
or U6627 (N_6627,N_4358,N_5769);
xnor U6628 (N_6628,N_3158,N_5919);
or U6629 (N_6629,N_4094,N_4704);
or U6630 (N_6630,N_4453,N_5914);
or U6631 (N_6631,N_3767,N_5506);
nand U6632 (N_6632,N_4819,N_4030);
and U6633 (N_6633,N_5986,N_3204);
or U6634 (N_6634,N_5835,N_4727);
nand U6635 (N_6635,N_5075,N_3968);
and U6636 (N_6636,N_3540,N_5494);
nor U6637 (N_6637,N_3749,N_4503);
nand U6638 (N_6638,N_3834,N_3327);
or U6639 (N_6639,N_5922,N_3076);
and U6640 (N_6640,N_3803,N_4651);
and U6641 (N_6641,N_4915,N_4113);
and U6642 (N_6642,N_3056,N_4570);
or U6643 (N_6643,N_3124,N_4308);
and U6644 (N_6644,N_4038,N_5739);
and U6645 (N_6645,N_3194,N_5729);
nand U6646 (N_6646,N_5875,N_4787);
nor U6647 (N_6647,N_5411,N_3171);
nand U6648 (N_6648,N_5764,N_4678);
xor U6649 (N_6649,N_5184,N_3804);
xor U6650 (N_6650,N_3643,N_5996);
nor U6651 (N_6651,N_5432,N_3958);
nor U6652 (N_6652,N_4861,N_3862);
nor U6653 (N_6653,N_5868,N_3389);
and U6654 (N_6654,N_4356,N_5237);
and U6655 (N_6655,N_4568,N_4395);
or U6656 (N_6656,N_5686,N_5547);
xnor U6657 (N_6657,N_5342,N_4382);
nor U6658 (N_6658,N_3248,N_4372);
and U6659 (N_6659,N_4321,N_3272);
nor U6660 (N_6660,N_3018,N_4744);
or U6661 (N_6661,N_4640,N_5613);
or U6662 (N_6662,N_3231,N_3377);
nand U6663 (N_6663,N_5161,N_5165);
or U6664 (N_6664,N_4131,N_5105);
nand U6665 (N_6665,N_5557,N_3514);
or U6666 (N_6666,N_5434,N_5670);
and U6667 (N_6667,N_4468,N_5205);
and U6668 (N_6668,N_5704,N_3578);
and U6669 (N_6669,N_3262,N_3116);
and U6670 (N_6670,N_3562,N_4796);
nor U6671 (N_6671,N_3927,N_4181);
nor U6672 (N_6672,N_3045,N_5756);
or U6673 (N_6673,N_4906,N_5012);
or U6674 (N_6674,N_5427,N_3374);
nor U6675 (N_6675,N_3560,N_3720);
and U6676 (N_6676,N_3850,N_5430);
nand U6677 (N_6677,N_3260,N_4396);
xnor U6678 (N_6678,N_3039,N_4439);
nor U6679 (N_6679,N_4610,N_4563);
and U6680 (N_6680,N_5828,N_4158);
or U6681 (N_6681,N_4126,N_4522);
or U6682 (N_6682,N_4885,N_4999);
nor U6683 (N_6683,N_4202,N_4806);
and U6684 (N_6684,N_3273,N_4096);
and U6685 (N_6685,N_4662,N_4916);
or U6686 (N_6686,N_5500,N_5169);
and U6687 (N_6687,N_4883,N_4562);
nor U6688 (N_6688,N_4448,N_5412);
nor U6689 (N_6689,N_3383,N_5722);
or U6690 (N_6690,N_3941,N_4201);
nand U6691 (N_6691,N_4821,N_3453);
or U6692 (N_6692,N_5706,N_4997);
xnor U6693 (N_6693,N_3437,N_3835);
and U6694 (N_6694,N_5178,N_3690);
or U6695 (N_6695,N_4386,N_5467);
and U6696 (N_6696,N_3246,N_3410);
nor U6697 (N_6697,N_4031,N_5505);
nor U6698 (N_6698,N_3810,N_3489);
nor U6699 (N_6699,N_3085,N_3101);
xor U6700 (N_6700,N_3155,N_4873);
nand U6701 (N_6701,N_5780,N_3050);
nand U6702 (N_6702,N_4760,N_3161);
or U6703 (N_6703,N_3015,N_3376);
nor U6704 (N_6704,N_4010,N_4661);
and U6705 (N_6705,N_5649,N_4919);
and U6706 (N_6706,N_5809,N_4247);
nand U6707 (N_6707,N_3715,N_4575);
nor U6708 (N_6708,N_5501,N_3379);
nor U6709 (N_6709,N_5991,N_4074);
nor U6710 (N_6710,N_3523,N_5824);
nor U6711 (N_6711,N_3954,N_4437);
and U6712 (N_6712,N_5657,N_4972);
nand U6713 (N_6713,N_5508,N_4514);
and U6714 (N_6714,N_3364,N_5368);
and U6715 (N_6715,N_3792,N_3607);
or U6716 (N_6716,N_4340,N_3996);
and U6717 (N_6717,N_3960,N_5390);
and U6718 (N_6718,N_4366,N_5552);
xnor U6719 (N_6719,N_5832,N_5240);
and U6720 (N_6720,N_4843,N_5383);
or U6721 (N_6721,N_3832,N_3629);
nor U6722 (N_6722,N_4967,N_4469);
or U6723 (N_6723,N_4142,N_5865);
xnor U6724 (N_6724,N_5332,N_4432);
and U6725 (N_6725,N_5477,N_5513);
nand U6726 (N_6726,N_3754,N_5036);
or U6727 (N_6727,N_3866,N_4067);
nor U6728 (N_6728,N_5674,N_4962);
nand U6729 (N_6729,N_4317,N_5894);
nand U6730 (N_6730,N_3413,N_3187);
or U6731 (N_6731,N_3870,N_4206);
or U6732 (N_6732,N_3693,N_5930);
nor U6733 (N_6733,N_4676,N_4303);
xnor U6734 (N_6734,N_5175,N_5637);
nor U6735 (N_6735,N_3468,N_4313);
or U6736 (N_6736,N_5551,N_5999);
xnor U6737 (N_6737,N_4233,N_5787);
nand U6738 (N_6738,N_4217,N_4797);
nor U6739 (N_6739,N_4508,N_4743);
nand U6740 (N_6740,N_5344,N_3010);
and U6741 (N_6741,N_5584,N_4209);
or U6742 (N_6742,N_4136,N_5593);
nand U6743 (N_6743,N_5519,N_4552);
nor U6744 (N_6744,N_3371,N_4703);
xor U6745 (N_6745,N_5608,N_4341);
xnor U6746 (N_6746,N_3209,N_5448);
nand U6747 (N_6747,N_4392,N_4959);
nor U6748 (N_6748,N_4878,N_3676);
nand U6749 (N_6749,N_3330,N_3632);
nor U6750 (N_6750,N_3500,N_3066);
and U6751 (N_6751,N_3281,N_3856);
xor U6752 (N_6752,N_4371,N_5617);
and U6753 (N_6753,N_4853,N_3771);
nand U6754 (N_6754,N_3360,N_5520);
and U6755 (N_6755,N_4242,N_4497);
and U6756 (N_6756,N_3550,N_5943);
xnor U6757 (N_6757,N_4226,N_3692);
xnor U6758 (N_6758,N_5469,N_5339);
and U6759 (N_6759,N_3636,N_3561);
nand U6760 (N_6760,N_4803,N_3530);
and U6761 (N_6761,N_4975,N_3675);
or U6762 (N_6762,N_5321,N_5619);
nor U6763 (N_6763,N_4925,N_3639);
and U6764 (N_6764,N_5024,N_4108);
and U6765 (N_6765,N_5049,N_5749);
nor U6766 (N_6766,N_3285,N_3980);
and U6767 (N_6767,N_4152,N_5243);
or U6768 (N_6768,N_5208,N_5765);
or U6769 (N_6769,N_4277,N_3645);
or U6770 (N_6770,N_5784,N_5538);
nor U6771 (N_6771,N_4292,N_3141);
nand U6772 (N_6772,N_3526,N_5464);
nand U6773 (N_6773,N_5457,N_3006);
or U6774 (N_6774,N_3348,N_5018);
nor U6775 (N_6775,N_5590,N_3545);
xor U6776 (N_6776,N_3677,N_3007);
and U6777 (N_6777,N_4276,N_4109);
nand U6778 (N_6778,N_3711,N_4064);
nand U6779 (N_6779,N_5525,N_5853);
or U6780 (N_6780,N_4848,N_4807);
or U6781 (N_6781,N_3889,N_4095);
nor U6782 (N_6782,N_3342,N_4147);
nor U6783 (N_6783,N_5311,N_4464);
or U6784 (N_6784,N_5797,N_4140);
nand U6785 (N_6785,N_4200,N_5768);
nor U6786 (N_6786,N_3118,N_3517);
or U6787 (N_6787,N_4482,N_5189);
or U6788 (N_6788,N_3446,N_5330);
nand U6789 (N_6789,N_5944,N_4601);
nand U6790 (N_6790,N_4937,N_4527);
or U6791 (N_6791,N_5135,N_5804);
or U6792 (N_6792,N_4429,N_4764);
and U6793 (N_6793,N_4741,N_3658);
and U6794 (N_6794,N_3142,N_4035);
nor U6795 (N_6795,N_5144,N_4304);
nor U6796 (N_6796,N_5419,N_3995);
nand U6797 (N_6797,N_4577,N_5850);
nand U6798 (N_6798,N_4117,N_3881);
nand U6799 (N_6799,N_5094,N_3023);
or U6800 (N_6800,N_5805,N_5631);
nand U6801 (N_6801,N_4256,N_3623);
and U6802 (N_6802,N_5705,N_3218);
and U6803 (N_6803,N_3655,N_5627);
and U6804 (N_6804,N_5968,N_3652);
nand U6805 (N_6805,N_5099,N_4462);
or U6806 (N_6806,N_4492,N_4859);
nand U6807 (N_6807,N_4332,N_4073);
or U6808 (N_6808,N_4510,N_4377);
xnor U6809 (N_6809,N_5950,N_4705);
xnor U6810 (N_6810,N_3396,N_4680);
xor U6811 (N_6811,N_5267,N_4969);
nand U6812 (N_6812,N_4014,N_4770);
nand U6813 (N_6813,N_3033,N_5131);
nand U6814 (N_6814,N_3082,N_4911);
and U6815 (N_6815,N_3421,N_3763);
nor U6816 (N_6816,N_5402,N_3385);
or U6817 (N_6817,N_3321,N_4894);
or U6818 (N_6818,N_3268,N_4120);
nor U6819 (N_6819,N_3060,N_4171);
or U6820 (N_6820,N_5817,N_4747);
nand U6821 (N_6821,N_5622,N_4289);
nor U6822 (N_6822,N_5645,N_5200);
and U6823 (N_6823,N_4809,N_4087);
and U6824 (N_6824,N_5082,N_5386);
nor U6825 (N_6825,N_5313,N_5737);
nand U6826 (N_6826,N_4196,N_4280);
and U6827 (N_6827,N_5201,N_5994);
or U6828 (N_6828,N_3745,N_4406);
or U6829 (N_6829,N_3301,N_4884);
or U6830 (N_6830,N_5080,N_3125);
nor U6831 (N_6831,N_3476,N_5069);
nand U6832 (N_6832,N_4735,N_4451);
nand U6833 (N_6833,N_3622,N_3373);
xnor U6834 (N_6834,N_5147,N_5785);
or U6835 (N_6835,N_3455,N_4833);
nor U6836 (N_6836,N_4234,N_5509);
nand U6837 (N_6837,N_3098,N_3740);
and U6838 (N_6838,N_3998,N_4190);
or U6839 (N_6839,N_3577,N_4409);
or U6840 (N_6840,N_4758,N_5566);
nor U6841 (N_6841,N_5410,N_5725);
nor U6842 (N_6842,N_3604,N_5763);
nor U6843 (N_6843,N_3174,N_4795);
or U6844 (N_6844,N_5644,N_4928);
nand U6845 (N_6845,N_4295,N_5134);
xnor U6846 (N_6846,N_3774,N_3224);
or U6847 (N_6847,N_5129,N_3119);
nand U6848 (N_6848,N_3529,N_4421);
nand U6849 (N_6849,N_5902,N_5070);
or U6850 (N_6850,N_3254,N_4380);
and U6851 (N_6851,N_3600,N_5071);
xnor U6852 (N_6852,N_4052,N_5774);
nor U6853 (N_6853,N_5369,N_3880);
nand U6854 (N_6854,N_4996,N_5106);
and U6855 (N_6855,N_5790,N_3233);
nand U6856 (N_6856,N_4119,N_4964);
nand U6857 (N_6857,N_3912,N_4632);
xor U6858 (N_6858,N_5221,N_5295);
nand U6859 (N_6859,N_4143,N_3892);
nor U6860 (N_6860,N_3283,N_4576);
or U6861 (N_6861,N_4565,N_3471);
nand U6862 (N_6862,N_4663,N_3198);
and U6863 (N_6863,N_4635,N_4172);
nand U6864 (N_6864,N_4323,N_5382);
nand U6865 (N_6865,N_4153,N_3576);
nand U6866 (N_6866,N_4722,N_4656);
or U6867 (N_6867,N_3096,N_3375);
xnor U6868 (N_6868,N_5728,N_5974);
nand U6869 (N_6869,N_4270,N_5420);
or U6870 (N_6870,N_5640,N_5782);
and U6871 (N_6871,N_3678,N_4157);
nor U6872 (N_6872,N_3058,N_3226);
or U6873 (N_6873,N_5458,N_5002);
and U6874 (N_6874,N_4148,N_4660);
nor U6875 (N_6875,N_4901,N_4634);
and U6876 (N_6876,N_5269,N_4691);
and U6877 (N_6877,N_4536,N_5289);
or U6878 (N_6878,N_5093,N_4102);
and U6879 (N_6879,N_3160,N_3899);
nor U6880 (N_6880,N_5981,N_4427);
nor U6881 (N_6881,N_4693,N_4261);
or U6882 (N_6882,N_3548,N_4756);
and U6883 (N_6883,N_4379,N_5401);
xor U6884 (N_6884,N_5888,N_5795);
or U6885 (N_6885,N_5050,N_5194);
xnor U6886 (N_6886,N_5376,N_3332);
nand U6887 (N_6887,N_4057,N_3265);
nor U6888 (N_6888,N_4051,N_5179);
nor U6889 (N_6889,N_4642,N_3943);
and U6890 (N_6890,N_3239,N_3662);
and U6891 (N_6891,N_4302,N_5076);
nand U6892 (N_6892,N_3657,N_5516);
or U6893 (N_6893,N_5579,N_3153);
nor U6894 (N_6894,N_4757,N_4505);
xnor U6895 (N_6895,N_5098,N_4015);
and U6896 (N_6896,N_4231,N_5155);
nand U6897 (N_6897,N_3969,N_3016);
and U6898 (N_6898,N_5387,N_5499);
and U6899 (N_6899,N_5341,N_3963);
nor U6900 (N_6900,N_4941,N_5160);
nor U6901 (N_6901,N_5438,N_5537);
xnor U6902 (N_6902,N_4003,N_5334);
nor U6903 (N_6903,N_3391,N_3707);
or U6904 (N_6904,N_5815,N_5544);
or U6905 (N_6905,N_4034,N_3781);
nor U6906 (N_6906,N_5391,N_4987);
nand U6907 (N_6907,N_4720,N_4811);
or U6908 (N_6908,N_3926,N_3399);
nand U6909 (N_6909,N_5777,N_3975);
nor U6910 (N_6910,N_4408,N_3710);
nor U6911 (N_6911,N_4742,N_3154);
nor U6912 (N_6912,N_4808,N_4767);
nand U6913 (N_6913,N_3762,N_3819);
nor U6914 (N_6914,N_3641,N_5168);
xnor U6915 (N_6915,N_3556,N_3539);
or U6916 (N_6916,N_5744,N_5303);
xor U6917 (N_6917,N_3201,N_5308);
and U6918 (N_6918,N_3664,N_4900);
nor U6919 (N_6919,N_5307,N_4611);
nor U6920 (N_6920,N_4413,N_4191);
and U6921 (N_6921,N_4571,N_5453);
or U6922 (N_6922,N_3251,N_4090);
or U6923 (N_6923,N_3830,N_4765);
nor U6924 (N_6924,N_4115,N_3635);
nand U6925 (N_6925,N_5314,N_4465);
or U6926 (N_6926,N_5716,N_4324);
or U6927 (N_6927,N_3689,N_5150);
or U6928 (N_6928,N_5703,N_3276);
nor U6929 (N_6929,N_4871,N_3131);
nor U6930 (N_6930,N_3013,N_3136);
nor U6931 (N_6931,N_4367,N_3264);
nand U6932 (N_6932,N_5607,N_3400);
nor U6933 (N_6933,N_3439,N_5171);
nor U6934 (N_6934,N_3601,N_3719);
nand U6935 (N_6935,N_5418,N_3309);
nor U6936 (N_6936,N_5554,N_4135);
or U6937 (N_6937,N_3277,N_5399);
nor U6938 (N_6938,N_5691,N_5910);
or U6939 (N_6939,N_3516,N_4907);
and U6940 (N_6940,N_3479,N_3640);
nand U6941 (N_6941,N_5781,N_4252);
and U6942 (N_6942,N_3244,N_3436);
nor U6943 (N_6943,N_3551,N_4164);
nand U6944 (N_6944,N_4058,N_4548);
and U6945 (N_6945,N_4491,N_5498);
xnor U6946 (N_6946,N_5025,N_5522);
nor U6947 (N_6947,N_3157,N_4230);
nor U6948 (N_6948,N_3660,N_3176);
and U6949 (N_6949,N_3466,N_4249);
xor U6950 (N_6950,N_4511,N_4734);
and U6951 (N_6951,N_4127,N_3145);
and U6952 (N_6952,N_5638,N_3973);
or U6953 (N_6953,N_4961,N_4299);
nor U6954 (N_6954,N_3874,N_3217);
nand U6955 (N_6955,N_5405,N_5392);
and U6956 (N_6956,N_4075,N_4021);
and U6957 (N_6957,N_3694,N_5679);
nand U6958 (N_6958,N_4205,N_5192);
or U6959 (N_6959,N_5964,N_4618);
nor U6960 (N_6960,N_4645,N_5982);
nand U6961 (N_6961,N_4944,N_4180);
and U6962 (N_6962,N_3725,N_3708);
and U6963 (N_6963,N_5840,N_4296);
and U6964 (N_6964,N_3402,N_5056);
nor U6965 (N_6965,N_3368,N_3296);
nand U6966 (N_6966,N_4974,N_3403);
nor U6967 (N_6967,N_5437,N_3563);
or U6968 (N_6968,N_3760,N_3753);
or U6969 (N_6969,N_5931,N_3798);
xnor U6970 (N_6970,N_4541,N_5111);
nand U6971 (N_6971,N_4801,N_4011);
and U6972 (N_6972,N_4418,N_3790);
xor U6973 (N_6973,N_5107,N_4268);
nand U6974 (N_6974,N_3432,N_3011);
nor U6975 (N_6975,N_3267,N_4970);
nor U6976 (N_6976,N_3310,N_4751);
or U6977 (N_6977,N_5681,N_3811);
nand U6978 (N_6978,N_3303,N_4644);
xnor U6979 (N_6979,N_5844,N_4921);
nor U6980 (N_6980,N_4532,N_4804);
or U6981 (N_6981,N_5470,N_5379);
and U6982 (N_6982,N_5122,N_4537);
and U6983 (N_6983,N_3502,N_3670);
or U6984 (N_6984,N_4118,N_4251);
and U6985 (N_6985,N_3543,N_5655);
or U6986 (N_6986,N_4876,N_3779);
nand U6987 (N_6987,N_5748,N_3698);
and U6988 (N_6988,N_5087,N_5960);
and U6989 (N_6989,N_5310,N_3906);
nor U6990 (N_6990,N_3190,N_3602);
nand U6991 (N_6991,N_3438,N_3827);
xor U6992 (N_6992,N_4597,N_4520);
xnor U6993 (N_6993,N_5385,N_3003);
nor U6994 (N_6994,N_3955,N_4723);
nor U6995 (N_6995,N_3959,N_3419);
nor U6996 (N_6996,N_4449,N_5062);
and U6997 (N_6997,N_4993,N_3182);
or U6998 (N_6998,N_3916,N_3067);
or U6999 (N_6999,N_5436,N_4777);
or U7000 (N_7000,N_5288,N_5783);
nand U7001 (N_7001,N_3213,N_4621);
nand U7002 (N_7002,N_4817,N_3922);
nand U7003 (N_7003,N_3851,N_4609);
or U7004 (N_7004,N_5374,N_4490);
nand U7005 (N_7005,N_3908,N_4842);
xor U7006 (N_7006,N_4284,N_4017);
nor U7007 (N_7007,N_5481,N_5750);
and U7008 (N_7008,N_3363,N_3838);
nor U7009 (N_7009,N_3737,N_3343);
and U7010 (N_7010,N_3415,N_3836);
nor U7011 (N_7011,N_3165,N_5064);
nand U7012 (N_7012,N_3188,N_4667);
nor U7013 (N_7013,N_5454,N_3409);
nor U7014 (N_7014,N_3948,N_5663);
or U7015 (N_7015,N_5413,N_4862);
nor U7016 (N_7016,N_4227,N_3173);
nand U7017 (N_7017,N_3126,N_5896);
nor U7018 (N_7018,N_5945,N_5897);
or U7019 (N_7019,N_4414,N_5615);
and U7020 (N_7020,N_3491,N_4359);
or U7021 (N_7021,N_3605,N_4898);
nor U7022 (N_7022,N_3405,N_3472);
nor U7023 (N_7023,N_4841,N_4434);
nor U7024 (N_7024,N_4431,N_5424);
nand U7025 (N_7025,N_4368,N_5114);
nor U7026 (N_7026,N_3351,N_4902);
nand U7027 (N_7027,N_4780,N_4966);
nand U7028 (N_7028,N_5350,N_5416);
and U7029 (N_7029,N_4519,N_3741);
and U7030 (N_7030,N_5493,N_4506);
or U7031 (N_7031,N_4047,N_5305);
xor U7032 (N_7032,N_4920,N_3427);
xnor U7033 (N_7033,N_4952,N_5900);
nand U7034 (N_7034,N_4553,N_4086);
and U7035 (N_7035,N_5364,N_5736);
xor U7036 (N_7036,N_4590,N_5546);
nor U7037 (N_7037,N_3035,N_4023);
and U7038 (N_7038,N_5035,N_5867);
nor U7039 (N_7039,N_3886,N_4827);
nor U7040 (N_7040,N_4799,N_4749);
xnor U7041 (N_7041,N_5485,N_5834);
or U7042 (N_7042,N_4216,N_5271);
or U7043 (N_7043,N_3022,N_4888);
and U7044 (N_7044,N_3993,N_5027);
nor U7045 (N_7045,N_3966,N_3032);
nand U7046 (N_7046,N_5055,N_5393);
xnor U7047 (N_7047,N_5081,N_5177);
nand U7048 (N_7048,N_3184,N_5972);
or U7049 (N_7049,N_5004,N_4805);
or U7050 (N_7050,N_5381,N_5126);
nor U7051 (N_7051,N_3423,N_5231);
nor U7052 (N_7052,N_5372,N_5898);
nor U7053 (N_7053,N_4711,N_3593);
nor U7054 (N_7054,N_4339,N_5259);
nand U7055 (N_7055,N_5770,N_4745);
or U7056 (N_7056,N_3840,N_5863);
nor U7057 (N_7057,N_4240,N_5806);
nand U7058 (N_7058,N_3002,N_4788);
and U7059 (N_7059,N_3845,N_4710);
and U7060 (N_7060,N_4480,N_3867);
and U7061 (N_7061,N_5257,N_3524);
nand U7062 (N_7062,N_4971,N_5141);
nand U7063 (N_7063,N_5316,N_4282);
xor U7064 (N_7064,N_3054,N_5447);
and U7065 (N_7065,N_3786,N_3297);
nor U7066 (N_7066,N_4105,N_4649);
and U7067 (N_7067,N_3618,N_3728);
nor U7068 (N_7068,N_3729,N_4390);
and U7069 (N_7069,N_3014,N_3947);
nand U7070 (N_7070,N_5395,N_5526);
or U7071 (N_7071,N_3817,N_4588);
and U7072 (N_7072,N_4297,N_3499);
nand U7073 (N_7073,N_4874,N_3295);
nand U7074 (N_7074,N_3923,N_4955);
nor U7075 (N_7075,N_5998,N_4245);
nor U7076 (N_7076,N_3554,N_5120);
nor U7077 (N_7077,N_4266,N_5230);
nand U7078 (N_7078,N_5104,N_4924);
nand U7079 (N_7079,N_4473,N_3271);
or U7080 (N_7080,N_5921,N_5848);
or U7081 (N_7081,N_3625,N_4957);
or U7082 (N_7082,N_4666,N_4696);
or U7083 (N_7083,N_4165,N_5667);
nor U7084 (N_7084,N_5626,N_4174);
and U7085 (N_7085,N_4080,N_5317);
and U7086 (N_7086,N_5417,N_4028);
nand U7087 (N_7087,N_4779,N_5838);
nor U7088 (N_7088,N_3735,N_5858);
nor U7089 (N_7089,N_5565,N_3346);
and U7090 (N_7090,N_3970,N_5067);
or U7091 (N_7091,N_3280,N_4746);
xnor U7092 (N_7092,N_4850,N_3931);
or U7093 (N_7093,N_4531,N_4012);
nand U7094 (N_7094,N_3610,N_4225);
nor U7095 (N_7095,N_3898,N_5190);
nand U7096 (N_7096,N_3109,N_5503);
xor U7097 (N_7097,N_4454,N_5444);
xnor U7098 (N_7098,N_3477,N_5345);
nand U7099 (N_7099,N_5601,N_5191);
and U7100 (N_7100,N_3773,N_3877);
and U7101 (N_7101,N_5535,N_3169);
and U7102 (N_7102,N_3630,N_5668);
nor U7103 (N_7103,N_4272,N_3279);
or U7104 (N_7104,N_3913,N_5874);
nor U7105 (N_7105,N_4542,N_4489);
or U7106 (N_7106,N_5013,N_3901);
or U7107 (N_7107,N_3230,N_5987);
xor U7108 (N_7108,N_5133,N_4897);
nor U7109 (N_7109,N_3884,N_4455);
nor U7110 (N_7110,N_5976,N_4223);
nor U7111 (N_7111,N_4566,N_4435);
and U7112 (N_7112,N_4378,N_5855);
or U7113 (N_7113,N_4740,N_4203);
nor U7114 (N_7114,N_4041,N_5491);
and U7115 (N_7115,N_3580,N_5103);
or U7116 (N_7116,N_4653,N_5270);
and U7117 (N_7117,N_3885,N_5048);
nand U7118 (N_7118,N_3837,N_3143);
or U7119 (N_7119,N_4309,N_3527);
nor U7120 (N_7120,N_4134,N_3149);
and U7121 (N_7121,N_4712,N_4477);
nor U7122 (N_7122,N_3206,N_4188);
or U7123 (N_7123,N_4246,N_4384);
xnor U7124 (N_7124,N_4555,N_3663);
and U7125 (N_7125,N_4016,N_5992);
and U7126 (N_7126,N_5934,N_3608);
nor U7127 (N_7127,N_3249,N_5326);
or U7128 (N_7128,N_5636,N_5008);
and U7129 (N_7129,N_5250,N_5571);
nand U7130 (N_7130,N_5074,N_4738);
nand U7131 (N_7131,N_3848,N_5406);
and U7132 (N_7132,N_5426,N_5925);
and U7133 (N_7133,N_4048,N_4071);
and U7134 (N_7134,N_5852,N_5359);
or U7135 (N_7135,N_4065,N_3240);
nor U7136 (N_7136,N_5043,N_3235);
and U7137 (N_7137,N_5015,N_5885);
and U7138 (N_7138,N_3921,N_5726);
and U7139 (N_7139,N_4144,N_5583);
nor U7140 (N_7140,N_3809,N_5199);
or U7141 (N_7141,N_5738,N_3594);
nand U7142 (N_7142,N_4316,N_5675);
nand U7143 (N_7143,N_5673,N_3597);
or U7144 (N_7144,N_5849,N_4288);
xor U7145 (N_7145,N_4248,N_3129);
nor U7146 (N_7146,N_5688,N_3994);
nor U7147 (N_7147,N_4232,N_3667);
nor U7148 (N_7148,N_3785,N_5882);
and U7149 (N_7149,N_4291,N_5066);
nand U7150 (N_7150,N_4433,N_5818);
nor U7151 (N_7151,N_4655,N_3717);
xor U7152 (N_7152,N_4353,N_4985);
nor U7153 (N_7153,N_3868,N_3616);
nand U7154 (N_7154,N_3528,N_5913);
and U7155 (N_7155,N_5196,N_5983);
or U7156 (N_7156,N_5188,N_3147);
nor U7157 (N_7157,N_4671,N_5949);
nand U7158 (N_7158,N_5349,N_5089);
nand U7159 (N_7159,N_3784,N_5564);
and U7160 (N_7160,N_3915,N_3300);
and U7161 (N_7161,N_4345,N_4837);
nor U7162 (N_7162,N_5492,N_4373);
nand U7163 (N_7163,N_3772,N_5892);
or U7164 (N_7164,N_5445,N_3957);
nand U7165 (N_7165,N_5664,N_3166);
nand U7166 (N_7166,N_5719,N_4945);
nor U7167 (N_7167,N_3444,N_5370);
nor U7168 (N_7168,N_4348,N_4816);
nand U7169 (N_7169,N_5929,N_5610);
nor U7170 (N_7170,N_3355,N_3111);
and U7171 (N_7171,N_3108,N_3461);
nor U7172 (N_7172,N_5978,N_5876);
or U7173 (N_7173,N_4337,N_3484);
xnor U7174 (N_7174,N_5366,N_4810);
and U7175 (N_7175,N_5278,N_3282);
and U7176 (N_7176,N_3875,N_4443);
or U7177 (N_7177,N_3812,N_4419);
nand U7178 (N_7178,N_3000,N_5380);
or U7179 (N_7179,N_5666,N_5367);
xnor U7180 (N_7180,N_4736,N_5496);
nor U7181 (N_7181,N_3977,N_3907);
xor U7182 (N_7182,N_5085,N_3706);
and U7183 (N_7183,N_3714,N_3317);
nand U7184 (N_7184,N_3925,N_4259);
nand U7185 (N_7185,N_3953,N_4631);
nor U7186 (N_7186,N_4098,N_4547);
nand U7187 (N_7187,N_4852,N_3470);
nor U7188 (N_7188,N_3486,N_4472);
and U7189 (N_7189,N_4496,N_4162);
xor U7190 (N_7190,N_4385,N_4005);
xnor U7191 (N_7191,N_4178,N_3864);
or U7192 (N_7192,N_5148,N_5889);
nor U7193 (N_7193,N_3747,N_4839);
nor U7194 (N_7194,N_4831,N_4210);
nor U7195 (N_7195,N_5174,N_3337);
nor U7196 (N_7196,N_4875,N_4818);
nand U7197 (N_7197,N_3270,N_4184);
nand U7198 (N_7198,N_3197,N_3797);
or U7199 (N_7199,N_3181,N_4024);
or U7200 (N_7200,N_5864,N_3429);
nor U7201 (N_7201,N_5651,N_4910);
xnor U7202 (N_7202,N_4689,N_3730);
nand U7203 (N_7203,N_5620,N_3780);
nand U7204 (N_7204,N_4199,N_3935);
nand U7205 (N_7205,N_3976,N_3822);
and U7206 (N_7206,N_4625,N_3589);
nor U7207 (N_7207,N_4082,N_5743);
nand U7208 (N_7208,N_3537,N_5229);
and U7209 (N_7209,N_5702,N_5263);
or U7210 (N_7210,N_3638,N_5042);
nand U7211 (N_7211,N_4387,N_4260);
nor U7212 (N_7212,N_5935,N_4056);
or U7213 (N_7213,N_5721,N_3241);
or U7214 (N_7214,N_4325,N_5468);
nor U7215 (N_7215,N_3843,N_5760);
nor U7216 (N_7216,N_5794,N_3945);
xor U7217 (N_7217,N_5324,N_4383);
nor U7218 (N_7218,N_3269,N_4097);
and U7219 (N_7219,N_4315,N_5761);
nand U7220 (N_7220,N_4721,N_5127);
nor U7221 (N_7221,N_4319,N_4401);
or U7222 (N_7222,N_3291,N_3216);
or U7223 (N_7223,N_5952,N_5883);
or U7224 (N_7224,N_4476,N_4605);
and U7225 (N_7225,N_4336,N_3199);
xnor U7226 (N_7226,N_5762,N_5214);
xor U7227 (N_7227,N_5635,N_4943);
or U7228 (N_7228,N_3558,N_5866);
nand U7229 (N_7229,N_4446,N_4914);
or U7230 (N_7230,N_5959,N_4792);
and U7231 (N_7231,N_5909,N_5901);
nand U7232 (N_7232,N_4106,N_4798);
nor U7233 (N_7233,N_3200,N_5005);
and U7234 (N_7234,N_3956,N_4545);
nor U7235 (N_7235,N_3869,N_5958);
xnor U7236 (N_7236,N_5483,N_4283);
and U7237 (N_7237,N_4046,N_4682);
nand U7238 (N_7238,N_3178,N_4675);
xor U7239 (N_7239,N_4849,N_3020);
or U7240 (N_7240,N_3102,N_4869);
nand U7241 (N_7241,N_5283,N_3222);
nand U7242 (N_7242,N_3609,N_5791);
and U7243 (N_7243,N_3247,N_3536);
and U7244 (N_7244,N_4054,N_4037);
or U7245 (N_7245,N_4561,N_4753);
and U7246 (N_7246,N_3258,N_4731);
or U7247 (N_7247,N_3069,N_5879);
xnor U7248 (N_7248,N_4394,N_5502);
nand U7249 (N_7249,N_3128,N_4375);
and U7250 (N_7250,N_4923,N_5459);
and U7251 (N_7251,N_5938,N_5315);
and U7252 (N_7252,N_5354,N_5532);
nand U7253 (N_7253,N_4020,N_4275);
and U7254 (N_7254,N_5559,N_3207);
or U7255 (N_7255,N_4265,N_5451);
nand U7256 (N_7256,N_3553,N_3356);
nor U7257 (N_7257,N_3839,N_5236);
xnor U7258 (N_7258,N_4500,N_4572);
nand U7259 (N_7259,N_5158,N_5407);
or U7260 (N_7260,N_4530,N_3932);
nor U7261 (N_7261,N_5710,N_4305);
nand U7262 (N_7262,N_3782,N_4800);
xnor U7263 (N_7263,N_3454,N_5203);
nor U7264 (N_7264,N_3202,N_3680);
or U7265 (N_7265,N_3298,N_4388);
or U7266 (N_7266,N_4669,N_5038);
or U7267 (N_7267,N_3483,N_4461);
nor U7268 (N_7268,N_5176,N_4620);
and U7269 (N_7269,N_5814,N_5803);
or U7270 (N_7270,N_5115,N_3095);
nor U7271 (N_7271,N_3731,N_5621);
nand U7272 (N_7272,N_4867,N_3229);
xnor U7273 (N_7273,N_3619,N_5182);
and U7274 (N_7274,N_5857,N_3335);
nand U7275 (N_7275,N_5878,N_3193);
xor U7276 (N_7276,N_5595,N_5941);
or U7277 (N_7277,N_5833,N_3196);
and U7278 (N_7278,N_3459,N_5078);
nor U7279 (N_7279,N_4009,N_5643);
or U7280 (N_7280,N_3083,N_5100);
xnor U7281 (N_7281,N_5400,N_3588);
nor U7282 (N_7282,N_3120,N_5588);
nand U7283 (N_7283,N_3305,N_4960);
or U7284 (N_7284,N_5272,N_3284);
or U7285 (N_7285,N_4312,N_3392);
or U7286 (N_7286,N_4549,N_4979);
nand U7287 (N_7287,N_5641,N_5146);
and U7288 (N_7288,N_3924,N_4285);
nand U7289 (N_7289,N_5562,N_4823);
nor U7290 (N_7290,N_3148,N_3612);
and U7291 (N_7291,N_3750,N_4081);
nor U7292 (N_7292,N_4717,N_3451);
and U7293 (N_7293,N_5633,N_4290);
and U7294 (N_7294,N_5860,N_5034);
or U7295 (N_7295,N_4151,N_4027);
nor U7296 (N_7296,N_5123,N_3596);
and U7297 (N_7297,N_4150,N_4889);
xor U7298 (N_7298,N_5138,N_5300);
nor U7299 (N_7299,N_4857,N_3475);
nor U7300 (N_7300,N_3621,N_4596);
nand U7301 (N_7301,N_5534,N_5713);
nand U7302 (N_7302,N_3752,N_3441);
or U7303 (N_7303,N_4525,N_5575);
or U7304 (N_7304,N_5193,N_3089);
nand U7305 (N_7305,N_5180,N_5132);
and U7306 (N_7306,N_4330,N_3911);
nand U7307 (N_7307,N_3208,N_4204);
or U7308 (N_7308,N_4781,N_3575);
nor U7309 (N_7309,N_5258,N_3572);
or U7310 (N_7310,N_5260,N_3791);
nor U7311 (N_7311,N_5045,N_4361);
nor U7312 (N_7312,N_3494,N_5186);
nor U7313 (N_7313,N_4033,N_4132);
and U7314 (N_7314,N_4197,N_5473);
nand U7315 (N_7315,N_3065,N_5304);
xor U7316 (N_7316,N_4863,N_5287);
nand U7317 (N_7317,N_5343,N_4182);
or U7318 (N_7318,N_4982,N_4329);
or U7319 (N_7319,N_5731,N_4652);
and U7320 (N_7320,N_3999,N_5527);
nor U7321 (N_7321,N_5044,N_4834);
or U7322 (N_7322,N_4287,N_3219);
xnor U7323 (N_7323,N_5484,N_4125);
or U7324 (N_7324,N_5198,N_5338);
or U7325 (N_7325,N_4538,N_3979);
nand U7326 (N_7326,N_3896,N_5630);
xor U7327 (N_7327,N_3807,N_4062);
nand U7328 (N_7328,N_5415,N_5478);
nor U7329 (N_7329,N_5294,N_5775);
and U7330 (N_7330,N_4254,N_4269);
or U7331 (N_7331,N_4866,N_5530);
nand U7332 (N_7332,N_5238,N_5047);
and U7333 (N_7333,N_4748,N_3390);
or U7334 (N_7334,N_4825,N_5409);
and U7335 (N_7335,N_5859,N_3879);
and U7336 (N_7336,N_5439,N_5528);
xnor U7337 (N_7337,N_3299,N_5088);
and U7338 (N_7338,N_3695,N_5598);
or U7339 (N_7339,N_4554,N_4255);
or U7340 (N_7340,N_5059,N_5421);
or U7341 (N_7341,N_4306,N_4802);
nand U7342 (N_7342,N_4835,N_5061);
nor U7343 (N_7343,N_4346,N_4617);
nor U7344 (N_7344,N_3650,N_4176);
and U7345 (N_7345,N_3697,N_3164);
nor U7346 (N_7346,N_5137,N_5109);
xor U7347 (N_7347,N_3367,N_4754);
and U7348 (N_7348,N_4351,N_3313);
and U7349 (N_7349,N_3038,N_4893);
xnor U7350 (N_7350,N_5656,N_3990);
or U7351 (N_7351,N_4529,N_4310);
nor U7352 (N_7352,N_3473,N_3722);
or U7353 (N_7353,N_3991,N_3557);
nand U7354 (N_7354,N_3642,N_3378);
xnor U7355 (N_7355,N_3852,N_5741);
nor U7356 (N_7356,N_5092,N_3666);
or U7357 (N_7357,N_5862,N_4932);
and U7358 (N_7358,N_4235,N_4100);
and U7359 (N_7359,N_4674,N_4257);
nor U7360 (N_7360,N_5219,N_3464);
and U7361 (N_7361,N_3236,N_4829);
or U7362 (N_7362,N_5572,N_5798);
nor U7363 (N_7363,N_4163,N_3878);
nor U7364 (N_7364,N_3191,N_5296);
and U7365 (N_7365,N_4089,N_3988);
and U7366 (N_7366,N_3751,N_4471);
nand U7367 (N_7367,N_3474,N_5441);
nand U7368 (N_7368,N_4488,N_5953);
and U7369 (N_7369,N_4949,N_5293);
and U7370 (N_7370,N_5977,N_4546);
and U7371 (N_7371,N_5507,N_3107);
nand U7372 (N_7372,N_4836,N_5542);
nand U7373 (N_7373,N_4936,N_5280);
and U7374 (N_7374,N_3433,N_4681);
and U7375 (N_7375,N_4938,N_3133);
and U7376 (N_7376,N_3072,N_5204);
and U7377 (N_7377,N_3549,N_3435);
or U7378 (N_7378,N_3904,N_5923);
xnor U7379 (N_7379,N_3005,N_4690);
and U7380 (N_7380,N_3341,N_5113);
and U7381 (N_7381,N_5217,N_3876);
nand U7382 (N_7382,N_3691,N_5033);
or U7383 (N_7383,N_4350,N_5079);
nor U7384 (N_7384,N_4423,N_5265);
and U7385 (N_7385,N_3463,N_3103);
and U7386 (N_7386,N_3381,N_4886);
nor U7387 (N_7387,N_4882,N_3505);
nand U7388 (N_7388,N_5077,N_5046);
nor U7389 (N_7389,N_3078,N_3130);
xor U7390 (N_7390,N_3595,N_4442);
and U7391 (N_7391,N_3344,N_3930);
or U7392 (N_7392,N_4956,N_4534);
and U7393 (N_7393,N_4708,N_3949);
and U7394 (N_7394,N_5594,N_4700);
nand U7395 (N_7395,N_3985,N_5906);
and U7396 (N_7396,N_3656,N_3401);
xor U7397 (N_7397,N_4766,N_5578);
and U7398 (N_7398,N_4908,N_5632);
nand U7399 (N_7399,N_4929,N_4487);
nand U7400 (N_7400,N_5893,N_5335);
nand U7401 (N_7401,N_5647,N_5097);
xor U7402 (N_7402,N_3748,N_5912);
nand U7403 (N_7403,N_3776,N_5363);
nand U7404 (N_7404,N_3081,N_3027);
or U7405 (N_7405,N_4393,N_5117);
nor U7406 (N_7406,N_3962,N_5461);
nor U7407 (N_7407,N_5751,N_4718);
nand U7408 (N_7408,N_4400,N_5709);
xor U7409 (N_7409,N_3865,N_4814);
nor U7410 (N_7410,N_3366,N_4726);
nor U7411 (N_7411,N_5460,N_3412);
or U7412 (N_7412,N_3393,N_5671);
or U7413 (N_7413,N_5654,N_4521);
nor U7414 (N_7414,N_3311,N_3789);
and U7415 (N_7415,N_3684,N_4481);
nor U7416 (N_7416,N_4612,N_3192);
or U7417 (N_7417,N_4352,N_4354);
and U7418 (N_7418,N_5058,N_4513);
nor U7419 (N_7419,N_3900,N_5140);
xor U7420 (N_7420,N_5839,N_4733);
or U7421 (N_7421,N_3936,N_4855);
or U7422 (N_7422,N_3761,N_3939);
or U7423 (N_7423,N_3286,N_4786);
and U7424 (N_7424,N_3289,N_3017);
nor U7425 (N_7425,N_5290,N_5403);
and U7426 (N_7426,N_5802,N_3617);
nor U7427 (N_7427,N_5373,N_5531);
nor U7428 (N_7428,N_3511,N_3653);
nand U7429 (N_7429,N_3525,N_5948);
xnor U7430 (N_7430,N_3765,N_3112);
and U7431 (N_7431,N_4701,N_4763);
nand U7432 (N_7432,N_4986,N_5711);
xor U7433 (N_7433,N_3634,N_3318);
xor U7434 (N_7434,N_5206,N_4606);
xor U7435 (N_7435,N_5365,N_5997);
and U7436 (N_7436,N_4101,N_4732);
and U7437 (N_7437,N_4646,N_5776);
and U7438 (N_7438,N_3624,N_4398);
nor U7439 (N_7439,N_4535,N_5581);
xor U7440 (N_7440,N_4585,N_5072);
and U7441 (N_7441,N_5128,N_5577);
and U7442 (N_7442,N_5291,N_3029);
and U7443 (N_7443,N_5299,N_5926);
nor U7444 (N_7444,N_3336,N_5431);
and U7445 (N_7445,N_5360,N_4456);
nor U7446 (N_7446,N_3501,N_5545);
xnor U7447 (N_7447,N_5352,N_5486);
nand U7448 (N_7448,N_4528,N_5940);
xnor U7449 (N_7449,N_5358,N_5336);
nor U7450 (N_7450,N_3938,N_3493);
xor U7451 (N_7451,N_5916,N_4043);
or U7452 (N_7452,N_3833,N_4001);
nand U7453 (N_7453,N_3031,N_5877);
or U7454 (N_7454,N_4019,N_4128);
or U7455 (N_7455,N_5003,N_3211);
nor U7456 (N_7456,N_4524,N_4614);
and U7457 (N_7457,N_4498,N_5973);
and U7458 (N_7458,N_5662,N_4092);
and U7459 (N_7459,N_3215,N_4619);
or U7460 (N_7460,N_5540,N_3308);
nand U7461 (N_7461,N_4250,N_5576);
and U7462 (N_7462,N_5218,N_3146);
nand U7463 (N_7463,N_5497,N_5276);
and U7464 (N_7464,N_5533,N_5811);
or U7465 (N_7465,N_3951,N_4050);
nor U7466 (N_7466,N_5110,N_5555);
or U7467 (N_7467,N_3788,N_4374);
nand U7468 (N_7468,N_3316,N_5216);
nand U7469 (N_7469,N_4598,N_4133);
or U7470 (N_7470,N_3061,N_4643);
nand U7471 (N_7471,N_5197,N_5353);
or U7472 (N_7472,N_5273,N_4457);
nor U7473 (N_7473,N_3611,N_5512);
and U7474 (N_7474,N_4129,N_3333);
or U7475 (N_7475,N_3252,N_4930);
nand U7476 (N_7476,N_5599,N_5472);
or U7477 (N_7477,N_5515,N_3758);
and U7478 (N_7478,N_4220,N_4342);
nor U7479 (N_7479,N_3534,N_5692);
nor U7480 (N_7480,N_4399,N_3214);
xnor U7481 (N_7481,N_3829,N_4116);
xnor U7482 (N_7482,N_3644,N_5480);
or U7483 (N_7483,N_4328,N_4360);
nand U7484 (N_7484,N_4856,N_3846);
or U7485 (N_7485,N_4426,N_5946);
and U7486 (N_7486,N_5020,N_4219);
or U7487 (N_7487,N_3104,N_4698);
nand U7488 (N_7488,N_4630,N_3971);
nor U7489 (N_7489,N_5266,N_4935);
and U7490 (N_7490,N_5690,N_4870);
nor U7491 (N_7491,N_4584,N_3928);
or U7492 (N_7492,N_5954,N_3097);
nor U7493 (N_7493,N_3591,N_5474);
nand U7494 (N_7494,N_5235,N_4007);
xor U7495 (N_7495,N_5831,N_5261);
nand U7496 (N_7496,N_5052,N_4587);
xnor U7497 (N_7497,N_4772,N_5837);
or U7498 (N_7498,N_3673,N_5592);
nand U7499 (N_7499,N_4402,N_5083);
or U7500 (N_7500,N_3248,N_3690);
nand U7501 (N_7501,N_5069,N_5390);
xnor U7502 (N_7502,N_5647,N_3066);
and U7503 (N_7503,N_5815,N_4406);
nor U7504 (N_7504,N_5316,N_3214);
nor U7505 (N_7505,N_5838,N_5446);
nand U7506 (N_7506,N_3406,N_3553);
nand U7507 (N_7507,N_3204,N_3968);
nor U7508 (N_7508,N_4893,N_5183);
or U7509 (N_7509,N_4051,N_3804);
or U7510 (N_7510,N_3252,N_4387);
and U7511 (N_7511,N_5525,N_3193);
or U7512 (N_7512,N_3088,N_3093);
nand U7513 (N_7513,N_5617,N_4250);
nor U7514 (N_7514,N_3395,N_5881);
nand U7515 (N_7515,N_4277,N_5790);
xnor U7516 (N_7516,N_3293,N_4480);
or U7517 (N_7517,N_3045,N_5721);
and U7518 (N_7518,N_4059,N_3386);
nor U7519 (N_7519,N_3447,N_5287);
or U7520 (N_7520,N_5147,N_4547);
or U7521 (N_7521,N_3236,N_5942);
or U7522 (N_7522,N_3646,N_5265);
and U7523 (N_7523,N_4494,N_4716);
nor U7524 (N_7524,N_3718,N_5708);
nand U7525 (N_7525,N_4278,N_5809);
nor U7526 (N_7526,N_3689,N_3823);
nand U7527 (N_7527,N_3224,N_3573);
nand U7528 (N_7528,N_5448,N_4639);
xor U7529 (N_7529,N_4670,N_4459);
and U7530 (N_7530,N_4958,N_5515);
and U7531 (N_7531,N_4744,N_4141);
nor U7532 (N_7532,N_3774,N_3697);
nor U7533 (N_7533,N_5288,N_3854);
nand U7534 (N_7534,N_3480,N_3930);
nor U7535 (N_7535,N_4103,N_5635);
nor U7536 (N_7536,N_4992,N_3320);
and U7537 (N_7537,N_5607,N_5355);
or U7538 (N_7538,N_5967,N_5066);
nor U7539 (N_7539,N_3182,N_3950);
nor U7540 (N_7540,N_3447,N_3917);
xnor U7541 (N_7541,N_3313,N_4772);
or U7542 (N_7542,N_3397,N_5602);
nor U7543 (N_7543,N_5194,N_3035);
and U7544 (N_7544,N_4225,N_3462);
or U7545 (N_7545,N_3225,N_5072);
xnor U7546 (N_7546,N_5639,N_4975);
or U7547 (N_7547,N_4426,N_5549);
xor U7548 (N_7548,N_4100,N_3985);
nor U7549 (N_7549,N_4785,N_3717);
and U7550 (N_7550,N_5759,N_5154);
and U7551 (N_7551,N_5768,N_4151);
xnor U7552 (N_7552,N_4476,N_4720);
nand U7553 (N_7553,N_4417,N_5623);
nand U7554 (N_7554,N_5122,N_3030);
or U7555 (N_7555,N_5316,N_4572);
nor U7556 (N_7556,N_3324,N_4126);
and U7557 (N_7557,N_3490,N_3923);
nor U7558 (N_7558,N_3814,N_3965);
or U7559 (N_7559,N_5395,N_5114);
nand U7560 (N_7560,N_3551,N_5035);
or U7561 (N_7561,N_3222,N_3929);
nor U7562 (N_7562,N_4354,N_5177);
or U7563 (N_7563,N_4080,N_5431);
and U7564 (N_7564,N_4162,N_4295);
nor U7565 (N_7565,N_3906,N_5797);
nand U7566 (N_7566,N_5103,N_3853);
and U7567 (N_7567,N_3824,N_4672);
and U7568 (N_7568,N_5160,N_3039);
nor U7569 (N_7569,N_4155,N_3071);
xnor U7570 (N_7570,N_5535,N_3673);
xnor U7571 (N_7571,N_4325,N_4810);
nor U7572 (N_7572,N_5253,N_5173);
nor U7573 (N_7573,N_3490,N_4233);
nor U7574 (N_7574,N_3915,N_5969);
or U7575 (N_7575,N_4781,N_5191);
nor U7576 (N_7576,N_4572,N_3782);
and U7577 (N_7577,N_5644,N_5116);
nor U7578 (N_7578,N_4532,N_4304);
nand U7579 (N_7579,N_5150,N_3797);
and U7580 (N_7580,N_5894,N_5557);
or U7581 (N_7581,N_4269,N_4627);
nand U7582 (N_7582,N_3795,N_4016);
xor U7583 (N_7583,N_5251,N_5286);
nand U7584 (N_7584,N_5577,N_3548);
and U7585 (N_7585,N_4668,N_3374);
and U7586 (N_7586,N_4262,N_3951);
nand U7587 (N_7587,N_4090,N_3163);
xnor U7588 (N_7588,N_5769,N_5012);
or U7589 (N_7589,N_5343,N_5172);
xnor U7590 (N_7590,N_3765,N_4707);
nand U7591 (N_7591,N_3967,N_3977);
nand U7592 (N_7592,N_4260,N_5561);
or U7593 (N_7593,N_5567,N_3385);
nand U7594 (N_7594,N_3732,N_3782);
or U7595 (N_7595,N_3782,N_5721);
nand U7596 (N_7596,N_3260,N_5044);
xor U7597 (N_7597,N_3058,N_5374);
xor U7598 (N_7598,N_3957,N_3488);
nor U7599 (N_7599,N_3197,N_5163);
or U7600 (N_7600,N_3111,N_5611);
and U7601 (N_7601,N_4906,N_3821);
or U7602 (N_7602,N_5104,N_3895);
and U7603 (N_7603,N_4929,N_5695);
and U7604 (N_7604,N_3347,N_3911);
or U7605 (N_7605,N_5155,N_4531);
xor U7606 (N_7606,N_4065,N_4391);
nor U7607 (N_7607,N_4554,N_3430);
nor U7608 (N_7608,N_4005,N_5830);
nand U7609 (N_7609,N_3919,N_3543);
nor U7610 (N_7610,N_4417,N_3883);
or U7611 (N_7611,N_5002,N_5313);
nand U7612 (N_7612,N_5581,N_4699);
nor U7613 (N_7613,N_3473,N_3329);
xnor U7614 (N_7614,N_4920,N_5854);
nand U7615 (N_7615,N_5734,N_3331);
or U7616 (N_7616,N_5396,N_4546);
or U7617 (N_7617,N_5279,N_4533);
and U7618 (N_7618,N_5632,N_4452);
or U7619 (N_7619,N_4090,N_5564);
or U7620 (N_7620,N_5681,N_3670);
nor U7621 (N_7621,N_4225,N_3213);
nand U7622 (N_7622,N_3227,N_4452);
nand U7623 (N_7623,N_3980,N_3407);
nand U7624 (N_7624,N_4087,N_3365);
and U7625 (N_7625,N_5343,N_4808);
or U7626 (N_7626,N_5096,N_4141);
nor U7627 (N_7627,N_3972,N_4567);
or U7628 (N_7628,N_4990,N_5390);
and U7629 (N_7629,N_3706,N_4514);
nor U7630 (N_7630,N_5814,N_4947);
nor U7631 (N_7631,N_5025,N_3281);
xor U7632 (N_7632,N_4557,N_5063);
nor U7633 (N_7633,N_4611,N_5395);
nand U7634 (N_7634,N_5865,N_3586);
nor U7635 (N_7635,N_3446,N_5854);
or U7636 (N_7636,N_4514,N_4881);
and U7637 (N_7637,N_4743,N_5503);
nor U7638 (N_7638,N_4667,N_3366);
or U7639 (N_7639,N_4152,N_5730);
and U7640 (N_7640,N_5903,N_3986);
xnor U7641 (N_7641,N_4640,N_3832);
nor U7642 (N_7642,N_3443,N_3922);
xor U7643 (N_7643,N_5185,N_4928);
xnor U7644 (N_7644,N_4179,N_4940);
nor U7645 (N_7645,N_3488,N_4958);
xor U7646 (N_7646,N_3306,N_4298);
nand U7647 (N_7647,N_5544,N_4787);
nor U7648 (N_7648,N_5667,N_4642);
nand U7649 (N_7649,N_3606,N_3226);
xor U7650 (N_7650,N_3887,N_5658);
and U7651 (N_7651,N_4695,N_5799);
or U7652 (N_7652,N_3202,N_5820);
xnor U7653 (N_7653,N_5144,N_4132);
or U7654 (N_7654,N_5487,N_5882);
xnor U7655 (N_7655,N_4497,N_3156);
nor U7656 (N_7656,N_4817,N_5416);
and U7657 (N_7657,N_4159,N_5449);
and U7658 (N_7658,N_5167,N_3274);
nand U7659 (N_7659,N_5140,N_3347);
nor U7660 (N_7660,N_3506,N_4043);
nor U7661 (N_7661,N_4498,N_3173);
and U7662 (N_7662,N_4186,N_5898);
or U7663 (N_7663,N_3442,N_3326);
nand U7664 (N_7664,N_5926,N_4658);
or U7665 (N_7665,N_3648,N_5191);
or U7666 (N_7666,N_5413,N_4802);
and U7667 (N_7667,N_3827,N_4054);
or U7668 (N_7668,N_5240,N_5006);
and U7669 (N_7669,N_4779,N_3081);
or U7670 (N_7670,N_4594,N_3969);
and U7671 (N_7671,N_4815,N_4414);
nand U7672 (N_7672,N_3547,N_3457);
xnor U7673 (N_7673,N_4696,N_3077);
nand U7674 (N_7674,N_5182,N_3152);
xnor U7675 (N_7675,N_5734,N_5859);
or U7676 (N_7676,N_3054,N_5454);
or U7677 (N_7677,N_5177,N_5155);
and U7678 (N_7678,N_3361,N_4047);
and U7679 (N_7679,N_3984,N_3909);
nor U7680 (N_7680,N_5610,N_5255);
or U7681 (N_7681,N_3243,N_5578);
nand U7682 (N_7682,N_5100,N_3424);
nor U7683 (N_7683,N_3068,N_3701);
nor U7684 (N_7684,N_4219,N_5182);
or U7685 (N_7685,N_5738,N_5476);
nor U7686 (N_7686,N_4696,N_3109);
or U7687 (N_7687,N_3446,N_5049);
and U7688 (N_7688,N_5146,N_3488);
and U7689 (N_7689,N_3899,N_5421);
nand U7690 (N_7690,N_5304,N_4752);
nand U7691 (N_7691,N_5463,N_3379);
xor U7692 (N_7692,N_3950,N_3053);
or U7693 (N_7693,N_5375,N_4232);
or U7694 (N_7694,N_3776,N_3391);
nand U7695 (N_7695,N_3412,N_4270);
and U7696 (N_7696,N_4383,N_3472);
or U7697 (N_7697,N_5891,N_3060);
or U7698 (N_7698,N_4432,N_5454);
and U7699 (N_7699,N_3105,N_4870);
or U7700 (N_7700,N_4927,N_5282);
and U7701 (N_7701,N_3013,N_5233);
nor U7702 (N_7702,N_5433,N_4513);
xnor U7703 (N_7703,N_4894,N_3129);
or U7704 (N_7704,N_5895,N_3870);
nand U7705 (N_7705,N_3607,N_4256);
and U7706 (N_7706,N_3964,N_4960);
nor U7707 (N_7707,N_5183,N_4234);
xor U7708 (N_7708,N_5878,N_3715);
nor U7709 (N_7709,N_5277,N_4109);
nor U7710 (N_7710,N_3103,N_5264);
nand U7711 (N_7711,N_5061,N_3344);
xor U7712 (N_7712,N_4409,N_5362);
nor U7713 (N_7713,N_3505,N_5881);
nor U7714 (N_7714,N_4043,N_5538);
or U7715 (N_7715,N_4942,N_5307);
or U7716 (N_7716,N_5161,N_5155);
nand U7717 (N_7717,N_3452,N_5670);
nor U7718 (N_7718,N_5908,N_5927);
or U7719 (N_7719,N_4859,N_5862);
nor U7720 (N_7720,N_3560,N_5711);
and U7721 (N_7721,N_3984,N_3466);
or U7722 (N_7722,N_3309,N_3828);
nand U7723 (N_7723,N_5246,N_4265);
and U7724 (N_7724,N_4757,N_3760);
nand U7725 (N_7725,N_4456,N_5642);
nor U7726 (N_7726,N_5608,N_5841);
nor U7727 (N_7727,N_5938,N_4262);
nand U7728 (N_7728,N_5419,N_5135);
xnor U7729 (N_7729,N_3246,N_5428);
or U7730 (N_7730,N_4773,N_3437);
or U7731 (N_7731,N_4125,N_4580);
nor U7732 (N_7732,N_3455,N_4692);
nor U7733 (N_7733,N_4885,N_4131);
nor U7734 (N_7734,N_3698,N_5197);
or U7735 (N_7735,N_5189,N_5147);
or U7736 (N_7736,N_3694,N_4896);
nand U7737 (N_7737,N_4433,N_5055);
nor U7738 (N_7738,N_5768,N_4420);
nand U7739 (N_7739,N_3287,N_5041);
and U7740 (N_7740,N_4079,N_3346);
and U7741 (N_7741,N_3102,N_3409);
xnor U7742 (N_7742,N_3058,N_3221);
nand U7743 (N_7743,N_5467,N_5937);
nand U7744 (N_7744,N_3089,N_3857);
xor U7745 (N_7745,N_5371,N_3688);
nor U7746 (N_7746,N_3449,N_4983);
or U7747 (N_7747,N_4700,N_3547);
and U7748 (N_7748,N_4387,N_3382);
or U7749 (N_7749,N_5317,N_3809);
nand U7750 (N_7750,N_5945,N_5999);
nor U7751 (N_7751,N_4540,N_5389);
nor U7752 (N_7752,N_3386,N_5010);
xnor U7753 (N_7753,N_3035,N_5877);
or U7754 (N_7754,N_5918,N_4878);
nor U7755 (N_7755,N_5119,N_5556);
or U7756 (N_7756,N_3294,N_5930);
nand U7757 (N_7757,N_4318,N_4440);
nor U7758 (N_7758,N_3398,N_3553);
nor U7759 (N_7759,N_4738,N_3105);
nor U7760 (N_7760,N_4252,N_3002);
or U7761 (N_7761,N_3347,N_4262);
and U7762 (N_7762,N_5436,N_5689);
xnor U7763 (N_7763,N_4976,N_4389);
and U7764 (N_7764,N_4182,N_3540);
or U7765 (N_7765,N_3544,N_5742);
and U7766 (N_7766,N_4292,N_3442);
nand U7767 (N_7767,N_3278,N_3649);
nor U7768 (N_7768,N_5197,N_4565);
nor U7769 (N_7769,N_5535,N_4516);
or U7770 (N_7770,N_3275,N_4550);
and U7771 (N_7771,N_5024,N_3840);
nand U7772 (N_7772,N_3588,N_5745);
xor U7773 (N_7773,N_5664,N_3437);
or U7774 (N_7774,N_4805,N_4113);
nor U7775 (N_7775,N_5775,N_4384);
nor U7776 (N_7776,N_5058,N_4813);
xor U7777 (N_7777,N_5170,N_3424);
nand U7778 (N_7778,N_5098,N_4636);
nor U7779 (N_7779,N_5379,N_5378);
and U7780 (N_7780,N_4725,N_3282);
and U7781 (N_7781,N_4846,N_5277);
nor U7782 (N_7782,N_5873,N_5773);
nand U7783 (N_7783,N_3951,N_5356);
and U7784 (N_7784,N_3580,N_3817);
or U7785 (N_7785,N_3148,N_5544);
and U7786 (N_7786,N_4619,N_4006);
and U7787 (N_7787,N_3282,N_5820);
or U7788 (N_7788,N_3730,N_5266);
nand U7789 (N_7789,N_5596,N_5284);
or U7790 (N_7790,N_5114,N_5522);
or U7791 (N_7791,N_5409,N_3932);
nor U7792 (N_7792,N_5498,N_3452);
nor U7793 (N_7793,N_5303,N_5290);
and U7794 (N_7794,N_5790,N_4689);
xor U7795 (N_7795,N_5262,N_4635);
and U7796 (N_7796,N_5475,N_4134);
and U7797 (N_7797,N_5725,N_4445);
and U7798 (N_7798,N_5017,N_3428);
nand U7799 (N_7799,N_5821,N_4586);
xnor U7800 (N_7800,N_5766,N_3731);
and U7801 (N_7801,N_5308,N_3515);
nand U7802 (N_7802,N_3267,N_3920);
xnor U7803 (N_7803,N_3089,N_3619);
nor U7804 (N_7804,N_3247,N_4370);
and U7805 (N_7805,N_3948,N_5644);
nand U7806 (N_7806,N_5902,N_5562);
or U7807 (N_7807,N_3486,N_3480);
nand U7808 (N_7808,N_4850,N_4546);
and U7809 (N_7809,N_3875,N_5510);
nand U7810 (N_7810,N_4558,N_3868);
or U7811 (N_7811,N_5464,N_5344);
nor U7812 (N_7812,N_4489,N_4948);
nand U7813 (N_7813,N_4829,N_4725);
nor U7814 (N_7814,N_5585,N_5481);
nor U7815 (N_7815,N_3927,N_4049);
nand U7816 (N_7816,N_4631,N_4852);
and U7817 (N_7817,N_3546,N_3750);
or U7818 (N_7818,N_5491,N_3907);
nor U7819 (N_7819,N_5685,N_4583);
xnor U7820 (N_7820,N_3594,N_5663);
and U7821 (N_7821,N_3425,N_3732);
nor U7822 (N_7822,N_4121,N_4971);
nor U7823 (N_7823,N_5088,N_5550);
or U7824 (N_7824,N_3034,N_4956);
nand U7825 (N_7825,N_3574,N_3536);
and U7826 (N_7826,N_4150,N_3457);
xor U7827 (N_7827,N_4680,N_5420);
and U7828 (N_7828,N_5074,N_3944);
nand U7829 (N_7829,N_5398,N_5811);
and U7830 (N_7830,N_4861,N_3109);
and U7831 (N_7831,N_5052,N_4619);
and U7832 (N_7832,N_5947,N_5082);
nor U7833 (N_7833,N_3564,N_5614);
and U7834 (N_7834,N_3507,N_3770);
and U7835 (N_7835,N_4841,N_4119);
or U7836 (N_7836,N_3722,N_4149);
nand U7837 (N_7837,N_3561,N_5158);
nand U7838 (N_7838,N_3852,N_4936);
nor U7839 (N_7839,N_3675,N_5506);
nand U7840 (N_7840,N_3764,N_5225);
nor U7841 (N_7841,N_4747,N_3754);
xnor U7842 (N_7842,N_3782,N_3866);
nor U7843 (N_7843,N_5234,N_4594);
xor U7844 (N_7844,N_4416,N_5101);
and U7845 (N_7845,N_5943,N_4346);
xor U7846 (N_7846,N_4473,N_5919);
or U7847 (N_7847,N_3099,N_5659);
and U7848 (N_7848,N_5153,N_5629);
nand U7849 (N_7849,N_5468,N_4414);
xor U7850 (N_7850,N_4457,N_3505);
nand U7851 (N_7851,N_3611,N_3089);
nand U7852 (N_7852,N_3310,N_5032);
nor U7853 (N_7853,N_5005,N_3840);
or U7854 (N_7854,N_5197,N_5371);
nand U7855 (N_7855,N_3348,N_4586);
nor U7856 (N_7856,N_4993,N_5260);
and U7857 (N_7857,N_3345,N_5929);
nand U7858 (N_7858,N_3340,N_4998);
nor U7859 (N_7859,N_3905,N_3359);
xnor U7860 (N_7860,N_5899,N_4248);
and U7861 (N_7861,N_3577,N_5372);
and U7862 (N_7862,N_4830,N_4502);
or U7863 (N_7863,N_4213,N_5985);
nor U7864 (N_7864,N_5692,N_3807);
nor U7865 (N_7865,N_5616,N_3224);
or U7866 (N_7866,N_5113,N_4940);
nor U7867 (N_7867,N_4521,N_5520);
and U7868 (N_7868,N_5897,N_5934);
nand U7869 (N_7869,N_4142,N_3577);
or U7870 (N_7870,N_5131,N_4376);
or U7871 (N_7871,N_4507,N_5900);
and U7872 (N_7872,N_4578,N_4465);
nand U7873 (N_7873,N_5268,N_3332);
and U7874 (N_7874,N_4563,N_4633);
and U7875 (N_7875,N_3635,N_4231);
and U7876 (N_7876,N_4009,N_5324);
and U7877 (N_7877,N_3736,N_5665);
xnor U7878 (N_7878,N_5103,N_4603);
or U7879 (N_7879,N_4405,N_4889);
nor U7880 (N_7880,N_5787,N_5177);
or U7881 (N_7881,N_5778,N_5798);
or U7882 (N_7882,N_3153,N_3952);
xor U7883 (N_7883,N_4613,N_4421);
nand U7884 (N_7884,N_5931,N_5651);
and U7885 (N_7885,N_3862,N_4966);
nor U7886 (N_7886,N_4905,N_4222);
and U7887 (N_7887,N_3617,N_5829);
and U7888 (N_7888,N_3297,N_4149);
nor U7889 (N_7889,N_4121,N_5676);
nand U7890 (N_7890,N_5731,N_5468);
nor U7891 (N_7891,N_4357,N_5618);
or U7892 (N_7892,N_4355,N_3391);
nor U7893 (N_7893,N_3830,N_4923);
and U7894 (N_7894,N_3020,N_4190);
and U7895 (N_7895,N_5675,N_3158);
and U7896 (N_7896,N_5941,N_5005);
nor U7897 (N_7897,N_4861,N_3674);
nand U7898 (N_7898,N_4563,N_4202);
nor U7899 (N_7899,N_3818,N_4235);
or U7900 (N_7900,N_4409,N_3433);
nand U7901 (N_7901,N_4247,N_5146);
nor U7902 (N_7902,N_3503,N_5938);
nand U7903 (N_7903,N_4652,N_5649);
nand U7904 (N_7904,N_5725,N_4595);
and U7905 (N_7905,N_4530,N_4715);
or U7906 (N_7906,N_4481,N_5027);
nand U7907 (N_7907,N_4856,N_3355);
nor U7908 (N_7908,N_3352,N_5507);
nor U7909 (N_7909,N_3522,N_3415);
nor U7910 (N_7910,N_5824,N_5607);
and U7911 (N_7911,N_4987,N_5330);
and U7912 (N_7912,N_3209,N_5718);
and U7913 (N_7913,N_3284,N_5762);
or U7914 (N_7914,N_3677,N_5116);
nor U7915 (N_7915,N_5813,N_3306);
or U7916 (N_7916,N_3774,N_4783);
nor U7917 (N_7917,N_3322,N_5633);
nand U7918 (N_7918,N_4684,N_4958);
nor U7919 (N_7919,N_3225,N_4826);
and U7920 (N_7920,N_5835,N_3247);
nand U7921 (N_7921,N_3625,N_3822);
or U7922 (N_7922,N_4857,N_5516);
nand U7923 (N_7923,N_4089,N_5403);
or U7924 (N_7924,N_4042,N_3956);
nand U7925 (N_7925,N_3596,N_3647);
or U7926 (N_7926,N_4438,N_4263);
xnor U7927 (N_7927,N_4778,N_4859);
nand U7928 (N_7928,N_5235,N_4224);
nand U7929 (N_7929,N_3875,N_4860);
nand U7930 (N_7930,N_5001,N_3845);
and U7931 (N_7931,N_5465,N_5122);
or U7932 (N_7932,N_5217,N_4183);
and U7933 (N_7933,N_3183,N_5179);
nand U7934 (N_7934,N_4312,N_4652);
xor U7935 (N_7935,N_3805,N_4817);
and U7936 (N_7936,N_4562,N_5346);
or U7937 (N_7937,N_5544,N_4333);
or U7938 (N_7938,N_5955,N_3334);
nor U7939 (N_7939,N_3676,N_3450);
or U7940 (N_7940,N_5744,N_5464);
nand U7941 (N_7941,N_5494,N_4109);
or U7942 (N_7942,N_4789,N_4936);
nor U7943 (N_7943,N_4956,N_4732);
xnor U7944 (N_7944,N_4566,N_4020);
nor U7945 (N_7945,N_3692,N_5977);
xnor U7946 (N_7946,N_5476,N_5821);
or U7947 (N_7947,N_5039,N_3842);
nand U7948 (N_7948,N_5230,N_5999);
and U7949 (N_7949,N_3076,N_4253);
and U7950 (N_7950,N_5249,N_3885);
and U7951 (N_7951,N_4149,N_3052);
or U7952 (N_7952,N_5784,N_5566);
nor U7953 (N_7953,N_3750,N_4374);
or U7954 (N_7954,N_4722,N_5060);
xnor U7955 (N_7955,N_5390,N_4174);
and U7956 (N_7956,N_3474,N_4315);
xor U7957 (N_7957,N_4026,N_3522);
nand U7958 (N_7958,N_5864,N_3312);
or U7959 (N_7959,N_3535,N_3161);
nand U7960 (N_7960,N_5720,N_4709);
or U7961 (N_7961,N_4930,N_3282);
nor U7962 (N_7962,N_4842,N_5713);
and U7963 (N_7963,N_3994,N_3865);
or U7964 (N_7964,N_4164,N_3302);
nand U7965 (N_7965,N_5311,N_3853);
nand U7966 (N_7966,N_5825,N_5295);
and U7967 (N_7967,N_4941,N_4360);
nor U7968 (N_7968,N_3437,N_4815);
and U7969 (N_7969,N_3779,N_3770);
or U7970 (N_7970,N_5776,N_3674);
and U7971 (N_7971,N_3475,N_5949);
or U7972 (N_7972,N_5014,N_3218);
nor U7973 (N_7973,N_3244,N_5579);
and U7974 (N_7974,N_3381,N_4713);
or U7975 (N_7975,N_3456,N_4587);
xnor U7976 (N_7976,N_3477,N_3150);
nand U7977 (N_7977,N_5870,N_5685);
and U7978 (N_7978,N_4291,N_5159);
nand U7979 (N_7979,N_3261,N_5200);
or U7980 (N_7980,N_3288,N_4825);
nor U7981 (N_7981,N_4165,N_5084);
or U7982 (N_7982,N_3803,N_3607);
or U7983 (N_7983,N_4078,N_5443);
nor U7984 (N_7984,N_5289,N_5268);
or U7985 (N_7985,N_3721,N_3210);
nor U7986 (N_7986,N_3488,N_5503);
or U7987 (N_7987,N_3981,N_4529);
and U7988 (N_7988,N_4489,N_3356);
nand U7989 (N_7989,N_4178,N_3332);
nor U7990 (N_7990,N_4403,N_5524);
nor U7991 (N_7991,N_3380,N_3158);
xnor U7992 (N_7992,N_5210,N_4166);
xor U7993 (N_7993,N_4424,N_4149);
and U7994 (N_7994,N_5194,N_5801);
and U7995 (N_7995,N_5673,N_4750);
or U7996 (N_7996,N_3317,N_4426);
or U7997 (N_7997,N_4959,N_4730);
nand U7998 (N_7998,N_4854,N_5659);
nor U7999 (N_7999,N_4895,N_4870);
or U8000 (N_8000,N_5375,N_3078);
xor U8001 (N_8001,N_4831,N_3759);
and U8002 (N_8002,N_5333,N_3683);
and U8003 (N_8003,N_3260,N_3507);
nor U8004 (N_8004,N_4730,N_3898);
nand U8005 (N_8005,N_5964,N_4396);
xor U8006 (N_8006,N_4833,N_5330);
or U8007 (N_8007,N_4607,N_3188);
nor U8008 (N_8008,N_4198,N_3859);
or U8009 (N_8009,N_4372,N_3144);
or U8010 (N_8010,N_4160,N_5614);
and U8011 (N_8011,N_5850,N_4469);
nand U8012 (N_8012,N_4724,N_3909);
or U8013 (N_8013,N_5933,N_4296);
nand U8014 (N_8014,N_5246,N_3340);
and U8015 (N_8015,N_5332,N_3767);
and U8016 (N_8016,N_3179,N_3032);
and U8017 (N_8017,N_5394,N_5648);
or U8018 (N_8018,N_5499,N_4879);
nand U8019 (N_8019,N_5722,N_5225);
or U8020 (N_8020,N_4321,N_3657);
and U8021 (N_8021,N_3374,N_5224);
nand U8022 (N_8022,N_3443,N_4222);
nand U8023 (N_8023,N_5141,N_5309);
and U8024 (N_8024,N_3894,N_5603);
nand U8025 (N_8025,N_3966,N_3077);
nor U8026 (N_8026,N_3631,N_3798);
nand U8027 (N_8027,N_3910,N_3560);
or U8028 (N_8028,N_4248,N_5070);
or U8029 (N_8029,N_5723,N_5086);
or U8030 (N_8030,N_4040,N_5881);
and U8031 (N_8031,N_4475,N_5859);
or U8032 (N_8032,N_3047,N_3169);
nor U8033 (N_8033,N_5732,N_5508);
xor U8034 (N_8034,N_3843,N_3078);
and U8035 (N_8035,N_5754,N_5392);
nand U8036 (N_8036,N_5225,N_5389);
nand U8037 (N_8037,N_5214,N_5859);
or U8038 (N_8038,N_3953,N_5190);
nand U8039 (N_8039,N_5134,N_4934);
nand U8040 (N_8040,N_5205,N_3483);
nand U8041 (N_8041,N_4234,N_5500);
or U8042 (N_8042,N_5961,N_3355);
or U8043 (N_8043,N_4130,N_4220);
nand U8044 (N_8044,N_3328,N_5853);
and U8045 (N_8045,N_3259,N_4008);
nor U8046 (N_8046,N_5641,N_5411);
nor U8047 (N_8047,N_5946,N_4246);
xnor U8048 (N_8048,N_4856,N_4265);
or U8049 (N_8049,N_4657,N_4522);
and U8050 (N_8050,N_5274,N_5811);
nand U8051 (N_8051,N_4374,N_4811);
and U8052 (N_8052,N_3212,N_5101);
or U8053 (N_8053,N_4164,N_4988);
nand U8054 (N_8054,N_5744,N_5892);
nor U8055 (N_8055,N_3805,N_5290);
nor U8056 (N_8056,N_5309,N_3316);
and U8057 (N_8057,N_3188,N_4453);
and U8058 (N_8058,N_3682,N_3160);
nand U8059 (N_8059,N_5493,N_5016);
nand U8060 (N_8060,N_3049,N_5850);
nand U8061 (N_8061,N_4857,N_4943);
xnor U8062 (N_8062,N_4627,N_3191);
or U8063 (N_8063,N_4612,N_5329);
nor U8064 (N_8064,N_4726,N_4338);
nand U8065 (N_8065,N_3667,N_3616);
nand U8066 (N_8066,N_5187,N_4646);
nor U8067 (N_8067,N_4678,N_4561);
or U8068 (N_8068,N_4766,N_4534);
nor U8069 (N_8069,N_5652,N_5692);
nand U8070 (N_8070,N_3138,N_4351);
nor U8071 (N_8071,N_3800,N_3544);
nor U8072 (N_8072,N_5600,N_5806);
nand U8073 (N_8073,N_5031,N_3742);
and U8074 (N_8074,N_4101,N_3396);
nand U8075 (N_8075,N_5606,N_4838);
xnor U8076 (N_8076,N_3619,N_5041);
and U8077 (N_8077,N_4481,N_3134);
or U8078 (N_8078,N_4036,N_4149);
nor U8079 (N_8079,N_5695,N_3149);
and U8080 (N_8080,N_5087,N_3815);
and U8081 (N_8081,N_5770,N_4031);
and U8082 (N_8082,N_4946,N_4819);
nor U8083 (N_8083,N_3892,N_3826);
nor U8084 (N_8084,N_4727,N_5489);
and U8085 (N_8085,N_5981,N_4328);
or U8086 (N_8086,N_4268,N_5500);
and U8087 (N_8087,N_4351,N_5272);
or U8088 (N_8088,N_3485,N_3693);
nor U8089 (N_8089,N_3133,N_3934);
and U8090 (N_8090,N_4507,N_3796);
xnor U8091 (N_8091,N_3450,N_5775);
nor U8092 (N_8092,N_3572,N_3307);
or U8093 (N_8093,N_4072,N_3172);
or U8094 (N_8094,N_3426,N_5533);
nor U8095 (N_8095,N_5901,N_5930);
or U8096 (N_8096,N_3058,N_4905);
nor U8097 (N_8097,N_4264,N_5423);
or U8098 (N_8098,N_4035,N_5018);
and U8099 (N_8099,N_4673,N_4195);
nand U8100 (N_8100,N_5560,N_4856);
and U8101 (N_8101,N_3943,N_3248);
nand U8102 (N_8102,N_5639,N_4488);
nand U8103 (N_8103,N_5440,N_3136);
nand U8104 (N_8104,N_5964,N_5904);
or U8105 (N_8105,N_3270,N_4335);
and U8106 (N_8106,N_5762,N_5607);
or U8107 (N_8107,N_3042,N_3087);
nor U8108 (N_8108,N_3219,N_3596);
and U8109 (N_8109,N_3355,N_3100);
and U8110 (N_8110,N_5615,N_4703);
nand U8111 (N_8111,N_3247,N_4339);
and U8112 (N_8112,N_5164,N_3209);
xnor U8113 (N_8113,N_3867,N_4771);
xor U8114 (N_8114,N_5195,N_3509);
or U8115 (N_8115,N_5287,N_4518);
nor U8116 (N_8116,N_5102,N_5133);
nand U8117 (N_8117,N_5662,N_4619);
nor U8118 (N_8118,N_5824,N_5577);
nor U8119 (N_8119,N_3087,N_5594);
nand U8120 (N_8120,N_4704,N_5398);
xor U8121 (N_8121,N_3728,N_5507);
and U8122 (N_8122,N_4949,N_3974);
nor U8123 (N_8123,N_4192,N_5398);
nor U8124 (N_8124,N_4003,N_5963);
or U8125 (N_8125,N_5446,N_4708);
and U8126 (N_8126,N_3205,N_5873);
and U8127 (N_8127,N_3786,N_5270);
nor U8128 (N_8128,N_4934,N_5184);
and U8129 (N_8129,N_5402,N_4447);
nor U8130 (N_8130,N_3188,N_4620);
or U8131 (N_8131,N_3549,N_5079);
nor U8132 (N_8132,N_3088,N_3233);
nor U8133 (N_8133,N_5430,N_4088);
and U8134 (N_8134,N_5980,N_4322);
or U8135 (N_8135,N_5870,N_4428);
or U8136 (N_8136,N_5657,N_4980);
or U8137 (N_8137,N_3348,N_5854);
and U8138 (N_8138,N_5960,N_4453);
or U8139 (N_8139,N_4337,N_3727);
nor U8140 (N_8140,N_3718,N_4489);
nand U8141 (N_8141,N_5109,N_3265);
nor U8142 (N_8142,N_3652,N_4913);
and U8143 (N_8143,N_3214,N_5579);
nand U8144 (N_8144,N_4337,N_5046);
or U8145 (N_8145,N_3041,N_4857);
xor U8146 (N_8146,N_5391,N_5238);
xor U8147 (N_8147,N_4992,N_4092);
or U8148 (N_8148,N_4284,N_5773);
nand U8149 (N_8149,N_4250,N_3274);
nor U8150 (N_8150,N_3975,N_3222);
or U8151 (N_8151,N_5076,N_3082);
or U8152 (N_8152,N_3513,N_4863);
nand U8153 (N_8153,N_4721,N_4575);
and U8154 (N_8154,N_5272,N_3840);
nand U8155 (N_8155,N_5142,N_4753);
nor U8156 (N_8156,N_5115,N_4325);
and U8157 (N_8157,N_3989,N_3922);
nand U8158 (N_8158,N_4160,N_4478);
or U8159 (N_8159,N_3576,N_4336);
or U8160 (N_8160,N_5442,N_5859);
or U8161 (N_8161,N_3239,N_5617);
xnor U8162 (N_8162,N_5025,N_5206);
nor U8163 (N_8163,N_4223,N_5553);
nor U8164 (N_8164,N_3808,N_5144);
nor U8165 (N_8165,N_4805,N_3609);
nor U8166 (N_8166,N_4696,N_5678);
nor U8167 (N_8167,N_4912,N_4393);
xnor U8168 (N_8168,N_4955,N_5642);
or U8169 (N_8169,N_3086,N_4877);
xor U8170 (N_8170,N_5014,N_3606);
and U8171 (N_8171,N_3941,N_3820);
nand U8172 (N_8172,N_3541,N_5835);
nor U8173 (N_8173,N_5953,N_3033);
and U8174 (N_8174,N_3303,N_5863);
and U8175 (N_8175,N_4331,N_5012);
nor U8176 (N_8176,N_3528,N_3649);
nand U8177 (N_8177,N_5650,N_5355);
xnor U8178 (N_8178,N_3039,N_5049);
and U8179 (N_8179,N_5601,N_4678);
nor U8180 (N_8180,N_5432,N_4865);
or U8181 (N_8181,N_3632,N_5350);
nor U8182 (N_8182,N_3444,N_3722);
and U8183 (N_8183,N_3414,N_5342);
or U8184 (N_8184,N_5575,N_5686);
nor U8185 (N_8185,N_5138,N_4305);
or U8186 (N_8186,N_3264,N_3186);
nor U8187 (N_8187,N_3688,N_4316);
nor U8188 (N_8188,N_4743,N_5464);
and U8189 (N_8189,N_4131,N_3993);
nand U8190 (N_8190,N_5853,N_5041);
nand U8191 (N_8191,N_3624,N_5884);
nor U8192 (N_8192,N_3236,N_5519);
or U8193 (N_8193,N_4428,N_4409);
or U8194 (N_8194,N_4247,N_4495);
and U8195 (N_8195,N_4898,N_4511);
and U8196 (N_8196,N_4420,N_4521);
xnor U8197 (N_8197,N_5138,N_5609);
nor U8198 (N_8198,N_5551,N_4975);
or U8199 (N_8199,N_4132,N_5552);
nand U8200 (N_8200,N_4001,N_4080);
and U8201 (N_8201,N_4414,N_5370);
or U8202 (N_8202,N_5932,N_3904);
and U8203 (N_8203,N_4492,N_5593);
nor U8204 (N_8204,N_3079,N_3600);
and U8205 (N_8205,N_5626,N_5249);
and U8206 (N_8206,N_5885,N_4895);
nor U8207 (N_8207,N_5400,N_4747);
xnor U8208 (N_8208,N_4880,N_4662);
nand U8209 (N_8209,N_3640,N_4079);
nor U8210 (N_8210,N_4451,N_5337);
nor U8211 (N_8211,N_5440,N_3917);
and U8212 (N_8212,N_4604,N_3774);
nor U8213 (N_8213,N_5289,N_5131);
nand U8214 (N_8214,N_4854,N_4073);
nand U8215 (N_8215,N_4322,N_3821);
xnor U8216 (N_8216,N_3893,N_4384);
and U8217 (N_8217,N_3552,N_5768);
nor U8218 (N_8218,N_3927,N_4804);
nor U8219 (N_8219,N_3190,N_3636);
xnor U8220 (N_8220,N_3638,N_4259);
nor U8221 (N_8221,N_5152,N_4979);
nor U8222 (N_8222,N_3580,N_3067);
or U8223 (N_8223,N_4502,N_3452);
nand U8224 (N_8224,N_4386,N_3335);
nor U8225 (N_8225,N_3063,N_4325);
nand U8226 (N_8226,N_3236,N_4747);
nand U8227 (N_8227,N_4981,N_3910);
nor U8228 (N_8228,N_5830,N_3863);
xnor U8229 (N_8229,N_5924,N_4673);
nor U8230 (N_8230,N_3682,N_3695);
nand U8231 (N_8231,N_3370,N_5924);
and U8232 (N_8232,N_3124,N_5429);
nand U8233 (N_8233,N_3828,N_5801);
nand U8234 (N_8234,N_4874,N_5668);
and U8235 (N_8235,N_4604,N_5405);
nor U8236 (N_8236,N_5026,N_3388);
or U8237 (N_8237,N_5659,N_5203);
or U8238 (N_8238,N_4980,N_3776);
nand U8239 (N_8239,N_5260,N_5981);
nor U8240 (N_8240,N_3157,N_3776);
xnor U8241 (N_8241,N_4286,N_3761);
nand U8242 (N_8242,N_5707,N_3126);
nand U8243 (N_8243,N_3398,N_3064);
nand U8244 (N_8244,N_4107,N_3262);
nor U8245 (N_8245,N_5117,N_3635);
and U8246 (N_8246,N_4024,N_5376);
xor U8247 (N_8247,N_3365,N_5089);
nor U8248 (N_8248,N_4125,N_3033);
and U8249 (N_8249,N_5182,N_5001);
nand U8250 (N_8250,N_5465,N_4284);
nor U8251 (N_8251,N_3140,N_5140);
or U8252 (N_8252,N_4897,N_3365);
nand U8253 (N_8253,N_3008,N_5939);
and U8254 (N_8254,N_4231,N_3397);
and U8255 (N_8255,N_5761,N_3327);
nand U8256 (N_8256,N_3891,N_5432);
or U8257 (N_8257,N_5577,N_4926);
nor U8258 (N_8258,N_3383,N_3487);
and U8259 (N_8259,N_4124,N_5454);
and U8260 (N_8260,N_5485,N_4297);
or U8261 (N_8261,N_4230,N_5646);
nand U8262 (N_8262,N_3158,N_5102);
or U8263 (N_8263,N_4730,N_3621);
and U8264 (N_8264,N_4958,N_4377);
nand U8265 (N_8265,N_5227,N_5063);
and U8266 (N_8266,N_3622,N_5329);
nor U8267 (N_8267,N_3885,N_3181);
xnor U8268 (N_8268,N_5298,N_5664);
or U8269 (N_8269,N_4061,N_5549);
nand U8270 (N_8270,N_4628,N_3552);
xnor U8271 (N_8271,N_3596,N_3773);
nand U8272 (N_8272,N_4895,N_4952);
nand U8273 (N_8273,N_3463,N_4915);
nor U8274 (N_8274,N_4055,N_4870);
and U8275 (N_8275,N_3215,N_4969);
or U8276 (N_8276,N_3830,N_4284);
nand U8277 (N_8277,N_4013,N_3895);
and U8278 (N_8278,N_4950,N_3424);
or U8279 (N_8279,N_5842,N_5884);
nor U8280 (N_8280,N_3058,N_5076);
and U8281 (N_8281,N_3952,N_4947);
nor U8282 (N_8282,N_4829,N_5135);
and U8283 (N_8283,N_5433,N_4542);
or U8284 (N_8284,N_4478,N_5604);
nor U8285 (N_8285,N_5111,N_5375);
nor U8286 (N_8286,N_5172,N_4129);
nand U8287 (N_8287,N_4965,N_3007);
nand U8288 (N_8288,N_5625,N_4270);
or U8289 (N_8289,N_4975,N_5997);
or U8290 (N_8290,N_5740,N_5589);
and U8291 (N_8291,N_4549,N_3976);
nand U8292 (N_8292,N_5856,N_3474);
nand U8293 (N_8293,N_4055,N_3154);
nand U8294 (N_8294,N_5603,N_5050);
xor U8295 (N_8295,N_5952,N_5566);
nor U8296 (N_8296,N_4961,N_5513);
xnor U8297 (N_8297,N_4213,N_3520);
xor U8298 (N_8298,N_5571,N_4097);
nand U8299 (N_8299,N_3312,N_4181);
or U8300 (N_8300,N_4246,N_4712);
nor U8301 (N_8301,N_3353,N_5223);
nor U8302 (N_8302,N_5903,N_5263);
nor U8303 (N_8303,N_3870,N_5792);
nor U8304 (N_8304,N_5444,N_4658);
or U8305 (N_8305,N_3118,N_5738);
nor U8306 (N_8306,N_5118,N_3250);
nor U8307 (N_8307,N_5136,N_3001);
nand U8308 (N_8308,N_4453,N_4534);
and U8309 (N_8309,N_4687,N_4929);
nand U8310 (N_8310,N_5987,N_3952);
and U8311 (N_8311,N_3597,N_3365);
and U8312 (N_8312,N_4453,N_5759);
nand U8313 (N_8313,N_5193,N_4845);
nand U8314 (N_8314,N_5750,N_3853);
nor U8315 (N_8315,N_4588,N_5078);
nor U8316 (N_8316,N_4452,N_5556);
nor U8317 (N_8317,N_5824,N_5467);
nand U8318 (N_8318,N_3625,N_4751);
or U8319 (N_8319,N_3112,N_5761);
nand U8320 (N_8320,N_3294,N_5569);
nor U8321 (N_8321,N_3448,N_3833);
nor U8322 (N_8322,N_4476,N_5245);
and U8323 (N_8323,N_3058,N_5206);
xnor U8324 (N_8324,N_5014,N_3800);
and U8325 (N_8325,N_5905,N_3062);
nand U8326 (N_8326,N_5104,N_5963);
nor U8327 (N_8327,N_4506,N_4706);
or U8328 (N_8328,N_4775,N_5001);
and U8329 (N_8329,N_3798,N_4996);
and U8330 (N_8330,N_3438,N_4632);
xor U8331 (N_8331,N_4808,N_4636);
xnor U8332 (N_8332,N_3347,N_4459);
or U8333 (N_8333,N_4206,N_3885);
and U8334 (N_8334,N_5977,N_4680);
nand U8335 (N_8335,N_3554,N_4146);
or U8336 (N_8336,N_3616,N_5822);
nor U8337 (N_8337,N_3420,N_3533);
or U8338 (N_8338,N_5370,N_5489);
xor U8339 (N_8339,N_3480,N_5866);
or U8340 (N_8340,N_3403,N_3389);
or U8341 (N_8341,N_4484,N_5417);
and U8342 (N_8342,N_4566,N_4255);
nand U8343 (N_8343,N_3815,N_5166);
nand U8344 (N_8344,N_5461,N_3089);
nor U8345 (N_8345,N_4124,N_4712);
or U8346 (N_8346,N_4289,N_3706);
and U8347 (N_8347,N_4850,N_5874);
nand U8348 (N_8348,N_4402,N_3261);
xor U8349 (N_8349,N_3573,N_3389);
and U8350 (N_8350,N_5894,N_4947);
nand U8351 (N_8351,N_3524,N_5275);
or U8352 (N_8352,N_5876,N_3446);
and U8353 (N_8353,N_3403,N_3975);
and U8354 (N_8354,N_4934,N_3812);
or U8355 (N_8355,N_5667,N_4732);
nor U8356 (N_8356,N_4617,N_4056);
nand U8357 (N_8357,N_4397,N_3170);
or U8358 (N_8358,N_5079,N_5644);
or U8359 (N_8359,N_3371,N_4119);
nand U8360 (N_8360,N_4631,N_5637);
or U8361 (N_8361,N_5759,N_4610);
nor U8362 (N_8362,N_3715,N_3637);
nor U8363 (N_8363,N_3599,N_5574);
or U8364 (N_8364,N_5521,N_5127);
or U8365 (N_8365,N_3631,N_3767);
xnor U8366 (N_8366,N_4749,N_4757);
nor U8367 (N_8367,N_3942,N_4608);
or U8368 (N_8368,N_5218,N_5248);
and U8369 (N_8369,N_5579,N_4137);
or U8370 (N_8370,N_5333,N_5317);
nand U8371 (N_8371,N_5634,N_3110);
and U8372 (N_8372,N_3840,N_4720);
or U8373 (N_8373,N_4424,N_5348);
nor U8374 (N_8374,N_5804,N_3428);
or U8375 (N_8375,N_4519,N_3972);
and U8376 (N_8376,N_5897,N_4612);
xnor U8377 (N_8377,N_3884,N_5513);
nand U8378 (N_8378,N_4115,N_3617);
nand U8379 (N_8379,N_5962,N_4429);
xnor U8380 (N_8380,N_3108,N_5527);
or U8381 (N_8381,N_4966,N_5070);
nand U8382 (N_8382,N_3727,N_5502);
nor U8383 (N_8383,N_4228,N_5169);
nor U8384 (N_8384,N_3010,N_3895);
xnor U8385 (N_8385,N_4283,N_4340);
and U8386 (N_8386,N_3681,N_5010);
nor U8387 (N_8387,N_3220,N_4679);
nand U8388 (N_8388,N_3512,N_3598);
nand U8389 (N_8389,N_3848,N_4422);
nor U8390 (N_8390,N_4433,N_5900);
and U8391 (N_8391,N_4727,N_5501);
or U8392 (N_8392,N_3701,N_4880);
nand U8393 (N_8393,N_3167,N_3388);
nand U8394 (N_8394,N_4460,N_5603);
nor U8395 (N_8395,N_3156,N_4834);
or U8396 (N_8396,N_3605,N_3404);
and U8397 (N_8397,N_5675,N_4486);
and U8398 (N_8398,N_5455,N_3764);
nand U8399 (N_8399,N_3189,N_3017);
and U8400 (N_8400,N_4951,N_4763);
xnor U8401 (N_8401,N_3569,N_4834);
nor U8402 (N_8402,N_4216,N_4141);
nor U8403 (N_8403,N_3124,N_3543);
or U8404 (N_8404,N_4762,N_5478);
nand U8405 (N_8405,N_4973,N_5460);
or U8406 (N_8406,N_5690,N_4970);
and U8407 (N_8407,N_5981,N_3744);
or U8408 (N_8408,N_3502,N_3321);
nand U8409 (N_8409,N_4434,N_4739);
nor U8410 (N_8410,N_5089,N_5401);
nor U8411 (N_8411,N_4564,N_5512);
or U8412 (N_8412,N_4447,N_5464);
xnor U8413 (N_8413,N_4491,N_5953);
nand U8414 (N_8414,N_3009,N_4768);
or U8415 (N_8415,N_4530,N_4795);
and U8416 (N_8416,N_4990,N_3496);
nor U8417 (N_8417,N_3242,N_4148);
or U8418 (N_8418,N_5451,N_5230);
or U8419 (N_8419,N_4134,N_5456);
xnor U8420 (N_8420,N_3672,N_4087);
xor U8421 (N_8421,N_5529,N_5973);
or U8422 (N_8422,N_3475,N_5649);
or U8423 (N_8423,N_5480,N_4866);
and U8424 (N_8424,N_5937,N_3502);
or U8425 (N_8425,N_4688,N_5067);
nor U8426 (N_8426,N_4275,N_3774);
and U8427 (N_8427,N_3202,N_3588);
nor U8428 (N_8428,N_3386,N_3875);
nor U8429 (N_8429,N_3585,N_5609);
nor U8430 (N_8430,N_3899,N_3630);
and U8431 (N_8431,N_4317,N_3069);
nand U8432 (N_8432,N_4418,N_5453);
xnor U8433 (N_8433,N_4839,N_3400);
xnor U8434 (N_8434,N_3130,N_4340);
nor U8435 (N_8435,N_5720,N_4487);
nand U8436 (N_8436,N_3407,N_5693);
nor U8437 (N_8437,N_4849,N_3990);
or U8438 (N_8438,N_5552,N_4648);
nor U8439 (N_8439,N_3230,N_3468);
nor U8440 (N_8440,N_5594,N_4259);
and U8441 (N_8441,N_3196,N_4675);
xor U8442 (N_8442,N_3943,N_5892);
nor U8443 (N_8443,N_4592,N_4890);
or U8444 (N_8444,N_5133,N_4448);
xnor U8445 (N_8445,N_3715,N_4764);
nor U8446 (N_8446,N_5918,N_4467);
and U8447 (N_8447,N_4255,N_4887);
nand U8448 (N_8448,N_3788,N_5139);
nor U8449 (N_8449,N_5031,N_5710);
nor U8450 (N_8450,N_4915,N_3647);
xnor U8451 (N_8451,N_5849,N_3787);
nor U8452 (N_8452,N_3528,N_3690);
or U8453 (N_8453,N_5517,N_3861);
nand U8454 (N_8454,N_5946,N_4997);
nor U8455 (N_8455,N_4169,N_5003);
xnor U8456 (N_8456,N_4730,N_5556);
or U8457 (N_8457,N_3067,N_5259);
and U8458 (N_8458,N_5045,N_5987);
and U8459 (N_8459,N_5011,N_3065);
nand U8460 (N_8460,N_4229,N_4855);
nand U8461 (N_8461,N_3507,N_4689);
nor U8462 (N_8462,N_5884,N_4075);
or U8463 (N_8463,N_3408,N_4169);
nand U8464 (N_8464,N_5156,N_4695);
or U8465 (N_8465,N_3934,N_4195);
nand U8466 (N_8466,N_5550,N_3263);
and U8467 (N_8467,N_4198,N_5162);
or U8468 (N_8468,N_3537,N_5412);
nand U8469 (N_8469,N_4302,N_5155);
nand U8470 (N_8470,N_4802,N_5762);
nor U8471 (N_8471,N_5607,N_3483);
nand U8472 (N_8472,N_5342,N_5021);
and U8473 (N_8473,N_3427,N_3001);
and U8474 (N_8474,N_4464,N_5760);
nor U8475 (N_8475,N_4913,N_4633);
nand U8476 (N_8476,N_4286,N_5056);
and U8477 (N_8477,N_3504,N_5630);
or U8478 (N_8478,N_5700,N_3794);
nand U8479 (N_8479,N_5453,N_4805);
or U8480 (N_8480,N_3826,N_4643);
or U8481 (N_8481,N_3855,N_3379);
and U8482 (N_8482,N_5689,N_3316);
xnor U8483 (N_8483,N_5377,N_3058);
and U8484 (N_8484,N_4561,N_4190);
xnor U8485 (N_8485,N_3126,N_5764);
nand U8486 (N_8486,N_5935,N_4786);
and U8487 (N_8487,N_3853,N_5514);
nand U8488 (N_8488,N_4751,N_5607);
and U8489 (N_8489,N_3913,N_5902);
nand U8490 (N_8490,N_5339,N_5438);
or U8491 (N_8491,N_5180,N_5838);
nor U8492 (N_8492,N_4066,N_5201);
or U8493 (N_8493,N_5213,N_3803);
nand U8494 (N_8494,N_5665,N_4785);
nor U8495 (N_8495,N_4889,N_5864);
and U8496 (N_8496,N_5023,N_3681);
nand U8497 (N_8497,N_5437,N_5753);
and U8498 (N_8498,N_3837,N_4182);
or U8499 (N_8499,N_3763,N_4413);
nor U8500 (N_8500,N_3757,N_4221);
or U8501 (N_8501,N_4563,N_5721);
nand U8502 (N_8502,N_3613,N_4097);
xor U8503 (N_8503,N_3589,N_4537);
nand U8504 (N_8504,N_5468,N_5000);
nor U8505 (N_8505,N_3006,N_4635);
xor U8506 (N_8506,N_5569,N_5805);
nor U8507 (N_8507,N_4025,N_3534);
nor U8508 (N_8508,N_4033,N_5662);
nor U8509 (N_8509,N_4039,N_5186);
nor U8510 (N_8510,N_4086,N_4935);
nand U8511 (N_8511,N_3752,N_5956);
or U8512 (N_8512,N_5770,N_5893);
nor U8513 (N_8513,N_3619,N_4157);
and U8514 (N_8514,N_3915,N_4488);
nor U8515 (N_8515,N_5658,N_3090);
and U8516 (N_8516,N_4344,N_4602);
or U8517 (N_8517,N_3676,N_3129);
or U8518 (N_8518,N_3079,N_3457);
and U8519 (N_8519,N_3599,N_4586);
xnor U8520 (N_8520,N_5808,N_4034);
nor U8521 (N_8521,N_5083,N_4877);
xnor U8522 (N_8522,N_3034,N_3097);
nand U8523 (N_8523,N_5222,N_5397);
or U8524 (N_8524,N_3411,N_3530);
or U8525 (N_8525,N_3249,N_4229);
and U8526 (N_8526,N_5131,N_4074);
nand U8527 (N_8527,N_3974,N_5233);
or U8528 (N_8528,N_3506,N_3708);
and U8529 (N_8529,N_4389,N_3329);
nand U8530 (N_8530,N_4597,N_4838);
nor U8531 (N_8531,N_5821,N_3076);
nand U8532 (N_8532,N_3391,N_3111);
nand U8533 (N_8533,N_5148,N_5102);
and U8534 (N_8534,N_3939,N_5305);
nor U8535 (N_8535,N_3848,N_5734);
xor U8536 (N_8536,N_3363,N_5643);
and U8537 (N_8537,N_4780,N_5177);
or U8538 (N_8538,N_3254,N_4141);
nand U8539 (N_8539,N_3954,N_5159);
xor U8540 (N_8540,N_5296,N_5365);
and U8541 (N_8541,N_5931,N_3129);
or U8542 (N_8542,N_3606,N_3116);
and U8543 (N_8543,N_5946,N_4044);
nand U8544 (N_8544,N_4644,N_5194);
and U8545 (N_8545,N_4673,N_3182);
nand U8546 (N_8546,N_3961,N_5253);
nand U8547 (N_8547,N_4554,N_3743);
nor U8548 (N_8548,N_5573,N_3724);
nor U8549 (N_8549,N_3137,N_5504);
or U8550 (N_8550,N_4338,N_4265);
and U8551 (N_8551,N_3629,N_4983);
nor U8552 (N_8552,N_3088,N_5425);
nand U8553 (N_8553,N_3104,N_4171);
and U8554 (N_8554,N_4125,N_3147);
nand U8555 (N_8555,N_3297,N_4526);
or U8556 (N_8556,N_4032,N_3153);
xnor U8557 (N_8557,N_4890,N_4216);
nor U8558 (N_8558,N_5212,N_3923);
xnor U8559 (N_8559,N_5559,N_3724);
xor U8560 (N_8560,N_3616,N_5289);
nand U8561 (N_8561,N_4553,N_4209);
or U8562 (N_8562,N_4325,N_3000);
nor U8563 (N_8563,N_3722,N_3571);
and U8564 (N_8564,N_5805,N_5733);
and U8565 (N_8565,N_3486,N_3917);
nor U8566 (N_8566,N_5298,N_4137);
xnor U8567 (N_8567,N_4342,N_3724);
xor U8568 (N_8568,N_3192,N_5796);
nand U8569 (N_8569,N_4436,N_5939);
and U8570 (N_8570,N_5100,N_4724);
nand U8571 (N_8571,N_5101,N_4329);
nand U8572 (N_8572,N_5065,N_5002);
nor U8573 (N_8573,N_3581,N_3356);
or U8574 (N_8574,N_4686,N_5790);
nand U8575 (N_8575,N_3205,N_5895);
and U8576 (N_8576,N_4079,N_3459);
and U8577 (N_8577,N_3762,N_4814);
and U8578 (N_8578,N_3919,N_5900);
and U8579 (N_8579,N_5544,N_4313);
and U8580 (N_8580,N_3607,N_4291);
nand U8581 (N_8581,N_5562,N_5577);
or U8582 (N_8582,N_4233,N_3032);
xnor U8583 (N_8583,N_4984,N_5952);
or U8584 (N_8584,N_4861,N_3287);
or U8585 (N_8585,N_3391,N_4356);
nand U8586 (N_8586,N_3579,N_5395);
nand U8587 (N_8587,N_4303,N_5774);
xnor U8588 (N_8588,N_5931,N_4781);
or U8589 (N_8589,N_4174,N_4773);
or U8590 (N_8590,N_3639,N_4094);
and U8591 (N_8591,N_5338,N_4822);
nand U8592 (N_8592,N_5197,N_3390);
and U8593 (N_8593,N_4862,N_4983);
nand U8594 (N_8594,N_5720,N_4206);
or U8595 (N_8595,N_5089,N_3043);
and U8596 (N_8596,N_4688,N_5204);
xor U8597 (N_8597,N_5286,N_4691);
or U8598 (N_8598,N_4357,N_4441);
nand U8599 (N_8599,N_4114,N_3957);
xnor U8600 (N_8600,N_4789,N_3667);
nor U8601 (N_8601,N_4286,N_4665);
nand U8602 (N_8602,N_3601,N_4638);
and U8603 (N_8603,N_5246,N_5994);
or U8604 (N_8604,N_4189,N_3944);
or U8605 (N_8605,N_5101,N_4985);
and U8606 (N_8606,N_3417,N_4072);
xnor U8607 (N_8607,N_3853,N_5059);
or U8608 (N_8608,N_3189,N_5572);
nor U8609 (N_8609,N_4246,N_3402);
nor U8610 (N_8610,N_5930,N_3531);
or U8611 (N_8611,N_5450,N_4629);
xnor U8612 (N_8612,N_4075,N_4683);
or U8613 (N_8613,N_4759,N_4660);
or U8614 (N_8614,N_4527,N_5362);
nor U8615 (N_8615,N_5413,N_5924);
or U8616 (N_8616,N_3282,N_4323);
nand U8617 (N_8617,N_3498,N_5621);
or U8618 (N_8618,N_5736,N_5249);
nor U8619 (N_8619,N_3215,N_4470);
nand U8620 (N_8620,N_5687,N_5668);
nand U8621 (N_8621,N_3150,N_4876);
nor U8622 (N_8622,N_3181,N_4574);
nand U8623 (N_8623,N_3624,N_5441);
and U8624 (N_8624,N_5298,N_3657);
nor U8625 (N_8625,N_4089,N_4469);
xnor U8626 (N_8626,N_4650,N_5934);
and U8627 (N_8627,N_4954,N_5157);
and U8628 (N_8628,N_4641,N_3784);
or U8629 (N_8629,N_3037,N_5856);
xnor U8630 (N_8630,N_3400,N_3623);
and U8631 (N_8631,N_3740,N_4474);
or U8632 (N_8632,N_3097,N_5891);
nor U8633 (N_8633,N_5738,N_4370);
or U8634 (N_8634,N_4343,N_3816);
or U8635 (N_8635,N_3128,N_5721);
nor U8636 (N_8636,N_4754,N_3454);
nand U8637 (N_8637,N_5963,N_4853);
nand U8638 (N_8638,N_4533,N_5214);
or U8639 (N_8639,N_3697,N_4252);
or U8640 (N_8640,N_4816,N_3787);
or U8641 (N_8641,N_5941,N_5357);
nor U8642 (N_8642,N_3463,N_3962);
nor U8643 (N_8643,N_5021,N_5205);
nand U8644 (N_8644,N_4397,N_5706);
nand U8645 (N_8645,N_4310,N_5003);
and U8646 (N_8646,N_5259,N_4644);
nor U8647 (N_8647,N_5777,N_4533);
and U8648 (N_8648,N_5935,N_3041);
or U8649 (N_8649,N_3942,N_3109);
nor U8650 (N_8650,N_4501,N_3069);
nor U8651 (N_8651,N_5300,N_5500);
nor U8652 (N_8652,N_4154,N_5947);
nor U8653 (N_8653,N_3397,N_4462);
and U8654 (N_8654,N_3430,N_3784);
xnor U8655 (N_8655,N_3461,N_4219);
or U8656 (N_8656,N_3580,N_4444);
or U8657 (N_8657,N_4577,N_4674);
or U8658 (N_8658,N_5634,N_4738);
nor U8659 (N_8659,N_3277,N_3839);
nor U8660 (N_8660,N_3107,N_5315);
nand U8661 (N_8661,N_5484,N_4921);
or U8662 (N_8662,N_4932,N_4790);
or U8663 (N_8663,N_4921,N_3233);
xor U8664 (N_8664,N_5398,N_4870);
nand U8665 (N_8665,N_3302,N_3481);
nor U8666 (N_8666,N_3755,N_5280);
or U8667 (N_8667,N_4986,N_4709);
nand U8668 (N_8668,N_4800,N_4097);
nand U8669 (N_8669,N_4010,N_5264);
and U8670 (N_8670,N_5784,N_4999);
xor U8671 (N_8671,N_5088,N_3353);
or U8672 (N_8672,N_5526,N_5205);
xnor U8673 (N_8673,N_3617,N_5991);
nand U8674 (N_8674,N_5207,N_5096);
nor U8675 (N_8675,N_3368,N_5987);
nand U8676 (N_8676,N_5726,N_5043);
nand U8677 (N_8677,N_5267,N_5861);
xor U8678 (N_8678,N_4386,N_3456);
nand U8679 (N_8679,N_3927,N_3992);
nand U8680 (N_8680,N_3395,N_5831);
and U8681 (N_8681,N_3091,N_3607);
and U8682 (N_8682,N_5663,N_4960);
and U8683 (N_8683,N_3759,N_4305);
nor U8684 (N_8684,N_5760,N_4536);
nand U8685 (N_8685,N_5345,N_3191);
or U8686 (N_8686,N_4633,N_5442);
nor U8687 (N_8687,N_4750,N_4009);
or U8688 (N_8688,N_5535,N_3421);
or U8689 (N_8689,N_4426,N_5669);
and U8690 (N_8690,N_4471,N_4213);
or U8691 (N_8691,N_5026,N_3785);
and U8692 (N_8692,N_3050,N_4342);
and U8693 (N_8693,N_5795,N_4960);
or U8694 (N_8694,N_4986,N_3365);
or U8695 (N_8695,N_4986,N_3938);
or U8696 (N_8696,N_5506,N_3614);
nor U8697 (N_8697,N_3553,N_3564);
and U8698 (N_8698,N_4792,N_4803);
nor U8699 (N_8699,N_3210,N_3169);
nor U8700 (N_8700,N_5124,N_4882);
nand U8701 (N_8701,N_4103,N_3553);
nor U8702 (N_8702,N_5893,N_4642);
and U8703 (N_8703,N_3582,N_3109);
xor U8704 (N_8704,N_5971,N_5214);
or U8705 (N_8705,N_3880,N_5090);
and U8706 (N_8706,N_5669,N_5414);
and U8707 (N_8707,N_3490,N_5911);
and U8708 (N_8708,N_5183,N_3191);
and U8709 (N_8709,N_3390,N_5287);
or U8710 (N_8710,N_3826,N_5927);
or U8711 (N_8711,N_5280,N_4858);
and U8712 (N_8712,N_5134,N_5450);
nor U8713 (N_8713,N_4221,N_4855);
nor U8714 (N_8714,N_5813,N_3746);
xor U8715 (N_8715,N_4533,N_3757);
and U8716 (N_8716,N_4644,N_4986);
nand U8717 (N_8717,N_3715,N_4540);
nor U8718 (N_8718,N_4185,N_3216);
or U8719 (N_8719,N_5134,N_3246);
and U8720 (N_8720,N_4006,N_5447);
xnor U8721 (N_8721,N_5023,N_5208);
nor U8722 (N_8722,N_4592,N_5015);
nand U8723 (N_8723,N_3970,N_3348);
and U8724 (N_8724,N_4195,N_3031);
nand U8725 (N_8725,N_4768,N_3573);
nor U8726 (N_8726,N_4085,N_4805);
or U8727 (N_8727,N_3842,N_4055);
and U8728 (N_8728,N_3961,N_3314);
nor U8729 (N_8729,N_4444,N_4337);
or U8730 (N_8730,N_3872,N_5616);
nor U8731 (N_8731,N_3907,N_4483);
xnor U8732 (N_8732,N_5384,N_4384);
and U8733 (N_8733,N_3182,N_3528);
nor U8734 (N_8734,N_4634,N_3061);
and U8735 (N_8735,N_3419,N_5152);
or U8736 (N_8736,N_3875,N_5517);
or U8737 (N_8737,N_4845,N_3351);
nand U8738 (N_8738,N_4200,N_3343);
and U8739 (N_8739,N_4286,N_4545);
or U8740 (N_8740,N_4655,N_4187);
nand U8741 (N_8741,N_3908,N_4128);
nor U8742 (N_8742,N_5646,N_5709);
nand U8743 (N_8743,N_4702,N_5504);
or U8744 (N_8744,N_3804,N_5119);
and U8745 (N_8745,N_5212,N_5469);
and U8746 (N_8746,N_4441,N_5287);
or U8747 (N_8747,N_5521,N_5186);
xor U8748 (N_8748,N_3518,N_3708);
nand U8749 (N_8749,N_3747,N_5485);
and U8750 (N_8750,N_4447,N_4744);
xnor U8751 (N_8751,N_3037,N_3140);
or U8752 (N_8752,N_3195,N_5869);
and U8753 (N_8753,N_4532,N_5722);
nor U8754 (N_8754,N_5179,N_3061);
and U8755 (N_8755,N_3104,N_5606);
or U8756 (N_8756,N_5672,N_4793);
nor U8757 (N_8757,N_3652,N_4748);
nand U8758 (N_8758,N_4020,N_4262);
or U8759 (N_8759,N_3437,N_3266);
nand U8760 (N_8760,N_4239,N_5623);
xnor U8761 (N_8761,N_5878,N_5936);
nand U8762 (N_8762,N_5442,N_4765);
nand U8763 (N_8763,N_5924,N_4869);
nand U8764 (N_8764,N_5815,N_4156);
or U8765 (N_8765,N_5341,N_3587);
or U8766 (N_8766,N_3246,N_3620);
nor U8767 (N_8767,N_5075,N_5938);
and U8768 (N_8768,N_5655,N_3439);
nand U8769 (N_8769,N_5396,N_4785);
nor U8770 (N_8770,N_4555,N_4775);
or U8771 (N_8771,N_5709,N_4878);
and U8772 (N_8772,N_4789,N_4367);
nor U8773 (N_8773,N_3218,N_5544);
and U8774 (N_8774,N_3225,N_4042);
and U8775 (N_8775,N_4111,N_4511);
nor U8776 (N_8776,N_3755,N_3561);
or U8777 (N_8777,N_3007,N_5813);
and U8778 (N_8778,N_5707,N_3637);
nand U8779 (N_8779,N_5335,N_3858);
nor U8780 (N_8780,N_3577,N_4716);
or U8781 (N_8781,N_3582,N_5843);
or U8782 (N_8782,N_3881,N_5218);
nand U8783 (N_8783,N_4129,N_4771);
and U8784 (N_8784,N_3904,N_5332);
nor U8785 (N_8785,N_4796,N_4180);
nand U8786 (N_8786,N_5533,N_4622);
xnor U8787 (N_8787,N_5767,N_4997);
or U8788 (N_8788,N_4633,N_3689);
and U8789 (N_8789,N_4943,N_3759);
and U8790 (N_8790,N_3500,N_5835);
nor U8791 (N_8791,N_3704,N_5028);
xnor U8792 (N_8792,N_5269,N_3964);
and U8793 (N_8793,N_3694,N_3414);
or U8794 (N_8794,N_5237,N_5401);
nand U8795 (N_8795,N_3579,N_4857);
and U8796 (N_8796,N_5260,N_4416);
nor U8797 (N_8797,N_4347,N_3062);
nor U8798 (N_8798,N_3897,N_4866);
nand U8799 (N_8799,N_5949,N_4341);
nor U8800 (N_8800,N_5540,N_3231);
nor U8801 (N_8801,N_4856,N_4337);
nor U8802 (N_8802,N_4328,N_4420);
xor U8803 (N_8803,N_5116,N_3515);
or U8804 (N_8804,N_4773,N_5284);
and U8805 (N_8805,N_3163,N_5565);
nor U8806 (N_8806,N_5825,N_4966);
nand U8807 (N_8807,N_3768,N_5567);
nand U8808 (N_8808,N_4041,N_5098);
xnor U8809 (N_8809,N_3176,N_5390);
nor U8810 (N_8810,N_5452,N_4540);
and U8811 (N_8811,N_4357,N_3373);
nor U8812 (N_8812,N_4776,N_4155);
and U8813 (N_8813,N_3779,N_5823);
nand U8814 (N_8814,N_4435,N_4564);
nor U8815 (N_8815,N_5384,N_5140);
or U8816 (N_8816,N_5544,N_4033);
nor U8817 (N_8817,N_3127,N_3109);
or U8818 (N_8818,N_3919,N_3094);
xor U8819 (N_8819,N_3859,N_3162);
or U8820 (N_8820,N_3416,N_4361);
nor U8821 (N_8821,N_4992,N_4742);
and U8822 (N_8822,N_4516,N_4430);
nor U8823 (N_8823,N_3292,N_4512);
xnor U8824 (N_8824,N_4949,N_4057);
nand U8825 (N_8825,N_3592,N_4961);
or U8826 (N_8826,N_3761,N_3604);
nand U8827 (N_8827,N_5240,N_3268);
nor U8828 (N_8828,N_5404,N_5012);
xnor U8829 (N_8829,N_3627,N_3634);
nand U8830 (N_8830,N_5064,N_4724);
or U8831 (N_8831,N_3051,N_5356);
xor U8832 (N_8832,N_5014,N_4242);
or U8833 (N_8833,N_3812,N_5857);
nor U8834 (N_8834,N_5241,N_4685);
and U8835 (N_8835,N_4259,N_4731);
and U8836 (N_8836,N_5881,N_4853);
xnor U8837 (N_8837,N_3351,N_3254);
and U8838 (N_8838,N_5877,N_4521);
nand U8839 (N_8839,N_5133,N_5068);
nor U8840 (N_8840,N_3196,N_3473);
nor U8841 (N_8841,N_4117,N_4824);
nand U8842 (N_8842,N_5421,N_4104);
or U8843 (N_8843,N_5193,N_4508);
nand U8844 (N_8844,N_3759,N_5558);
and U8845 (N_8845,N_4266,N_3205);
or U8846 (N_8846,N_3882,N_3017);
nor U8847 (N_8847,N_3628,N_5939);
and U8848 (N_8848,N_4133,N_4922);
xnor U8849 (N_8849,N_4149,N_4752);
or U8850 (N_8850,N_5370,N_4990);
nand U8851 (N_8851,N_4218,N_4875);
nor U8852 (N_8852,N_3548,N_5211);
nor U8853 (N_8853,N_3828,N_3946);
and U8854 (N_8854,N_5813,N_4232);
or U8855 (N_8855,N_3628,N_3996);
or U8856 (N_8856,N_3824,N_3043);
nand U8857 (N_8857,N_3108,N_4214);
nor U8858 (N_8858,N_4780,N_3616);
or U8859 (N_8859,N_5998,N_4449);
or U8860 (N_8860,N_4667,N_3721);
and U8861 (N_8861,N_3762,N_3113);
nor U8862 (N_8862,N_5761,N_5232);
nor U8863 (N_8863,N_4833,N_3691);
nor U8864 (N_8864,N_5007,N_5198);
and U8865 (N_8865,N_3390,N_4448);
or U8866 (N_8866,N_4604,N_5350);
and U8867 (N_8867,N_4732,N_5435);
and U8868 (N_8868,N_4502,N_4594);
nand U8869 (N_8869,N_4077,N_3061);
xnor U8870 (N_8870,N_4551,N_3926);
and U8871 (N_8871,N_5019,N_5785);
nor U8872 (N_8872,N_5475,N_5138);
nand U8873 (N_8873,N_5675,N_3775);
xor U8874 (N_8874,N_4067,N_3657);
nand U8875 (N_8875,N_3816,N_4489);
or U8876 (N_8876,N_4406,N_3474);
xnor U8877 (N_8877,N_5454,N_4452);
nand U8878 (N_8878,N_3090,N_5495);
nand U8879 (N_8879,N_4497,N_5804);
or U8880 (N_8880,N_5527,N_3700);
or U8881 (N_8881,N_3321,N_5227);
nor U8882 (N_8882,N_3195,N_4842);
nor U8883 (N_8883,N_5602,N_4728);
nor U8884 (N_8884,N_4432,N_3001);
and U8885 (N_8885,N_5158,N_5467);
and U8886 (N_8886,N_5196,N_5361);
nand U8887 (N_8887,N_5799,N_5526);
and U8888 (N_8888,N_4072,N_5316);
nand U8889 (N_8889,N_3432,N_5207);
nor U8890 (N_8890,N_4307,N_5351);
or U8891 (N_8891,N_4100,N_3168);
and U8892 (N_8892,N_5901,N_4341);
nand U8893 (N_8893,N_5509,N_5270);
or U8894 (N_8894,N_4018,N_3571);
nand U8895 (N_8895,N_5689,N_3795);
and U8896 (N_8896,N_4768,N_4703);
xor U8897 (N_8897,N_5882,N_4782);
xnor U8898 (N_8898,N_5491,N_4934);
nand U8899 (N_8899,N_5960,N_4887);
and U8900 (N_8900,N_3834,N_3894);
nor U8901 (N_8901,N_4823,N_5843);
nor U8902 (N_8902,N_3644,N_3704);
nand U8903 (N_8903,N_5895,N_4449);
nor U8904 (N_8904,N_4357,N_3847);
nor U8905 (N_8905,N_3776,N_3246);
xor U8906 (N_8906,N_5078,N_5220);
xnor U8907 (N_8907,N_3155,N_3584);
or U8908 (N_8908,N_5845,N_3052);
xnor U8909 (N_8909,N_3255,N_4845);
nor U8910 (N_8910,N_4198,N_4568);
and U8911 (N_8911,N_4316,N_5482);
nor U8912 (N_8912,N_5641,N_5837);
and U8913 (N_8913,N_4523,N_3339);
or U8914 (N_8914,N_3179,N_5934);
and U8915 (N_8915,N_3097,N_4592);
and U8916 (N_8916,N_4164,N_4852);
nor U8917 (N_8917,N_3664,N_5521);
nand U8918 (N_8918,N_5231,N_5840);
nand U8919 (N_8919,N_4715,N_5506);
nand U8920 (N_8920,N_5522,N_4382);
nor U8921 (N_8921,N_5748,N_4285);
xnor U8922 (N_8922,N_3863,N_5138);
and U8923 (N_8923,N_5129,N_4426);
xor U8924 (N_8924,N_4404,N_3109);
and U8925 (N_8925,N_3142,N_5081);
nand U8926 (N_8926,N_4885,N_5586);
or U8927 (N_8927,N_3553,N_4270);
xnor U8928 (N_8928,N_4659,N_4101);
nor U8929 (N_8929,N_3381,N_3909);
or U8930 (N_8930,N_3153,N_3206);
xnor U8931 (N_8931,N_5550,N_4430);
and U8932 (N_8932,N_5101,N_5976);
or U8933 (N_8933,N_5371,N_5807);
nor U8934 (N_8934,N_3971,N_3179);
nand U8935 (N_8935,N_3980,N_5910);
nor U8936 (N_8936,N_4169,N_5694);
xor U8937 (N_8937,N_3145,N_3048);
nand U8938 (N_8938,N_5058,N_5042);
xnor U8939 (N_8939,N_5104,N_5842);
nand U8940 (N_8940,N_4934,N_4047);
and U8941 (N_8941,N_5422,N_5659);
nand U8942 (N_8942,N_5978,N_4509);
and U8943 (N_8943,N_5909,N_5009);
and U8944 (N_8944,N_5432,N_3767);
nor U8945 (N_8945,N_5367,N_4560);
and U8946 (N_8946,N_3273,N_3530);
and U8947 (N_8947,N_5563,N_4478);
nand U8948 (N_8948,N_3023,N_3000);
or U8949 (N_8949,N_5999,N_4187);
xnor U8950 (N_8950,N_5373,N_3701);
and U8951 (N_8951,N_5704,N_3739);
xnor U8952 (N_8952,N_4147,N_3502);
nand U8953 (N_8953,N_3036,N_3339);
xor U8954 (N_8954,N_4976,N_4369);
nand U8955 (N_8955,N_4521,N_4726);
or U8956 (N_8956,N_5461,N_5878);
nand U8957 (N_8957,N_3999,N_4693);
or U8958 (N_8958,N_4279,N_5637);
nand U8959 (N_8959,N_3247,N_4038);
nor U8960 (N_8960,N_5903,N_4596);
and U8961 (N_8961,N_5136,N_3035);
nor U8962 (N_8962,N_5057,N_3257);
or U8963 (N_8963,N_3952,N_5420);
xnor U8964 (N_8964,N_5707,N_3193);
and U8965 (N_8965,N_3051,N_4428);
and U8966 (N_8966,N_4589,N_3382);
and U8967 (N_8967,N_3025,N_4758);
nor U8968 (N_8968,N_5905,N_5359);
and U8969 (N_8969,N_5563,N_4918);
nand U8970 (N_8970,N_3166,N_5213);
or U8971 (N_8971,N_5951,N_4616);
nand U8972 (N_8972,N_4465,N_3437);
nand U8973 (N_8973,N_4903,N_4886);
nor U8974 (N_8974,N_5673,N_3216);
nand U8975 (N_8975,N_4758,N_4514);
nor U8976 (N_8976,N_3869,N_4296);
xnor U8977 (N_8977,N_4075,N_4216);
nand U8978 (N_8978,N_5947,N_4292);
or U8979 (N_8979,N_3983,N_5664);
and U8980 (N_8980,N_3346,N_4302);
or U8981 (N_8981,N_3837,N_3371);
or U8982 (N_8982,N_3539,N_5308);
or U8983 (N_8983,N_5475,N_4215);
and U8984 (N_8984,N_4677,N_3514);
nand U8985 (N_8985,N_3988,N_5328);
nand U8986 (N_8986,N_4294,N_5887);
and U8987 (N_8987,N_4131,N_4972);
or U8988 (N_8988,N_3579,N_3668);
nor U8989 (N_8989,N_3095,N_5982);
and U8990 (N_8990,N_3529,N_5268);
xor U8991 (N_8991,N_3396,N_5011);
and U8992 (N_8992,N_5437,N_5936);
nand U8993 (N_8993,N_3129,N_3789);
or U8994 (N_8994,N_5375,N_5133);
nor U8995 (N_8995,N_3579,N_5635);
nand U8996 (N_8996,N_4366,N_5281);
nor U8997 (N_8997,N_4542,N_5985);
or U8998 (N_8998,N_3333,N_3301);
xor U8999 (N_8999,N_5254,N_5212);
and U9000 (N_9000,N_6160,N_8772);
nand U9001 (N_9001,N_7050,N_7797);
or U9002 (N_9002,N_7568,N_7625);
nor U9003 (N_9003,N_7972,N_7722);
nand U9004 (N_9004,N_6055,N_6524);
nand U9005 (N_9005,N_7369,N_8504);
and U9006 (N_9006,N_8102,N_6768);
and U9007 (N_9007,N_8325,N_8139);
nor U9008 (N_9008,N_8180,N_7839);
or U9009 (N_9009,N_6361,N_6909);
or U9010 (N_9010,N_6156,N_7206);
nand U9011 (N_9011,N_8917,N_7899);
or U9012 (N_9012,N_8719,N_8488);
and U9013 (N_9013,N_7274,N_8999);
nor U9014 (N_9014,N_8873,N_8882);
and U9015 (N_9015,N_8644,N_8057);
and U9016 (N_9016,N_7575,N_8854);
xnor U9017 (N_9017,N_8577,N_7278);
nand U9018 (N_9018,N_7370,N_8932);
nor U9019 (N_9019,N_7407,N_6362);
and U9020 (N_9020,N_8731,N_7216);
nor U9021 (N_9021,N_8828,N_7923);
xor U9022 (N_9022,N_6318,N_7467);
xnor U9023 (N_9023,N_6371,N_6283);
nand U9024 (N_9024,N_8331,N_6015);
and U9025 (N_9025,N_6612,N_7900);
nor U9026 (N_9026,N_8847,N_7310);
nand U9027 (N_9027,N_8483,N_8538);
and U9028 (N_9028,N_7306,N_6672);
or U9029 (N_9029,N_6916,N_7685);
or U9030 (N_9030,N_6086,N_8654);
nor U9031 (N_9031,N_7411,N_7836);
or U9032 (N_9032,N_6713,N_6546);
xnor U9033 (N_9033,N_7189,N_6796);
nor U9034 (N_9034,N_6609,N_6323);
or U9035 (N_9035,N_7191,N_8991);
nand U9036 (N_9036,N_7237,N_6252);
or U9037 (N_9037,N_6985,N_7680);
nor U9038 (N_9038,N_8142,N_6516);
and U9039 (N_9039,N_8175,N_7466);
and U9040 (N_9040,N_6913,N_6358);
or U9041 (N_9041,N_6892,N_7672);
and U9042 (N_9042,N_7412,N_7666);
and U9043 (N_9043,N_6510,N_8894);
nor U9044 (N_9044,N_8702,N_8899);
xor U9045 (N_9045,N_8652,N_7400);
and U9046 (N_9046,N_6726,N_6474);
nor U9047 (N_9047,N_7249,N_7589);
nor U9048 (N_9048,N_6421,N_6057);
nand U9049 (N_9049,N_6821,N_8086);
and U9050 (N_9050,N_7626,N_7435);
nand U9051 (N_9051,N_8145,N_8388);
nor U9052 (N_9052,N_6236,N_8759);
or U9053 (N_9053,N_6306,N_6836);
nand U9054 (N_9054,N_8448,N_7176);
nor U9055 (N_9055,N_7288,N_7069);
nand U9056 (N_9056,N_7955,N_6861);
and U9057 (N_9057,N_7503,N_7173);
xnor U9058 (N_9058,N_8919,N_8144);
or U9059 (N_9059,N_8682,N_8558);
nor U9060 (N_9060,N_8512,N_6042);
nand U9061 (N_9061,N_7147,N_6158);
and U9062 (N_9062,N_6813,N_8259);
and U9063 (N_9063,N_7422,N_8440);
xnor U9064 (N_9064,N_8713,N_6235);
nor U9065 (N_9065,N_7227,N_8510);
or U9066 (N_9066,N_8327,N_8027);
or U9067 (N_9067,N_8303,N_6711);
and U9068 (N_9068,N_6037,N_6248);
and U9069 (N_9069,N_7989,N_7280);
xor U9070 (N_9070,N_7507,N_8755);
nor U9071 (N_9071,N_7064,N_7226);
nor U9072 (N_9072,N_8569,N_7220);
nand U9073 (N_9073,N_6506,N_8306);
and U9074 (N_9074,N_6325,N_8422);
or U9075 (N_9075,N_6418,N_7408);
xnor U9076 (N_9076,N_6354,N_8414);
nor U9077 (N_9077,N_7322,N_7809);
nor U9078 (N_9078,N_8640,N_7596);
or U9079 (N_9079,N_6563,N_6071);
and U9080 (N_9080,N_8585,N_6584);
nand U9081 (N_9081,N_6380,N_8870);
nand U9082 (N_9082,N_8760,N_7070);
xnor U9083 (N_9083,N_7477,N_8253);
nor U9084 (N_9084,N_7590,N_8628);
or U9085 (N_9085,N_6171,N_8801);
nand U9086 (N_9086,N_8466,N_8354);
nand U9087 (N_9087,N_6435,N_8505);
and U9088 (N_9088,N_7952,N_6538);
or U9089 (N_9089,N_7663,N_6389);
or U9090 (N_9090,N_6949,N_7832);
nand U9091 (N_9091,N_7451,N_8594);
nand U9092 (N_9092,N_6844,N_8220);
nand U9093 (N_9093,N_6787,N_6062);
and U9094 (N_9094,N_6113,N_8468);
nor U9095 (N_9095,N_6603,N_8231);
xor U9096 (N_9096,N_8951,N_7442);
or U9097 (N_9097,N_7617,N_8093);
or U9098 (N_9098,N_6050,N_7326);
nor U9099 (N_9099,N_6995,N_6274);
or U9100 (N_9100,N_7366,N_8288);
or U9101 (N_9101,N_7481,N_8452);
xor U9102 (N_9102,N_7582,N_7183);
and U9103 (N_9103,N_7533,N_7072);
nand U9104 (N_9104,N_7787,N_8861);
or U9105 (N_9105,N_8007,N_7434);
and U9106 (N_9106,N_8823,N_6479);
and U9107 (N_9107,N_6356,N_8211);
nand U9108 (N_9108,N_8243,N_7891);
nor U9109 (N_9109,N_6219,N_7356);
or U9110 (N_9110,N_8202,N_6558);
xor U9111 (N_9111,N_7478,N_8263);
nand U9112 (N_9112,N_7460,N_7855);
nand U9113 (N_9113,N_6781,N_7750);
nor U9114 (N_9114,N_7986,N_8112);
nand U9115 (N_9115,N_7565,N_8345);
and U9116 (N_9116,N_6571,N_8790);
and U9117 (N_9117,N_6394,N_6937);
and U9118 (N_9118,N_8246,N_6905);
nand U9119 (N_9119,N_8580,N_8547);
nand U9120 (N_9120,N_6551,N_6674);
nor U9121 (N_9121,N_8517,N_6815);
nand U9122 (N_9122,N_6072,N_8081);
or U9123 (N_9123,N_8878,N_8537);
and U9124 (N_9124,N_7027,N_7002);
nand U9125 (N_9125,N_8542,N_7324);
or U9126 (N_9126,N_7962,N_8099);
nand U9127 (N_9127,N_6379,N_6972);
or U9128 (N_9128,N_7627,N_6760);
and U9129 (N_9129,N_6999,N_8565);
nor U9130 (N_9130,N_8972,N_8437);
nor U9131 (N_9131,N_7689,N_7656);
nor U9132 (N_9132,N_7530,N_6253);
and U9133 (N_9133,N_7806,N_8756);
nand U9134 (N_9134,N_8276,N_7420);
nand U9135 (N_9135,N_7062,N_6777);
and U9136 (N_9136,N_7464,N_8025);
nand U9137 (N_9137,N_6216,N_7242);
or U9138 (N_9138,N_8578,N_7188);
nor U9139 (N_9139,N_6877,N_7009);
and U9140 (N_9140,N_7522,N_6381);
and U9141 (N_9141,N_7441,N_8219);
and U9142 (N_9142,N_7840,N_8681);
or U9143 (N_9143,N_8834,N_8379);
or U9144 (N_9144,N_6695,N_7785);
or U9145 (N_9145,N_6540,N_6289);
nand U9146 (N_9146,N_6302,N_8582);
nand U9147 (N_9147,N_8796,N_6124);
or U9148 (N_9148,N_6297,N_6691);
nand U9149 (N_9149,N_7704,N_8725);
or U9150 (N_9150,N_8011,N_8970);
nor U9151 (N_9151,N_6148,N_7379);
nor U9152 (N_9152,N_7543,N_6973);
nand U9153 (N_9153,N_8778,N_6974);
nor U9154 (N_9154,N_7992,N_7592);
xnor U9155 (N_9155,N_6264,N_8138);
xnor U9156 (N_9156,N_7375,N_8430);
nor U9157 (N_9157,N_8741,N_7098);
and U9158 (N_9158,N_8927,N_6218);
nand U9159 (N_9159,N_8619,N_6876);
xnor U9160 (N_9160,N_6754,N_6854);
and U9161 (N_9161,N_7544,N_8450);
or U9162 (N_9162,N_8267,N_7246);
and U9163 (N_9163,N_6519,N_6491);
nor U9164 (N_9164,N_7710,N_6317);
and U9165 (N_9165,N_8529,N_7788);
xnor U9166 (N_9166,N_7929,N_7223);
xnor U9167 (N_9167,N_7706,N_6620);
or U9168 (N_9168,N_7395,N_6707);
nand U9169 (N_9169,N_6560,N_7194);
nor U9170 (N_9170,N_6133,N_8050);
and U9171 (N_9171,N_7684,N_7117);
xnor U9172 (N_9172,N_7723,N_6775);
xnor U9173 (N_9173,N_7184,N_6508);
nand U9174 (N_9174,N_8104,N_6220);
and U9175 (N_9175,N_7336,N_6975);
or U9176 (N_9176,N_7107,N_7372);
or U9177 (N_9177,N_7525,N_7059);
xor U9178 (N_9178,N_8680,N_6803);
nand U9179 (N_9179,N_7971,N_8995);
xnor U9180 (N_9180,N_7866,N_7462);
nor U9181 (N_9181,N_6522,N_8297);
nor U9182 (N_9182,N_7388,N_6445);
nor U9183 (N_9183,N_6893,N_7595);
and U9184 (N_9184,N_7028,N_8123);
or U9185 (N_9185,N_8645,N_8397);
and U9186 (N_9186,N_6463,N_8261);
nor U9187 (N_9187,N_6030,N_8234);
nor U9188 (N_9188,N_7837,N_6338);
nand U9189 (N_9189,N_8819,N_6756);
and U9190 (N_9190,N_6614,N_6805);
or U9191 (N_9191,N_7160,N_6322);
or U9192 (N_9192,N_6583,N_6799);
and U9193 (N_9193,N_8735,N_8302);
and U9194 (N_9194,N_6135,N_7045);
or U9195 (N_9195,N_7798,N_8914);
and U9196 (N_9196,N_8453,N_7550);
or U9197 (N_9197,N_7861,N_7032);
nand U9198 (N_9198,N_6376,N_7344);
nor U9199 (N_9199,N_6616,N_8903);
or U9200 (N_9200,N_7739,N_6428);
nor U9201 (N_9201,N_8475,N_6301);
and U9202 (N_9202,N_6458,N_8378);
and U9203 (N_9203,N_6308,N_6336);
or U9204 (N_9204,N_6555,N_6083);
or U9205 (N_9205,N_7000,N_7579);
or U9206 (N_9206,N_7919,N_6554);
nor U9207 (N_9207,N_6618,N_6542);
nand U9208 (N_9208,N_8833,N_8807);
nand U9209 (N_9209,N_7951,N_8674);
nand U9210 (N_9210,N_7129,N_8190);
or U9211 (N_9211,N_6065,N_8028);
xnor U9212 (N_9212,N_8496,N_8181);
nor U9213 (N_9213,N_6493,N_7413);
or U9214 (N_9214,N_7082,N_8309);
nand U9215 (N_9215,N_6820,N_8372);
and U9216 (N_9216,N_7588,N_8410);
nand U9217 (N_9217,N_7250,N_6259);
and U9218 (N_9218,N_6696,N_6517);
nand U9219 (N_9219,N_6058,N_7692);
or U9220 (N_9220,N_7964,N_8848);
nor U9221 (N_9221,N_8922,N_7882);
nand U9222 (N_9222,N_7865,N_7529);
nand U9223 (N_9223,N_7851,N_8767);
or U9224 (N_9224,N_8736,N_8387);
or U9225 (N_9225,N_7316,N_7283);
nand U9226 (N_9226,N_8831,N_8636);
nor U9227 (N_9227,N_8194,N_7734);
xnor U9228 (N_9228,N_6925,N_6249);
and U9229 (N_9229,N_7470,N_6214);
nor U9230 (N_9230,N_8940,N_6272);
nor U9231 (N_9231,N_7264,N_7038);
nand U9232 (N_9232,N_7586,N_8479);
and U9233 (N_9233,N_7204,N_7755);
nor U9234 (N_9234,N_7248,N_8635);
nand U9235 (N_9235,N_8366,N_7300);
and U9236 (N_9236,N_7404,N_6592);
nand U9237 (N_9237,N_6332,N_8618);
and U9238 (N_9238,N_6500,N_7872);
and U9239 (N_9239,N_8295,N_7262);
and U9240 (N_9240,N_8715,N_6675);
and U9241 (N_9241,N_7824,N_6211);
nor U9242 (N_9242,N_8408,N_6265);
nor U9243 (N_9243,N_6473,N_7368);
nor U9244 (N_9244,N_6221,N_6978);
or U9245 (N_9245,N_6879,N_7385);
nand U9246 (N_9246,N_7124,N_7635);
and U9247 (N_9247,N_8771,N_8507);
nand U9248 (N_9248,N_7528,N_6898);
or U9249 (N_9249,N_8324,N_8258);
or U9250 (N_9250,N_8762,N_8183);
nor U9251 (N_9251,N_8147,N_6848);
nor U9252 (N_9252,N_7217,N_6686);
nor U9253 (N_9253,N_6929,N_6596);
nor U9254 (N_9254,N_6926,N_8390);
nand U9255 (N_9255,N_8318,N_7505);
nor U9256 (N_9256,N_6009,N_7122);
nand U9257 (N_9257,N_6339,N_6823);
and U9258 (N_9258,N_8403,N_6683);
or U9259 (N_9259,N_6528,N_8374);
nor U9260 (N_9260,N_7558,N_7901);
nand U9261 (N_9261,N_6122,N_6650);
nand U9262 (N_9262,N_7396,N_6868);
or U9263 (N_9263,N_7658,N_6964);
and U9264 (N_9264,N_7431,N_7615);
nor U9265 (N_9265,N_8096,N_8359);
nor U9266 (N_9266,N_6484,N_8129);
nand U9267 (N_9267,N_8954,N_6134);
or U9268 (N_9268,N_8885,N_6128);
and U9269 (N_9269,N_8633,N_7591);
and U9270 (N_9270,N_6550,N_6780);
nand U9271 (N_9271,N_8737,N_6901);
nor U9272 (N_9272,N_6088,N_7023);
and U9273 (N_9273,N_8315,N_6087);
or U9274 (N_9274,N_6636,N_8843);
nand U9275 (N_9275,N_7611,N_6740);
nor U9276 (N_9276,N_8369,N_6600);
and U9277 (N_9277,N_6416,N_7709);
nand U9278 (N_9278,N_8552,N_7287);
nor U9279 (N_9279,N_8699,N_6988);
and U9280 (N_9280,N_7454,N_6941);
and U9281 (N_9281,N_6193,N_8776);
and U9282 (N_9282,N_8126,N_8791);
nand U9283 (N_9283,N_7687,N_6569);
and U9284 (N_9284,N_6657,N_8272);
and U9285 (N_9285,N_8988,N_7143);
nand U9286 (N_9286,N_6606,N_6127);
or U9287 (N_9287,N_6002,N_6315);
or U9288 (N_9288,N_6677,N_8581);
nand U9289 (N_9289,N_7125,N_6039);
or U9290 (N_9290,N_7931,N_8486);
and U9291 (N_9291,N_7337,N_7508);
nand U9292 (N_9292,N_6477,N_7608);
nor U9293 (N_9293,N_7162,N_8605);
and U9294 (N_9294,N_6783,N_7128);
nor U9295 (N_9295,N_7081,N_6933);
or U9296 (N_9296,N_6429,N_8458);
or U9297 (N_9297,N_8465,N_8852);
or U9298 (N_9298,N_6897,N_6722);
nor U9299 (N_9299,N_6702,N_8709);
or U9300 (N_9300,N_6690,N_8607);
or U9301 (N_9301,N_7948,N_8056);
or U9302 (N_9302,N_8394,N_8171);
or U9303 (N_9303,N_8376,N_7234);
nor U9304 (N_9304,N_8809,N_6367);
nor U9305 (N_9305,N_6172,N_6291);
and U9306 (N_9306,N_7051,N_6948);
and U9307 (N_9307,N_7736,N_7646);
nand U9308 (N_9308,N_6132,N_6281);
or U9309 (N_9309,N_8269,N_6968);
nand U9310 (N_9310,N_7294,N_6446);
nor U9311 (N_9311,N_6589,N_6655);
or U9312 (N_9312,N_6212,N_6883);
nor U9313 (N_9313,N_6635,N_6912);
nor U9314 (N_9314,N_6544,N_8199);
xor U9315 (N_9315,N_7593,N_6226);
and U9316 (N_9316,N_6142,N_7996);
and U9317 (N_9317,N_8985,N_6910);
and U9318 (N_9318,N_7893,N_7281);
and U9319 (N_9319,N_7569,N_7376);
nor U9320 (N_9320,N_6952,N_8881);
nand U9321 (N_9321,N_8395,N_6454);
nor U9322 (N_9322,N_6492,N_7202);
nand U9323 (N_9323,N_8184,N_7137);
xnor U9324 (N_9324,N_6859,N_8602);
nand U9325 (N_9325,N_8212,N_6424);
or U9326 (N_9326,N_8469,N_6449);
nor U9327 (N_9327,N_7843,N_6374);
or U9328 (N_9328,N_7796,N_7762);
nand U9329 (N_9329,N_7229,N_7105);
and U9330 (N_9330,N_7780,N_7940);
nor U9331 (N_9331,N_6241,N_8773);
and U9332 (N_9332,N_8810,N_8621);
nor U9333 (N_9333,N_7517,N_7917);
nand U9334 (N_9334,N_7152,N_7485);
nand U9335 (N_9335,N_8856,N_6460);
xnor U9336 (N_9336,N_8895,N_6478);
or U9337 (N_9337,N_8247,N_7988);
or U9338 (N_9338,N_6947,N_8751);
and U9339 (N_9339,N_8285,N_8103);
nand U9340 (N_9340,N_6224,N_8244);
nand U9341 (N_9341,N_6811,N_6673);
nor U9342 (N_9342,N_6772,N_7711);
nand U9343 (N_9343,N_8412,N_6628);
or U9344 (N_9344,N_8033,N_8849);
or U9345 (N_9345,N_6577,N_8067);
nor U9346 (N_9346,N_7885,N_7016);
nand U9347 (N_9347,N_8049,N_6881);
nor U9348 (N_9348,N_8035,N_8655);
nor U9349 (N_9349,N_6076,N_7610);
nor U9350 (N_9350,N_8941,N_8131);
nor U9351 (N_9351,N_7136,N_6044);
nand U9352 (N_9352,N_7773,N_7382);
or U9353 (N_9353,N_8548,N_7488);
nand U9354 (N_9354,N_8814,N_6716);
or U9355 (N_9355,N_7609,N_7506);
or U9356 (N_9356,N_8423,N_8158);
and U9357 (N_9357,N_8222,N_8508);
or U9358 (N_9358,N_7682,N_8764);
nor U9359 (N_9359,N_6979,N_6335);
nand U9360 (N_9360,N_7857,N_7458);
or U9361 (N_9361,N_7386,N_6669);
and U9362 (N_9362,N_7604,N_7812);
nor U9363 (N_9363,N_6918,N_7500);
and U9364 (N_9364,N_8799,N_6299);
nor U9365 (N_9365,N_7121,N_7677);
or U9366 (N_9366,N_6348,N_8428);
nor U9367 (N_9367,N_6333,N_7426);
nand U9368 (N_9368,N_8141,N_6017);
xnor U9369 (N_9369,N_8019,N_8584);
nand U9370 (N_9370,N_7638,N_8720);
or U9371 (N_9371,N_8143,N_7922);
nand U9372 (N_9372,N_8738,N_8884);
nor U9373 (N_9373,N_6061,N_6209);
and U9374 (N_9374,N_6806,N_8038);
nor U9375 (N_9375,N_8723,N_6074);
nor U9376 (N_9376,N_8313,N_6422);
or U9377 (N_9377,N_8962,N_6415);
xor U9378 (N_9378,N_6543,N_8705);
xnor U9379 (N_9379,N_6295,N_6194);
nor U9380 (N_9380,N_7650,N_6029);
nor U9381 (N_9381,N_6668,N_7390);
nor U9382 (N_9382,N_7871,N_6334);
and U9383 (N_9383,N_7738,N_7945);
and U9384 (N_9384,N_6043,N_6643);
nor U9385 (N_9385,N_7555,N_8030);
or U9386 (N_9386,N_7698,N_8206);
nand U9387 (N_9387,N_8631,N_7425);
nor U9388 (N_9388,N_8996,N_8010);
or U9389 (N_9389,N_8714,N_8770);
and U9390 (N_9390,N_8800,N_6426);
or U9391 (N_9391,N_8887,N_7559);
nand U9392 (N_9392,N_6033,N_7149);
and U9393 (N_9393,N_6035,N_6147);
nand U9394 (N_9394,N_7104,N_7203);
or U9395 (N_9395,N_6621,N_7157);
nor U9396 (N_9396,N_6094,N_8939);
nand U9397 (N_9397,N_6110,N_7066);
nand U9398 (N_9398,N_7954,N_8868);
nand U9399 (N_9399,N_6397,N_6237);
or U9400 (N_9400,N_7239,N_8511);
and U9401 (N_9401,N_6159,N_7093);
or U9402 (N_9402,N_6104,N_6206);
or U9403 (N_9403,N_8808,N_8227);
nand U9404 (N_9404,N_7660,N_8346);
or U9405 (N_9405,N_7793,N_8958);
xnor U9406 (N_9406,N_6203,N_7889);
nand U9407 (N_9407,N_6273,N_8877);
or U9408 (N_9408,N_7571,N_6700);
nand U9409 (N_9409,N_8566,N_6645);
and U9410 (N_9410,N_7106,N_7083);
nor U9411 (N_9411,N_7959,N_6305);
or U9412 (N_9412,N_6090,N_7903);
nor U9413 (N_9413,N_7979,N_8984);
and U9414 (N_9414,N_8509,N_8442);
nor U9415 (N_9415,N_6835,N_6932);
or U9416 (N_9416,N_8685,N_7599);
and U9417 (N_9417,N_8162,N_6649);
nor U9418 (N_9418,N_8140,N_6860);
nand U9419 (N_9419,N_7717,N_8338);
and U9420 (N_9420,N_6863,N_7332);
nand U9421 (N_9421,N_6732,N_7346);
or U9422 (N_9422,N_6945,N_6842);
or U9423 (N_9423,N_7409,N_7381);
nor U9424 (N_9424,N_7108,N_6640);
xnor U9425 (N_9425,N_8524,N_7743);
nand U9426 (N_9426,N_8763,N_7833);
nor U9427 (N_9427,N_8842,N_8530);
nand U9428 (N_9428,N_8935,N_7662);
xnor U9429 (N_9429,N_8721,N_8789);
nand U9430 (N_9430,N_6439,N_8484);
nand U9431 (N_9431,N_7041,N_8471);
or U9432 (N_9432,N_6312,N_6387);
and U9433 (N_9433,N_8238,N_6024);
or U9434 (N_9434,N_7694,N_8840);
nor U9435 (N_9435,N_8664,N_7078);
or U9436 (N_9436,N_7146,N_6195);
xnor U9437 (N_9437,N_6795,N_6392);
nor U9438 (N_9438,N_7270,N_6007);
nor U9439 (N_9439,N_6247,N_7010);
xnor U9440 (N_9440,N_8400,N_7724);
or U9441 (N_9441,N_8615,N_7873);
nor U9442 (N_9442,N_6277,N_6111);
nand U9443 (N_9443,N_6630,N_6566);
nand U9444 (N_9444,N_6204,N_7718);
nand U9445 (N_9445,N_8716,N_7004);
and U9446 (N_9446,N_6143,N_8293);
or U9447 (N_9447,N_7999,N_6369);
xor U9448 (N_9448,N_7699,N_8463);
nor U9449 (N_9449,N_8196,N_6911);
nand U9450 (N_9450,N_6935,N_6067);
nor U9451 (N_9451,N_7037,N_7612);
xnor U9452 (N_9452,N_6984,N_8097);
and U9453 (N_9453,N_6644,N_7540);
and U9454 (N_9454,N_8462,N_8931);
nand U9455 (N_9455,N_8945,N_8797);
xnor U9456 (N_9456,N_6032,N_6785);
or U9457 (N_9457,N_6404,N_8975);
or U9458 (N_9458,N_8850,N_7934);
nor U9459 (N_9459,N_7632,N_8706);
or U9460 (N_9460,N_8311,N_7181);
or U9461 (N_9461,N_8784,N_8678);
or U9462 (N_9462,N_6018,N_8107);
and U9463 (N_9463,N_8865,N_8226);
and U9464 (N_9464,N_8560,N_8963);
nand U9465 (N_9465,N_6364,N_6331);
xnor U9466 (N_9466,N_6438,N_7443);
nand U9467 (N_9467,N_8382,N_7991);
nand U9468 (N_9468,N_7970,N_6958);
nor U9469 (N_9469,N_6232,N_8929);
nor U9470 (N_9470,N_7536,N_7317);
nand U9471 (N_9471,N_7207,N_6816);
nor U9472 (N_9472,N_6174,N_8473);
or U9473 (N_9473,N_8229,N_7080);
xor U9474 (N_9474,N_7055,N_7564);
nand U9475 (N_9475,N_8740,N_7523);
nand U9476 (N_9476,N_6792,N_7842);
nand U9477 (N_9477,N_8924,N_8389);
or U9478 (N_9478,N_8075,N_7212);
nand U9479 (N_9479,N_8824,N_8623);
nand U9480 (N_9480,N_8911,N_8816);
nand U9481 (N_9481,N_8696,N_7577);
or U9482 (N_9482,N_7583,N_8660);
nand U9483 (N_9483,N_6080,N_8750);
nor U9484 (N_9484,N_8955,N_7896);
nand U9485 (N_9485,N_7043,N_8912);
nor U9486 (N_9486,N_7325,N_6300);
nand U9487 (N_9487,N_8900,N_8296);
nor U9488 (N_9488,N_7097,N_8950);
nor U9489 (N_9489,N_8441,N_8079);
and U9490 (N_9490,N_7667,N_7133);
nand U9491 (N_9491,N_7005,N_7163);
nor U9492 (N_9492,N_7261,N_7665);
and U9493 (N_9493,N_6742,N_7144);
nand U9494 (N_9494,N_7534,N_7730);
nand U9495 (N_9495,N_7410,N_8905);
and U9496 (N_9496,N_7418,N_8225);
nor U9497 (N_9497,N_7349,N_6243);
and U9498 (N_9498,N_6192,N_6282);
nand U9499 (N_9499,N_8377,N_8349);
nor U9500 (N_9500,N_6576,N_7818);
and U9501 (N_9501,N_7265,N_8490);
nor U9502 (N_9502,N_7924,N_8059);
or U9503 (N_9503,N_8031,N_6810);
nand U9504 (N_9504,N_8961,N_6553);
nor U9505 (N_9505,N_7077,N_6730);
or U9506 (N_9506,N_8150,N_7701);
or U9507 (N_9507,N_6504,N_6370);
nand U9508 (N_9508,N_7044,N_6874);
nor U9509 (N_9509,N_7021,N_7065);
or U9510 (N_9510,N_6279,N_6485);
nand U9511 (N_9511,N_6774,N_7878);
or U9512 (N_9512,N_6658,N_6001);
or U9513 (N_9513,N_6116,N_7487);
and U9514 (N_9514,N_6663,N_7636);
xor U9515 (N_9515,N_7777,N_7920);
and U9516 (N_9516,N_7664,N_8535);
nand U9517 (N_9517,N_8314,N_8676);
nor U9518 (N_9518,N_8693,N_8083);
or U9519 (N_9519,N_8907,N_6840);
nor U9520 (N_9520,N_7118,N_6961);
nand U9521 (N_9521,N_8047,N_8657);
or U9522 (N_9522,N_8053,N_7562);
xor U9523 (N_9523,N_8456,N_7469);
and U9524 (N_9524,N_8255,N_8671);
nand U9525 (N_9525,N_8500,N_6494);
and U9526 (N_9526,N_6286,N_6465);
and U9527 (N_9527,N_7854,N_8151);
nor U9528 (N_9528,N_8606,N_7981);
and U9529 (N_9529,N_7088,N_6851);
and U9530 (N_9530,N_7232,N_8451);
nand U9531 (N_9531,N_7888,N_8245);
nor U9532 (N_9532,N_7127,N_8557);
nand U9533 (N_9533,N_7247,N_6587);
nor U9534 (N_9534,N_7289,N_8017);
or U9535 (N_9535,N_8210,N_8990);
and U9536 (N_9536,N_6971,N_8622);
xor U9537 (N_9537,N_6712,N_7419);
or U9538 (N_9538,N_7006,N_8289);
nor U9539 (N_9539,N_8804,N_7776);
or U9540 (N_9540,N_6400,N_8639);
nor U9541 (N_9541,N_6081,N_7126);
or U9542 (N_9542,N_7414,N_6350);
nor U9543 (N_9543,N_7823,N_8248);
and U9544 (N_9544,N_6790,N_7729);
xnor U9545 (N_9545,N_7230,N_8064);
nand U9546 (N_9546,N_7867,N_7576);
nor U9547 (N_9547,N_7630,N_8616);
and U9548 (N_9548,N_8587,N_8426);
and U9549 (N_9549,N_6895,N_6373);
nor U9550 (N_9550,N_8108,N_7111);
and U9551 (N_9551,N_6904,N_7048);
nor U9552 (N_9552,N_6254,N_7298);
nor U9553 (N_9553,N_7875,N_7803);
nor U9554 (N_9554,N_8967,N_6118);
and U9555 (N_9555,N_8375,N_7405);
or U9556 (N_9556,N_7047,N_6593);
nor U9557 (N_9557,N_7360,N_7218);
nor U9558 (N_9558,N_6028,N_8734);
nor U9559 (N_9559,N_6040,N_8957);
and U9560 (N_9560,N_7502,N_6855);
or U9561 (N_9561,N_8034,N_7084);
nor U9562 (N_9562,N_7847,N_7319);
nand U9563 (N_9563,N_6646,N_6222);
or U9564 (N_9564,N_7728,N_8420);
or U9565 (N_9565,N_8332,N_7033);
and U9566 (N_9566,N_8046,N_7392);
or U9567 (N_9567,N_8305,N_8658);
nand U9568 (N_9568,N_8677,N_8921);
and U9569 (N_9569,N_7156,N_8915);
and U9570 (N_9570,N_7879,N_8687);
nand U9571 (N_9571,N_6169,N_8916);
nand U9572 (N_9572,N_8707,N_8391);
nor U9573 (N_9573,N_6886,N_7737);
nor U9574 (N_9574,N_8284,N_7770);
nor U9575 (N_9575,N_6048,N_6157);
nand U9576 (N_9576,N_6434,N_7095);
nor U9577 (N_9577,N_7740,N_8817);
or U9578 (N_9578,N_8055,N_8662);
nor U9579 (N_9579,N_8977,N_6954);
and U9580 (N_9580,N_7892,N_8948);
nor U9581 (N_9581,N_7150,N_6575);
nor U9582 (N_9582,N_8251,N_7584);
nor U9583 (N_9583,N_7956,N_6936);
xnor U9584 (N_9584,N_7794,N_7200);
nand U9585 (N_9585,N_6873,N_8312);
or U9586 (N_9586,N_6831,N_6763);
nand U9587 (N_9587,N_8686,N_6099);
nor U9588 (N_9588,N_8883,N_6951);
or U9589 (N_9589,N_6580,N_7166);
nor U9590 (N_9590,N_8614,N_8209);
and U9591 (N_9591,N_6022,N_8396);
and U9592 (N_9592,N_7613,N_8891);
or U9593 (N_9593,N_8532,N_6520);
and U9594 (N_9594,N_8564,N_7515);
nand U9595 (N_9595,N_7902,N_7199);
nor U9596 (N_9596,N_7915,N_6200);
and U9597 (N_9597,N_6676,N_6687);
or U9598 (N_9598,N_7479,N_7815);
and U9599 (N_9599,N_8812,N_6767);
nand U9600 (N_9600,N_8937,N_6098);
nand U9601 (N_9601,N_6980,N_6561);
nor U9602 (N_9602,N_6482,N_6849);
xor U9603 (N_9603,N_8482,N_8003);
xor U9604 (N_9604,N_7208,N_7046);
and U9605 (N_9605,N_7026,N_7383);
nor U9606 (N_9606,N_7277,N_7241);
and U9607 (N_9607,N_6705,N_8641);
or U9608 (N_9608,N_6284,N_6639);
or U9609 (N_9609,N_8859,N_7686);
nor U9610 (N_9610,N_6266,N_6451);
or U9611 (N_9611,N_6987,N_6256);
nor U9612 (N_9612,N_7090,N_6016);
nor U9613 (N_9613,N_8411,N_8563);
or U9614 (N_9614,N_8553,N_8586);
and U9615 (N_9615,N_7950,N_8117);
or U9616 (N_9616,N_7894,N_6215);
nor U9617 (N_9617,N_6574,N_8022);
nand U9618 (N_9618,N_7552,N_6699);
xnor U9619 (N_9619,N_6483,N_6518);
or U9620 (N_9620,N_8193,N_8149);
or U9621 (N_9621,N_7765,N_8820);
and U9622 (N_9622,N_7675,N_6534);
nor U9623 (N_9623,N_8084,N_8637);
and U9624 (N_9624,N_7659,N_6068);
or U9625 (N_9625,N_8610,N_8956);
or U9626 (N_9626,N_7030,N_8646);
nand U9627 (N_9627,N_8531,N_7708);
nand U9628 (N_9628,N_7233,N_7279);
or U9629 (N_9629,N_7049,N_6920);
and U9630 (N_9630,N_6884,N_6662);
or U9631 (N_9631,N_6659,N_8822);
and U9632 (N_9632,N_6101,N_6131);
or U9633 (N_9633,N_8335,N_6010);
and U9634 (N_9634,N_8134,N_6814);
or U9635 (N_9635,N_6180,N_8768);
and U9636 (N_9636,N_8792,N_6870);
nor U9637 (N_9637,N_8858,N_6697);
and U9638 (N_9638,N_8172,N_6013);
nand U9639 (N_9639,N_7886,N_8300);
or U9640 (N_9640,N_6233,N_8892);
or U9641 (N_9641,N_8384,N_8197);
nor U9642 (N_9642,N_6549,N_7171);
or U9643 (N_9643,N_8039,N_7643);
nor U9644 (N_9644,N_8307,N_7532);
or U9645 (N_9645,N_7139,N_7389);
or U9646 (N_9646,N_6667,N_6393);
xnor U9647 (N_9647,N_8065,N_7101);
and U9648 (N_9648,N_7141,N_8683);
or U9649 (N_9649,N_7953,N_6826);
or U9650 (N_9650,N_6413,N_8722);
nor U9651 (N_9651,N_8205,N_8691);
and U9652 (N_9652,N_8947,N_7130);
and U9653 (N_9653,N_6340,N_8846);
nor U9654 (N_9654,N_6251,N_8670);
or U9655 (N_9655,N_7594,N_7681);
or U9656 (N_9656,N_7267,N_7185);
and U9657 (N_9657,N_7444,N_6631);
nand U9658 (N_9658,N_8133,N_6977);
nand U9659 (N_9659,N_6488,N_7228);
nor U9660 (N_9660,N_8477,N_8459);
and U9661 (N_9661,N_8866,N_6625);
nor U9662 (N_9662,N_6515,N_8058);
xor U9663 (N_9663,N_7348,N_6710);
nand U9664 (N_9664,N_7829,N_8579);
xor U9665 (N_9665,N_8880,N_8447);
nor U9666 (N_9666,N_7161,N_8651);
nand U9667 (N_9667,N_8514,N_6347);
xnor U9668 (N_9668,N_8562,N_6121);
nand U9669 (N_9669,N_8968,N_7884);
nor U9670 (N_9670,N_6368,N_7911);
and U9671 (N_9671,N_8597,N_8213);
or U9672 (N_9672,N_6020,N_7671);
nand U9673 (N_9673,N_7690,N_6150);
and U9674 (N_9674,N_7804,N_8237);
nand U9675 (N_9675,N_8994,N_6225);
or U9676 (N_9676,N_6559,N_8115);
and U9677 (N_9677,N_7845,N_6466);
nor U9678 (N_9678,N_6417,N_6782);
nand U9679 (N_9679,N_7455,N_6942);
nand U9680 (N_9680,N_8228,N_6521);
nand U9681 (N_9681,N_8669,N_7427);
and U9682 (N_9682,N_8130,N_8946);
or U9683 (N_9683,N_6309,N_6967);
nor U9684 (N_9684,N_8419,N_8457);
or U9685 (N_9685,N_7151,N_7273);
and U9686 (N_9686,N_7096,N_8001);
xor U9687 (N_9687,N_8758,N_7791);
and U9688 (N_9688,N_6337,N_7678);
nand U9689 (N_9689,N_6208,N_7748);
nor U9690 (N_9690,N_6229,N_8528);
or U9691 (N_9691,N_6144,N_7340);
and U9692 (N_9692,N_8592,N_7222);
or U9693 (N_9693,N_7932,N_8165);
nand U9694 (N_9694,N_6623,N_6390);
and U9695 (N_9695,N_7997,N_6809);
and U9696 (N_9696,N_6100,N_6862);
or U9697 (N_9697,N_6986,N_7961);
xnor U9698 (N_9698,N_8043,N_8348);
nand U9699 (N_9699,N_7086,N_6619);
or U9700 (N_9700,N_7020,N_7484);
or U9701 (N_9701,N_8029,N_8684);
nor U9702 (N_9702,N_7099,N_7974);
and U9703 (N_9703,N_6183,N_7058);
nor U9704 (N_9704,N_6923,N_6125);
nand U9705 (N_9705,N_8886,N_8015);
and U9706 (N_9706,N_7707,N_6959);
or U9707 (N_9707,N_6755,N_7211);
and U9708 (N_9708,N_7567,N_7359);
nand U9709 (N_9709,N_7909,N_8061);
or U9710 (N_9710,N_6950,N_7712);
nand U9711 (N_9711,N_8598,N_6095);
nand U9712 (N_9712,N_6864,N_7014);
nand U9713 (N_9713,N_6149,N_6784);
nor U9714 (N_9714,N_6296,N_7980);
and U9715 (N_9715,N_6178,N_8726);
nor U9716 (N_9716,N_8392,N_6341);
xor U9717 (N_9717,N_7939,N_6262);
nor U9718 (N_9718,N_7252,N_8830);
or U9719 (N_9719,N_7304,N_7852);
and U9720 (N_9720,N_6078,N_6012);
nand U9721 (N_9721,N_7499,N_8926);
nand U9722 (N_9722,N_6153,N_7828);
xnor U9723 (N_9723,N_8550,N_7123);
nor U9724 (N_9724,N_8266,N_7456);
nor U9725 (N_9725,N_6271,N_7351);
nor U9726 (N_9726,N_7813,N_7056);
and U9727 (N_9727,N_6704,N_6060);
and U9728 (N_9728,N_6151,N_7966);
or U9729 (N_9729,N_6678,N_6996);
or U9730 (N_9730,N_6410,N_6899);
and U9731 (N_9731,N_6261,N_7497);
nor U9732 (N_9732,N_8012,N_8275);
nor U9733 (N_9733,N_6779,N_7749);
and U9734 (N_9734,N_8443,N_8694);
nand U9735 (N_9735,N_8777,N_6314);
xor U9736 (N_9736,N_7744,N_7007);
nor U9737 (N_9737,N_6476,N_6066);
nand U9738 (N_9738,N_6915,N_7285);
xor U9739 (N_9739,N_8166,N_8973);
or U9740 (N_9740,N_8368,N_6586);
xor U9741 (N_9741,N_8152,N_6383);
nand U9742 (N_9742,N_8282,N_6182);
xnor U9743 (N_9743,N_7448,N_6089);
and U9744 (N_9744,N_8188,N_8987);
nor U9745 (N_9745,N_8704,N_6495);
nand U9746 (N_9746,N_6773,N_6461);
nand U9747 (N_9747,N_8406,N_6197);
nand U9748 (N_9748,N_8733,N_8665);
or U9749 (N_9749,N_6939,N_8409);
nor U9750 (N_9750,N_7061,N_6955);
nor U9751 (N_9751,N_8413,N_7965);
and U9752 (N_9752,N_8690,N_8802);
nand U9753 (N_9753,N_7361,N_6902);
or U9754 (N_9754,N_7697,N_7398);
nor U9755 (N_9755,N_6378,N_7624);
xor U9756 (N_9756,N_6470,N_6719);
or U9757 (N_9757,N_6396,N_8236);
xnor U9758 (N_9758,N_6351,N_8876);
or U9759 (N_9759,N_7358,N_6807);
and U9760 (N_9760,N_8005,N_8161);
nor U9761 (N_9761,N_7913,N_6801);
and U9762 (N_9762,N_6352,N_6731);
nand U9763 (N_9763,N_8173,N_7994);
nand U9764 (N_9764,N_6829,N_7769);
nor U9765 (N_9765,N_8575,N_8381);
nor U9766 (N_9766,N_6298,N_6185);
nor U9767 (N_9767,N_7040,N_8109);
and U9768 (N_9768,N_8952,N_7538);
and U9769 (N_9769,N_6709,N_7214);
nand U9770 (N_9770,N_7063,N_7657);
nor U9771 (N_9771,N_8753,N_8527);
nor U9772 (N_9772,N_6103,N_6749);
nor U9773 (N_9773,N_7178,N_7012);
nand U9774 (N_9774,N_7547,N_7362);
or U9775 (N_9775,N_8634,N_7245);
nand U9776 (N_9776,N_8249,N_7013);
nor U9777 (N_9777,N_7365,N_8089);
nor U9778 (N_9778,N_7341,N_8208);
nand U9779 (N_9779,N_7468,N_8224);
nand U9780 (N_9780,N_8106,N_8936);
nor U9781 (N_9781,N_6375,N_6353);
nand U9782 (N_9782,N_7071,N_8570);
and U9783 (N_9783,N_8841,N_8179);
nor U9784 (N_9784,N_7860,N_7034);
and U9785 (N_9785,N_6427,N_8630);
nor U9786 (N_9786,N_6199,N_7423);
and U9787 (N_9787,N_6885,N_6059);
xor U9788 (N_9788,N_8520,N_6822);
nor U9789 (N_9789,N_7856,N_6498);
nand U9790 (N_9790,N_7259,N_8980);
nor U9791 (N_9791,N_6377,N_7883);
nand U9792 (N_9792,N_7926,N_8747);
nand U9793 (N_9793,N_7482,N_8698);
or U9794 (N_9794,N_7841,N_6223);
or U9795 (N_9795,N_8174,N_6747);
nor U9796 (N_9796,N_7768,N_8088);
xor U9797 (N_9797,N_6547,N_6671);
xnor U9798 (N_9798,N_7679,N_6857);
nor U9799 (N_9799,N_8024,N_6698);
or U9800 (N_9800,N_8320,N_7364);
and U9801 (N_9801,N_8127,N_8177);
nor U9802 (N_9802,N_7076,N_8663);
or U9803 (N_9803,N_6847,N_6102);
nor U9804 (N_9804,N_6647,N_6051);
and U9805 (N_9805,N_7637,N_7572);
and U9806 (N_9806,N_8274,N_8002);
or U9807 (N_9807,N_8365,N_7802);
nor U9808 (N_9808,N_6268,N_6946);
and U9809 (N_9809,N_8230,N_6496);
or U9810 (N_9810,N_8794,N_8708);
nand U9811 (N_9811,N_6744,N_6615);
nor U9812 (N_9812,N_8330,N_6692);
and U9813 (N_9813,N_6591,N_8114);
nor U9814 (N_9814,N_7695,N_7510);
nor U9815 (N_9815,N_8077,N_6956);
and U9816 (N_9816,N_6173,N_7355);
and U9817 (N_9817,N_7542,N_7269);
and U9818 (N_9818,N_7563,N_6841);
nor U9819 (N_9819,N_7880,N_8187);
or U9820 (N_9820,N_6391,N_7373);
xor U9821 (N_9821,N_6242,N_6014);
nor U9822 (N_9822,N_6581,N_8832);
nor U9823 (N_9823,N_7696,N_7983);
nand U9824 (N_9824,N_7312,N_8087);
or U9825 (N_9825,N_8974,N_8105);
nor U9826 (N_9826,N_7721,N_7976);
nand U9827 (N_9827,N_7774,N_7822);
nor U9828 (N_9828,N_7017,N_6867);
nor U9829 (N_9829,N_7440,N_7792);
nor U9830 (N_9830,N_8596,N_8254);
nor U9831 (N_9831,N_6793,N_8119);
xnor U9832 (N_9832,N_7674,N_7767);
nor U9833 (N_9833,N_8746,N_7557);
nand U9834 (N_9834,N_8901,N_6263);
nor U9835 (N_9835,N_7606,N_8360);
and U9836 (N_9836,N_6850,N_7471);
nand U9837 (N_9837,N_8006,N_7642);
or U9838 (N_9838,N_7713,N_7616);
xor U9839 (N_9839,N_6633,N_6539);
xor U9840 (N_9840,N_6409,N_6319);
or U9841 (N_9841,N_8417,N_6287);
and U9842 (N_9842,N_7135,N_6152);
xor U9843 (N_9843,N_8018,N_8168);
nor U9844 (N_9844,N_7402,N_7541);
nand U9845 (N_9845,N_6170,N_8513);
and U9846 (N_9846,N_7371,N_6441);
and U9847 (N_9847,N_7984,N_7741);
nand U9848 (N_9848,N_7949,N_7334);
nor U9849 (N_9849,N_6924,N_7874);
nand U9850 (N_9850,N_7182,N_7190);
nor U9851 (N_9851,N_6430,N_6303);
or U9852 (N_9852,N_7132,N_7169);
and U9853 (N_9853,N_8350,N_6189);
nand U9854 (N_9854,N_8233,N_6346);
nand U9855 (N_9855,N_6622,N_8169);
and U9856 (N_9856,N_6680,N_6761);
nor U9857 (N_9857,N_7520,N_8860);
or U9858 (N_9858,N_7158,N_8906);
nand U9859 (N_9859,N_6708,N_7445);
xor U9860 (N_9860,N_7321,N_8599);
nand U9861 (N_9861,N_7783,N_6210);
nand U9862 (N_9862,N_7714,N_7619);
or U9863 (N_9863,N_7439,N_7008);
nand U9864 (N_9864,N_8062,N_8659);
nor U9865 (N_9865,N_8608,N_6856);
nand U9866 (N_9866,N_6789,N_7838);
or U9867 (N_9867,N_6599,N_7719);
nor U9868 (N_9868,N_7683,N_6579);
nand U9869 (N_9869,N_6903,N_7378);
and U9870 (N_9870,N_7174,N_7240);
nand U9871 (N_9871,N_7639,N_6993);
nor U9872 (N_9872,N_7938,N_7927);
or U9873 (N_9873,N_7179,N_8111);
nand U9874 (N_9874,N_6459,N_7333);
xnor U9875 (N_9875,N_8319,N_6714);
and U9876 (N_9876,N_6927,N_7197);
nand U9877 (N_9877,N_8074,N_6838);
and U9878 (N_9878,N_7311,N_7772);
or U9879 (N_9879,N_6443,N_7089);
and U9880 (N_9880,N_8976,N_7819);
xnor U9881 (N_9881,N_7215,N_8435);
xnor U9882 (N_9882,N_8867,N_6843);
nand U9883 (N_9883,N_7193,N_8515);
and U9884 (N_9884,N_6344,N_8668);
or U9885 (N_9885,N_8666,N_6091);
nand U9886 (N_9886,N_8533,N_7238);
or U9887 (N_9887,N_7148,N_6490);
nand U9888 (N_9888,N_8026,N_6468);
and U9889 (N_9889,N_6276,N_8415);
and U9890 (N_9890,N_6313,N_6734);
and U9891 (N_9891,N_7219,N_6565);
nand U9892 (N_9892,N_7025,N_6648);
nor U9893 (N_9893,N_7180,N_8076);
nand U9894 (N_9894,N_7103,N_7585);
nor U9895 (N_9895,N_7921,N_6766);
nor U9896 (N_9896,N_7566,N_7196);
nand U9897 (N_9897,N_7601,N_8460);
nand U9898 (N_9898,N_6845,N_8536);
nor U9899 (N_9899,N_6982,N_8559);
or U9900 (N_9900,N_6234,N_8000);
nor U9901 (N_9901,N_7597,N_6052);
and U9902 (N_9902,N_8835,N_6207);
or U9903 (N_9903,N_6721,N_6191);
and U9904 (N_9904,N_8481,N_6728);
or U9905 (N_9905,N_7570,N_7655);
or U9906 (N_9906,N_8439,N_6293);
and U9907 (N_9907,N_6041,N_7995);
and U9908 (N_9908,N_8434,N_8672);
and U9909 (N_9909,N_7483,N_8781);
nand U9910 (N_9910,N_6681,N_8624);
nand U9911 (N_9911,N_7944,N_7509);
and U9912 (N_9912,N_7391,N_8356);
and U9913 (N_9913,N_7116,N_6693);
xor U9914 (N_9914,N_6743,N_6634);
nor U9915 (N_9915,N_6244,N_7476);
nor U9916 (N_9916,N_6733,N_6475);
nand U9917 (N_9917,N_8729,N_7168);
nor U9918 (N_9918,N_7430,N_7758);
and U9919 (N_9919,N_8821,N_6327);
nor U9920 (N_9920,N_6187,N_6736);
or U9921 (N_9921,N_7620,N_8604);
nand U9922 (N_9922,N_6656,N_7377);
or U9923 (N_9923,N_7862,N_8113);
nor U9924 (N_9924,N_8904,N_6399);
nor U9925 (N_9925,N_6930,N_6786);
xor U9926 (N_9926,N_6326,N_8574);
nand U9927 (N_9927,N_6003,N_7786);
nand U9928 (N_9928,N_6045,N_7958);
nand U9929 (N_9929,N_8979,N_7303);
and U9930 (N_9930,N_6503,N_8090);
nand U9931 (N_9931,N_8642,N_6117);
and U9932 (N_9932,N_6231,N_7263);
nand U9933 (N_9933,N_8908,N_6703);
nor U9934 (N_9934,N_7908,N_6355);
nor U9935 (N_9935,N_8710,N_7153);
or U9936 (N_9936,N_7928,N_6651);
nor U9937 (N_9937,N_6938,N_6919);
nand U9938 (N_9938,N_6328,N_7969);
or U9939 (N_9939,N_7827,N_6006);
nor U9940 (N_9940,N_8241,N_7560);
or U9941 (N_9941,N_6038,N_6349);
and U9942 (N_9942,N_6718,N_6205);
nand U9943 (N_9943,N_6880,N_7990);
xnor U9944 (N_9944,N_6752,N_6990);
nand U9945 (N_9945,N_7282,N_6545);
and U9946 (N_9946,N_7459,N_7731);
nor U9947 (N_9947,N_7314,N_7323);
nand U9948 (N_9948,N_6866,N_8798);
nand U9949 (N_9949,N_6595,N_6981);
nand U9950 (N_9950,N_8857,N_8544);
or U9951 (N_9951,N_8703,N_6228);
nor U9952 (N_9952,N_8752,N_6075);
and U9953 (N_9953,N_8281,N_8576);
or U9954 (N_9954,N_6240,N_8480);
nand U9955 (N_9955,N_6943,N_6457);
and U9956 (N_9956,N_6727,N_7644);
or U9957 (N_9957,N_6998,N_8765);
or U9958 (N_9958,N_8492,N_7347);
and U9959 (N_9959,N_8279,N_8124);
nor U9960 (N_9960,N_6398,N_6130);
nor U9961 (N_9961,N_8551,N_7490);
nand U9962 (N_9962,N_6983,N_7075);
and U9963 (N_9963,N_7820,N_6278);
xor U9964 (N_9964,N_8216,N_8357);
and U9965 (N_9965,N_7031,N_7302);
nor U9966 (N_9966,N_8045,N_6177);
nand U9967 (N_9967,N_6401,N_8429);
xnor U9968 (N_9968,N_6720,N_6921);
nand U9969 (N_9969,N_8371,N_7489);
nand U9970 (N_9970,N_8526,N_6198);
or U9971 (N_9971,N_8170,N_8650);
nand U9972 (N_9972,N_8863,N_6624);
nor U9973 (N_9973,N_7401,N_8491);
nor U9974 (N_9974,N_6825,N_6137);
nand U9975 (N_9975,N_6552,N_8054);
or U9976 (N_9976,N_8793,N_6887);
nand U9977 (N_9977,N_8783,N_8934);
xnor U9978 (N_9978,N_7835,N_8534);
and U9979 (N_9979,N_8370,N_7752);
nand U9980 (N_9980,N_7475,N_7094);
nor U9981 (N_9981,N_7501,N_6526);
and U9982 (N_9982,N_6320,N_6757);
xor U9983 (N_9983,N_6164,N_8648);
or U9984 (N_9984,N_7556,N_7651);
nor U9985 (N_9985,N_8521,N_7275);
or U9986 (N_9986,N_7973,N_6928);
or U9987 (N_9987,N_7876,N_6564);
nor U9988 (N_9988,N_8294,N_6788);
nand U9989 (N_9989,N_6808,N_7175);
nand U9990 (N_9990,N_7452,N_6568);
nor U9991 (N_9991,N_7789,N_8393);
xor U9992 (N_9992,N_8432,N_6097);
and U9993 (N_9993,N_6395,N_6324);
nand U9994 (N_9994,N_8780,N_8749);
and U9995 (N_9995,N_6227,N_7870);
nor U9996 (N_9996,N_8092,N_8653);
and U9997 (N_9997,N_6865,N_7977);
or U9998 (N_9998,N_8098,N_7293);
nand U9999 (N_9999,N_8519,N_8070);
nor U10000 (N_10000,N_7531,N_7881);
xor U10001 (N_10001,N_6345,N_6436);
xnor U10002 (N_10002,N_7784,N_8836);
nand U10003 (N_10003,N_7548,N_6196);
nor U10004 (N_10004,N_6513,N_6069);
nor U10005 (N_10005,N_6762,N_8806);
and U10006 (N_10006,N_6452,N_6250);
or U10007 (N_10007,N_7024,N_7640);
nand U10008 (N_10008,N_6034,N_7198);
or U10009 (N_10009,N_6997,N_8203);
nand U10010 (N_10010,N_6878,N_6053);
nor U10011 (N_10011,N_6556,N_7631);
and U10012 (N_10012,N_8568,N_7916);
nand U10013 (N_10013,N_7327,N_8815);
nor U10014 (N_10014,N_7449,N_8060);
or U10015 (N_10015,N_7268,N_7308);
xnor U10016 (N_10016,N_8341,N_7676);
nand U10017 (N_10017,N_7299,N_7957);
and U10018 (N_10018,N_6894,N_8427);
nor U10019 (N_10019,N_6109,N_6765);
xnor U10020 (N_10020,N_6818,N_7112);
nor U10021 (N_10021,N_8163,N_8643);
nor U10022 (N_10022,N_8125,N_6382);
nand U10023 (N_10023,N_7761,N_7415);
nor U10024 (N_10024,N_6246,N_6023);
nand U10025 (N_10025,N_7271,N_8221);
xor U10026 (N_10026,N_6481,N_7848);
xnor U10027 (N_10027,N_8590,N_8775);
and U10028 (N_10028,N_8405,N_7811);
xor U10029 (N_10029,N_7527,N_6464);
and U10030 (N_10030,N_7292,N_6960);
nand U10031 (N_10031,N_8037,N_6944);
xnor U10032 (N_10032,N_6685,N_7331);
or U10033 (N_10033,N_6129,N_6162);
or U10034 (N_10034,N_6608,N_6267);
or U10035 (N_10035,N_6962,N_7256);
nor U10036 (N_10036,N_7438,N_6063);
nor U10037 (N_10037,N_6027,N_6047);
nand U10038 (N_10038,N_6626,N_8364);
xnor U10039 (N_10039,N_8337,N_7201);
and U10040 (N_10040,N_7808,N_6689);
or U10041 (N_10041,N_7907,N_6828);
nand U10042 (N_10042,N_6567,N_7453);
or U10043 (N_10043,N_8156,N_6450);
or U10044 (N_10044,N_7330,N_8160);
nor U10045 (N_10045,N_8467,N_8497);
and U10046 (N_10046,N_8617,N_7669);
nor U10047 (N_10047,N_8013,N_8889);
or U10048 (N_10048,N_6512,N_7428);
or U10049 (N_10049,N_6359,N_7521);
or U10050 (N_10050,N_7887,N_7140);
or U10051 (N_10051,N_7429,N_7057);
nand U10052 (N_10052,N_6717,N_7895);
nor U10053 (N_10053,N_8298,N_6384);
nand U10054 (N_10054,N_8301,N_8522);
xnor U10055 (N_10055,N_7073,N_7473);
and U10056 (N_10056,N_7535,N_7100);
and U10057 (N_10057,N_6501,N_6188);
nor U10058 (N_10058,N_8191,N_6238);
nand U10059 (N_10059,N_6402,N_6969);
nand U10060 (N_10060,N_6419,N_6408);
nor U10061 (N_10061,N_6403,N_7380);
or U10062 (N_10062,N_6582,N_7764);
nand U10063 (N_10063,N_7224,N_8869);
nand U10064 (N_10064,N_7904,N_6269);
xor U10065 (N_10065,N_8688,N_8438);
and U10066 (N_10066,N_8157,N_6145);
and U10067 (N_10067,N_8262,N_7814);
nor U10068 (N_10068,N_6138,N_8268);
nand U10069 (N_10069,N_6906,N_8270);
nor U10070 (N_10070,N_7580,N_7119);
nor U10071 (N_10071,N_7231,N_6741);
or U10072 (N_10072,N_7011,N_8499);
nor U10073 (N_10073,N_8476,N_6907);
nor U10074 (N_10074,N_8786,N_8036);
or U10075 (N_10075,N_6486,N_7474);
and U10076 (N_10076,N_6529,N_8016);
or U10077 (N_10077,N_7910,N_8609);
or U10078 (N_10078,N_8629,N_6085);
or U10079 (N_10079,N_7493,N_8591);
and U10080 (N_10080,N_7001,N_7192);
or U10081 (N_10081,N_6642,N_6084);
or U10082 (N_10082,N_6432,N_8692);
and U10083 (N_10083,N_8489,N_6965);
nand U10084 (N_10084,N_8101,N_8813);
or U10085 (N_10085,N_6239,N_6386);
nor U10086 (N_10086,N_8845,N_7433);
nor U10087 (N_10087,N_7120,N_7235);
xor U10088 (N_10088,N_6316,N_7742);
or U10089 (N_10089,N_7436,N_7914);
and U10090 (N_10090,N_7859,N_6896);
or U10091 (N_10091,N_6753,N_7496);
nand U10092 (N_10092,N_8250,N_7622);
or U10093 (N_10093,N_8235,N_6385);
nor U10094 (N_10094,N_8986,N_7614);
and U10095 (N_10095,N_6412,N_6453);
or U10096 (N_10096,N_6610,N_6970);
xnor U10097 (N_10097,N_6940,N_6119);
and U10098 (N_10098,N_8278,N_7424);
and U10099 (N_10099,N_8310,N_8023);
and U10100 (N_10100,N_7756,N_6570);
nor U10101 (N_10101,N_7504,N_6230);
and U10102 (N_10102,N_7276,N_7253);
and U10103 (N_10103,N_7763,N_8164);
nand U10104 (N_10104,N_8795,N_8239);
nand U10105 (N_10105,N_6819,N_7830);
nor U10106 (N_10106,N_8252,N_8516);
or U10107 (N_10107,N_8072,N_8063);
and U10108 (N_10108,N_6798,N_7703);
xnor U10109 (N_10109,N_8769,N_6105);
and U10110 (N_10110,N_8135,N_6585);
nor U10111 (N_10111,N_7858,N_8573);
nand U10112 (N_10112,N_7399,N_8277);
nand U10113 (N_10113,N_7946,N_7771);
nor U10114 (N_10114,N_8910,N_7587);
or U10115 (N_10115,N_8603,N_6537);
or U10116 (N_10116,N_8627,N_7975);
or U10117 (N_10117,N_8913,N_6627);
nor U10118 (N_10118,N_8978,N_7546);
and U10119 (N_10119,N_6738,N_6632);
nand U10120 (N_10120,N_6963,N_8137);
and U10121 (N_10121,N_8571,N_8727);
nor U10122 (N_10122,N_8701,N_8082);
or U10123 (N_10123,N_6106,N_8803);
or U10124 (N_10124,N_8418,N_6005);
nand U10125 (N_10125,N_6746,N_6290);
nor U10126 (N_10126,N_7315,N_8993);
or U10127 (N_10127,N_7800,N_7732);
nor U10128 (N_10128,N_6360,N_6953);
xor U10129 (N_10129,N_8788,N_6533);
nand U10130 (N_10130,N_7260,N_8110);
nor U10131 (N_10131,N_8923,N_7406);
or U10132 (N_10132,N_7726,N_7022);
or U10133 (N_10133,N_7727,N_7978);
nand U10134 (N_10134,N_8472,N_6858);
xnor U10135 (N_10135,N_6388,N_8898);
or U10136 (N_10136,N_7746,N_6852);
nand U10137 (N_10137,N_8425,N_7164);
nor U10138 (N_10138,N_6363,N_6557);
nand U10139 (N_10139,N_6653,N_6480);
xor U10140 (N_10140,N_7313,N_8539);
and U10141 (N_10141,N_7301,N_7195);
and U10142 (N_10142,N_6629,N_7258);
nor U10143 (N_10143,N_6285,N_8555);
nor U10144 (N_10144,N_8265,N_7186);
and U10145 (N_10145,N_7524,N_8818);
nor U10146 (N_10146,N_8543,N_7834);
nand U10147 (N_10147,N_6523,N_8766);
and U10148 (N_10148,N_8122,N_7831);
or U10149 (N_10149,N_7760,N_7213);
xor U10150 (N_10150,N_8198,N_6872);
or U10151 (N_10151,N_6769,N_8455);
or U10152 (N_10152,N_8020,N_6800);
or U10153 (N_10153,N_8154,N_6092);
nor U10154 (N_10154,N_6637,N_8291);
nand U10155 (N_10155,N_8626,N_8260);
and U10156 (N_10156,N_7936,N_8782);
nand U10157 (N_10157,N_7947,N_7019);
xnor U10158 (N_10158,N_6175,N_7826);
nor U10159 (N_10159,N_7633,N_8875);
nor U10160 (N_10160,N_8257,N_7754);
nand U10161 (N_10161,N_6357,N_7581);
xnor U10162 (N_10162,N_8148,N_7985);
and U10163 (N_10163,N_7751,N_8827);
and U10164 (N_10164,N_7131,N_6292);
or U10165 (N_10165,N_8897,N_8839);
nor U10166 (N_10166,N_6433,N_6407);
nand U10167 (N_10167,N_6176,N_8742);
nor U10168 (N_10168,N_8971,N_6126);
nand U10169 (N_10169,N_6511,N_6664);
and U10170 (N_10170,N_8051,N_6694);
nand U10171 (N_10171,N_7015,N_8401);
nor U10172 (N_10172,N_7039,N_8078);
and U10173 (N_10173,N_6472,N_8256);
nor U10174 (N_10174,N_6469,N_6532);
nand U10175 (N_10175,N_8048,N_8004);
or U10176 (N_10176,N_6917,N_7930);
and U10177 (N_10177,N_6890,N_8572);
nand U10178 (N_10178,N_7177,N_8864);
nor U10179 (N_10179,N_7801,N_7807);
or U10180 (N_10180,N_6751,N_6405);
and U10181 (N_10181,N_6070,N_6329);
xnor U10182 (N_10182,N_6163,N_7918);
and U10183 (N_10183,N_6054,N_6573);
xnor U10184 (N_10184,N_8811,N_7447);
nand U10185 (N_10185,N_6343,N_6096);
or U10186 (N_10186,N_6181,N_7561);
or U10187 (N_10187,N_6739,N_8805);
nand U10188 (N_10188,N_6190,N_8712);
or U10189 (N_10189,N_7353,N_6770);
nand U10190 (N_10190,N_6462,N_8207);
nand U10191 (N_10191,N_7421,N_7757);
nor U10192 (N_10192,N_7998,N_8398);
and U10193 (N_10193,N_8549,N_8632);
nor U10194 (N_10194,N_6270,N_6992);
or U10195 (N_10195,N_6008,N_7465);
and U10196 (N_10196,N_8094,N_8474);
or U10197 (N_10197,N_6112,N_7446);
nand U10198 (N_10198,N_6525,N_7649);
nor U10199 (N_10199,N_7554,N_7225);
or U10200 (N_10200,N_8155,N_7394);
nor U10201 (N_10201,N_7154,N_7085);
nor U10202 (N_10202,N_8449,N_6288);
nor U10203 (N_10203,N_7350,N_7868);
xnor U10204 (N_10204,N_8321,N_7805);
nand U10205 (N_10205,N_6994,N_7309);
and U10206 (N_10206,N_8589,N_6514);
and U10207 (N_10207,N_8997,N_7715);
or U10208 (N_10208,N_7933,N_8120);
or U10209 (N_10209,N_7778,N_7912);
nand U10210 (N_10210,N_8373,N_8204);
nor U10211 (N_10211,N_7654,N_7343);
nand U10212 (N_10212,N_6342,N_7766);
nand U10213 (N_10213,N_8290,N_8351);
nand U10214 (N_10214,N_7821,N_7155);
nor U10215 (N_10215,N_6679,N_7087);
nor U10216 (N_10216,N_8186,N_6853);
or U10217 (N_10217,N_8855,N_6764);
xor U10218 (N_10218,N_8304,N_8960);
xor U10219 (N_10219,N_7053,N_7272);
and U10220 (N_10220,N_7668,N_8717);
nor U10221 (N_10221,N_8322,N_6723);
nor U10222 (N_10222,N_8595,N_7747);
nor U10223 (N_10223,N_8132,N_8287);
and U10224 (N_10224,N_8787,N_8100);
nand U10225 (N_10225,N_7693,N_7251);
nor U10226 (N_10226,N_8611,N_7036);
or U10227 (N_10227,N_8981,N_8052);
nor U10228 (N_10228,N_7357,N_7138);
or U10229 (N_10229,N_6804,N_8896);
nand U10230 (N_10230,N_7652,N_8943);
or U10231 (N_10231,N_7578,N_6745);
and U10232 (N_10232,N_7782,N_7745);
nor U10233 (N_10233,N_6049,N_6682);
or U10234 (N_10234,N_6976,N_6846);
and U10235 (N_10235,N_8890,N_6406);
or U10236 (N_10236,N_8661,N_6304);
or U10237 (N_10237,N_7209,N_7457);
nand U10238 (N_10238,N_8445,N_7079);
and U10239 (N_10239,N_7342,N_6425);
nand U10240 (N_10240,N_7142,N_8380);
nor U10241 (N_10241,N_8273,N_7397);
and U10242 (N_10242,N_7691,N_6706);
and U10243 (N_10243,N_8404,N_6735);
xnor U10244 (N_10244,N_6026,N_8779);
and U10245 (N_10245,N_7735,N_7720);
and U10246 (N_10246,N_8159,N_7628);
nand U10247 (N_10247,N_8128,N_7670);
nand U10248 (N_10248,N_7673,N_8844);
nor U10249 (N_10249,N_7254,N_7495);
and U10250 (N_10250,N_6827,N_7799);
nand U10251 (N_10251,N_8561,N_6365);
nand U10252 (N_10252,N_7114,N_7054);
or U10253 (N_10253,N_6019,N_7110);
and U10254 (N_10254,N_8317,N_7603);
nor U10255 (N_10255,N_7167,N_7113);
or U10256 (N_10256,N_6531,N_7290);
or U10257 (N_10257,N_6184,N_6093);
or U10258 (N_10258,N_8567,N_8711);
nor U10259 (N_10259,N_7134,N_7210);
or U10260 (N_10260,N_7297,N_8323);
nand U10261 (N_10261,N_6139,N_7318);
nor U10262 (N_10262,N_7987,N_8928);
and U10263 (N_10263,N_6136,N_7537);
nor U10264 (N_10264,N_6505,N_8044);
xor U10265 (N_10265,N_8021,N_6217);
and U10266 (N_10266,N_6701,N_8066);
and U10267 (N_10267,N_8785,N_7172);
and U10268 (N_10268,N_7480,N_7091);
nor U10269 (N_10269,N_7968,N_6487);
nor U10270 (N_10270,N_6791,N_8909);
nand U10271 (N_10271,N_7159,N_7367);
and U10272 (N_10272,N_6107,N_7549);
or U10273 (N_10273,N_8761,N_7035);
or U10274 (N_10274,N_8217,N_8340);
or U10275 (N_10275,N_6824,N_8436);
nor U10276 (N_10276,N_8367,N_7853);
nor U10277 (N_10277,N_8336,N_8176);
nand U10278 (N_10278,N_6448,N_7463);
xnor U10279 (N_10279,N_7491,N_6875);
xor U10280 (N_10280,N_7284,N_8431);
and U10281 (N_10281,N_6578,N_8748);
nand U10282 (N_10282,N_8407,N_7042);
nand U10283 (N_10283,N_7753,N_8071);
xor U10284 (N_10284,N_6155,N_8399);
nor U10285 (N_10285,N_8362,N_6830);
nor U10286 (N_10286,N_7551,N_6715);
xnor U10287 (N_10287,N_8556,N_6046);
and U10288 (N_10288,N_8872,N_6036);
nor U10289 (N_10289,N_6602,N_8918);
nor U10290 (N_10290,N_8554,N_8424);
nor U10291 (N_10291,N_7526,N_6165);
xnor U10292 (N_10292,N_7363,N_6590);
nand U10293 (N_10293,N_7877,N_6079);
nor U10294 (N_10294,N_8862,N_6638);
or U10295 (N_10295,N_8942,N_7967);
or U10296 (N_10296,N_8264,N_8040);
nand U10297 (N_10297,N_8953,N_6082);
nor U10298 (N_10298,N_8743,N_6601);
nor U10299 (N_10299,N_6166,N_6922);
or U10300 (N_10300,N_7863,N_6617);
xnor U10301 (N_10301,N_6750,N_6245);
xnor U10302 (N_10302,N_8334,N_7943);
or U10303 (N_10303,N_6837,N_6991);
and U10304 (N_10304,N_7255,N_8757);
nand U10305 (N_10305,N_8523,N_8085);
xor U10306 (N_10306,N_6891,N_8200);
nand U10307 (N_10307,N_6497,N_7494);
and U10308 (N_10308,N_7759,N_8280);
nor U10309 (N_10309,N_6611,N_6834);
nand U10310 (N_10310,N_7982,N_7067);
nand U10311 (N_10311,N_7329,N_8983);
xnor U10312 (N_10312,N_6442,N_7629);
nand U10313 (N_10313,N_8032,N_6771);
or U10314 (N_10314,N_7029,N_8182);
and U10315 (N_10315,N_7187,N_6330);
xnor U10316 (N_10316,N_6652,N_8308);
nor U10317 (N_10317,N_8433,N_8718);
nor U10318 (N_10318,N_8944,N_8283);
and U10319 (N_10319,N_6797,N_6934);
and U10320 (N_10320,N_6000,N_8153);
nor U10321 (N_10321,N_7795,N_7387);
nand U10322 (N_10322,N_8920,N_8498);
and U10323 (N_10323,N_6794,N_7937);
or U10324 (N_10324,N_7352,N_7553);
or U10325 (N_10325,N_6889,N_8146);
nand U10326 (N_10326,N_8009,N_6141);
xor U10327 (N_10327,N_6455,N_8342);
nor U10328 (N_10328,N_6420,N_6725);
nor U10329 (N_10329,N_8339,N_8829);
or U10330 (N_10330,N_7074,N_7700);
and U10331 (N_10331,N_6871,N_7849);
nor U10332 (N_10332,N_6431,N_8888);
nor U10333 (N_10333,N_8601,N_7716);
xor U10334 (N_10334,N_8739,N_6729);
and U10335 (N_10335,N_8647,N_8195);
nor U10336 (N_10336,N_6914,N_7890);
nor U10337 (N_10337,N_6833,N_8837);
nor U10338 (N_10338,N_6467,N_8825);
nand U10339 (N_10339,N_7492,N_7472);
xor U10340 (N_10340,N_8965,N_7295);
nand U10341 (N_10341,N_7941,N_7328);
xnor U10342 (N_10342,N_8386,N_8745);
or U10343 (N_10343,N_7513,N_7607);
nand U10344 (N_10344,N_7648,N_7864);
nor U10345 (N_10345,N_7846,N_8292);
or U10346 (N_10346,N_8333,N_8416);
nor U10347 (N_10347,N_8008,N_7338);
nand U10348 (N_10348,N_7653,N_6064);
or U10349 (N_10349,N_8625,N_8638);
or U10350 (N_10350,N_8732,N_6507);
nand U10351 (N_10351,N_7244,N_7602);
nand U10352 (N_10352,N_7257,N_6931);
nand U10353 (N_10353,N_6025,N_8506);
or U10354 (N_10354,N_8933,N_7993);
nor U10355 (N_10355,N_6021,N_6654);
nand U10356 (N_10356,N_8541,N_8902);
or U10357 (N_10357,N_6605,N_7018);
and U10358 (N_10358,N_8073,N_8502);
nand U10359 (N_10359,N_6572,N_6444);
nor U10360 (N_10360,N_8485,N_6280);
nand U10361 (N_10361,N_8495,N_8620);
or U10362 (N_10362,N_6527,N_8593);
nand U10363 (N_10363,N_6502,N_8214);
xor U10364 (N_10364,N_7519,N_8600);
or U10365 (N_10365,N_8874,N_6108);
nor U10366 (N_10366,N_6414,N_7825);
xnor U10367 (N_10367,N_6471,N_7925);
nand U10368 (N_10368,N_8893,N_7450);
nor U10369 (N_10369,N_6908,N_6604);
and U10370 (N_10370,N_8189,N_6275);
xnor U10371 (N_10371,N_7498,N_7115);
nor U10372 (N_10372,N_8744,N_6989);
nand U10373 (N_10373,N_6724,N_7960);
nand U10374 (N_10374,N_8992,N_6869);
and U10375 (N_10375,N_7461,N_6535);
or U10376 (N_10376,N_7102,N_8697);
or U10377 (N_10377,N_8080,N_6737);
or U10378 (N_10378,N_8851,N_8118);
nor U10379 (N_10379,N_8344,N_6011);
nand U10380 (N_10380,N_6411,N_6688);
or U10381 (N_10381,N_6372,N_6588);
or U10382 (N_10382,N_7705,N_6186);
nor U10383 (N_10383,N_7810,N_6154);
nand U10384 (N_10384,N_6530,N_6660);
nand U10385 (N_10385,N_7170,N_6423);
nand U10386 (N_10386,N_8446,N_7598);
or U10387 (N_10387,N_8464,N_8675);
nand U10388 (N_10388,N_8724,N_7897);
nor U10389 (N_10389,N_7374,N_8136);
nor U10390 (N_10390,N_6666,N_8612);
nand U10391 (N_10391,N_7702,N_8998);
nor U10392 (N_10392,N_6213,N_8041);
or U10393 (N_10393,N_6817,N_8949);
xor U10394 (N_10394,N_8421,N_8385);
xnor U10395 (N_10395,N_6120,N_8069);
and U10396 (N_10396,N_7844,N_8583);
nand U10397 (N_10397,N_8656,N_8470);
or U10398 (N_10398,N_6670,N_6562);
and U10399 (N_10399,N_6146,N_7205);
xor U10400 (N_10400,N_7286,N_6123);
and U10401 (N_10401,N_7688,N_6056);
or U10402 (N_10402,N_8454,N_8178);
nand U10403 (N_10403,N_7345,N_8091);
and U10404 (N_10404,N_7905,N_8728);
nand U10405 (N_10405,N_7775,N_7092);
or U10406 (N_10406,N_8487,N_8116);
and U10407 (N_10407,N_7354,N_8223);
nand U10408 (N_10408,N_6598,N_7335);
xor U10409 (N_10409,N_6257,N_8014);
nand U10410 (N_10410,N_8525,N_8667);
or U10411 (N_10411,N_8299,N_8546);
and U10412 (N_10412,N_8185,N_7518);
nand U10413 (N_10413,N_6839,N_8355);
and U10414 (N_10414,N_6665,N_8871);
and U10415 (N_10415,N_8700,N_7339);
nand U10416 (N_10416,N_7869,N_7512);
and U10417 (N_10417,N_7437,N_7068);
or U10418 (N_10418,N_7545,N_6597);
and U10419 (N_10419,N_6031,N_6140);
and U10420 (N_10420,N_7963,N_6321);
and U10421 (N_10421,N_8402,N_7003);
or U10422 (N_10422,N_7641,N_8192);
nand U10423 (N_10423,N_8679,N_6179);
nand U10424 (N_10424,N_7898,N_6437);
nand U10425 (N_10425,N_7291,N_8215);
nand U10426 (N_10426,N_7486,N_6114);
nor U10427 (N_10427,N_6310,N_8232);
xor U10428 (N_10428,N_8673,N_8461);
nand U10429 (N_10429,N_7647,N_8444);
nand U10430 (N_10430,N_7296,N_8966);
or U10431 (N_10431,N_6812,N_6366);
and U10432 (N_10432,N_7221,N_8353);
nor U10433 (N_10433,N_7779,N_6077);
or U10434 (N_10434,N_7733,N_7417);
nand U10435 (N_10435,N_6778,N_7432);
nor U10436 (N_10436,N_7052,N_8201);
nor U10437 (N_10437,N_8613,N_7236);
or U10438 (N_10438,N_6776,N_7416);
and U10439 (N_10439,N_6489,N_8838);
nor U10440 (N_10440,N_8329,N_6548);
nand U10441 (N_10441,N_8343,N_8588);
and U10442 (N_10442,N_8218,N_7574);
and U10443 (N_10443,N_7645,N_8240);
nor U10444 (N_10444,N_7539,N_7935);
nor U10445 (N_10445,N_8493,N_7573);
and U10446 (N_10446,N_6900,N_7109);
or U10447 (N_10447,N_8271,N_8695);
nor U10448 (N_10448,N_6882,N_6613);
xor U10449 (N_10449,N_7623,N_8503);
and U10450 (N_10450,N_7781,N_7600);
nand U10451 (N_10451,N_7145,N_8938);
nand U10452 (N_10452,N_6447,N_6607);
nor U10453 (N_10453,N_7243,N_8853);
nor U10454 (N_10454,N_8730,N_8774);
nand U10455 (N_10455,N_8545,N_8494);
and U10456 (N_10456,N_6966,N_8361);
and U10457 (N_10457,N_8518,N_6167);
nand U10458 (N_10458,N_8358,N_8326);
or U10459 (N_10459,N_8328,N_8501);
nor U10460 (N_10460,N_7403,N_8121);
and U10461 (N_10461,N_8363,N_7817);
xnor U10462 (N_10462,N_7634,N_8095);
nor U10463 (N_10463,N_7511,N_6161);
nor U10464 (N_10464,N_8316,N_7307);
or U10465 (N_10465,N_7618,N_8347);
and U10466 (N_10466,N_8930,N_6957);
nor U10467 (N_10467,N_6202,N_7621);
xnor U10468 (N_10468,N_6260,N_6888);
and U10469 (N_10469,N_7393,N_8989);
or U10470 (N_10470,N_6509,N_6440);
or U10471 (N_10471,N_8042,N_7514);
nand U10472 (N_10472,N_6748,N_7725);
nand U10473 (N_10473,N_8879,N_8826);
nand U10474 (N_10474,N_6255,N_7384);
nor U10475 (N_10475,N_7165,N_6684);
nor U10476 (N_10476,N_6759,N_8959);
nor U10477 (N_10477,N_6641,N_8352);
or U10478 (N_10478,N_6115,N_8286);
nor U10479 (N_10479,N_8964,N_6168);
xnor U10480 (N_10480,N_7266,N_6456);
nor U10481 (N_10481,N_7605,N_7816);
xnor U10482 (N_10482,N_7790,N_8754);
and U10483 (N_10483,N_7320,N_6661);
nor U10484 (N_10484,N_7942,N_6201);
or U10485 (N_10485,N_6541,N_7060);
and U10486 (N_10486,N_6307,N_6594);
nand U10487 (N_10487,N_7516,N_6536);
xnor U10488 (N_10488,N_8167,N_8689);
nor U10489 (N_10489,N_7906,N_6758);
nand U10490 (N_10490,N_8478,N_6832);
nand U10491 (N_10491,N_6802,N_8925);
xor U10492 (N_10492,N_7305,N_7661);
or U10493 (N_10493,N_8969,N_8383);
or U10494 (N_10494,N_6004,N_8649);
or U10495 (N_10495,N_8242,N_7850);
or U10496 (N_10496,N_8540,N_8068);
and U10497 (N_10497,N_6499,N_6258);
nand U10498 (N_10498,N_6311,N_8982);
or U10499 (N_10499,N_6073,N_6294);
or U10500 (N_10500,N_8164,N_8500);
nand U10501 (N_10501,N_7785,N_8921);
xor U10502 (N_10502,N_6751,N_6041);
nand U10503 (N_10503,N_6289,N_6677);
nand U10504 (N_10504,N_6368,N_6933);
or U10505 (N_10505,N_6203,N_8035);
xor U10506 (N_10506,N_7522,N_8984);
nand U10507 (N_10507,N_8999,N_6613);
or U10508 (N_10508,N_7622,N_7914);
xnor U10509 (N_10509,N_7890,N_6716);
and U10510 (N_10510,N_8778,N_7323);
or U10511 (N_10511,N_7847,N_8937);
and U10512 (N_10512,N_7583,N_7198);
nand U10513 (N_10513,N_6887,N_8606);
or U10514 (N_10514,N_7014,N_7552);
nor U10515 (N_10515,N_7165,N_8525);
xor U10516 (N_10516,N_6713,N_7376);
or U10517 (N_10517,N_7138,N_7757);
xnor U10518 (N_10518,N_7961,N_8986);
nand U10519 (N_10519,N_6502,N_7428);
nand U10520 (N_10520,N_7741,N_7226);
or U10521 (N_10521,N_6407,N_7957);
or U10522 (N_10522,N_6890,N_8201);
and U10523 (N_10523,N_7340,N_7208);
and U10524 (N_10524,N_6179,N_7280);
nand U10525 (N_10525,N_8343,N_6165);
xor U10526 (N_10526,N_7514,N_7874);
or U10527 (N_10527,N_6888,N_6735);
nand U10528 (N_10528,N_6398,N_8934);
nand U10529 (N_10529,N_6777,N_6684);
and U10530 (N_10530,N_7076,N_6652);
nor U10531 (N_10531,N_6619,N_6697);
and U10532 (N_10532,N_6725,N_6017);
xor U10533 (N_10533,N_6009,N_7387);
nor U10534 (N_10534,N_8198,N_6468);
or U10535 (N_10535,N_8178,N_6426);
nor U10536 (N_10536,N_8605,N_6096);
and U10537 (N_10537,N_6955,N_7711);
nor U10538 (N_10538,N_8583,N_6303);
or U10539 (N_10539,N_6261,N_8247);
or U10540 (N_10540,N_6556,N_7195);
nor U10541 (N_10541,N_8307,N_6771);
nand U10542 (N_10542,N_7005,N_8279);
or U10543 (N_10543,N_7275,N_8881);
nand U10544 (N_10544,N_6295,N_8301);
xnor U10545 (N_10545,N_7228,N_8572);
nand U10546 (N_10546,N_6920,N_7991);
nor U10547 (N_10547,N_7490,N_7080);
nand U10548 (N_10548,N_6258,N_7865);
nand U10549 (N_10549,N_6900,N_7668);
nand U10550 (N_10550,N_6058,N_8267);
or U10551 (N_10551,N_6858,N_8893);
nand U10552 (N_10552,N_8292,N_7445);
or U10553 (N_10553,N_6642,N_7104);
and U10554 (N_10554,N_8016,N_7648);
and U10555 (N_10555,N_6706,N_8651);
or U10556 (N_10556,N_6968,N_6934);
nor U10557 (N_10557,N_7649,N_7297);
nand U10558 (N_10558,N_7616,N_8074);
or U10559 (N_10559,N_6040,N_8722);
and U10560 (N_10560,N_7143,N_7253);
nand U10561 (N_10561,N_8179,N_6967);
or U10562 (N_10562,N_7440,N_8808);
nand U10563 (N_10563,N_8477,N_8347);
nand U10564 (N_10564,N_7763,N_8662);
or U10565 (N_10565,N_7476,N_7714);
nor U10566 (N_10566,N_6180,N_6936);
xor U10567 (N_10567,N_8584,N_7919);
nor U10568 (N_10568,N_7690,N_8612);
nand U10569 (N_10569,N_8580,N_6290);
or U10570 (N_10570,N_8369,N_8663);
nand U10571 (N_10571,N_8697,N_8794);
nand U10572 (N_10572,N_6616,N_8706);
nor U10573 (N_10573,N_7493,N_7253);
or U10574 (N_10574,N_6445,N_8091);
and U10575 (N_10575,N_7418,N_6098);
or U10576 (N_10576,N_8172,N_7462);
or U10577 (N_10577,N_8005,N_6913);
or U10578 (N_10578,N_6703,N_7288);
or U10579 (N_10579,N_6107,N_8554);
and U10580 (N_10580,N_7876,N_7608);
and U10581 (N_10581,N_8298,N_8645);
nor U10582 (N_10582,N_8339,N_7582);
xnor U10583 (N_10583,N_6996,N_7989);
and U10584 (N_10584,N_6754,N_7090);
nand U10585 (N_10585,N_6576,N_7508);
and U10586 (N_10586,N_7009,N_6736);
and U10587 (N_10587,N_7964,N_8493);
or U10588 (N_10588,N_8205,N_6833);
xor U10589 (N_10589,N_8489,N_6975);
nor U10590 (N_10590,N_6856,N_7716);
nor U10591 (N_10591,N_8026,N_6539);
and U10592 (N_10592,N_6537,N_8226);
nand U10593 (N_10593,N_7375,N_6319);
or U10594 (N_10594,N_7125,N_8755);
or U10595 (N_10595,N_7391,N_7408);
or U10596 (N_10596,N_8320,N_7978);
or U10597 (N_10597,N_8203,N_6236);
xnor U10598 (N_10598,N_7754,N_8666);
or U10599 (N_10599,N_7355,N_7961);
xnor U10600 (N_10600,N_6400,N_7678);
or U10601 (N_10601,N_7855,N_8809);
xor U10602 (N_10602,N_6125,N_8490);
nand U10603 (N_10603,N_7648,N_8029);
nor U10604 (N_10604,N_8422,N_8205);
or U10605 (N_10605,N_8441,N_6352);
or U10606 (N_10606,N_8687,N_7722);
nand U10607 (N_10607,N_8206,N_8312);
and U10608 (N_10608,N_7903,N_8492);
xnor U10609 (N_10609,N_8515,N_7169);
or U10610 (N_10610,N_6686,N_8226);
nand U10611 (N_10611,N_8753,N_6591);
xnor U10612 (N_10612,N_6903,N_8163);
nand U10613 (N_10613,N_8908,N_6305);
nor U10614 (N_10614,N_7571,N_6681);
and U10615 (N_10615,N_6169,N_7309);
and U10616 (N_10616,N_8725,N_8480);
or U10617 (N_10617,N_6310,N_6381);
or U10618 (N_10618,N_6908,N_8074);
nand U10619 (N_10619,N_7160,N_6832);
and U10620 (N_10620,N_8709,N_8949);
and U10621 (N_10621,N_8527,N_8685);
nand U10622 (N_10622,N_7969,N_7856);
or U10623 (N_10623,N_6986,N_6673);
nor U10624 (N_10624,N_8868,N_8045);
and U10625 (N_10625,N_6476,N_7021);
nor U10626 (N_10626,N_7333,N_8505);
nand U10627 (N_10627,N_7338,N_8277);
or U10628 (N_10628,N_8510,N_7486);
or U10629 (N_10629,N_7618,N_8254);
or U10630 (N_10630,N_8520,N_6323);
and U10631 (N_10631,N_8299,N_8767);
and U10632 (N_10632,N_7110,N_6264);
nand U10633 (N_10633,N_6263,N_8163);
xnor U10634 (N_10634,N_8860,N_8204);
and U10635 (N_10635,N_6969,N_8194);
or U10636 (N_10636,N_8772,N_6385);
and U10637 (N_10637,N_6802,N_8701);
or U10638 (N_10638,N_6121,N_6398);
xor U10639 (N_10639,N_7633,N_7017);
or U10640 (N_10640,N_8558,N_8423);
nor U10641 (N_10641,N_7001,N_8373);
xnor U10642 (N_10642,N_6304,N_7324);
nor U10643 (N_10643,N_7477,N_6879);
xnor U10644 (N_10644,N_8005,N_6379);
nand U10645 (N_10645,N_7159,N_7914);
or U10646 (N_10646,N_6966,N_8319);
xor U10647 (N_10647,N_8802,N_6338);
and U10648 (N_10648,N_6481,N_7982);
or U10649 (N_10649,N_8274,N_6294);
or U10650 (N_10650,N_6121,N_6426);
nor U10651 (N_10651,N_6338,N_6596);
and U10652 (N_10652,N_6948,N_7682);
and U10653 (N_10653,N_6984,N_8185);
nor U10654 (N_10654,N_8915,N_6560);
nor U10655 (N_10655,N_8233,N_6860);
or U10656 (N_10656,N_8004,N_6968);
xor U10657 (N_10657,N_7823,N_6006);
nor U10658 (N_10658,N_7402,N_7946);
or U10659 (N_10659,N_8029,N_6866);
or U10660 (N_10660,N_7583,N_8167);
nor U10661 (N_10661,N_7893,N_7849);
nor U10662 (N_10662,N_7972,N_8766);
nor U10663 (N_10663,N_6118,N_7832);
nand U10664 (N_10664,N_7440,N_6310);
and U10665 (N_10665,N_8546,N_6781);
nand U10666 (N_10666,N_8634,N_7949);
xor U10667 (N_10667,N_8380,N_7507);
and U10668 (N_10668,N_6860,N_7848);
and U10669 (N_10669,N_8594,N_6856);
or U10670 (N_10670,N_8557,N_7322);
nand U10671 (N_10671,N_7151,N_7803);
nand U10672 (N_10672,N_7416,N_7925);
nand U10673 (N_10673,N_7377,N_6747);
and U10674 (N_10674,N_6521,N_8558);
and U10675 (N_10675,N_8005,N_6124);
nor U10676 (N_10676,N_8805,N_6291);
and U10677 (N_10677,N_6363,N_8517);
and U10678 (N_10678,N_8350,N_6477);
and U10679 (N_10679,N_6772,N_8282);
nor U10680 (N_10680,N_6420,N_7176);
xnor U10681 (N_10681,N_6656,N_7022);
nor U10682 (N_10682,N_7077,N_6494);
nand U10683 (N_10683,N_6795,N_8067);
or U10684 (N_10684,N_7929,N_6113);
nor U10685 (N_10685,N_8072,N_7156);
nor U10686 (N_10686,N_6212,N_7738);
nor U10687 (N_10687,N_8578,N_6651);
nand U10688 (N_10688,N_6474,N_8390);
or U10689 (N_10689,N_8053,N_7876);
nand U10690 (N_10690,N_7803,N_8801);
and U10691 (N_10691,N_6070,N_7545);
and U10692 (N_10692,N_8049,N_7089);
nand U10693 (N_10693,N_8880,N_8040);
or U10694 (N_10694,N_7988,N_8987);
nor U10695 (N_10695,N_8012,N_8142);
or U10696 (N_10696,N_6211,N_7583);
or U10697 (N_10697,N_6933,N_6031);
nor U10698 (N_10698,N_8143,N_8479);
nand U10699 (N_10699,N_7313,N_6264);
and U10700 (N_10700,N_6440,N_7930);
or U10701 (N_10701,N_7707,N_7951);
or U10702 (N_10702,N_8627,N_8717);
nand U10703 (N_10703,N_8228,N_6063);
nor U10704 (N_10704,N_6476,N_6959);
nand U10705 (N_10705,N_7786,N_6232);
nor U10706 (N_10706,N_8609,N_8144);
or U10707 (N_10707,N_7079,N_8957);
nand U10708 (N_10708,N_8357,N_6825);
or U10709 (N_10709,N_7424,N_6262);
or U10710 (N_10710,N_8147,N_8052);
or U10711 (N_10711,N_8399,N_6015);
nor U10712 (N_10712,N_6188,N_6263);
nand U10713 (N_10713,N_6230,N_6930);
or U10714 (N_10714,N_8979,N_7231);
nand U10715 (N_10715,N_8725,N_8236);
nor U10716 (N_10716,N_8811,N_8196);
and U10717 (N_10717,N_7121,N_8426);
and U10718 (N_10718,N_6100,N_7475);
nand U10719 (N_10719,N_6205,N_8253);
or U10720 (N_10720,N_8155,N_8256);
or U10721 (N_10721,N_7174,N_7351);
nand U10722 (N_10722,N_7025,N_6624);
and U10723 (N_10723,N_7281,N_8063);
nor U10724 (N_10724,N_6636,N_7133);
or U10725 (N_10725,N_7757,N_8740);
or U10726 (N_10726,N_6637,N_7259);
nand U10727 (N_10727,N_8234,N_8483);
nor U10728 (N_10728,N_6347,N_6720);
nor U10729 (N_10729,N_8202,N_8512);
and U10730 (N_10730,N_6623,N_6728);
and U10731 (N_10731,N_6876,N_7112);
nor U10732 (N_10732,N_8732,N_6938);
nor U10733 (N_10733,N_8936,N_6939);
nor U10734 (N_10734,N_6754,N_8496);
and U10735 (N_10735,N_7026,N_7664);
nand U10736 (N_10736,N_7316,N_7699);
xor U10737 (N_10737,N_7520,N_6653);
nand U10738 (N_10738,N_8990,N_6322);
or U10739 (N_10739,N_6747,N_8065);
nor U10740 (N_10740,N_7668,N_7730);
nand U10741 (N_10741,N_7488,N_7386);
and U10742 (N_10742,N_6082,N_6307);
nor U10743 (N_10743,N_6914,N_6037);
or U10744 (N_10744,N_7497,N_8829);
nand U10745 (N_10745,N_8737,N_7826);
nor U10746 (N_10746,N_8056,N_6335);
nand U10747 (N_10747,N_6302,N_6468);
nor U10748 (N_10748,N_7472,N_6866);
nor U10749 (N_10749,N_7266,N_8040);
xnor U10750 (N_10750,N_6659,N_8624);
xor U10751 (N_10751,N_8088,N_6840);
nor U10752 (N_10752,N_8346,N_7489);
nor U10753 (N_10753,N_8739,N_6982);
and U10754 (N_10754,N_7191,N_7483);
nand U10755 (N_10755,N_6181,N_8785);
xnor U10756 (N_10756,N_6469,N_6337);
xnor U10757 (N_10757,N_7163,N_6754);
and U10758 (N_10758,N_8995,N_6149);
or U10759 (N_10759,N_8796,N_7055);
and U10760 (N_10760,N_6183,N_7338);
and U10761 (N_10761,N_7400,N_8563);
nand U10762 (N_10762,N_8585,N_6042);
nand U10763 (N_10763,N_6351,N_8159);
nor U10764 (N_10764,N_7616,N_7638);
or U10765 (N_10765,N_6329,N_6306);
xnor U10766 (N_10766,N_6697,N_6233);
or U10767 (N_10767,N_8636,N_7422);
nor U10768 (N_10768,N_7873,N_6579);
nand U10769 (N_10769,N_6287,N_7279);
and U10770 (N_10770,N_7437,N_6580);
nand U10771 (N_10771,N_6771,N_7000);
nor U10772 (N_10772,N_6252,N_8089);
nand U10773 (N_10773,N_6130,N_6330);
and U10774 (N_10774,N_6748,N_7022);
and U10775 (N_10775,N_7884,N_7226);
or U10776 (N_10776,N_8118,N_7907);
or U10777 (N_10777,N_6021,N_7196);
nand U10778 (N_10778,N_6736,N_7193);
nand U10779 (N_10779,N_7968,N_8868);
xor U10780 (N_10780,N_6475,N_7669);
and U10781 (N_10781,N_6095,N_7819);
nand U10782 (N_10782,N_7534,N_8471);
or U10783 (N_10783,N_8916,N_8374);
nor U10784 (N_10784,N_8155,N_8338);
and U10785 (N_10785,N_7402,N_8632);
xor U10786 (N_10786,N_8228,N_7360);
or U10787 (N_10787,N_6288,N_7738);
or U10788 (N_10788,N_7467,N_8624);
nand U10789 (N_10789,N_6330,N_8517);
xor U10790 (N_10790,N_8306,N_6754);
or U10791 (N_10791,N_7186,N_8791);
xnor U10792 (N_10792,N_6935,N_6172);
nor U10793 (N_10793,N_7178,N_7637);
nor U10794 (N_10794,N_7650,N_7535);
nand U10795 (N_10795,N_7369,N_8107);
or U10796 (N_10796,N_8331,N_8622);
or U10797 (N_10797,N_8711,N_8732);
nand U10798 (N_10798,N_6534,N_6427);
nand U10799 (N_10799,N_7345,N_7052);
or U10800 (N_10800,N_6009,N_8806);
xor U10801 (N_10801,N_7564,N_8787);
and U10802 (N_10802,N_6587,N_8849);
and U10803 (N_10803,N_7505,N_7616);
or U10804 (N_10804,N_6859,N_8222);
nand U10805 (N_10805,N_8417,N_8988);
xnor U10806 (N_10806,N_6832,N_7253);
nor U10807 (N_10807,N_7612,N_6174);
or U10808 (N_10808,N_7838,N_8391);
nand U10809 (N_10809,N_7570,N_7471);
or U10810 (N_10810,N_6254,N_7616);
nand U10811 (N_10811,N_7933,N_6264);
nand U10812 (N_10812,N_8757,N_6046);
nand U10813 (N_10813,N_7332,N_8943);
and U10814 (N_10814,N_6736,N_6569);
nand U10815 (N_10815,N_6218,N_8426);
nand U10816 (N_10816,N_7130,N_8692);
and U10817 (N_10817,N_8260,N_8168);
xnor U10818 (N_10818,N_6447,N_8739);
nor U10819 (N_10819,N_6939,N_8654);
nand U10820 (N_10820,N_8423,N_8925);
nor U10821 (N_10821,N_7035,N_7538);
and U10822 (N_10822,N_7558,N_6383);
nand U10823 (N_10823,N_8222,N_6558);
nor U10824 (N_10824,N_8063,N_7289);
or U10825 (N_10825,N_8898,N_8509);
nor U10826 (N_10826,N_7887,N_8639);
and U10827 (N_10827,N_7993,N_7962);
or U10828 (N_10828,N_7808,N_8637);
nor U10829 (N_10829,N_8983,N_7302);
nand U10830 (N_10830,N_8304,N_7573);
nor U10831 (N_10831,N_7609,N_6671);
and U10832 (N_10832,N_8450,N_7563);
nor U10833 (N_10833,N_8218,N_8396);
nand U10834 (N_10834,N_8320,N_8671);
nand U10835 (N_10835,N_6737,N_6033);
nand U10836 (N_10836,N_6252,N_7227);
nand U10837 (N_10837,N_6190,N_7608);
nor U10838 (N_10838,N_6842,N_8777);
and U10839 (N_10839,N_6978,N_6188);
and U10840 (N_10840,N_8438,N_7974);
xnor U10841 (N_10841,N_6731,N_7424);
or U10842 (N_10842,N_8173,N_6505);
or U10843 (N_10843,N_6517,N_6619);
nor U10844 (N_10844,N_8448,N_7607);
or U10845 (N_10845,N_7542,N_8841);
xor U10846 (N_10846,N_6085,N_7716);
and U10847 (N_10847,N_6503,N_7558);
or U10848 (N_10848,N_8144,N_6364);
nand U10849 (N_10849,N_7351,N_6673);
nand U10850 (N_10850,N_6201,N_6711);
nand U10851 (N_10851,N_8606,N_7105);
and U10852 (N_10852,N_6828,N_6033);
or U10853 (N_10853,N_6382,N_8619);
nor U10854 (N_10854,N_6109,N_7881);
nor U10855 (N_10855,N_7067,N_6948);
nand U10856 (N_10856,N_7826,N_8817);
nor U10857 (N_10857,N_6794,N_7991);
and U10858 (N_10858,N_8865,N_8309);
or U10859 (N_10859,N_8329,N_8794);
or U10860 (N_10860,N_7480,N_6246);
xor U10861 (N_10861,N_8289,N_7659);
nand U10862 (N_10862,N_6876,N_6164);
or U10863 (N_10863,N_6969,N_6747);
or U10864 (N_10864,N_8196,N_8635);
nor U10865 (N_10865,N_8950,N_6210);
or U10866 (N_10866,N_8710,N_8773);
xor U10867 (N_10867,N_7513,N_7880);
nor U10868 (N_10868,N_7944,N_7994);
or U10869 (N_10869,N_7061,N_8924);
and U10870 (N_10870,N_8243,N_7838);
nand U10871 (N_10871,N_7022,N_6680);
and U10872 (N_10872,N_8639,N_8714);
xor U10873 (N_10873,N_8054,N_6895);
nor U10874 (N_10874,N_6359,N_6506);
nand U10875 (N_10875,N_6725,N_8311);
or U10876 (N_10876,N_6576,N_6598);
xor U10877 (N_10877,N_8510,N_8299);
nor U10878 (N_10878,N_6606,N_8704);
nor U10879 (N_10879,N_6801,N_7233);
nor U10880 (N_10880,N_8013,N_7122);
nor U10881 (N_10881,N_6992,N_6197);
and U10882 (N_10882,N_8037,N_8169);
and U10883 (N_10883,N_6995,N_7027);
xor U10884 (N_10884,N_7019,N_8223);
and U10885 (N_10885,N_8618,N_7838);
nor U10886 (N_10886,N_7734,N_6205);
nor U10887 (N_10887,N_8534,N_7327);
nand U10888 (N_10888,N_7093,N_8601);
or U10889 (N_10889,N_6631,N_7942);
or U10890 (N_10890,N_7789,N_8127);
xnor U10891 (N_10891,N_8866,N_7050);
nor U10892 (N_10892,N_8207,N_7370);
and U10893 (N_10893,N_7542,N_6157);
or U10894 (N_10894,N_7091,N_6581);
xor U10895 (N_10895,N_8104,N_8515);
nand U10896 (N_10896,N_6457,N_8585);
nor U10897 (N_10897,N_6871,N_8555);
and U10898 (N_10898,N_7399,N_7316);
or U10899 (N_10899,N_6267,N_6280);
nand U10900 (N_10900,N_8768,N_6000);
or U10901 (N_10901,N_6567,N_7735);
and U10902 (N_10902,N_8647,N_8260);
nand U10903 (N_10903,N_8361,N_7654);
nand U10904 (N_10904,N_8409,N_8929);
and U10905 (N_10905,N_8967,N_6857);
and U10906 (N_10906,N_6512,N_8881);
nand U10907 (N_10907,N_8771,N_7232);
or U10908 (N_10908,N_6663,N_8454);
xnor U10909 (N_10909,N_6608,N_6640);
or U10910 (N_10910,N_7064,N_6375);
nand U10911 (N_10911,N_8209,N_7394);
or U10912 (N_10912,N_7348,N_8944);
nor U10913 (N_10913,N_8545,N_8290);
and U10914 (N_10914,N_7823,N_8289);
or U10915 (N_10915,N_8456,N_7574);
nand U10916 (N_10916,N_6244,N_7813);
xnor U10917 (N_10917,N_8832,N_8543);
or U10918 (N_10918,N_6014,N_6635);
nor U10919 (N_10919,N_6464,N_6576);
nand U10920 (N_10920,N_7040,N_8507);
nand U10921 (N_10921,N_6992,N_6808);
or U10922 (N_10922,N_7909,N_7140);
xnor U10923 (N_10923,N_7686,N_7967);
or U10924 (N_10924,N_8887,N_7204);
nand U10925 (N_10925,N_6756,N_8930);
nor U10926 (N_10926,N_8358,N_7670);
or U10927 (N_10927,N_6575,N_8377);
nand U10928 (N_10928,N_8985,N_7243);
or U10929 (N_10929,N_8392,N_6521);
or U10930 (N_10930,N_7248,N_8951);
or U10931 (N_10931,N_8262,N_8854);
nor U10932 (N_10932,N_8560,N_7669);
nor U10933 (N_10933,N_7059,N_7581);
or U10934 (N_10934,N_8110,N_6506);
or U10935 (N_10935,N_7223,N_6456);
and U10936 (N_10936,N_7491,N_8594);
xnor U10937 (N_10937,N_6145,N_7303);
nor U10938 (N_10938,N_7317,N_7496);
and U10939 (N_10939,N_6417,N_8609);
nand U10940 (N_10940,N_7533,N_8256);
nand U10941 (N_10941,N_6911,N_7823);
or U10942 (N_10942,N_8955,N_7133);
and U10943 (N_10943,N_7823,N_7317);
or U10944 (N_10944,N_8202,N_6370);
nand U10945 (N_10945,N_6186,N_7029);
and U10946 (N_10946,N_6156,N_6201);
or U10947 (N_10947,N_6368,N_8724);
nor U10948 (N_10948,N_7875,N_7279);
and U10949 (N_10949,N_6170,N_8861);
nor U10950 (N_10950,N_7184,N_7752);
nor U10951 (N_10951,N_7976,N_8681);
or U10952 (N_10952,N_8570,N_8457);
or U10953 (N_10953,N_8633,N_6795);
nand U10954 (N_10954,N_8483,N_6549);
or U10955 (N_10955,N_7582,N_6516);
and U10956 (N_10956,N_6499,N_7167);
nand U10957 (N_10957,N_8309,N_7740);
nor U10958 (N_10958,N_8259,N_7728);
nor U10959 (N_10959,N_6191,N_6043);
and U10960 (N_10960,N_8774,N_6091);
and U10961 (N_10961,N_7921,N_7384);
or U10962 (N_10962,N_7184,N_6119);
nor U10963 (N_10963,N_6227,N_8767);
nand U10964 (N_10964,N_8321,N_8878);
or U10965 (N_10965,N_8062,N_7902);
nor U10966 (N_10966,N_8943,N_6310);
nor U10967 (N_10967,N_6385,N_6333);
nand U10968 (N_10968,N_7382,N_7423);
and U10969 (N_10969,N_8498,N_8836);
and U10970 (N_10970,N_8349,N_7136);
or U10971 (N_10971,N_6547,N_6842);
nor U10972 (N_10972,N_8507,N_7030);
or U10973 (N_10973,N_7471,N_6674);
nor U10974 (N_10974,N_8353,N_7812);
and U10975 (N_10975,N_8365,N_7704);
nand U10976 (N_10976,N_6354,N_7897);
or U10977 (N_10977,N_8979,N_8018);
nor U10978 (N_10978,N_6123,N_8005);
nor U10979 (N_10979,N_7242,N_6452);
or U10980 (N_10980,N_6981,N_6785);
and U10981 (N_10981,N_7125,N_6965);
or U10982 (N_10982,N_7800,N_8929);
nand U10983 (N_10983,N_6334,N_8333);
xnor U10984 (N_10984,N_7566,N_6717);
and U10985 (N_10985,N_7063,N_6333);
or U10986 (N_10986,N_6826,N_8375);
and U10987 (N_10987,N_8990,N_6328);
and U10988 (N_10988,N_7318,N_7825);
nand U10989 (N_10989,N_6039,N_8268);
or U10990 (N_10990,N_6041,N_8905);
and U10991 (N_10991,N_7784,N_7006);
and U10992 (N_10992,N_6885,N_7920);
or U10993 (N_10993,N_6018,N_7924);
or U10994 (N_10994,N_6029,N_8778);
xor U10995 (N_10995,N_8432,N_8369);
or U10996 (N_10996,N_6095,N_8693);
nand U10997 (N_10997,N_6773,N_8418);
nand U10998 (N_10998,N_7936,N_8309);
nor U10999 (N_10999,N_7164,N_6044);
nand U11000 (N_11000,N_7255,N_8689);
or U11001 (N_11001,N_8826,N_7606);
nand U11002 (N_11002,N_7071,N_8719);
or U11003 (N_11003,N_7157,N_7456);
nand U11004 (N_11004,N_7152,N_8186);
nor U11005 (N_11005,N_7441,N_6976);
nand U11006 (N_11006,N_7749,N_8704);
nor U11007 (N_11007,N_8094,N_7133);
and U11008 (N_11008,N_8544,N_7973);
or U11009 (N_11009,N_7502,N_7503);
xnor U11010 (N_11010,N_7956,N_6736);
nand U11011 (N_11011,N_7391,N_6930);
nor U11012 (N_11012,N_6493,N_7387);
xor U11013 (N_11013,N_6977,N_7721);
nor U11014 (N_11014,N_7469,N_6265);
nand U11015 (N_11015,N_7747,N_7270);
and U11016 (N_11016,N_6152,N_6558);
xor U11017 (N_11017,N_7763,N_7547);
or U11018 (N_11018,N_7776,N_7053);
or U11019 (N_11019,N_6214,N_7409);
nand U11020 (N_11020,N_6371,N_8502);
or U11021 (N_11021,N_6408,N_8918);
and U11022 (N_11022,N_7907,N_8267);
nor U11023 (N_11023,N_7528,N_6827);
and U11024 (N_11024,N_6220,N_6908);
xnor U11025 (N_11025,N_8528,N_8039);
and U11026 (N_11026,N_7646,N_8114);
or U11027 (N_11027,N_6808,N_6949);
or U11028 (N_11028,N_6033,N_8876);
and U11029 (N_11029,N_7895,N_6035);
and U11030 (N_11030,N_7277,N_6976);
and U11031 (N_11031,N_6951,N_8011);
or U11032 (N_11032,N_8891,N_6806);
nor U11033 (N_11033,N_7457,N_6303);
nand U11034 (N_11034,N_8584,N_8438);
and U11035 (N_11035,N_8679,N_8741);
nand U11036 (N_11036,N_6438,N_6412);
nand U11037 (N_11037,N_8449,N_6901);
nor U11038 (N_11038,N_6772,N_8325);
nor U11039 (N_11039,N_7653,N_8665);
or U11040 (N_11040,N_8724,N_7260);
and U11041 (N_11041,N_6607,N_7367);
nand U11042 (N_11042,N_8628,N_6055);
or U11043 (N_11043,N_7184,N_7960);
and U11044 (N_11044,N_8415,N_6025);
xnor U11045 (N_11045,N_8834,N_7539);
or U11046 (N_11046,N_6566,N_7862);
nand U11047 (N_11047,N_7866,N_6550);
and U11048 (N_11048,N_7831,N_8162);
and U11049 (N_11049,N_7825,N_7005);
and U11050 (N_11050,N_7926,N_6015);
or U11051 (N_11051,N_7698,N_8769);
and U11052 (N_11052,N_7260,N_7917);
and U11053 (N_11053,N_7832,N_6494);
or U11054 (N_11054,N_7776,N_7190);
nand U11055 (N_11055,N_7240,N_7336);
nand U11056 (N_11056,N_8325,N_6226);
nand U11057 (N_11057,N_7999,N_6269);
or U11058 (N_11058,N_7375,N_8236);
xor U11059 (N_11059,N_6042,N_7956);
nor U11060 (N_11060,N_8433,N_7093);
or U11061 (N_11061,N_7405,N_8742);
nor U11062 (N_11062,N_8527,N_8699);
nand U11063 (N_11063,N_7475,N_6238);
or U11064 (N_11064,N_8338,N_8492);
nor U11065 (N_11065,N_6696,N_8797);
nor U11066 (N_11066,N_6314,N_6748);
nand U11067 (N_11067,N_6343,N_7835);
nand U11068 (N_11068,N_6247,N_8069);
and U11069 (N_11069,N_7892,N_6729);
or U11070 (N_11070,N_8398,N_7271);
and U11071 (N_11071,N_6642,N_7860);
nand U11072 (N_11072,N_7026,N_6314);
nand U11073 (N_11073,N_7606,N_6239);
or U11074 (N_11074,N_7275,N_6469);
xor U11075 (N_11075,N_8861,N_6244);
and U11076 (N_11076,N_6063,N_8355);
nor U11077 (N_11077,N_7041,N_7494);
or U11078 (N_11078,N_6923,N_6575);
or U11079 (N_11079,N_8113,N_6760);
or U11080 (N_11080,N_6288,N_6009);
nand U11081 (N_11081,N_8315,N_7495);
nor U11082 (N_11082,N_7351,N_6945);
or U11083 (N_11083,N_8255,N_6940);
xor U11084 (N_11084,N_6737,N_6138);
nor U11085 (N_11085,N_7544,N_8231);
or U11086 (N_11086,N_6437,N_6131);
nor U11087 (N_11087,N_6116,N_8631);
xor U11088 (N_11088,N_7745,N_8968);
xor U11089 (N_11089,N_7078,N_7618);
and U11090 (N_11090,N_8869,N_6935);
and U11091 (N_11091,N_6578,N_7914);
or U11092 (N_11092,N_7041,N_7404);
xnor U11093 (N_11093,N_8083,N_7749);
or U11094 (N_11094,N_7660,N_6748);
and U11095 (N_11095,N_7439,N_7838);
or U11096 (N_11096,N_7041,N_8235);
and U11097 (N_11097,N_6714,N_7514);
nor U11098 (N_11098,N_8472,N_8858);
nor U11099 (N_11099,N_7759,N_7426);
and U11100 (N_11100,N_7364,N_6389);
nor U11101 (N_11101,N_6820,N_6057);
nand U11102 (N_11102,N_6092,N_8566);
nor U11103 (N_11103,N_6621,N_8602);
and U11104 (N_11104,N_8899,N_6915);
or U11105 (N_11105,N_8374,N_6296);
nand U11106 (N_11106,N_7454,N_7750);
nand U11107 (N_11107,N_7707,N_6147);
and U11108 (N_11108,N_6894,N_6692);
nand U11109 (N_11109,N_8103,N_6920);
or U11110 (N_11110,N_6185,N_8060);
and U11111 (N_11111,N_8799,N_6599);
or U11112 (N_11112,N_7935,N_6803);
and U11113 (N_11113,N_8046,N_7301);
and U11114 (N_11114,N_8156,N_6763);
xor U11115 (N_11115,N_6083,N_7792);
nor U11116 (N_11116,N_8314,N_6098);
or U11117 (N_11117,N_7868,N_8720);
nor U11118 (N_11118,N_7217,N_8549);
nor U11119 (N_11119,N_8631,N_6649);
nand U11120 (N_11120,N_6055,N_8244);
nand U11121 (N_11121,N_8748,N_6648);
nor U11122 (N_11122,N_8355,N_6123);
and U11123 (N_11123,N_6431,N_8056);
nor U11124 (N_11124,N_8170,N_6625);
or U11125 (N_11125,N_8880,N_7585);
and U11126 (N_11126,N_8097,N_6838);
xnor U11127 (N_11127,N_7377,N_7361);
and U11128 (N_11128,N_7611,N_6712);
nor U11129 (N_11129,N_7474,N_6696);
and U11130 (N_11130,N_7875,N_7263);
nand U11131 (N_11131,N_7498,N_6988);
and U11132 (N_11132,N_7687,N_6298);
nor U11133 (N_11133,N_7042,N_6389);
nor U11134 (N_11134,N_8967,N_6685);
and U11135 (N_11135,N_7285,N_6525);
nand U11136 (N_11136,N_7248,N_7146);
nand U11137 (N_11137,N_8703,N_8306);
and U11138 (N_11138,N_7033,N_6093);
nand U11139 (N_11139,N_8322,N_8128);
xnor U11140 (N_11140,N_6238,N_6137);
nand U11141 (N_11141,N_7550,N_7050);
or U11142 (N_11142,N_8622,N_8176);
and U11143 (N_11143,N_6592,N_7215);
nor U11144 (N_11144,N_7935,N_6812);
and U11145 (N_11145,N_8222,N_7749);
nand U11146 (N_11146,N_6723,N_7005);
nand U11147 (N_11147,N_8247,N_7333);
nor U11148 (N_11148,N_7126,N_8208);
and U11149 (N_11149,N_8821,N_6878);
or U11150 (N_11150,N_7927,N_6897);
nand U11151 (N_11151,N_8073,N_6031);
and U11152 (N_11152,N_7046,N_8842);
xnor U11153 (N_11153,N_7401,N_7141);
nor U11154 (N_11154,N_6938,N_7500);
or U11155 (N_11155,N_7968,N_7112);
nor U11156 (N_11156,N_7523,N_8341);
nor U11157 (N_11157,N_6975,N_6562);
nor U11158 (N_11158,N_8182,N_6943);
nor U11159 (N_11159,N_6657,N_6747);
or U11160 (N_11160,N_6939,N_6211);
nand U11161 (N_11161,N_7215,N_7066);
and U11162 (N_11162,N_6555,N_8492);
or U11163 (N_11163,N_8708,N_8045);
xnor U11164 (N_11164,N_8554,N_8215);
nor U11165 (N_11165,N_7699,N_7809);
nor U11166 (N_11166,N_8387,N_8152);
and U11167 (N_11167,N_8119,N_8251);
and U11168 (N_11168,N_6365,N_8974);
nand U11169 (N_11169,N_7235,N_7203);
nand U11170 (N_11170,N_6632,N_7610);
or U11171 (N_11171,N_6391,N_8382);
nand U11172 (N_11172,N_7885,N_8150);
nor U11173 (N_11173,N_6962,N_7548);
nand U11174 (N_11174,N_6800,N_7420);
xnor U11175 (N_11175,N_7711,N_8104);
nand U11176 (N_11176,N_6913,N_7513);
nor U11177 (N_11177,N_8238,N_6720);
and U11178 (N_11178,N_8240,N_6009);
nand U11179 (N_11179,N_7007,N_7174);
nand U11180 (N_11180,N_7337,N_8306);
nor U11181 (N_11181,N_7480,N_7725);
and U11182 (N_11182,N_8053,N_7866);
and U11183 (N_11183,N_6752,N_7492);
xor U11184 (N_11184,N_7971,N_6913);
xor U11185 (N_11185,N_7673,N_7583);
and U11186 (N_11186,N_8014,N_6772);
and U11187 (N_11187,N_7810,N_8770);
nor U11188 (N_11188,N_7010,N_6957);
nand U11189 (N_11189,N_6172,N_7178);
or U11190 (N_11190,N_6605,N_6872);
or U11191 (N_11191,N_8998,N_8394);
or U11192 (N_11192,N_7912,N_6542);
nand U11193 (N_11193,N_6032,N_7721);
nand U11194 (N_11194,N_7154,N_8310);
nand U11195 (N_11195,N_6222,N_6234);
and U11196 (N_11196,N_7178,N_6805);
nor U11197 (N_11197,N_7169,N_7228);
nor U11198 (N_11198,N_6382,N_7302);
nor U11199 (N_11199,N_7289,N_7438);
and U11200 (N_11200,N_6062,N_8918);
nand U11201 (N_11201,N_7078,N_8979);
and U11202 (N_11202,N_7881,N_6026);
or U11203 (N_11203,N_8371,N_7510);
nand U11204 (N_11204,N_8941,N_6391);
and U11205 (N_11205,N_7930,N_8913);
nand U11206 (N_11206,N_6577,N_6074);
nand U11207 (N_11207,N_7239,N_6220);
nor U11208 (N_11208,N_8812,N_8933);
nor U11209 (N_11209,N_8563,N_7858);
or U11210 (N_11210,N_8803,N_8516);
or U11211 (N_11211,N_7459,N_8783);
and U11212 (N_11212,N_7163,N_8352);
or U11213 (N_11213,N_8316,N_6934);
nor U11214 (N_11214,N_7168,N_8410);
or U11215 (N_11215,N_8617,N_8628);
nor U11216 (N_11216,N_7609,N_8352);
and U11217 (N_11217,N_8601,N_8243);
xor U11218 (N_11218,N_8037,N_8318);
nand U11219 (N_11219,N_6952,N_6315);
and U11220 (N_11220,N_7330,N_6660);
and U11221 (N_11221,N_8816,N_7307);
xnor U11222 (N_11222,N_7915,N_7163);
and U11223 (N_11223,N_6672,N_7778);
nor U11224 (N_11224,N_7088,N_7556);
xnor U11225 (N_11225,N_8140,N_6623);
nand U11226 (N_11226,N_7372,N_8337);
and U11227 (N_11227,N_6109,N_6613);
nor U11228 (N_11228,N_8179,N_7518);
nand U11229 (N_11229,N_6894,N_7141);
nor U11230 (N_11230,N_8989,N_6603);
xnor U11231 (N_11231,N_7075,N_7764);
nor U11232 (N_11232,N_8755,N_7659);
nor U11233 (N_11233,N_7738,N_8315);
and U11234 (N_11234,N_7227,N_6166);
xor U11235 (N_11235,N_7110,N_7737);
xnor U11236 (N_11236,N_8328,N_6630);
xnor U11237 (N_11237,N_6443,N_8798);
or U11238 (N_11238,N_7720,N_7200);
nor U11239 (N_11239,N_7620,N_8927);
nand U11240 (N_11240,N_6684,N_7709);
nand U11241 (N_11241,N_7127,N_6937);
or U11242 (N_11242,N_8155,N_7753);
or U11243 (N_11243,N_7073,N_7513);
or U11244 (N_11244,N_7936,N_7159);
nor U11245 (N_11245,N_6659,N_6840);
nor U11246 (N_11246,N_6189,N_6389);
xnor U11247 (N_11247,N_8516,N_8215);
or U11248 (N_11248,N_6095,N_6968);
and U11249 (N_11249,N_8847,N_8315);
nor U11250 (N_11250,N_7285,N_8663);
nand U11251 (N_11251,N_6013,N_8139);
nor U11252 (N_11252,N_6095,N_8103);
nand U11253 (N_11253,N_7190,N_7531);
nor U11254 (N_11254,N_8169,N_8893);
nor U11255 (N_11255,N_6572,N_6079);
nand U11256 (N_11256,N_7852,N_8934);
or U11257 (N_11257,N_6037,N_8686);
and U11258 (N_11258,N_8245,N_6739);
xnor U11259 (N_11259,N_8120,N_8049);
nor U11260 (N_11260,N_8450,N_8298);
nand U11261 (N_11261,N_7042,N_8972);
or U11262 (N_11262,N_8069,N_6607);
nor U11263 (N_11263,N_6543,N_6020);
nor U11264 (N_11264,N_8488,N_8487);
nor U11265 (N_11265,N_8102,N_6540);
and U11266 (N_11266,N_7339,N_7310);
and U11267 (N_11267,N_6719,N_6643);
and U11268 (N_11268,N_8770,N_6464);
or U11269 (N_11269,N_8941,N_8340);
nor U11270 (N_11270,N_6539,N_7976);
or U11271 (N_11271,N_7403,N_7119);
nor U11272 (N_11272,N_8236,N_7269);
or U11273 (N_11273,N_7113,N_8931);
nand U11274 (N_11274,N_6717,N_7636);
or U11275 (N_11275,N_8622,N_8518);
nand U11276 (N_11276,N_6952,N_8344);
or U11277 (N_11277,N_7514,N_6895);
and U11278 (N_11278,N_8645,N_7933);
and U11279 (N_11279,N_7510,N_7928);
or U11280 (N_11280,N_8803,N_6420);
or U11281 (N_11281,N_7596,N_7458);
and U11282 (N_11282,N_8703,N_8279);
nand U11283 (N_11283,N_8168,N_7726);
xor U11284 (N_11284,N_6538,N_6443);
or U11285 (N_11285,N_7032,N_6413);
nand U11286 (N_11286,N_7266,N_7941);
or U11287 (N_11287,N_7267,N_8358);
nor U11288 (N_11288,N_6330,N_7198);
and U11289 (N_11289,N_6359,N_6995);
nand U11290 (N_11290,N_6338,N_6859);
xor U11291 (N_11291,N_7852,N_7331);
nand U11292 (N_11292,N_8074,N_8753);
and U11293 (N_11293,N_8830,N_6393);
or U11294 (N_11294,N_7528,N_7934);
and U11295 (N_11295,N_6825,N_7000);
nand U11296 (N_11296,N_7654,N_7278);
xnor U11297 (N_11297,N_6293,N_6386);
and U11298 (N_11298,N_7669,N_6418);
and U11299 (N_11299,N_7897,N_7008);
or U11300 (N_11300,N_8265,N_7766);
nand U11301 (N_11301,N_8957,N_6557);
and U11302 (N_11302,N_7480,N_7790);
or U11303 (N_11303,N_7392,N_7739);
or U11304 (N_11304,N_8100,N_6422);
and U11305 (N_11305,N_8078,N_6114);
nor U11306 (N_11306,N_6882,N_6323);
or U11307 (N_11307,N_8712,N_8694);
or U11308 (N_11308,N_7874,N_6713);
and U11309 (N_11309,N_8555,N_8122);
xnor U11310 (N_11310,N_8046,N_7105);
or U11311 (N_11311,N_8823,N_6483);
or U11312 (N_11312,N_7280,N_6291);
nand U11313 (N_11313,N_7150,N_6222);
xnor U11314 (N_11314,N_7786,N_6356);
nand U11315 (N_11315,N_7213,N_7073);
or U11316 (N_11316,N_8924,N_8144);
xnor U11317 (N_11317,N_8505,N_8033);
xor U11318 (N_11318,N_7212,N_7488);
nand U11319 (N_11319,N_7538,N_8866);
and U11320 (N_11320,N_6477,N_8780);
nand U11321 (N_11321,N_8563,N_7081);
or U11322 (N_11322,N_7280,N_8996);
xor U11323 (N_11323,N_8763,N_6513);
and U11324 (N_11324,N_7465,N_7190);
nand U11325 (N_11325,N_8221,N_6571);
nor U11326 (N_11326,N_6802,N_7648);
nand U11327 (N_11327,N_8118,N_6679);
nand U11328 (N_11328,N_7799,N_7302);
nor U11329 (N_11329,N_8015,N_8376);
nand U11330 (N_11330,N_6344,N_6608);
nor U11331 (N_11331,N_6588,N_6152);
or U11332 (N_11332,N_8675,N_7413);
and U11333 (N_11333,N_7653,N_6111);
xnor U11334 (N_11334,N_6005,N_7751);
and U11335 (N_11335,N_6576,N_6757);
or U11336 (N_11336,N_8005,N_7956);
nor U11337 (N_11337,N_7381,N_6043);
xor U11338 (N_11338,N_8816,N_7857);
and U11339 (N_11339,N_7198,N_6959);
or U11340 (N_11340,N_8381,N_8092);
and U11341 (N_11341,N_8017,N_7028);
and U11342 (N_11342,N_6610,N_7090);
or U11343 (N_11343,N_7303,N_6873);
and U11344 (N_11344,N_7227,N_6408);
or U11345 (N_11345,N_7973,N_8779);
nor U11346 (N_11346,N_6986,N_6912);
xnor U11347 (N_11347,N_7914,N_8786);
nand U11348 (N_11348,N_6070,N_7034);
nand U11349 (N_11349,N_7160,N_8511);
and U11350 (N_11350,N_7969,N_8711);
nand U11351 (N_11351,N_6098,N_8019);
or U11352 (N_11352,N_6370,N_7067);
or U11353 (N_11353,N_6108,N_7108);
nand U11354 (N_11354,N_7696,N_8721);
xor U11355 (N_11355,N_6748,N_8582);
xnor U11356 (N_11356,N_6765,N_6790);
nor U11357 (N_11357,N_8517,N_7703);
or U11358 (N_11358,N_6377,N_6333);
nand U11359 (N_11359,N_8946,N_7461);
nand U11360 (N_11360,N_6703,N_6636);
nor U11361 (N_11361,N_7579,N_7738);
or U11362 (N_11362,N_6022,N_6522);
and U11363 (N_11363,N_7786,N_6405);
nor U11364 (N_11364,N_6347,N_6725);
or U11365 (N_11365,N_6859,N_7841);
nor U11366 (N_11366,N_7244,N_8880);
nor U11367 (N_11367,N_6309,N_7632);
nor U11368 (N_11368,N_6252,N_6747);
or U11369 (N_11369,N_8648,N_7639);
xnor U11370 (N_11370,N_6686,N_7586);
nor U11371 (N_11371,N_7987,N_6870);
nor U11372 (N_11372,N_7440,N_7369);
and U11373 (N_11373,N_6178,N_6254);
and U11374 (N_11374,N_8402,N_6871);
nand U11375 (N_11375,N_8343,N_8063);
and U11376 (N_11376,N_8119,N_7964);
nor U11377 (N_11377,N_7201,N_7927);
or U11378 (N_11378,N_7708,N_8760);
xor U11379 (N_11379,N_7765,N_6433);
nor U11380 (N_11380,N_6378,N_8910);
nor U11381 (N_11381,N_6627,N_7924);
nand U11382 (N_11382,N_7032,N_7457);
nor U11383 (N_11383,N_7464,N_6397);
nor U11384 (N_11384,N_8252,N_8330);
and U11385 (N_11385,N_6671,N_6257);
nor U11386 (N_11386,N_6839,N_6399);
nor U11387 (N_11387,N_7898,N_7402);
xor U11388 (N_11388,N_8522,N_6703);
and U11389 (N_11389,N_8793,N_6807);
nand U11390 (N_11390,N_6598,N_7247);
and U11391 (N_11391,N_6137,N_6027);
nor U11392 (N_11392,N_7738,N_6967);
nand U11393 (N_11393,N_8259,N_6346);
nand U11394 (N_11394,N_8135,N_6090);
and U11395 (N_11395,N_7461,N_8868);
or U11396 (N_11396,N_6394,N_7609);
nor U11397 (N_11397,N_8988,N_6270);
nand U11398 (N_11398,N_7405,N_6319);
nand U11399 (N_11399,N_8229,N_8455);
nor U11400 (N_11400,N_8817,N_8659);
and U11401 (N_11401,N_6058,N_8099);
and U11402 (N_11402,N_7620,N_6597);
nand U11403 (N_11403,N_6021,N_6794);
or U11404 (N_11404,N_6047,N_7005);
and U11405 (N_11405,N_6563,N_6342);
nor U11406 (N_11406,N_8681,N_7219);
and U11407 (N_11407,N_6071,N_6012);
nor U11408 (N_11408,N_6009,N_8232);
and U11409 (N_11409,N_6806,N_7058);
nand U11410 (N_11410,N_8040,N_6557);
and U11411 (N_11411,N_8918,N_8041);
nand U11412 (N_11412,N_6910,N_7038);
and U11413 (N_11413,N_6516,N_6649);
nor U11414 (N_11414,N_6672,N_8880);
and U11415 (N_11415,N_6489,N_8287);
and U11416 (N_11416,N_8399,N_7109);
or U11417 (N_11417,N_7337,N_7289);
or U11418 (N_11418,N_6325,N_6403);
or U11419 (N_11419,N_8370,N_6134);
nor U11420 (N_11420,N_8453,N_7231);
xnor U11421 (N_11421,N_8011,N_6920);
and U11422 (N_11422,N_6585,N_8019);
or U11423 (N_11423,N_7736,N_6048);
xnor U11424 (N_11424,N_8862,N_6291);
nor U11425 (N_11425,N_8701,N_6205);
or U11426 (N_11426,N_7643,N_8822);
nand U11427 (N_11427,N_6834,N_8548);
xor U11428 (N_11428,N_6807,N_8103);
xnor U11429 (N_11429,N_7211,N_7740);
and U11430 (N_11430,N_6434,N_8987);
nand U11431 (N_11431,N_6665,N_7618);
nor U11432 (N_11432,N_7232,N_7490);
or U11433 (N_11433,N_8783,N_7656);
nor U11434 (N_11434,N_8697,N_6289);
and U11435 (N_11435,N_7324,N_8573);
nand U11436 (N_11436,N_7477,N_6981);
and U11437 (N_11437,N_7715,N_6243);
nand U11438 (N_11438,N_7200,N_6505);
or U11439 (N_11439,N_8400,N_6216);
and U11440 (N_11440,N_8409,N_6462);
nand U11441 (N_11441,N_8930,N_6034);
nand U11442 (N_11442,N_7242,N_7947);
nand U11443 (N_11443,N_6465,N_6169);
nand U11444 (N_11444,N_6979,N_7757);
nor U11445 (N_11445,N_6439,N_6199);
and U11446 (N_11446,N_8722,N_7332);
and U11447 (N_11447,N_8404,N_6806);
or U11448 (N_11448,N_7964,N_8001);
or U11449 (N_11449,N_6692,N_7311);
nor U11450 (N_11450,N_6322,N_7549);
nand U11451 (N_11451,N_7654,N_8255);
and U11452 (N_11452,N_8199,N_6105);
and U11453 (N_11453,N_8419,N_7457);
nand U11454 (N_11454,N_8711,N_7687);
and U11455 (N_11455,N_7740,N_6572);
xnor U11456 (N_11456,N_6932,N_7550);
or U11457 (N_11457,N_8205,N_6810);
or U11458 (N_11458,N_6613,N_8088);
xnor U11459 (N_11459,N_6697,N_6388);
or U11460 (N_11460,N_7752,N_6242);
and U11461 (N_11461,N_7587,N_6516);
and U11462 (N_11462,N_6322,N_8355);
xnor U11463 (N_11463,N_6505,N_7032);
nor U11464 (N_11464,N_8071,N_7607);
nand U11465 (N_11465,N_7464,N_7476);
nor U11466 (N_11466,N_8901,N_6967);
nand U11467 (N_11467,N_8392,N_8542);
and U11468 (N_11468,N_7910,N_6277);
nand U11469 (N_11469,N_6095,N_8732);
and U11470 (N_11470,N_7132,N_8228);
or U11471 (N_11471,N_6973,N_8985);
nor U11472 (N_11472,N_6261,N_8224);
and U11473 (N_11473,N_8050,N_6125);
nor U11474 (N_11474,N_7410,N_8174);
or U11475 (N_11475,N_6099,N_6528);
nand U11476 (N_11476,N_6548,N_8460);
nand U11477 (N_11477,N_8642,N_8989);
nand U11478 (N_11478,N_8947,N_8787);
or U11479 (N_11479,N_7339,N_6138);
or U11480 (N_11480,N_6395,N_6400);
nor U11481 (N_11481,N_7502,N_6798);
xnor U11482 (N_11482,N_6075,N_8001);
and U11483 (N_11483,N_8215,N_8222);
and U11484 (N_11484,N_6676,N_8314);
nand U11485 (N_11485,N_6653,N_7726);
and U11486 (N_11486,N_6866,N_7288);
or U11487 (N_11487,N_7025,N_8910);
and U11488 (N_11488,N_6785,N_6792);
nand U11489 (N_11489,N_6008,N_8866);
nand U11490 (N_11490,N_7159,N_7376);
nor U11491 (N_11491,N_7353,N_7361);
and U11492 (N_11492,N_7796,N_7884);
xor U11493 (N_11493,N_7665,N_8682);
or U11494 (N_11494,N_7307,N_7039);
nor U11495 (N_11495,N_8415,N_8385);
nand U11496 (N_11496,N_7241,N_7004);
xor U11497 (N_11497,N_7385,N_7570);
and U11498 (N_11498,N_7917,N_7183);
nor U11499 (N_11499,N_7442,N_7669);
and U11500 (N_11500,N_6964,N_6290);
or U11501 (N_11501,N_7962,N_6070);
xnor U11502 (N_11502,N_8874,N_7429);
nand U11503 (N_11503,N_6383,N_8009);
nor U11504 (N_11504,N_6131,N_7712);
nor U11505 (N_11505,N_7049,N_6756);
nor U11506 (N_11506,N_8709,N_8995);
nand U11507 (N_11507,N_8647,N_7264);
or U11508 (N_11508,N_6098,N_7129);
nor U11509 (N_11509,N_7946,N_6616);
nor U11510 (N_11510,N_7696,N_6145);
nor U11511 (N_11511,N_8769,N_7091);
or U11512 (N_11512,N_6172,N_7595);
nor U11513 (N_11513,N_6164,N_8227);
nor U11514 (N_11514,N_7533,N_7045);
and U11515 (N_11515,N_6053,N_7568);
or U11516 (N_11516,N_8206,N_8774);
or U11517 (N_11517,N_8186,N_6006);
nor U11518 (N_11518,N_7438,N_7750);
or U11519 (N_11519,N_8717,N_7667);
or U11520 (N_11520,N_6666,N_8774);
or U11521 (N_11521,N_8738,N_7388);
or U11522 (N_11522,N_8551,N_7251);
nand U11523 (N_11523,N_6075,N_7139);
and U11524 (N_11524,N_7505,N_7198);
nand U11525 (N_11525,N_6686,N_6380);
nand U11526 (N_11526,N_7650,N_6007);
and U11527 (N_11527,N_7459,N_7160);
nor U11528 (N_11528,N_7806,N_7575);
nor U11529 (N_11529,N_8170,N_6596);
nor U11530 (N_11530,N_6386,N_6144);
nor U11531 (N_11531,N_8206,N_6122);
nand U11532 (N_11532,N_8189,N_6990);
nand U11533 (N_11533,N_6791,N_7273);
or U11534 (N_11534,N_8567,N_6984);
and U11535 (N_11535,N_7279,N_7291);
nor U11536 (N_11536,N_7978,N_6779);
nor U11537 (N_11537,N_7785,N_6264);
xnor U11538 (N_11538,N_6524,N_6780);
and U11539 (N_11539,N_8162,N_8937);
or U11540 (N_11540,N_8195,N_6631);
nor U11541 (N_11541,N_7048,N_7403);
nor U11542 (N_11542,N_8914,N_7036);
or U11543 (N_11543,N_6955,N_8012);
nor U11544 (N_11544,N_8238,N_7498);
nor U11545 (N_11545,N_7826,N_6479);
xor U11546 (N_11546,N_7450,N_6549);
xnor U11547 (N_11547,N_6896,N_6207);
and U11548 (N_11548,N_6587,N_6633);
and U11549 (N_11549,N_8203,N_6556);
nand U11550 (N_11550,N_6099,N_6972);
nand U11551 (N_11551,N_6029,N_6067);
or U11552 (N_11552,N_6803,N_6971);
nand U11553 (N_11553,N_6313,N_7953);
or U11554 (N_11554,N_6618,N_7564);
and U11555 (N_11555,N_8256,N_7334);
or U11556 (N_11556,N_7076,N_6873);
and U11557 (N_11557,N_8873,N_8642);
or U11558 (N_11558,N_6367,N_8035);
nand U11559 (N_11559,N_6405,N_7114);
or U11560 (N_11560,N_7549,N_8825);
nand U11561 (N_11561,N_8742,N_7374);
nand U11562 (N_11562,N_7856,N_6676);
nand U11563 (N_11563,N_7350,N_8432);
nor U11564 (N_11564,N_6135,N_6741);
nand U11565 (N_11565,N_6547,N_8024);
nor U11566 (N_11566,N_8994,N_7036);
nor U11567 (N_11567,N_7208,N_7293);
nor U11568 (N_11568,N_7488,N_6982);
nor U11569 (N_11569,N_8640,N_8856);
nor U11570 (N_11570,N_6887,N_8386);
nor U11571 (N_11571,N_6416,N_7112);
nor U11572 (N_11572,N_6587,N_6008);
and U11573 (N_11573,N_8191,N_7732);
xnor U11574 (N_11574,N_7265,N_7506);
xnor U11575 (N_11575,N_6844,N_6885);
nand U11576 (N_11576,N_8073,N_7126);
and U11577 (N_11577,N_8211,N_8550);
nand U11578 (N_11578,N_6492,N_6253);
and U11579 (N_11579,N_8344,N_8351);
nor U11580 (N_11580,N_7059,N_8507);
nor U11581 (N_11581,N_6597,N_6034);
or U11582 (N_11582,N_7297,N_7598);
and U11583 (N_11583,N_6741,N_7661);
nor U11584 (N_11584,N_6853,N_7124);
and U11585 (N_11585,N_6399,N_8439);
or U11586 (N_11586,N_8600,N_8922);
xnor U11587 (N_11587,N_6586,N_6388);
and U11588 (N_11588,N_8799,N_7832);
or U11589 (N_11589,N_7668,N_7852);
and U11590 (N_11590,N_7566,N_7378);
nor U11591 (N_11591,N_8776,N_7422);
nand U11592 (N_11592,N_6970,N_6722);
nor U11593 (N_11593,N_6193,N_7153);
xnor U11594 (N_11594,N_6935,N_8520);
and U11595 (N_11595,N_8467,N_8594);
or U11596 (N_11596,N_8741,N_6736);
nor U11597 (N_11597,N_7808,N_8956);
xnor U11598 (N_11598,N_8007,N_8370);
nand U11599 (N_11599,N_8056,N_7725);
and U11600 (N_11600,N_8795,N_7942);
xor U11601 (N_11601,N_8246,N_8557);
nand U11602 (N_11602,N_8341,N_6910);
nor U11603 (N_11603,N_6706,N_6680);
nand U11604 (N_11604,N_7703,N_7901);
nor U11605 (N_11605,N_7042,N_6589);
nand U11606 (N_11606,N_6929,N_8821);
and U11607 (N_11607,N_7317,N_6519);
xnor U11608 (N_11608,N_6416,N_8452);
or U11609 (N_11609,N_8933,N_6795);
xor U11610 (N_11610,N_8392,N_7807);
nor U11611 (N_11611,N_7538,N_7353);
and U11612 (N_11612,N_6820,N_6408);
nor U11613 (N_11613,N_7804,N_6857);
and U11614 (N_11614,N_7858,N_7003);
or U11615 (N_11615,N_8643,N_8796);
nand U11616 (N_11616,N_6336,N_8290);
or U11617 (N_11617,N_8055,N_8698);
and U11618 (N_11618,N_6050,N_8328);
nand U11619 (N_11619,N_6695,N_7983);
nand U11620 (N_11620,N_8192,N_6520);
or U11621 (N_11621,N_6478,N_6714);
and U11622 (N_11622,N_6184,N_6419);
nand U11623 (N_11623,N_8561,N_7459);
nor U11624 (N_11624,N_6914,N_6224);
xnor U11625 (N_11625,N_7107,N_7226);
xor U11626 (N_11626,N_6354,N_8827);
nor U11627 (N_11627,N_6194,N_6144);
or U11628 (N_11628,N_7225,N_8657);
or U11629 (N_11629,N_6942,N_7960);
nor U11630 (N_11630,N_7397,N_7685);
and U11631 (N_11631,N_6413,N_8478);
and U11632 (N_11632,N_7801,N_8493);
nand U11633 (N_11633,N_8749,N_6305);
or U11634 (N_11634,N_7371,N_7244);
nand U11635 (N_11635,N_8177,N_6973);
nand U11636 (N_11636,N_6132,N_7435);
nand U11637 (N_11637,N_7040,N_6702);
and U11638 (N_11638,N_8296,N_8153);
nand U11639 (N_11639,N_7562,N_6793);
nand U11640 (N_11640,N_7069,N_8579);
nor U11641 (N_11641,N_6570,N_6364);
nor U11642 (N_11642,N_8865,N_8677);
and U11643 (N_11643,N_8722,N_7069);
nand U11644 (N_11644,N_6686,N_7456);
or U11645 (N_11645,N_8552,N_6096);
nor U11646 (N_11646,N_8361,N_7489);
and U11647 (N_11647,N_6448,N_7012);
and U11648 (N_11648,N_6707,N_6035);
nor U11649 (N_11649,N_7005,N_7411);
nand U11650 (N_11650,N_6002,N_6545);
and U11651 (N_11651,N_7922,N_6043);
xnor U11652 (N_11652,N_8905,N_8371);
nand U11653 (N_11653,N_8647,N_7164);
nor U11654 (N_11654,N_8784,N_6547);
nand U11655 (N_11655,N_8470,N_6727);
or U11656 (N_11656,N_7529,N_6718);
or U11657 (N_11657,N_6723,N_6424);
nand U11658 (N_11658,N_6844,N_6731);
nor U11659 (N_11659,N_6890,N_8627);
or U11660 (N_11660,N_6682,N_8229);
and U11661 (N_11661,N_6366,N_7586);
or U11662 (N_11662,N_7691,N_7851);
and U11663 (N_11663,N_8337,N_7580);
nand U11664 (N_11664,N_6957,N_8691);
and U11665 (N_11665,N_7024,N_6614);
nor U11666 (N_11666,N_8747,N_7185);
and U11667 (N_11667,N_8472,N_7667);
and U11668 (N_11668,N_7610,N_6950);
nor U11669 (N_11669,N_8038,N_8516);
or U11670 (N_11670,N_7725,N_6725);
xor U11671 (N_11671,N_6610,N_6746);
xor U11672 (N_11672,N_7401,N_6569);
nand U11673 (N_11673,N_6535,N_7760);
nand U11674 (N_11674,N_6304,N_7629);
nand U11675 (N_11675,N_6693,N_8588);
nand U11676 (N_11676,N_7583,N_6790);
nand U11677 (N_11677,N_6598,N_6348);
or U11678 (N_11678,N_7560,N_6371);
and U11679 (N_11679,N_7736,N_8294);
xnor U11680 (N_11680,N_8697,N_8095);
or U11681 (N_11681,N_8058,N_7788);
xnor U11682 (N_11682,N_6196,N_6885);
nor U11683 (N_11683,N_7811,N_6051);
and U11684 (N_11684,N_8195,N_6805);
nor U11685 (N_11685,N_7470,N_6692);
and U11686 (N_11686,N_8645,N_7081);
xor U11687 (N_11687,N_8021,N_6274);
and U11688 (N_11688,N_6344,N_6751);
and U11689 (N_11689,N_6031,N_8162);
nor U11690 (N_11690,N_7421,N_6148);
nand U11691 (N_11691,N_8074,N_7871);
nor U11692 (N_11692,N_8015,N_8389);
and U11693 (N_11693,N_7157,N_8940);
and U11694 (N_11694,N_6685,N_6729);
or U11695 (N_11695,N_8705,N_8350);
nand U11696 (N_11696,N_6990,N_8874);
and U11697 (N_11697,N_6429,N_7796);
nor U11698 (N_11698,N_7571,N_8287);
and U11699 (N_11699,N_6645,N_6726);
or U11700 (N_11700,N_8776,N_6206);
and U11701 (N_11701,N_6898,N_7510);
or U11702 (N_11702,N_6695,N_6250);
or U11703 (N_11703,N_6495,N_8140);
nor U11704 (N_11704,N_8187,N_8564);
and U11705 (N_11705,N_7063,N_7376);
and U11706 (N_11706,N_8215,N_6834);
or U11707 (N_11707,N_7508,N_8877);
and U11708 (N_11708,N_8367,N_7680);
xnor U11709 (N_11709,N_7027,N_6139);
and U11710 (N_11710,N_7463,N_8443);
nor U11711 (N_11711,N_7952,N_6482);
nor U11712 (N_11712,N_8108,N_6272);
xor U11713 (N_11713,N_7466,N_8410);
or U11714 (N_11714,N_8600,N_8071);
and U11715 (N_11715,N_8916,N_8232);
nand U11716 (N_11716,N_8594,N_8213);
nand U11717 (N_11717,N_8742,N_6415);
nor U11718 (N_11718,N_8744,N_7500);
and U11719 (N_11719,N_6204,N_8106);
and U11720 (N_11720,N_7953,N_6036);
and U11721 (N_11721,N_7794,N_8599);
nor U11722 (N_11722,N_7770,N_8183);
and U11723 (N_11723,N_7371,N_7460);
nand U11724 (N_11724,N_6363,N_7631);
or U11725 (N_11725,N_6376,N_6610);
and U11726 (N_11726,N_8086,N_7396);
nor U11727 (N_11727,N_8027,N_8751);
or U11728 (N_11728,N_6946,N_6542);
and U11729 (N_11729,N_6472,N_6715);
or U11730 (N_11730,N_8589,N_6184);
or U11731 (N_11731,N_7769,N_6684);
and U11732 (N_11732,N_7782,N_7760);
nand U11733 (N_11733,N_6705,N_7892);
or U11734 (N_11734,N_8865,N_6825);
nand U11735 (N_11735,N_8996,N_8851);
and U11736 (N_11736,N_7069,N_8860);
and U11737 (N_11737,N_8628,N_6608);
nand U11738 (N_11738,N_6138,N_7512);
or U11739 (N_11739,N_7383,N_7370);
nand U11740 (N_11740,N_6072,N_8301);
or U11741 (N_11741,N_7710,N_6877);
or U11742 (N_11742,N_6917,N_7575);
nor U11743 (N_11743,N_8047,N_8592);
nor U11744 (N_11744,N_7142,N_8064);
or U11745 (N_11745,N_6911,N_8608);
or U11746 (N_11746,N_8157,N_7732);
nand U11747 (N_11747,N_8920,N_7317);
nor U11748 (N_11748,N_8335,N_8686);
and U11749 (N_11749,N_6231,N_6344);
nor U11750 (N_11750,N_6246,N_8827);
or U11751 (N_11751,N_8561,N_8429);
nor U11752 (N_11752,N_8727,N_7829);
and U11753 (N_11753,N_8265,N_6095);
nor U11754 (N_11754,N_7727,N_6338);
nor U11755 (N_11755,N_7597,N_7137);
or U11756 (N_11756,N_7247,N_7784);
and U11757 (N_11757,N_8031,N_8897);
or U11758 (N_11758,N_8180,N_8216);
nor U11759 (N_11759,N_6213,N_6253);
and U11760 (N_11760,N_6083,N_8156);
or U11761 (N_11761,N_8050,N_8860);
and U11762 (N_11762,N_7628,N_7198);
xor U11763 (N_11763,N_8297,N_8887);
and U11764 (N_11764,N_7189,N_7568);
and U11765 (N_11765,N_6810,N_7088);
nand U11766 (N_11766,N_8530,N_7267);
nand U11767 (N_11767,N_8570,N_7900);
and U11768 (N_11768,N_6369,N_7138);
nand U11769 (N_11769,N_7179,N_6921);
and U11770 (N_11770,N_8626,N_7596);
and U11771 (N_11771,N_8312,N_7493);
nand U11772 (N_11772,N_6022,N_7517);
nor U11773 (N_11773,N_7604,N_6500);
or U11774 (N_11774,N_8702,N_6716);
and U11775 (N_11775,N_7710,N_8997);
or U11776 (N_11776,N_7627,N_7086);
and U11777 (N_11777,N_7472,N_6084);
xor U11778 (N_11778,N_6882,N_7520);
nor U11779 (N_11779,N_8007,N_8215);
nand U11780 (N_11780,N_8468,N_8516);
or U11781 (N_11781,N_6467,N_8558);
or U11782 (N_11782,N_8360,N_7557);
or U11783 (N_11783,N_6693,N_6586);
nand U11784 (N_11784,N_8271,N_6127);
or U11785 (N_11785,N_7848,N_6189);
or U11786 (N_11786,N_7446,N_7068);
or U11787 (N_11787,N_8118,N_8687);
and U11788 (N_11788,N_8624,N_6787);
or U11789 (N_11789,N_6170,N_6744);
xor U11790 (N_11790,N_7701,N_8033);
or U11791 (N_11791,N_8402,N_8309);
nor U11792 (N_11792,N_6242,N_7135);
or U11793 (N_11793,N_7311,N_6856);
nor U11794 (N_11794,N_7155,N_6571);
xnor U11795 (N_11795,N_8725,N_6857);
nand U11796 (N_11796,N_6679,N_7933);
or U11797 (N_11797,N_7468,N_6049);
or U11798 (N_11798,N_8368,N_6941);
nor U11799 (N_11799,N_7034,N_7342);
and U11800 (N_11800,N_7084,N_6664);
xnor U11801 (N_11801,N_6034,N_6084);
and U11802 (N_11802,N_8711,N_7704);
nor U11803 (N_11803,N_7240,N_7347);
and U11804 (N_11804,N_6244,N_6764);
or U11805 (N_11805,N_8952,N_7057);
or U11806 (N_11806,N_6450,N_7773);
and U11807 (N_11807,N_6988,N_8615);
or U11808 (N_11808,N_6925,N_8732);
nor U11809 (N_11809,N_6653,N_6258);
or U11810 (N_11810,N_7248,N_7228);
nor U11811 (N_11811,N_6087,N_7600);
nor U11812 (N_11812,N_7796,N_7961);
nor U11813 (N_11813,N_8509,N_6351);
or U11814 (N_11814,N_7938,N_8672);
and U11815 (N_11815,N_8598,N_8971);
nand U11816 (N_11816,N_6522,N_7177);
nand U11817 (N_11817,N_7003,N_6371);
xnor U11818 (N_11818,N_7965,N_7040);
nand U11819 (N_11819,N_6301,N_8313);
nor U11820 (N_11820,N_6096,N_6703);
or U11821 (N_11821,N_7979,N_8100);
nand U11822 (N_11822,N_7019,N_6574);
or U11823 (N_11823,N_6737,N_8796);
or U11824 (N_11824,N_8967,N_8259);
and U11825 (N_11825,N_7474,N_8586);
nand U11826 (N_11826,N_6777,N_6764);
and U11827 (N_11827,N_6176,N_8386);
or U11828 (N_11828,N_6434,N_7632);
and U11829 (N_11829,N_8348,N_8341);
or U11830 (N_11830,N_8722,N_6796);
or U11831 (N_11831,N_6817,N_7407);
and U11832 (N_11832,N_8258,N_8768);
and U11833 (N_11833,N_8612,N_8929);
and U11834 (N_11834,N_6512,N_7824);
nor U11835 (N_11835,N_8697,N_8015);
or U11836 (N_11836,N_6706,N_8249);
and U11837 (N_11837,N_7232,N_6424);
nand U11838 (N_11838,N_6190,N_7044);
or U11839 (N_11839,N_7849,N_6437);
nor U11840 (N_11840,N_6297,N_7946);
nand U11841 (N_11841,N_8909,N_8300);
nor U11842 (N_11842,N_6871,N_6472);
or U11843 (N_11843,N_8654,N_8284);
xor U11844 (N_11844,N_8774,N_8454);
nor U11845 (N_11845,N_7140,N_6062);
nor U11846 (N_11846,N_6023,N_7364);
nand U11847 (N_11847,N_8989,N_6292);
and U11848 (N_11848,N_6707,N_8242);
nor U11849 (N_11849,N_6286,N_8546);
nand U11850 (N_11850,N_7578,N_8408);
and U11851 (N_11851,N_7417,N_6383);
xor U11852 (N_11852,N_8865,N_6538);
nor U11853 (N_11853,N_6580,N_6337);
xnor U11854 (N_11854,N_6150,N_7780);
and U11855 (N_11855,N_7791,N_6463);
nor U11856 (N_11856,N_8700,N_7506);
xor U11857 (N_11857,N_6363,N_6372);
nand U11858 (N_11858,N_8062,N_7068);
xnor U11859 (N_11859,N_6759,N_6035);
xor U11860 (N_11860,N_6752,N_7588);
nor U11861 (N_11861,N_8116,N_7503);
nor U11862 (N_11862,N_7069,N_7468);
or U11863 (N_11863,N_8107,N_7592);
or U11864 (N_11864,N_8844,N_6526);
nand U11865 (N_11865,N_6090,N_7449);
xnor U11866 (N_11866,N_8132,N_8401);
and U11867 (N_11867,N_6954,N_8816);
nand U11868 (N_11868,N_7392,N_6598);
nand U11869 (N_11869,N_8076,N_6034);
nand U11870 (N_11870,N_8633,N_8019);
nor U11871 (N_11871,N_7775,N_8000);
nand U11872 (N_11872,N_7703,N_8222);
or U11873 (N_11873,N_7042,N_8824);
nand U11874 (N_11874,N_6527,N_8357);
xor U11875 (N_11875,N_6421,N_7912);
nor U11876 (N_11876,N_7416,N_8048);
xnor U11877 (N_11877,N_6216,N_8424);
nor U11878 (N_11878,N_7332,N_6024);
and U11879 (N_11879,N_6561,N_7498);
or U11880 (N_11880,N_8082,N_6795);
nand U11881 (N_11881,N_8275,N_6827);
nor U11882 (N_11882,N_6491,N_8621);
nand U11883 (N_11883,N_6245,N_6852);
or U11884 (N_11884,N_7404,N_7606);
xnor U11885 (N_11885,N_8222,N_6060);
and U11886 (N_11886,N_8199,N_7752);
and U11887 (N_11887,N_6893,N_8388);
nor U11888 (N_11888,N_6020,N_7345);
nor U11889 (N_11889,N_6706,N_8634);
nand U11890 (N_11890,N_6296,N_7727);
and U11891 (N_11891,N_8952,N_8168);
or U11892 (N_11892,N_8787,N_6583);
or U11893 (N_11893,N_6744,N_7163);
or U11894 (N_11894,N_7657,N_6466);
nor U11895 (N_11895,N_6311,N_8329);
xnor U11896 (N_11896,N_8235,N_8350);
nand U11897 (N_11897,N_7404,N_7111);
xor U11898 (N_11898,N_7244,N_8421);
and U11899 (N_11899,N_7411,N_8139);
or U11900 (N_11900,N_6277,N_8724);
nor U11901 (N_11901,N_7714,N_7305);
and U11902 (N_11902,N_8319,N_7468);
and U11903 (N_11903,N_6354,N_8940);
and U11904 (N_11904,N_7078,N_6280);
and U11905 (N_11905,N_7718,N_6656);
nand U11906 (N_11906,N_7797,N_8918);
xnor U11907 (N_11907,N_8582,N_7406);
and U11908 (N_11908,N_6906,N_8682);
or U11909 (N_11909,N_7810,N_7039);
or U11910 (N_11910,N_8811,N_6224);
nand U11911 (N_11911,N_6392,N_6072);
and U11912 (N_11912,N_6652,N_7747);
nand U11913 (N_11913,N_7729,N_8171);
nor U11914 (N_11914,N_6451,N_6624);
xnor U11915 (N_11915,N_7910,N_7171);
or U11916 (N_11916,N_8251,N_8040);
xnor U11917 (N_11917,N_8017,N_8811);
nand U11918 (N_11918,N_8628,N_6928);
nand U11919 (N_11919,N_8769,N_7732);
nand U11920 (N_11920,N_8653,N_8124);
nand U11921 (N_11921,N_6910,N_8947);
nor U11922 (N_11922,N_6405,N_8638);
nand U11923 (N_11923,N_7387,N_6838);
nand U11924 (N_11924,N_8256,N_8481);
or U11925 (N_11925,N_8406,N_6447);
nand U11926 (N_11926,N_6987,N_7647);
nor U11927 (N_11927,N_6970,N_8999);
nor U11928 (N_11928,N_7232,N_7367);
nor U11929 (N_11929,N_8811,N_7898);
and U11930 (N_11930,N_7317,N_8080);
or U11931 (N_11931,N_6737,N_8632);
or U11932 (N_11932,N_7339,N_7483);
or U11933 (N_11933,N_7796,N_6043);
nand U11934 (N_11934,N_6386,N_8809);
or U11935 (N_11935,N_8162,N_6170);
or U11936 (N_11936,N_7237,N_7579);
xnor U11937 (N_11937,N_6044,N_7981);
and U11938 (N_11938,N_7533,N_6700);
and U11939 (N_11939,N_6119,N_6602);
nor U11940 (N_11940,N_7528,N_8760);
nor U11941 (N_11941,N_8997,N_8474);
or U11942 (N_11942,N_6516,N_8036);
nand U11943 (N_11943,N_6635,N_6128);
nand U11944 (N_11944,N_8258,N_7264);
or U11945 (N_11945,N_8935,N_7614);
nand U11946 (N_11946,N_6101,N_7350);
nor U11947 (N_11947,N_7689,N_6008);
nand U11948 (N_11948,N_7447,N_7092);
nor U11949 (N_11949,N_6118,N_7342);
nand U11950 (N_11950,N_7523,N_6864);
nand U11951 (N_11951,N_7446,N_8938);
and U11952 (N_11952,N_6025,N_6803);
and U11953 (N_11953,N_7559,N_8137);
xnor U11954 (N_11954,N_6714,N_6390);
nand U11955 (N_11955,N_6050,N_7968);
or U11956 (N_11956,N_6821,N_8786);
xnor U11957 (N_11957,N_6569,N_6866);
nand U11958 (N_11958,N_6180,N_8979);
nor U11959 (N_11959,N_7527,N_7455);
nor U11960 (N_11960,N_7676,N_8526);
nor U11961 (N_11961,N_7962,N_7304);
or U11962 (N_11962,N_7712,N_7819);
or U11963 (N_11963,N_8114,N_8421);
or U11964 (N_11964,N_8617,N_6712);
or U11965 (N_11965,N_7924,N_7808);
and U11966 (N_11966,N_6257,N_7644);
or U11967 (N_11967,N_8052,N_6895);
and U11968 (N_11968,N_7153,N_7485);
nor U11969 (N_11969,N_6970,N_6156);
nand U11970 (N_11970,N_8297,N_8114);
nor U11971 (N_11971,N_6420,N_6324);
nand U11972 (N_11972,N_7620,N_7074);
nor U11973 (N_11973,N_6577,N_8709);
nor U11974 (N_11974,N_7192,N_6234);
and U11975 (N_11975,N_8089,N_8994);
and U11976 (N_11976,N_8233,N_8830);
nor U11977 (N_11977,N_7965,N_6573);
and U11978 (N_11978,N_6512,N_8574);
nor U11979 (N_11979,N_8981,N_6169);
and U11980 (N_11980,N_6452,N_6884);
and U11981 (N_11981,N_6893,N_7419);
nand U11982 (N_11982,N_8108,N_7069);
nand U11983 (N_11983,N_6606,N_7273);
or U11984 (N_11984,N_8879,N_7269);
and U11985 (N_11985,N_8705,N_6664);
xor U11986 (N_11986,N_6906,N_8860);
or U11987 (N_11987,N_8931,N_8226);
or U11988 (N_11988,N_8225,N_6712);
xnor U11989 (N_11989,N_7664,N_7514);
nand U11990 (N_11990,N_7017,N_6345);
nor U11991 (N_11991,N_7896,N_7138);
nand U11992 (N_11992,N_7696,N_8452);
nand U11993 (N_11993,N_8332,N_7416);
nor U11994 (N_11994,N_8788,N_7350);
or U11995 (N_11995,N_7028,N_7844);
or U11996 (N_11996,N_7122,N_6179);
nand U11997 (N_11997,N_7410,N_7498);
and U11998 (N_11998,N_8932,N_8792);
nor U11999 (N_11999,N_8130,N_7677);
or U12000 (N_12000,N_10808,N_11057);
nor U12001 (N_12001,N_11814,N_11031);
or U12002 (N_12002,N_10852,N_9882);
or U12003 (N_12003,N_10855,N_10011);
nor U12004 (N_12004,N_11952,N_10655);
nand U12005 (N_12005,N_9071,N_10724);
and U12006 (N_12006,N_10822,N_11136);
or U12007 (N_12007,N_11511,N_10305);
nand U12008 (N_12008,N_10609,N_9262);
nand U12009 (N_12009,N_11968,N_11769);
or U12010 (N_12010,N_10806,N_10232);
or U12011 (N_12011,N_11732,N_9860);
nor U12012 (N_12012,N_10897,N_9880);
nor U12013 (N_12013,N_11830,N_10255);
xor U12014 (N_12014,N_11274,N_11464);
nand U12015 (N_12015,N_9053,N_9593);
nand U12016 (N_12016,N_9640,N_10361);
nor U12017 (N_12017,N_10846,N_11240);
nand U12018 (N_12018,N_9259,N_10797);
nand U12019 (N_12019,N_9775,N_10439);
nor U12020 (N_12020,N_10621,N_11226);
nand U12021 (N_12021,N_9258,N_10673);
and U12022 (N_12022,N_10737,N_11495);
nand U12023 (N_12023,N_11823,N_9854);
xor U12024 (N_12024,N_9572,N_9715);
nor U12025 (N_12025,N_11561,N_9445);
nor U12026 (N_12026,N_11522,N_9012);
nor U12027 (N_12027,N_10747,N_9198);
nand U12028 (N_12028,N_9250,N_11775);
nor U12029 (N_12029,N_10519,N_11251);
nand U12030 (N_12030,N_9865,N_10710);
or U12031 (N_12031,N_10031,N_10311);
nor U12032 (N_12032,N_10900,N_9584);
nor U12033 (N_12033,N_10283,N_9828);
nor U12034 (N_12034,N_9273,N_11314);
nand U12035 (N_12035,N_11633,N_10496);
nand U12036 (N_12036,N_11883,N_9580);
nor U12037 (N_12037,N_9106,N_11677);
and U12038 (N_12038,N_9402,N_9834);
nand U12039 (N_12039,N_9404,N_11438);
nor U12040 (N_12040,N_10974,N_9490);
nand U12041 (N_12041,N_11743,N_9643);
and U12042 (N_12042,N_10869,N_11216);
nor U12043 (N_12043,N_11540,N_11075);
nor U12044 (N_12044,N_10201,N_10442);
xnor U12045 (N_12045,N_9306,N_11369);
nand U12046 (N_12046,N_10330,N_9059);
nand U12047 (N_12047,N_11704,N_10105);
nor U12048 (N_12048,N_10642,N_11861);
or U12049 (N_12049,N_9528,N_10707);
and U12050 (N_12050,N_11010,N_10340);
and U12051 (N_12051,N_9628,N_9808);
and U12052 (N_12052,N_10478,N_11526);
nor U12053 (N_12053,N_10677,N_10353);
and U12054 (N_12054,N_9830,N_10564);
nand U12055 (N_12055,N_9845,N_11407);
nand U12056 (N_12056,N_11552,N_10896);
or U12057 (N_12057,N_10607,N_9017);
or U12058 (N_12058,N_11070,N_9417);
nor U12059 (N_12059,N_11080,N_11686);
and U12060 (N_12060,N_10946,N_9850);
nor U12061 (N_12061,N_11019,N_9129);
or U12062 (N_12062,N_10804,N_11728);
nand U12063 (N_12063,N_9015,N_11772);
nand U12064 (N_12064,N_10202,N_11213);
nand U12065 (N_12065,N_10921,N_11364);
nor U12066 (N_12066,N_9183,N_10613);
nor U12067 (N_12067,N_9203,N_9214);
and U12068 (N_12068,N_11727,N_9756);
xor U12069 (N_12069,N_10187,N_11268);
nor U12070 (N_12070,N_11864,N_9669);
and U12071 (N_12071,N_10507,N_11544);
xnor U12072 (N_12072,N_10004,N_9261);
xor U12073 (N_12073,N_9900,N_9476);
or U12074 (N_12074,N_11286,N_11058);
or U12075 (N_12075,N_9581,N_10840);
and U12076 (N_12076,N_10799,N_9178);
and U12077 (N_12077,N_11731,N_11916);
nor U12078 (N_12078,N_10690,N_11917);
nand U12079 (N_12079,N_9181,N_9057);
nand U12080 (N_12080,N_11486,N_10835);
or U12081 (N_12081,N_9534,N_9690);
or U12082 (N_12082,N_10739,N_9758);
or U12083 (N_12083,N_10731,N_9994);
nand U12084 (N_12084,N_11073,N_11559);
xnor U12085 (N_12085,N_9199,N_10887);
xnor U12086 (N_12086,N_9356,N_11648);
and U12087 (N_12087,N_11386,N_10837);
and U12088 (N_12088,N_10604,N_10743);
nor U12089 (N_12089,N_9942,N_10438);
nor U12090 (N_12090,N_11037,N_11970);
and U12091 (N_12091,N_10375,N_10148);
nand U12092 (N_12092,N_9153,N_10476);
nand U12093 (N_12093,N_9403,N_9541);
nor U12094 (N_12094,N_9998,N_11718);
nand U12095 (N_12095,N_10220,N_11990);
nand U12096 (N_12096,N_9915,N_9531);
and U12097 (N_12097,N_10050,N_9410);
nand U12098 (N_12098,N_9216,N_10516);
xnor U12099 (N_12099,N_9038,N_10877);
nand U12100 (N_12100,N_9896,N_10864);
or U12101 (N_12101,N_9884,N_10112);
or U12102 (N_12102,N_11191,N_9113);
nor U12103 (N_12103,N_10640,N_9759);
or U12104 (N_12104,N_10966,N_11660);
nand U12105 (N_12105,N_10553,N_10858);
and U12106 (N_12106,N_9036,N_9163);
and U12107 (N_12107,N_11105,N_11340);
or U12108 (N_12108,N_9702,N_9603);
and U12109 (N_12109,N_9815,N_10461);
nand U12110 (N_12110,N_11184,N_11549);
nor U12111 (N_12111,N_9026,N_9475);
nor U12112 (N_12112,N_9268,N_9116);
nor U12113 (N_12113,N_9137,N_11889);
xnor U12114 (N_12114,N_9708,N_10007);
xnor U12115 (N_12115,N_11168,N_10230);
or U12116 (N_12116,N_9844,N_10178);
and U12117 (N_12117,N_10076,N_10001);
nor U12118 (N_12118,N_9256,N_9753);
or U12119 (N_12119,N_11420,N_10394);
or U12120 (N_12120,N_9792,N_9206);
and U12121 (N_12121,N_9033,N_10793);
and U12122 (N_12122,N_11385,N_11289);
and U12123 (N_12123,N_9633,N_10063);
nand U12124 (N_12124,N_9149,N_10458);
or U12125 (N_12125,N_11809,N_11798);
and U12126 (N_12126,N_10087,N_9656);
nand U12127 (N_12127,N_11455,N_11338);
or U12128 (N_12128,N_9504,N_11311);
xnor U12129 (N_12129,N_11187,N_9095);
and U12130 (N_12130,N_9427,N_11817);
nand U12131 (N_12131,N_10121,N_9468);
or U12132 (N_12132,N_11389,N_11611);
or U12133 (N_12133,N_9735,N_11770);
nand U12134 (N_12134,N_10693,N_9184);
nor U12135 (N_12135,N_9174,N_11481);
nor U12136 (N_12136,N_10585,N_11965);
and U12137 (N_12137,N_10164,N_10410);
xor U12138 (N_12138,N_11343,N_11974);
nand U12139 (N_12139,N_9147,N_11606);
or U12140 (N_12140,N_11713,N_10990);
xor U12141 (N_12141,N_10997,N_9619);
nor U12142 (N_12142,N_10061,N_10696);
nor U12143 (N_12143,N_9964,N_11394);
nand U12144 (N_12144,N_10853,N_10975);
and U12145 (N_12145,N_11285,N_11902);
nor U12146 (N_12146,N_11282,N_10815);
or U12147 (N_12147,N_9704,N_11129);
xor U12148 (N_12148,N_11962,N_9355);
nor U12149 (N_12149,N_9207,N_10297);
or U12150 (N_12150,N_11708,N_9368);
nand U12151 (N_12151,N_11987,N_11937);
nor U12152 (N_12152,N_9571,N_10985);
xnor U12153 (N_12153,N_10376,N_9500);
nand U12154 (N_12154,N_10615,N_11160);
xnor U12155 (N_12155,N_11147,N_10069);
or U12156 (N_12156,N_11752,N_9966);
nand U12157 (N_12157,N_9002,N_9725);
nor U12158 (N_12158,N_11118,N_11178);
nor U12159 (N_12159,N_10191,N_9892);
xnor U12160 (N_12160,N_11177,N_10278);
nor U12161 (N_12161,N_9151,N_10522);
nand U12162 (N_12162,N_10108,N_10198);
or U12163 (N_12163,N_11395,N_11207);
nor U12164 (N_12164,N_11113,N_9350);
or U12165 (N_12165,N_11875,N_10792);
nor U12166 (N_12166,N_11319,N_9709);
or U12167 (N_12167,N_10433,N_10650);
nand U12168 (N_12168,N_11847,N_9312);
xnor U12169 (N_12169,N_10116,N_9721);
or U12170 (N_12170,N_10943,N_10536);
nor U12171 (N_12171,N_9561,N_11026);
nand U12172 (N_12172,N_9888,N_9379);
nand U12173 (N_12173,N_10598,N_9622);
or U12174 (N_12174,N_10090,N_10068);
nand U12175 (N_12175,N_11567,N_11765);
and U12176 (N_12176,N_9343,N_10531);
nand U12177 (N_12177,N_10666,N_10923);
nor U12178 (N_12178,N_9952,N_11664);
and U12179 (N_12179,N_9659,N_9825);
nand U12180 (N_12180,N_9076,N_10322);
nand U12181 (N_12181,N_9511,N_10735);
xor U12182 (N_12182,N_9873,N_11796);
and U12183 (N_12183,N_10493,N_10711);
or U12184 (N_12184,N_11405,N_10557);
nand U12185 (N_12185,N_11346,N_10346);
xor U12186 (N_12186,N_10406,N_9540);
nand U12187 (N_12187,N_10929,N_9663);
or U12188 (N_12188,N_11739,N_10571);
nand U12189 (N_12189,N_10776,N_9069);
nor U12190 (N_12190,N_9270,N_11297);
nor U12191 (N_12191,N_10251,N_11662);
or U12192 (N_12192,N_10633,N_10427);
nand U12193 (N_12193,N_11276,N_9722);
nand U12194 (N_12194,N_10654,N_10794);
and U12195 (N_12195,N_9143,N_11487);
nand U12196 (N_12196,N_10714,N_9978);
nand U12197 (N_12197,N_11503,N_11201);
nand U12198 (N_12198,N_9887,N_11806);
nand U12199 (N_12199,N_10634,N_10931);
or U12200 (N_12200,N_9728,N_9448);
nand U12201 (N_12201,N_9227,N_10344);
nand U12202 (N_12202,N_10916,N_9255);
or U12203 (N_12203,N_10502,N_10168);
and U12204 (N_12204,N_11423,N_11306);
or U12205 (N_12205,N_10072,N_11292);
nand U12206 (N_12206,N_9464,N_10740);
nand U12207 (N_12207,N_11335,N_11563);
nor U12208 (N_12208,N_10398,N_11746);
or U12209 (N_12209,N_10382,N_9085);
or U12210 (N_12210,N_11398,N_11763);
or U12211 (N_12211,N_11195,N_9634);
nand U12212 (N_12212,N_10554,N_9245);
and U12213 (N_12213,N_10078,N_9586);
or U12214 (N_12214,N_10071,N_10608);
nand U12215 (N_12215,N_11930,N_11542);
or U12216 (N_12216,N_9326,N_10810);
xor U12217 (N_12217,N_11933,N_9107);
nand U12218 (N_12218,N_9956,N_11397);
and U12219 (N_12219,N_11500,N_10378);
or U12220 (N_12220,N_10142,N_11138);
nor U12221 (N_12221,N_10430,N_9311);
or U12222 (N_12222,N_11032,N_9347);
and U12223 (N_12223,N_10390,N_10092);
or U12224 (N_12224,N_11923,N_9724);
or U12225 (N_12225,N_9883,N_9167);
and U12226 (N_12226,N_9201,N_10345);
xnor U12227 (N_12227,N_9565,N_10998);
nor U12228 (N_12228,N_10592,N_11706);
or U12229 (N_12229,N_10863,N_9861);
and U12230 (N_12230,N_9526,N_9078);
nor U12231 (N_12231,N_10182,N_9631);
or U12232 (N_12232,N_9960,N_10367);
and U12233 (N_12233,N_10995,N_9931);
xor U12234 (N_12234,N_10880,N_10014);
or U12235 (N_12235,N_10448,N_9943);
and U12236 (N_12236,N_9569,N_10495);
or U12237 (N_12237,N_11801,N_9682);
xor U12238 (N_12238,N_11810,N_9176);
nand U12239 (N_12239,N_10039,N_11803);
nor U12240 (N_12240,N_9824,N_11279);
and U12241 (N_12241,N_11624,N_9717);
and U12242 (N_12242,N_11734,N_9155);
xor U12243 (N_12243,N_10996,N_10159);
xor U12244 (N_12244,N_11538,N_10002);
nand U12245 (N_12245,N_11625,N_10936);
nor U12246 (N_12246,N_11988,N_11961);
nand U12247 (N_12247,N_10280,N_11891);
or U12248 (N_12248,N_11610,N_10948);
nor U12249 (N_12249,N_11493,N_11152);
and U12250 (N_12250,N_11556,N_11555);
nand U12251 (N_12251,N_11034,N_10579);
and U12252 (N_12252,N_11926,N_11211);
nand U12253 (N_12253,N_9139,N_9662);
nand U12254 (N_12254,N_10184,N_10088);
nand U12255 (N_12255,N_10817,N_11277);
and U12256 (N_12256,N_11247,N_11403);
nor U12257 (N_12257,N_11218,N_11554);
and U12258 (N_12258,N_10415,N_11482);
and U12259 (N_12259,N_10578,N_10147);
xor U12260 (N_12260,N_10813,N_10140);
xnor U12261 (N_12261,N_10662,N_9380);
or U12262 (N_12262,N_10243,N_9388);
and U12263 (N_12263,N_9009,N_10027);
or U12264 (N_12264,N_9703,N_9301);
or U12265 (N_12265,N_11248,N_9186);
nor U12266 (N_12266,N_11776,N_9171);
or U12267 (N_12267,N_10132,N_10194);
and U12268 (N_12268,N_10901,N_9290);
or U12269 (N_12269,N_11782,N_11571);
or U12270 (N_12270,N_11509,N_10883);
nand U12271 (N_12271,N_11997,N_10567);
or U12272 (N_12272,N_10778,N_9164);
nor U12273 (N_12273,N_10755,N_11125);
nor U12274 (N_12274,N_11049,N_10447);
and U12275 (N_12275,N_11408,N_11504);
and U12276 (N_12276,N_11741,N_10919);
xor U12277 (N_12277,N_10606,N_9228);
or U12278 (N_12278,N_11264,N_11936);
nor U12279 (N_12279,N_10079,N_9805);
or U12280 (N_12280,N_11954,N_9160);
nor U12281 (N_12281,N_10138,N_11885);
nand U12282 (N_12282,N_10023,N_11558);
and U12283 (N_12283,N_11579,N_9816);
nor U12284 (N_12284,N_9418,N_11128);
or U12285 (N_12285,N_10774,N_10304);
and U12286 (N_12286,N_10437,N_10521);
nand U12287 (N_12287,N_10588,N_11827);
and U12288 (N_12288,N_9336,N_9332);
or U12289 (N_12289,N_11384,N_9800);
and U12290 (N_12290,N_11618,N_9434);
and U12291 (N_12291,N_11905,N_9415);
nor U12292 (N_12292,N_11716,N_11760);
nor U12293 (N_12293,N_11622,N_9063);
and U12294 (N_12294,N_11516,N_9393);
nand U12295 (N_12295,N_10440,N_9617);
nand U12296 (N_12296,N_11257,N_9197);
or U12297 (N_12297,N_10189,N_10547);
xor U12298 (N_12298,N_10208,N_10209);
and U12299 (N_12299,N_10844,N_11094);
nand U12300 (N_12300,N_11278,N_9140);
and U12301 (N_12301,N_9713,N_10722);
nand U12302 (N_12302,N_11171,N_10094);
nor U12303 (N_12303,N_11533,N_11904);
nor U12304 (N_12304,N_10485,N_11043);
and U12305 (N_12305,N_10572,N_10498);
and U12306 (N_12306,N_9831,N_9544);
and U12307 (N_12307,N_9676,N_11192);
nand U12308 (N_12308,N_9718,N_10221);
nand U12309 (N_12309,N_9909,N_11460);
and U12310 (N_12310,N_9419,N_10101);
and U12311 (N_12311,N_10653,N_11020);
nor U12312 (N_12312,N_9436,N_9723);
nand U12313 (N_12313,N_9179,N_9443);
or U12314 (N_12314,N_11698,N_11259);
xor U12315 (N_12315,N_11528,N_10399);
nor U12316 (N_12316,N_11273,N_9185);
or U12317 (N_12317,N_11644,N_10980);
nand U12318 (N_12318,N_10871,N_9649);
nor U12319 (N_12319,N_10161,N_10040);
and U12320 (N_12320,N_10436,N_11893);
or U12321 (N_12321,N_11015,N_11222);
xor U12322 (N_12322,N_9734,N_9019);
nor U12323 (N_12323,N_11508,N_10411);
and U12324 (N_12324,N_11252,N_9452);
and U12325 (N_12325,N_9212,N_10492);
nand U12326 (N_12326,N_10273,N_11215);
and U12327 (N_12327,N_9486,N_10867);
nand U12328 (N_12328,N_10669,N_9832);
and U12329 (N_12329,N_10645,N_10020);
and U12330 (N_12330,N_9670,N_10821);
and U12331 (N_12331,N_9247,N_9499);
xor U12332 (N_12332,N_11095,N_9519);
nor U12333 (N_12333,N_10825,N_10918);
nor U12334 (N_12334,N_9190,N_9503);
and U12335 (N_12335,N_11960,N_10300);
or U12336 (N_12336,N_10082,N_9736);
and U12337 (N_12337,N_9602,N_11059);
xnor U12338 (N_12338,N_10667,N_10573);
nor U12339 (N_12339,N_9836,N_11242);
nand U12340 (N_12340,N_9008,N_9077);
nand U12341 (N_12341,N_10888,N_11060);
or U12342 (N_12342,N_11159,N_10527);
or U12343 (N_12343,N_10917,N_11836);
nor U12344 (N_12344,N_11354,N_11229);
or U12345 (N_12345,N_9241,N_11869);
or U12346 (N_12346,N_9927,N_11149);
and U12347 (N_12347,N_10356,N_9322);
and U12348 (N_12348,N_11236,N_10876);
and U12349 (N_12349,N_11413,N_11468);
or U12350 (N_12350,N_9745,N_9283);
nand U12351 (N_12351,N_10380,N_11947);
nand U12352 (N_12352,N_9141,N_9447);
xnor U12353 (N_12353,N_9983,N_9922);
nor U12354 (N_12354,N_9570,N_10558);
or U12355 (N_12355,N_11725,N_10316);
xor U12356 (N_12356,N_10757,N_9778);
nand U12357 (N_12357,N_10246,N_10152);
or U12358 (N_12358,N_10351,N_9678);
nand U12359 (N_12359,N_10083,N_10017);
and U12360 (N_12360,N_11953,N_9453);
and U12361 (N_12361,N_9835,N_11726);
or U12362 (N_12362,N_11946,N_11223);
nor U12363 (N_12363,N_9296,N_10355);
or U12364 (N_12364,N_9848,N_9108);
nor U12365 (N_12365,N_11183,N_10686);
and U12366 (N_12366,N_9683,N_11999);
or U12367 (N_12367,N_9472,N_11233);
or U12368 (N_12368,N_9578,N_10474);
and U12369 (N_12369,N_11994,N_10704);
or U12370 (N_12370,N_11944,N_11519);
nand U12371 (N_12371,N_10234,N_9914);
nand U12372 (N_12372,N_11733,N_10548);
or U12373 (N_12373,N_11196,N_10036);
nor U12374 (N_12374,N_11269,N_11368);
nand U12375 (N_12375,N_11174,N_11860);
and U12376 (N_12376,N_10497,N_9408);
or U12377 (N_12377,N_11811,N_10773);
xor U12378 (N_12378,N_10983,N_11707);
nand U12379 (N_12379,N_11002,N_11890);
and U12380 (N_12380,N_9016,N_11584);
nand U12381 (N_12381,N_10056,N_9269);
and U12382 (N_12382,N_11913,N_9196);
nand U12383 (N_12383,N_9604,N_9665);
xor U12384 (N_12384,N_11941,N_10387);
nand U12385 (N_12385,N_10525,N_10894);
xnor U12386 (N_12386,N_11497,N_9849);
or U12387 (N_12387,N_11723,N_9599);
or U12388 (N_12388,N_9547,N_11022);
or U12389 (N_12389,N_9609,N_11047);
nand U12390 (N_12390,N_9958,N_10197);
or U12391 (N_12391,N_11646,N_10032);
and U12392 (N_12392,N_10245,N_10183);
xnor U12393 (N_12393,N_11266,N_9986);
xnor U12394 (N_12394,N_11449,N_11055);
or U12395 (N_12395,N_10679,N_10229);
nor U12396 (N_12396,N_10672,N_11599);
nor U12397 (N_12397,N_11454,N_10008);
and U12398 (N_12398,N_11690,N_11432);
nand U12399 (N_12399,N_11347,N_9652);
nand U12400 (N_12400,N_9871,N_9325);
or U12401 (N_12401,N_10293,N_11176);
nand U12402 (N_12402,N_10593,N_9248);
nor U12403 (N_12403,N_11761,N_11615);
or U12404 (N_12404,N_11906,N_9058);
and U12405 (N_12405,N_9866,N_11967);
and U12406 (N_12406,N_10620,N_10196);
or U12407 (N_12407,N_11682,N_9093);
nand U12408 (N_12408,N_11907,N_11474);
xnor U12409 (N_12409,N_10003,N_11357);
and U12410 (N_12410,N_9237,N_11383);
nor U12411 (N_12411,N_10911,N_9488);
and U12412 (N_12412,N_9507,N_10018);
and U12413 (N_12413,N_9737,N_9689);
xnor U12414 (N_12414,N_11576,N_9050);
nand U12415 (N_12415,N_9560,N_9902);
nand U12416 (N_12416,N_11607,N_10359);
or U12417 (N_12417,N_10253,N_9574);
nand U12418 (N_12418,N_10319,N_9889);
nand U12419 (N_12419,N_11463,N_10421);
or U12420 (N_12420,N_11832,N_9697);
nor U12421 (N_12421,N_11443,N_9329);
nand U12422 (N_12422,N_10590,N_11410);
or U12423 (N_12423,N_10185,N_11284);
nand U12424 (N_12424,N_11425,N_11310);
and U12425 (N_12425,N_10335,N_10716);
and U12426 (N_12426,N_11756,N_9298);
or U12427 (N_12427,N_9668,N_10016);
nor U12428 (N_12428,N_9299,N_10524);
nand U12429 (N_12429,N_10694,N_10156);
nand U12430 (N_12430,N_11843,N_11399);
xor U12431 (N_12431,N_10317,N_10227);
or U12432 (N_12432,N_10123,N_10816);
xor U12433 (N_12433,N_10733,N_11172);
nand U12434 (N_12434,N_11744,N_10104);
or U12435 (N_12435,N_9286,N_9360);
or U12436 (N_12436,N_11896,N_11067);
nand U12437 (N_12437,N_10641,N_10472);
and U12438 (N_12438,N_9099,N_9877);
and U12439 (N_12439,N_9980,N_11681);
or U12440 (N_12440,N_11689,N_9309);
and U12441 (N_12441,N_9707,N_10396);
nand U12442 (N_12442,N_11632,N_9799);
and U12443 (N_12443,N_11079,N_9246);
and U12444 (N_12444,N_11754,N_11370);
and U12445 (N_12445,N_10429,N_9542);
and U12446 (N_12446,N_10523,N_9772);
and U12447 (N_12447,N_10131,N_11507);
nand U12448 (N_12448,N_9949,N_9451);
nor U12449 (N_12449,N_9591,N_11780);
or U12450 (N_12450,N_10632,N_9905);
and U12451 (N_12451,N_9249,N_11390);
or U12452 (N_12452,N_11345,N_11378);
xnor U12453 (N_12453,N_9794,N_10179);
and U12454 (N_12454,N_10383,N_9991);
nor U12455 (N_12455,N_11181,N_11948);
and U12456 (N_12456,N_11773,N_11298);
xnor U12457 (N_12457,N_10586,N_11461);
xor U12458 (N_12458,N_10700,N_9316);
nand U12459 (N_12459,N_11759,N_11749);
and U12460 (N_12460,N_9134,N_9411);
nor U12461 (N_12461,N_9520,N_11626);
nor U12462 (N_12462,N_10687,N_11139);
or U12463 (N_12463,N_10265,N_11200);
or U12464 (N_12464,N_10796,N_9231);
nand U12465 (N_12465,N_11206,N_11560);
and U12466 (N_12466,N_11417,N_9293);
nand U12467 (N_12467,N_10093,N_11914);
and U12468 (N_12468,N_11392,N_10885);
and U12469 (N_12469,N_10260,N_9456);
nand U12470 (N_12470,N_10689,N_10569);
and U12471 (N_12471,N_10884,N_10708);
xor U12472 (N_12472,N_9750,N_11702);
or U12473 (N_12473,N_10832,N_11294);
or U12474 (N_12474,N_10765,N_10589);
or U12475 (N_12475,N_10624,N_10807);
and U12476 (N_12476,N_11230,N_10169);
nor U12477 (N_12477,N_9097,N_9789);
nand U12478 (N_12478,N_10528,N_9119);
nor U12479 (N_12479,N_10950,N_10659);
and U12480 (N_12480,N_11878,N_9467);
and U12481 (N_12481,N_11642,N_10057);
xor U12482 (N_12482,N_11793,N_9525);
nand U12483 (N_12483,N_9573,N_11376);
or U12484 (N_12484,N_11331,N_10803);
nor U12485 (N_12485,N_9615,N_11373);
xor U12486 (N_12486,N_11098,N_10978);
and U12487 (N_12487,N_11121,N_10879);
nand U12488 (N_12488,N_11078,N_9442);
nor U12489 (N_12489,N_9006,N_11107);
or U12490 (N_12490,N_9509,N_9474);
and U12491 (N_12491,N_10294,N_10172);
and U12492 (N_12492,N_9973,N_11865);
nor U12493 (N_12493,N_9688,N_11912);
and U12494 (N_12494,N_10904,N_11038);
or U12495 (N_12495,N_10418,N_9390);
nand U12496 (N_12496,N_10787,N_9345);
or U12497 (N_12497,N_9940,N_10186);
nand U12498 (N_12498,N_9564,N_10712);
nand U12499 (N_12499,N_10479,N_9660);
nor U12500 (N_12500,N_11938,N_11547);
nand U12501 (N_12501,N_11422,N_11643);
nand U12502 (N_12502,N_9202,N_11712);
xnor U12503 (N_12503,N_11748,N_11258);
nor U12504 (N_12504,N_9366,N_10318);
and U12505 (N_12505,N_10125,N_11472);
and U12506 (N_12506,N_9483,N_10504);
or U12507 (N_12507,N_10499,N_9135);
nor U12508 (N_12508,N_10199,N_9576);
nand U12509 (N_12509,N_9897,N_9876);
and U12510 (N_12510,N_10977,N_10828);
nor U12511 (N_12511,N_11777,N_10697);
nand U12512 (N_12512,N_9118,N_11785);
nand U12513 (N_12513,N_11097,N_10772);
or U12514 (N_12514,N_11868,N_10241);
or U12515 (N_12515,N_11220,N_9052);
or U12516 (N_12516,N_9802,N_9821);
or U12517 (N_12517,N_9933,N_11573);
xnor U12518 (N_12518,N_10959,N_10420);
and U12519 (N_12519,N_10055,N_11301);
xnor U12520 (N_12520,N_11989,N_9730);
nor U12521 (N_12521,N_9251,N_11597);
and U12522 (N_12522,N_11036,N_10738);
nand U12523 (N_12523,N_9305,N_11774);
nand U12524 (N_12524,N_10193,N_10428);
and U12525 (N_12525,N_11825,N_11006);
nor U12526 (N_12526,N_11028,N_10886);
and U12527 (N_12527,N_10575,N_11874);
and U12528 (N_12528,N_10944,N_11421);
nand U12529 (N_12529,N_10222,N_10514);
or U12530 (N_12530,N_9046,N_11525);
nand U12531 (N_12531,N_9597,N_11465);
nor U12532 (N_12532,N_11155,N_11456);
and U12533 (N_12533,N_9780,N_10922);
and U12534 (N_12534,N_10725,N_11452);
or U12535 (N_12535,N_9323,N_11871);
and U12536 (N_12536,N_9754,N_11023);
or U12537 (N_12537,N_9793,N_11521);
nand U12538 (N_12538,N_10584,N_11077);
xnor U12539 (N_12539,N_10798,N_10166);
nor U12540 (N_12540,N_10301,N_10644);
and U12541 (N_12541,N_9492,N_11908);
xor U12542 (N_12542,N_9522,N_10422);
nor U12543 (N_12543,N_11973,N_10129);
xnor U12544 (N_12544,N_11447,N_10216);
or U12545 (N_12545,N_9223,N_11033);
or U12546 (N_12546,N_11979,N_10377);
nor U12547 (N_12547,N_10635,N_11683);
nor U12548 (N_12548,N_9045,N_9813);
and U12549 (N_12549,N_11666,N_10336);
nor U12550 (N_12550,N_10425,N_11688);
nor U12551 (N_12551,N_9477,N_10533);
and U12552 (N_12552,N_9044,N_10818);
nor U12553 (N_12553,N_11480,N_10480);
or U12554 (N_12554,N_9030,N_11009);
or U12555 (N_12555,N_11543,N_11484);
nand U12556 (N_12556,N_10705,N_9755);
and U12557 (N_12557,N_9537,N_10664);
nand U12558 (N_12558,N_10307,N_9177);
nand U12559 (N_12559,N_9878,N_11362);
nor U12560 (N_12560,N_10518,N_11605);
and U12561 (N_12561,N_9867,N_11135);
nand U12562 (N_12562,N_10562,N_11835);
nand U12563 (N_12563,N_9369,N_11641);
nand U12564 (N_12564,N_11270,N_11123);
or U12565 (N_12565,N_9493,N_9658);
or U12566 (N_12566,N_11824,N_9685);
and U12567 (N_12567,N_11453,N_10254);
or U12568 (N_12568,N_10914,N_11530);
nand U12569 (N_12569,N_10468,N_9126);
and U12570 (N_12570,N_9224,N_11303);
nand U12571 (N_12571,N_11048,N_9075);
and U12572 (N_12572,N_9444,N_11478);
or U12573 (N_12573,N_11637,N_11720);
nor U12574 (N_12574,N_9625,N_11603);
and U12575 (N_12575,N_10790,N_9400);
and U12576 (N_12576,N_9079,N_9916);
and U12577 (N_12577,N_10403,N_11256);
or U12578 (N_12578,N_9105,N_10431);
nand U12579 (N_12579,N_10715,N_10482);
nor U12580 (N_12580,N_10648,N_11104);
nand U12581 (N_12581,N_9801,N_11355);
or U12582 (N_12582,N_9953,N_9773);
nand U12583 (N_12583,N_9068,N_9406);
or U12584 (N_12584,N_9766,N_9040);
nor U12585 (N_12585,N_11764,N_11700);
and U12586 (N_12586,N_10982,N_11379);
nand U12587 (N_12587,N_11431,N_9635);
xnor U12588 (N_12588,N_10252,N_10576);
nand U12589 (N_12589,N_10559,N_11789);
or U12590 (N_12590,N_11100,N_10006);
or U12591 (N_12591,N_11580,N_10839);
xor U12592 (N_12592,N_10702,N_9020);
nor U12593 (N_12593,N_11040,N_9005);
or U12594 (N_12594,N_10013,N_11583);
nor U12595 (N_12595,N_9837,N_10475);
and U12596 (N_12596,N_9967,N_10934);
and U12597 (N_12597,N_9340,N_11807);
xnor U12598 (N_12598,N_10158,N_10637);
and U12599 (N_12599,N_9985,N_11124);
nor U12600 (N_12600,N_11588,N_11828);
and U12601 (N_12601,N_9691,N_11513);
xnor U12602 (N_12602,N_11365,N_11175);
and U12603 (N_12603,N_11235,N_9606);
or U12604 (N_12604,N_10405,N_10683);
nor U12605 (N_12605,N_10848,N_10306);
or U12606 (N_12606,N_11352,N_9536);
and U12607 (N_12607,N_10473,N_9729);
nor U12608 (N_12608,N_10048,N_9950);
nand U12609 (N_12609,N_9822,N_11494);
or U12610 (N_12610,N_11550,N_11877);
nand U12611 (N_12611,N_9162,N_10960);
or U12612 (N_12612,N_9655,N_10099);
or U12613 (N_12613,N_9784,N_10126);
nor U12614 (N_12614,N_9731,N_11065);
or U12615 (N_12615,N_10021,N_10534);
and U12616 (N_12616,N_11388,N_10370);
and U12617 (N_12617,N_10270,N_9928);
nand U12618 (N_12618,N_9743,N_10477);
or U12619 (N_12619,N_10552,N_11173);
and U12620 (N_12620,N_10928,N_9412);
and U12621 (N_12621,N_11859,N_11185);
xor U12622 (N_12622,N_10895,N_10267);
nand U12623 (N_12623,N_9138,N_9761);
or U12624 (N_12624,N_9829,N_11645);
or U12625 (N_12625,N_11227,N_11411);
or U12626 (N_12626,N_10250,N_9487);
nor U12627 (N_12627,N_9626,N_10719);
and U12628 (N_12628,N_9485,N_10034);
and U12629 (N_12629,N_9727,N_10195);
nor U12630 (N_12630,N_9532,N_9292);
and U12631 (N_12631,N_10899,N_9502);
nand U12632 (N_12632,N_10540,N_10402);
nand U12633 (N_12633,N_10616,N_10713);
and U12634 (N_12634,N_10325,N_11344);
and U12635 (N_12635,N_10784,N_11265);
or U12636 (N_12636,N_10120,N_11071);
or U12637 (N_12637,N_10217,N_10652);
nand U12638 (N_12638,N_11332,N_10935);
and U12639 (N_12639,N_11161,N_10856);
nor U12640 (N_12640,N_9235,N_9747);
or U12641 (N_12641,N_9583,N_9891);
nand U12642 (N_12642,N_11483,N_10970);
nand U12643 (N_12643,N_11730,N_11490);
nand U12644 (N_12644,N_9239,N_10591);
nor U12645 (N_12645,N_10969,N_10460);
and U12646 (N_12646,N_11356,N_11924);
and U12647 (N_12647,N_10371,N_10058);
nand U12648 (N_12648,N_9568,N_9779);
and U12649 (N_12649,N_10012,N_10908);
nor U12650 (N_12650,N_10249,N_11360);
nor U12651 (N_12651,N_9620,N_9895);
nor U12652 (N_12652,N_9354,N_9338);
nor U12653 (N_12653,N_9995,N_11450);
nand U12654 (N_12654,N_10107,N_11131);
nor U12655 (N_12655,N_9204,N_10500);
nand U12656 (N_12656,N_10688,N_11092);
nand U12657 (N_12657,N_10862,N_11085);
or U12658 (N_12658,N_9131,N_10910);
nor U12659 (N_12659,N_11088,N_9518);
or U12660 (N_12660,N_10313,N_10085);
and U12661 (N_12661,N_9847,N_11241);
xnor U12662 (N_12662,N_10544,N_9387);
nor U12663 (N_12663,N_9996,N_11684);
and U12664 (N_12664,N_10647,N_9462);
and U12665 (N_12665,N_11382,N_11590);
or U12666 (N_12666,N_9701,N_11246);
and U12667 (N_12667,N_9760,N_9804);
nor U12668 (N_12668,N_9324,N_10758);
nor U12669 (N_12669,N_11245,N_9130);
nand U12670 (N_12670,N_10854,N_10729);
nor U12671 (N_12671,N_11087,N_11108);
or U12672 (N_12672,N_11485,N_9111);
or U12673 (N_12673,N_11302,N_10834);
or U12674 (N_12674,N_11562,N_10721);
xor U12675 (N_12675,N_10423,N_9263);
nor U12676 (N_12676,N_10113,N_10651);
or U12677 (N_12677,N_9820,N_10992);
nand U12678 (N_12678,N_10210,N_11722);
nand U12679 (N_12679,N_10981,N_9074);
nor U12680 (N_12680,N_10053,N_9607);
nand U12681 (N_12681,N_11661,N_11815);
or U12682 (N_12682,N_9230,N_11616);
nand U12683 (N_12683,N_10860,N_10341);
or U12684 (N_12684,N_11143,N_9875);
nor U12685 (N_12685,N_10565,N_10329);
nand U12686 (N_12686,N_10363,N_11565);
nand U12687 (N_12687,N_9070,N_10889);
nand U12688 (N_12688,N_11011,N_10117);
nor U12689 (N_12689,N_10045,N_9274);
and U12690 (N_12690,N_9460,N_10913);
and U12691 (N_12691,N_10111,N_9275);
xor U12692 (N_12692,N_9208,N_11694);
nor U12693 (N_12693,N_11329,N_9826);
or U12694 (N_12694,N_10947,N_9657);
nand U12695 (N_12695,N_10226,N_9929);
xor U12696 (N_12696,N_9321,N_11876);
and U12697 (N_12697,N_9358,N_10259);
nand U12698 (N_12698,N_9384,N_9563);
and U12699 (N_12699,N_9217,N_9279);
or U12700 (N_12700,N_10509,N_9254);
nor U12701 (N_12701,N_10211,N_10366);
nor U12702 (N_12702,N_9339,N_11054);
or U12703 (N_12703,N_11090,N_10751);
and U12704 (N_12704,N_11320,N_9304);
nand U12705 (N_12705,N_9439,N_11056);
nor U12706 (N_12706,N_10044,N_9240);
nand U12707 (N_12707,N_11167,N_9976);
xnor U12708 (N_12708,N_10391,N_9548);
or U12709 (N_12709,N_11813,N_11404);
nor U12710 (N_12710,N_11596,N_9797);
or U12711 (N_12711,N_10701,N_11029);
or U12712 (N_12712,N_9935,N_9109);
or U12713 (N_12713,N_10656,N_11654);
and U12714 (N_12714,N_11190,N_11679);
xnor U12715 (N_12715,N_9310,N_10176);
xnor U12716 (N_12716,N_9225,N_10955);
and U12717 (N_12717,N_9706,N_10503);
and U12718 (N_12718,N_9514,N_9552);
and U12719 (N_12719,N_10150,N_9535);
nor U12720 (N_12720,N_11995,N_9923);
nor U12721 (N_12721,N_9025,N_9021);
or U12722 (N_12722,N_10723,N_9749);
or U12723 (N_12723,N_10801,N_10354);
and U12724 (N_12724,N_9182,N_10443);
and U12725 (N_12725,N_10972,N_11884);
nor U12726 (N_12726,N_9945,N_10882);
or U12727 (N_12727,N_9638,N_9809);
nor U12728 (N_12728,N_11050,N_9925);
and U12729 (N_12729,N_10788,N_9232);
nand U12730 (N_12730,N_11154,N_9710);
or U12731 (N_12731,N_10225,N_11587);
nor U12732 (N_12732,N_10732,N_10459);
nor U12733 (N_12733,N_11581,N_10752);
or U12734 (N_12734,N_9067,N_9610);
xnor U12735 (N_12735,N_10276,N_11441);
and U12736 (N_12736,N_9977,N_11738);
and U12737 (N_12737,N_9466,N_10550);
or U12738 (N_12738,N_9315,N_11969);
xnor U12739 (N_12739,N_11134,N_9211);
xnor U12740 (N_12740,N_10360,N_11153);
nor U12741 (N_12741,N_9859,N_10035);
and U12742 (N_12742,N_10845,N_9297);
and U12743 (N_12743,N_10829,N_10115);
nor U12744 (N_12744,N_9303,N_11371);
or U12745 (N_12745,N_9313,N_10369);
nor U12746 (N_12746,N_9533,N_10568);
nor U12747 (N_12747,N_11076,N_9752);
nor U12748 (N_12748,N_9851,N_11204);
nor U12749 (N_12749,N_10236,N_9192);
xnor U12750 (N_12750,N_10597,N_11210);
or U12751 (N_12751,N_10781,N_9060);
nand U12752 (N_12752,N_11000,N_9327);
or U12753 (N_12753,N_9551,N_11313);
or U12754 (N_12754,N_10930,N_11863);
and U12755 (N_12755,N_11445,N_9788);
or U12756 (N_12756,N_10455,N_11524);
nand U12757 (N_12757,N_10906,N_10263);
xnor U12758 (N_12758,N_9605,N_10000);
and U12759 (N_12759,N_10905,N_9142);
and U12760 (N_12760,N_11669,N_11374);
nor U12761 (N_12761,N_9144,N_11950);
and U12762 (N_12762,N_10279,N_11024);
or U12763 (N_12763,N_10703,N_11021);
nor U12764 (N_12764,N_11670,N_11719);
nand U12765 (N_12765,N_11249,N_10205);
or U12766 (N_12766,N_10824,N_10891);
or U12767 (N_12767,N_9031,N_11359);
nand U12768 (N_12768,N_11695,N_11437);
or U12769 (N_12769,N_10795,N_10320);
and U12770 (N_12770,N_9763,N_11433);
or U12771 (N_12771,N_11870,N_9629);
nand U12772 (N_12772,N_10520,N_10529);
xnor U12773 (N_12773,N_11221,N_11091);
or U12774 (N_12774,N_9947,N_11459);
and U12775 (N_12775,N_11442,N_10999);
or U12776 (N_12776,N_9524,N_10097);
or U12777 (N_12777,N_9041,N_10971);
or U12778 (N_12778,N_11372,N_10691);
and U12779 (N_12779,N_10517,N_9919);
or U12780 (N_12780,N_10933,N_11663);
nand U12781 (N_12781,N_11735,N_10401);
or U12782 (N_12782,N_10699,N_10332);
and U12783 (N_12783,N_10450,N_10095);
and U12784 (N_12784,N_10051,N_10228);
nand U12785 (N_12785,N_11342,N_11959);
nand U12786 (N_12786,N_11272,N_9396);
nor U12787 (N_12787,N_9173,N_9422);
nor U12788 (N_12788,N_11505,N_11214);
nand U12789 (N_12789,N_11671,N_9621);
nand U12790 (N_12790,N_9014,N_11897);
nand U12791 (N_12791,N_11471,N_10661);
and U12792 (N_12792,N_11145,N_11820);
nand U12793 (N_12793,N_9446,N_9785);
or U12794 (N_12794,N_11971,N_9716);
nor U12795 (N_12795,N_9482,N_10820);
nor U12796 (N_12796,N_9963,N_9220);
or U12797 (N_12797,N_9553,N_11697);
or U12798 (N_12798,N_11012,N_10046);
nor U12799 (N_12799,N_9146,N_11578);
and U12800 (N_12800,N_11535,N_11647);
or U12801 (N_12801,N_11110,N_9630);
xnor U12802 (N_12802,N_9671,N_11797);
nand U12803 (N_12803,N_9122,N_9252);
and U12804 (N_12804,N_10766,N_9455);
nor U12805 (N_12805,N_11721,N_10266);
xnor U12806 (N_12806,N_10709,N_10312);
nand U12807 (N_12807,N_9767,N_9065);
nor U12808 (N_12808,N_9911,N_11955);
nor U12809 (N_12809,N_10486,N_11601);
nor U12810 (N_12810,N_10932,N_11652);
nor U12811 (N_12811,N_10494,N_10441);
nor U12812 (N_12812,N_9762,N_11387);
nand U12813 (N_12813,N_11658,N_10483);
and U12814 (N_12814,N_9971,N_10692);
or U12815 (N_12815,N_9280,N_10487);
and U12816 (N_12816,N_9817,N_9435);
and U12817 (N_12817,N_10466,N_9397);
nand U12818 (N_12818,N_9917,N_10649);
nand U12819 (N_12819,N_9974,N_11784);
or U12820 (N_12820,N_10133,N_11163);
nor U12821 (N_12821,N_10281,N_9972);
nor U12822 (N_12822,N_11699,N_9567);
nor U12823 (N_12823,N_10501,N_10764);
nor U12824 (N_12824,N_11881,N_10903);
nor U12825 (N_12825,N_11260,N_10264);
xnor U12826 (N_12826,N_10233,N_11348);
nand U12827 (N_12827,N_11322,N_11910);
nor U12828 (N_12828,N_9376,N_10838);
and U12829 (N_12829,N_10154,N_10812);
nor U12830 (N_12830,N_11539,N_11194);
nor U12831 (N_12831,N_9244,N_9372);
or U12832 (N_12832,N_11418,N_10392);
or U12833 (N_12833,N_9926,N_10993);
or U12834 (N_12834,N_11862,N_10949);
nand U12835 (N_12835,N_9295,N_9092);
and U12836 (N_12836,N_9786,N_11262);
nand U12837 (N_12837,N_11209,N_9698);
or U12838 (N_12838,N_9776,N_11768);
or U12839 (N_12839,N_9084,N_9238);
or U12840 (N_12840,N_10357,N_9064);
and U12841 (N_12841,N_11102,N_11546);
nand U12842 (N_12842,N_9011,N_9864);
nor U12843 (N_12843,N_9981,N_11617);
and U12844 (N_12844,N_9645,N_10098);
nor U12845 (N_12845,N_10358,N_10510);
nand U12846 (N_12846,N_9102,N_9700);
xnor U12847 (N_12847,N_10286,N_11203);
nand U12848 (N_12848,N_9159,N_9037);
and U12849 (N_12849,N_9539,N_9684);
nand U12850 (N_12850,N_9592,N_10295);
nand U12851 (N_12851,N_9613,N_9253);
or U12852 (N_12852,N_9365,N_11841);
nand U12853 (N_12853,N_11499,N_10872);
and U12854 (N_12854,N_11409,N_10555);
or U12855 (N_12855,N_11180,N_10556);
or U12856 (N_12856,N_10749,N_10005);
nor U12857 (N_12857,N_11151,N_9267);
nand U12858 (N_12858,N_11613,N_10122);
and U12859 (N_12859,N_11496,N_10851);
or U12860 (N_12860,N_11244,N_11170);
and U12861 (N_12861,N_11589,N_10890);
nand U12862 (N_12862,N_9394,N_11261);
or U12863 (N_12863,N_11939,N_11312);
nor U12864 (N_12864,N_9080,N_9962);
nor U12865 (N_12865,N_11834,N_10275);
nand U12866 (N_12866,N_10618,N_10902);
nor U12867 (N_12867,N_9104,N_10861);
or U12868 (N_12868,N_10678,N_10771);
and U12869 (N_12869,N_9627,N_11115);
nand U12870 (N_12870,N_11638,N_11986);
nor U12871 (N_12871,N_9579,N_11915);
or U12872 (N_12872,N_11925,N_9145);
nand U12873 (N_12873,N_9614,N_10583);
nand U12874 (N_12874,N_9608,N_9618);
and U12875 (N_12875,N_10636,N_11851);
and U12876 (N_12876,N_10026,N_9470);
xnor U12877 (N_12877,N_10538,N_10291);
nand U12878 (N_12878,N_10434,N_10269);
nand U12879 (N_12879,N_10537,N_10407);
nand U12880 (N_12880,N_11127,N_11435);
and U12881 (N_12881,N_11401,N_9556);
and U12882 (N_12882,N_11595,N_11030);
or U12883 (N_12883,N_10349,N_10874);
or U12884 (N_12884,N_10814,N_10135);
or U12885 (N_12885,N_11488,N_11072);
and U12886 (N_12886,N_11975,N_9494);
nand U12887 (N_12887,N_10762,N_11802);
nand U12888 (N_12888,N_10759,N_9951);
and U12889 (N_12889,N_10951,N_11321);
or U12890 (N_12890,N_11157,N_9328);
xor U12891 (N_12891,N_9459,N_11572);
nor U12892 (N_12892,N_10049,N_11288);
and U12893 (N_12893,N_11934,N_9842);
nor U12894 (N_12894,N_9024,N_9992);
xor U12895 (N_12895,N_9948,N_9803);
nor U12896 (N_12896,N_10785,N_11854);
xor U12897 (N_12897,N_10768,N_9349);
or U12898 (N_12898,N_11132,N_10389);
or U12899 (N_12899,N_10775,N_11198);
nand U12900 (N_12900,N_9999,N_10337);
nand U12901 (N_12901,N_10118,N_9637);
or U12902 (N_12902,N_11532,N_9770);
nor U12903 (N_12903,N_11672,N_10754);
or U12904 (N_12904,N_9673,N_11424);
xnor U12905 (N_12905,N_10077,N_11839);
xnor U12906 (N_12906,N_11186,N_11783);
nor U12907 (N_12907,N_11978,N_9765);
nand U12908 (N_12908,N_10298,N_10025);
nor U12909 (N_12909,N_11846,N_9538);
nor U12910 (N_12910,N_10173,N_10779);
or U12911 (N_12911,N_9667,N_9352);
or U12912 (N_12912,N_11363,N_11639);
and U12913 (N_12913,N_11771,N_9508);
and U12914 (N_12914,N_11715,N_9242);
nand U12915 (N_12915,N_10847,N_9200);
nor U12916 (N_12916,N_9440,N_11976);
or U12917 (N_12917,N_10881,N_9523);
and U12918 (N_12918,N_9901,N_10033);
nor U12919 (N_12919,N_11366,N_10842);
nor U12920 (N_12920,N_9029,N_9582);
or U12921 (N_12921,N_11586,N_10445);
and U12922 (N_12922,N_9062,N_11212);
and U12923 (N_12923,N_11293,N_10412);
or U12924 (N_12924,N_11680,N_11705);
and U12925 (N_12925,N_10109,N_9838);
nor U12926 (N_12926,N_10212,N_9291);
nor U12927 (N_12927,N_11566,N_10600);
nand U12928 (N_12928,N_11812,N_11502);
or U12929 (N_12929,N_9154,N_10258);
nor U12930 (N_12930,N_9284,N_11133);
and U12931 (N_12931,N_9346,N_10231);
and U12932 (N_12932,N_11112,N_11315);
and U12933 (N_12933,N_11842,N_11845);
nand U12934 (N_12934,N_11512,N_10962);
nand U12935 (N_12935,N_9205,N_10419);
xor U12936 (N_12936,N_11271,N_10155);
and U12937 (N_12937,N_9150,N_10760);
nor U12938 (N_12938,N_9133,N_11158);
or U12939 (N_12939,N_11808,N_11867);
nor U12940 (N_12940,N_11419,N_11899);
or U12941 (N_12941,N_11856,N_9257);
or U12942 (N_12942,N_9399,N_9392);
and U12943 (N_12943,N_10491,N_11239);
or U12944 (N_12944,N_10446,N_11436);
xor U12945 (N_12945,N_9094,N_9677);
and U12946 (N_12946,N_10397,N_9425);
nand U12947 (N_12947,N_9272,N_9598);
nand U12948 (N_12948,N_10561,N_10167);
xor U12949 (N_12949,N_11709,N_11142);
or U12950 (N_12950,N_9066,N_10343);
and U12951 (N_12951,N_11900,N_10629);
nor U12952 (N_12952,N_10989,N_11609);
nand U12953 (N_12953,N_11391,N_11848);
nand U12954 (N_12954,N_11932,N_10171);
or U12955 (N_12955,N_9997,N_10244);
or U12956 (N_12956,N_10850,N_11014);
nand U12957 (N_12957,N_11296,N_9912);
nand U12958 (N_12958,N_10745,N_10365);
nor U12959 (N_12959,N_9746,N_11568);
nand U12960 (N_12960,N_10362,N_11448);
and U12961 (N_12961,N_9843,N_10506);
and U12962 (N_12962,N_9732,N_9236);
nor U12963 (N_12963,N_11659,N_10404);
and U12964 (N_12964,N_11758,N_9035);
or U12965 (N_12965,N_9777,N_9032);
nand U12966 (N_12966,N_11527,N_9913);
and U12967 (N_12967,N_10742,N_9807);
nand U12968 (N_12968,N_9219,N_11872);
and U12969 (N_12969,N_9879,N_11330);
or U12970 (N_12970,N_10802,N_11017);
nor U12971 (N_12971,N_10984,N_9308);
or U12972 (N_12972,N_9932,N_9771);
or U12973 (N_12973,N_9812,N_10602);
nor U12974 (N_12974,N_9342,N_10973);
or U12975 (N_12975,N_11458,N_9714);
or U12976 (N_12976,N_10663,N_10248);
or U12977 (N_12977,N_9437,N_11243);
and U12978 (N_12978,N_10456,N_9648);
xor U12979 (N_12979,N_9333,N_11958);
or U12980 (N_12980,N_11692,N_9557);
and U12981 (N_12981,N_11353,N_10819);
and U12982 (N_12982,N_10512,N_10009);
and U12983 (N_12983,N_9791,N_11325);
or U12984 (N_12984,N_11283,N_10388);
and U12985 (N_12985,N_10915,N_9169);
nor U12986 (N_12986,N_9562,N_10015);
or U12987 (N_12987,N_9096,N_9679);
nor U12988 (N_12988,N_11400,N_11545);
and U12989 (N_12989,N_11980,N_10308);
nand U12990 (N_12990,N_11737,N_9910);
nor U12991 (N_12991,N_9344,N_9429);
and U12992 (N_12992,N_11619,N_11119);
nand U12993 (N_12993,N_10628,N_9740);
nor U12994 (N_12994,N_11255,N_11081);
and U12995 (N_12995,N_11711,N_9506);
and U12996 (N_12996,N_9549,N_9692);
nand U12997 (N_12997,N_10065,N_10513);
nor U12998 (N_12998,N_9330,N_10130);
and U12999 (N_12999,N_9480,N_9946);
and U13000 (N_13000,N_11473,N_10595);
nor U13001 (N_13001,N_11520,N_9351);
nor U13002 (N_13002,N_9432,N_9090);
nor U13003 (N_13003,N_10414,N_9007);
nand U13004 (N_13004,N_10625,N_10782);
xor U13005 (N_13005,N_11786,N_9478);
xnor U13006 (N_13006,N_9194,N_10268);
or U13007 (N_13007,N_9022,N_10988);
nand U13008 (N_13008,N_11762,N_9013);
xor U13009 (N_13009,N_11833,N_10299);
nor U13010 (N_13010,N_10698,N_10596);
and U13011 (N_13011,N_11724,N_9961);
nand U13012 (N_13012,N_10282,N_11477);
or U13013 (N_13013,N_11981,N_10614);
and U13014 (N_13014,N_10452,N_11840);
or U13015 (N_13015,N_10684,N_10417);
nor U13016 (N_13016,N_10741,N_10893);
and U13017 (N_13017,N_10060,N_11794);
nand U13018 (N_13018,N_9768,N_11822);
and U13019 (N_13019,N_11064,N_11879);
nor U13020 (N_13020,N_9989,N_9193);
and U13021 (N_13021,N_9103,N_11130);
nor U13022 (N_13022,N_10809,N_9170);
nor U13023 (N_13023,N_9782,N_11324);
and U13024 (N_13024,N_9441,N_10599);
nor U13025 (N_13025,N_9039,N_11074);
nand U13026 (N_13026,N_9924,N_9229);
or U13027 (N_13027,N_9282,N_9168);
or U13028 (N_13028,N_11182,N_11998);
or U13029 (N_13029,N_9975,N_10967);
nor U13030 (N_13030,N_11287,N_10639);
nor U13031 (N_13031,N_9423,N_10239);
or U13032 (N_13032,N_9385,N_9371);
and U13033 (N_13033,N_9501,N_11594);
and U13034 (N_13034,N_11318,N_10218);
and U13035 (N_13035,N_11710,N_10953);
and U13036 (N_13036,N_10665,N_11281);
nand U13037 (N_13037,N_10551,N_9271);
and U13038 (N_13038,N_10717,N_11895);
and U13039 (N_13039,N_10481,N_9383);
xnor U13040 (N_13040,N_9738,N_9449);
nand U13041 (N_13041,N_10261,N_11821);
and U13042 (N_13042,N_9124,N_9450);
or U13043 (N_13043,N_9127,N_9642);
nor U13044 (N_13044,N_9521,N_10062);
or U13045 (N_13045,N_10348,N_9087);
nor U13046 (N_13046,N_10515,N_9855);
and U13047 (N_13047,N_9457,N_10309);
or U13048 (N_13048,N_10866,N_9215);
xnor U13049 (N_13049,N_10424,N_10145);
and U13050 (N_13050,N_11858,N_11742);
or U13051 (N_13051,N_10327,N_9611);
nor U13052 (N_13052,N_11451,N_10213);
nor U13053 (N_13053,N_11016,N_11630);
and U13054 (N_13054,N_9515,N_11691);
xor U13055 (N_13055,N_11767,N_11412);
nand U13056 (N_13056,N_11446,N_10786);
xnor U13057 (N_13057,N_10767,N_10029);
nor U13058 (N_13058,N_10413,N_9641);
nor U13059 (N_13059,N_9497,N_9868);
or U13060 (N_13060,N_10449,N_9739);
nor U13061 (N_13061,N_10271,N_10611);
nor U13062 (N_13062,N_11600,N_11898);
and U13063 (N_13063,N_9000,N_10157);
xnor U13064 (N_13064,N_10451,N_10462);
nand U13065 (N_13065,N_11254,N_11062);
or U13066 (N_13066,N_11945,N_10165);
xor U13067 (N_13067,N_11857,N_9937);
xnor U13068 (N_13068,N_9416,N_10753);
nor U13069 (N_13069,N_9693,N_10470);
nand U13070 (N_13070,N_9517,N_10761);
nand U13071 (N_13071,N_10646,N_11592);
xnor U13072 (N_13072,N_10287,N_10898);
and U13073 (N_13073,N_10631,N_10965);
nand U13074 (N_13074,N_9195,N_11231);
nor U13075 (N_13075,N_9302,N_11219);
or U13076 (N_13076,N_11674,N_9357);
nor U13077 (N_13077,N_10162,N_10865);
nor U13078 (N_13078,N_11337,N_9420);
nor U13079 (N_13079,N_10623,N_9681);
and U13080 (N_13080,N_11792,N_11205);
nor U13081 (N_13081,N_10331,N_10096);
nand U13082 (N_13082,N_11013,N_11234);
nand U13083 (N_13083,N_9921,N_11156);
or U13084 (N_13084,N_10127,N_11574);
or U13085 (N_13085,N_11634,N_9362);
or U13086 (N_13086,N_11406,N_10067);
or U13087 (N_13087,N_10610,N_10177);
nand U13088 (N_13088,N_9904,N_11326);
xnor U13089 (N_13089,N_11375,N_10945);
and U13090 (N_13090,N_9226,N_9939);
or U13091 (N_13091,N_10695,N_9051);
or U13092 (N_13092,N_10532,N_11003);
nand U13093 (N_13093,N_10435,N_11612);
nor U13094 (N_13094,N_10823,N_10160);
and U13095 (N_13095,N_10566,N_11517);
nor U13096 (N_13096,N_11892,N_9317);
nor U13097 (N_13097,N_10826,N_10334);
nor U13098 (N_13098,N_10373,N_10857);
xnor U13099 (N_13099,N_10368,N_10783);
nand U13100 (N_13100,N_11591,N_9320);
xnor U13101 (N_13101,N_9654,N_9156);
nand U13102 (N_13102,N_10789,N_11275);
nor U13103 (N_13103,N_9790,N_9840);
nor U13104 (N_13104,N_11476,N_11120);
nand U13105 (N_13105,N_10175,N_11920);
nand U13106 (N_13106,N_9664,N_11819);
nor U13107 (N_13107,N_10326,N_10393);
nor U13108 (N_13108,N_9121,N_9529);
and U13109 (N_13109,N_11179,N_10323);
or U13110 (N_13110,N_10626,N_11651);
and U13111 (N_13111,N_11850,N_9587);
or U13112 (N_13112,N_11299,N_9157);
nand U13113 (N_13113,N_9495,N_11745);
nor U13114 (N_13114,N_9166,N_11949);
and U13115 (N_13115,N_11308,N_11685);
nor U13116 (N_13116,N_9091,N_9370);
and U13117 (N_13117,N_11199,N_10581);
and U13118 (N_13118,N_10010,N_9968);
nor U13119 (N_13119,N_9596,N_9696);
nand U13120 (N_13120,N_9984,N_11025);
and U13121 (N_13121,N_9413,N_10549);
nand U13122 (N_13122,N_10991,N_9675);
and U13123 (N_13123,N_10570,N_11929);
nand U13124 (N_13124,N_10075,N_10285);
xnor U13125 (N_13125,N_9970,N_11046);
nor U13126 (N_13126,N_11816,N_9375);
nor U13127 (N_13127,N_11093,N_11402);
or U13128 (N_13128,N_10878,N_9277);
or U13129 (N_13129,N_9276,N_9686);
or U13130 (N_13130,N_9438,N_11018);
xnor U13131 (N_13131,N_9191,N_11778);
nand U13132 (N_13132,N_11621,N_11253);
or U13133 (N_13133,N_11687,N_11109);
xor U13134 (N_13134,N_11614,N_11627);
nor U13135 (N_13135,N_11304,N_10976);
and U13136 (N_13136,N_10505,N_11942);
nor U13137 (N_13137,N_10128,N_11779);
nor U13138 (N_13138,N_10041,N_10214);
nand U13139 (N_13139,N_11585,N_10257);
or U13140 (N_13140,N_10605,N_9918);
xnor U13141 (N_13141,N_11541,N_11781);
nand U13142 (N_13142,N_10103,N_9288);
or U13143 (N_13143,N_9281,N_10938);
or U13144 (N_13144,N_11536,N_9757);
and U13145 (N_13145,N_9632,N_10859);
or U13146 (N_13146,N_10453,N_10748);
xnor U13147 (N_13147,N_11829,N_10907);
or U13148 (N_13148,N_11966,N_11657);
nand U13149 (N_13149,N_10203,N_9846);
or U13150 (N_13150,N_11084,N_9431);
nor U13151 (N_13151,N_10490,N_10409);
or U13152 (N_13152,N_11146,N_11602);
nand U13153 (N_13153,N_9741,N_9774);
and U13154 (N_13154,N_10964,N_11434);
nand U13155 (N_13155,N_10685,N_9787);
xnor U13156 (N_13156,N_11757,N_10744);
nand U13157 (N_13157,N_11714,N_11309);
nor U13158 (N_13158,N_9115,N_11649);
or U13159 (N_13159,N_9862,N_9841);
or U13160 (N_13160,N_10019,N_9110);
and U13161 (N_13161,N_11650,N_11202);
or U13162 (N_13162,N_10303,N_10454);
nor U13163 (N_13163,N_11501,N_10763);
and U13164 (N_13164,N_9624,N_10756);
xnor U13165 (N_13165,N_10030,N_10219);
xnor U13166 (N_13166,N_11852,N_11665);
and U13167 (N_13167,N_11300,N_11996);
nor U13168 (N_13168,N_9335,N_10350);
nand U13169 (N_13169,N_10728,N_11655);
nand U13170 (N_13170,N_9589,N_9421);
and U13171 (N_13171,N_11316,N_11964);
nand U13172 (N_13172,N_11066,N_10080);
xor U13173 (N_13173,N_11921,N_9128);
xor U13174 (N_13174,N_11295,N_10100);
xor U13175 (N_13175,N_11396,N_10315);
nand U13176 (N_13176,N_11701,N_10047);
or U13177 (N_13177,N_9381,N_11537);
nand U13178 (N_13178,N_11523,N_11086);
xnor U13179 (N_13179,N_11569,N_10920);
and U13180 (N_13180,N_11623,N_10296);
nor U13181 (N_13181,N_11089,N_10381);
and U13182 (N_13182,N_10875,N_11148);
or U13183 (N_13183,N_10994,N_9600);
or U13184 (N_13184,N_9577,N_9188);
nand U13185 (N_13185,N_9132,N_9510);
xnor U13186 (N_13186,N_10941,N_11818);
and U13187 (N_13187,N_11551,N_9484);
and U13188 (N_13188,N_9496,N_11290);
nor U13189 (N_13189,N_9260,N_10577);
nor U13190 (N_13190,N_10444,N_9318);
nor U13191 (N_13191,N_10134,N_10730);
xor U13192 (N_13192,N_10769,N_10939);
nand U13193 (N_13193,N_11992,N_9870);
and U13194 (N_13194,N_9898,N_10235);
nand U13195 (N_13195,N_10206,N_11991);
and U13196 (N_13196,N_10660,N_9027);
or U13197 (N_13197,N_11675,N_10682);
nor U13198 (N_13198,N_9559,N_11162);
and U13199 (N_13199,N_9530,N_11333);
or U13200 (N_13200,N_9424,N_9695);
nand U13201 (N_13201,N_11150,N_9004);
and U13202 (N_13202,N_10237,N_11140);
or U13203 (N_13203,N_10321,N_9674);
nor U13204 (N_13204,N_10114,N_11328);
nor U13205 (N_13205,N_11061,N_9266);
nand U13206 (N_13206,N_11426,N_9651);
nor U13207 (N_13207,N_10734,N_9373);
nor U13208 (N_13208,N_9112,N_11919);
and U13209 (N_13209,N_9158,N_10811);
nor U13210 (N_13210,N_10680,N_11766);
nor U13211 (N_13211,N_10181,N_11636);
nand U13212 (N_13212,N_10043,N_10963);
or U13213 (N_13213,N_10909,N_11004);
nor U13214 (N_13214,N_10726,N_10638);
nor U13215 (N_13215,N_9957,N_9733);
and U13216 (N_13216,N_9906,N_11927);
nand U13217 (N_13217,N_9827,N_10238);
nand U13218 (N_13218,N_9426,N_10511);
xor U13219 (N_13219,N_9863,N_9428);
nand U13220 (N_13220,N_10535,N_11492);
or U13221 (N_13221,N_9489,N_11416);
xor U13222 (N_13222,N_11880,N_9938);
nor U13223 (N_13223,N_10052,N_11635);
xnor U13224 (N_13224,N_9048,N_11126);
xor U13225 (N_13225,N_10290,N_11957);
xnor U13226 (N_13226,N_11101,N_11640);
nor U13227 (N_13227,N_11901,N_9481);
and U13228 (N_13228,N_11350,N_9982);
and U13229 (N_13229,N_11188,N_10408);
nor U13230 (N_13230,N_9010,N_11339);
nand U13231 (N_13231,N_9334,N_10668);
or U13232 (N_13232,N_9341,N_11928);
and U13233 (N_13233,N_9222,N_10542);
nor U13234 (N_13234,N_11039,N_9666);
and U13235 (N_13235,N_9433,N_11415);
nand U13236 (N_13236,N_9210,N_10284);
nand U13237 (N_13237,N_11855,N_10028);
nor U13238 (N_13238,N_10968,N_9623);
or U13239 (N_13239,N_11985,N_10223);
nor U13240 (N_13240,N_10925,N_11117);
and U13241 (N_13241,N_10059,N_10926);
nor U13242 (N_13242,N_10457,N_10622);
or U13243 (N_13243,N_11736,N_9857);
or U13244 (N_13244,N_9213,N_11972);
and U13245 (N_13245,N_10868,N_10146);
nor U13246 (N_13246,N_9941,N_10718);
or U13247 (N_13247,N_9711,N_10681);
nor U13248 (N_13248,N_10188,N_11534);
nor U13249 (N_13249,N_10545,N_11667);
and U13250 (N_13250,N_11575,N_11886);
nor U13251 (N_13251,N_9516,N_10215);
nor U13252 (N_13252,N_11069,N_9378);
or U13253 (N_13253,N_10153,N_9001);
and U13254 (N_13254,N_11656,N_11439);
nand U13255 (N_13255,N_9694,N_10746);
nand U13256 (N_13256,N_10084,N_10374);
or U13257 (N_13257,N_11631,N_10927);
and U13258 (N_13258,N_11729,N_10124);
and U13259 (N_13259,N_9811,N_11804);
nand U13260 (N_13260,N_10957,N_10091);
xor U13261 (N_13261,N_11358,N_9233);
and U13262 (N_13262,N_9479,N_9043);
or U13263 (N_13263,N_9221,N_9120);
nor U13264 (N_13264,N_9028,N_9853);
or U13265 (N_13265,N_9086,N_10488);
or U13266 (N_13266,N_10256,N_9218);
nor U13267 (N_13267,N_10314,N_9712);
nor U13268 (N_13268,N_11570,N_10541);
nand U13269 (N_13269,N_11678,N_11164);
nor U13270 (N_13270,N_9348,N_10956);
xor U13271 (N_13271,N_9136,N_9751);
and U13272 (N_13272,N_10144,N_9100);
and U13273 (N_13273,N_9314,N_9458);
nor U13274 (N_13274,N_10539,N_9823);
or U13275 (N_13275,N_9363,N_10831);
or U13276 (N_13276,N_9639,N_11035);
and U13277 (N_13277,N_9243,N_10432);
xor U13278 (N_13278,N_10924,N_10870);
nand U13279 (N_13279,N_9594,N_9264);
nand U13280 (N_13280,N_9798,N_9796);
nor U13281 (N_13281,N_9165,N_9890);
and U13282 (N_13282,N_11041,N_11515);
nor U13283 (N_13283,N_9175,N_10137);
nand U13284 (N_13284,N_11122,N_9856);
or U13285 (N_13285,N_9395,N_10274);
nor U13286 (N_13286,N_9908,N_11510);
xor U13287 (N_13287,N_10777,N_10833);
nand U13288 (N_13288,N_11250,N_10670);
and U13289 (N_13289,N_11693,N_11197);
nor U13290 (N_13290,N_11629,N_10526);
or U13291 (N_13291,N_11103,N_9172);
nand U13292 (N_13292,N_11457,N_9764);
and U13293 (N_13293,N_9612,N_10489);
nand U13294 (N_13294,N_11873,N_9114);
nand U13295 (N_13295,N_11628,N_11341);
and U13296 (N_13296,N_9818,N_10352);
nor U13297 (N_13297,N_9285,N_10042);
or U13298 (N_13298,N_9545,N_11479);
nor U13299 (N_13299,N_11144,N_10986);
and U13300 (N_13300,N_10912,N_9894);
nor U13301 (N_13301,N_11008,N_9719);
or U13302 (N_13302,N_10272,N_10574);
xnor U13303 (N_13303,N_9098,N_9505);
or U13304 (N_13304,N_9491,N_10180);
nor U13305 (N_13305,N_11238,N_11751);
or U13306 (N_13306,N_10706,N_11498);
xnor U13307 (N_13307,N_9180,N_10302);
nand U13308 (N_13308,N_11844,N_9407);
nand U13309 (N_13309,N_9899,N_11042);
and U13310 (N_13310,N_10364,N_9289);
and U13311 (N_13311,N_10338,N_9377);
xnor U13312 (N_13312,N_9337,N_11351);
nor U13313 (N_13313,N_10119,N_11099);
nand U13314 (N_13314,N_9287,N_11673);
or U13315 (N_13315,N_9944,N_10954);
nand U13316 (N_13316,N_11106,N_9810);
nand U13317 (N_13317,N_11894,N_10979);
nor U13318 (N_13318,N_11267,N_9513);
nor U13319 (N_13319,N_11430,N_10727);
or U13320 (N_13320,N_9319,N_10089);
or U13321 (N_13321,N_9089,N_11977);
or U13322 (N_13322,N_9806,N_9959);
xnor U13323 (N_13323,N_10560,N_11208);
nor U13324 (N_13324,N_10416,N_11826);
nand U13325 (N_13325,N_9934,N_10070);
nor U13326 (N_13326,N_11334,N_11787);
or U13327 (N_13327,N_9498,N_10942);
and U13328 (N_13328,N_9852,N_9543);
and U13329 (N_13329,N_11676,N_10720);
nor U13330 (N_13330,N_11489,N_11604);
nor U13331 (N_13331,N_11083,N_9430);
or U13332 (N_13332,N_9278,N_10224);
nor U13333 (N_13333,N_9081,N_11361);
nand U13334 (N_13334,N_9034,N_11467);
xnor U13335 (N_13335,N_11703,N_11943);
nor U13336 (N_13336,N_9881,N_9636);
or U13337 (N_13337,N_11307,N_10612);
and U13338 (N_13338,N_10463,N_10024);
nand U13339 (N_13339,N_9072,N_9473);
xnor U13340 (N_13340,N_11531,N_9550);
nor U13341 (N_13341,N_11982,N_10580);
and U13342 (N_13342,N_9874,N_11116);
and U13343 (N_13343,N_11557,N_9555);
and U13344 (N_13344,N_9361,N_11470);
or U13345 (N_13345,N_9885,N_11564);
and U13346 (N_13346,N_11166,N_9647);
xor U13347 (N_13347,N_11027,N_10395);
xnor U13348 (N_13348,N_9653,N_10836);
nor U13349 (N_13349,N_11838,N_11805);
or U13350 (N_13350,N_9554,N_9088);
nor U13351 (N_13351,N_9819,N_10508);
or U13352 (N_13352,N_10892,N_9398);
nor U13353 (N_13353,N_11377,N_9082);
nor U13354 (N_13354,N_11747,N_9546);
or U13355 (N_13355,N_10619,N_10469);
nor U13356 (N_13356,N_11444,N_10601);
xor U13357 (N_13357,N_11217,N_11593);
nand U13358 (N_13358,N_9527,N_9644);
and U13359 (N_13359,N_10149,N_11440);
or U13360 (N_13360,N_11336,N_11963);
or U13361 (N_13361,N_10277,N_9463);
and U13362 (N_13362,N_9988,N_11653);
nor U13363 (N_13363,N_10151,N_11045);
nor U13364 (N_13364,N_10736,N_9101);
and U13365 (N_13365,N_9409,N_11940);
or U13366 (N_13366,N_11189,N_10333);
nand U13367 (N_13367,N_9353,N_10192);
nor U13368 (N_13368,N_11007,N_10830);
or U13369 (N_13369,N_9389,N_11237);
nand U13370 (N_13370,N_10143,N_9054);
xnor U13371 (N_13371,N_10658,N_9558);
nor U13372 (N_13372,N_11349,N_11068);
nand U13373 (N_13373,N_11529,N_9744);
or U13374 (N_13374,N_11951,N_10141);
nand U13375 (N_13375,N_11169,N_9401);
nand U13376 (N_13376,N_10800,N_11063);
and U13377 (N_13377,N_10106,N_11323);
or U13378 (N_13378,N_9265,N_10262);
nand U13379 (N_13379,N_9414,N_11052);
and U13380 (N_13380,N_10204,N_11935);
or U13381 (N_13381,N_9769,N_10022);
nand U13382 (N_13382,N_11918,N_9907);
nand U13383 (N_13383,N_9187,N_11696);
or U13384 (N_13384,N_9294,N_11956);
nand U13385 (N_13385,N_9680,N_10170);
or U13386 (N_13386,N_10750,N_9073);
nand U13387 (N_13387,N_10102,N_9003);
nand U13388 (N_13388,N_10289,N_10037);
nand U13389 (N_13389,N_10086,N_10038);
or U13390 (N_13390,N_9839,N_11381);
nor U13391 (N_13391,N_10543,N_10464);
or U13392 (N_13392,N_11427,N_11831);
nand U13393 (N_13393,N_10675,N_9595);
and U13394 (N_13394,N_11491,N_10074);
or U13395 (N_13395,N_11225,N_10467);
nand U13396 (N_13396,N_9566,N_10937);
xor U13397 (N_13397,N_11114,N_11228);
nand U13398 (N_13398,N_10240,N_11305);
xor U13399 (N_13399,N_9359,N_9987);
and U13400 (N_13400,N_9125,N_10465);
and U13401 (N_13401,N_10207,N_10310);
nand U13402 (N_13402,N_9374,N_10630);
nand U13403 (N_13403,N_9367,N_10676);
nor U13404 (N_13404,N_9616,N_9661);
nor U13405 (N_13405,N_11668,N_10174);
or U13406 (N_13406,N_11888,N_11909);
or U13407 (N_13407,N_11853,N_9047);
and U13408 (N_13408,N_11317,N_10066);
nor U13409 (N_13409,N_9148,N_11922);
nand U13410 (N_13410,N_10958,N_9042);
and U13411 (N_13411,N_11141,N_9189);
xor U13412 (N_13412,N_10247,N_10952);
nor U13413 (N_13413,N_9979,N_9461);
nand U13414 (N_13414,N_11051,N_11475);
nor U13415 (N_13415,N_10770,N_10587);
or U13416 (N_13416,N_9405,N_10484);
and U13417 (N_13417,N_11791,N_10372);
and U13418 (N_13418,N_9386,N_11514);
or U13419 (N_13419,N_11469,N_9965);
and U13420 (N_13420,N_9699,N_9391);
nand U13421 (N_13421,N_11740,N_9234);
or U13422 (N_13422,N_11044,N_10200);
nor U13423 (N_13423,N_10288,N_9726);
and U13424 (N_13424,N_9575,N_10843);
and U13425 (N_13425,N_10657,N_9936);
nand U13426 (N_13426,N_11993,N_10530);
nand U13427 (N_13427,N_10400,N_9930);
nor U13428 (N_13428,N_10379,N_9650);
nand U13429 (N_13429,N_9969,N_10292);
and U13430 (N_13430,N_9055,N_9781);
nand U13431 (N_13431,N_9903,N_9471);
nor U13432 (N_13432,N_11984,N_9920);
or U13433 (N_13433,N_9382,N_11866);
nand U13434 (N_13434,N_11882,N_10139);
and U13435 (N_13435,N_9018,N_11462);
and U13436 (N_13436,N_9886,N_9585);
nor U13437 (N_13437,N_10849,N_11750);
or U13438 (N_13438,N_10339,N_11005);
nand U13439 (N_13439,N_9364,N_11263);
nor U13440 (N_13440,N_11849,N_11053);
nor U13441 (N_13441,N_9161,N_11582);
nor U13442 (N_13442,N_9454,N_10546);
or U13443 (N_13443,N_9858,N_11790);
nor U13444 (N_13444,N_9833,N_10643);
nand U13445 (N_13445,N_10471,N_11795);
nand U13446 (N_13446,N_10940,N_9307);
nor U13447 (N_13447,N_9742,N_9783);
nand U13448 (N_13448,N_9209,N_10617);
nor U13449 (N_13449,N_9588,N_9117);
nor U13450 (N_13450,N_9023,N_9056);
nor U13451 (N_13451,N_10780,N_11506);
nand U13452 (N_13452,N_10163,N_11414);
and U13453 (N_13453,N_11429,N_9814);
nor U13454 (N_13454,N_9123,N_11165);
or U13455 (N_13455,N_10627,N_10805);
nor U13456 (N_13456,N_9954,N_10328);
or U13457 (N_13457,N_11280,N_10385);
and U13458 (N_13458,N_11620,N_10242);
or U13459 (N_13459,N_11428,N_10674);
nor U13460 (N_13460,N_10827,N_11001);
or U13461 (N_13461,N_10324,N_11291);
and U13462 (N_13462,N_9512,N_10190);
or U13463 (N_13463,N_9601,N_10426);
nor U13464 (N_13464,N_9955,N_10136);
and U13465 (N_13465,N_9687,N_10671);
nand U13466 (N_13466,N_10594,N_11799);
nand U13467 (N_13467,N_11466,N_10054);
nor U13468 (N_13468,N_9893,N_11608);
nand U13469 (N_13469,N_10064,N_9300);
and U13470 (N_13470,N_9152,N_11800);
nand U13471 (N_13471,N_10563,N_9872);
or U13472 (N_13472,N_10342,N_10961);
or U13473 (N_13473,N_10384,N_10603);
nor U13474 (N_13474,N_10110,N_9331);
xnor U13475 (N_13475,N_11082,N_10873);
nor U13476 (N_13476,N_9590,N_11911);
nand U13477 (N_13477,N_11837,N_11137);
xnor U13478 (N_13478,N_11380,N_11598);
xor U13479 (N_13479,N_11327,N_11224);
nand U13480 (N_13480,N_9990,N_11518);
and U13481 (N_13481,N_9748,N_10791);
or U13482 (N_13482,N_10582,N_9469);
nor U13483 (N_13483,N_9993,N_11903);
and U13484 (N_13484,N_11553,N_11096);
nand U13485 (N_13485,N_9646,N_9705);
and U13486 (N_13486,N_11983,N_10841);
or U13487 (N_13487,N_11577,N_9465);
nor U13488 (N_13488,N_9795,N_11788);
xor U13489 (N_13489,N_10987,N_9672);
and U13490 (N_13490,N_10081,N_11393);
and U13491 (N_13491,N_9049,N_11931);
nand U13492 (N_13492,N_11193,N_9083);
nand U13493 (N_13493,N_10386,N_10347);
and U13494 (N_13494,N_11232,N_11367);
and U13495 (N_13495,N_11753,N_9869);
and U13496 (N_13496,N_11111,N_9061);
or U13497 (N_13497,N_11755,N_9720);
xor U13498 (N_13498,N_10073,N_11548);
and U13499 (N_13499,N_11887,N_11717);
xor U13500 (N_13500,N_11344,N_11925);
or U13501 (N_13501,N_10858,N_9588);
nor U13502 (N_13502,N_10282,N_11154);
nor U13503 (N_13503,N_11669,N_9423);
and U13504 (N_13504,N_9781,N_11017);
nand U13505 (N_13505,N_11926,N_9505);
nand U13506 (N_13506,N_11681,N_10850);
or U13507 (N_13507,N_9823,N_11487);
nor U13508 (N_13508,N_11402,N_11340);
nand U13509 (N_13509,N_11588,N_9915);
nand U13510 (N_13510,N_10390,N_11775);
and U13511 (N_13511,N_9010,N_9245);
nor U13512 (N_13512,N_11750,N_11403);
and U13513 (N_13513,N_10669,N_10706);
or U13514 (N_13514,N_10505,N_11073);
nor U13515 (N_13515,N_9828,N_9472);
nand U13516 (N_13516,N_9269,N_10818);
xor U13517 (N_13517,N_9550,N_11847);
and U13518 (N_13518,N_11305,N_9451);
or U13519 (N_13519,N_11870,N_9586);
nor U13520 (N_13520,N_9266,N_10783);
or U13521 (N_13521,N_10007,N_11305);
or U13522 (N_13522,N_10978,N_11519);
nor U13523 (N_13523,N_11612,N_10228);
or U13524 (N_13524,N_9581,N_10430);
xor U13525 (N_13525,N_11006,N_9609);
nor U13526 (N_13526,N_10519,N_9437);
and U13527 (N_13527,N_9986,N_10289);
nand U13528 (N_13528,N_11238,N_9260);
xor U13529 (N_13529,N_10496,N_9738);
or U13530 (N_13530,N_9724,N_11407);
nand U13531 (N_13531,N_9094,N_9553);
nand U13532 (N_13532,N_11630,N_11055);
xor U13533 (N_13533,N_11074,N_11931);
and U13534 (N_13534,N_10387,N_11510);
nand U13535 (N_13535,N_9919,N_9308);
nand U13536 (N_13536,N_9044,N_11308);
and U13537 (N_13537,N_9823,N_11469);
nand U13538 (N_13538,N_9763,N_9163);
nor U13539 (N_13539,N_10320,N_10084);
and U13540 (N_13540,N_11755,N_9318);
nor U13541 (N_13541,N_11531,N_9623);
nor U13542 (N_13542,N_10265,N_9406);
or U13543 (N_13543,N_10441,N_10738);
nor U13544 (N_13544,N_10804,N_9016);
nor U13545 (N_13545,N_10174,N_10678);
nor U13546 (N_13546,N_10640,N_9679);
xnor U13547 (N_13547,N_11639,N_10805);
or U13548 (N_13548,N_11382,N_10973);
nor U13549 (N_13549,N_10116,N_9154);
xnor U13550 (N_13550,N_9160,N_9752);
nor U13551 (N_13551,N_10339,N_10444);
nor U13552 (N_13552,N_11583,N_11396);
nor U13553 (N_13553,N_10171,N_10649);
nand U13554 (N_13554,N_10070,N_10467);
and U13555 (N_13555,N_10418,N_9765);
and U13556 (N_13556,N_10743,N_10197);
xor U13557 (N_13557,N_10874,N_11758);
nand U13558 (N_13558,N_10857,N_10957);
xor U13559 (N_13559,N_11003,N_10456);
xnor U13560 (N_13560,N_10572,N_9877);
nand U13561 (N_13561,N_11608,N_11896);
nor U13562 (N_13562,N_10019,N_11189);
xor U13563 (N_13563,N_11123,N_10857);
and U13564 (N_13564,N_9244,N_10495);
and U13565 (N_13565,N_10623,N_9545);
or U13566 (N_13566,N_9859,N_11796);
and U13567 (N_13567,N_9821,N_9187);
and U13568 (N_13568,N_9877,N_10422);
and U13569 (N_13569,N_10883,N_9465);
nor U13570 (N_13570,N_11508,N_11771);
and U13571 (N_13571,N_10290,N_11926);
nor U13572 (N_13572,N_11891,N_10737);
xor U13573 (N_13573,N_9372,N_11617);
or U13574 (N_13574,N_10037,N_11989);
xnor U13575 (N_13575,N_10768,N_10464);
and U13576 (N_13576,N_10902,N_10137);
and U13577 (N_13577,N_10437,N_9047);
or U13578 (N_13578,N_10420,N_10776);
nand U13579 (N_13579,N_9280,N_10450);
nand U13580 (N_13580,N_9392,N_10675);
nor U13581 (N_13581,N_9718,N_9540);
nand U13582 (N_13582,N_9050,N_11670);
or U13583 (N_13583,N_9960,N_10467);
and U13584 (N_13584,N_9652,N_11780);
xor U13585 (N_13585,N_11848,N_10946);
nand U13586 (N_13586,N_11644,N_11664);
nand U13587 (N_13587,N_10570,N_11182);
xor U13588 (N_13588,N_10029,N_9391);
or U13589 (N_13589,N_11314,N_9278);
nand U13590 (N_13590,N_11659,N_10920);
or U13591 (N_13591,N_11114,N_10426);
nand U13592 (N_13592,N_11178,N_9232);
or U13593 (N_13593,N_11327,N_11471);
nand U13594 (N_13594,N_11304,N_11420);
xor U13595 (N_13595,N_11730,N_9359);
nand U13596 (N_13596,N_11186,N_11353);
xor U13597 (N_13597,N_9441,N_9452);
nand U13598 (N_13598,N_10834,N_10308);
nand U13599 (N_13599,N_10790,N_9643);
nor U13600 (N_13600,N_11043,N_11004);
nor U13601 (N_13601,N_10955,N_11119);
and U13602 (N_13602,N_11524,N_11134);
or U13603 (N_13603,N_9710,N_10836);
nor U13604 (N_13604,N_11940,N_9381);
or U13605 (N_13605,N_10936,N_9628);
nor U13606 (N_13606,N_10414,N_11081);
nor U13607 (N_13607,N_9855,N_10444);
nor U13608 (N_13608,N_11028,N_11306);
or U13609 (N_13609,N_9095,N_9249);
xor U13610 (N_13610,N_10954,N_11028);
nor U13611 (N_13611,N_11820,N_10814);
or U13612 (N_13612,N_9049,N_10283);
nor U13613 (N_13613,N_11922,N_11567);
or U13614 (N_13614,N_11316,N_10378);
or U13615 (N_13615,N_10096,N_11254);
and U13616 (N_13616,N_10058,N_9832);
or U13617 (N_13617,N_11819,N_9669);
nor U13618 (N_13618,N_10791,N_10656);
or U13619 (N_13619,N_9295,N_9485);
and U13620 (N_13620,N_11724,N_11082);
and U13621 (N_13621,N_10319,N_9516);
nand U13622 (N_13622,N_11985,N_10653);
and U13623 (N_13623,N_11266,N_10805);
nand U13624 (N_13624,N_10138,N_10824);
nor U13625 (N_13625,N_10268,N_10812);
nor U13626 (N_13626,N_11554,N_11256);
and U13627 (N_13627,N_10418,N_9986);
xor U13628 (N_13628,N_10997,N_9005);
nor U13629 (N_13629,N_10301,N_10266);
or U13630 (N_13630,N_9915,N_10257);
and U13631 (N_13631,N_11655,N_10216);
nand U13632 (N_13632,N_9382,N_10363);
nand U13633 (N_13633,N_9031,N_9748);
and U13634 (N_13634,N_11617,N_9926);
and U13635 (N_13635,N_9137,N_10819);
and U13636 (N_13636,N_11610,N_10613);
nor U13637 (N_13637,N_10791,N_11786);
and U13638 (N_13638,N_10617,N_11414);
or U13639 (N_13639,N_10923,N_11403);
and U13640 (N_13640,N_11202,N_9134);
nand U13641 (N_13641,N_9915,N_10659);
and U13642 (N_13642,N_9281,N_10430);
nand U13643 (N_13643,N_10445,N_9726);
nor U13644 (N_13644,N_9201,N_11465);
xor U13645 (N_13645,N_10512,N_10213);
xnor U13646 (N_13646,N_10511,N_10944);
or U13647 (N_13647,N_9566,N_11792);
nand U13648 (N_13648,N_9975,N_9493);
xnor U13649 (N_13649,N_10576,N_11584);
and U13650 (N_13650,N_10556,N_10413);
and U13651 (N_13651,N_9761,N_10275);
nand U13652 (N_13652,N_10945,N_9756);
nor U13653 (N_13653,N_9038,N_9353);
nand U13654 (N_13654,N_9643,N_10274);
nor U13655 (N_13655,N_10334,N_11421);
or U13656 (N_13656,N_11267,N_11437);
nand U13657 (N_13657,N_11751,N_11174);
nor U13658 (N_13658,N_9308,N_11717);
or U13659 (N_13659,N_10513,N_11366);
nor U13660 (N_13660,N_11671,N_11140);
and U13661 (N_13661,N_9677,N_11789);
xor U13662 (N_13662,N_10397,N_10124);
and U13663 (N_13663,N_9362,N_10956);
nand U13664 (N_13664,N_11122,N_9877);
and U13665 (N_13665,N_10460,N_10798);
and U13666 (N_13666,N_9245,N_11128);
or U13667 (N_13667,N_10911,N_11213);
or U13668 (N_13668,N_9537,N_9291);
nand U13669 (N_13669,N_11386,N_9437);
xnor U13670 (N_13670,N_10559,N_9172);
and U13671 (N_13671,N_10395,N_11447);
nor U13672 (N_13672,N_9044,N_9635);
nand U13673 (N_13673,N_9088,N_11355);
and U13674 (N_13674,N_11847,N_9612);
nor U13675 (N_13675,N_9083,N_10997);
and U13676 (N_13676,N_9710,N_9857);
nor U13677 (N_13677,N_10966,N_10139);
nand U13678 (N_13678,N_10514,N_11746);
and U13679 (N_13679,N_10244,N_9991);
nor U13680 (N_13680,N_11916,N_10414);
nor U13681 (N_13681,N_11646,N_9722);
nor U13682 (N_13682,N_10835,N_10906);
xnor U13683 (N_13683,N_11925,N_10295);
and U13684 (N_13684,N_11473,N_11161);
nor U13685 (N_13685,N_11588,N_9951);
and U13686 (N_13686,N_10233,N_10109);
nor U13687 (N_13687,N_11295,N_10745);
nor U13688 (N_13688,N_11679,N_11115);
nor U13689 (N_13689,N_10851,N_11679);
and U13690 (N_13690,N_10759,N_9112);
and U13691 (N_13691,N_9908,N_10018);
or U13692 (N_13692,N_11435,N_10865);
and U13693 (N_13693,N_11175,N_11980);
nor U13694 (N_13694,N_11953,N_10689);
or U13695 (N_13695,N_10154,N_10272);
nand U13696 (N_13696,N_11660,N_11873);
or U13697 (N_13697,N_11165,N_10062);
and U13698 (N_13698,N_10575,N_10394);
nand U13699 (N_13699,N_11330,N_10767);
xor U13700 (N_13700,N_10949,N_9988);
nand U13701 (N_13701,N_9902,N_11371);
nand U13702 (N_13702,N_10895,N_11107);
and U13703 (N_13703,N_10620,N_10700);
and U13704 (N_13704,N_11626,N_9249);
and U13705 (N_13705,N_9756,N_9469);
nand U13706 (N_13706,N_10203,N_10904);
and U13707 (N_13707,N_10638,N_10308);
nand U13708 (N_13708,N_11564,N_9720);
xor U13709 (N_13709,N_11404,N_9592);
or U13710 (N_13710,N_9982,N_9641);
and U13711 (N_13711,N_10153,N_10103);
nor U13712 (N_13712,N_11320,N_10944);
or U13713 (N_13713,N_11732,N_11254);
nand U13714 (N_13714,N_9554,N_9139);
nand U13715 (N_13715,N_10751,N_11622);
xnor U13716 (N_13716,N_9919,N_9277);
and U13717 (N_13717,N_11202,N_9015);
nor U13718 (N_13718,N_10798,N_11622);
or U13719 (N_13719,N_9533,N_10097);
and U13720 (N_13720,N_9340,N_9677);
nand U13721 (N_13721,N_9061,N_10277);
xor U13722 (N_13722,N_10088,N_9828);
and U13723 (N_13723,N_10759,N_10054);
nor U13724 (N_13724,N_11980,N_10825);
nand U13725 (N_13725,N_10062,N_10521);
nor U13726 (N_13726,N_11848,N_10106);
and U13727 (N_13727,N_10115,N_11130);
and U13728 (N_13728,N_11780,N_10514);
and U13729 (N_13729,N_9375,N_9184);
and U13730 (N_13730,N_10360,N_10835);
nand U13731 (N_13731,N_10364,N_9872);
xor U13732 (N_13732,N_11421,N_9233);
nand U13733 (N_13733,N_10605,N_11843);
and U13734 (N_13734,N_10369,N_9858);
and U13735 (N_13735,N_9269,N_9492);
or U13736 (N_13736,N_10240,N_9944);
nor U13737 (N_13737,N_10630,N_11140);
or U13738 (N_13738,N_11360,N_9344);
nand U13739 (N_13739,N_9275,N_10125);
and U13740 (N_13740,N_9705,N_11992);
nand U13741 (N_13741,N_10906,N_11264);
nor U13742 (N_13742,N_10129,N_9222);
and U13743 (N_13743,N_10900,N_9229);
or U13744 (N_13744,N_10429,N_9278);
xor U13745 (N_13745,N_11772,N_10512);
nor U13746 (N_13746,N_11884,N_11619);
or U13747 (N_13747,N_9743,N_10014);
nand U13748 (N_13748,N_9677,N_11012);
nand U13749 (N_13749,N_10544,N_10523);
nor U13750 (N_13750,N_9212,N_10133);
nand U13751 (N_13751,N_9940,N_10160);
and U13752 (N_13752,N_9326,N_11047);
or U13753 (N_13753,N_9528,N_9769);
nor U13754 (N_13754,N_11811,N_11749);
or U13755 (N_13755,N_9922,N_9339);
nor U13756 (N_13756,N_10837,N_9001);
and U13757 (N_13757,N_11298,N_11155);
nand U13758 (N_13758,N_11683,N_11681);
and U13759 (N_13759,N_9020,N_10040);
nor U13760 (N_13760,N_11603,N_9647);
or U13761 (N_13761,N_10017,N_9594);
and U13762 (N_13762,N_11190,N_9991);
and U13763 (N_13763,N_11295,N_11428);
nor U13764 (N_13764,N_10334,N_11209);
xor U13765 (N_13765,N_11962,N_11585);
xnor U13766 (N_13766,N_10577,N_9367);
and U13767 (N_13767,N_11383,N_10169);
nor U13768 (N_13768,N_9824,N_10386);
nor U13769 (N_13769,N_11364,N_11947);
nor U13770 (N_13770,N_9198,N_10652);
and U13771 (N_13771,N_11234,N_10352);
nand U13772 (N_13772,N_10561,N_10172);
nor U13773 (N_13773,N_9560,N_9104);
nor U13774 (N_13774,N_11281,N_11995);
and U13775 (N_13775,N_9997,N_11078);
nand U13776 (N_13776,N_11465,N_9355);
or U13777 (N_13777,N_10322,N_10098);
xnor U13778 (N_13778,N_10268,N_10630);
and U13779 (N_13779,N_10696,N_10621);
nand U13780 (N_13780,N_9361,N_10129);
nand U13781 (N_13781,N_10399,N_10426);
nand U13782 (N_13782,N_9237,N_11750);
and U13783 (N_13783,N_10837,N_9844);
nor U13784 (N_13784,N_10449,N_10757);
nor U13785 (N_13785,N_10883,N_10366);
xor U13786 (N_13786,N_11709,N_9526);
nand U13787 (N_13787,N_11851,N_10419);
xor U13788 (N_13788,N_9356,N_9746);
nor U13789 (N_13789,N_9743,N_11903);
nor U13790 (N_13790,N_10821,N_9141);
and U13791 (N_13791,N_11418,N_11479);
or U13792 (N_13792,N_11894,N_11242);
or U13793 (N_13793,N_9870,N_10908);
nand U13794 (N_13794,N_9247,N_11145);
nand U13795 (N_13795,N_11225,N_11815);
nor U13796 (N_13796,N_11616,N_11277);
xnor U13797 (N_13797,N_11549,N_9187);
xor U13798 (N_13798,N_10447,N_11837);
or U13799 (N_13799,N_11926,N_11985);
nor U13800 (N_13800,N_9595,N_11654);
or U13801 (N_13801,N_11164,N_9815);
nand U13802 (N_13802,N_10104,N_10809);
nand U13803 (N_13803,N_11777,N_10134);
nor U13804 (N_13804,N_11488,N_9413);
nor U13805 (N_13805,N_10404,N_10954);
nand U13806 (N_13806,N_11910,N_9270);
nor U13807 (N_13807,N_9199,N_10634);
or U13808 (N_13808,N_10525,N_11467);
and U13809 (N_13809,N_11338,N_10471);
nor U13810 (N_13810,N_9621,N_9890);
and U13811 (N_13811,N_11938,N_9613);
and U13812 (N_13812,N_9432,N_11499);
or U13813 (N_13813,N_11666,N_11247);
and U13814 (N_13814,N_10408,N_10187);
xnor U13815 (N_13815,N_10811,N_9128);
and U13816 (N_13816,N_11810,N_11676);
nor U13817 (N_13817,N_11925,N_10928);
or U13818 (N_13818,N_9782,N_10272);
xor U13819 (N_13819,N_9094,N_11260);
nand U13820 (N_13820,N_10439,N_11592);
nand U13821 (N_13821,N_11249,N_11021);
and U13822 (N_13822,N_9037,N_10475);
nand U13823 (N_13823,N_11023,N_10955);
and U13824 (N_13824,N_9294,N_9997);
and U13825 (N_13825,N_9024,N_9484);
and U13826 (N_13826,N_11668,N_9336);
or U13827 (N_13827,N_11813,N_10873);
nand U13828 (N_13828,N_9040,N_10804);
nand U13829 (N_13829,N_10452,N_11524);
nor U13830 (N_13830,N_10563,N_11187);
and U13831 (N_13831,N_10033,N_10057);
nor U13832 (N_13832,N_11367,N_11969);
nand U13833 (N_13833,N_9515,N_10635);
or U13834 (N_13834,N_9182,N_9597);
nor U13835 (N_13835,N_9024,N_9253);
and U13836 (N_13836,N_9362,N_11999);
xor U13837 (N_13837,N_11834,N_9987);
nor U13838 (N_13838,N_9237,N_11235);
nand U13839 (N_13839,N_9614,N_10915);
xor U13840 (N_13840,N_10688,N_11063);
nand U13841 (N_13841,N_11094,N_11980);
or U13842 (N_13842,N_10029,N_9500);
and U13843 (N_13843,N_10420,N_9419);
nand U13844 (N_13844,N_10444,N_9691);
nor U13845 (N_13845,N_9124,N_10225);
nand U13846 (N_13846,N_11305,N_9353);
nand U13847 (N_13847,N_11653,N_9984);
or U13848 (N_13848,N_11051,N_11184);
nand U13849 (N_13849,N_9788,N_11384);
nor U13850 (N_13850,N_9318,N_11058);
nand U13851 (N_13851,N_10268,N_11304);
nand U13852 (N_13852,N_11445,N_10874);
nand U13853 (N_13853,N_9465,N_10989);
or U13854 (N_13854,N_11823,N_9978);
nand U13855 (N_13855,N_11408,N_9691);
or U13856 (N_13856,N_11173,N_9435);
or U13857 (N_13857,N_10100,N_9525);
or U13858 (N_13858,N_11370,N_9735);
and U13859 (N_13859,N_9007,N_11989);
nor U13860 (N_13860,N_10545,N_9565);
nand U13861 (N_13861,N_11349,N_11920);
or U13862 (N_13862,N_9753,N_9795);
and U13863 (N_13863,N_11758,N_10035);
or U13864 (N_13864,N_11346,N_10008);
nor U13865 (N_13865,N_11803,N_9149);
or U13866 (N_13866,N_10927,N_9742);
or U13867 (N_13867,N_9317,N_9851);
nand U13868 (N_13868,N_9717,N_9490);
nand U13869 (N_13869,N_10443,N_9043);
nand U13870 (N_13870,N_9033,N_10605);
nand U13871 (N_13871,N_10726,N_11984);
and U13872 (N_13872,N_10627,N_9934);
or U13873 (N_13873,N_11011,N_10175);
or U13874 (N_13874,N_9175,N_11358);
or U13875 (N_13875,N_11141,N_10031);
nor U13876 (N_13876,N_11893,N_9177);
nor U13877 (N_13877,N_10626,N_11572);
nand U13878 (N_13878,N_11723,N_11425);
nor U13879 (N_13879,N_9185,N_9252);
nor U13880 (N_13880,N_10245,N_10325);
nand U13881 (N_13881,N_9592,N_9049);
xor U13882 (N_13882,N_9889,N_9800);
xnor U13883 (N_13883,N_9278,N_11666);
or U13884 (N_13884,N_9177,N_11154);
nand U13885 (N_13885,N_10983,N_9840);
nand U13886 (N_13886,N_11215,N_9344);
or U13887 (N_13887,N_10166,N_9864);
nand U13888 (N_13888,N_11904,N_10075);
nand U13889 (N_13889,N_9679,N_10806);
nand U13890 (N_13890,N_9913,N_10718);
and U13891 (N_13891,N_10011,N_9563);
nand U13892 (N_13892,N_9409,N_10688);
or U13893 (N_13893,N_10912,N_11438);
and U13894 (N_13894,N_10140,N_10915);
nor U13895 (N_13895,N_9682,N_11475);
nand U13896 (N_13896,N_10909,N_11250);
nand U13897 (N_13897,N_9224,N_11796);
xor U13898 (N_13898,N_11791,N_11959);
nor U13899 (N_13899,N_9701,N_9442);
or U13900 (N_13900,N_10129,N_9024);
xnor U13901 (N_13901,N_10638,N_11350);
nor U13902 (N_13902,N_11325,N_9434);
nand U13903 (N_13903,N_10033,N_9446);
and U13904 (N_13904,N_11972,N_9949);
or U13905 (N_13905,N_9830,N_10271);
nand U13906 (N_13906,N_11548,N_10948);
nor U13907 (N_13907,N_11598,N_9871);
nor U13908 (N_13908,N_9327,N_10753);
xnor U13909 (N_13909,N_10868,N_10067);
and U13910 (N_13910,N_9006,N_10239);
nand U13911 (N_13911,N_11011,N_10273);
nor U13912 (N_13912,N_10913,N_9586);
nor U13913 (N_13913,N_10676,N_10626);
xor U13914 (N_13914,N_11439,N_10881);
or U13915 (N_13915,N_10999,N_9691);
nor U13916 (N_13916,N_11381,N_11970);
or U13917 (N_13917,N_9212,N_11530);
nor U13918 (N_13918,N_10145,N_9117);
nand U13919 (N_13919,N_11822,N_11693);
nand U13920 (N_13920,N_11326,N_10547);
and U13921 (N_13921,N_9538,N_9602);
nor U13922 (N_13922,N_10963,N_11552);
nand U13923 (N_13923,N_11185,N_11424);
and U13924 (N_13924,N_9460,N_9734);
and U13925 (N_13925,N_9145,N_11680);
xnor U13926 (N_13926,N_9260,N_11023);
and U13927 (N_13927,N_9022,N_11808);
and U13928 (N_13928,N_9093,N_11451);
nand U13929 (N_13929,N_10672,N_10333);
or U13930 (N_13930,N_10108,N_11483);
or U13931 (N_13931,N_10514,N_10236);
and U13932 (N_13932,N_10747,N_9476);
or U13933 (N_13933,N_10743,N_9151);
nor U13934 (N_13934,N_11569,N_11516);
or U13935 (N_13935,N_9286,N_11308);
nor U13936 (N_13936,N_11333,N_9723);
nor U13937 (N_13937,N_9372,N_11519);
nand U13938 (N_13938,N_11922,N_10115);
or U13939 (N_13939,N_11866,N_10646);
or U13940 (N_13940,N_10720,N_10762);
nand U13941 (N_13941,N_10355,N_10863);
and U13942 (N_13942,N_9896,N_11569);
nand U13943 (N_13943,N_11786,N_10924);
or U13944 (N_13944,N_9752,N_10769);
nand U13945 (N_13945,N_11711,N_9291);
nor U13946 (N_13946,N_11646,N_9801);
and U13947 (N_13947,N_10191,N_9425);
nand U13948 (N_13948,N_11496,N_9427);
or U13949 (N_13949,N_11899,N_10634);
xnor U13950 (N_13950,N_11033,N_9586);
nand U13951 (N_13951,N_10221,N_11894);
nor U13952 (N_13952,N_11651,N_9704);
nand U13953 (N_13953,N_10316,N_11875);
or U13954 (N_13954,N_11102,N_9114);
nor U13955 (N_13955,N_10949,N_10203);
or U13956 (N_13956,N_9233,N_10025);
and U13957 (N_13957,N_10554,N_11693);
xnor U13958 (N_13958,N_10545,N_9051);
nor U13959 (N_13959,N_9941,N_10371);
and U13960 (N_13960,N_11027,N_11016);
nand U13961 (N_13961,N_9503,N_11342);
nor U13962 (N_13962,N_11717,N_10226);
nand U13963 (N_13963,N_11162,N_9254);
or U13964 (N_13964,N_9706,N_9745);
nand U13965 (N_13965,N_11266,N_11585);
nor U13966 (N_13966,N_10770,N_10867);
nand U13967 (N_13967,N_9132,N_9691);
xor U13968 (N_13968,N_10658,N_9837);
and U13969 (N_13969,N_11027,N_11794);
and U13970 (N_13970,N_10123,N_11826);
nor U13971 (N_13971,N_9276,N_11676);
and U13972 (N_13972,N_9733,N_10857);
and U13973 (N_13973,N_10934,N_11049);
nor U13974 (N_13974,N_11640,N_10282);
xnor U13975 (N_13975,N_10998,N_10407);
or U13976 (N_13976,N_9078,N_9366);
nor U13977 (N_13977,N_9057,N_11110);
or U13978 (N_13978,N_11584,N_10200);
nor U13979 (N_13979,N_10744,N_11839);
nand U13980 (N_13980,N_11247,N_10516);
or U13981 (N_13981,N_9499,N_9953);
nand U13982 (N_13982,N_11210,N_10941);
xor U13983 (N_13983,N_10275,N_9111);
nand U13984 (N_13984,N_10182,N_11717);
nor U13985 (N_13985,N_10009,N_11561);
nor U13986 (N_13986,N_9877,N_9396);
nand U13987 (N_13987,N_9131,N_11913);
nor U13988 (N_13988,N_10368,N_10695);
or U13989 (N_13989,N_10846,N_9658);
nor U13990 (N_13990,N_11641,N_11944);
nand U13991 (N_13991,N_9523,N_10577);
or U13992 (N_13992,N_9581,N_9139);
or U13993 (N_13993,N_10613,N_9513);
or U13994 (N_13994,N_11260,N_9457);
xnor U13995 (N_13995,N_11498,N_9614);
and U13996 (N_13996,N_11771,N_11998);
and U13997 (N_13997,N_10233,N_9337);
and U13998 (N_13998,N_11023,N_11895);
and U13999 (N_13999,N_11981,N_9863);
and U14000 (N_14000,N_9786,N_9279);
or U14001 (N_14001,N_10057,N_11013);
and U14002 (N_14002,N_11591,N_11300);
nand U14003 (N_14003,N_9243,N_11571);
nor U14004 (N_14004,N_11426,N_10696);
nand U14005 (N_14005,N_11390,N_10421);
and U14006 (N_14006,N_9759,N_11510);
nor U14007 (N_14007,N_9352,N_11248);
nand U14008 (N_14008,N_10753,N_10277);
and U14009 (N_14009,N_10831,N_11151);
and U14010 (N_14010,N_9149,N_9216);
and U14011 (N_14011,N_9137,N_11364);
or U14012 (N_14012,N_11590,N_10454);
or U14013 (N_14013,N_11414,N_9437);
nor U14014 (N_14014,N_9658,N_9853);
and U14015 (N_14015,N_11221,N_9092);
and U14016 (N_14016,N_11949,N_10118);
nor U14017 (N_14017,N_9267,N_11101);
or U14018 (N_14018,N_11686,N_10913);
and U14019 (N_14019,N_11782,N_10430);
and U14020 (N_14020,N_11251,N_11186);
and U14021 (N_14021,N_9883,N_11285);
and U14022 (N_14022,N_10894,N_11694);
nor U14023 (N_14023,N_9515,N_9495);
xnor U14024 (N_14024,N_11788,N_10888);
or U14025 (N_14025,N_11814,N_9780);
nor U14026 (N_14026,N_10574,N_9543);
xor U14027 (N_14027,N_11064,N_10565);
and U14028 (N_14028,N_10792,N_11196);
nand U14029 (N_14029,N_11847,N_10701);
nand U14030 (N_14030,N_11167,N_9575);
nand U14031 (N_14031,N_9294,N_10554);
and U14032 (N_14032,N_10231,N_10991);
or U14033 (N_14033,N_10734,N_9261);
nand U14034 (N_14034,N_10422,N_10570);
nor U14035 (N_14035,N_9388,N_9025);
or U14036 (N_14036,N_11076,N_10802);
nor U14037 (N_14037,N_11241,N_11334);
and U14038 (N_14038,N_10050,N_10018);
and U14039 (N_14039,N_9208,N_11732);
nand U14040 (N_14040,N_11812,N_9161);
and U14041 (N_14041,N_9786,N_11263);
nand U14042 (N_14042,N_9668,N_11382);
nor U14043 (N_14043,N_11013,N_10331);
and U14044 (N_14044,N_10845,N_11945);
nand U14045 (N_14045,N_11626,N_10616);
or U14046 (N_14046,N_10394,N_10133);
or U14047 (N_14047,N_11062,N_9906);
nor U14048 (N_14048,N_9045,N_10658);
and U14049 (N_14049,N_11797,N_9578);
and U14050 (N_14050,N_11199,N_10792);
or U14051 (N_14051,N_11707,N_10442);
nor U14052 (N_14052,N_11130,N_11745);
and U14053 (N_14053,N_11804,N_10614);
or U14054 (N_14054,N_10685,N_9327);
nor U14055 (N_14055,N_11856,N_10644);
nor U14056 (N_14056,N_9675,N_10068);
nand U14057 (N_14057,N_11639,N_11182);
and U14058 (N_14058,N_10904,N_10330);
or U14059 (N_14059,N_11001,N_10517);
nor U14060 (N_14060,N_11510,N_10732);
nand U14061 (N_14061,N_11501,N_11360);
and U14062 (N_14062,N_11752,N_11641);
nand U14063 (N_14063,N_9406,N_9783);
nor U14064 (N_14064,N_11782,N_11767);
nand U14065 (N_14065,N_9392,N_11869);
and U14066 (N_14066,N_9693,N_11431);
or U14067 (N_14067,N_10598,N_9441);
or U14068 (N_14068,N_11739,N_10713);
and U14069 (N_14069,N_11015,N_9811);
nor U14070 (N_14070,N_11690,N_10122);
or U14071 (N_14071,N_10474,N_11118);
xnor U14072 (N_14072,N_11293,N_11383);
or U14073 (N_14073,N_11160,N_10643);
or U14074 (N_14074,N_10391,N_9527);
or U14075 (N_14075,N_11046,N_10473);
xnor U14076 (N_14076,N_11656,N_9413);
and U14077 (N_14077,N_9338,N_11298);
xnor U14078 (N_14078,N_11580,N_9674);
nor U14079 (N_14079,N_9631,N_11236);
nor U14080 (N_14080,N_10502,N_9678);
and U14081 (N_14081,N_11149,N_9560);
and U14082 (N_14082,N_10523,N_10833);
nor U14083 (N_14083,N_10351,N_9441);
nor U14084 (N_14084,N_10880,N_10487);
and U14085 (N_14085,N_9765,N_9508);
nor U14086 (N_14086,N_11281,N_11243);
or U14087 (N_14087,N_9240,N_9432);
nand U14088 (N_14088,N_10351,N_9461);
nor U14089 (N_14089,N_10806,N_11614);
and U14090 (N_14090,N_11928,N_11529);
xor U14091 (N_14091,N_10513,N_11522);
nor U14092 (N_14092,N_10481,N_11063);
and U14093 (N_14093,N_10523,N_9992);
nand U14094 (N_14094,N_9683,N_9687);
xnor U14095 (N_14095,N_9321,N_11506);
nor U14096 (N_14096,N_9214,N_11734);
nand U14097 (N_14097,N_11604,N_11855);
xor U14098 (N_14098,N_9809,N_9436);
nor U14099 (N_14099,N_10379,N_11808);
xor U14100 (N_14100,N_10277,N_11268);
nand U14101 (N_14101,N_11833,N_11993);
nand U14102 (N_14102,N_11750,N_10627);
nor U14103 (N_14103,N_9294,N_9274);
nand U14104 (N_14104,N_10129,N_11215);
and U14105 (N_14105,N_11387,N_11192);
nor U14106 (N_14106,N_10675,N_11728);
nand U14107 (N_14107,N_11932,N_9800);
xor U14108 (N_14108,N_9119,N_10541);
xnor U14109 (N_14109,N_11470,N_11011);
nor U14110 (N_14110,N_10764,N_9153);
nand U14111 (N_14111,N_10065,N_11350);
xor U14112 (N_14112,N_11396,N_10357);
and U14113 (N_14113,N_10085,N_11682);
nand U14114 (N_14114,N_9197,N_10574);
nand U14115 (N_14115,N_9425,N_10344);
and U14116 (N_14116,N_11325,N_9997);
nor U14117 (N_14117,N_10487,N_9717);
nand U14118 (N_14118,N_11548,N_9475);
or U14119 (N_14119,N_11010,N_9692);
and U14120 (N_14120,N_10109,N_9725);
and U14121 (N_14121,N_10928,N_9661);
nand U14122 (N_14122,N_9779,N_9681);
or U14123 (N_14123,N_9623,N_10841);
nand U14124 (N_14124,N_11518,N_11245);
and U14125 (N_14125,N_10090,N_10945);
nand U14126 (N_14126,N_10212,N_11955);
or U14127 (N_14127,N_9368,N_9081);
nand U14128 (N_14128,N_9545,N_11098);
nor U14129 (N_14129,N_9880,N_11097);
nor U14130 (N_14130,N_11406,N_9568);
nor U14131 (N_14131,N_11227,N_9701);
and U14132 (N_14132,N_9469,N_10697);
nor U14133 (N_14133,N_9116,N_9788);
nor U14134 (N_14134,N_10209,N_11501);
nand U14135 (N_14135,N_11807,N_9366);
and U14136 (N_14136,N_11641,N_10129);
nor U14137 (N_14137,N_9557,N_10303);
and U14138 (N_14138,N_9934,N_10897);
and U14139 (N_14139,N_11591,N_10678);
nor U14140 (N_14140,N_10449,N_11127);
nand U14141 (N_14141,N_9658,N_10821);
nand U14142 (N_14142,N_10234,N_11148);
nor U14143 (N_14143,N_10937,N_11192);
or U14144 (N_14144,N_9946,N_11995);
nand U14145 (N_14145,N_11824,N_10201);
and U14146 (N_14146,N_10483,N_9604);
and U14147 (N_14147,N_9215,N_10897);
xnor U14148 (N_14148,N_10582,N_9003);
nor U14149 (N_14149,N_10902,N_11169);
and U14150 (N_14150,N_10951,N_11178);
or U14151 (N_14151,N_11469,N_10130);
and U14152 (N_14152,N_10144,N_10205);
or U14153 (N_14153,N_11695,N_9669);
xor U14154 (N_14154,N_9641,N_10256);
and U14155 (N_14155,N_10623,N_9879);
nand U14156 (N_14156,N_9443,N_11756);
nand U14157 (N_14157,N_11376,N_11838);
or U14158 (N_14158,N_9967,N_9304);
or U14159 (N_14159,N_11799,N_10201);
or U14160 (N_14160,N_10279,N_10153);
xnor U14161 (N_14161,N_9478,N_11005);
xnor U14162 (N_14162,N_10872,N_11965);
xor U14163 (N_14163,N_9214,N_10784);
or U14164 (N_14164,N_10373,N_10313);
or U14165 (N_14165,N_9759,N_11856);
and U14166 (N_14166,N_10396,N_11504);
nor U14167 (N_14167,N_9123,N_11866);
and U14168 (N_14168,N_11156,N_9886);
nor U14169 (N_14169,N_10921,N_11674);
and U14170 (N_14170,N_11494,N_11177);
nor U14171 (N_14171,N_9521,N_10683);
nor U14172 (N_14172,N_11456,N_9104);
nor U14173 (N_14173,N_10437,N_10118);
or U14174 (N_14174,N_10475,N_9717);
xnor U14175 (N_14175,N_9368,N_11852);
nand U14176 (N_14176,N_11045,N_9247);
nor U14177 (N_14177,N_10280,N_11861);
or U14178 (N_14178,N_10060,N_11500);
nand U14179 (N_14179,N_11645,N_9746);
xnor U14180 (N_14180,N_9144,N_9394);
and U14181 (N_14181,N_11610,N_11692);
nand U14182 (N_14182,N_11717,N_11278);
xor U14183 (N_14183,N_11578,N_11548);
nor U14184 (N_14184,N_10347,N_9552);
nand U14185 (N_14185,N_9421,N_9166);
nor U14186 (N_14186,N_9113,N_9349);
xnor U14187 (N_14187,N_11725,N_11080);
xor U14188 (N_14188,N_10929,N_10157);
xor U14189 (N_14189,N_11610,N_9625);
or U14190 (N_14190,N_10935,N_9625);
and U14191 (N_14191,N_11147,N_9739);
and U14192 (N_14192,N_11388,N_9045);
or U14193 (N_14193,N_11898,N_10058);
nand U14194 (N_14194,N_11979,N_10921);
nand U14195 (N_14195,N_11173,N_9308);
and U14196 (N_14196,N_9270,N_9866);
nand U14197 (N_14197,N_9191,N_11689);
and U14198 (N_14198,N_11938,N_10684);
or U14199 (N_14199,N_10078,N_10902);
and U14200 (N_14200,N_10580,N_11412);
nand U14201 (N_14201,N_10008,N_11374);
nor U14202 (N_14202,N_9266,N_9559);
or U14203 (N_14203,N_11487,N_9247);
or U14204 (N_14204,N_11185,N_11976);
nand U14205 (N_14205,N_11593,N_11441);
nor U14206 (N_14206,N_10397,N_9523);
nand U14207 (N_14207,N_11914,N_9756);
nand U14208 (N_14208,N_11680,N_9494);
nand U14209 (N_14209,N_11921,N_9083);
and U14210 (N_14210,N_11304,N_10771);
or U14211 (N_14211,N_11761,N_9200);
and U14212 (N_14212,N_10694,N_9381);
xnor U14213 (N_14213,N_11907,N_10215);
nor U14214 (N_14214,N_11543,N_9658);
xnor U14215 (N_14215,N_9926,N_11731);
nand U14216 (N_14216,N_10015,N_9589);
or U14217 (N_14217,N_11517,N_9541);
or U14218 (N_14218,N_9093,N_11580);
nand U14219 (N_14219,N_10247,N_9031);
nor U14220 (N_14220,N_11077,N_11374);
nor U14221 (N_14221,N_9960,N_9959);
nand U14222 (N_14222,N_11920,N_11432);
nand U14223 (N_14223,N_10558,N_11618);
nor U14224 (N_14224,N_11227,N_10704);
and U14225 (N_14225,N_9916,N_11965);
or U14226 (N_14226,N_9417,N_11048);
or U14227 (N_14227,N_11617,N_11996);
or U14228 (N_14228,N_9635,N_9732);
nand U14229 (N_14229,N_10959,N_10563);
and U14230 (N_14230,N_9938,N_9671);
xnor U14231 (N_14231,N_11367,N_11029);
nor U14232 (N_14232,N_9963,N_9663);
and U14233 (N_14233,N_11973,N_10598);
and U14234 (N_14234,N_11396,N_9313);
and U14235 (N_14235,N_9988,N_10865);
or U14236 (N_14236,N_9009,N_10145);
nor U14237 (N_14237,N_11784,N_9866);
nor U14238 (N_14238,N_11962,N_10570);
or U14239 (N_14239,N_10600,N_11170);
and U14240 (N_14240,N_10196,N_10179);
and U14241 (N_14241,N_10220,N_9564);
and U14242 (N_14242,N_10551,N_11749);
nor U14243 (N_14243,N_9312,N_9567);
nor U14244 (N_14244,N_11043,N_9489);
xnor U14245 (N_14245,N_11713,N_11880);
xnor U14246 (N_14246,N_11792,N_10252);
and U14247 (N_14247,N_10287,N_10539);
or U14248 (N_14248,N_11347,N_10590);
or U14249 (N_14249,N_9647,N_10092);
and U14250 (N_14250,N_9908,N_11080);
or U14251 (N_14251,N_11351,N_11686);
nand U14252 (N_14252,N_9610,N_10359);
nor U14253 (N_14253,N_9444,N_10508);
nand U14254 (N_14254,N_10946,N_10856);
or U14255 (N_14255,N_9133,N_10800);
and U14256 (N_14256,N_9512,N_11578);
nand U14257 (N_14257,N_11218,N_10151);
nor U14258 (N_14258,N_10115,N_10511);
nand U14259 (N_14259,N_9944,N_11342);
or U14260 (N_14260,N_9973,N_9265);
or U14261 (N_14261,N_9157,N_10477);
nor U14262 (N_14262,N_10236,N_9473);
nor U14263 (N_14263,N_10573,N_11591);
nand U14264 (N_14264,N_9052,N_11939);
nor U14265 (N_14265,N_10115,N_10554);
xnor U14266 (N_14266,N_11531,N_9880);
nor U14267 (N_14267,N_11495,N_9556);
xnor U14268 (N_14268,N_10911,N_10982);
nand U14269 (N_14269,N_10587,N_11092);
and U14270 (N_14270,N_10251,N_9913);
and U14271 (N_14271,N_11701,N_9538);
or U14272 (N_14272,N_9995,N_11936);
nand U14273 (N_14273,N_10454,N_11357);
or U14274 (N_14274,N_10942,N_10533);
and U14275 (N_14275,N_9152,N_9483);
or U14276 (N_14276,N_11885,N_10458);
or U14277 (N_14277,N_9459,N_9915);
nor U14278 (N_14278,N_10262,N_10436);
nor U14279 (N_14279,N_9993,N_10325);
nor U14280 (N_14280,N_11009,N_11805);
or U14281 (N_14281,N_10012,N_10131);
and U14282 (N_14282,N_10055,N_11285);
xnor U14283 (N_14283,N_9824,N_10042);
or U14284 (N_14284,N_9179,N_9485);
and U14285 (N_14285,N_9086,N_11829);
or U14286 (N_14286,N_10193,N_9571);
or U14287 (N_14287,N_9161,N_10128);
or U14288 (N_14288,N_10367,N_11197);
nor U14289 (N_14289,N_11699,N_10583);
nand U14290 (N_14290,N_11723,N_11360);
nand U14291 (N_14291,N_9901,N_10365);
nor U14292 (N_14292,N_9891,N_10683);
or U14293 (N_14293,N_11932,N_11850);
nor U14294 (N_14294,N_11873,N_10304);
nor U14295 (N_14295,N_10239,N_10571);
nor U14296 (N_14296,N_9800,N_10449);
nor U14297 (N_14297,N_10298,N_10159);
nor U14298 (N_14298,N_10735,N_9364);
and U14299 (N_14299,N_11432,N_11434);
and U14300 (N_14300,N_10252,N_10422);
nand U14301 (N_14301,N_9025,N_11990);
nand U14302 (N_14302,N_11481,N_11658);
and U14303 (N_14303,N_11089,N_9248);
nor U14304 (N_14304,N_10133,N_10302);
and U14305 (N_14305,N_10830,N_9358);
xor U14306 (N_14306,N_11574,N_9156);
nand U14307 (N_14307,N_10899,N_10608);
nor U14308 (N_14308,N_11454,N_10518);
nor U14309 (N_14309,N_9271,N_11506);
and U14310 (N_14310,N_10850,N_11646);
and U14311 (N_14311,N_11525,N_11285);
and U14312 (N_14312,N_11075,N_11203);
nor U14313 (N_14313,N_11756,N_11422);
nor U14314 (N_14314,N_10943,N_11429);
nand U14315 (N_14315,N_10283,N_9592);
nand U14316 (N_14316,N_9412,N_10507);
nor U14317 (N_14317,N_10043,N_11832);
nand U14318 (N_14318,N_9565,N_11032);
or U14319 (N_14319,N_10585,N_9593);
or U14320 (N_14320,N_10549,N_11970);
nor U14321 (N_14321,N_9921,N_9447);
nand U14322 (N_14322,N_11278,N_11054);
nor U14323 (N_14323,N_9738,N_10580);
and U14324 (N_14324,N_10095,N_10679);
and U14325 (N_14325,N_9255,N_11102);
and U14326 (N_14326,N_11138,N_9634);
and U14327 (N_14327,N_11515,N_9679);
or U14328 (N_14328,N_9013,N_9953);
nand U14329 (N_14329,N_9512,N_11835);
or U14330 (N_14330,N_11482,N_10049);
nor U14331 (N_14331,N_10644,N_11075);
nor U14332 (N_14332,N_10936,N_10329);
and U14333 (N_14333,N_9195,N_9794);
xor U14334 (N_14334,N_11691,N_10271);
nor U14335 (N_14335,N_10882,N_10915);
xor U14336 (N_14336,N_10884,N_11760);
nor U14337 (N_14337,N_11517,N_9883);
nand U14338 (N_14338,N_9828,N_10638);
nor U14339 (N_14339,N_10305,N_10921);
nor U14340 (N_14340,N_11798,N_10866);
or U14341 (N_14341,N_9404,N_10876);
nor U14342 (N_14342,N_11250,N_10251);
nor U14343 (N_14343,N_11854,N_11646);
nor U14344 (N_14344,N_11503,N_11428);
and U14345 (N_14345,N_9234,N_9917);
nor U14346 (N_14346,N_10433,N_9789);
nand U14347 (N_14347,N_10525,N_9161);
and U14348 (N_14348,N_10092,N_11278);
nor U14349 (N_14349,N_11426,N_9738);
nand U14350 (N_14350,N_11475,N_9415);
or U14351 (N_14351,N_10240,N_11302);
nor U14352 (N_14352,N_11555,N_11592);
and U14353 (N_14353,N_11079,N_11716);
xnor U14354 (N_14354,N_10654,N_10082);
xor U14355 (N_14355,N_10047,N_9615);
xnor U14356 (N_14356,N_10363,N_10769);
or U14357 (N_14357,N_11346,N_9145);
nor U14358 (N_14358,N_10797,N_11577);
or U14359 (N_14359,N_10032,N_10121);
or U14360 (N_14360,N_11057,N_10297);
nor U14361 (N_14361,N_10187,N_9109);
or U14362 (N_14362,N_9776,N_10484);
and U14363 (N_14363,N_11625,N_10421);
nor U14364 (N_14364,N_10208,N_9242);
nand U14365 (N_14365,N_10067,N_11157);
and U14366 (N_14366,N_11405,N_10152);
nand U14367 (N_14367,N_10234,N_9897);
or U14368 (N_14368,N_9441,N_11664);
nor U14369 (N_14369,N_11022,N_10783);
nor U14370 (N_14370,N_11735,N_11748);
or U14371 (N_14371,N_10211,N_11481);
or U14372 (N_14372,N_9740,N_11354);
and U14373 (N_14373,N_11132,N_9759);
or U14374 (N_14374,N_10359,N_9386);
and U14375 (N_14375,N_9211,N_11203);
nand U14376 (N_14376,N_9701,N_11199);
or U14377 (N_14377,N_11682,N_11262);
or U14378 (N_14378,N_10119,N_11792);
nor U14379 (N_14379,N_10407,N_9701);
or U14380 (N_14380,N_11231,N_9624);
or U14381 (N_14381,N_11936,N_11035);
and U14382 (N_14382,N_11780,N_11072);
nor U14383 (N_14383,N_9738,N_9386);
and U14384 (N_14384,N_9675,N_9476);
nand U14385 (N_14385,N_10226,N_11112);
nand U14386 (N_14386,N_9006,N_10985);
nor U14387 (N_14387,N_10549,N_9015);
and U14388 (N_14388,N_11626,N_11782);
nor U14389 (N_14389,N_10513,N_10690);
or U14390 (N_14390,N_9090,N_10073);
and U14391 (N_14391,N_11210,N_11302);
or U14392 (N_14392,N_10034,N_11140);
nand U14393 (N_14393,N_11413,N_9572);
nand U14394 (N_14394,N_9880,N_10878);
nand U14395 (N_14395,N_9135,N_10560);
nor U14396 (N_14396,N_10360,N_10629);
and U14397 (N_14397,N_9675,N_9112);
or U14398 (N_14398,N_10495,N_11925);
or U14399 (N_14399,N_11387,N_9511);
nor U14400 (N_14400,N_10442,N_10668);
nor U14401 (N_14401,N_9112,N_11145);
nor U14402 (N_14402,N_10749,N_10176);
xnor U14403 (N_14403,N_11423,N_11104);
nand U14404 (N_14404,N_11481,N_9853);
and U14405 (N_14405,N_10136,N_10607);
and U14406 (N_14406,N_9641,N_9137);
nand U14407 (N_14407,N_9167,N_10562);
nor U14408 (N_14408,N_11830,N_11552);
nand U14409 (N_14409,N_10089,N_11171);
or U14410 (N_14410,N_10220,N_10743);
nand U14411 (N_14411,N_10717,N_10208);
or U14412 (N_14412,N_9281,N_10361);
nor U14413 (N_14413,N_11522,N_9233);
nor U14414 (N_14414,N_10918,N_10248);
nand U14415 (N_14415,N_9269,N_10200);
nand U14416 (N_14416,N_11346,N_11266);
or U14417 (N_14417,N_11620,N_11743);
and U14418 (N_14418,N_11549,N_9320);
xnor U14419 (N_14419,N_9971,N_11058);
nand U14420 (N_14420,N_10992,N_11613);
nand U14421 (N_14421,N_10123,N_10777);
or U14422 (N_14422,N_9823,N_10289);
and U14423 (N_14423,N_10309,N_10360);
and U14424 (N_14424,N_10911,N_11901);
or U14425 (N_14425,N_9732,N_11633);
nand U14426 (N_14426,N_10745,N_9742);
nor U14427 (N_14427,N_9237,N_9912);
or U14428 (N_14428,N_10917,N_11493);
and U14429 (N_14429,N_10722,N_10053);
or U14430 (N_14430,N_9894,N_9720);
or U14431 (N_14431,N_9574,N_11643);
or U14432 (N_14432,N_9861,N_9655);
xnor U14433 (N_14433,N_10317,N_9004);
nor U14434 (N_14434,N_9404,N_11568);
nor U14435 (N_14435,N_10872,N_10492);
and U14436 (N_14436,N_9656,N_11830);
or U14437 (N_14437,N_11733,N_9353);
or U14438 (N_14438,N_9906,N_11819);
or U14439 (N_14439,N_11047,N_10623);
nand U14440 (N_14440,N_10927,N_11693);
nand U14441 (N_14441,N_11569,N_11927);
or U14442 (N_14442,N_10404,N_10859);
and U14443 (N_14443,N_10585,N_11013);
nor U14444 (N_14444,N_11831,N_9056);
nand U14445 (N_14445,N_10529,N_10272);
or U14446 (N_14446,N_10701,N_10410);
xnor U14447 (N_14447,N_10973,N_9345);
and U14448 (N_14448,N_10979,N_9202);
xnor U14449 (N_14449,N_10047,N_11306);
nor U14450 (N_14450,N_11343,N_9926);
or U14451 (N_14451,N_9051,N_9289);
and U14452 (N_14452,N_9687,N_11170);
and U14453 (N_14453,N_9371,N_10648);
nor U14454 (N_14454,N_9871,N_11130);
and U14455 (N_14455,N_9532,N_9120);
and U14456 (N_14456,N_10957,N_9572);
nand U14457 (N_14457,N_10051,N_10954);
nand U14458 (N_14458,N_10819,N_11593);
nor U14459 (N_14459,N_11065,N_10973);
and U14460 (N_14460,N_11534,N_10704);
xnor U14461 (N_14461,N_11719,N_10966);
nor U14462 (N_14462,N_9824,N_10174);
and U14463 (N_14463,N_9502,N_10621);
xnor U14464 (N_14464,N_9441,N_9169);
nor U14465 (N_14465,N_9435,N_11755);
or U14466 (N_14466,N_10798,N_11800);
or U14467 (N_14467,N_10735,N_11189);
xnor U14468 (N_14468,N_10501,N_11908);
and U14469 (N_14469,N_10397,N_11881);
or U14470 (N_14470,N_11596,N_11103);
and U14471 (N_14471,N_10822,N_10938);
or U14472 (N_14472,N_9502,N_10189);
or U14473 (N_14473,N_9784,N_10739);
or U14474 (N_14474,N_11816,N_9530);
and U14475 (N_14475,N_11774,N_9713);
nand U14476 (N_14476,N_10240,N_9982);
and U14477 (N_14477,N_9715,N_11489);
nor U14478 (N_14478,N_10708,N_10003);
xnor U14479 (N_14479,N_10225,N_11954);
xor U14480 (N_14480,N_9162,N_9558);
nand U14481 (N_14481,N_9569,N_10597);
nor U14482 (N_14482,N_11532,N_9481);
nand U14483 (N_14483,N_11228,N_11338);
nor U14484 (N_14484,N_9591,N_11492);
nand U14485 (N_14485,N_9197,N_10074);
or U14486 (N_14486,N_10849,N_9249);
and U14487 (N_14487,N_10273,N_10292);
or U14488 (N_14488,N_11976,N_11357);
nor U14489 (N_14489,N_11266,N_11933);
nand U14490 (N_14490,N_11165,N_11397);
nand U14491 (N_14491,N_11113,N_10256);
and U14492 (N_14492,N_10459,N_11325);
or U14493 (N_14493,N_9368,N_9216);
or U14494 (N_14494,N_10873,N_11844);
nand U14495 (N_14495,N_9492,N_10259);
xnor U14496 (N_14496,N_9769,N_9233);
nand U14497 (N_14497,N_10020,N_9986);
nor U14498 (N_14498,N_11208,N_11310);
or U14499 (N_14499,N_10366,N_11875);
nor U14500 (N_14500,N_11165,N_11439);
nor U14501 (N_14501,N_11270,N_10123);
nor U14502 (N_14502,N_9706,N_11455);
or U14503 (N_14503,N_9331,N_10583);
nor U14504 (N_14504,N_9019,N_9851);
and U14505 (N_14505,N_11456,N_10203);
nor U14506 (N_14506,N_9796,N_9080);
xnor U14507 (N_14507,N_9815,N_9207);
nand U14508 (N_14508,N_11923,N_11694);
nand U14509 (N_14509,N_10227,N_10553);
nand U14510 (N_14510,N_11361,N_10716);
nand U14511 (N_14511,N_9717,N_11411);
nor U14512 (N_14512,N_10519,N_11542);
nor U14513 (N_14513,N_10346,N_11494);
and U14514 (N_14514,N_11057,N_9969);
nand U14515 (N_14515,N_10975,N_10100);
xnor U14516 (N_14516,N_10007,N_9712);
nand U14517 (N_14517,N_11641,N_9435);
nand U14518 (N_14518,N_10270,N_9676);
xnor U14519 (N_14519,N_11153,N_11620);
or U14520 (N_14520,N_10579,N_9740);
nand U14521 (N_14521,N_9027,N_11331);
nand U14522 (N_14522,N_9425,N_10862);
and U14523 (N_14523,N_11514,N_11918);
and U14524 (N_14524,N_10216,N_9580);
or U14525 (N_14525,N_11439,N_9764);
nor U14526 (N_14526,N_9729,N_11382);
nor U14527 (N_14527,N_11073,N_10906);
or U14528 (N_14528,N_10691,N_11559);
and U14529 (N_14529,N_10732,N_10473);
or U14530 (N_14530,N_10898,N_11902);
and U14531 (N_14531,N_11773,N_11764);
nor U14532 (N_14532,N_11660,N_10743);
or U14533 (N_14533,N_10010,N_9152);
nand U14534 (N_14534,N_11544,N_11673);
nor U14535 (N_14535,N_9439,N_11124);
or U14536 (N_14536,N_9138,N_9742);
nor U14537 (N_14537,N_10101,N_10072);
and U14538 (N_14538,N_11058,N_11738);
nor U14539 (N_14539,N_9045,N_10982);
nand U14540 (N_14540,N_9413,N_11555);
nand U14541 (N_14541,N_10950,N_10652);
and U14542 (N_14542,N_10018,N_9257);
and U14543 (N_14543,N_10128,N_9030);
xor U14544 (N_14544,N_11380,N_9054);
nor U14545 (N_14545,N_10107,N_11447);
nor U14546 (N_14546,N_10122,N_11235);
or U14547 (N_14547,N_9171,N_9911);
nand U14548 (N_14548,N_11548,N_10036);
or U14549 (N_14549,N_10324,N_11361);
nand U14550 (N_14550,N_9885,N_10710);
and U14551 (N_14551,N_11169,N_9019);
and U14552 (N_14552,N_11722,N_9441);
nor U14553 (N_14553,N_10941,N_9114);
nor U14554 (N_14554,N_9273,N_9658);
nand U14555 (N_14555,N_10279,N_10938);
nand U14556 (N_14556,N_11520,N_10208);
nand U14557 (N_14557,N_10516,N_9778);
and U14558 (N_14558,N_10024,N_9512);
or U14559 (N_14559,N_9217,N_9871);
or U14560 (N_14560,N_11640,N_10865);
nor U14561 (N_14561,N_9949,N_10029);
nand U14562 (N_14562,N_9812,N_9335);
nand U14563 (N_14563,N_9483,N_10289);
nor U14564 (N_14564,N_11839,N_9345);
nor U14565 (N_14565,N_10649,N_9822);
or U14566 (N_14566,N_9397,N_10529);
nand U14567 (N_14567,N_10542,N_10500);
nand U14568 (N_14568,N_11281,N_11277);
nand U14569 (N_14569,N_10100,N_9770);
and U14570 (N_14570,N_10432,N_9488);
nand U14571 (N_14571,N_10368,N_11244);
or U14572 (N_14572,N_10449,N_9194);
and U14573 (N_14573,N_10578,N_10721);
nor U14574 (N_14574,N_9092,N_11245);
and U14575 (N_14575,N_10340,N_9377);
and U14576 (N_14576,N_10774,N_10194);
or U14577 (N_14577,N_10742,N_9928);
nand U14578 (N_14578,N_10468,N_11311);
nand U14579 (N_14579,N_10011,N_10768);
nand U14580 (N_14580,N_11633,N_11732);
or U14581 (N_14581,N_10934,N_11009);
nand U14582 (N_14582,N_10486,N_11782);
nor U14583 (N_14583,N_10050,N_9242);
xnor U14584 (N_14584,N_10205,N_11696);
nand U14585 (N_14585,N_9413,N_10063);
nand U14586 (N_14586,N_9035,N_11392);
nor U14587 (N_14587,N_11809,N_9761);
xnor U14588 (N_14588,N_10947,N_10785);
or U14589 (N_14589,N_11251,N_11581);
nand U14590 (N_14590,N_9381,N_11251);
xor U14591 (N_14591,N_10536,N_9086);
or U14592 (N_14592,N_9765,N_11469);
nor U14593 (N_14593,N_10507,N_9641);
nor U14594 (N_14594,N_10616,N_11796);
nor U14595 (N_14595,N_10535,N_10122);
nand U14596 (N_14596,N_9978,N_11628);
or U14597 (N_14597,N_9509,N_9448);
nand U14598 (N_14598,N_10529,N_11420);
and U14599 (N_14599,N_9157,N_10285);
nor U14600 (N_14600,N_10548,N_10140);
nand U14601 (N_14601,N_10683,N_10808);
and U14602 (N_14602,N_10441,N_9168);
and U14603 (N_14603,N_11531,N_9263);
nor U14604 (N_14604,N_11613,N_9599);
nor U14605 (N_14605,N_10141,N_9080);
or U14606 (N_14606,N_10051,N_9350);
or U14607 (N_14607,N_10384,N_9176);
xnor U14608 (N_14608,N_10772,N_9995);
nand U14609 (N_14609,N_10122,N_11612);
and U14610 (N_14610,N_10298,N_11508);
nand U14611 (N_14611,N_9408,N_11637);
and U14612 (N_14612,N_10392,N_9917);
and U14613 (N_14613,N_10657,N_9334);
or U14614 (N_14614,N_11869,N_10511);
xor U14615 (N_14615,N_9145,N_9782);
or U14616 (N_14616,N_11986,N_10724);
nor U14617 (N_14617,N_11166,N_9374);
or U14618 (N_14618,N_9170,N_11874);
nand U14619 (N_14619,N_11257,N_9895);
or U14620 (N_14620,N_10296,N_9741);
and U14621 (N_14621,N_11016,N_11415);
and U14622 (N_14622,N_11155,N_9911);
and U14623 (N_14623,N_10192,N_11788);
nor U14624 (N_14624,N_11195,N_9072);
and U14625 (N_14625,N_11288,N_9467);
nand U14626 (N_14626,N_9800,N_11058);
nor U14627 (N_14627,N_11714,N_10817);
nand U14628 (N_14628,N_9145,N_9832);
and U14629 (N_14629,N_11971,N_9139);
nand U14630 (N_14630,N_11910,N_10096);
nor U14631 (N_14631,N_10242,N_9136);
xnor U14632 (N_14632,N_9267,N_10380);
and U14633 (N_14633,N_10105,N_11236);
and U14634 (N_14634,N_9512,N_9319);
and U14635 (N_14635,N_10681,N_9247);
nor U14636 (N_14636,N_11020,N_11032);
and U14637 (N_14637,N_11376,N_9604);
and U14638 (N_14638,N_9193,N_11192);
nor U14639 (N_14639,N_10101,N_10598);
and U14640 (N_14640,N_9254,N_10930);
and U14641 (N_14641,N_10784,N_10545);
xor U14642 (N_14642,N_10518,N_9576);
nor U14643 (N_14643,N_11800,N_10875);
and U14644 (N_14644,N_9208,N_10906);
and U14645 (N_14645,N_10007,N_11044);
or U14646 (N_14646,N_10503,N_11530);
and U14647 (N_14647,N_9560,N_10621);
or U14648 (N_14648,N_9188,N_11109);
nand U14649 (N_14649,N_11869,N_9296);
nand U14650 (N_14650,N_11552,N_11981);
or U14651 (N_14651,N_9663,N_9120);
and U14652 (N_14652,N_11240,N_9209);
nor U14653 (N_14653,N_11966,N_11366);
nor U14654 (N_14654,N_11822,N_9422);
and U14655 (N_14655,N_9058,N_10912);
or U14656 (N_14656,N_9989,N_10807);
nand U14657 (N_14657,N_10428,N_11187);
nor U14658 (N_14658,N_10978,N_11114);
xor U14659 (N_14659,N_9487,N_10219);
or U14660 (N_14660,N_9913,N_10825);
nand U14661 (N_14661,N_9338,N_9912);
nand U14662 (N_14662,N_9685,N_9426);
nand U14663 (N_14663,N_10648,N_10661);
nor U14664 (N_14664,N_11212,N_9989);
or U14665 (N_14665,N_9361,N_11293);
nor U14666 (N_14666,N_11734,N_9066);
xnor U14667 (N_14667,N_10259,N_9657);
nor U14668 (N_14668,N_9402,N_11593);
or U14669 (N_14669,N_10503,N_9196);
nand U14670 (N_14670,N_10250,N_10688);
and U14671 (N_14671,N_9955,N_10204);
nor U14672 (N_14672,N_9956,N_10313);
nor U14673 (N_14673,N_9664,N_11883);
or U14674 (N_14674,N_10496,N_9676);
nand U14675 (N_14675,N_11911,N_10422);
nand U14676 (N_14676,N_9982,N_11500);
nand U14677 (N_14677,N_10553,N_11752);
or U14678 (N_14678,N_9481,N_10941);
and U14679 (N_14679,N_10835,N_10438);
nor U14680 (N_14680,N_10643,N_10443);
xor U14681 (N_14681,N_9156,N_10186);
xnor U14682 (N_14682,N_9187,N_11278);
xor U14683 (N_14683,N_10424,N_9371);
or U14684 (N_14684,N_9769,N_9867);
nand U14685 (N_14685,N_11297,N_10121);
nor U14686 (N_14686,N_10390,N_9115);
or U14687 (N_14687,N_9038,N_11645);
xor U14688 (N_14688,N_10887,N_10131);
or U14689 (N_14689,N_10101,N_10876);
nor U14690 (N_14690,N_10686,N_9991);
xnor U14691 (N_14691,N_9662,N_10520);
and U14692 (N_14692,N_9600,N_9367);
nor U14693 (N_14693,N_10339,N_10367);
nor U14694 (N_14694,N_11257,N_11572);
and U14695 (N_14695,N_9839,N_11664);
nand U14696 (N_14696,N_11467,N_10919);
nand U14697 (N_14697,N_10690,N_9425);
nand U14698 (N_14698,N_10678,N_11624);
nand U14699 (N_14699,N_11338,N_10747);
nand U14700 (N_14700,N_9259,N_10920);
nor U14701 (N_14701,N_9939,N_10510);
nor U14702 (N_14702,N_9779,N_9045);
or U14703 (N_14703,N_11728,N_9806);
nor U14704 (N_14704,N_10755,N_10986);
and U14705 (N_14705,N_11851,N_10466);
nor U14706 (N_14706,N_11620,N_9161);
nand U14707 (N_14707,N_11885,N_9176);
nand U14708 (N_14708,N_11742,N_9823);
nor U14709 (N_14709,N_9879,N_9301);
and U14710 (N_14710,N_10058,N_11013);
nand U14711 (N_14711,N_11962,N_9616);
or U14712 (N_14712,N_9046,N_11447);
xor U14713 (N_14713,N_9797,N_9842);
or U14714 (N_14714,N_10907,N_11560);
xor U14715 (N_14715,N_9632,N_9599);
nand U14716 (N_14716,N_9470,N_11183);
or U14717 (N_14717,N_9461,N_9229);
nor U14718 (N_14718,N_9707,N_10129);
nand U14719 (N_14719,N_11182,N_9899);
or U14720 (N_14720,N_11148,N_9218);
nor U14721 (N_14721,N_9056,N_10125);
nand U14722 (N_14722,N_11673,N_9957);
nand U14723 (N_14723,N_9381,N_10388);
nor U14724 (N_14724,N_10246,N_11387);
and U14725 (N_14725,N_10156,N_9948);
nor U14726 (N_14726,N_11202,N_10217);
or U14727 (N_14727,N_10269,N_9033);
xor U14728 (N_14728,N_10578,N_9225);
nand U14729 (N_14729,N_10899,N_10458);
nor U14730 (N_14730,N_9323,N_10835);
or U14731 (N_14731,N_9304,N_10821);
xnor U14732 (N_14732,N_9721,N_11418);
xor U14733 (N_14733,N_9596,N_9137);
nor U14734 (N_14734,N_11251,N_9627);
and U14735 (N_14735,N_10757,N_10951);
nand U14736 (N_14736,N_10931,N_11539);
nand U14737 (N_14737,N_11095,N_11203);
and U14738 (N_14738,N_11617,N_10174);
nand U14739 (N_14739,N_11876,N_10985);
or U14740 (N_14740,N_9936,N_10543);
and U14741 (N_14741,N_11513,N_9656);
nor U14742 (N_14742,N_9663,N_10893);
and U14743 (N_14743,N_10138,N_9156);
or U14744 (N_14744,N_10921,N_9048);
nand U14745 (N_14745,N_9444,N_11371);
nor U14746 (N_14746,N_10205,N_11606);
nand U14747 (N_14747,N_11357,N_9498);
and U14748 (N_14748,N_10973,N_11111);
or U14749 (N_14749,N_10921,N_10918);
or U14750 (N_14750,N_9272,N_11488);
nand U14751 (N_14751,N_9391,N_10052);
and U14752 (N_14752,N_11792,N_10106);
nor U14753 (N_14753,N_10388,N_10479);
and U14754 (N_14754,N_10325,N_9187);
or U14755 (N_14755,N_11885,N_11804);
nand U14756 (N_14756,N_10918,N_11910);
xor U14757 (N_14757,N_10737,N_10646);
and U14758 (N_14758,N_11934,N_9451);
nand U14759 (N_14759,N_11040,N_10776);
nand U14760 (N_14760,N_9661,N_9906);
nand U14761 (N_14761,N_9769,N_10472);
and U14762 (N_14762,N_9936,N_11541);
nor U14763 (N_14763,N_10205,N_9938);
or U14764 (N_14764,N_11478,N_11059);
or U14765 (N_14765,N_11022,N_11902);
or U14766 (N_14766,N_11514,N_11945);
nand U14767 (N_14767,N_10744,N_10349);
nand U14768 (N_14768,N_10629,N_10501);
nand U14769 (N_14769,N_11896,N_10396);
xor U14770 (N_14770,N_9265,N_11692);
and U14771 (N_14771,N_9553,N_9044);
and U14772 (N_14772,N_11354,N_10363);
and U14773 (N_14773,N_9981,N_11834);
or U14774 (N_14774,N_10410,N_9305);
nand U14775 (N_14775,N_11458,N_10104);
or U14776 (N_14776,N_9090,N_11851);
xnor U14777 (N_14777,N_11747,N_9251);
nand U14778 (N_14778,N_9269,N_9216);
xor U14779 (N_14779,N_11148,N_11385);
nor U14780 (N_14780,N_11287,N_11327);
nor U14781 (N_14781,N_9028,N_11254);
xor U14782 (N_14782,N_10634,N_9094);
nor U14783 (N_14783,N_9412,N_9269);
nor U14784 (N_14784,N_9113,N_9039);
or U14785 (N_14785,N_11118,N_10152);
and U14786 (N_14786,N_11038,N_11952);
or U14787 (N_14787,N_10023,N_10557);
xnor U14788 (N_14788,N_9031,N_11471);
or U14789 (N_14789,N_9546,N_9063);
nor U14790 (N_14790,N_9475,N_11737);
nor U14791 (N_14791,N_11267,N_9801);
nor U14792 (N_14792,N_11159,N_11681);
or U14793 (N_14793,N_9502,N_10850);
xnor U14794 (N_14794,N_9823,N_10307);
nor U14795 (N_14795,N_10854,N_10652);
nor U14796 (N_14796,N_9418,N_11465);
nor U14797 (N_14797,N_10587,N_9441);
nand U14798 (N_14798,N_10630,N_9570);
and U14799 (N_14799,N_10792,N_9882);
xnor U14800 (N_14800,N_11451,N_11446);
and U14801 (N_14801,N_10557,N_11419);
and U14802 (N_14802,N_9967,N_10621);
nor U14803 (N_14803,N_11462,N_10431);
or U14804 (N_14804,N_10221,N_10276);
nand U14805 (N_14805,N_10562,N_10394);
nand U14806 (N_14806,N_10656,N_11779);
nor U14807 (N_14807,N_9644,N_10542);
nor U14808 (N_14808,N_9135,N_9024);
and U14809 (N_14809,N_11506,N_10045);
nand U14810 (N_14810,N_9026,N_9299);
or U14811 (N_14811,N_9114,N_10418);
and U14812 (N_14812,N_10474,N_10707);
and U14813 (N_14813,N_11311,N_10114);
or U14814 (N_14814,N_10326,N_9163);
and U14815 (N_14815,N_9743,N_11566);
or U14816 (N_14816,N_10254,N_10375);
or U14817 (N_14817,N_10969,N_10101);
or U14818 (N_14818,N_11988,N_10315);
and U14819 (N_14819,N_11308,N_9838);
or U14820 (N_14820,N_11753,N_10139);
nor U14821 (N_14821,N_11851,N_11498);
nand U14822 (N_14822,N_10414,N_10350);
nor U14823 (N_14823,N_11014,N_9556);
nand U14824 (N_14824,N_9008,N_11615);
nand U14825 (N_14825,N_11934,N_10868);
and U14826 (N_14826,N_10277,N_10159);
and U14827 (N_14827,N_11442,N_9136);
nand U14828 (N_14828,N_11945,N_10644);
nand U14829 (N_14829,N_11964,N_11162);
nor U14830 (N_14830,N_10038,N_10737);
and U14831 (N_14831,N_11567,N_11581);
xor U14832 (N_14832,N_10154,N_9913);
nor U14833 (N_14833,N_9050,N_10149);
nor U14834 (N_14834,N_9916,N_10605);
xnor U14835 (N_14835,N_11753,N_10736);
or U14836 (N_14836,N_9785,N_9919);
nor U14837 (N_14837,N_9698,N_9800);
nand U14838 (N_14838,N_10530,N_11355);
and U14839 (N_14839,N_11039,N_11459);
xor U14840 (N_14840,N_11203,N_10404);
xor U14841 (N_14841,N_10939,N_11640);
or U14842 (N_14842,N_9541,N_11608);
or U14843 (N_14843,N_9471,N_9173);
nor U14844 (N_14844,N_9135,N_10669);
nor U14845 (N_14845,N_9410,N_10442);
and U14846 (N_14846,N_9052,N_10910);
and U14847 (N_14847,N_11772,N_11658);
xnor U14848 (N_14848,N_9572,N_9957);
or U14849 (N_14849,N_11918,N_9315);
nor U14850 (N_14850,N_9300,N_9048);
nand U14851 (N_14851,N_11145,N_11369);
and U14852 (N_14852,N_10866,N_10998);
nor U14853 (N_14853,N_10330,N_10504);
and U14854 (N_14854,N_9370,N_10129);
nor U14855 (N_14855,N_10110,N_11761);
or U14856 (N_14856,N_10744,N_10618);
nor U14857 (N_14857,N_11152,N_11774);
nor U14858 (N_14858,N_9892,N_10911);
or U14859 (N_14859,N_9389,N_11238);
and U14860 (N_14860,N_9933,N_9514);
nand U14861 (N_14861,N_9225,N_9055);
nor U14862 (N_14862,N_10434,N_9448);
or U14863 (N_14863,N_9846,N_11088);
nor U14864 (N_14864,N_10211,N_9252);
nand U14865 (N_14865,N_11910,N_11724);
xor U14866 (N_14866,N_9815,N_10826);
nor U14867 (N_14867,N_11744,N_9741);
nand U14868 (N_14868,N_10853,N_11747);
xor U14869 (N_14869,N_11391,N_11565);
and U14870 (N_14870,N_11822,N_10052);
and U14871 (N_14871,N_11127,N_11431);
nor U14872 (N_14872,N_9160,N_9766);
or U14873 (N_14873,N_10692,N_9508);
and U14874 (N_14874,N_9801,N_9556);
nand U14875 (N_14875,N_11688,N_9452);
nor U14876 (N_14876,N_10329,N_9481);
or U14877 (N_14877,N_9680,N_11696);
and U14878 (N_14878,N_11421,N_11926);
nand U14879 (N_14879,N_10656,N_11987);
nand U14880 (N_14880,N_10252,N_9453);
and U14881 (N_14881,N_10402,N_10463);
and U14882 (N_14882,N_11858,N_9794);
nand U14883 (N_14883,N_9618,N_11154);
or U14884 (N_14884,N_10713,N_11837);
or U14885 (N_14885,N_10798,N_9129);
nor U14886 (N_14886,N_11185,N_11575);
or U14887 (N_14887,N_11276,N_11939);
and U14888 (N_14888,N_9809,N_11015);
nor U14889 (N_14889,N_9572,N_10372);
nand U14890 (N_14890,N_9479,N_10558);
and U14891 (N_14891,N_9604,N_10113);
xnor U14892 (N_14892,N_10562,N_9305);
nor U14893 (N_14893,N_9347,N_11496);
and U14894 (N_14894,N_10787,N_9850);
nor U14895 (N_14895,N_9651,N_9665);
nand U14896 (N_14896,N_9666,N_9194);
or U14897 (N_14897,N_9295,N_11485);
or U14898 (N_14898,N_9798,N_9938);
nand U14899 (N_14899,N_10326,N_11649);
xor U14900 (N_14900,N_11121,N_9002);
xor U14901 (N_14901,N_11510,N_9129);
and U14902 (N_14902,N_9374,N_11949);
and U14903 (N_14903,N_10777,N_9945);
xor U14904 (N_14904,N_9391,N_9833);
and U14905 (N_14905,N_11649,N_11785);
nand U14906 (N_14906,N_11050,N_9088);
nor U14907 (N_14907,N_9572,N_11832);
or U14908 (N_14908,N_11854,N_11359);
nor U14909 (N_14909,N_10623,N_11613);
xor U14910 (N_14910,N_9547,N_11980);
or U14911 (N_14911,N_10263,N_10269);
nor U14912 (N_14912,N_10603,N_10057);
nor U14913 (N_14913,N_11261,N_11204);
xnor U14914 (N_14914,N_10270,N_11238);
and U14915 (N_14915,N_9972,N_9768);
xor U14916 (N_14916,N_11112,N_10382);
nor U14917 (N_14917,N_10567,N_11361);
nor U14918 (N_14918,N_11279,N_10974);
and U14919 (N_14919,N_9071,N_10988);
nor U14920 (N_14920,N_11369,N_9059);
nor U14921 (N_14921,N_11882,N_10368);
xnor U14922 (N_14922,N_11348,N_9705);
nand U14923 (N_14923,N_9289,N_10717);
nand U14924 (N_14924,N_11475,N_10213);
nor U14925 (N_14925,N_9207,N_11565);
nand U14926 (N_14926,N_10377,N_9791);
nand U14927 (N_14927,N_10362,N_11764);
nor U14928 (N_14928,N_11063,N_10298);
nand U14929 (N_14929,N_11621,N_10818);
and U14930 (N_14930,N_11836,N_10549);
nor U14931 (N_14931,N_10413,N_10908);
nor U14932 (N_14932,N_9832,N_10557);
nand U14933 (N_14933,N_10032,N_9254);
or U14934 (N_14934,N_9277,N_10439);
nor U14935 (N_14935,N_10337,N_10654);
and U14936 (N_14936,N_11248,N_11910);
or U14937 (N_14937,N_9822,N_11860);
xnor U14938 (N_14938,N_9449,N_11494);
and U14939 (N_14939,N_10672,N_11389);
and U14940 (N_14940,N_9009,N_11264);
and U14941 (N_14941,N_11797,N_9620);
or U14942 (N_14942,N_9365,N_11210);
nor U14943 (N_14943,N_9896,N_11557);
nor U14944 (N_14944,N_9781,N_9564);
or U14945 (N_14945,N_10526,N_11161);
or U14946 (N_14946,N_10015,N_11943);
and U14947 (N_14947,N_9061,N_9833);
nand U14948 (N_14948,N_10882,N_11194);
nand U14949 (N_14949,N_9762,N_10411);
and U14950 (N_14950,N_9896,N_10985);
and U14951 (N_14951,N_10313,N_10166);
or U14952 (N_14952,N_11819,N_10951);
nor U14953 (N_14953,N_9001,N_9510);
xnor U14954 (N_14954,N_9974,N_9264);
nand U14955 (N_14955,N_9079,N_9272);
nand U14956 (N_14956,N_10282,N_9541);
nand U14957 (N_14957,N_10688,N_10610);
nand U14958 (N_14958,N_11075,N_9740);
or U14959 (N_14959,N_11996,N_11850);
or U14960 (N_14960,N_11552,N_11577);
nand U14961 (N_14961,N_9048,N_11266);
nor U14962 (N_14962,N_10706,N_11777);
xnor U14963 (N_14963,N_11629,N_11600);
nor U14964 (N_14964,N_11928,N_10440);
nor U14965 (N_14965,N_11016,N_9512);
nor U14966 (N_14966,N_10583,N_9179);
nand U14967 (N_14967,N_11183,N_11759);
nand U14968 (N_14968,N_11320,N_9940);
and U14969 (N_14969,N_10651,N_11925);
or U14970 (N_14970,N_10643,N_11537);
xnor U14971 (N_14971,N_10730,N_11371);
nor U14972 (N_14972,N_10750,N_11891);
nor U14973 (N_14973,N_10102,N_10480);
or U14974 (N_14974,N_10149,N_10729);
nand U14975 (N_14975,N_9743,N_11625);
nor U14976 (N_14976,N_10489,N_9145);
nor U14977 (N_14977,N_9104,N_10864);
nand U14978 (N_14978,N_9304,N_11735);
nor U14979 (N_14979,N_9861,N_10483);
nand U14980 (N_14980,N_10927,N_10319);
nor U14981 (N_14981,N_11878,N_11817);
nand U14982 (N_14982,N_11811,N_10643);
or U14983 (N_14983,N_11126,N_9755);
nor U14984 (N_14984,N_10488,N_11645);
nand U14985 (N_14985,N_9929,N_9275);
nand U14986 (N_14986,N_11032,N_9934);
nand U14987 (N_14987,N_10094,N_11701);
nor U14988 (N_14988,N_9273,N_10711);
nand U14989 (N_14989,N_9300,N_11385);
nor U14990 (N_14990,N_9146,N_9337);
or U14991 (N_14991,N_11663,N_9593);
nor U14992 (N_14992,N_10556,N_9712);
or U14993 (N_14993,N_9106,N_10714);
nor U14994 (N_14994,N_10012,N_10735);
and U14995 (N_14995,N_9748,N_9938);
nand U14996 (N_14996,N_10135,N_9623);
and U14997 (N_14997,N_10989,N_9192);
or U14998 (N_14998,N_9545,N_9697);
or U14999 (N_14999,N_9432,N_10242);
nor UO_0 (O_0,N_13959,N_12600);
nand UO_1 (O_1,N_13978,N_13113);
or UO_2 (O_2,N_13599,N_14161);
xnor UO_3 (O_3,N_14268,N_12213);
nand UO_4 (O_4,N_13748,N_13092);
nand UO_5 (O_5,N_12215,N_14746);
and UO_6 (O_6,N_14734,N_13646);
nor UO_7 (O_7,N_12671,N_13015);
xnor UO_8 (O_8,N_12329,N_14551);
or UO_9 (O_9,N_13665,N_14825);
and UO_10 (O_10,N_13543,N_14406);
or UO_11 (O_11,N_12682,N_13107);
nor UO_12 (O_12,N_14656,N_13289);
nand UO_13 (O_13,N_12366,N_12577);
nand UO_14 (O_14,N_12390,N_12833);
nor UO_15 (O_15,N_14378,N_14590);
nor UO_16 (O_16,N_14120,N_14547);
or UO_17 (O_17,N_13782,N_13935);
xnor UO_18 (O_18,N_14178,N_12327);
or UO_19 (O_19,N_13409,N_14413);
and UO_20 (O_20,N_12207,N_13727);
or UO_21 (O_21,N_13290,N_14070);
nor UO_22 (O_22,N_13279,N_12744);
or UO_23 (O_23,N_14117,N_13282);
nand UO_24 (O_24,N_13122,N_14335);
and UO_25 (O_25,N_12546,N_13733);
nand UO_26 (O_26,N_13298,N_12801);
or UO_27 (O_27,N_13336,N_12898);
and UO_28 (O_28,N_14211,N_14663);
nand UO_29 (O_29,N_14486,N_14035);
nand UO_30 (O_30,N_12344,N_13096);
or UO_31 (O_31,N_12512,N_12268);
and UO_32 (O_32,N_13189,N_12129);
and UO_33 (O_33,N_14855,N_13213);
or UO_34 (O_34,N_13652,N_14971);
nand UO_35 (O_35,N_13264,N_12084);
and UO_36 (O_36,N_12638,N_14505);
or UO_37 (O_37,N_12325,N_14146);
and UO_38 (O_38,N_12654,N_13559);
or UO_39 (O_39,N_14031,N_14341);
and UO_40 (O_40,N_13094,N_14124);
nand UO_41 (O_41,N_14735,N_12515);
nor UO_42 (O_42,N_14201,N_13453);
nand UO_43 (O_43,N_12653,N_13544);
nand UO_44 (O_44,N_12594,N_13839);
or UO_45 (O_45,N_13754,N_13204);
nand UO_46 (O_46,N_13831,N_12246);
nor UO_47 (O_47,N_13603,N_13238);
or UO_48 (O_48,N_13498,N_14476);
or UO_49 (O_49,N_13155,N_14611);
xor UO_50 (O_50,N_13191,N_13140);
and UO_51 (O_51,N_12857,N_12460);
nand UO_52 (O_52,N_12032,N_14078);
xnor UO_53 (O_53,N_12995,N_14732);
nor UO_54 (O_54,N_14087,N_13322);
and UO_55 (O_55,N_14275,N_12306);
xnor UO_56 (O_56,N_14381,N_13358);
and UO_57 (O_57,N_14299,N_14941);
xnor UO_58 (O_58,N_14755,N_14664);
nor UO_59 (O_59,N_13896,N_14456);
nand UO_60 (O_60,N_14500,N_12700);
or UO_61 (O_61,N_14581,N_12558);
and UO_62 (O_62,N_12205,N_13593);
and UO_63 (O_63,N_14319,N_12054);
or UO_64 (O_64,N_14577,N_14262);
and UO_65 (O_65,N_12364,N_14959);
and UO_66 (O_66,N_12313,N_12738);
nand UO_67 (O_67,N_14502,N_12373);
or UO_68 (O_68,N_12858,N_14974);
or UO_69 (O_69,N_14968,N_12230);
xnor UO_70 (O_70,N_14585,N_12878);
xnor UO_71 (O_71,N_13390,N_12873);
and UO_72 (O_72,N_13542,N_14294);
or UO_73 (O_73,N_14243,N_12647);
nand UO_74 (O_74,N_13654,N_12191);
nand UO_75 (O_75,N_13458,N_14565);
nor UO_76 (O_76,N_12667,N_12828);
and UO_77 (O_77,N_13971,N_13635);
nor UO_78 (O_78,N_12384,N_14858);
nor UO_79 (O_79,N_13497,N_14228);
or UO_80 (O_80,N_12848,N_13234);
nand UO_81 (O_81,N_13442,N_13979);
nand UO_82 (O_82,N_14127,N_12776);
nand UO_83 (O_83,N_13469,N_13031);
nand UO_84 (O_84,N_12935,N_14730);
nor UO_85 (O_85,N_12061,N_14556);
nand UO_86 (O_86,N_12825,N_13487);
and UO_87 (O_87,N_13074,N_14007);
nor UO_88 (O_88,N_13731,N_12122);
nor UO_89 (O_89,N_13346,N_14793);
nand UO_90 (O_90,N_12971,N_13965);
nand UO_91 (O_91,N_14754,N_13243);
nor UO_92 (O_92,N_14434,N_12637);
or UO_93 (O_93,N_12049,N_14284);
or UO_94 (O_94,N_12754,N_12714);
and UO_95 (O_95,N_14153,N_14155);
or UO_96 (O_96,N_13779,N_13580);
and UO_97 (O_97,N_12245,N_12928);
nand UO_98 (O_98,N_14163,N_12830);
nor UO_99 (O_99,N_14699,N_13997);
or UO_100 (O_100,N_12798,N_12285);
or UO_101 (O_101,N_14894,N_12936);
and UO_102 (O_102,N_12768,N_12255);
or UO_103 (O_103,N_14308,N_14792);
and UO_104 (O_104,N_13633,N_13172);
nor UO_105 (O_105,N_13156,N_14644);
nor UO_106 (O_106,N_13833,N_13974);
and UO_107 (O_107,N_13832,N_14379);
nand UO_108 (O_108,N_12144,N_13202);
or UO_109 (O_109,N_13014,N_12818);
nand UO_110 (O_110,N_14318,N_13389);
nand UO_111 (O_111,N_12314,N_14890);
nand UO_112 (O_112,N_13317,N_13843);
or UO_113 (O_113,N_13925,N_12094);
and UO_114 (O_114,N_12254,N_12326);
nor UO_115 (O_115,N_12757,N_13527);
and UO_116 (O_116,N_14900,N_12787);
and UO_117 (O_117,N_13129,N_14451);
nor UO_118 (O_118,N_14952,N_13802);
nand UO_119 (O_119,N_13132,N_14784);
and UO_120 (O_120,N_13115,N_13364);
nand UO_121 (O_121,N_12549,N_12186);
or UO_122 (O_122,N_14179,N_12605);
nand UO_123 (O_123,N_13316,N_13570);
nand UO_124 (O_124,N_13299,N_14753);
nor UO_125 (O_125,N_12089,N_14295);
nand UO_126 (O_126,N_13471,N_12752);
and UO_127 (O_127,N_14956,N_13809);
or UO_128 (O_128,N_14189,N_13973);
nor UO_129 (O_129,N_14237,N_13569);
nor UO_130 (O_130,N_14978,N_13319);
nand UO_131 (O_131,N_13626,N_13144);
nand UO_132 (O_132,N_14516,N_13340);
nand UO_133 (O_133,N_14705,N_14857);
xor UO_134 (O_134,N_13632,N_14367);
nor UO_135 (O_135,N_12553,N_12824);
and UO_136 (O_136,N_13003,N_13105);
nand UO_137 (O_137,N_12079,N_12575);
or UO_138 (O_138,N_13110,N_14336);
nor UO_139 (O_139,N_13566,N_14122);
and UO_140 (O_140,N_14427,N_12118);
nor UO_141 (O_141,N_14386,N_13605);
xor UO_142 (O_142,N_13434,N_14036);
nand UO_143 (O_143,N_13022,N_12680);
or UO_144 (O_144,N_14643,N_14404);
nand UO_145 (O_145,N_14786,N_12911);
and UO_146 (O_146,N_13584,N_12424);
and UO_147 (O_147,N_12713,N_13499);
nand UO_148 (O_148,N_13417,N_12781);
nor UO_149 (O_149,N_12222,N_14926);
or UO_150 (O_150,N_13511,N_13670);
xnor UO_151 (O_151,N_13478,N_14655);
and UO_152 (O_152,N_14853,N_14954);
nand UO_153 (O_153,N_14029,N_14396);
xor UO_154 (O_154,N_14492,N_13255);
or UO_155 (O_155,N_13787,N_12992);
and UO_156 (O_156,N_12426,N_14553);
or UO_157 (O_157,N_13987,N_12674);
nor UO_158 (O_158,N_12634,N_13119);
and UO_159 (O_159,N_14447,N_14095);
nor UO_160 (O_160,N_12349,N_13966);
and UO_161 (O_161,N_13445,N_13529);
nand UO_162 (O_162,N_13021,N_12448);
nor UO_163 (O_163,N_14241,N_14706);
nor UO_164 (O_164,N_13009,N_14554);
nor UO_165 (O_165,N_13806,N_13112);
nor UO_166 (O_166,N_12906,N_12339);
nor UO_167 (O_167,N_12291,N_12778);
and UO_168 (O_168,N_12739,N_13516);
and UO_169 (O_169,N_12888,N_13993);
nand UO_170 (O_170,N_12405,N_12095);
nor UO_171 (O_171,N_12136,N_14250);
nor UO_172 (O_172,N_14364,N_13372);
nand UO_173 (O_173,N_13175,N_13373);
nand UO_174 (O_174,N_12815,N_13900);
and UO_175 (O_175,N_12444,N_13791);
xor UO_176 (O_176,N_14116,N_14843);
nor UO_177 (O_177,N_14651,N_13099);
and UO_178 (O_178,N_14313,N_13315);
nand UO_179 (O_179,N_13909,N_12636);
or UO_180 (O_180,N_13361,N_12529);
nor UO_181 (O_181,N_12492,N_14046);
and UO_182 (O_182,N_12821,N_14795);
nor UO_183 (O_183,N_13607,N_13276);
nor UO_184 (O_184,N_14158,N_12035);
nand UO_185 (O_185,N_12792,N_13065);
and UO_186 (O_186,N_13089,N_12038);
or UO_187 (O_187,N_13734,N_13206);
and UO_188 (O_188,N_13784,N_12080);
and UO_189 (O_189,N_12606,N_14722);
and UO_190 (O_190,N_13045,N_14809);
nand UO_191 (O_191,N_14756,N_13352);
and UO_192 (O_192,N_13715,N_13781);
nand UO_193 (O_193,N_14563,N_13455);
and UO_194 (O_194,N_12323,N_14258);
nand UO_195 (O_195,N_12350,N_13232);
nor UO_196 (O_196,N_12056,N_13100);
nor UO_197 (O_197,N_12475,N_13981);
and UO_198 (O_198,N_12181,N_14869);
or UO_199 (O_199,N_13735,N_12124);
or UO_200 (O_200,N_14854,N_14052);
or UO_201 (O_201,N_14414,N_14454);
or UO_202 (O_202,N_13047,N_13248);
or UO_203 (O_203,N_12474,N_12839);
nor UO_204 (O_204,N_14707,N_14626);
nand UO_205 (O_205,N_14353,N_13746);
nand UO_206 (O_206,N_14600,N_13157);
or UO_207 (O_207,N_12946,N_14226);
nand UO_208 (O_208,N_12498,N_13994);
nor UO_209 (O_209,N_14860,N_14444);
or UO_210 (O_210,N_14215,N_14397);
nor UO_211 (O_211,N_13610,N_14824);
or UO_212 (O_212,N_12272,N_12321);
and UO_213 (O_213,N_13771,N_12704);
or UO_214 (O_214,N_13126,N_13533);
nand UO_215 (O_215,N_14647,N_13522);
or UO_216 (O_216,N_13291,N_13583);
or UO_217 (O_217,N_14708,N_14879);
or UO_218 (O_218,N_13812,N_13293);
or UO_219 (O_219,N_14519,N_13464);
nand UO_220 (O_220,N_12661,N_13770);
and UO_221 (O_221,N_12319,N_14607);
and UO_222 (O_222,N_13148,N_14162);
or UO_223 (O_223,N_13999,N_13850);
nand UO_224 (O_224,N_13338,N_14909);
or UO_225 (O_225,N_12114,N_13167);
nor UO_226 (O_226,N_12286,N_13363);
nor UO_227 (O_227,N_14069,N_12520);
or UO_228 (O_228,N_13852,N_14485);
xnor UO_229 (O_229,N_12915,N_12484);
xnor UO_230 (O_230,N_13829,N_13972);
or UO_231 (O_231,N_14443,N_14330);
or UO_232 (O_232,N_14641,N_13795);
and UO_233 (O_233,N_14936,N_12889);
and UO_234 (O_234,N_13117,N_12335);
and UO_235 (O_235,N_13944,N_14420);
or UO_236 (O_236,N_14468,N_13165);
or UO_237 (O_237,N_12678,N_14667);
or UO_238 (O_238,N_13086,N_12297);
or UO_239 (O_239,N_14895,N_13035);
or UO_240 (O_240,N_14230,N_14967);
or UO_241 (O_241,N_14180,N_13524);
nor UO_242 (O_242,N_13630,N_13922);
nand UO_243 (O_243,N_14957,N_14614);
nor UO_244 (O_244,N_12531,N_14040);
nor UO_245 (O_245,N_13413,N_12648);
nor UO_246 (O_246,N_13309,N_13354);
and UO_247 (O_247,N_12380,N_13058);
or UO_248 (O_248,N_13300,N_13668);
nor UO_249 (O_249,N_14467,N_12176);
or UO_250 (O_250,N_12208,N_14888);
nand UO_251 (O_251,N_12470,N_12456);
nor UO_252 (O_252,N_12891,N_12694);
or UO_253 (O_253,N_13307,N_14982);
and UO_254 (O_254,N_14359,N_12237);
nor UO_255 (O_255,N_14132,N_14453);
nor UO_256 (O_256,N_12951,N_12371);
nand UO_257 (O_257,N_13881,N_14334);
or UO_258 (O_258,N_14244,N_14441);
nor UO_259 (O_259,N_14701,N_14488);
and UO_260 (O_260,N_14238,N_14912);
and UO_261 (O_261,N_13173,N_14597);
nand UO_262 (O_262,N_14576,N_12773);
nand UO_263 (O_263,N_12289,N_14043);
and UO_264 (O_264,N_12625,N_12287);
or UO_265 (O_265,N_13328,N_12609);
or UO_266 (O_266,N_13486,N_13465);
and UO_267 (O_267,N_14586,N_12423);
nand UO_268 (O_268,N_12864,N_13220);
nor UO_269 (O_269,N_12188,N_13637);
nand UO_270 (O_270,N_14817,N_12265);
xnor UO_271 (O_271,N_13722,N_14415);
nand UO_272 (O_272,N_13656,N_14355);
xor UO_273 (O_273,N_14921,N_14839);
nand UO_274 (O_274,N_14812,N_12696);
nor UO_275 (O_275,N_13466,N_13163);
or UO_276 (O_276,N_14963,N_12722);
nand UO_277 (O_277,N_12775,N_12155);
and UO_278 (O_278,N_12536,N_14797);
or UO_279 (O_279,N_14431,N_12949);
nand UO_280 (O_280,N_13828,N_12855);
nand UO_281 (O_281,N_14645,N_14955);
and UO_282 (O_282,N_14739,N_14806);
nor UO_283 (O_283,N_12903,N_14901);
and UO_284 (O_284,N_12395,N_13483);
and UO_285 (O_285,N_13258,N_14992);
and UO_286 (O_286,N_14933,N_12379);
or UO_287 (O_287,N_12964,N_14990);
nand UO_288 (O_288,N_14693,N_12378);
and UO_289 (O_289,N_12708,N_14712);
or UO_290 (O_290,N_12042,N_13918);
and UO_291 (O_291,N_13397,N_13990);
nand UO_292 (O_292,N_12764,N_12175);
nand UO_293 (O_293,N_14961,N_14629);
nor UO_294 (O_294,N_13899,N_12202);
nor UO_295 (O_295,N_14008,N_14851);
nand UO_296 (O_296,N_12440,N_12487);
and UO_297 (O_297,N_12619,N_13071);
and UO_298 (O_298,N_12877,N_12590);
nor UO_299 (O_299,N_13391,N_13263);
and UO_300 (O_300,N_13756,N_13636);
and UO_301 (O_301,N_12970,N_14481);
nand UO_302 (O_302,N_14970,N_13326);
nand UO_303 (O_303,N_12733,N_12585);
and UO_304 (O_304,N_13568,N_14183);
and UO_305 (O_305,N_14836,N_13788);
and UO_306 (O_306,N_13621,N_14966);
nor UO_307 (O_307,N_13208,N_13484);
nor UO_308 (O_308,N_12257,N_12206);
xnor UO_309 (O_309,N_13379,N_12169);
and UO_310 (O_310,N_14167,N_14062);
nand UO_311 (O_311,N_13893,N_12802);
and UO_312 (O_312,N_12088,N_12510);
and UO_313 (O_313,N_14572,N_13749);
or UO_314 (O_314,N_13716,N_14616);
nand UO_315 (O_315,N_12357,N_13018);
nand UO_316 (O_316,N_12058,N_12576);
nand UO_317 (O_317,N_12358,N_14526);
nand UO_318 (O_318,N_12179,N_14994);
nand UO_319 (O_319,N_12142,N_13026);
nor UO_320 (O_320,N_14993,N_12140);
nand UO_321 (O_321,N_13101,N_13500);
or UO_322 (O_322,N_14061,N_12547);
nand UO_323 (O_323,N_14939,N_13414);
or UO_324 (O_324,N_13286,N_14717);
and UO_325 (O_325,N_14818,N_13153);
and UO_326 (O_326,N_12774,N_12106);
and UO_327 (O_327,N_14653,N_14896);
or UO_328 (O_328,N_12641,N_12737);
and UO_329 (O_329,N_13676,N_12865);
nand UO_330 (O_330,N_12132,N_13764);
or UO_331 (O_331,N_13171,N_12770);
and UO_332 (O_332,N_12897,N_14249);
or UO_333 (O_333,N_14401,N_13368);
or UO_334 (O_334,N_12893,N_12248);
nand UO_335 (O_335,N_13154,N_12218);
xor UO_336 (O_336,N_14491,N_12659);
nor UO_337 (O_337,N_14361,N_13851);
and UO_338 (O_338,N_14752,N_14587);
nand UO_339 (O_339,N_14579,N_13640);
or UO_340 (O_340,N_14130,N_12279);
nor UO_341 (O_341,N_14835,N_13842);
nor UO_342 (O_342,N_13392,N_13714);
or UO_343 (O_343,N_12309,N_12077);
nand UO_344 (O_344,N_12642,N_13267);
nor UO_345 (O_345,N_14018,N_12073);
and UO_346 (O_346,N_12952,N_12806);
nor UO_347 (O_347,N_14648,N_13878);
nand UO_348 (O_348,N_14410,N_13555);
nand UO_349 (O_349,N_13526,N_14542);
xnor UO_350 (O_350,N_13460,N_14908);
nor UO_351 (O_351,N_13785,N_13349);
nor UO_352 (O_352,N_12779,N_12087);
and UO_353 (O_353,N_14710,N_12672);
xnor UO_354 (O_354,N_12416,N_12355);
nand UO_355 (O_355,N_14068,N_14079);
or UO_356 (O_356,N_14141,N_12288);
and UO_357 (O_357,N_14170,N_14004);
nand UO_358 (O_358,N_14125,N_14202);
xor UO_359 (O_359,N_12699,N_13590);
and UO_360 (O_360,N_14603,N_12715);
nand UO_361 (O_361,N_13989,N_13147);
and UO_362 (O_362,N_14339,N_14814);
nand UO_363 (O_363,N_13701,N_12530);
nand UO_364 (O_364,N_14066,N_12559);
and UO_365 (O_365,N_14640,N_12324);
or UO_366 (O_366,N_12710,N_13507);
xor UO_367 (O_367,N_14919,N_14474);
and UO_368 (O_368,N_13273,N_12428);
nand UO_369 (O_369,N_14515,N_14609);
nand UO_370 (O_370,N_14652,N_12102);
xor UO_371 (O_371,N_12040,N_13216);
nor UO_372 (O_372,N_12973,N_14915);
nand UO_373 (O_373,N_12281,N_13532);
nor UO_374 (O_374,N_13970,N_12103);
or UO_375 (O_375,N_14140,N_14425);
and UO_376 (O_376,N_14271,N_12356);
nor UO_377 (O_377,N_13313,N_12716);
and UO_378 (O_378,N_13446,N_12535);
or UO_379 (O_379,N_12514,N_13182);
nor UO_380 (O_380,N_13027,N_13535);
nand UO_381 (O_381,N_12243,N_12771);
and UO_382 (O_382,N_13149,N_13864);
and UO_383 (O_383,N_13166,N_14395);
and UO_384 (O_384,N_13565,N_14343);
or UO_385 (O_385,N_13744,N_12948);
xor UO_386 (O_386,N_13639,N_13671);
nor UO_387 (O_387,N_12210,N_12723);
and UO_388 (O_388,N_14157,N_12068);
and UO_389 (O_389,N_12227,N_12432);
or UO_390 (O_390,N_14219,N_12919);
nand UO_391 (O_391,N_13139,N_13061);
and UO_392 (O_392,N_14612,N_14276);
and UO_393 (O_393,N_14235,N_14801);
nand UO_394 (O_394,N_14214,N_14139);
and UO_395 (O_395,N_12029,N_13116);
nand UO_396 (O_396,N_14882,N_13075);
and UO_397 (O_397,N_14385,N_13327);
nor UO_398 (O_398,N_13675,N_13692);
and UO_399 (O_399,N_13333,N_13585);
nand UO_400 (O_400,N_12011,N_14002);
and UO_401 (O_401,N_14665,N_13721);
or UO_402 (O_402,N_14914,N_12616);
and UO_403 (O_403,N_13564,N_14274);
nand UO_404 (O_404,N_12601,N_13287);
and UO_405 (O_405,N_12209,N_14151);
nor UO_406 (O_406,N_14077,N_14104);
or UO_407 (O_407,N_13314,N_12985);
or UO_408 (O_408,N_12668,N_12250);
and UO_409 (O_409,N_13310,N_12702);
nor UO_410 (O_410,N_14884,N_12564);
nand UO_411 (O_411,N_12701,N_13509);
or UO_412 (O_412,N_14159,N_13203);
nor UO_413 (O_413,N_12216,N_14511);
nand UO_414 (O_414,N_14679,N_12322);
or UO_415 (O_415,N_13385,N_12490);
or UO_416 (O_416,N_14398,N_13597);
and UO_417 (O_417,N_13143,N_13353);
and UO_418 (O_418,N_12522,N_12196);
nand UO_419 (O_419,N_12747,N_12067);
nor UO_420 (O_420,N_14771,N_14246);
nor UO_421 (O_421,N_12278,N_14538);
or UO_422 (O_422,N_12308,N_12938);
and UO_423 (O_423,N_14833,N_13684);
or UO_424 (O_424,N_12471,N_14777);
and UO_425 (O_425,N_13595,N_12883);
or UO_426 (O_426,N_14234,N_13384);
xor UO_427 (O_427,N_14723,N_14370);
or UO_428 (O_428,N_14015,N_12057);
nand UO_429 (O_429,N_12683,N_12370);
nand UO_430 (O_430,N_14631,N_13647);
nand UO_431 (O_431,N_12957,N_13013);
and UO_432 (O_432,N_13717,N_12840);
nor UO_433 (O_433,N_13888,N_12099);
xnor UO_434 (O_434,N_13412,N_13728);
nand UO_435 (O_435,N_14439,N_13142);
and UO_436 (O_436,N_13755,N_14412);
nand UO_437 (O_437,N_13423,N_12532);
nand UO_438 (O_438,N_13660,N_13098);
nor UO_439 (O_439,N_14862,N_14583);
or UO_440 (O_440,N_13266,N_13247);
nor UO_441 (O_441,N_14568,N_14164);
xnor UO_442 (O_442,N_12832,N_13774);
nand UO_443 (O_443,N_13662,N_13907);
or UO_444 (O_444,N_13194,N_14711);
or UO_445 (O_445,N_13275,N_14156);
or UO_446 (O_446,N_12860,N_12697);
or UO_447 (O_447,N_13673,N_13421);
and UO_448 (O_448,N_14889,N_12837);
and UO_449 (O_449,N_12586,N_14056);
xor UO_450 (O_450,N_13007,N_12203);
or UO_451 (O_451,N_14662,N_13252);
and UO_452 (O_452,N_13049,N_12381);
and UO_453 (O_453,N_12736,N_12582);
nor UO_454 (O_454,N_13927,N_12506);
nor UO_455 (O_455,N_14075,N_12958);
nand UO_456 (O_456,N_12902,N_14528);
nor UO_457 (O_457,N_13934,N_13548);
nor UO_458 (O_458,N_14826,N_12273);
and UO_459 (O_459,N_13554,N_13847);
and UO_460 (O_460,N_12611,N_12622);
and UO_461 (O_461,N_13841,N_12811);
or UO_462 (O_462,N_14521,N_14977);
xor UO_463 (O_463,N_13708,N_13561);
nand UO_464 (O_464,N_14023,N_14152);
nor UO_465 (O_465,N_12657,N_14424);
nor UO_466 (O_466,N_14113,N_12411);
xor UO_467 (O_467,N_13254,N_12527);
nand UO_468 (O_468,N_12336,N_13719);
or UO_469 (O_469,N_13520,N_14298);
nand UO_470 (O_470,N_12856,N_14205);
nor UO_471 (O_471,N_13056,N_14009);
xor UO_472 (O_472,N_12910,N_14346);
nor UO_473 (O_473,N_12725,N_12508);
or UO_474 (O_474,N_14314,N_14751);
or UO_475 (O_475,N_14269,N_12167);
nand UO_476 (O_476,N_13050,N_13270);
nand UO_477 (O_477,N_13622,N_12195);
or UO_478 (O_478,N_12660,N_13849);
or UO_479 (O_479,N_13669,N_14976);
and UO_480 (O_480,N_12748,N_14144);
nand UO_481 (O_481,N_14091,N_12503);
or UO_482 (O_482,N_13810,N_14975);
nand UO_483 (O_483,N_12987,N_14744);
nor UO_484 (O_484,N_12465,N_14863);
nand UO_485 (O_485,N_13926,N_14014);
nor UO_486 (O_486,N_14910,N_13631);
or UO_487 (O_487,N_14017,N_14695);
nor UO_488 (O_488,N_13135,N_13482);
nand UO_489 (O_489,N_12413,N_14807);
nand UO_490 (O_490,N_13800,N_13371);
nor UO_491 (O_491,N_13020,N_13547);
or UO_492 (O_492,N_12125,N_14991);
or UO_493 (O_493,N_13415,N_12190);
nand UO_494 (O_494,N_13920,N_13619);
xnor UO_495 (O_495,N_14462,N_13803);
or UO_496 (O_496,N_13052,N_14608);
and UO_497 (O_497,N_12879,N_13808);
nand UO_498 (O_498,N_13943,N_12495);
nand UO_499 (O_499,N_12310,N_14736);
or UO_500 (O_500,N_12563,N_14630);
and UO_501 (O_501,N_12219,N_12211);
and UO_502 (O_502,N_13347,N_14749);
and UO_503 (O_503,N_14293,N_12302);
and UO_504 (O_504,N_12720,N_14168);
nor UO_505 (O_505,N_13877,N_13948);
nor UO_506 (O_506,N_13001,N_13470);
nor UO_507 (O_507,N_13283,N_14536);
xor UO_508 (O_508,N_13396,N_12859);
nor UO_509 (O_509,N_14514,N_12134);
xor UO_510 (O_510,N_13898,N_14845);
or UO_511 (O_511,N_12317,N_13477);
or UO_512 (O_512,N_13295,N_12153);
or UO_513 (O_513,N_14721,N_12063);
nand UO_514 (O_514,N_12162,N_14844);
or UO_515 (O_515,N_14302,N_12756);
or UO_516 (O_516,N_14868,N_13259);
nor UO_517 (O_517,N_14489,N_14392);
nor UO_518 (O_518,N_14770,N_14621);
nand UO_519 (O_519,N_14634,N_14622);
nor UO_520 (O_520,N_12446,N_14633);
or UO_521 (O_521,N_13223,N_13146);
and UO_522 (O_522,N_12165,N_12296);
nor UO_523 (O_523,N_13917,N_14032);
and UO_524 (O_524,N_12746,N_14709);
or UO_525 (O_525,N_12969,N_12480);
or UO_526 (O_526,N_14333,N_13740);
or UO_527 (O_527,N_14738,N_12711);
and UO_528 (O_528,N_13694,N_12555);
and UO_529 (O_529,N_12123,N_13059);
nand UO_530 (O_530,N_12131,N_12603);
or UO_531 (O_531,N_14272,N_14632);
or UO_532 (O_532,N_12795,N_12817);
nor UO_533 (O_533,N_12868,N_13758);
nor UO_534 (O_534,N_13955,N_12024);
and UO_535 (O_535,N_13932,N_14848);
or UO_536 (O_536,N_14494,N_14400);
nand UO_537 (O_537,N_14074,N_14165);
and UO_538 (O_538,N_13271,N_13625);
xor UO_539 (O_539,N_14450,N_14535);
and UO_540 (O_540,N_12097,N_12295);
nor UO_541 (O_541,N_13538,N_13905);
and UO_542 (O_542,N_13854,N_12305);
or UO_543 (O_543,N_13941,N_14076);
or UO_544 (O_544,N_14192,N_13064);
nand UO_545 (O_545,N_13010,N_12628);
nor UO_546 (O_546,N_12831,N_14864);
nor UO_547 (O_547,N_13219,N_13377);
nand UO_548 (O_548,N_13950,N_13545);
and UO_549 (O_549,N_12796,N_14886);
xnor UO_550 (O_550,N_12043,N_12164);
and UO_551 (O_551,N_14000,N_12613);
or UO_552 (O_552,N_14593,N_13591);
and UO_553 (O_553,N_12021,N_14509);
and UO_554 (O_554,N_12908,N_12627);
nor UO_555 (O_555,N_14147,N_14995);
or UO_556 (O_556,N_12312,N_14935);
nand UO_557 (O_557,N_14768,N_12588);
nand UO_558 (O_558,N_14432,N_13737);
and UO_559 (O_559,N_13751,N_12518);
or UO_560 (O_560,N_12421,N_13296);
nor UO_561 (O_561,N_12462,N_14042);
nor UO_562 (O_562,N_13030,N_13792);
nor UO_563 (O_563,N_14027,N_14761);
nand UO_564 (O_564,N_12566,N_13091);
nor UO_565 (O_565,N_12942,N_12731);
or UO_566 (O_566,N_13304,N_12743);
nand UO_567 (O_567,N_13231,N_14904);
nor UO_568 (O_568,N_14578,N_13724);
or UO_569 (O_569,N_13120,N_13503);
nand UO_570 (O_570,N_13747,N_14217);
nand UO_571 (O_571,N_12793,N_13285);
xor UO_572 (O_572,N_14323,N_12742);
nor UO_573 (O_573,N_13663,N_13138);
nand UO_574 (O_574,N_13016,N_12709);
xnor UO_575 (O_575,N_13856,N_13992);
or UO_576 (O_576,N_12342,N_14907);
or UO_577 (O_577,N_13383,N_13474);
xor UO_578 (O_578,N_12429,N_12658);
or UO_579 (O_579,N_13616,N_14448);
nand UO_580 (O_580,N_12183,N_13042);
or UO_581 (O_581,N_13645,N_14596);
nand UO_582 (O_582,N_13515,N_12461);
or UO_583 (O_583,N_14852,N_12387);
nor UO_584 (O_584,N_13761,N_13738);
nor UO_585 (O_585,N_13106,N_13023);
nand UO_586 (O_586,N_14880,N_14123);
nor UO_587 (O_587,N_12008,N_13677);
nor UO_588 (O_588,N_12881,N_14064);
or UO_589 (O_589,N_13121,N_14650);
xnor UO_590 (O_590,N_13152,N_12500);
xnor UO_591 (O_591,N_12415,N_13505);
nor UO_592 (O_592,N_12543,N_14716);
or UO_593 (O_593,N_14329,N_14737);
xor UO_594 (O_594,N_14969,N_12092);
and UO_595 (O_595,N_14310,N_14037);
xnor UO_596 (O_596,N_12695,N_14376);
or UO_597 (O_597,N_12085,N_13688);
nor UO_598 (O_598,N_12863,N_14725);
xor UO_599 (O_599,N_12224,N_13127);
nand UO_600 (O_600,N_14986,N_14479);
nand UO_601 (O_601,N_14877,N_14022);
nor UO_602 (O_602,N_14794,N_13485);
and UO_603 (O_603,N_12780,N_12398);
nor UO_604 (O_604,N_14639,N_12759);
and UO_605 (O_605,N_13872,N_14331);
and UO_606 (O_606,N_13814,N_14360);
nand UO_607 (O_607,N_13325,N_13573);
or UO_608 (O_608,N_12141,N_14490);
or UO_609 (O_609,N_13318,N_13217);
nand UO_610 (O_610,N_13991,N_14210);
nand UO_611 (O_611,N_14252,N_14372);
nand UO_612 (O_612,N_13159,N_13947);
and UO_613 (O_613,N_14071,N_12353);
nand UO_614 (O_614,N_13790,N_13807);
nand UO_615 (O_615,N_13627,N_13575);
and UO_616 (O_616,N_14757,N_12220);
or UO_617 (O_617,N_13426,N_14800);
or UO_618 (O_618,N_13975,N_13211);
xnor UO_619 (O_619,N_12784,N_12345);
and UO_620 (O_620,N_14947,N_12318);
nand UO_621 (O_621,N_13174,N_12025);
or UO_622 (O_622,N_12909,N_12442);
xnor UO_623 (O_623,N_14150,N_14187);
nor UO_624 (O_624,N_14544,N_12260);
nor UO_625 (O_625,N_12133,N_13815);
or UO_626 (O_626,N_13680,N_13225);
nand UO_627 (O_627,N_12650,N_14767);
nand UO_628 (O_628,N_14517,N_12293);
or UO_629 (O_629,N_12604,N_12835);
and UO_630 (O_630,N_14898,N_13084);
nor UO_631 (O_631,N_12509,N_12916);
nor UO_632 (O_632,N_13468,N_13408);
or UO_633 (O_633,N_13438,N_13448);
nor UO_634 (O_634,N_14393,N_12808);
xnor UO_635 (O_635,N_12282,N_14106);
and UO_636 (O_636,N_13574,N_12689);
and UO_637 (O_637,N_14200,N_14290);
or UO_638 (O_638,N_12457,N_13012);
nor UO_639 (O_639,N_13080,N_14883);
nand UO_640 (O_640,N_12392,N_12809);
nor UO_641 (O_641,N_12554,N_13118);
and UO_642 (O_642,N_13480,N_14247);
nand UO_643 (O_643,N_14601,N_14841);
or UO_644 (O_644,N_12401,N_13967);
nand UO_645 (O_645,N_14126,N_13043);
and UO_646 (O_646,N_14464,N_13301);
nand UO_647 (O_647,N_14866,N_12292);
nor UO_648 (O_648,N_14615,N_13265);
nand UO_649 (O_649,N_12920,N_12198);
nand UO_650 (O_650,N_13874,N_12184);
or UO_651 (O_651,N_13638,N_12006);
nand UO_652 (O_652,N_12418,N_12486);
nand UO_653 (O_653,N_12414,N_13718);
and UO_654 (O_654,N_14186,N_13125);
or UO_655 (O_655,N_13109,N_14774);
and UO_656 (O_656,N_12934,N_14764);
xnor UO_657 (O_657,N_14575,N_12351);
and UO_658 (O_658,N_12315,N_13903);
or UO_659 (O_659,N_13961,N_14913);
and UO_660 (O_660,N_14198,N_12963);
nand UO_661 (O_661,N_14452,N_13750);
nor UO_662 (O_662,N_12372,N_12472);
or UO_663 (O_663,N_14038,N_12688);
or UO_664 (O_664,N_13370,N_13709);
nand UO_665 (O_665,N_12538,N_14109);
and UO_666 (O_666,N_14870,N_12051);
or UO_667 (O_667,N_13348,N_14092);
and UO_668 (O_668,N_12238,N_12376);
and UO_669 (O_669,N_12290,N_12729);
and UO_670 (O_670,N_13062,N_12330);
nor UO_671 (O_671,N_14459,N_13355);
nand UO_672 (O_672,N_13916,N_12074);
xnor UO_673 (O_673,N_12823,N_13777);
nand UO_674 (O_674,N_13995,N_12076);
xor UO_675 (O_675,N_13343,N_14529);
nor UO_676 (O_676,N_12455,N_12965);
or UO_677 (O_677,N_12541,N_12034);
xor UO_678 (O_678,N_13339,N_12482);
xor UO_679 (O_679,N_14671,N_13294);
nand UO_680 (O_680,N_13381,N_14311);
or UO_681 (O_681,N_14524,N_14222);
and UO_682 (O_682,N_14937,N_12252);
nand UO_683 (O_683,N_12849,N_13226);
nand UO_684 (O_684,N_12403,N_14932);
nor UO_685 (O_685,N_12244,N_14110);
nor UO_686 (O_686,N_13906,N_13452);
nand UO_687 (O_687,N_13376,N_12229);
and UO_688 (O_688,N_14566,N_13817);
xor UO_689 (O_689,N_14033,N_12912);
nand UO_690 (O_690,N_14740,N_13763);
nand UO_691 (O_691,N_13196,N_14685);
xnor UO_692 (O_692,N_13686,N_13804);
nor UO_693 (O_693,N_13501,N_13103);
and UO_694 (O_694,N_14465,N_13891);
or UO_695 (O_695,N_13977,N_12562);
nand UO_696 (O_696,N_14264,N_12896);
or UO_697 (O_697,N_14567,N_14949);
or UO_698 (O_698,N_12721,N_13151);
and UO_699 (O_699,N_13441,N_13508);
nand UO_700 (O_700,N_12055,N_14582);
nand UO_701 (O_701,N_14160,N_13865);
nand UO_702 (O_702,N_14137,N_14368);
nor UO_703 (O_703,N_14798,N_13169);
nor UO_704 (O_704,N_13179,N_14902);
or UO_705 (O_705,N_13685,N_14559);
nor UO_706 (O_706,N_13230,N_13983);
or UO_707 (O_707,N_13367,N_13181);
and UO_708 (O_708,N_14666,N_13783);
nor UO_709 (O_709,N_13063,N_14498);
or UO_710 (O_710,N_13521,N_12464);
or UO_711 (O_711,N_14304,N_12172);
and UO_712 (O_712,N_14897,N_13960);
or UO_713 (O_713,N_13551,N_13456);
or UO_714 (O_714,N_14384,N_12187);
or UO_715 (O_715,N_14696,N_12769);
and UO_716 (O_716,N_13613,N_13246);
nand UO_717 (O_717,N_13366,N_14541);
nand UO_718 (O_718,N_12573,N_14101);
or UO_719 (O_719,N_13072,N_12100);
nand UO_720 (O_720,N_13177,N_14714);
xor UO_721 (O_721,N_13743,N_13822);
xnor UO_722 (O_722,N_12918,N_13518);
or UO_723 (O_723,N_12091,N_13914);
or UO_724 (O_724,N_14111,N_14849);
nor UO_725 (O_725,N_12705,N_14428);
nand UO_726 (O_726,N_13546,N_13819);
xnor UO_727 (O_727,N_12333,N_12193);
or UO_728 (O_728,N_12128,N_12065);
nor UO_729 (O_729,N_13150,N_14690);
nor UO_730 (O_730,N_12567,N_12649);
xnor UO_731 (O_731,N_13553,N_13628);
nor UO_732 (O_732,N_12045,N_12568);
nand UO_733 (O_733,N_14417,N_14166);
or UO_734 (O_734,N_13674,N_14661);
nor UO_735 (O_735,N_13418,N_14118);
or UO_736 (O_736,N_14682,N_14316);
nor UO_737 (O_737,N_14688,N_13281);
or UO_738 (O_738,N_14537,N_13053);
nand UO_739 (O_739,N_14260,N_14742);
nor UO_740 (O_740,N_12812,N_13188);
nor UO_741 (O_741,N_13840,N_12467);
and UO_742 (O_742,N_13620,N_14703);
xor UO_743 (O_743,N_14487,N_13393);
nor UO_744 (O_744,N_14059,N_14923);
nand UO_745 (O_745,N_12360,N_13429);
nor UO_746 (O_746,N_14446,N_12986);
and UO_747 (O_747,N_13161,N_14856);
xnor UO_748 (O_748,N_14728,N_13093);
nor UO_749 (O_749,N_13519,N_14466);
nand UO_750 (O_750,N_14047,N_12267);
xor UO_751 (O_751,N_13337,N_12256);
and UO_752 (O_752,N_13915,N_14660);
and UO_753 (O_753,N_14019,N_12334);
and UO_754 (O_754,N_13577,N_12537);
nor UO_755 (O_755,N_12875,N_14267);
xnor UO_756 (O_756,N_12620,N_12138);
nand UO_757 (O_757,N_13302,N_12762);
nor UO_758 (O_758,N_14697,N_13732);
nor UO_759 (O_759,N_13996,N_14759);
and UO_760 (O_760,N_13528,N_13939);
nand UO_761 (O_761,N_14558,N_14321);
xnor UO_762 (O_762,N_13329,N_12931);
nor UO_763 (O_763,N_13811,N_13419);
nand UO_764 (O_764,N_13614,N_13957);
or UO_765 (O_765,N_13936,N_13956);
nand UO_766 (O_766,N_14980,N_12929);
nand UO_767 (O_767,N_13857,N_14248);
xor UO_768 (O_768,N_13942,N_13892);
and UO_769 (O_769,N_13463,N_14903);
nor UO_770 (O_770,N_12941,N_12599);
and UO_771 (O_771,N_14382,N_14054);
nand UO_772 (O_772,N_14831,N_12788);
and UO_773 (O_773,N_12437,N_12383);
and UO_774 (O_774,N_14546,N_13704);
and UO_775 (O_775,N_14503,N_14785);
nor UO_776 (O_776,N_14927,N_12348);
nor UO_777 (O_777,N_12212,N_13678);
and UO_778 (O_778,N_12884,N_12895);
and UO_779 (O_779,N_12505,N_13178);
nand UO_780 (O_780,N_12525,N_14365);
nor UO_781 (O_781,N_13687,N_12137);
or UO_782 (O_782,N_12961,N_13713);
nand UO_783 (O_783,N_14430,N_13958);
nand UO_784 (O_784,N_14273,N_12477);
and UO_785 (O_785,N_12434,N_13904);
and UO_786 (O_786,N_12939,N_12652);
xor UO_787 (O_787,N_14965,N_12200);
nand UO_788 (O_788,N_14327,N_14520);
nand UO_789 (O_789,N_13540,N_13837);
and UO_790 (O_790,N_14548,N_12610);
or UO_791 (O_791,N_14115,N_14340);
and UO_792 (O_792,N_12669,N_12119);
and UO_793 (O_793,N_14377,N_14196);
or UO_794 (O_794,N_12847,N_12059);
nand UO_795 (O_795,N_12679,N_14407);
nor UO_796 (O_796,N_13651,N_14700);
xnor UO_797 (O_797,N_12121,N_14822);
nand UO_798 (O_798,N_12443,N_14184);
nor UO_799 (O_799,N_14387,N_14480);
and UO_800 (O_800,N_12251,N_13581);
and UO_801 (O_801,N_14922,N_12347);
and UO_802 (O_802,N_13183,N_13222);
and UO_803 (O_803,N_12404,N_13923);
or UO_804 (O_804,N_14277,N_13332);
or UO_805 (O_805,N_13838,N_12684);
nand UO_806 (O_806,N_14637,N_13435);
nand UO_807 (O_807,N_12732,N_12887);
xor UO_808 (O_808,N_12201,N_14338);
xnor UO_809 (O_809,N_13742,N_14471);
and UO_810 (O_810,N_14649,N_12814);
or UO_811 (O_811,N_13481,N_13491);
nor UO_812 (O_812,N_12107,N_13280);
or UO_813 (O_813,N_12105,N_12249);
nor UO_814 (O_814,N_12953,N_14433);
or UO_815 (O_815,N_12872,N_14501);
and UO_816 (O_816,N_14591,N_14108);
nor UO_817 (O_817,N_14371,N_13846);
and UO_818 (O_818,N_13879,N_12284);
and UO_819 (O_819,N_12846,N_12170);
and UO_820 (O_820,N_14987,N_12861);
and UO_821 (O_821,N_13825,N_14188);
xor UO_822 (O_822,N_12685,N_13131);
xor UO_823 (O_823,N_14351,N_12845);
nor UO_824 (O_824,N_14475,N_14620);
nor UO_825 (O_825,N_14772,N_12352);
xnor UO_826 (O_826,N_14203,N_12015);
and UO_827 (O_827,N_12981,N_13786);
nor UO_828 (O_828,N_14677,N_13606);
and UO_829 (O_829,N_12081,N_14906);
xor UO_830 (O_830,N_13488,N_14307);
nand UO_831 (O_831,N_13940,N_14478);
nand UO_832 (O_832,N_12340,N_13695);
or UO_833 (O_833,N_14646,N_14438);
xnor UO_834 (O_834,N_14613,N_14747);
nand UO_835 (O_835,N_13214,N_12499);
or UO_836 (O_836,N_13087,N_12419);
nand UO_837 (O_837,N_13550,N_12569);
nand UO_838 (O_838,N_14112,N_13440);
nand UO_839 (O_839,N_12944,N_14325);
nor UO_840 (O_840,N_12745,N_12235);
and UO_841 (O_841,N_14416,N_12740);
or UO_842 (O_842,N_13504,N_14745);
nor UO_843 (O_843,N_12886,N_14020);
or UO_844 (O_844,N_12385,N_14349);
nor UO_845 (O_845,N_14850,N_12320);
nand UO_846 (O_846,N_13040,N_12800);
and UO_847 (O_847,N_14972,N_13897);
and UO_848 (O_848,N_13705,N_14673);
nand UO_849 (O_849,N_14766,N_13437);
or UO_850 (O_850,N_12152,N_12822);
nor UO_851 (O_851,N_12018,N_14605);
and UO_852 (O_852,N_13563,N_14564);
nand UO_853 (O_853,N_14129,N_14231);
nand UO_854 (O_854,N_14374,N_13321);
nand UO_855 (O_855,N_13911,N_14460);
or UO_856 (O_856,N_13720,N_13073);
or UO_857 (O_857,N_14686,N_13380);
nor UO_858 (O_858,N_13712,N_13170);
nand UO_859 (O_859,N_14861,N_14216);
xor UO_860 (O_860,N_14729,N_13576);
nand UO_861 (O_861,N_12452,N_12261);
and UO_862 (O_862,N_12354,N_12819);
nor UO_863 (O_863,N_13141,N_12177);
nor UO_864 (O_864,N_13845,N_13160);
and UO_865 (O_865,N_13928,N_14507);
and UO_866 (O_866,N_13186,N_14946);
nand UO_867 (O_867,N_12033,N_13885);
and UO_868 (O_868,N_14455,N_14028);
or UO_869 (O_869,N_13443,N_14253);
nand UO_870 (O_870,N_12478,N_13726);
nand UO_871 (O_871,N_14638,N_13233);
and UO_872 (O_872,N_12519,N_14024);
nand UO_873 (O_873,N_13866,N_12785);
nand UO_874 (O_874,N_13244,N_14172);
nand UO_875 (O_875,N_12571,N_14195);
or UO_876 (O_876,N_12892,N_12111);
nand UO_877 (O_877,N_12583,N_13218);
xnor UO_878 (O_878,N_14128,N_13820);
and UO_879 (O_879,N_14097,N_12767);
nor UO_880 (O_880,N_14309,N_14929);
and UO_881 (O_881,N_12496,N_13054);
xor UO_882 (O_882,N_14874,N_12597);
or UO_883 (O_883,N_13476,N_13530);
xnor UO_884 (O_884,N_14571,N_12494);
and UO_885 (O_885,N_12662,N_13297);
nor UO_886 (O_886,N_13697,N_14405);
nand UO_887 (O_887,N_13439,N_14204);
or UO_888 (O_888,N_13827,N_12675);
or UO_889 (O_889,N_12988,N_13506);
or UO_890 (O_890,N_13335,N_14421);
nor UO_891 (O_891,N_12407,N_14121);
or UO_892 (O_892,N_13420,N_14628);
nor UO_893 (O_893,N_12922,N_12266);
nor UO_894 (O_894,N_14539,N_12180);
or UO_895 (O_895,N_14748,N_12996);
nor UO_896 (O_896,N_14678,N_14998);
and UO_897 (O_897,N_13824,N_12540);
or UO_898 (O_898,N_13902,N_14694);
nand UO_899 (O_899,N_13008,N_12493);
and UO_900 (O_900,N_12890,N_14057);
and UO_901 (O_901,N_13272,N_14847);
xor UO_902 (O_902,N_14182,N_12947);
nand UO_903 (O_903,N_14805,N_12027);
xnor UO_904 (O_904,N_12584,N_12989);
and UO_905 (O_905,N_14808,N_12990);
nor UO_906 (O_906,N_14287,N_12901);
and UO_907 (O_907,N_13661,N_14363);
or UO_908 (O_908,N_14181,N_13341);
nand UO_909 (O_909,N_14011,N_12850);
and UO_910 (O_910,N_12417,N_13324);
and UO_911 (O_911,N_14297,N_14096);
nand UO_912 (O_912,N_13375,N_12014);
nor UO_913 (O_913,N_13765,N_14291);
and UO_914 (O_914,N_14102,N_12790);
and UO_915 (O_915,N_12408,N_12972);
or UO_916 (O_916,N_14719,N_12120);
or UO_917 (O_917,N_12834,N_13292);
nand UO_918 (O_918,N_12724,N_14718);
nand UO_919 (O_919,N_14905,N_14282);
nor UO_920 (O_920,N_14263,N_12984);
nor UO_921 (O_921,N_14483,N_13180);
and UO_922 (O_922,N_14251,N_14283);
xnor UO_923 (O_923,N_13473,N_14383);
and UO_924 (O_924,N_12631,N_13951);
or UO_925 (O_925,N_14442,N_14114);
or UO_926 (O_926,N_12221,N_14684);
and UO_927 (O_927,N_12427,N_14245);
or UO_928 (O_928,N_14865,N_14962);
xor UO_929 (O_929,N_14148,N_14394);
and UO_930 (O_930,N_12023,N_13436);
nand UO_931 (O_931,N_13048,N_13587);
nand UO_932 (O_932,N_12459,N_12149);
nand UO_933 (O_933,N_13197,N_12528);
nand UO_934 (O_934,N_14846,N_14676);
nor UO_935 (O_935,N_12075,N_14704);
nor UO_936 (O_936,N_13736,N_14080);
or UO_937 (O_937,N_14837,N_14422);
nor UO_938 (O_938,N_13288,N_14867);
nand UO_939 (O_939,N_12827,N_14804);
nor UO_940 (O_940,N_12253,N_12974);
nor UO_941 (O_941,N_13799,N_12453);
or UO_942 (O_942,N_14973,N_13360);
or UO_943 (O_943,N_12854,N_13502);
or UO_944 (O_944,N_14440,N_14493);
and UO_945 (O_945,N_12925,N_14143);
nand UO_946 (O_946,N_12026,N_12943);
nor UO_947 (O_947,N_14829,N_12396);
nor UO_948 (O_948,N_14680,N_14067);
and UO_949 (O_949,N_14082,N_12761);
nand UO_950 (O_950,N_12002,N_14099);
or UO_951 (O_951,N_12017,N_14296);
or UO_952 (O_952,N_13467,N_14357);
and UO_953 (O_953,N_12194,N_14306);
xor UO_954 (O_954,N_14021,N_14816);
nor UO_955 (O_955,N_12692,N_12885);
nand UO_956 (O_956,N_12670,N_14610);
and UO_957 (O_957,N_14783,N_12146);
xor UO_958 (O_958,N_13848,N_14518);
nand UO_959 (O_959,N_13571,N_12328);
nor UO_960 (O_960,N_13410,N_12010);
and UO_961 (O_961,N_12926,N_14669);
nand UO_962 (O_962,N_14743,N_12117);
nor UO_963 (O_963,N_14016,N_13425);
nand UO_964 (O_964,N_12676,N_12488);
nor UO_965 (O_965,N_13422,N_12980);
and UO_966 (O_966,N_12703,N_14045);
and UO_967 (O_967,N_12578,N_14899);
xor UO_968 (O_968,N_13775,N_13185);
nand UO_969 (O_969,N_14435,N_14821);
or UO_970 (O_970,N_14240,N_12090);
and UO_971 (O_971,N_13834,N_14918);
xor UO_972 (O_972,N_13629,N_12816);
or UO_973 (O_973,N_12690,N_12369);
or UO_974 (O_974,N_14177,N_13552);
nor UO_975 (O_975,N_14773,N_14780);
nand UO_976 (O_976,N_13130,N_14588);
xor UO_977 (O_977,N_13005,N_13794);
nor UO_978 (O_978,N_12791,N_13895);
nor UO_979 (O_979,N_14458,N_12270);
and UO_980 (O_980,N_12937,N_12420);
xnor UO_981 (O_981,N_13198,N_14916);
or UO_982 (O_982,N_13725,N_12580);
xor UO_983 (O_983,N_13345,N_13858);
xnor UO_984 (O_984,N_14654,N_12083);
nor UO_985 (O_985,N_12593,N_14119);
nor UO_986 (O_986,N_13407,N_12361);
or UO_987 (O_987,N_13432,N_12003);
and UO_988 (O_988,N_12664,N_13402);
and UO_989 (O_989,N_12048,N_12629);
and UO_990 (O_990,N_14403,N_12240);
and UO_991 (O_991,N_12226,N_14224);
nor UO_992 (O_992,N_14573,N_14171);
or UO_993 (O_993,N_12005,N_13821);
and UO_994 (O_994,N_13404,N_13162);
and UO_995 (O_995,N_14227,N_12071);
nand UO_996 (O_996,N_13773,N_13873);
and UO_997 (O_997,N_12968,N_13805);
and UO_998 (O_998,N_13168,N_14557);
nor UO_999 (O_999,N_13600,N_14058);
nand UO_1000 (O_1000,N_12592,N_14041);
nor UO_1001 (O_1001,N_12805,N_12570);
and UO_1002 (O_1002,N_12217,N_14025);
and UO_1003 (O_1003,N_12157,N_14324);
or UO_1004 (O_1004,N_14911,N_13766);
or UO_1005 (O_1005,N_12539,N_13088);
xnor UO_1006 (O_1006,N_12311,N_14328);
or UO_1007 (O_1007,N_13615,N_12526);
and UO_1008 (O_1008,N_14419,N_13513);
xor UO_1009 (O_1009,N_14034,N_14259);
and UO_1010 (O_1010,N_12019,N_14819);
nand UO_1011 (O_1011,N_13365,N_14332);
or UO_1012 (O_1012,N_12402,N_14463);
nor UO_1013 (O_1013,N_12560,N_12955);
nand UO_1014 (O_1014,N_14984,N_13883);
nand UO_1015 (O_1015,N_12734,N_12375);
nor UO_1016 (O_1016,N_14602,N_12797);
nand UO_1017 (O_1017,N_13741,N_14138);
and UO_1018 (O_1018,N_14827,N_14191);
and UO_1019 (O_1019,N_13887,N_14261);
or UO_1020 (O_1020,N_13207,N_13427);
nand UO_1021 (O_1021,N_13760,N_14429);
nand UO_1022 (O_1022,N_14940,N_13562);
xnor UO_1023 (O_1023,N_14149,N_12145);
xnor UO_1024 (O_1024,N_13602,N_13730);
nand UO_1025 (O_1025,N_13269,N_13205);
or UO_1026 (O_1026,N_12135,N_14691);
xnor UO_1027 (O_1027,N_13369,N_14681);
nand UO_1028 (O_1028,N_14423,N_14229);
nor UO_1029 (O_1029,N_14872,N_13201);
nand UO_1030 (O_1030,N_14348,N_14532);
or UO_1031 (O_1031,N_12013,N_12728);
xor UO_1032 (O_1032,N_14473,N_14934);
xor UO_1033 (O_1033,N_12608,N_14223);
nor UO_1034 (O_1034,N_12481,N_14674);
nand UO_1035 (O_1035,N_13517,N_12225);
nand UO_1036 (O_1036,N_13311,N_12645);
nand UO_1037 (O_1037,N_13251,N_13032);
nand UO_1038 (O_1038,N_14220,N_14225);
nand UO_1039 (O_1039,N_13798,N_12497);
nor UO_1040 (O_1040,N_13549,N_14760);
and UO_1041 (O_1041,N_12913,N_12735);
nand UO_1042 (O_1042,N_14342,N_13889);
or UO_1043 (O_1043,N_12727,N_12533);
and UO_1044 (O_1044,N_14236,N_14834);
or UO_1045 (O_1045,N_12687,N_13305);
and UO_1046 (O_1046,N_12468,N_13095);
and UO_1047 (O_1047,N_12607,N_13946);
nor UO_1048 (O_1048,N_12168,N_14702);
nand UO_1049 (O_1049,N_14733,N_14731);
nand UO_1050 (O_1050,N_12618,N_13536);
nor UO_1051 (O_1051,N_12874,N_12862);
or UO_1052 (O_1052,N_13209,N_13876);
xor UO_1053 (O_1053,N_13123,N_14683);
nand UO_1054 (O_1054,N_13921,N_14769);
xnor UO_1055 (O_1055,N_14527,N_14051);
nand UO_1056 (O_1056,N_12016,N_13350);
nand UO_1057 (O_1057,N_13871,N_13933);
or UO_1058 (O_1058,N_14232,N_12450);
and UO_1059 (O_1059,N_13250,N_14049);
nand UO_1060 (O_1060,N_12521,N_12341);
and UO_1061 (O_1061,N_14142,N_12617);
nand UO_1062 (O_1062,N_12706,N_12007);
nor UO_1063 (O_1063,N_13494,N_12445);
and UO_1064 (O_1064,N_13534,N_14925);
nand UO_1065 (O_1065,N_14266,N_14409);
and UO_1066 (O_1066,N_14606,N_13757);
or UO_1067 (O_1067,N_14053,N_12718);
or UO_1068 (O_1068,N_12435,N_12298);
and UO_1069 (O_1069,N_14169,N_14322);
or UO_1070 (O_1070,N_12640,N_12501);
nand UO_1071 (O_1071,N_14873,N_12765);
or UO_1072 (O_1072,N_13249,N_12719);
or UO_1073 (O_1073,N_14803,N_14689);
or UO_1074 (O_1074,N_14006,N_12550);
nor UO_1075 (O_1075,N_14345,N_14242);
nand UO_1076 (O_1076,N_14208,N_12060);
xor UO_1077 (O_1077,N_14550,N_13424);
nor UO_1078 (O_1078,N_12030,N_13759);
nand UO_1079 (O_1079,N_13919,N_14776);
xor UO_1080 (O_1080,N_12004,N_14482);
and UO_1081 (O_1081,N_14672,N_13980);
or UO_1082 (O_1082,N_14131,N_13963);
nor UO_1083 (O_1083,N_13449,N_14185);
xnor UO_1084 (O_1084,N_13457,N_12001);
nor UO_1085 (O_1085,N_12476,N_13356);
and UO_1086 (O_1086,N_13908,N_12274);
nor UO_1087 (O_1087,N_13672,N_12612);
xor UO_1088 (O_1088,N_13556,N_14418);
nor UO_1089 (O_1089,N_14213,N_14778);
or UO_1090 (O_1090,N_14218,N_13066);
nand UO_1091 (O_1091,N_13830,N_14530);
and UO_1092 (O_1092,N_13985,N_13081);
nand UO_1093 (O_1093,N_14985,N_14084);
nand UO_1094 (O_1094,N_13046,N_12665);
or UO_1095 (O_1095,N_14088,N_14255);
nand UO_1096 (O_1096,N_14552,N_14617);
and UO_1097 (O_1097,N_12978,N_14495);
and UO_1098 (O_1098,N_13472,N_12882);
nor UO_1099 (O_1099,N_13634,N_12171);
nor UO_1100 (O_1100,N_13929,N_12259);
xor UO_1101 (O_1101,N_13262,N_12156);
nor UO_1102 (O_1102,N_14779,N_13886);
and UO_1103 (O_1103,N_14692,N_13303);
nor UO_1104 (O_1104,N_12663,N_14470);
and UO_1105 (O_1105,N_14598,N_14930);
and UO_1106 (O_1106,N_12945,N_12441);
nand UO_1107 (O_1107,N_13362,N_14893);
or UO_1108 (O_1108,N_14315,N_13976);
xnor UO_1109 (O_1109,N_12596,N_14472);
and UO_1110 (O_1110,N_12921,N_13862);
nand UO_1111 (O_1111,N_12803,N_13187);
or UO_1112 (O_1112,N_14657,N_14943);
or UO_1113 (O_1113,N_12000,N_14436);
xor UO_1114 (O_1114,N_12192,N_13489);
or UO_1115 (O_1115,N_12994,N_14081);
and UO_1116 (O_1116,N_12098,N_13772);
nor UO_1117 (O_1117,N_13702,N_13539);
nor UO_1118 (O_1118,N_12483,N_13039);
nand UO_1119 (O_1119,N_12178,N_14931);
nand UO_1120 (O_1120,N_13068,N_12750);
and UO_1121 (O_1121,N_13558,N_14670);
nand UO_1122 (O_1122,N_14658,N_13306);
nor UO_1123 (O_1123,N_12523,N_13618);
nand UO_1124 (O_1124,N_14477,N_13260);
xor UO_1125 (O_1125,N_12374,N_12189);
or UO_1126 (O_1126,N_13598,N_12624);
and UO_1127 (O_1127,N_14545,N_14280);
nor UO_1128 (O_1128,N_12009,N_12954);
nand UO_1129 (O_1129,N_12485,N_14668);
and UO_1130 (O_1130,N_12041,N_13077);
nor UO_1131 (O_1131,N_14832,N_14469);
or UO_1132 (O_1132,N_14775,N_13253);
nand UO_1133 (O_1133,N_13691,N_13768);
xnor UO_1134 (O_1134,N_13493,N_14762);
nand UO_1135 (O_1135,N_12572,N_12677);
nand UO_1136 (O_1136,N_12548,N_13357);
and UO_1137 (O_1137,N_14176,N_13085);
or UO_1138 (O_1138,N_12976,N_12386);
nor UO_1139 (O_1139,N_12425,N_13024);
and UO_1140 (O_1140,N_12940,N_13572);
xor UO_1141 (O_1141,N_12993,N_12112);
nor UO_1142 (O_1142,N_14618,N_14983);
nand UO_1143 (O_1143,N_12962,N_12064);
nor UO_1144 (O_1144,N_12093,N_14281);
or UO_1145 (O_1145,N_12726,N_13986);
nor UO_1146 (O_1146,N_12126,N_12491);
nand UO_1147 (O_1147,N_12626,N_14107);
nand UO_1148 (O_1148,N_12232,N_12050);
nand UO_1149 (O_1149,N_12241,N_13256);
nor UO_1150 (O_1150,N_13753,N_12086);
xnor UO_1151 (O_1151,N_13644,N_12504);
xor UO_1152 (O_1152,N_12367,N_12182);
and UO_1153 (O_1153,N_13931,N_12151);
or UO_1154 (O_1154,N_12439,N_13586);
and UO_1155 (O_1155,N_14979,N_14012);
nor UO_1156 (O_1156,N_12632,N_12643);
or UO_1157 (O_1157,N_13707,N_12894);
or UO_1158 (O_1158,N_12579,N_13334);
or UO_1159 (O_1159,N_12595,N_12096);
xor UO_1160 (O_1160,N_12907,N_13869);
and UO_1161 (O_1161,N_12644,N_13962);
nor UO_1162 (O_1162,N_14636,N_14337);
and UO_1163 (O_1163,N_12469,N_13395);
nand UO_1164 (O_1164,N_13102,N_12116);
or UO_1165 (O_1165,N_13767,N_12956);
or UO_1166 (O_1166,N_12950,N_14063);
nand UO_1167 (O_1167,N_14875,N_12967);
or UO_1168 (O_1168,N_14303,N_14174);
and UO_1169 (O_1169,N_14001,N_13912);
nand UO_1170 (O_1170,N_13560,N_13589);
nand UO_1171 (O_1171,N_13284,N_14199);
nor UO_1172 (O_1172,N_14624,N_12870);
nor UO_1173 (O_1173,N_12104,N_13133);
and UO_1174 (O_1174,N_14437,N_13078);
and UO_1175 (O_1175,N_12927,N_12489);
and UO_1176 (O_1176,N_12614,N_14635);
xor UO_1177 (O_1177,N_12242,N_13588);
xnor UO_1178 (O_1178,N_12933,N_12438);
nor UO_1179 (O_1179,N_14562,N_13320);
nor UO_1180 (O_1180,N_12900,N_13664);
nor UO_1181 (O_1181,N_13945,N_13592);
or UO_1182 (O_1182,N_13789,N_12866);
nor UO_1183 (O_1183,N_12905,N_13523);
nand UO_1184 (O_1184,N_12544,N_12751);
and UO_1185 (O_1185,N_13344,N_14533);
or UO_1186 (O_1186,N_14256,N_12589);
nor UO_1187 (O_1187,N_13657,N_12686);
and UO_1188 (O_1188,N_13044,N_14950);
and UO_1189 (O_1189,N_14881,N_13459);
and UO_1190 (O_1190,N_12069,N_14823);
or UO_1191 (O_1191,N_13475,N_13537);
nor UO_1192 (O_1192,N_12382,N_12012);
nand UO_1193 (O_1193,N_12410,N_14154);
or UO_1194 (O_1194,N_14871,N_12028);
and UO_1195 (O_1195,N_12960,N_13382);
nor UO_1196 (O_1196,N_13323,N_13210);
and UO_1197 (O_1197,N_13374,N_13433);
nand UO_1198 (O_1198,N_13242,N_12807);
nand UO_1199 (O_1199,N_13859,N_14787);
or UO_1200 (O_1200,N_12020,N_14917);
or UO_1201 (O_1201,N_13215,N_14312);
and UO_1202 (O_1202,N_13034,N_13752);
xnor UO_1203 (O_1203,N_12712,N_12110);
or UO_1204 (O_1204,N_12829,N_14859);
xnor UO_1205 (O_1205,N_13378,N_14300);
or UO_1206 (O_1206,N_12174,N_12148);
and UO_1207 (O_1207,N_12066,N_13002);
nor UO_1208 (O_1208,N_13579,N_14445);
nor UO_1209 (O_1209,N_14522,N_14085);
nand UO_1210 (O_1210,N_14050,N_14958);
xor UO_1211 (O_1211,N_12377,N_14305);
nor UO_1212 (O_1212,N_13111,N_13776);
nor UO_1213 (O_1213,N_13541,N_12810);
or UO_1214 (O_1214,N_12391,N_14233);
nor UO_1215 (O_1215,N_13495,N_12389);
nand UO_1216 (O_1216,N_13257,N_13124);
and UO_1217 (O_1217,N_13190,N_14569);
xnor UO_1218 (O_1218,N_14892,N_14525);
nor UO_1219 (O_1219,N_12615,N_13004);
nand UO_1220 (O_1220,N_12581,N_14820);
and UO_1221 (O_1221,N_12109,N_14549);
nor UO_1222 (O_1222,N_12046,N_12838);
and UO_1223 (O_1223,N_14944,N_14506);
and UO_1224 (O_1224,N_12786,N_14510);
xor UO_1225 (O_1225,N_12214,N_13057);
or UO_1226 (O_1226,N_14100,N_12070);
xor UO_1227 (O_1227,N_13028,N_14555);
or UO_1228 (O_1228,N_13643,N_13041);
nor UO_1229 (O_1229,N_13681,N_14103);
nor UO_1230 (O_1230,N_13608,N_12633);
nand UO_1231 (O_1231,N_12772,N_14951);
or UO_1232 (O_1232,N_12552,N_12651);
and UO_1233 (O_1233,N_12078,N_14193);
nand UO_1234 (O_1234,N_14715,N_12666);
nor UO_1235 (O_1235,N_14145,N_12307);
and UO_1236 (O_1236,N_12923,N_14891);
and UO_1237 (O_1237,N_14782,N_12031);
or UO_1238 (O_1238,N_13769,N_13890);
and UO_1239 (O_1239,N_12299,N_14358);
nand UO_1240 (O_1240,N_13954,N_12574);
or UO_1241 (O_1241,N_12161,N_12799);
nand UO_1242 (O_1242,N_13836,N_12899);
nand UO_1243 (O_1243,N_14411,N_14964);
and UO_1244 (O_1244,N_13184,N_12160);
nand UO_1245 (O_1245,N_13952,N_12707);
nand UO_1246 (O_1246,N_14265,N_12269);
and UO_1247 (O_1247,N_14320,N_13706);
and UO_1248 (O_1248,N_12454,N_13083);
or UO_1249 (O_1249,N_14508,N_12565);
nor UO_1250 (O_1250,N_12062,N_13025);
or UO_1251 (O_1251,N_13398,N_13450);
xor UO_1252 (O_1252,N_13176,N_14885);
and UO_1253 (O_1253,N_12204,N_13394);
nand UO_1254 (O_1254,N_12999,N_13145);
and UO_1255 (O_1255,N_12463,N_13038);
nand UO_1256 (O_1256,N_12139,N_13648);
and UO_1257 (O_1257,N_14484,N_12159);
and UO_1258 (O_1258,N_13875,N_13241);
nand UO_1259 (O_1259,N_12263,N_14496);
and UO_1260 (O_1260,N_12983,N_13860);
nand UO_1261 (O_1261,N_13659,N_13399);
nor UO_1262 (O_1262,N_13612,N_14399);
and UO_1263 (O_1263,N_14828,N_13693);
and UO_1264 (O_1264,N_14799,N_14724);
nand UO_1265 (O_1265,N_13268,N_12199);
and UO_1266 (O_1266,N_12346,N_13624);
or UO_1267 (O_1267,N_13229,N_12368);
or UO_1268 (O_1268,N_12036,N_13882);
and UO_1269 (O_1269,N_12451,N_14030);
and UO_1270 (O_1270,N_12869,N_12044);
nor UO_1271 (O_1271,N_12115,N_14802);
and UO_1272 (O_1272,N_14197,N_14953);
nor UO_1273 (O_1273,N_12303,N_12557);
nand UO_1274 (O_1274,N_12022,N_13682);
xnor UO_1275 (O_1275,N_14457,N_14543);
or UO_1276 (O_1276,N_14512,N_13594);
nand UO_1277 (O_1277,N_13596,N_14840);
and UO_1278 (O_1278,N_14698,N_13953);
or UO_1279 (O_1279,N_12163,N_13212);
or UO_1280 (O_1280,N_12431,N_14513);
xor UO_1281 (O_1281,N_13797,N_13261);
xor UO_1282 (O_1282,N_13405,N_13649);
nor UO_1283 (O_1283,N_13274,N_12130);
xor UO_1284 (O_1284,N_12591,N_14326);
nor UO_1285 (O_1285,N_14073,N_13134);
or UO_1286 (O_1286,N_13451,N_14813);
nor UO_1287 (O_1287,N_14981,N_12630);
nand UO_1288 (O_1288,N_13937,N_12820);
nand UO_1289 (O_1289,N_14426,N_14838);
nand UO_1290 (O_1290,N_12247,N_14194);
xnor UO_1291 (O_1291,N_13308,N_13745);
or UO_1292 (O_1292,N_14175,N_14534);
nor UO_1293 (O_1293,N_12763,N_14402);
xor UO_1294 (O_1294,N_13431,N_13076);
nand UO_1295 (O_1295,N_13813,N_13312);
and UO_1296 (O_1296,N_14221,N_14344);
and UO_1297 (O_1297,N_13411,N_12277);
and UO_1298 (O_1298,N_12332,N_14072);
nor UO_1299 (O_1299,N_12991,N_13051);
nand UO_1300 (O_1300,N_12101,N_14212);
and UO_1301 (O_1301,N_12507,N_12449);
nor UO_1302 (O_1302,N_12783,N_14960);
or UO_1303 (O_1303,N_12394,N_13235);
or UO_1304 (O_1304,N_14301,N_12639);
nand UO_1305 (O_1305,N_12108,N_13582);
xnor UO_1306 (O_1306,N_14570,N_12966);
nor UO_1307 (O_1307,N_12502,N_13351);
nand UO_1308 (O_1308,N_12338,N_13793);
or UO_1309 (O_1309,N_14781,N_12871);
nor UO_1310 (O_1310,N_12082,N_13531);
or UO_1311 (O_1311,N_12914,N_12646);
nor UO_1312 (O_1312,N_12447,N_14098);
nor UO_1313 (O_1313,N_13910,N_14763);
nand UO_1314 (O_1314,N_13195,N_14136);
nor UO_1315 (O_1315,N_12621,N_13403);
nand UO_1316 (O_1316,N_12422,N_14356);
xor UO_1317 (O_1317,N_13128,N_14830);
and UO_1318 (O_1318,N_12975,N_12362);
or UO_1319 (O_1319,N_14133,N_12053);
nand UO_1320 (O_1320,N_12343,N_12545);
and UO_1321 (O_1321,N_12623,N_12717);
nand UO_1322 (O_1322,N_14135,N_13136);
nand UO_1323 (O_1323,N_12880,N_12239);
nor UO_1324 (O_1324,N_12777,N_12513);
and UO_1325 (O_1325,N_12542,N_12602);
xor UO_1326 (O_1326,N_12359,N_13447);
nand UO_1327 (O_1327,N_14938,N_13104);
or UO_1328 (O_1328,N_13033,N_14375);
nand UO_1329 (O_1329,N_12534,N_13867);
nor UO_1330 (O_1330,N_12561,N_14948);
and UO_1331 (O_1331,N_12826,N_13193);
nand UO_1332 (O_1332,N_14540,N_14659);
and UO_1333 (O_1333,N_12166,N_14623);
nand UO_1334 (O_1334,N_13388,N_14997);
and UO_1335 (O_1335,N_14604,N_14350);
xnor UO_1336 (O_1336,N_13611,N_14094);
and UO_1337 (O_1337,N_14369,N_12766);
nor UO_1338 (O_1338,N_13342,N_14044);
xor UO_1339 (O_1339,N_13228,N_12047);
nor UO_1340 (O_1340,N_12852,N_12409);
or UO_1341 (O_1341,N_13729,N_12301);
nor UO_1342 (O_1342,N_12406,N_12294);
and UO_1343 (O_1343,N_13069,N_13227);
or UO_1344 (O_1344,N_12052,N_12113);
nand UO_1345 (O_1345,N_14595,N_13200);
nor UO_1346 (O_1346,N_12233,N_13863);
nand UO_1347 (O_1347,N_13880,N_13969);
or UO_1348 (O_1348,N_13137,N_13623);
and UO_1349 (O_1349,N_12813,N_14390);
or UO_1350 (O_1350,N_14574,N_12691);
and UO_1351 (O_1351,N_12598,N_13998);
xnor UO_1352 (O_1352,N_12127,N_13601);
or UO_1353 (O_1353,N_13861,N_14239);
nand UO_1354 (O_1354,N_13236,N_12275);
nand UO_1355 (O_1355,N_13930,N_13461);
nor UO_1356 (O_1356,N_12234,N_14389);
or UO_1357 (O_1357,N_14086,N_14988);
or UO_1358 (O_1358,N_13617,N_12393);
nor UO_1359 (O_1359,N_14347,N_12998);
or UO_1360 (O_1360,N_14687,N_12412);
or UO_1361 (O_1361,N_13655,N_12749);
and UO_1362 (O_1362,N_12197,N_13199);
and UO_1363 (O_1363,N_12258,N_12458);
and UO_1364 (O_1364,N_12280,N_12388);
or UO_1365 (O_1365,N_12158,N_13667);
or UO_1366 (O_1366,N_14408,N_13604);
nor UO_1367 (O_1367,N_13097,N_13011);
or UO_1368 (O_1368,N_13082,N_12516);
nor UO_1369 (O_1369,N_14366,N_13796);
nand UO_1370 (O_1370,N_13924,N_13067);
nand UO_1371 (O_1371,N_13492,N_14592);
nor UO_1372 (O_1372,N_12851,N_14727);
nor UO_1373 (O_1373,N_13826,N_14625);
nor UO_1374 (O_1374,N_12173,N_14619);
or UO_1375 (O_1375,N_13984,N_13982);
or UO_1376 (O_1376,N_12400,N_13658);
or UO_1377 (O_1377,N_14675,N_14497);
nor UO_1378 (O_1378,N_12635,N_12524);
nor UO_1379 (O_1379,N_12841,N_14811);
xor UO_1380 (O_1380,N_13968,N_14388);
nand UO_1381 (O_1381,N_14594,N_13108);
nand UO_1382 (O_1382,N_12693,N_14134);
and UO_1383 (O_1383,N_14060,N_12316);
and UO_1384 (O_1384,N_14815,N_13823);
and UO_1385 (O_1385,N_14999,N_14642);
nor UO_1386 (O_1386,N_14209,N_14090);
and UO_1387 (O_1387,N_13164,N_14207);
and UO_1388 (O_1388,N_13400,N_14206);
or UO_1389 (O_1389,N_12397,N_12517);
xnor UO_1390 (O_1390,N_12271,N_12154);
xnor UO_1391 (O_1391,N_12147,N_12979);
and UO_1392 (O_1392,N_14055,N_13090);
or UO_1393 (O_1393,N_13240,N_13454);
or UO_1394 (O_1394,N_14005,N_13723);
nand UO_1395 (O_1395,N_12730,N_13844);
nand UO_1396 (O_1396,N_13055,N_13938);
or UO_1397 (O_1397,N_13578,N_12977);
xor UO_1398 (O_1398,N_14523,N_12236);
or UO_1399 (O_1399,N_13387,N_12755);
and UO_1400 (O_1400,N_12072,N_13000);
nor UO_1401 (O_1401,N_13462,N_14720);
or UO_1402 (O_1402,N_14083,N_13496);
or UO_1403 (O_1403,N_12673,N_13988);
nor UO_1404 (O_1404,N_13245,N_13359);
or UO_1405 (O_1405,N_13884,N_12276);
nand UO_1406 (O_1406,N_12804,N_14362);
nand UO_1407 (O_1407,N_12185,N_14924);
xor UO_1408 (O_1408,N_12479,N_13444);
xor UO_1409 (O_1409,N_14789,N_13653);
xnor UO_1410 (O_1410,N_13710,N_13816);
or UO_1411 (O_1411,N_14531,N_14449);
or UO_1412 (O_1412,N_12300,N_13567);
nor UO_1413 (O_1413,N_13158,N_14713);
xnor UO_1414 (O_1414,N_13696,N_14942);
nand UO_1415 (O_1415,N_14048,N_14887);
or UO_1416 (O_1416,N_12997,N_13609);
xor UO_1417 (O_1417,N_13221,N_13699);
nand UO_1418 (O_1418,N_12836,N_13017);
nor UO_1419 (O_1419,N_14039,N_14561);
nand UO_1420 (O_1420,N_13641,N_14584);
nand UO_1421 (O_1421,N_13868,N_14173);
or UO_1422 (O_1422,N_13060,N_14627);
xnor UO_1423 (O_1423,N_12231,N_12433);
nor UO_1424 (O_1424,N_12228,N_13278);
and UO_1425 (O_1425,N_14928,N_13835);
nor UO_1426 (O_1426,N_13428,N_14810);
and UO_1427 (O_1427,N_13006,N_13853);
nor UO_1428 (O_1428,N_13700,N_13224);
nand UO_1429 (O_1429,N_13330,N_12655);
or UO_1430 (O_1430,N_14876,N_12511);
or UO_1431 (O_1431,N_12436,N_13490);
and UO_1432 (O_1432,N_14278,N_13818);
and UO_1433 (O_1433,N_13277,N_14065);
nand UO_1434 (O_1434,N_13711,N_13239);
and UO_1435 (O_1435,N_13114,N_14945);
and UO_1436 (O_1436,N_12741,N_12843);
or UO_1437 (O_1437,N_14013,N_14288);
and UO_1438 (O_1438,N_12758,N_12262);
nand UO_1439 (O_1439,N_13901,N_13019);
nor UO_1440 (O_1440,N_13036,N_13870);
nand UO_1441 (O_1441,N_13430,N_13894);
nand UO_1442 (O_1442,N_14842,N_13510);
nand UO_1443 (O_1443,N_12853,N_12331);
and UO_1444 (O_1444,N_14105,N_13514);
nor UO_1445 (O_1445,N_12337,N_13913);
nand UO_1446 (O_1446,N_12930,N_13703);
or UO_1447 (O_1447,N_13666,N_14791);
and UO_1448 (O_1448,N_14750,N_14560);
nor UO_1449 (O_1449,N_14391,N_14010);
nand UO_1450 (O_1450,N_13762,N_14589);
nor UO_1451 (O_1451,N_13557,N_14599);
and UO_1452 (O_1452,N_13386,N_13689);
xnor UO_1453 (O_1453,N_12904,N_13331);
nor UO_1454 (O_1454,N_14920,N_13964);
and UO_1455 (O_1455,N_14190,N_12150);
nand UO_1456 (O_1456,N_14254,N_12363);
or UO_1457 (O_1457,N_13029,N_14790);
nand UO_1458 (O_1458,N_14292,N_12466);
nor UO_1459 (O_1459,N_13679,N_13801);
and UO_1460 (O_1460,N_13650,N_12304);
or UO_1461 (O_1461,N_14352,N_12587);
nand UO_1462 (O_1462,N_14317,N_12556);
nor UO_1463 (O_1463,N_14796,N_12789);
or UO_1464 (O_1464,N_14279,N_12959);
and UO_1465 (O_1465,N_14788,N_13739);
and UO_1466 (O_1466,N_14286,N_12867);
xor UO_1467 (O_1467,N_13037,N_13780);
or UO_1468 (O_1468,N_12794,N_14741);
nand UO_1469 (O_1469,N_12365,N_13525);
or UO_1470 (O_1470,N_14726,N_12698);
nand UO_1471 (O_1471,N_12551,N_13479);
and UO_1472 (O_1472,N_14989,N_12656);
nand UO_1473 (O_1473,N_14089,N_13070);
nor UO_1474 (O_1474,N_13406,N_12782);
xor UO_1475 (O_1475,N_14373,N_13683);
nand UO_1476 (O_1476,N_12844,N_12681);
or UO_1477 (O_1477,N_14504,N_13401);
nand UO_1478 (O_1478,N_14765,N_12143);
or UO_1479 (O_1479,N_12039,N_12283);
nor UO_1480 (O_1480,N_14878,N_14003);
xor UO_1481 (O_1481,N_12932,N_14026);
and UO_1482 (O_1482,N_12753,N_12473);
nand UO_1483 (O_1483,N_13690,N_13512);
nand UO_1484 (O_1484,N_12876,N_13949);
nand UO_1485 (O_1485,N_14270,N_14758);
or UO_1486 (O_1486,N_13079,N_14499);
nand UO_1487 (O_1487,N_14996,N_12917);
or UO_1488 (O_1488,N_12982,N_14461);
and UO_1489 (O_1489,N_12264,N_14257);
nor UO_1490 (O_1490,N_14580,N_13642);
nor UO_1491 (O_1491,N_12842,N_14289);
or UO_1492 (O_1492,N_13416,N_12399);
or UO_1493 (O_1493,N_14093,N_14380);
or UO_1494 (O_1494,N_12760,N_13778);
nor UO_1495 (O_1495,N_12223,N_13237);
nor UO_1496 (O_1496,N_13192,N_13855);
nand UO_1497 (O_1497,N_12037,N_12430);
xor UO_1498 (O_1498,N_14285,N_12924);
and UO_1499 (O_1499,N_13698,N_14354);
and UO_1500 (O_1500,N_14274,N_12238);
nor UO_1501 (O_1501,N_14163,N_12325);
nor UO_1502 (O_1502,N_13599,N_12826);
or UO_1503 (O_1503,N_12188,N_14033);
xor UO_1504 (O_1504,N_14210,N_12901);
or UO_1505 (O_1505,N_12967,N_12613);
nor UO_1506 (O_1506,N_13708,N_12026);
nor UO_1507 (O_1507,N_14585,N_13864);
nand UO_1508 (O_1508,N_14303,N_14372);
and UO_1509 (O_1509,N_12869,N_13644);
and UO_1510 (O_1510,N_13889,N_12424);
or UO_1511 (O_1511,N_12094,N_14540);
nor UO_1512 (O_1512,N_14649,N_13729);
and UO_1513 (O_1513,N_13079,N_14353);
and UO_1514 (O_1514,N_12943,N_14660);
or UO_1515 (O_1515,N_14796,N_12074);
nor UO_1516 (O_1516,N_12054,N_13345);
nand UO_1517 (O_1517,N_13860,N_14564);
nand UO_1518 (O_1518,N_13119,N_13927);
or UO_1519 (O_1519,N_14966,N_13096);
xnor UO_1520 (O_1520,N_14837,N_12943);
xor UO_1521 (O_1521,N_13595,N_12042);
or UO_1522 (O_1522,N_12879,N_14861);
nor UO_1523 (O_1523,N_13556,N_13442);
and UO_1524 (O_1524,N_12996,N_13711);
xnor UO_1525 (O_1525,N_12934,N_13362);
nor UO_1526 (O_1526,N_13919,N_14205);
nor UO_1527 (O_1527,N_14595,N_13239);
and UO_1528 (O_1528,N_12096,N_13663);
nand UO_1529 (O_1529,N_14708,N_14656);
and UO_1530 (O_1530,N_14975,N_12923);
or UO_1531 (O_1531,N_13314,N_13299);
or UO_1532 (O_1532,N_12019,N_12696);
nor UO_1533 (O_1533,N_12464,N_14985);
xnor UO_1534 (O_1534,N_13277,N_14502);
and UO_1535 (O_1535,N_13541,N_13805);
and UO_1536 (O_1536,N_14030,N_13609);
nor UO_1537 (O_1537,N_14837,N_12700);
nor UO_1538 (O_1538,N_12956,N_12797);
or UO_1539 (O_1539,N_12793,N_13816);
and UO_1540 (O_1540,N_13232,N_14241);
nand UO_1541 (O_1541,N_12919,N_12728);
nand UO_1542 (O_1542,N_14568,N_12687);
nand UO_1543 (O_1543,N_13933,N_14892);
nand UO_1544 (O_1544,N_14492,N_14191);
nor UO_1545 (O_1545,N_13000,N_13489);
and UO_1546 (O_1546,N_14309,N_12270);
nand UO_1547 (O_1547,N_12259,N_12464);
or UO_1548 (O_1548,N_12093,N_12339);
nor UO_1549 (O_1549,N_14749,N_14720);
nand UO_1550 (O_1550,N_13583,N_13852);
xor UO_1551 (O_1551,N_12571,N_14937);
or UO_1552 (O_1552,N_14029,N_12328);
and UO_1553 (O_1553,N_13945,N_12840);
nor UO_1554 (O_1554,N_14770,N_14244);
nand UO_1555 (O_1555,N_13580,N_14855);
or UO_1556 (O_1556,N_12951,N_14747);
nand UO_1557 (O_1557,N_14168,N_14343);
and UO_1558 (O_1558,N_13465,N_13524);
and UO_1559 (O_1559,N_14915,N_14761);
nor UO_1560 (O_1560,N_12087,N_14412);
xnor UO_1561 (O_1561,N_14065,N_12850);
or UO_1562 (O_1562,N_13455,N_13136);
and UO_1563 (O_1563,N_12484,N_13127);
nand UO_1564 (O_1564,N_12278,N_14361);
nor UO_1565 (O_1565,N_14519,N_12936);
xnor UO_1566 (O_1566,N_12631,N_12562);
nand UO_1567 (O_1567,N_12035,N_14524);
nand UO_1568 (O_1568,N_13892,N_14499);
nor UO_1569 (O_1569,N_12173,N_14160);
and UO_1570 (O_1570,N_12723,N_13014);
or UO_1571 (O_1571,N_12970,N_14827);
and UO_1572 (O_1572,N_12106,N_14899);
nor UO_1573 (O_1573,N_12306,N_14759);
or UO_1574 (O_1574,N_12517,N_13502);
nand UO_1575 (O_1575,N_13609,N_13645);
and UO_1576 (O_1576,N_14467,N_13137);
nand UO_1577 (O_1577,N_12373,N_14294);
or UO_1578 (O_1578,N_13010,N_13244);
or UO_1579 (O_1579,N_12413,N_12758);
or UO_1580 (O_1580,N_12092,N_12026);
nand UO_1581 (O_1581,N_14322,N_14244);
nand UO_1582 (O_1582,N_14548,N_13678);
nor UO_1583 (O_1583,N_14869,N_13554);
and UO_1584 (O_1584,N_14673,N_12062);
or UO_1585 (O_1585,N_12259,N_13315);
or UO_1586 (O_1586,N_12092,N_14303);
nand UO_1587 (O_1587,N_13036,N_13587);
and UO_1588 (O_1588,N_14699,N_14492);
nand UO_1589 (O_1589,N_12902,N_14822);
or UO_1590 (O_1590,N_12066,N_12092);
or UO_1591 (O_1591,N_14703,N_13852);
and UO_1592 (O_1592,N_13782,N_14674);
and UO_1593 (O_1593,N_12913,N_13909);
xor UO_1594 (O_1594,N_14782,N_12166);
nor UO_1595 (O_1595,N_12460,N_12464);
nor UO_1596 (O_1596,N_13114,N_13672);
nand UO_1597 (O_1597,N_14873,N_13007);
and UO_1598 (O_1598,N_12099,N_14358);
nor UO_1599 (O_1599,N_12425,N_14717);
nand UO_1600 (O_1600,N_12070,N_12885);
nor UO_1601 (O_1601,N_12603,N_12674);
or UO_1602 (O_1602,N_13639,N_12427);
and UO_1603 (O_1603,N_13354,N_13666);
xor UO_1604 (O_1604,N_13468,N_14713);
or UO_1605 (O_1605,N_12375,N_13343);
nor UO_1606 (O_1606,N_13734,N_14086);
nor UO_1607 (O_1607,N_13188,N_13257);
and UO_1608 (O_1608,N_12310,N_13696);
nor UO_1609 (O_1609,N_14227,N_12555);
nand UO_1610 (O_1610,N_13644,N_14182);
nand UO_1611 (O_1611,N_13710,N_12466);
and UO_1612 (O_1612,N_14467,N_12168);
nand UO_1613 (O_1613,N_14179,N_12581);
nand UO_1614 (O_1614,N_13836,N_14247);
and UO_1615 (O_1615,N_14629,N_14128);
and UO_1616 (O_1616,N_12740,N_12421);
nor UO_1617 (O_1617,N_13340,N_13887);
and UO_1618 (O_1618,N_12807,N_12985);
nand UO_1619 (O_1619,N_12063,N_12168);
nor UO_1620 (O_1620,N_14335,N_13003);
or UO_1621 (O_1621,N_12650,N_14168);
and UO_1622 (O_1622,N_13882,N_14241);
or UO_1623 (O_1623,N_13851,N_14374);
nor UO_1624 (O_1624,N_14459,N_14863);
and UO_1625 (O_1625,N_14865,N_13500);
and UO_1626 (O_1626,N_14702,N_12965);
or UO_1627 (O_1627,N_14220,N_14129);
and UO_1628 (O_1628,N_13366,N_14947);
nor UO_1629 (O_1629,N_13437,N_13676);
nor UO_1630 (O_1630,N_13429,N_12927);
xnor UO_1631 (O_1631,N_12208,N_13417);
and UO_1632 (O_1632,N_14633,N_13966);
or UO_1633 (O_1633,N_14711,N_14018);
nor UO_1634 (O_1634,N_12546,N_12164);
or UO_1635 (O_1635,N_13681,N_13215);
and UO_1636 (O_1636,N_13634,N_13671);
nand UO_1637 (O_1637,N_13467,N_13458);
nand UO_1638 (O_1638,N_12089,N_12820);
nand UO_1639 (O_1639,N_13956,N_13726);
or UO_1640 (O_1640,N_13163,N_14537);
and UO_1641 (O_1641,N_14801,N_13487);
or UO_1642 (O_1642,N_12935,N_12677);
nand UO_1643 (O_1643,N_12009,N_12124);
or UO_1644 (O_1644,N_14698,N_14523);
or UO_1645 (O_1645,N_12817,N_13718);
nor UO_1646 (O_1646,N_14835,N_13728);
or UO_1647 (O_1647,N_13462,N_12715);
nor UO_1648 (O_1648,N_12386,N_13352);
xor UO_1649 (O_1649,N_13641,N_13814);
xnor UO_1650 (O_1650,N_12589,N_12040);
nor UO_1651 (O_1651,N_14384,N_12945);
and UO_1652 (O_1652,N_12120,N_12989);
and UO_1653 (O_1653,N_12839,N_14684);
nor UO_1654 (O_1654,N_13991,N_14436);
or UO_1655 (O_1655,N_14248,N_13722);
or UO_1656 (O_1656,N_12716,N_14379);
and UO_1657 (O_1657,N_14260,N_12396);
nand UO_1658 (O_1658,N_12643,N_12327);
or UO_1659 (O_1659,N_13591,N_12691);
nand UO_1660 (O_1660,N_14738,N_12058);
nor UO_1661 (O_1661,N_13665,N_12016);
xnor UO_1662 (O_1662,N_14798,N_14620);
or UO_1663 (O_1663,N_14273,N_14680);
xor UO_1664 (O_1664,N_13487,N_14919);
nand UO_1665 (O_1665,N_13827,N_14137);
and UO_1666 (O_1666,N_12468,N_13170);
xnor UO_1667 (O_1667,N_13060,N_12879);
or UO_1668 (O_1668,N_12977,N_14795);
and UO_1669 (O_1669,N_12295,N_12734);
nor UO_1670 (O_1670,N_13722,N_13803);
xor UO_1671 (O_1671,N_12435,N_14168);
and UO_1672 (O_1672,N_13446,N_12722);
nand UO_1673 (O_1673,N_12985,N_14928);
or UO_1674 (O_1674,N_12194,N_13890);
or UO_1675 (O_1675,N_13442,N_14709);
xor UO_1676 (O_1676,N_12828,N_13201);
or UO_1677 (O_1677,N_12524,N_14093);
nand UO_1678 (O_1678,N_12638,N_12756);
nand UO_1679 (O_1679,N_13256,N_13212);
or UO_1680 (O_1680,N_14592,N_12878);
and UO_1681 (O_1681,N_12530,N_12222);
and UO_1682 (O_1682,N_14870,N_12197);
or UO_1683 (O_1683,N_14667,N_12199);
nand UO_1684 (O_1684,N_12810,N_12718);
nor UO_1685 (O_1685,N_14149,N_14398);
nor UO_1686 (O_1686,N_12962,N_14633);
or UO_1687 (O_1687,N_14535,N_14168);
nand UO_1688 (O_1688,N_14931,N_12131);
and UO_1689 (O_1689,N_13107,N_13457);
and UO_1690 (O_1690,N_14607,N_14770);
nor UO_1691 (O_1691,N_14834,N_12055);
or UO_1692 (O_1692,N_12305,N_12714);
or UO_1693 (O_1693,N_13049,N_14551);
nand UO_1694 (O_1694,N_14766,N_14316);
nor UO_1695 (O_1695,N_14934,N_14406);
nand UO_1696 (O_1696,N_12569,N_12605);
nor UO_1697 (O_1697,N_12567,N_13913);
nor UO_1698 (O_1698,N_14745,N_14330);
nand UO_1699 (O_1699,N_12056,N_14283);
or UO_1700 (O_1700,N_12447,N_14843);
and UO_1701 (O_1701,N_14391,N_12122);
nand UO_1702 (O_1702,N_14991,N_12147);
nor UO_1703 (O_1703,N_14077,N_12251);
nor UO_1704 (O_1704,N_12969,N_14889);
nor UO_1705 (O_1705,N_12355,N_14471);
nor UO_1706 (O_1706,N_13496,N_14536);
xor UO_1707 (O_1707,N_14980,N_14470);
nand UO_1708 (O_1708,N_13008,N_14194);
and UO_1709 (O_1709,N_13492,N_14458);
nand UO_1710 (O_1710,N_14960,N_14177);
and UO_1711 (O_1711,N_14416,N_12287);
or UO_1712 (O_1712,N_13953,N_13910);
and UO_1713 (O_1713,N_12659,N_12385);
xor UO_1714 (O_1714,N_14955,N_13634);
and UO_1715 (O_1715,N_13052,N_14114);
nor UO_1716 (O_1716,N_12131,N_12013);
and UO_1717 (O_1717,N_12742,N_13700);
and UO_1718 (O_1718,N_13284,N_13177);
nor UO_1719 (O_1719,N_12521,N_13088);
and UO_1720 (O_1720,N_14680,N_12561);
nor UO_1721 (O_1721,N_13128,N_13484);
nor UO_1722 (O_1722,N_14178,N_13764);
nor UO_1723 (O_1723,N_14464,N_13366);
nand UO_1724 (O_1724,N_14729,N_12445);
and UO_1725 (O_1725,N_12281,N_12366);
or UO_1726 (O_1726,N_14823,N_14227);
and UO_1727 (O_1727,N_12814,N_12021);
nor UO_1728 (O_1728,N_12921,N_13958);
nand UO_1729 (O_1729,N_14993,N_14002);
or UO_1730 (O_1730,N_12064,N_13438);
or UO_1731 (O_1731,N_12819,N_12995);
and UO_1732 (O_1732,N_14462,N_14076);
or UO_1733 (O_1733,N_14146,N_14852);
nand UO_1734 (O_1734,N_12752,N_13924);
or UO_1735 (O_1735,N_14408,N_12097);
and UO_1736 (O_1736,N_12297,N_12686);
nor UO_1737 (O_1737,N_13380,N_14440);
nor UO_1738 (O_1738,N_14175,N_13365);
nand UO_1739 (O_1739,N_13982,N_13751);
or UO_1740 (O_1740,N_12782,N_13034);
and UO_1741 (O_1741,N_13027,N_12169);
nor UO_1742 (O_1742,N_14700,N_14024);
nor UO_1743 (O_1743,N_12876,N_14868);
and UO_1744 (O_1744,N_12123,N_13335);
nor UO_1745 (O_1745,N_14210,N_12783);
and UO_1746 (O_1746,N_14204,N_14640);
nor UO_1747 (O_1747,N_14364,N_14361);
xor UO_1748 (O_1748,N_13621,N_14802);
and UO_1749 (O_1749,N_12726,N_12825);
xor UO_1750 (O_1750,N_13628,N_12707);
and UO_1751 (O_1751,N_13533,N_13212);
and UO_1752 (O_1752,N_13822,N_13328);
nor UO_1753 (O_1753,N_12066,N_14061);
xor UO_1754 (O_1754,N_14944,N_13782);
or UO_1755 (O_1755,N_13798,N_14730);
nor UO_1756 (O_1756,N_12153,N_14555);
nand UO_1757 (O_1757,N_14815,N_13992);
or UO_1758 (O_1758,N_14048,N_14381);
or UO_1759 (O_1759,N_13483,N_14257);
nor UO_1760 (O_1760,N_14843,N_14278);
and UO_1761 (O_1761,N_13217,N_14697);
nor UO_1762 (O_1762,N_14275,N_13783);
and UO_1763 (O_1763,N_13521,N_14175);
nor UO_1764 (O_1764,N_14976,N_12583);
and UO_1765 (O_1765,N_13342,N_14393);
or UO_1766 (O_1766,N_12151,N_12004);
nor UO_1767 (O_1767,N_13888,N_12025);
or UO_1768 (O_1768,N_12466,N_13732);
and UO_1769 (O_1769,N_14654,N_12595);
or UO_1770 (O_1770,N_14746,N_14875);
nand UO_1771 (O_1771,N_12242,N_14212);
and UO_1772 (O_1772,N_14319,N_13543);
nor UO_1773 (O_1773,N_13575,N_13202);
and UO_1774 (O_1774,N_12775,N_12734);
and UO_1775 (O_1775,N_13547,N_13212);
and UO_1776 (O_1776,N_12127,N_14425);
and UO_1777 (O_1777,N_12942,N_13290);
and UO_1778 (O_1778,N_13345,N_14518);
nand UO_1779 (O_1779,N_14200,N_14996);
and UO_1780 (O_1780,N_12559,N_13531);
or UO_1781 (O_1781,N_13041,N_13363);
or UO_1782 (O_1782,N_13459,N_12033);
and UO_1783 (O_1783,N_13980,N_13262);
nor UO_1784 (O_1784,N_13510,N_14567);
or UO_1785 (O_1785,N_13354,N_14354);
and UO_1786 (O_1786,N_14447,N_14290);
and UO_1787 (O_1787,N_13834,N_14181);
nand UO_1788 (O_1788,N_14101,N_14823);
nor UO_1789 (O_1789,N_13898,N_14413);
nand UO_1790 (O_1790,N_13767,N_12935);
nor UO_1791 (O_1791,N_14018,N_12576);
nand UO_1792 (O_1792,N_13595,N_14499);
nand UO_1793 (O_1793,N_12277,N_12203);
nand UO_1794 (O_1794,N_14438,N_12558);
nand UO_1795 (O_1795,N_14570,N_12905);
and UO_1796 (O_1796,N_13639,N_13256);
nor UO_1797 (O_1797,N_12443,N_13688);
and UO_1798 (O_1798,N_14854,N_13133);
and UO_1799 (O_1799,N_14123,N_12694);
or UO_1800 (O_1800,N_13990,N_12355);
xnor UO_1801 (O_1801,N_14461,N_14167);
or UO_1802 (O_1802,N_12210,N_13735);
xnor UO_1803 (O_1803,N_14310,N_13502);
xnor UO_1804 (O_1804,N_13370,N_13628);
or UO_1805 (O_1805,N_14642,N_14471);
nor UO_1806 (O_1806,N_12628,N_14530);
and UO_1807 (O_1807,N_12914,N_14459);
or UO_1808 (O_1808,N_13443,N_13578);
and UO_1809 (O_1809,N_13803,N_14552);
nor UO_1810 (O_1810,N_12744,N_14533);
or UO_1811 (O_1811,N_12359,N_14446);
nor UO_1812 (O_1812,N_14883,N_13258);
or UO_1813 (O_1813,N_12440,N_13703);
or UO_1814 (O_1814,N_13660,N_13212);
and UO_1815 (O_1815,N_12626,N_12773);
and UO_1816 (O_1816,N_13370,N_13096);
nor UO_1817 (O_1817,N_13517,N_14127);
nor UO_1818 (O_1818,N_14582,N_12805);
nand UO_1819 (O_1819,N_12321,N_13730);
nor UO_1820 (O_1820,N_14043,N_12505);
nand UO_1821 (O_1821,N_12628,N_13486);
and UO_1822 (O_1822,N_14996,N_13957);
or UO_1823 (O_1823,N_12775,N_13042);
xor UO_1824 (O_1824,N_14299,N_13994);
nand UO_1825 (O_1825,N_13453,N_14838);
nand UO_1826 (O_1826,N_12168,N_14545);
nor UO_1827 (O_1827,N_13652,N_12045);
or UO_1828 (O_1828,N_12618,N_14433);
xnor UO_1829 (O_1829,N_12020,N_12164);
and UO_1830 (O_1830,N_12861,N_14038);
nor UO_1831 (O_1831,N_13932,N_14382);
nand UO_1832 (O_1832,N_13499,N_13913);
nand UO_1833 (O_1833,N_14515,N_12923);
or UO_1834 (O_1834,N_12643,N_14491);
nand UO_1835 (O_1835,N_12276,N_13986);
and UO_1836 (O_1836,N_12766,N_12911);
and UO_1837 (O_1837,N_13052,N_12680);
and UO_1838 (O_1838,N_14712,N_14030);
nand UO_1839 (O_1839,N_13600,N_12023);
and UO_1840 (O_1840,N_12025,N_12383);
and UO_1841 (O_1841,N_14505,N_14724);
or UO_1842 (O_1842,N_13653,N_14715);
or UO_1843 (O_1843,N_13900,N_14165);
or UO_1844 (O_1844,N_14441,N_14620);
or UO_1845 (O_1845,N_12339,N_13052);
xor UO_1846 (O_1846,N_14427,N_14551);
nand UO_1847 (O_1847,N_14655,N_13206);
nand UO_1848 (O_1848,N_13773,N_12749);
nor UO_1849 (O_1849,N_14974,N_14891);
or UO_1850 (O_1850,N_12299,N_13294);
xor UO_1851 (O_1851,N_14754,N_14139);
and UO_1852 (O_1852,N_14598,N_13021);
nor UO_1853 (O_1853,N_14298,N_12422);
nor UO_1854 (O_1854,N_12139,N_12788);
nand UO_1855 (O_1855,N_12968,N_13322);
nor UO_1856 (O_1856,N_13610,N_13340);
nand UO_1857 (O_1857,N_12765,N_14721);
or UO_1858 (O_1858,N_12779,N_13934);
xor UO_1859 (O_1859,N_13986,N_12538);
nand UO_1860 (O_1860,N_12506,N_14368);
nand UO_1861 (O_1861,N_13409,N_12649);
and UO_1862 (O_1862,N_14046,N_12431);
or UO_1863 (O_1863,N_12986,N_13618);
nor UO_1864 (O_1864,N_12636,N_12612);
nand UO_1865 (O_1865,N_13680,N_13490);
or UO_1866 (O_1866,N_12824,N_13502);
nand UO_1867 (O_1867,N_13320,N_13661);
and UO_1868 (O_1868,N_12155,N_14387);
nand UO_1869 (O_1869,N_12889,N_13394);
or UO_1870 (O_1870,N_12203,N_13281);
xnor UO_1871 (O_1871,N_13901,N_13013);
and UO_1872 (O_1872,N_12390,N_12886);
and UO_1873 (O_1873,N_13484,N_12119);
or UO_1874 (O_1874,N_14938,N_12046);
nor UO_1875 (O_1875,N_14450,N_14211);
nor UO_1876 (O_1876,N_12825,N_14126);
nand UO_1877 (O_1877,N_13251,N_14189);
nor UO_1878 (O_1878,N_14174,N_12841);
and UO_1879 (O_1879,N_13499,N_12401);
or UO_1880 (O_1880,N_14542,N_14973);
nand UO_1881 (O_1881,N_14875,N_12329);
and UO_1882 (O_1882,N_14336,N_14647);
nand UO_1883 (O_1883,N_14508,N_13499);
or UO_1884 (O_1884,N_13012,N_13675);
and UO_1885 (O_1885,N_12338,N_12348);
and UO_1886 (O_1886,N_13544,N_13669);
and UO_1887 (O_1887,N_13844,N_14582);
nand UO_1888 (O_1888,N_14699,N_12724);
and UO_1889 (O_1889,N_13819,N_13505);
nand UO_1890 (O_1890,N_14154,N_13800);
nor UO_1891 (O_1891,N_12955,N_14073);
and UO_1892 (O_1892,N_13108,N_12786);
and UO_1893 (O_1893,N_14416,N_14418);
and UO_1894 (O_1894,N_13660,N_13881);
or UO_1895 (O_1895,N_12851,N_13787);
and UO_1896 (O_1896,N_12815,N_12559);
or UO_1897 (O_1897,N_14050,N_14550);
nand UO_1898 (O_1898,N_14745,N_13254);
nand UO_1899 (O_1899,N_13890,N_12107);
and UO_1900 (O_1900,N_12505,N_13223);
nand UO_1901 (O_1901,N_14760,N_12961);
and UO_1902 (O_1902,N_13202,N_14097);
and UO_1903 (O_1903,N_12611,N_13304);
nor UO_1904 (O_1904,N_14168,N_14772);
or UO_1905 (O_1905,N_14503,N_12654);
nand UO_1906 (O_1906,N_12494,N_13131);
nand UO_1907 (O_1907,N_12894,N_13803);
or UO_1908 (O_1908,N_12004,N_14466);
and UO_1909 (O_1909,N_14954,N_14552);
nand UO_1910 (O_1910,N_12051,N_13590);
or UO_1911 (O_1911,N_12858,N_13449);
or UO_1912 (O_1912,N_13974,N_12907);
nor UO_1913 (O_1913,N_12634,N_13423);
and UO_1914 (O_1914,N_12612,N_13614);
and UO_1915 (O_1915,N_14312,N_14428);
xnor UO_1916 (O_1916,N_13045,N_13551);
nor UO_1917 (O_1917,N_13750,N_14177);
xnor UO_1918 (O_1918,N_13886,N_13557);
nand UO_1919 (O_1919,N_14322,N_12016);
xnor UO_1920 (O_1920,N_13495,N_13020);
nor UO_1921 (O_1921,N_13237,N_13358);
xor UO_1922 (O_1922,N_13670,N_13795);
nand UO_1923 (O_1923,N_14275,N_13533);
nor UO_1924 (O_1924,N_13052,N_14962);
nand UO_1925 (O_1925,N_13803,N_14134);
xor UO_1926 (O_1926,N_12552,N_12162);
nor UO_1927 (O_1927,N_12141,N_13763);
or UO_1928 (O_1928,N_14354,N_14360);
nand UO_1929 (O_1929,N_14857,N_13903);
xor UO_1930 (O_1930,N_14221,N_14763);
or UO_1931 (O_1931,N_13875,N_13475);
or UO_1932 (O_1932,N_13029,N_14775);
or UO_1933 (O_1933,N_13835,N_13642);
xnor UO_1934 (O_1934,N_12181,N_13421);
nor UO_1935 (O_1935,N_12929,N_13680);
and UO_1936 (O_1936,N_14100,N_14142);
and UO_1937 (O_1937,N_13778,N_13534);
and UO_1938 (O_1938,N_12936,N_13493);
or UO_1939 (O_1939,N_14167,N_12150);
and UO_1940 (O_1940,N_13543,N_13266);
or UO_1941 (O_1941,N_13666,N_14480);
nor UO_1942 (O_1942,N_12928,N_14857);
nor UO_1943 (O_1943,N_12298,N_12153);
nand UO_1944 (O_1944,N_14829,N_14210);
nor UO_1945 (O_1945,N_13435,N_13854);
nor UO_1946 (O_1946,N_12163,N_14615);
xnor UO_1947 (O_1947,N_12515,N_13365);
nand UO_1948 (O_1948,N_13789,N_13769);
nand UO_1949 (O_1949,N_14270,N_13590);
and UO_1950 (O_1950,N_14710,N_12236);
or UO_1951 (O_1951,N_12052,N_12000);
nand UO_1952 (O_1952,N_13322,N_13867);
nor UO_1953 (O_1953,N_13842,N_13496);
or UO_1954 (O_1954,N_14641,N_13174);
nor UO_1955 (O_1955,N_12760,N_14944);
or UO_1956 (O_1956,N_13570,N_14248);
or UO_1957 (O_1957,N_13998,N_14179);
nand UO_1958 (O_1958,N_14267,N_14181);
or UO_1959 (O_1959,N_14067,N_13182);
nor UO_1960 (O_1960,N_13818,N_13793);
and UO_1961 (O_1961,N_14446,N_12639);
nand UO_1962 (O_1962,N_14818,N_12669);
xor UO_1963 (O_1963,N_13019,N_14620);
xor UO_1964 (O_1964,N_14013,N_12407);
or UO_1965 (O_1965,N_12394,N_13813);
nand UO_1966 (O_1966,N_12340,N_12756);
or UO_1967 (O_1967,N_12809,N_13072);
nor UO_1968 (O_1968,N_14464,N_12539);
xor UO_1969 (O_1969,N_12658,N_12176);
nand UO_1970 (O_1970,N_13400,N_14641);
or UO_1971 (O_1971,N_14710,N_12313);
nand UO_1972 (O_1972,N_13598,N_12379);
nor UO_1973 (O_1973,N_13113,N_14830);
and UO_1974 (O_1974,N_13705,N_13696);
nor UO_1975 (O_1975,N_12439,N_12463);
xor UO_1976 (O_1976,N_14798,N_13367);
nand UO_1977 (O_1977,N_12664,N_14879);
nor UO_1978 (O_1978,N_14345,N_13857);
and UO_1979 (O_1979,N_12063,N_14227);
xor UO_1980 (O_1980,N_12550,N_13095);
nand UO_1981 (O_1981,N_12511,N_13700);
nor UO_1982 (O_1982,N_14348,N_12175);
or UO_1983 (O_1983,N_12914,N_12959);
nor UO_1984 (O_1984,N_13303,N_12357);
and UO_1985 (O_1985,N_13788,N_12693);
or UO_1986 (O_1986,N_13252,N_12499);
or UO_1987 (O_1987,N_14757,N_13539);
nor UO_1988 (O_1988,N_14419,N_12171);
nand UO_1989 (O_1989,N_12412,N_14467);
xnor UO_1990 (O_1990,N_12678,N_13149);
or UO_1991 (O_1991,N_12628,N_13235);
or UO_1992 (O_1992,N_14071,N_13719);
nor UO_1993 (O_1993,N_12373,N_13696);
xnor UO_1994 (O_1994,N_12368,N_13274);
and UO_1995 (O_1995,N_14212,N_14235);
and UO_1996 (O_1996,N_12547,N_12157);
nor UO_1997 (O_1997,N_14285,N_13817);
nor UO_1998 (O_1998,N_12738,N_12801);
or UO_1999 (O_1999,N_13103,N_14988);
endmodule