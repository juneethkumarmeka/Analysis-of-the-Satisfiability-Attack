module basic_750_5000_1000_5_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_18,In_618);
nand U1 (N_1,In_442,In_651);
and U2 (N_2,In_690,In_472);
or U3 (N_3,In_231,In_272);
and U4 (N_4,In_702,In_417);
nand U5 (N_5,In_587,In_218);
nand U6 (N_6,In_739,In_674);
or U7 (N_7,In_515,In_467);
or U8 (N_8,In_224,In_216);
or U9 (N_9,In_341,In_443);
nand U10 (N_10,In_3,In_196);
or U11 (N_11,In_697,In_323);
nand U12 (N_12,In_726,In_320);
or U13 (N_13,In_409,In_38);
and U14 (N_14,In_124,In_448);
and U15 (N_15,In_423,In_584);
or U16 (N_16,In_355,In_680);
and U17 (N_17,In_556,In_292);
nor U18 (N_18,In_92,In_172);
nand U19 (N_19,In_376,In_159);
nor U20 (N_20,In_247,In_549);
or U21 (N_21,In_644,In_568);
or U22 (N_22,In_570,In_386);
nor U23 (N_23,In_678,In_508);
xor U24 (N_24,In_712,In_6);
or U25 (N_25,In_184,In_45);
or U26 (N_26,In_478,In_366);
or U27 (N_27,In_668,In_527);
or U28 (N_28,In_368,In_748);
nor U29 (N_29,In_483,In_40);
nand U30 (N_30,In_377,In_462);
and U31 (N_31,In_270,In_707);
nor U32 (N_32,In_44,In_378);
or U33 (N_33,In_264,In_497);
or U34 (N_34,In_717,In_153);
nor U35 (N_35,In_275,In_276);
or U36 (N_36,In_689,In_609);
and U37 (N_37,In_435,In_491);
or U38 (N_38,In_607,In_724);
nand U39 (N_39,In_234,In_273);
nor U40 (N_40,In_107,In_173);
and U41 (N_41,In_164,In_634);
or U42 (N_42,In_715,In_295);
nor U43 (N_43,In_594,In_572);
nor U44 (N_44,In_490,In_670);
xnor U45 (N_45,In_104,In_242);
nand U46 (N_46,In_83,In_130);
nor U47 (N_47,In_461,In_676);
nor U48 (N_48,In_420,In_387);
and U49 (N_49,In_743,In_639);
and U50 (N_50,In_625,In_460);
nand U51 (N_51,In_672,In_400);
and U52 (N_52,In_551,In_226);
or U53 (N_53,In_21,In_220);
or U54 (N_54,In_694,In_727);
or U55 (N_55,In_330,In_326);
nor U56 (N_56,In_26,In_359);
nor U57 (N_57,In_468,In_314);
or U58 (N_58,In_471,In_313);
or U59 (N_59,In_201,In_561);
nand U60 (N_60,In_682,In_582);
nand U61 (N_61,In_64,In_266);
nor U62 (N_62,In_654,In_42);
nand U63 (N_63,In_48,In_39);
nand U64 (N_64,In_532,In_170);
nand U65 (N_65,In_202,In_66);
and U66 (N_66,In_631,In_97);
and U67 (N_67,In_494,In_134);
and U68 (N_68,In_565,In_392);
or U69 (N_69,In_8,In_28);
nor U70 (N_70,In_362,In_518);
nand U71 (N_71,In_206,In_681);
nor U72 (N_72,In_113,In_641);
nor U73 (N_73,In_536,In_627);
and U74 (N_74,In_289,In_391);
and U75 (N_75,In_127,In_431);
nor U76 (N_76,In_58,In_426);
nor U77 (N_77,In_211,In_236);
and U78 (N_78,In_685,In_575);
nand U79 (N_79,In_734,In_333);
or U80 (N_80,In_517,In_335);
xor U81 (N_81,In_354,In_297);
and U82 (N_82,In_439,In_597);
nand U83 (N_83,In_611,In_353);
and U84 (N_84,In_412,In_165);
and U85 (N_85,In_719,In_5);
nor U86 (N_86,In_732,In_598);
nand U87 (N_87,In_339,In_123);
nand U88 (N_88,In_336,In_505);
nand U89 (N_89,In_31,In_208);
nand U90 (N_90,In_194,In_160);
or U91 (N_91,In_480,In_51);
or U92 (N_92,In_293,In_129);
and U93 (N_93,In_604,In_139);
xor U94 (N_94,In_344,In_161);
nor U95 (N_95,In_630,In_301);
nand U96 (N_96,In_658,In_262);
or U97 (N_97,In_521,In_503);
or U98 (N_98,In_195,In_285);
or U99 (N_99,In_253,In_605);
nor U100 (N_100,In_119,In_4);
nand U101 (N_101,In_327,In_351);
nand U102 (N_102,In_610,In_349);
or U103 (N_103,In_70,In_1);
nor U104 (N_104,In_176,In_288);
and U105 (N_105,In_553,In_512);
nor U106 (N_106,In_80,In_539);
and U107 (N_107,In_402,In_519);
xnor U108 (N_108,In_413,In_722);
nand U109 (N_109,In_464,In_151);
nor U110 (N_110,In_398,In_615);
nand U111 (N_111,In_374,In_736);
nand U112 (N_112,In_576,In_32);
or U113 (N_113,In_267,In_514);
or U114 (N_114,In_542,In_408);
nand U115 (N_115,In_259,In_25);
and U116 (N_116,In_621,In_473);
nand U117 (N_117,In_571,In_269);
xnor U118 (N_118,In_217,In_188);
xnor U119 (N_119,In_233,In_701);
or U120 (N_120,In_158,In_533);
or U121 (N_121,In_662,In_200);
nor U122 (N_122,In_683,In_733);
nand U123 (N_123,In_283,In_248);
or U124 (N_124,In_452,In_171);
or U125 (N_125,In_9,In_197);
nor U126 (N_126,In_177,In_738);
nor U127 (N_127,In_401,In_495);
or U128 (N_128,In_13,In_309);
or U129 (N_129,In_65,In_746);
or U130 (N_130,In_310,In_530);
or U131 (N_131,In_69,In_73);
nand U132 (N_132,In_181,In_227);
or U133 (N_133,In_50,In_82);
or U134 (N_134,In_579,In_692);
or U135 (N_135,In_96,In_688);
and U136 (N_136,In_718,In_235);
or U137 (N_137,In_440,In_745);
and U138 (N_138,In_659,In_588);
and U139 (N_139,In_63,In_255);
or U140 (N_140,In_241,In_559);
and U141 (N_141,In_524,In_528);
and U142 (N_142,In_302,In_535);
or U143 (N_143,In_457,In_406);
nand U144 (N_144,In_221,In_147);
nor U145 (N_145,In_15,In_585);
or U146 (N_146,In_245,In_135);
nand U147 (N_147,In_703,In_257);
nor U148 (N_148,In_741,In_470);
and U149 (N_149,In_237,In_175);
and U150 (N_150,In_540,In_223);
nand U151 (N_151,In_671,In_543);
nand U152 (N_152,In_370,In_493);
or U153 (N_153,In_602,In_300);
nor U154 (N_154,In_414,In_531);
nor U155 (N_155,In_101,In_586);
or U156 (N_156,In_338,In_581);
nand U157 (N_157,In_404,In_268);
nor U158 (N_158,In_74,In_463);
xnor U159 (N_159,In_99,In_282);
nand U160 (N_160,In_729,In_81);
or U161 (N_161,In_477,In_251);
nand U162 (N_162,In_312,In_510);
nand U163 (N_163,In_466,In_422);
or U164 (N_164,In_663,In_459);
and U165 (N_165,In_169,In_204);
and U166 (N_166,In_429,In_122);
nand U167 (N_167,In_589,In_385);
or U168 (N_168,In_279,In_669);
or U169 (N_169,In_277,In_705);
or U170 (N_170,In_254,In_30);
and U171 (N_171,In_361,In_198);
and U172 (N_172,In_507,In_437);
nor U173 (N_173,In_150,In_140);
nand U174 (N_174,In_436,In_620);
and U175 (N_175,In_128,In_428);
or U176 (N_176,In_445,In_555);
and U177 (N_177,In_501,In_450);
or U178 (N_178,In_447,In_560);
nand U179 (N_179,In_695,In_619);
or U180 (N_180,In_421,In_290);
and U181 (N_181,In_444,In_324);
or U182 (N_182,In_382,In_192);
or U183 (N_183,In_121,In_388);
or U184 (N_184,In_486,In_375);
or U185 (N_185,In_731,In_603);
or U186 (N_186,In_263,In_182);
or U187 (N_187,In_210,In_416);
and U188 (N_188,In_496,In_108);
nand U189 (N_189,In_427,In_744);
nor U190 (N_190,In_43,In_72);
nor U191 (N_191,In_281,In_29);
or U192 (N_192,In_433,In_156);
and U193 (N_193,In_93,In_133);
nor U194 (N_194,In_479,In_166);
or U195 (N_195,In_713,In_145);
and U196 (N_196,In_612,In_229);
and U197 (N_197,In_306,In_296);
and U198 (N_198,In_723,In_642);
nor U199 (N_199,In_638,In_183);
and U200 (N_200,In_95,In_365);
nor U201 (N_201,In_381,In_213);
and U202 (N_202,In_469,In_499);
or U203 (N_203,In_316,In_57);
nand U204 (N_204,In_89,In_189);
nor U205 (N_205,In_53,In_547);
nor U206 (N_206,In_23,In_574);
and U207 (N_207,In_686,In_661);
or U208 (N_208,In_67,In_343);
nor U209 (N_209,In_606,In_68);
or U210 (N_210,In_474,In_632);
nor U211 (N_211,In_525,In_673);
or U212 (N_212,In_60,In_308);
nand U213 (N_213,In_737,In_541);
nand U214 (N_214,In_645,In_284);
or U215 (N_215,In_481,In_360);
and U216 (N_216,In_432,In_256);
and U217 (N_217,In_307,In_199);
or U218 (N_218,In_449,In_71);
nor U219 (N_219,In_46,In_347);
nor U220 (N_220,In_520,In_476);
or U221 (N_221,In_185,In_329);
and U222 (N_222,In_334,In_693);
and U223 (N_223,In_389,In_465);
or U224 (N_224,In_337,In_600);
or U225 (N_225,In_367,In_35);
nor U226 (N_226,In_305,In_578);
nor U227 (N_227,In_10,In_131);
or U228 (N_228,In_274,In_657);
and U229 (N_229,In_434,In_643);
nor U230 (N_230,In_0,In_438);
and U231 (N_231,In_14,In_22);
nor U232 (N_232,In_315,In_411);
or U233 (N_233,In_506,In_407);
or U234 (N_234,In_114,In_526);
nor U235 (N_235,In_577,In_637);
nor U236 (N_236,In_191,In_394);
nor U237 (N_237,In_656,In_509);
nor U238 (N_238,In_149,In_118);
and U239 (N_239,In_714,In_655);
nand U240 (N_240,In_280,In_34);
and U241 (N_241,In_348,In_174);
nor U242 (N_242,In_544,In_54);
and U243 (N_243,In_552,In_91);
nor U244 (N_244,In_325,In_397);
and U245 (N_245,In_356,In_61);
and U246 (N_246,In_358,In_554);
nand U247 (N_247,In_390,In_487);
nand U248 (N_248,In_332,In_679);
or U249 (N_249,In_212,In_137);
nand U250 (N_250,In_340,In_109);
xor U251 (N_251,In_345,In_700);
nand U252 (N_252,In_614,In_425);
nor U253 (N_253,In_529,In_163);
nand U254 (N_254,In_331,In_317);
or U255 (N_255,In_371,In_522);
and U256 (N_256,In_155,In_225);
nor U257 (N_257,In_157,In_500);
and U258 (N_258,In_239,In_110);
nand U259 (N_259,In_168,In_143);
and U260 (N_260,In_492,In_484);
nand U261 (N_261,In_567,In_278);
nand U262 (N_262,In_311,In_249);
or U263 (N_263,In_418,In_37);
and U264 (N_264,In_294,In_410);
and U265 (N_265,In_593,In_105);
or U266 (N_266,In_62,In_260);
nand U267 (N_267,In_318,In_115);
and U268 (N_268,In_246,In_190);
nand U269 (N_269,In_677,In_77);
nor U270 (N_270,In_564,In_395);
nand U271 (N_271,In_342,In_291);
nor U272 (N_272,In_142,In_304);
or U273 (N_273,In_728,In_652);
nand U274 (N_274,In_569,In_106);
nor U275 (N_275,In_187,In_384);
nand U276 (N_276,In_55,In_243);
nor U277 (N_277,In_94,In_238);
nand U278 (N_278,In_740,In_120);
and U279 (N_279,In_271,In_403);
nand U280 (N_280,In_592,In_558);
nand U281 (N_281,In_747,In_380);
or U282 (N_282,In_502,In_87);
or U283 (N_283,In_511,In_125);
and U284 (N_284,In_446,In_222);
or U285 (N_285,In_322,In_148);
or U286 (N_286,In_504,In_207);
nand U287 (N_287,In_430,In_710);
nor U288 (N_288,In_100,In_516);
and U289 (N_289,In_696,In_11);
nor U290 (N_290,In_141,In_383);
nand U291 (N_291,In_583,In_219);
nand U292 (N_292,In_49,In_52);
nand U293 (N_293,In_636,In_405);
nand U294 (N_294,In_179,In_666);
nand U295 (N_295,In_595,In_116);
or U296 (N_296,In_513,In_144);
and U297 (N_297,In_261,In_563);
nand U298 (N_298,In_441,In_84);
or U299 (N_299,In_616,In_653);
nor U300 (N_300,In_419,In_706);
nor U301 (N_301,In_485,In_244);
nand U302 (N_302,In_482,In_613);
nor U303 (N_303,In_458,In_649);
nand U304 (N_304,In_633,In_725);
and U305 (N_305,In_19,In_186);
nor U306 (N_306,In_146,In_178);
nor U307 (N_307,In_545,In_373);
or U308 (N_308,In_215,In_537);
nor U309 (N_309,In_675,In_629);
or U310 (N_310,In_455,In_36);
and U311 (N_311,In_691,In_103);
or U312 (N_312,In_117,In_2);
and U313 (N_313,In_328,In_20);
nor U314 (N_314,In_232,In_475);
and U315 (N_315,In_372,In_321);
nor U316 (N_316,In_730,In_580);
nand U317 (N_317,In_180,In_566);
or U318 (N_318,In_287,In_489);
and U319 (N_319,In_228,In_646);
nor U320 (N_320,In_667,In_709);
nand U321 (N_321,In_350,In_687);
and U322 (N_322,In_59,In_534);
or U323 (N_323,In_154,In_17);
or U324 (N_324,In_699,In_88);
or U325 (N_325,In_623,In_399);
nand U326 (N_326,In_162,In_152);
and U327 (N_327,In_665,In_599);
and U328 (N_328,In_635,In_363);
nor U329 (N_329,In_742,In_205);
nand U330 (N_330,In_265,In_711);
and U331 (N_331,In_193,In_573);
nor U332 (N_332,In_456,In_102);
and U333 (N_333,In_240,In_650);
or U334 (N_334,In_749,In_548);
or U335 (N_335,In_590,In_454);
nor U336 (N_336,In_258,In_85);
nand U337 (N_337,In_498,In_346);
and U338 (N_338,In_252,In_47);
nand U339 (N_339,In_298,In_488);
nor U340 (N_340,In_628,In_601);
nor U341 (N_341,In_319,In_209);
nand U342 (N_342,In_698,In_640);
or U343 (N_343,In_214,In_112);
nand U344 (N_344,In_352,In_286);
nor U345 (N_345,In_720,In_617);
nor U346 (N_346,In_12,In_704);
nor U347 (N_347,In_86,In_299);
and U348 (N_348,In_557,In_79);
nor U349 (N_349,In_203,In_369);
and U350 (N_350,In_75,In_24);
nand U351 (N_351,In_415,In_27);
nand U352 (N_352,In_379,In_664);
nand U353 (N_353,In_396,In_364);
and U354 (N_354,In_684,In_250);
and U355 (N_355,In_41,In_56);
nor U356 (N_356,In_132,In_562);
nor U357 (N_357,In_167,In_453);
and U358 (N_358,In_7,In_546);
nor U359 (N_359,In_357,In_647);
and U360 (N_360,In_424,In_660);
and U361 (N_361,In_735,In_538);
nand U362 (N_362,In_98,In_622);
and U363 (N_363,In_303,In_138);
or U364 (N_364,In_90,In_648);
nand U365 (N_365,In_626,In_78);
and U366 (N_366,In_608,In_716);
nand U367 (N_367,In_624,In_721);
or U368 (N_368,In_126,In_708);
nand U369 (N_369,In_76,In_591);
nand U370 (N_370,In_451,In_33);
nor U371 (N_371,In_136,In_550);
nand U372 (N_372,In_596,In_16);
or U373 (N_373,In_230,In_523);
nand U374 (N_374,In_393,In_111);
nor U375 (N_375,In_249,In_73);
or U376 (N_376,In_77,In_729);
and U377 (N_377,In_39,In_148);
nor U378 (N_378,In_683,In_625);
nand U379 (N_379,In_475,In_317);
and U380 (N_380,In_429,In_291);
nor U381 (N_381,In_294,In_273);
nor U382 (N_382,In_314,In_666);
or U383 (N_383,In_629,In_516);
nor U384 (N_384,In_589,In_42);
nor U385 (N_385,In_703,In_174);
or U386 (N_386,In_659,In_676);
nor U387 (N_387,In_260,In_313);
or U388 (N_388,In_148,In_414);
and U389 (N_389,In_220,In_341);
or U390 (N_390,In_389,In_372);
or U391 (N_391,In_0,In_641);
or U392 (N_392,In_137,In_4);
or U393 (N_393,In_465,In_476);
and U394 (N_394,In_705,In_289);
nor U395 (N_395,In_589,In_239);
nand U396 (N_396,In_513,In_649);
nor U397 (N_397,In_529,In_313);
and U398 (N_398,In_86,In_225);
and U399 (N_399,In_579,In_436);
nand U400 (N_400,In_704,In_332);
nor U401 (N_401,In_427,In_615);
and U402 (N_402,In_35,In_159);
nand U403 (N_403,In_288,In_686);
nand U404 (N_404,In_698,In_166);
and U405 (N_405,In_453,In_625);
or U406 (N_406,In_372,In_65);
nor U407 (N_407,In_435,In_632);
or U408 (N_408,In_91,In_583);
and U409 (N_409,In_59,In_697);
nand U410 (N_410,In_497,In_249);
nor U411 (N_411,In_476,In_298);
nand U412 (N_412,In_615,In_406);
nand U413 (N_413,In_576,In_104);
or U414 (N_414,In_749,In_597);
nand U415 (N_415,In_50,In_623);
or U416 (N_416,In_698,In_503);
and U417 (N_417,In_546,In_711);
nor U418 (N_418,In_427,In_80);
nand U419 (N_419,In_412,In_544);
and U420 (N_420,In_589,In_151);
and U421 (N_421,In_682,In_287);
nor U422 (N_422,In_624,In_414);
or U423 (N_423,In_25,In_313);
and U424 (N_424,In_449,In_51);
and U425 (N_425,In_427,In_711);
nor U426 (N_426,In_8,In_361);
nor U427 (N_427,In_626,In_362);
or U428 (N_428,In_257,In_725);
nor U429 (N_429,In_678,In_38);
or U430 (N_430,In_139,In_73);
nand U431 (N_431,In_116,In_386);
or U432 (N_432,In_72,In_308);
or U433 (N_433,In_183,In_38);
or U434 (N_434,In_236,In_112);
or U435 (N_435,In_704,In_421);
or U436 (N_436,In_304,In_705);
or U437 (N_437,In_286,In_130);
nand U438 (N_438,In_87,In_570);
or U439 (N_439,In_729,In_469);
nand U440 (N_440,In_643,In_499);
nor U441 (N_441,In_748,In_482);
or U442 (N_442,In_589,In_482);
xnor U443 (N_443,In_131,In_48);
or U444 (N_444,In_419,In_745);
or U445 (N_445,In_466,In_95);
nand U446 (N_446,In_445,In_304);
and U447 (N_447,In_91,In_6);
and U448 (N_448,In_641,In_22);
and U449 (N_449,In_577,In_338);
or U450 (N_450,In_343,In_509);
and U451 (N_451,In_466,In_227);
and U452 (N_452,In_622,In_618);
and U453 (N_453,In_558,In_475);
or U454 (N_454,In_257,In_347);
nand U455 (N_455,In_19,In_114);
or U456 (N_456,In_595,In_228);
nand U457 (N_457,In_472,In_39);
nand U458 (N_458,In_92,In_233);
nand U459 (N_459,In_91,In_67);
nand U460 (N_460,In_162,In_662);
nor U461 (N_461,In_603,In_605);
or U462 (N_462,In_595,In_15);
nor U463 (N_463,In_363,In_210);
and U464 (N_464,In_699,In_740);
or U465 (N_465,In_647,In_579);
or U466 (N_466,In_299,In_248);
nor U467 (N_467,In_730,In_686);
and U468 (N_468,In_670,In_472);
and U469 (N_469,In_480,In_723);
nor U470 (N_470,In_563,In_129);
nand U471 (N_471,In_340,In_354);
or U472 (N_472,In_588,In_548);
and U473 (N_473,In_690,In_255);
nand U474 (N_474,In_254,In_539);
and U475 (N_475,In_285,In_627);
nor U476 (N_476,In_682,In_316);
nor U477 (N_477,In_371,In_170);
nand U478 (N_478,In_383,In_551);
nand U479 (N_479,In_581,In_723);
and U480 (N_480,In_685,In_521);
or U481 (N_481,In_726,In_500);
nor U482 (N_482,In_709,In_3);
or U483 (N_483,In_229,In_663);
and U484 (N_484,In_144,In_442);
or U485 (N_485,In_76,In_220);
or U486 (N_486,In_691,In_168);
nor U487 (N_487,In_477,In_415);
and U488 (N_488,In_707,In_652);
nand U489 (N_489,In_664,In_663);
or U490 (N_490,In_355,In_682);
nand U491 (N_491,In_628,In_650);
or U492 (N_492,In_493,In_644);
or U493 (N_493,In_59,In_164);
nor U494 (N_494,In_498,In_597);
or U495 (N_495,In_275,In_736);
nor U496 (N_496,In_541,In_177);
and U497 (N_497,In_583,In_49);
nand U498 (N_498,In_440,In_467);
nand U499 (N_499,In_334,In_569);
and U500 (N_500,In_31,In_368);
and U501 (N_501,In_364,In_537);
nor U502 (N_502,In_469,In_382);
nand U503 (N_503,In_420,In_16);
nand U504 (N_504,In_365,In_349);
nor U505 (N_505,In_550,In_727);
nand U506 (N_506,In_426,In_635);
nor U507 (N_507,In_467,In_278);
or U508 (N_508,In_475,In_336);
and U509 (N_509,In_117,In_268);
nor U510 (N_510,In_634,In_246);
or U511 (N_511,In_136,In_707);
nand U512 (N_512,In_96,In_283);
nand U513 (N_513,In_688,In_588);
nor U514 (N_514,In_737,In_742);
or U515 (N_515,In_410,In_321);
xor U516 (N_516,In_47,In_740);
nand U517 (N_517,In_3,In_494);
nand U518 (N_518,In_726,In_401);
nor U519 (N_519,In_86,In_234);
or U520 (N_520,In_694,In_127);
nor U521 (N_521,In_72,In_661);
and U522 (N_522,In_268,In_347);
nand U523 (N_523,In_558,In_310);
nand U524 (N_524,In_495,In_517);
nand U525 (N_525,In_430,In_597);
or U526 (N_526,In_280,In_515);
nor U527 (N_527,In_69,In_60);
nor U528 (N_528,In_230,In_181);
or U529 (N_529,In_731,In_703);
or U530 (N_530,In_534,In_276);
nand U531 (N_531,In_183,In_674);
nand U532 (N_532,In_408,In_498);
nand U533 (N_533,In_637,In_548);
nand U534 (N_534,In_237,In_654);
and U535 (N_535,In_628,In_161);
and U536 (N_536,In_724,In_246);
nand U537 (N_537,In_533,In_206);
nand U538 (N_538,In_394,In_7);
nor U539 (N_539,In_219,In_615);
or U540 (N_540,In_395,In_728);
or U541 (N_541,In_482,In_734);
and U542 (N_542,In_3,In_675);
nand U543 (N_543,In_213,In_251);
nand U544 (N_544,In_8,In_29);
or U545 (N_545,In_344,In_397);
or U546 (N_546,In_625,In_712);
and U547 (N_547,In_529,In_685);
and U548 (N_548,In_417,In_186);
and U549 (N_549,In_18,In_213);
nand U550 (N_550,In_476,In_97);
and U551 (N_551,In_389,In_203);
and U552 (N_552,In_472,In_21);
or U553 (N_553,In_375,In_417);
nor U554 (N_554,In_284,In_124);
nand U555 (N_555,In_141,In_62);
nand U556 (N_556,In_171,In_721);
nor U557 (N_557,In_122,In_590);
or U558 (N_558,In_278,In_29);
and U559 (N_559,In_628,In_479);
nor U560 (N_560,In_241,In_81);
or U561 (N_561,In_571,In_150);
nand U562 (N_562,In_686,In_167);
and U563 (N_563,In_511,In_102);
and U564 (N_564,In_51,In_526);
or U565 (N_565,In_4,In_350);
and U566 (N_566,In_96,In_681);
or U567 (N_567,In_407,In_64);
nand U568 (N_568,In_314,In_603);
or U569 (N_569,In_405,In_73);
nand U570 (N_570,In_474,In_596);
or U571 (N_571,In_529,In_326);
nor U572 (N_572,In_46,In_298);
nor U573 (N_573,In_427,In_520);
and U574 (N_574,In_226,In_231);
or U575 (N_575,In_18,In_273);
nor U576 (N_576,In_578,In_243);
or U577 (N_577,In_491,In_359);
nand U578 (N_578,In_97,In_346);
or U579 (N_579,In_404,In_452);
and U580 (N_580,In_486,In_5);
or U581 (N_581,In_158,In_99);
nand U582 (N_582,In_568,In_70);
or U583 (N_583,In_498,In_62);
nand U584 (N_584,In_399,In_293);
and U585 (N_585,In_245,In_723);
or U586 (N_586,In_121,In_621);
or U587 (N_587,In_89,In_665);
nand U588 (N_588,In_70,In_170);
nor U589 (N_589,In_100,In_155);
or U590 (N_590,In_320,In_670);
nor U591 (N_591,In_501,In_203);
and U592 (N_592,In_93,In_728);
or U593 (N_593,In_404,In_263);
nor U594 (N_594,In_554,In_465);
nor U595 (N_595,In_421,In_259);
or U596 (N_596,In_356,In_123);
nor U597 (N_597,In_490,In_101);
and U598 (N_598,In_506,In_74);
nor U599 (N_599,In_329,In_215);
nor U600 (N_600,In_350,In_77);
and U601 (N_601,In_641,In_48);
nand U602 (N_602,In_285,In_283);
nor U603 (N_603,In_407,In_627);
and U604 (N_604,In_538,In_38);
or U605 (N_605,In_682,In_375);
nand U606 (N_606,In_499,In_431);
or U607 (N_607,In_540,In_423);
xor U608 (N_608,In_659,In_484);
and U609 (N_609,In_184,In_57);
nand U610 (N_610,In_6,In_72);
nand U611 (N_611,In_490,In_244);
or U612 (N_612,In_348,In_617);
or U613 (N_613,In_717,In_4);
or U614 (N_614,In_234,In_336);
or U615 (N_615,In_573,In_527);
or U616 (N_616,In_745,In_138);
nor U617 (N_617,In_277,In_417);
or U618 (N_618,In_8,In_295);
xor U619 (N_619,In_620,In_190);
or U620 (N_620,In_722,In_671);
nor U621 (N_621,In_192,In_632);
nor U622 (N_622,In_598,In_717);
or U623 (N_623,In_571,In_124);
and U624 (N_624,In_434,In_77);
or U625 (N_625,In_56,In_184);
and U626 (N_626,In_518,In_495);
or U627 (N_627,In_1,In_43);
and U628 (N_628,In_345,In_740);
nand U629 (N_629,In_130,In_152);
nor U630 (N_630,In_354,In_198);
nand U631 (N_631,In_632,In_77);
or U632 (N_632,In_260,In_363);
nand U633 (N_633,In_163,In_72);
xnor U634 (N_634,In_740,In_518);
nand U635 (N_635,In_592,In_24);
and U636 (N_636,In_383,In_397);
nor U637 (N_637,In_326,In_458);
and U638 (N_638,In_437,In_15);
nor U639 (N_639,In_466,In_308);
nor U640 (N_640,In_170,In_42);
nand U641 (N_641,In_552,In_346);
nor U642 (N_642,In_475,In_540);
and U643 (N_643,In_82,In_194);
nand U644 (N_644,In_101,In_721);
nor U645 (N_645,In_68,In_417);
nor U646 (N_646,In_427,In_356);
and U647 (N_647,In_90,In_229);
nand U648 (N_648,In_140,In_463);
nand U649 (N_649,In_686,In_439);
or U650 (N_650,In_645,In_220);
and U651 (N_651,In_424,In_300);
nor U652 (N_652,In_66,In_451);
or U653 (N_653,In_186,In_288);
nand U654 (N_654,In_733,In_40);
or U655 (N_655,In_534,In_257);
nor U656 (N_656,In_13,In_167);
or U657 (N_657,In_171,In_689);
or U658 (N_658,In_323,In_244);
nand U659 (N_659,In_610,In_299);
and U660 (N_660,In_505,In_332);
or U661 (N_661,In_735,In_728);
or U662 (N_662,In_41,In_504);
and U663 (N_663,In_747,In_433);
nand U664 (N_664,In_265,In_99);
or U665 (N_665,In_274,In_257);
or U666 (N_666,In_402,In_306);
nand U667 (N_667,In_156,In_596);
nand U668 (N_668,In_678,In_223);
or U669 (N_669,In_675,In_386);
or U670 (N_670,In_478,In_541);
nand U671 (N_671,In_446,In_537);
nor U672 (N_672,In_235,In_71);
or U673 (N_673,In_526,In_600);
nor U674 (N_674,In_179,In_569);
or U675 (N_675,In_530,In_57);
and U676 (N_676,In_637,In_560);
and U677 (N_677,In_247,In_684);
or U678 (N_678,In_413,In_537);
or U679 (N_679,In_255,In_211);
or U680 (N_680,In_122,In_719);
nand U681 (N_681,In_369,In_29);
nor U682 (N_682,In_189,In_249);
and U683 (N_683,In_666,In_221);
nand U684 (N_684,In_221,In_102);
nor U685 (N_685,In_430,In_75);
nor U686 (N_686,In_283,In_43);
or U687 (N_687,In_487,In_385);
nand U688 (N_688,In_251,In_434);
nand U689 (N_689,In_724,In_411);
and U690 (N_690,In_25,In_189);
or U691 (N_691,In_498,In_218);
or U692 (N_692,In_386,In_193);
and U693 (N_693,In_533,In_23);
and U694 (N_694,In_240,In_315);
nand U695 (N_695,In_300,In_490);
nor U696 (N_696,In_306,In_707);
or U697 (N_697,In_165,In_136);
or U698 (N_698,In_536,In_618);
and U699 (N_699,In_508,In_627);
or U700 (N_700,In_246,In_300);
and U701 (N_701,In_46,In_535);
and U702 (N_702,In_472,In_728);
nor U703 (N_703,In_342,In_303);
or U704 (N_704,In_194,In_706);
xor U705 (N_705,In_706,In_413);
or U706 (N_706,In_49,In_167);
or U707 (N_707,In_192,In_644);
nor U708 (N_708,In_346,In_200);
and U709 (N_709,In_439,In_536);
or U710 (N_710,In_526,In_307);
nor U711 (N_711,In_75,In_303);
nor U712 (N_712,In_311,In_691);
and U713 (N_713,In_459,In_246);
or U714 (N_714,In_442,In_31);
nor U715 (N_715,In_394,In_716);
and U716 (N_716,In_304,In_257);
or U717 (N_717,In_102,In_283);
nand U718 (N_718,In_653,In_438);
nand U719 (N_719,In_418,In_464);
nand U720 (N_720,In_526,In_159);
and U721 (N_721,In_547,In_409);
nand U722 (N_722,In_130,In_627);
nand U723 (N_723,In_442,In_283);
and U724 (N_724,In_681,In_580);
or U725 (N_725,In_525,In_618);
and U726 (N_726,In_555,In_138);
or U727 (N_727,In_301,In_623);
or U728 (N_728,In_333,In_160);
nand U729 (N_729,In_292,In_695);
nand U730 (N_730,In_404,In_230);
and U731 (N_731,In_476,In_455);
nor U732 (N_732,In_448,In_724);
nor U733 (N_733,In_35,In_401);
nand U734 (N_734,In_444,In_211);
or U735 (N_735,In_727,In_280);
nor U736 (N_736,In_85,In_618);
and U737 (N_737,In_242,In_233);
nor U738 (N_738,In_168,In_164);
and U739 (N_739,In_319,In_217);
or U740 (N_740,In_55,In_472);
nand U741 (N_741,In_341,In_395);
or U742 (N_742,In_38,In_734);
nor U743 (N_743,In_670,In_402);
and U744 (N_744,In_477,In_592);
nor U745 (N_745,In_455,In_88);
and U746 (N_746,In_69,In_694);
nor U747 (N_747,In_239,In_70);
or U748 (N_748,In_489,In_652);
nor U749 (N_749,In_343,In_724);
nand U750 (N_750,In_171,In_285);
nand U751 (N_751,In_681,In_661);
nand U752 (N_752,In_489,In_85);
and U753 (N_753,In_111,In_207);
or U754 (N_754,In_89,In_99);
and U755 (N_755,In_75,In_669);
or U756 (N_756,In_492,In_37);
nor U757 (N_757,In_631,In_614);
nand U758 (N_758,In_119,In_38);
or U759 (N_759,In_35,In_166);
or U760 (N_760,In_671,In_124);
and U761 (N_761,In_281,In_83);
and U762 (N_762,In_274,In_198);
nand U763 (N_763,In_76,In_552);
and U764 (N_764,In_27,In_68);
nand U765 (N_765,In_198,In_141);
nor U766 (N_766,In_547,In_76);
nand U767 (N_767,In_389,In_129);
nor U768 (N_768,In_332,In_664);
nand U769 (N_769,In_158,In_180);
nor U770 (N_770,In_185,In_716);
and U771 (N_771,In_428,In_568);
or U772 (N_772,In_645,In_147);
nand U773 (N_773,In_18,In_652);
and U774 (N_774,In_371,In_400);
and U775 (N_775,In_342,In_587);
and U776 (N_776,In_244,In_164);
nor U777 (N_777,In_737,In_602);
and U778 (N_778,In_712,In_738);
nor U779 (N_779,In_268,In_472);
nand U780 (N_780,In_524,In_7);
nor U781 (N_781,In_481,In_523);
or U782 (N_782,In_686,In_259);
nand U783 (N_783,In_88,In_585);
nor U784 (N_784,In_663,In_466);
nor U785 (N_785,In_44,In_723);
and U786 (N_786,In_7,In_456);
and U787 (N_787,In_169,In_522);
nor U788 (N_788,In_111,In_460);
and U789 (N_789,In_274,In_285);
nand U790 (N_790,In_612,In_244);
nand U791 (N_791,In_303,In_699);
nand U792 (N_792,In_728,In_174);
or U793 (N_793,In_225,In_734);
nor U794 (N_794,In_1,In_675);
nor U795 (N_795,In_341,In_580);
nor U796 (N_796,In_219,In_131);
and U797 (N_797,In_554,In_289);
nand U798 (N_798,In_297,In_164);
nand U799 (N_799,In_477,In_632);
nor U800 (N_800,In_557,In_515);
nand U801 (N_801,In_310,In_88);
nand U802 (N_802,In_694,In_75);
nor U803 (N_803,In_370,In_338);
or U804 (N_804,In_377,In_719);
or U805 (N_805,In_189,In_459);
nor U806 (N_806,In_675,In_658);
and U807 (N_807,In_424,In_462);
nor U808 (N_808,In_549,In_545);
or U809 (N_809,In_448,In_723);
nor U810 (N_810,In_330,In_121);
xor U811 (N_811,In_295,In_666);
or U812 (N_812,In_301,In_727);
and U813 (N_813,In_113,In_688);
and U814 (N_814,In_578,In_87);
or U815 (N_815,In_339,In_8);
nand U816 (N_816,In_28,In_197);
nand U817 (N_817,In_716,In_603);
and U818 (N_818,In_716,In_436);
and U819 (N_819,In_376,In_47);
and U820 (N_820,In_69,In_457);
and U821 (N_821,In_578,In_198);
nor U822 (N_822,In_209,In_624);
and U823 (N_823,In_307,In_479);
nand U824 (N_824,In_417,In_359);
nor U825 (N_825,In_486,In_89);
or U826 (N_826,In_524,In_292);
xnor U827 (N_827,In_605,In_380);
nand U828 (N_828,In_553,In_711);
or U829 (N_829,In_166,In_323);
nor U830 (N_830,In_69,In_485);
and U831 (N_831,In_619,In_718);
nor U832 (N_832,In_56,In_125);
and U833 (N_833,In_148,In_125);
nor U834 (N_834,In_734,In_339);
and U835 (N_835,In_7,In_719);
nor U836 (N_836,In_345,In_514);
nand U837 (N_837,In_269,In_293);
or U838 (N_838,In_422,In_404);
or U839 (N_839,In_331,In_145);
and U840 (N_840,In_64,In_174);
and U841 (N_841,In_432,In_510);
and U842 (N_842,In_292,In_133);
and U843 (N_843,In_638,In_41);
or U844 (N_844,In_180,In_38);
or U845 (N_845,In_652,In_236);
nand U846 (N_846,In_738,In_655);
or U847 (N_847,In_5,In_127);
nand U848 (N_848,In_398,In_190);
and U849 (N_849,In_660,In_740);
nor U850 (N_850,In_60,In_278);
nand U851 (N_851,In_512,In_644);
nor U852 (N_852,In_626,In_637);
and U853 (N_853,In_698,In_571);
or U854 (N_854,In_328,In_544);
nor U855 (N_855,In_130,In_735);
and U856 (N_856,In_461,In_728);
and U857 (N_857,In_312,In_446);
or U858 (N_858,In_509,In_95);
nor U859 (N_859,In_254,In_13);
nor U860 (N_860,In_608,In_513);
nand U861 (N_861,In_21,In_5);
and U862 (N_862,In_294,In_162);
and U863 (N_863,In_319,In_473);
nor U864 (N_864,In_666,In_67);
or U865 (N_865,In_189,In_16);
or U866 (N_866,In_630,In_50);
and U867 (N_867,In_513,In_415);
and U868 (N_868,In_616,In_487);
or U869 (N_869,In_558,In_37);
nor U870 (N_870,In_563,In_487);
or U871 (N_871,In_442,In_116);
nor U872 (N_872,In_522,In_258);
nand U873 (N_873,In_729,In_747);
nor U874 (N_874,In_571,In_218);
nand U875 (N_875,In_296,In_165);
and U876 (N_876,In_195,In_156);
nand U877 (N_877,In_676,In_339);
nor U878 (N_878,In_405,In_593);
and U879 (N_879,In_356,In_68);
nand U880 (N_880,In_405,In_225);
and U881 (N_881,In_739,In_77);
nor U882 (N_882,In_420,In_169);
nor U883 (N_883,In_332,In_131);
nor U884 (N_884,In_707,In_217);
nand U885 (N_885,In_295,In_90);
nand U886 (N_886,In_87,In_161);
or U887 (N_887,In_639,In_470);
nand U888 (N_888,In_591,In_593);
nor U889 (N_889,In_566,In_469);
nand U890 (N_890,In_747,In_280);
nand U891 (N_891,In_397,In_234);
nor U892 (N_892,In_360,In_476);
nand U893 (N_893,In_37,In_414);
nand U894 (N_894,In_91,In_90);
and U895 (N_895,In_48,In_516);
nor U896 (N_896,In_317,In_428);
and U897 (N_897,In_162,In_397);
and U898 (N_898,In_685,In_572);
or U899 (N_899,In_442,In_83);
or U900 (N_900,In_224,In_480);
and U901 (N_901,In_352,In_49);
nand U902 (N_902,In_492,In_160);
and U903 (N_903,In_3,In_666);
nand U904 (N_904,In_491,In_626);
xor U905 (N_905,In_31,In_596);
nand U906 (N_906,In_349,In_42);
nand U907 (N_907,In_586,In_577);
nor U908 (N_908,In_352,In_0);
and U909 (N_909,In_416,In_550);
and U910 (N_910,In_406,In_1);
nor U911 (N_911,In_458,In_332);
and U912 (N_912,In_142,In_367);
nand U913 (N_913,In_275,In_318);
and U914 (N_914,In_142,In_314);
or U915 (N_915,In_442,In_701);
or U916 (N_916,In_388,In_307);
nor U917 (N_917,In_228,In_622);
or U918 (N_918,In_542,In_367);
or U919 (N_919,In_113,In_56);
nor U920 (N_920,In_300,In_291);
nand U921 (N_921,In_533,In_538);
nor U922 (N_922,In_365,In_433);
nor U923 (N_923,In_559,In_316);
nor U924 (N_924,In_640,In_121);
nor U925 (N_925,In_268,In_738);
and U926 (N_926,In_129,In_499);
and U927 (N_927,In_703,In_338);
or U928 (N_928,In_296,In_134);
and U929 (N_929,In_583,In_270);
and U930 (N_930,In_680,In_258);
or U931 (N_931,In_324,In_706);
or U932 (N_932,In_203,In_652);
and U933 (N_933,In_435,In_156);
and U934 (N_934,In_655,In_416);
nand U935 (N_935,In_382,In_33);
nor U936 (N_936,In_135,In_253);
or U937 (N_937,In_137,In_585);
nand U938 (N_938,In_56,In_49);
nand U939 (N_939,In_155,In_98);
and U940 (N_940,In_600,In_506);
nand U941 (N_941,In_509,In_510);
nor U942 (N_942,In_74,In_34);
nand U943 (N_943,In_112,In_256);
nor U944 (N_944,In_701,In_625);
and U945 (N_945,In_683,In_179);
nand U946 (N_946,In_509,In_43);
and U947 (N_947,In_286,In_624);
nor U948 (N_948,In_247,In_81);
nor U949 (N_949,In_588,In_431);
nand U950 (N_950,In_715,In_508);
nand U951 (N_951,In_220,In_296);
and U952 (N_952,In_107,In_128);
or U953 (N_953,In_613,In_305);
nand U954 (N_954,In_456,In_54);
or U955 (N_955,In_57,In_515);
nand U956 (N_956,In_394,In_343);
and U957 (N_957,In_327,In_245);
nand U958 (N_958,In_530,In_271);
and U959 (N_959,In_200,In_625);
and U960 (N_960,In_239,In_58);
nand U961 (N_961,In_382,In_455);
or U962 (N_962,In_376,In_744);
nor U963 (N_963,In_345,In_18);
and U964 (N_964,In_87,In_486);
nand U965 (N_965,In_740,In_248);
nor U966 (N_966,In_174,In_378);
xor U967 (N_967,In_680,In_253);
nand U968 (N_968,In_81,In_412);
and U969 (N_969,In_461,In_161);
nor U970 (N_970,In_684,In_413);
nand U971 (N_971,In_682,In_658);
nor U972 (N_972,In_278,In_355);
nand U973 (N_973,In_342,In_722);
and U974 (N_974,In_388,In_25);
nor U975 (N_975,In_647,In_44);
and U976 (N_976,In_690,In_205);
or U977 (N_977,In_348,In_298);
and U978 (N_978,In_335,In_337);
and U979 (N_979,In_440,In_652);
nor U980 (N_980,In_303,In_512);
and U981 (N_981,In_36,In_21);
nor U982 (N_982,In_233,In_462);
nand U983 (N_983,In_288,In_322);
or U984 (N_984,In_510,In_124);
nand U985 (N_985,In_164,In_553);
nor U986 (N_986,In_97,In_140);
nor U987 (N_987,In_562,In_678);
and U988 (N_988,In_467,In_107);
nand U989 (N_989,In_299,In_38);
and U990 (N_990,In_386,In_84);
and U991 (N_991,In_31,In_339);
and U992 (N_992,In_440,In_180);
or U993 (N_993,In_559,In_63);
nor U994 (N_994,In_497,In_513);
and U995 (N_995,In_718,In_108);
nor U996 (N_996,In_566,In_162);
nand U997 (N_997,In_122,In_562);
nor U998 (N_998,In_440,In_302);
or U999 (N_999,In_168,In_582);
and U1000 (N_1000,N_353,N_405);
nand U1001 (N_1001,N_46,N_293);
nand U1002 (N_1002,N_453,N_852);
xor U1003 (N_1003,N_845,N_724);
or U1004 (N_1004,N_422,N_135);
nand U1005 (N_1005,N_654,N_421);
nor U1006 (N_1006,N_31,N_496);
and U1007 (N_1007,N_419,N_344);
and U1008 (N_1008,N_793,N_837);
and U1009 (N_1009,N_139,N_786);
nor U1010 (N_1010,N_528,N_578);
nand U1011 (N_1011,N_36,N_318);
nor U1012 (N_1012,N_39,N_471);
nor U1013 (N_1013,N_708,N_533);
nand U1014 (N_1014,N_914,N_412);
nor U1015 (N_1015,N_427,N_362);
nor U1016 (N_1016,N_820,N_683);
xnor U1017 (N_1017,N_545,N_463);
and U1018 (N_1018,N_359,N_541);
nor U1019 (N_1019,N_785,N_704);
or U1020 (N_1020,N_870,N_464);
nand U1021 (N_1021,N_637,N_717);
nand U1022 (N_1022,N_896,N_180);
nand U1023 (N_1023,N_383,N_681);
nand U1024 (N_1024,N_977,N_238);
nor U1025 (N_1025,N_961,N_885);
and U1026 (N_1026,N_175,N_140);
nor U1027 (N_1027,N_286,N_466);
or U1028 (N_1028,N_842,N_354);
or U1029 (N_1029,N_160,N_342);
or U1030 (N_1030,N_282,N_571);
or U1031 (N_1031,N_984,N_397);
or U1032 (N_1032,N_592,N_289);
nand U1033 (N_1033,N_436,N_16);
nor U1034 (N_1034,N_410,N_61);
nand U1035 (N_1035,N_809,N_916);
or U1036 (N_1036,N_957,N_220);
and U1037 (N_1037,N_511,N_10);
nor U1038 (N_1038,N_983,N_875);
nor U1039 (N_1039,N_542,N_27);
and U1040 (N_1040,N_121,N_881);
or U1041 (N_1041,N_231,N_894);
nand U1042 (N_1042,N_259,N_271);
nor U1043 (N_1043,N_260,N_822);
and U1044 (N_1044,N_166,N_806);
nor U1045 (N_1045,N_742,N_168);
and U1046 (N_1046,N_304,N_653);
and U1047 (N_1047,N_905,N_561);
and U1048 (N_1048,N_538,N_426);
nor U1049 (N_1049,N_13,N_555);
nand U1050 (N_1050,N_937,N_425);
or U1051 (N_1051,N_150,N_442);
xnor U1052 (N_1052,N_931,N_367);
nand U1053 (N_1053,N_141,N_674);
nand U1054 (N_1054,N_660,N_727);
nor U1055 (N_1055,N_735,N_276);
nand U1056 (N_1056,N_262,N_940);
or U1057 (N_1057,N_156,N_67);
nor U1058 (N_1058,N_802,N_266);
nand U1059 (N_1059,N_366,N_715);
nand U1060 (N_1060,N_219,N_142);
nor U1061 (N_1061,N_115,N_668);
and U1062 (N_1062,N_756,N_672);
nor U1063 (N_1063,N_981,N_301);
nor U1064 (N_1064,N_759,N_402);
nor U1065 (N_1065,N_805,N_586);
nand U1066 (N_1066,N_41,N_853);
nor U1067 (N_1067,N_394,N_11);
nor U1068 (N_1068,N_192,N_546);
nor U1069 (N_1069,N_745,N_468);
and U1070 (N_1070,N_866,N_638);
and U1071 (N_1071,N_491,N_275);
and U1072 (N_1072,N_749,N_803);
nor U1073 (N_1073,N_146,N_165);
nand U1074 (N_1074,N_928,N_428);
nor U1075 (N_1075,N_54,N_549);
xor U1076 (N_1076,N_713,N_960);
or U1077 (N_1077,N_524,N_830);
or U1078 (N_1078,N_310,N_242);
and U1079 (N_1079,N_987,N_450);
or U1080 (N_1080,N_923,N_243);
and U1081 (N_1081,N_544,N_89);
and U1082 (N_1082,N_161,N_687);
or U1083 (N_1083,N_859,N_563);
or U1084 (N_1084,N_609,N_201);
nor U1085 (N_1085,N_66,N_57);
nor U1086 (N_1086,N_195,N_693);
xor U1087 (N_1087,N_514,N_955);
nor U1088 (N_1088,N_445,N_626);
nand U1089 (N_1089,N_663,N_157);
nand U1090 (N_1090,N_123,N_530);
and U1091 (N_1091,N_547,N_883);
nand U1092 (N_1092,N_413,N_677);
and U1093 (N_1093,N_936,N_839);
xor U1094 (N_1094,N_824,N_212);
and U1095 (N_1095,N_565,N_337);
and U1096 (N_1096,N_331,N_874);
nand U1097 (N_1097,N_732,N_50);
or U1098 (N_1098,N_574,N_840);
nor U1099 (N_1099,N_87,N_813);
or U1100 (N_1100,N_921,N_433);
xor U1101 (N_1101,N_227,N_700);
nor U1102 (N_1102,N_128,N_944);
nor U1103 (N_1103,N_373,N_296);
nor U1104 (N_1104,N_6,N_808);
nand U1105 (N_1105,N_313,N_652);
nor U1106 (N_1106,N_440,N_986);
nand U1107 (N_1107,N_409,N_593);
nor U1108 (N_1108,N_982,N_810);
or U1109 (N_1109,N_543,N_863);
nand U1110 (N_1110,N_850,N_945);
nor U1111 (N_1111,N_90,N_540);
and U1112 (N_1112,N_206,N_119);
nor U1113 (N_1113,N_927,N_392);
or U1114 (N_1114,N_284,N_203);
nor U1115 (N_1115,N_971,N_340);
nor U1116 (N_1116,N_692,N_489);
or U1117 (N_1117,N_278,N_671);
and U1118 (N_1118,N_964,N_216);
and U1119 (N_1119,N_181,N_188);
or U1120 (N_1120,N_688,N_457);
nand U1121 (N_1121,N_832,N_817);
nor U1122 (N_1122,N_886,N_795);
nor U1123 (N_1123,N_779,N_281);
nor U1124 (N_1124,N_416,N_300);
and U1125 (N_1125,N_209,N_920);
nand U1126 (N_1126,N_77,N_30);
or U1127 (N_1127,N_903,N_12);
or U1128 (N_1128,N_917,N_703);
nand U1129 (N_1129,N_694,N_689);
nand U1130 (N_1130,N_930,N_826);
and U1131 (N_1131,N_437,N_499);
nor U1132 (N_1132,N_163,N_629);
nand U1133 (N_1133,N_179,N_14);
or U1134 (N_1134,N_28,N_974);
or U1135 (N_1135,N_843,N_448);
xor U1136 (N_1136,N_909,N_241);
nor U1137 (N_1137,N_904,N_627);
or U1138 (N_1138,N_228,N_958);
nand U1139 (N_1139,N_603,N_125);
and U1140 (N_1140,N_835,N_919);
or U1141 (N_1141,N_531,N_420);
and U1142 (N_1142,N_218,N_579);
nor U1143 (N_1143,N_854,N_939);
nor U1144 (N_1144,N_49,N_458);
and U1145 (N_1145,N_942,N_235);
nor U1146 (N_1146,N_83,N_941);
and U1147 (N_1147,N_632,N_617);
nand U1148 (N_1148,N_104,N_967);
and U1149 (N_1149,N_43,N_486);
and U1150 (N_1150,N_605,N_82);
and U1151 (N_1151,N_208,N_539);
or U1152 (N_1152,N_746,N_666);
nor U1153 (N_1153,N_35,N_347);
nand U1154 (N_1154,N_762,N_72);
nand U1155 (N_1155,N_643,N_678);
nand U1156 (N_1156,N_40,N_370);
and U1157 (N_1157,N_709,N_37);
or U1158 (N_1158,N_829,N_773);
and U1159 (N_1159,N_225,N_947);
nand U1160 (N_1160,N_9,N_664);
and U1161 (N_1161,N_751,N_979);
nor U1162 (N_1162,N_473,N_583);
or U1163 (N_1163,N_312,N_601);
nor U1164 (N_1164,N_630,N_966);
nor U1165 (N_1165,N_730,N_645);
and U1166 (N_1166,N_294,N_116);
nand U1167 (N_1167,N_623,N_641);
nand U1168 (N_1168,N_484,N_815);
and U1169 (N_1169,N_34,N_145);
nor U1170 (N_1170,N_963,N_127);
or U1171 (N_1171,N_912,N_0);
and U1172 (N_1172,N_106,N_949);
and U1173 (N_1173,N_910,N_868);
nor U1174 (N_1174,N_96,N_189);
nand U1175 (N_1175,N_134,N_918);
or U1176 (N_1176,N_559,N_245);
or U1177 (N_1177,N_274,N_758);
and U1178 (N_1178,N_222,N_532);
xnor U1179 (N_1179,N_118,N_349);
and U1180 (N_1180,N_71,N_752);
or U1181 (N_1181,N_307,N_269);
nor U1182 (N_1182,N_60,N_887);
and U1183 (N_1183,N_807,N_505);
nand U1184 (N_1184,N_415,N_319);
or U1185 (N_1185,N_358,N_257);
nand U1186 (N_1186,N_952,N_679);
or U1187 (N_1187,N_714,N_953);
and U1188 (N_1188,N_595,N_577);
nand U1189 (N_1189,N_741,N_535);
and U1190 (N_1190,N_492,N_47);
nand U1191 (N_1191,N_495,N_298);
nor U1192 (N_1192,N_568,N_596);
or U1193 (N_1193,N_459,N_103);
nor U1194 (N_1194,N_816,N_512);
or U1195 (N_1195,N_314,N_120);
or U1196 (N_1196,N_465,N_92);
or U1197 (N_1197,N_232,N_285);
or U1198 (N_1198,N_556,N_44);
nand U1199 (N_1199,N_109,N_202);
or U1200 (N_1200,N_754,N_335);
nand U1201 (N_1201,N_330,N_787);
and U1202 (N_1202,N_333,N_283);
nor U1203 (N_1203,N_265,N_411);
nor U1204 (N_1204,N_833,N_508);
nand U1205 (N_1205,N_193,N_480);
and U1206 (N_1206,N_51,N_604);
or U1207 (N_1207,N_889,N_913);
nand U1208 (N_1208,N_934,N_174);
nand U1209 (N_1209,N_733,N_747);
and U1210 (N_1210,N_915,N_136);
and U1211 (N_1211,N_587,N_101);
nor U1212 (N_1212,N_521,N_256);
or U1213 (N_1213,N_110,N_53);
nor U1214 (N_1214,N_898,N_591);
and U1215 (N_1215,N_435,N_107);
nor U1216 (N_1216,N_871,N_761);
or U1217 (N_1217,N_778,N_764);
or U1218 (N_1218,N_226,N_736);
nor U1219 (N_1219,N_73,N_951);
nor U1220 (N_1220,N_847,N_959);
nor U1221 (N_1221,N_381,N_170);
and U1222 (N_1222,N_861,N_324);
and U1223 (N_1223,N_962,N_223);
and U1224 (N_1224,N_207,N_376);
or U1225 (N_1225,N_393,N_15);
nor U1226 (N_1226,N_562,N_607);
nand U1227 (N_1227,N_796,N_315);
nand U1228 (N_1228,N_551,N_444);
nor U1229 (N_1229,N_728,N_251);
or U1230 (N_1230,N_336,N_851);
and U1231 (N_1231,N_989,N_720);
and U1232 (N_1232,N_460,N_503);
nor U1233 (N_1233,N_738,N_299);
or U1234 (N_1234,N_548,N_650);
or U1235 (N_1235,N_608,N_569);
or U1236 (N_1236,N_84,N_701);
nand U1237 (N_1237,N_210,N_234);
nand U1238 (N_1238,N_352,N_321);
nor U1239 (N_1239,N_375,N_481);
nand U1240 (N_1240,N_661,N_613);
nor U1241 (N_1241,N_857,N_363);
or U1242 (N_1242,N_99,N_865);
or U1243 (N_1243,N_884,N_554);
nand U1244 (N_1244,N_472,N_599);
nor U1245 (N_1245,N_424,N_323);
or U1246 (N_1246,N_879,N_770);
nand U1247 (N_1247,N_902,N_476);
nand U1248 (N_1248,N_369,N_765);
and U1249 (N_1249,N_997,N_306);
or U1250 (N_1250,N_65,N_867);
nor U1251 (N_1251,N_792,N_311);
nor U1252 (N_1252,N_408,N_684);
or U1253 (N_1253,N_860,N_988);
and U1254 (N_1254,N_308,N_901);
nand U1255 (N_1255,N_838,N_911);
xor U1256 (N_1256,N_699,N_564);
or U1257 (N_1257,N_357,N_938);
and U1258 (N_1258,N_848,N_244);
nor U1259 (N_1259,N_976,N_753);
or U1260 (N_1260,N_552,N_527);
or U1261 (N_1261,N_483,N_446);
nand U1262 (N_1262,N_1,N_924);
nand U1263 (N_1263,N_173,N_954);
and U1264 (N_1264,N_522,N_113);
nor U1265 (N_1265,N_589,N_182);
nor U1266 (N_1266,N_734,N_814);
nor U1267 (N_1267,N_297,N_204);
nand U1268 (N_1268,N_343,N_836);
nor U1269 (N_1269,N_517,N_111);
nand U1270 (N_1270,N_164,N_526);
nor U1271 (N_1271,N_152,N_112);
or U1272 (N_1272,N_737,N_263);
or U1273 (N_1273,N_975,N_510);
and U1274 (N_1274,N_518,N_154);
nand U1275 (N_1275,N_615,N_825);
and U1276 (N_1276,N_614,N_162);
and U1277 (N_1277,N_804,N_731);
nand U1278 (N_1278,N_774,N_659);
and U1279 (N_1279,N_144,N_711);
or U1280 (N_1280,N_633,N_240);
nand U1281 (N_1281,N_58,N_519);
nand U1282 (N_1282,N_620,N_8);
nor U1283 (N_1283,N_827,N_469);
or U1284 (N_1284,N_869,N_598);
and U1285 (N_1285,N_662,N_648);
and U1286 (N_1286,N_504,N_788);
nor U1287 (N_1287,N_585,N_611);
and U1288 (N_1288,N_288,N_619);
nand U1289 (N_1289,N_434,N_996);
or U1290 (N_1290,N_943,N_280);
nor U1291 (N_1291,N_763,N_171);
and U1292 (N_1292,N_247,N_783);
nand U1293 (N_1293,N_794,N_249);
nand U1294 (N_1294,N_355,N_612);
nand U1295 (N_1295,N_777,N_167);
nor U1296 (N_1296,N_682,N_258);
nand U1297 (N_1297,N_775,N_237);
and U1298 (N_1298,N_341,N_224);
nor U1299 (N_1299,N_364,N_719);
or U1300 (N_1300,N_186,N_757);
nor U1301 (N_1301,N_86,N_441);
nor U1302 (N_1302,N_891,N_117);
nor U1303 (N_1303,N_864,N_279);
nand U1304 (N_1304,N_669,N_214);
nor U1305 (N_1305,N_339,N_130);
nor U1306 (N_1306,N_980,N_590);
nand U1307 (N_1307,N_725,N_573);
and U1308 (N_1308,N_716,N_382);
nand U1309 (N_1309,N_76,N_858);
nand U1310 (N_1310,N_926,N_685);
or U1311 (N_1311,N_584,N_769);
nand U1312 (N_1312,N_326,N_114);
nand U1313 (N_1313,N_270,N_70);
or U1314 (N_1314,N_236,N_197);
xnor U1315 (N_1315,N_994,N_823);
nor U1316 (N_1316,N_365,N_21);
nand U1317 (N_1317,N_991,N_190);
nor U1318 (N_1318,N_801,N_429);
or U1319 (N_1319,N_3,N_760);
nand U1320 (N_1320,N_187,N_147);
nand U1321 (N_1321,N_890,N_882);
or U1322 (N_1322,N_834,N_475);
or U1323 (N_1323,N_215,N_969);
nor U1324 (N_1324,N_819,N_766);
nor U1325 (N_1325,N_452,N_722);
nand U1326 (N_1326,N_430,N_217);
and U1327 (N_1327,N_378,N_122);
nor U1328 (N_1328,N_493,N_893);
or U1329 (N_1329,N_148,N_62);
or U1330 (N_1330,N_316,N_529);
nor U1331 (N_1331,N_635,N_702);
and U1332 (N_1332,N_396,N_649);
and U1333 (N_1333,N_895,N_970);
or U1334 (N_1334,N_345,N_566);
or U1335 (N_1335,N_291,N_932);
nor U1336 (N_1336,N_557,N_973);
nor U1337 (N_1337,N_246,N_948);
nor U1338 (N_1338,N_634,N_933);
xnor U1339 (N_1339,N_892,N_509);
and U1340 (N_1340,N_513,N_184);
nand U1341 (N_1341,N_550,N_407);
nor U1342 (N_1342,N_348,N_644);
and U1343 (N_1343,N_377,N_24);
and U1344 (N_1344,N_897,N_52);
nand U1345 (N_1345,N_610,N_800);
and U1346 (N_1346,N_59,N_621);
and U1347 (N_1347,N_91,N_368);
nand U1348 (N_1348,N_327,N_196);
nand U1349 (N_1349,N_516,N_131);
or U1350 (N_1350,N_443,N_501);
and U1351 (N_1351,N_85,N_25);
or U1352 (N_1352,N_560,N_177);
and U1353 (N_1353,N_213,N_755);
nor U1354 (N_1354,N_618,N_844);
nand U1355 (N_1355,N_477,N_178);
or U1356 (N_1356,N_799,N_506);
or U1357 (N_1357,N_42,N_64);
or U1358 (N_1358,N_811,N_273);
or U1359 (N_1359,N_482,N_137);
and U1360 (N_1360,N_474,N_386);
nor U1361 (N_1361,N_329,N_38);
or U1362 (N_1362,N_100,N_487);
and U1363 (N_1363,N_520,N_438);
and U1364 (N_1364,N_199,N_723);
or U1365 (N_1365,N_780,N_675);
nand U1366 (N_1366,N_726,N_697);
or U1367 (N_1367,N_384,N_581);
nand U1368 (N_1368,N_782,N_351);
nor U1369 (N_1369,N_79,N_995);
or U1370 (N_1370,N_705,N_153);
nor U1371 (N_1371,N_628,N_129);
nand U1372 (N_1372,N_124,N_48);
nor U1373 (N_1373,N_325,N_69);
and U1374 (N_1374,N_639,N_385);
nand U1375 (N_1375,N_401,N_906);
and U1376 (N_1376,N_309,N_230);
nand U1377 (N_1377,N_862,N_588);
or U1378 (N_1378,N_828,N_696);
and U1379 (N_1379,N_622,N_255);
nor U1380 (N_1380,N_387,N_277);
or U1381 (N_1381,N_254,N_972);
nor U1382 (N_1382,N_439,N_706);
nor U1383 (N_1383,N_461,N_400);
nor U1384 (N_1384,N_740,N_264);
or U1385 (N_1385,N_831,N_360);
or U1386 (N_1386,N_138,N_158);
and U1387 (N_1387,N_470,N_5);
or U1388 (N_1388,N_2,N_55);
or U1389 (N_1389,N_676,N_398);
or U1390 (N_1390,N_32,N_56);
nand U1391 (N_1391,N_536,N_292);
and U1392 (N_1392,N_102,N_462);
or U1393 (N_1393,N_371,N_695);
nand U1394 (N_1394,N_821,N_771);
and U1395 (N_1395,N_198,N_624);
or U1396 (N_1396,N_956,N_781);
and U1397 (N_1397,N_640,N_744);
and U1398 (N_1398,N_176,N_880);
or U1399 (N_1399,N_572,N_673);
nor U1400 (N_1400,N_567,N_18);
or U1401 (N_1401,N_332,N_431);
nand U1402 (N_1402,N_346,N_935);
or U1403 (N_1403,N_380,N_303);
nor U1404 (N_1404,N_88,N_797);
nand U1405 (N_1405,N_149,N_126);
nand U1406 (N_1406,N_748,N_374);
and U1407 (N_1407,N_185,N_575);
and U1408 (N_1408,N_582,N_108);
and U1409 (N_1409,N_594,N_143);
or U1410 (N_1410,N_272,N_743);
nor U1411 (N_1411,N_183,N_23);
and U1412 (N_1412,N_287,N_647);
or U1413 (N_1413,N_239,N_646);
and U1414 (N_1414,N_523,N_534);
nor U1415 (N_1415,N_93,N_22);
and U1416 (N_1416,N_818,N_328);
nor U1417 (N_1417,N_159,N_625);
or U1418 (N_1418,N_75,N_602);
nand U1419 (N_1419,N_784,N_670);
nand U1420 (N_1420,N_925,N_45);
nand U1421 (N_1421,N_657,N_391);
nor U1422 (N_1422,N_686,N_81);
or U1423 (N_1423,N_631,N_295);
or U1424 (N_1424,N_950,N_878);
and U1425 (N_1425,N_389,N_155);
and U1426 (N_1426,N_479,N_636);
and U1427 (N_1427,N_507,N_356);
nor U1428 (N_1428,N_372,N_302);
and U1429 (N_1429,N_403,N_406);
and U1430 (N_1430,N_261,N_388);
or U1431 (N_1431,N_710,N_965);
nor U1432 (N_1432,N_712,N_856);
and U1433 (N_1433,N_877,N_929);
and U1434 (N_1434,N_233,N_772);
and U1435 (N_1435,N_908,N_449);
and U1436 (N_1436,N_322,N_600);
nand U1437 (N_1437,N_80,N_390);
nor U1438 (N_1438,N_497,N_132);
and U1439 (N_1439,N_515,N_350);
nor U1440 (N_1440,N_338,N_899);
nand U1441 (N_1441,N_789,N_68);
and U1442 (N_1442,N_451,N_580);
and U1443 (N_1443,N_667,N_7);
or U1444 (N_1444,N_97,N_194);
nand U1445 (N_1445,N_525,N_211);
and U1446 (N_1446,N_907,N_498);
or U1447 (N_1447,N_846,N_798);
or U1448 (N_1448,N_200,N_485);
nand U1449 (N_1449,N_985,N_361);
nand U1450 (N_1450,N_305,N_691);
nand U1451 (N_1451,N_999,N_698);
and U1452 (N_1452,N_418,N_729);
nor U1453 (N_1453,N_978,N_454);
and U1454 (N_1454,N_767,N_399);
nand U1455 (N_1455,N_721,N_20);
or U1456 (N_1456,N_776,N_998);
or U1457 (N_1457,N_221,N_768);
and U1458 (N_1458,N_395,N_500);
nand U1459 (N_1459,N_447,N_320);
nand U1460 (N_1460,N_252,N_841);
or U1461 (N_1461,N_250,N_98);
nand U1462 (N_1462,N_290,N_873);
nor U1463 (N_1463,N_537,N_4);
and U1464 (N_1464,N_490,N_169);
nand U1465 (N_1465,N_133,N_191);
nor U1466 (N_1466,N_268,N_95);
or U1467 (N_1467,N_172,N_94);
xnor U1468 (N_1468,N_922,N_990);
or U1469 (N_1469,N_558,N_105);
and U1470 (N_1470,N_467,N_690);
or U1471 (N_1471,N_253,N_78);
nand U1472 (N_1472,N_750,N_379);
nor U1473 (N_1473,N_656,N_33);
nand U1474 (N_1474,N_26,N_946);
or U1475 (N_1475,N_665,N_488);
nand U1476 (N_1476,N_229,N_791);
and U1477 (N_1477,N_968,N_849);
nor U1478 (N_1478,N_456,N_248);
nand U1479 (N_1479,N_597,N_423);
or U1480 (N_1480,N_658,N_718);
and U1481 (N_1481,N_478,N_576);
xnor U1482 (N_1482,N_17,N_151);
nor U1483 (N_1483,N_205,N_29);
or U1484 (N_1484,N_707,N_992);
and U1485 (N_1485,N_655,N_900);
nand U1486 (N_1486,N_414,N_317);
and U1487 (N_1487,N_872,N_455);
nor U1488 (N_1488,N_570,N_888);
nor U1489 (N_1489,N_855,N_267);
nor U1490 (N_1490,N_553,N_680);
nor U1491 (N_1491,N_502,N_74);
nand U1492 (N_1492,N_63,N_651);
nand U1493 (N_1493,N_739,N_876);
or U1494 (N_1494,N_790,N_642);
and U1495 (N_1495,N_606,N_812);
nor U1496 (N_1496,N_432,N_19);
nand U1497 (N_1497,N_404,N_993);
nand U1498 (N_1498,N_494,N_334);
or U1499 (N_1499,N_417,N_616);
nand U1500 (N_1500,N_491,N_768);
or U1501 (N_1501,N_572,N_778);
and U1502 (N_1502,N_664,N_338);
nor U1503 (N_1503,N_591,N_573);
or U1504 (N_1504,N_196,N_468);
and U1505 (N_1505,N_752,N_744);
and U1506 (N_1506,N_48,N_954);
nand U1507 (N_1507,N_809,N_318);
nor U1508 (N_1508,N_187,N_972);
nor U1509 (N_1509,N_122,N_630);
or U1510 (N_1510,N_933,N_325);
and U1511 (N_1511,N_158,N_689);
or U1512 (N_1512,N_423,N_222);
or U1513 (N_1513,N_698,N_865);
and U1514 (N_1514,N_300,N_383);
and U1515 (N_1515,N_924,N_701);
or U1516 (N_1516,N_474,N_950);
or U1517 (N_1517,N_941,N_232);
nor U1518 (N_1518,N_369,N_205);
nor U1519 (N_1519,N_322,N_595);
nor U1520 (N_1520,N_392,N_835);
or U1521 (N_1521,N_275,N_942);
and U1522 (N_1522,N_696,N_288);
nand U1523 (N_1523,N_610,N_640);
nand U1524 (N_1524,N_569,N_598);
or U1525 (N_1525,N_83,N_440);
nand U1526 (N_1526,N_92,N_25);
nand U1527 (N_1527,N_521,N_577);
or U1528 (N_1528,N_566,N_812);
nand U1529 (N_1529,N_831,N_625);
nand U1530 (N_1530,N_493,N_848);
nand U1531 (N_1531,N_785,N_242);
nand U1532 (N_1532,N_384,N_643);
nand U1533 (N_1533,N_353,N_304);
or U1534 (N_1534,N_437,N_800);
and U1535 (N_1535,N_884,N_914);
nor U1536 (N_1536,N_699,N_8);
nand U1537 (N_1537,N_742,N_32);
nand U1538 (N_1538,N_340,N_515);
nor U1539 (N_1539,N_360,N_619);
and U1540 (N_1540,N_68,N_167);
nor U1541 (N_1541,N_352,N_327);
nand U1542 (N_1542,N_368,N_171);
nor U1543 (N_1543,N_665,N_680);
nand U1544 (N_1544,N_267,N_832);
and U1545 (N_1545,N_695,N_39);
and U1546 (N_1546,N_269,N_252);
or U1547 (N_1547,N_888,N_450);
and U1548 (N_1548,N_779,N_593);
or U1549 (N_1549,N_135,N_618);
nor U1550 (N_1550,N_693,N_884);
and U1551 (N_1551,N_166,N_280);
nand U1552 (N_1552,N_483,N_169);
nor U1553 (N_1553,N_297,N_723);
nand U1554 (N_1554,N_199,N_576);
nand U1555 (N_1555,N_34,N_464);
nand U1556 (N_1556,N_335,N_297);
nand U1557 (N_1557,N_133,N_530);
or U1558 (N_1558,N_643,N_767);
and U1559 (N_1559,N_983,N_535);
and U1560 (N_1560,N_87,N_820);
nor U1561 (N_1561,N_724,N_607);
or U1562 (N_1562,N_21,N_667);
and U1563 (N_1563,N_103,N_238);
nor U1564 (N_1564,N_31,N_230);
nand U1565 (N_1565,N_322,N_90);
and U1566 (N_1566,N_948,N_315);
nand U1567 (N_1567,N_479,N_597);
nor U1568 (N_1568,N_503,N_913);
or U1569 (N_1569,N_562,N_671);
or U1570 (N_1570,N_91,N_852);
nor U1571 (N_1571,N_391,N_827);
nand U1572 (N_1572,N_651,N_246);
xor U1573 (N_1573,N_386,N_264);
nor U1574 (N_1574,N_880,N_925);
and U1575 (N_1575,N_358,N_934);
and U1576 (N_1576,N_65,N_727);
nor U1577 (N_1577,N_123,N_91);
nand U1578 (N_1578,N_936,N_675);
or U1579 (N_1579,N_662,N_342);
nand U1580 (N_1580,N_467,N_894);
and U1581 (N_1581,N_691,N_79);
xor U1582 (N_1582,N_939,N_718);
xor U1583 (N_1583,N_312,N_294);
or U1584 (N_1584,N_305,N_784);
and U1585 (N_1585,N_331,N_969);
or U1586 (N_1586,N_965,N_781);
and U1587 (N_1587,N_525,N_610);
and U1588 (N_1588,N_868,N_446);
and U1589 (N_1589,N_785,N_63);
or U1590 (N_1590,N_729,N_199);
nor U1591 (N_1591,N_754,N_408);
and U1592 (N_1592,N_906,N_442);
and U1593 (N_1593,N_77,N_148);
nor U1594 (N_1594,N_557,N_46);
and U1595 (N_1595,N_872,N_599);
nor U1596 (N_1596,N_676,N_469);
nor U1597 (N_1597,N_156,N_132);
and U1598 (N_1598,N_847,N_175);
or U1599 (N_1599,N_836,N_662);
nor U1600 (N_1600,N_100,N_53);
nand U1601 (N_1601,N_988,N_558);
and U1602 (N_1602,N_77,N_584);
nor U1603 (N_1603,N_37,N_674);
nor U1604 (N_1604,N_301,N_756);
nand U1605 (N_1605,N_363,N_84);
nand U1606 (N_1606,N_173,N_637);
or U1607 (N_1607,N_888,N_115);
nor U1608 (N_1608,N_623,N_891);
or U1609 (N_1609,N_318,N_76);
nand U1610 (N_1610,N_384,N_435);
nor U1611 (N_1611,N_230,N_438);
nand U1612 (N_1612,N_455,N_376);
or U1613 (N_1613,N_230,N_237);
or U1614 (N_1614,N_143,N_970);
and U1615 (N_1615,N_692,N_52);
nand U1616 (N_1616,N_386,N_789);
and U1617 (N_1617,N_661,N_316);
or U1618 (N_1618,N_18,N_326);
and U1619 (N_1619,N_433,N_942);
or U1620 (N_1620,N_263,N_677);
nor U1621 (N_1621,N_879,N_52);
nand U1622 (N_1622,N_240,N_571);
nor U1623 (N_1623,N_270,N_596);
nand U1624 (N_1624,N_311,N_401);
nand U1625 (N_1625,N_945,N_213);
nand U1626 (N_1626,N_967,N_615);
or U1627 (N_1627,N_375,N_62);
nand U1628 (N_1628,N_542,N_455);
or U1629 (N_1629,N_888,N_59);
or U1630 (N_1630,N_544,N_209);
or U1631 (N_1631,N_280,N_829);
nor U1632 (N_1632,N_739,N_925);
nand U1633 (N_1633,N_291,N_227);
and U1634 (N_1634,N_213,N_412);
and U1635 (N_1635,N_617,N_654);
or U1636 (N_1636,N_743,N_988);
or U1637 (N_1637,N_761,N_104);
and U1638 (N_1638,N_967,N_447);
and U1639 (N_1639,N_748,N_636);
nand U1640 (N_1640,N_877,N_259);
nand U1641 (N_1641,N_534,N_600);
nand U1642 (N_1642,N_605,N_623);
and U1643 (N_1643,N_802,N_38);
nand U1644 (N_1644,N_468,N_481);
or U1645 (N_1645,N_677,N_748);
nor U1646 (N_1646,N_89,N_241);
or U1647 (N_1647,N_354,N_881);
or U1648 (N_1648,N_930,N_525);
xor U1649 (N_1649,N_85,N_739);
and U1650 (N_1650,N_703,N_926);
nand U1651 (N_1651,N_140,N_349);
nand U1652 (N_1652,N_41,N_666);
and U1653 (N_1653,N_55,N_742);
nor U1654 (N_1654,N_277,N_102);
and U1655 (N_1655,N_27,N_76);
nor U1656 (N_1656,N_901,N_568);
and U1657 (N_1657,N_594,N_238);
nor U1658 (N_1658,N_131,N_112);
or U1659 (N_1659,N_557,N_716);
or U1660 (N_1660,N_984,N_117);
or U1661 (N_1661,N_454,N_973);
or U1662 (N_1662,N_285,N_165);
or U1663 (N_1663,N_101,N_907);
and U1664 (N_1664,N_395,N_771);
or U1665 (N_1665,N_135,N_823);
nand U1666 (N_1666,N_803,N_505);
or U1667 (N_1667,N_897,N_493);
or U1668 (N_1668,N_499,N_353);
or U1669 (N_1669,N_524,N_375);
nand U1670 (N_1670,N_738,N_287);
or U1671 (N_1671,N_906,N_116);
nand U1672 (N_1672,N_681,N_675);
nand U1673 (N_1673,N_622,N_903);
or U1674 (N_1674,N_721,N_497);
and U1675 (N_1675,N_85,N_626);
and U1676 (N_1676,N_489,N_368);
nand U1677 (N_1677,N_453,N_330);
nor U1678 (N_1678,N_739,N_742);
nand U1679 (N_1679,N_801,N_241);
nor U1680 (N_1680,N_462,N_534);
nand U1681 (N_1681,N_300,N_725);
and U1682 (N_1682,N_265,N_896);
nor U1683 (N_1683,N_406,N_417);
nand U1684 (N_1684,N_638,N_524);
and U1685 (N_1685,N_537,N_761);
nand U1686 (N_1686,N_674,N_323);
nand U1687 (N_1687,N_781,N_678);
nand U1688 (N_1688,N_311,N_588);
and U1689 (N_1689,N_734,N_661);
nand U1690 (N_1690,N_8,N_615);
nand U1691 (N_1691,N_104,N_495);
and U1692 (N_1692,N_154,N_120);
nand U1693 (N_1693,N_365,N_203);
and U1694 (N_1694,N_678,N_72);
nor U1695 (N_1695,N_811,N_726);
nand U1696 (N_1696,N_240,N_499);
and U1697 (N_1697,N_681,N_114);
and U1698 (N_1698,N_602,N_186);
or U1699 (N_1699,N_359,N_59);
and U1700 (N_1700,N_599,N_509);
or U1701 (N_1701,N_780,N_283);
and U1702 (N_1702,N_97,N_597);
nand U1703 (N_1703,N_987,N_570);
and U1704 (N_1704,N_205,N_265);
nand U1705 (N_1705,N_60,N_782);
nor U1706 (N_1706,N_332,N_397);
nand U1707 (N_1707,N_392,N_148);
nor U1708 (N_1708,N_138,N_928);
nand U1709 (N_1709,N_682,N_51);
or U1710 (N_1710,N_60,N_590);
nand U1711 (N_1711,N_700,N_152);
and U1712 (N_1712,N_835,N_209);
nor U1713 (N_1713,N_580,N_386);
or U1714 (N_1714,N_229,N_10);
and U1715 (N_1715,N_18,N_922);
and U1716 (N_1716,N_746,N_968);
or U1717 (N_1717,N_501,N_615);
or U1718 (N_1718,N_628,N_652);
or U1719 (N_1719,N_385,N_284);
nor U1720 (N_1720,N_686,N_773);
nor U1721 (N_1721,N_56,N_679);
nor U1722 (N_1722,N_190,N_788);
and U1723 (N_1723,N_435,N_178);
or U1724 (N_1724,N_948,N_484);
nor U1725 (N_1725,N_838,N_297);
or U1726 (N_1726,N_290,N_106);
or U1727 (N_1727,N_709,N_185);
nor U1728 (N_1728,N_533,N_495);
or U1729 (N_1729,N_463,N_682);
and U1730 (N_1730,N_989,N_201);
or U1731 (N_1731,N_438,N_304);
nand U1732 (N_1732,N_849,N_315);
nand U1733 (N_1733,N_67,N_169);
nand U1734 (N_1734,N_471,N_271);
nor U1735 (N_1735,N_54,N_770);
or U1736 (N_1736,N_784,N_145);
nor U1737 (N_1737,N_148,N_347);
nand U1738 (N_1738,N_517,N_615);
and U1739 (N_1739,N_282,N_408);
or U1740 (N_1740,N_45,N_780);
nor U1741 (N_1741,N_177,N_538);
nor U1742 (N_1742,N_331,N_570);
or U1743 (N_1743,N_910,N_352);
nor U1744 (N_1744,N_144,N_503);
nand U1745 (N_1745,N_479,N_62);
or U1746 (N_1746,N_667,N_306);
or U1747 (N_1747,N_893,N_618);
nor U1748 (N_1748,N_631,N_101);
nand U1749 (N_1749,N_605,N_707);
nand U1750 (N_1750,N_863,N_567);
nand U1751 (N_1751,N_101,N_197);
nand U1752 (N_1752,N_102,N_963);
and U1753 (N_1753,N_540,N_776);
or U1754 (N_1754,N_33,N_896);
or U1755 (N_1755,N_856,N_384);
or U1756 (N_1756,N_9,N_971);
nor U1757 (N_1757,N_471,N_549);
nor U1758 (N_1758,N_127,N_971);
and U1759 (N_1759,N_922,N_196);
nand U1760 (N_1760,N_151,N_334);
and U1761 (N_1761,N_797,N_328);
or U1762 (N_1762,N_17,N_449);
or U1763 (N_1763,N_983,N_97);
and U1764 (N_1764,N_6,N_31);
or U1765 (N_1765,N_12,N_584);
nand U1766 (N_1766,N_448,N_649);
nor U1767 (N_1767,N_332,N_500);
nand U1768 (N_1768,N_946,N_42);
or U1769 (N_1769,N_625,N_316);
or U1770 (N_1770,N_736,N_55);
or U1771 (N_1771,N_953,N_291);
xnor U1772 (N_1772,N_956,N_657);
or U1773 (N_1773,N_836,N_888);
nand U1774 (N_1774,N_633,N_961);
and U1775 (N_1775,N_750,N_773);
nor U1776 (N_1776,N_238,N_983);
and U1777 (N_1777,N_618,N_753);
nor U1778 (N_1778,N_216,N_822);
or U1779 (N_1779,N_566,N_117);
or U1780 (N_1780,N_488,N_849);
xor U1781 (N_1781,N_185,N_17);
or U1782 (N_1782,N_283,N_239);
and U1783 (N_1783,N_782,N_407);
or U1784 (N_1784,N_363,N_748);
xor U1785 (N_1785,N_347,N_134);
nand U1786 (N_1786,N_837,N_994);
nand U1787 (N_1787,N_724,N_637);
nand U1788 (N_1788,N_298,N_481);
nor U1789 (N_1789,N_751,N_3);
and U1790 (N_1790,N_1,N_800);
nor U1791 (N_1791,N_647,N_826);
nand U1792 (N_1792,N_198,N_558);
nor U1793 (N_1793,N_455,N_215);
nand U1794 (N_1794,N_802,N_54);
or U1795 (N_1795,N_653,N_528);
and U1796 (N_1796,N_963,N_468);
xor U1797 (N_1797,N_892,N_461);
and U1798 (N_1798,N_591,N_391);
or U1799 (N_1799,N_908,N_943);
nand U1800 (N_1800,N_561,N_256);
and U1801 (N_1801,N_564,N_525);
and U1802 (N_1802,N_546,N_27);
and U1803 (N_1803,N_599,N_269);
nand U1804 (N_1804,N_166,N_405);
or U1805 (N_1805,N_666,N_139);
and U1806 (N_1806,N_280,N_685);
nor U1807 (N_1807,N_191,N_152);
or U1808 (N_1808,N_417,N_12);
nand U1809 (N_1809,N_936,N_815);
nand U1810 (N_1810,N_855,N_71);
and U1811 (N_1811,N_102,N_187);
nor U1812 (N_1812,N_406,N_851);
nor U1813 (N_1813,N_796,N_927);
xnor U1814 (N_1814,N_82,N_830);
nand U1815 (N_1815,N_515,N_509);
nand U1816 (N_1816,N_269,N_373);
nor U1817 (N_1817,N_948,N_614);
nand U1818 (N_1818,N_975,N_63);
nor U1819 (N_1819,N_389,N_170);
nor U1820 (N_1820,N_389,N_680);
and U1821 (N_1821,N_836,N_711);
and U1822 (N_1822,N_707,N_701);
nand U1823 (N_1823,N_398,N_420);
nand U1824 (N_1824,N_483,N_929);
or U1825 (N_1825,N_87,N_57);
and U1826 (N_1826,N_150,N_335);
nor U1827 (N_1827,N_739,N_423);
nor U1828 (N_1828,N_744,N_300);
nand U1829 (N_1829,N_647,N_618);
and U1830 (N_1830,N_786,N_282);
or U1831 (N_1831,N_727,N_346);
nand U1832 (N_1832,N_142,N_538);
and U1833 (N_1833,N_931,N_481);
and U1834 (N_1834,N_707,N_251);
or U1835 (N_1835,N_489,N_785);
and U1836 (N_1836,N_583,N_388);
nor U1837 (N_1837,N_411,N_174);
and U1838 (N_1838,N_60,N_740);
nand U1839 (N_1839,N_584,N_563);
xor U1840 (N_1840,N_858,N_534);
nor U1841 (N_1841,N_421,N_242);
nand U1842 (N_1842,N_786,N_739);
nor U1843 (N_1843,N_215,N_269);
and U1844 (N_1844,N_140,N_603);
and U1845 (N_1845,N_656,N_435);
or U1846 (N_1846,N_941,N_547);
nor U1847 (N_1847,N_66,N_903);
and U1848 (N_1848,N_911,N_951);
or U1849 (N_1849,N_659,N_259);
or U1850 (N_1850,N_786,N_491);
and U1851 (N_1851,N_830,N_118);
and U1852 (N_1852,N_759,N_401);
and U1853 (N_1853,N_310,N_291);
or U1854 (N_1854,N_288,N_583);
and U1855 (N_1855,N_485,N_955);
nand U1856 (N_1856,N_23,N_294);
or U1857 (N_1857,N_195,N_236);
or U1858 (N_1858,N_825,N_556);
and U1859 (N_1859,N_671,N_399);
or U1860 (N_1860,N_19,N_853);
or U1861 (N_1861,N_160,N_561);
nor U1862 (N_1862,N_347,N_399);
and U1863 (N_1863,N_224,N_363);
or U1864 (N_1864,N_643,N_130);
nand U1865 (N_1865,N_910,N_814);
or U1866 (N_1866,N_85,N_986);
or U1867 (N_1867,N_454,N_824);
or U1868 (N_1868,N_78,N_672);
and U1869 (N_1869,N_630,N_895);
nor U1870 (N_1870,N_434,N_756);
nand U1871 (N_1871,N_323,N_911);
nor U1872 (N_1872,N_758,N_15);
nor U1873 (N_1873,N_3,N_783);
nor U1874 (N_1874,N_743,N_676);
or U1875 (N_1875,N_54,N_929);
nand U1876 (N_1876,N_663,N_843);
or U1877 (N_1877,N_633,N_510);
and U1878 (N_1878,N_632,N_385);
nand U1879 (N_1879,N_146,N_936);
or U1880 (N_1880,N_37,N_394);
and U1881 (N_1881,N_96,N_754);
nand U1882 (N_1882,N_919,N_637);
or U1883 (N_1883,N_270,N_700);
and U1884 (N_1884,N_408,N_726);
or U1885 (N_1885,N_725,N_736);
and U1886 (N_1886,N_472,N_591);
nand U1887 (N_1887,N_620,N_617);
or U1888 (N_1888,N_195,N_635);
or U1889 (N_1889,N_470,N_873);
nor U1890 (N_1890,N_994,N_9);
and U1891 (N_1891,N_855,N_712);
nand U1892 (N_1892,N_27,N_375);
nand U1893 (N_1893,N_451,N_351);
nor U1894 (N_1894,N_537,N_609);
nor U1895 (N_1895,N_213,N_603);
and U1896 (N_1896,N_892,N_982);
nor U1897 (N_1897,N_89,N_182);
and U1898 (N_1898,N_417,N_492);
or U1899 (N_1899,N_753,N_838);
or U1900 (N_1900,N_40,N_640);
and U1901 (N_1901,N_312,N_72);
or U1902 (N_1902,N_898,N_712);
and U1903 (N_1903,N_483,N_122);
nand U1904 (N_1904,N_360,N_572);
or U1905 (N_1905,N_247,N_350);
or U1906 (N_1906,N_695,N_518);
and U1907 (N_1907,N_217,N_964);
and U1908 (N_1908,N_118,N_745);
or U1909 (N_1909,N_197,N_587);
nand U1910 (N_1910,N_349,N_638);
nor U1911 (N_1911,N_929,N_757);
xor U1912 (N_1912,N_306,N_705);
nand U1913 (N_1913,N_686,N_165);
nand U1914 (N_1914,N_205,N_734);
nand U1915 (N_1915,N_56,N_982);
nor U1916 (N_1916,N_735,N_716);
or U1917 (N_1917,N_822,N_858);
and U1918 (N_1918,N_248,N_415);
nand U1919 (N_1919,N_261,N_462);
or U1920 (N_1920,N_630,N_102);
and U1921 (N_1921,N_233,N_198);
and U1922 (N_1922,N_934,N_893);
or U1923 (N_1923,N_201,N_416);
or U1924 (N_1924,N_439,N_34);
or U1925 (N_1925,N_614,N_481);
and U1926 (N_1926,N_32,N_71);
nand U1927 (N_1927,N_579,N_17);
or U1928 (N_1928,N_942,N_809);
nand U1929 (N_1929,N_770,N_232);
and U1930 (N_1930,N_865,N_550);
and U1931 (N_1931,N_782,N_839);
or U1932 (N_1932,N_584,N_532);
and U1933 (N_1933,N_471,N_895);
nand U1934 (N_1934,N_820,N_672);
or U1935 (N_1935,N_567,N_187);
nand U1936 (N_1936,N_93,N_416);
and U1937 (N_1937,N_590,N_378);
or U1938 (N_1938,N_653,N_57);
nor U1939 (N_1939,N_987,N_699);
or U1940 (N_1940,N_952,N_12);
or U1941 (N_1941,N_862,N_596);
and U1942 (N_1942,N_137,N_392);
and U1943 (N_1943,N_418,N_178);
nor U1944 (N_1944,N_985,N_560);
and U1945 (N_1945,N_658,N_937);
nor U1946 (N_1946,N_347,N_860);
or U1947 (N_1947,N_255,N_250);
or U1948 (N_1948,N_264,N_927);
nand U1949 (N_1949,N_399,N_539);
or U1950 (N_1950,N_394,N_31);
or U1951 (N_1951,N_420,N_467);
nor U1952 (N_1952,N_822,N_380);
and U1953 (N_1953,N_558,N_944);
nand U1954 (N_1954,N_185,N_998);
or U1955 (N_1955,N_830,N_231);
and U1956 (N_1956,N_682,N_143);
and U1957 (N_1957,N_753,N_874);
or U1958 (N_1958,N_399,N_262);
nor U1959 (N_1959,N_364,N_958);
or U1960 (N_1960,N_328,N_593);
nor U1961 (N_1961,N_318,N_514);
or U1962 (N_1962,N_825,N_88);
or U1963 (N_1963,N_612,N_255);
nand U1964 (N_1964,N_452,N_569);
nand U1965 (N_1965,N_438,N_523);
or U1966 (N_1966,N_500,N_263);
or U1967 (N_1967,N_312,N_282);
and U1968 (N_1968,N_718,N_271);
nand U1969 (N_1969,N_533,N_389);
and U1970 (N_1970,N_999,N_910);
nor U1971 (N_1971,N_464,N_799);
nor U1972 (N_1972,N_51,N_476);
or U1973 (N_1973,N_679,N_50);
and U1974 (N_1974,N_853,N_36);
and U1975 (N_1975,N_559,N_677);
nor U1976 (N_1976,N_400,N_558);
or U1977 (N_1977,N_153,N_875);
or U1978 (N_1978,N_948,N_748);
nor U1979 (N_1979,N_93,N_598);
or U1980 (N_1980,N_369,N_21);
nand U1981 (N_1981,N_995,N_657);
or U1982 (N_1982,N_279,N_49);
and U1983 (N_1983,N_42,N_736);
or U1984 (N_1984,N_836,N_944);
or U1985 (N_1985,N_536,N_958);
nor U1986 (N_1986,N_746,N_946);
nand U1987 (N_1987,N_901,N_602);
and U1988 (N_1988,N_443,N_208);
nand U1989 (N_1989,N_966,N_953);
or U1990 (N_1990,N_320,N_521);
and U1991 (N_1991,N_53,N_451);
or U1992 (N_1992,N_170,N_667);
nor U1993 (N_1993,N_760,N_583);
and U1994 (N_1994,N_290,N_852);
nand U1995 (N_1995,N_626,N_518);
nor U1996 (N_1996,N_325,N_334);
nor U1997 (N_1997,N_193,N_826);
nand U1998 (N_1998,N_912,N_130);
or U1999 (N_1999,N_240,N_299);
and U2000 (N_2000,N_1198,N_1671);
nand U2001 (N_2001,N_1697,N_1229);
nor U2002 (N_2002,N_1819,N_1402);
or U2003 (N_2003,N_1812,N_1661);
and U2004 (N_2004,N_1392,N_1056);
nand U2005 (N_2005,N_1635,N_1658);
nor U2006 (N_2006,N_1904,N_1901);
or U2007 (N_2007,N_1617,N_1099);
and U2008 (N_2008,N_1467,N_1379);
and U2009 (N_2009,N_1835,N_1592);
nand U2010 (N_2010,N_1169,N_1751);
nor U2011 (N_2011,N_1763,N_1417);
and U2012 (N_2012,N_1456,N_1998);
nor U2013 (N_2013,N_1519,N_1807);
nand U2014 (N_2014,N_1016,N_1919);
nor U2015 (N_2015,N_1026,N_1504);
or U2016 (N_2016,N_1106,N_1712);
nand U2017 (N_2017,N_1801,N_1937);
nand U2018 (N_2018,N_1983,N_1348);
nand U2019 (N_2019,N_1657,N_1047);
nor U2020 (N_2020,N_1777,N_1875);
or U2021 (N_2021,N_1311,N_1072);
nor U2022 (N_2022,N_1925,N_1693);
and U2023 (N_2023,N_1742,N_1286);
nand U2024 (N_2024,N_1676,N_1060);
nand U2025 (N_2025,N_1158,N_1084);
nor U2026 (N_2026,N_1190,N_1911);
and U2027 (N_2027,N_1384,N_1791);
and U2028 (N_2028,N_1055,N_1065);
or U2029 (N_2029,N_1376,N_1769);
or U2030 (N_2030,N_1023,N_1648);
nand U2031 (N_2031,N_1424,N_1173);
nor U2032 (N_2032,N_1955,N_1864);
nand U2033 (N_2033,N_1339,N_1464);
nor U2034 (N_2034,N_1351,N_1009);
nor U2035 (N_2035,N_1122,N_1381);
and U2036 (N_2036,N_1189,N_1045);
nor U2037 (N_2037,N_1057,N_1269);
nor U2038 (N_2038,N_1775,N_1849);
nor U2039 (N_2039,N_1560,N_1618);
nor U2040 (N_2040,N_1188,N_1843);
or U2041 (N_2041,N_1015,N_1191);
and U2042 (N_2042,N_1215,N_1971);
nor U2043 (N_2043,N_1921,N_1789);
nand U2044 (N_2044,N_1880,N_1404);
nor U2045 (N_2045,N_1207,N_1529);
nor U2046 (N_2046,N_1884,N_1073);
and U2047 (N_2047,N_1991,N_1887);
or U2048 (N_2048,N_1956,N_1263);
nor U2049 (N_2049,N_1561,N_1347);
and U2050 (N_2050,N_1380,N_1494);
nor U2051 (N_2051,N_1407,N_1272);
or U2052 (N_2052,N_1240,N_1248);
or U2053 (N_2053,N_1876,N_1227);
or U2054 (N_2054,N_1214,N_1757);
or U2055 (N_2055,N_1936,N_1588);
nor U2056 (N_2056,N_1509,N_1116);
or U2057 (N_2057,N_1995,N_1946);
nand U2058 (N_2058,N_1639,N_1331);
nor U2059 (N_2059,N_1346,N_1458);
nor U2060 (N_2060,N_1759,N_1896);
or U2061 (N_2061,N_1054,N_1942);
nand U2062 (N_2062,N_1194,N_1077);
or U2063 (N_2063,N_1493,N_1014);
and U2064 (N_2064,N_1707,N_1206);
or U2065 (N_2065,N_1010,N_1360);
and U2066 (N_2066,N_1343,N_1480);
nand U2067 (N_2067,N_1913,N_1965);
and U2068 (N_2068,N_1502,N_1498);
nand U2069 (N_2069,N_1727,N_1290);
and U2070 (N_2070,N_1159,N_1933);
nand U2071 (N_2071,N_1692,N_1893);
nand U2072 (N_2072,N_1196,N_1069);
or U2073 (N_2073,N_1792,N_1950);
and U2074 (N_2074,N_1636,N_1974);
or U2075 (N_2075,N_1987,N_1066);
or U2076 (N_2076,N_1308,N_1886);
and U2077 (N_2077,N_1581,N_1938);
nor U2078 (N_2078,N_1916,N_1665);
nand U2079 (N_2079,N_1150,N_1575);
nor U2080 (N_2080,N_1545,N_1660);
or U2081 (N_2081,N_1681,N_1164);
and U2082 (N_2082,N_1328,N_1293);
and U2083 (N_2083,N_1868,N_1619);
nor U2084 (N_2084,N_1332,N_1976);
nor U2085 (N_2085,N_1341,N_1973);
nor U2086 (N_2086,N_1963,N_1064);
nand U2087 (N_2087,N_1964,N_1850);
nand U2088 (N_2088,N_1885,N_1684);
or U2089 (N_2089,N_1267,N_1059);
or U2090 (N_2090,N_1689,N_1553);
nand U2091 (N_2091,N_1770,N_1966);
nand U2092 (N_2092,N_1317,N_1972);
or U2093 (N_2093,N_1805,N_1871);
nand U2094 (N_2094,N_1912,N_1472);
nor U2095 (N_2095,N_1414,N_1860);
and U2096 (N_2096,N_1102,N_1113);
nor U2097 (N_2097,N_1434,N_1699);
nand U2098 (N_2098,N_1209,N_1626);
and U2099 (N_2099,N_1570,N_1898);
nor U2100 (N_2100,N_1910,N_1143);
nor U2101 (N_2101,N_1683,N_1601);
nand U2102 (N_2102,N_1841,N_1517);
or U2103 (N_2103,N_1748,N_1556);
nor U2104 (N_2104,N_1675,N_1283);
and U2105 (N_2105,N_1590,N_1802);
nand U2106 (N_2106,N_1643,N_1631);
nand U2107 (N_2107,N_1304,N_1908);
nand U2108 (N_2108,N_1285,N_1291);
or U2109 (N_2109,N_1958,N_1129);
nor U2110 (N_2110,N_1257,N_1473);
and U2111 (N_2111,N_1825,N_1366);
nor U2112 (N_2112,N_1305,N_1945);
or U2113 (N_2113,N_1422,N_1216);
or U2114 (N_2114,N_1610,N_1603);
nor U2115 (N_2115,N_1823,N_1217);
or U2116 (N_2116,N_1273,N_1221);
and U2117 (N_2117,N_1301,N_1829);
or U2118 (N_2118,N_1444,N_1922);
nor U2119 (N_2119,N_1852,N_1249);
nand U2120 (N_2120,N_1428,N_1337);
nand U2121 (N_2121,N_1262,N_1359);
nor U2122 (N_2122,N_1186,N_1320);
or U2123 (N_2123,N_1008,N_1572);
nand U2124 (N_2124,N_1862,N_1039);
and U2125 (N_2125,N_1142,N_1438);
and U2126 (N_2126,N_1951,N_1605);
xnor U2127 (N_2127,N_1416,N_1231);
or U2128 (N_2128,N_1947,N_1764);
or U2129 (N_2129,N_1342,N_1389);
and U2130 (N_2130,N_1754,N_1596);
nor U2131 (N_2131,N_1546,N_1753);
and U2132 (N_2132,N_1834,N_1411);
nand U2133 (N_2133,N_1507,N_1451);
or U2134 (N_2134,N_1799,N_1760);
nor U2135 (N_2135,N_1755,N_1388);
or U2136 (N_2136,N_1678,N_1637);
xor U2137 (N_2137,N_1461,N_1774);
nor U2138 (N_2138,N_1996,N_1481);
and U2139 (N_2139,N_1048,N_1356);
nand U2140 (N_2140,N_1729,N_1932);
or U2141 (N_2141,N_1446,N_1485);
and U2142 (N_2142,N_1747,N_1032);
and U2143 (N_2143,N_1824,N_1121);
nor U2144 (N_2144,N_1688,N_1490);
nand U2145 (N_2145,N_1147,N_1361);
nand U2146 (N_2146,N_1097,N_1583);
or U2147 (N_2147,N_1130,N_1846);
nand U2148 (N_2148,N_1704,N_1036);
and U2149 (N_2149,N_1365,N_1894);
nor U2150 (N_2150,N_1604,N_1144);
or U2151 (N_2151,N_1117,N_1653);
nor U2152 (N_2152,N_1810,N_1396);
nand U2153 (N_2153,N_1100,N_1149);
and U2154 (N_2154,N_1827,N_1953);
and U2155 (N_2155,N_1557,N_1355);
and U2156 (N_2156,N_1322,N_1132);
and U2157 (N_2157,N_1833,N_1203);
or U2158 (N_2158,N_1294,N_1644);
nor U2159 (N_2159,N_1749,N_1243);
or U2160 (N_2160,N_1061,N_1836);
nand U2161 (N_2161,N_1666,N_1436);
nand U2162 (N_2162,N_1703,N_1872);
or U2163 (N_2163,N_1078,N_1330);
or U2164 (N_2164,N_1195,N_1881);
and U2165 (N_2165,N_1315,N_1104);
or U2166 (N_2166,N_1528,N_1087);
nor U2167 (N_2167,N_1977,N_1027);
nor U2168 (N_2168,N_1784,N_1479);
nand U2169 (N_2169,N_1726,N_1210);
or U2170 (N_2170,N_1020,N_1353);
nand U2171 (N_2171,N_1238,N_1698);
nor U2172 (N_2172,N_1584,N_1620);
or U2173 (N_2173,N_1606,N_1177);
or U2174 (N_2174,N_1281,N_1165);
and U2175 (N_2175,N_1597,N_1335);
or U2176 (N_2176,N_1505,N_1489);
or U2177 (N_2177,N_1544,N_1591);
or U2178 (N_2178,N_1524,N_1861);
nand U2179 (N_2179,N_1741,N_1401);
nand U2180 (N_2180,N_1969,N_1928);
and U2181 (N_2181,N_1818,N_1705);
nand U2182 (N_2182,N_1838,N_1765);
nand U2183 (N_2183,N_1303,N_1718);
nand U2184 (N_2184,N_1041,N_1255);
nand U2185 (N_2185,N_1338,N_1562);
and U2186 (N_2186,N_1719,N_1029);
nand U2187 (N_2187,N_1773,N_1168);
and U2188 (N_2188,N_1200,N_1017);
nand U2189 (N_2189,N_1171,N_1419);
nor U2190 (N_2190,N_1462,N_1484);
nand U2191 (N_2191,N_1776,N_1199);
nand U2192 (N_2192,N_1649,N_1814);
or U2193 (N_2193,N_1559,N_1432);
nand U2194 (N_2194,N_1135,N_1090);
nand U2195 (N_2195,N_1003,N_1939);
nand U2196 (N_2196,N_1278,N_1975);
and U2197 (N_2197,N_1152,N_1882);
nor U2198 (N_2198,N_1319,N_1133);
and U2199 (N_2199,N_1264,N_1270);
or U2200 (N_2200,N_1670,N_1120);
or U2201 (N_2201,N_1526,N_1358);
nor U2202 (N_2202,N_1465,N_1442);
nand U2203 (N_2203,N_1161,N_1344);
and U2204 (N_2204,N_1970,N_1700);
nor U2205 (N_2205,N_1865,N_1107);
and U2206 (N_2206,N_1378,N_1992);
nor U2207 (N_2207,N_1382,N_1028);
nor U2208 (N_2208,N_1336,N_1074);
and U2209 (N_2209,N_1582,N_1426);
and U2210 (N_2210,N_1420,N_1923);
nor U2211 (N_2211,N_1326,N_1092);
nor U2212 (N_2212,N_1779,N_1540);
or U2213 (N_2213,N_1146,N_1433);
nor U2214 (N_2214,N_1793,N_1654);
nand U2215 (N_2215,N_1098,N_1744);
nand U2216 (N_2216,N_1141,N_1192);
and U2217 (N_2217,N_1312,N_1873);
or U2218 (N_2218,N_1445,N_1598);
and U2219 (N_2219,N_1226,N_1611);
nand U2220 (N_2220,N_1225,N_1869);
nand U2221 (N_2221,N_1762,N_1298);
or U2222 (N_2222,N_1443,N_1800);
nand U2223 (N_2223,N_1181,N_1521);
or U2224 (N_2224,N_1892,N_1174);
or U2225 (N_2225,N_1794,N_1131);
or U2226 (N_2226,N_1002,N_1112);
and U2227 (N_2227,N_1323,N_1577);
nor U2228 (N_2228,N_1275,N_1614);
nor U2229 (N_2229,N_1780,N_1448);
xnor U2230 (N_2230,N_1709,N_1329);
nand U2231 (N_2231,N_1542,N_1449);
nor U2232 (N_2232,N_1300,N_1806);
and U2233 (N_2233,N_1492,N_1115);
and U2234 (N_2234,N_1235,N_1390);
nand U2235 (N_2235,N_1567,N_1903);
and U2236 (N_2236,N_1728,N_1948);
nand U2237 (N_2237,N_1701,N_1364);
nand U2238 (N_2238,N_1687,N_1239);
nor U2239 (N_2239,N_1085,N_1926);
nand U2240 (N_2240,N_1576,N_1909);
or U2241 (N_2241,N_1418,N_1766);
nor U2242 (N_2242,N_1333,N_1080);
and U2243 (N_2243,N_1471,N_1035);
nand U2244 (N_2244,N_1110,N_1522);
nor U2245 (N_2245,N_1108,N_1713);
nor U2246 (N_2246,N_1091,N_1616);
nor U2247 (N_2247,N_1732,N_1645);
nor U2248 (N_2248,N_1883,N_1512);
xor U2249 (N_2249,N_1979,N_1790);
nor U2250 (N_2250,N_1525,N_1430);
nand U2251 (N_2251,N_1552,N_1310);
and U2252 (N_2252,N_1599,N_1877);
nand U2253 (N_2253,N_1822,N_1350);
and U2254 (N_2254,N_1224,N_1625);
and U2255 (N_2255,N_1393,N_1959);
or U2256 (N_2256,N_1372,N_1463);
nor U2257 (N_2257,N_1111,N_1566);
and U2258 (N_2258,N_1879,N_1482);
or U2259 (N_2259,N_1514,N_1564);
nand U2260 (N_2260,N_1737,N_1721);
and U2261 (N_2261,N_1523,N_1981);
nor U2262 (N_2262,N_1813,N_1568);
or U2263 (N_2263,N_1863,N_1673);
or U2264 (N_2264,N_1716,N_1984);
and U2265 (N_2265,N_1752,N_1232);
and U2266 (N_2266,N_1949,N_1474);
nor U2267 (N_2267,N_1828,N_1413);
or U2268 (N_2268,N_1000,N_1425);
or U2269 (N_2269,N_1044,N_1781);
nand U2270 (N_2270,N_1006,N_1837);
nor U2271 (N_2271,N_1313,N_1578);
nor U2272 (N_2272,N_1621,N_1175);
nor U2273 (N_2273,N_1415,N_1710);
nand U2274 (N_2274,N_1851,N_1105);
or U2275 (N_2275,N_1409,N_1600);
or U2276 (N_2276,N_1720,N_1798);
or U2277 (N_2277,N_1722,N_1857);
and U2278 (N_2278,N_1265,N_1237);
nand U2279 (N_2279,N_1162,N_1859);
nor U2280 (N_2280,N_1024,N_1076);
and U2281 (N_2281,N_1746,N_1202);
nor U2282 (N_2282,N_1993,N_1724);
or U2283 (N_2283,N_1031,N_1153);
or U2284 (N_2284,N_1037,N_1109);
nand U2285 (N_2285,N_1486,N_1797);
nand U2286 (N_2286,N_1758,N_1826);
nor U2287 (N_2287,N_1539,N_1651);
nor U2288 (N_2288,N_1367,N_1460);
nor U2289 (N_2289,N_1212,N_1469);
nand U2290 (N_2290,N_1624,N_1640);
nor U2291 (N_2291,N_1750,N_1292);
or U2292 (N_2292,N_1241,N_1371);
nor U2293 (N_2293,N_1589,N_1516);
nor U2294 (N_2294,N_1831,N_1488);
nor U2295 (N_2295,N_1391,N_1907);
nor U2296 (N_2296,N_1470,N_1230);
nand U2297 (N_2297,N_1483,N_1941);
or U2298 (N_2298,N_1520,N_1515);
and U2299 (N_2299,N_1848,N_1441);
and U2300 (N_2300,N_1609,N_1193);
and U2301 (N_2301,N_1134,N_1437);
nor U2302 (N_2302,N_1094,N_1145);
nand U2303 (N_2303,N_1088,N_1487);
and U2304 (N_2304,N_1325,N_1647);
nand U2305 (N_2305,N_1034,N_1408);
nand U2306 (N_2306,N_1623,N_1260);
or U2307 (N_2307,N_1538,N_1137);
nor U2308 (N_2308,N_1496,N_1821);
or U2309 (N_2309,N_1258,N_1050);
and U2310 (N_2310,N_1927,N_1246);
nor U2311 (N_2311,N_1287,N_1089);
nor U2312 (N_2312,N_1447,N_1354);
and U2313 (N_2313,N_1276,N_1247);
nor U2314 (N_2314,N_1554,N_1782);
or U2315 (N_2315,N_1030,N_1733);
nor U2316 (N_2316,N_1124,N_1254);
nor U2317 (N_2317,N_1767,N_1917);
and U2318 (N_2318,N_1691,N_1259);
nand U2319 (N_2319,N_1180,N_1204);
nand U2320 (N_2320,N_1920,N_1659);
and U2321 (N_2321,N_1250,N_1935);
or U2322 (N_2322,N_1271,N_1594);
and U2323 (N_2323,N_1565,N_1082);
nor U2324 (N_2324,N_1368,N_1761);
nor U2325 (N_2325,N_1058,N_1563);
and U2326 (N_2326,N_1682,N_1261);
nand U2327 (N_2327,N_1148,N_1155);
nor U2328 (N_2328,N_1399,N_1004);
xor U2329 (N_2329,N_1918,N_1160);
and U2330 (N_2330,N_1874,N_1569);
xnor U2331 (N_2331,N_1178,N_1674);
or U2332 (N_2332,N_1151,N_1213);
nor U2333 (N_2333,N_1547,N_1233);
and U2334 (N_2334,N_1400,N_1398);
and U2335 (N_2335,N_1655,N_1067);
nor U2336 (N_2336,N_1176,N_1468);
or U2337 (N_2337,N_1672,N_1550);
nand U2338 (N_2338,N_1349,N_1052);
and U2339 (N_2339,N_1988,N_1081);
nand U2340 (N_2340,N_1280,N_1220);
or U2341 (N_2341,N_1961,N_1531);
and U2342 (N_2342,N_1593,N_1585);
or U2343 (N_2343,N_1503,N_1680);
nor U2344 (N_2344,N_1967,N_1982);
or U2345 (N_2345,N_1394,N_1633);
and U2346 (N_2346,N_1499,N_1185);
nor U2347 (N_2347,N_1579,N_1439);
nor U2348 (N_2348,N_1466,N_1602);
nand U2349 (N_2349,N_1495,N_1702);
xor U2350 (N_2350,N_1043,N_1452);
nor U2351 (N_2351,N_1905,N_1622);
nor U2352 (N_2352,N_1357,N_1297);
nor U2353 (N_2353,N_1943,N_1352);
nor U2354 (N_2354,N_1299,N_1731);
or U2355 (N_2355,N_1435,N_1870);
or U2356 (N_2356,N_1652,N_1989);
or U2357 (N_2357,N_1978,N_1808);
or U2358 (N_2358,N_1811,N_1501);
nor U2359 (N_2359,N_1855,N_1628);
or U2360 (N_2360,N_1478,N_1431);
nor U2361 (N_2361,N_1662,N_1295);
nor U2362 (N_2362,N_1395,N_1075);
nand U2363 (N_2363,N_1960,N_1457);
and U2364 (N_2364,N_1236,N_1321);
and U2365 (N_2365,N_1796,N_1866);
nor U2366 (N_2366,N_1251,N_1128);
and U2367 (N_2367,N_1114,N_1079);
nand U2368 (N_2368,N_1980,N_1500);
and U2369 (N_2369,N_1208,N_1840);
or U2370 (N_2370,N_1685,N_1156);
or U2371 (N_2371,N_1815,N_1429);
or U2372 (N_2372,N_1634,N_1314);
and U2373 (N_2373,N_1891,N_1318);
nor U2374 (N_2374,N_1696,N_1093);
nor U2375 (N_2375,N_1668,N_1914);
nor U2376 (N_2376,N_1070,N_1005);
or U2377 (N_2377,N_1558,N_1218);
nand U2378 (N_2378,N_1316,N_1062);
nor U2379 (N_2379,N_1664,N_1809);
or U2380 (N_2380,N_1571,N_1387);
nor U2381 (N_2381,N_1453,N_1853);
nand U2382 (N_2382,N_1686,N_1650);
nand U2383 (N_2383,N_1656,N_1289);
and U2384 (N_2384,N_1049,N_1739);
nand U2385 (N_2385,N_1715,N_1786);
nand U2386 (N_2386,N_1535,N_1944);
nor U2387 (N_2387,N_1842,N_1440);
nor U2388 (N_2388,N_1580,N_1667);
or U2389 (N_2389,N_1530,N_1708);
or U2390 (N_2390,N_1101,N_1847);
or U2391 (N_2391,N_1804,N_1309);
or U2392 (N_2392,N_1244,N_1706);
nand U2393 (N_2393,N_1167,N_1491);
or U2394 (N_2394,N_1410,N_1126);
or U2395 (N_2395,N_1787,N_1253);
and U2396 (N_2396,N_1118,N_1427);
and U2397 (N_2397,N_1940,N_1362);
nor U2398 (N_2398,N_1679,N_1205);
and U2399 (N_2399,N_1086,N_1277);
nor U2400 (N_2400,N_1242,N_1228);
and U2401 (N_2401,N_1858,N_1022);
or U2402 (N_2402,N_1157,N_1856);
nor U2403 (N_2403,N_1513,N_1385);
or U2404 (N_2404,N_1771,N_1370);
nor U2405 (N_2405,N_1934,N_1324);
and U2406 (N_2406,N_1363,N_1574);
and U2407 (N_2407,N_1375,N_1476);
or U2408 (N_2408,N_1537,N_1138);
or U2409 (N_2409,N_1924,N_1071);
nand U2410 (N_2410,N_1033,N_1541);
nand U2411 (N_2411,N_1756,N_1340);
or U2412 (N_2412,N_1740,N_1383);
nand U2413 (N_2413,N_1123,N_1163);
or U2414 (N_2414,N_1586,N_1068);
or U2415 (N_2415,N_1182,N_1405);
and U2416 (N_2416,N_1629,N_1302);
and U2417 (N_2417,N_1477,N_1170);
and U2418 (N_2418,N_1268,N_1551);
nand U2419 (N_2419,N_1454,N_1245);
nor U2420 (N_2420,N_1252,N_1669);
nor U2421 (N_2421,N_1573,N_1397);
or U2422 (N_2422,N_1279,N_1990);
or U2423 (N_2423,N_1613,N_1345);
nand U2424 (N_2424,N_1897,N_1677);
nand U2425 (N_2425,N_1455,N_1536);
nor U2426 (N_2426,N_1638,N_1266);
nand U2427 (N_2427,N_1103,N_1377);
or U2428 (N_2428,N_1854,N_1930);
and U2429 (N_2429,N_1783,N_1717);
and U2430 (N_2430,N_1795,N_1906);
or U2431 (N_2431,N_1140,N_1136);
or U2432 (N_2432,N_1095,N_1051);
nand U2433 (N_2433,N_1040,N_1915);
xor U2434 (N_2434,N_1256,N_1608);
and U2435 (N_2435,N_1327,N_1369);
nor U2436 (N_2436,N_1888,N_1695);
nor U2437 (N_2437,N_1816,N_1723);
or U2438 (N_2438,N_1423,N_1053);
or U2439 (N_2439,N_1139,N_1820);
nand U2440 (N_2440,N_1296,N_1778);
nand U2441 (N_2441,N_1587,N_1197);
nor U2442 (N_2442,N_1817,N_1475);
nor U2443 (N_2443,N_1506,N_1902);
and U2444 (N_2444,N_1282,N_1497);
or U2445 (N_2445,N_1307,N_1125);
nand U2446 (N_2446,N_1038,N_1962);
nand U2447 (N_2447,N_1627,N_1952);
or U2448 (N_2448,N_1459,N_1690);
nor U2449 (N_2449,N_1895,N_1450);
nand U2450 (N_2450,N_1845,N_1994);
nand U2451 (N_2451,N_1042,N_1403);
and U2452 (N_2452,N_1007,N_1532);
nor U2453 (N_2453,N_1745,N_1839);
and U2454 (N_2454,N_1001,N_1694);
or U2455 (N_2455,N_1711,N_1890);
nor U2456 (N_2456,N_1012,N_1615);
nor U2457 (N_2457,N_1046,N_1096);
nor U2458 (N_2458,N_1201,N_1412);
nand U2459 (N_2459,N_1011,N_1612);
and U2460 (N_2460,N_1630,N_1641);
nor U2461 (N_2461,N_1288,N_1772);
nand U2462 (N_2462,N_1899,N_1714);
or U2463 (N_2463,N_1510,N_1548);
nand U2464 (N_2464,N_1595,N_1019);
nor U2465 (N_2465,N_1832,N_1844);
or U2466 (N_2466,N_1632,N_1889);
nand U2467 (N_2467,N_1968,N_1929);
or U2468 (N_2468,N_1274,N_1607);
and U2469 (N_2469,N_1527,N_1083);
or U2470 (N_2470,N_1985,N_1166);
or U2471 (N_2471,N_1127,N_1013);
and U2472 (N_2472,N_1986,N_1533);
nand U2473 (N_2473,N_1421,N_1154);
nand U2474 (N_2474,N_1179,N_1386);
and U2475 (N_2475,N_1730,N_1646);
nand U2476 (N_2476,N_1306,N_1768);
nand U2477 (N_2477,N_1997,N_1743);
or U2478 (N_2478,N_1867,N_1021);
nand U2479 (N_2479,N_1830,N_1508);
nand U2480 (N_2480,N_1025,N_1878);
nor U2481 (N_2481,N_1785,N_1725);
and U2482 (N_2482,N_1931,N_1211);
and U2483 (N_2483,N_1803,N_1223);
nor U2484 (N_2484,N_1183,N_1511);
or U2485 (N_2485,N_1172,N_1555);
or U2486 (N_2486,N_1406,N_1518);
or U2487 (N_2487,N_1374,N_1954);
nand U2488 (N_2488,N_1018,N_1534);
xnor U2489 (N_2489,N_1222,N_1119);
nor U2490 (N_2490,N_1549,N_1334);
nand U2491 (N_2491,N_1184,N_1219);
nor U2492 (N_2492,N_1900,N_1284);
nor U2493 (N_2493,N_1543,N_1063);
nand U2494 (N_2494,N_1373,N_1999);
or U2495 (N_2495,N_1234,N_1735);
nand U2496 (N_2496,N_1957,N_1736);
nand U2497 (N_2497,N_1187,N_1788);
nand U2498 (N_2498,N_1738,N_1663);
or U2499 (N_2499,N_1642,N_1734);
or U2500 (N_2500,N_1633,N_1043);
or U2501 (N_2501,N_1899,N_1139);
or U2502 (N_2502,N_1629,N_1851);
or U2503 (N_2503,N_1789,N_1299);
nor U2504 (N_2504,N_1580,N_1745);
xnor U2505 (N_2505,N_1669,N_1972);
nor U2506 (N_2506,N_1359,N_1160);
nand U2507 (N_2507,N_1456,N_1413);
nor U2508 (N_2508,N_1259,N_1623);
nand U2509 (N_2509,N_1143,N_1129);
and U2510 (N_2510,N_1539,N_1009);
nor U2511 (N_2511,N_1715,N_1432);
nand U2512 (N_2512,N_1257,N_1089);
nand U2513 (N_2513,N_1280,N_1482);
and U2514 (N_2514,N_1148,N_1902);
xor U2515 (N_2515,N_1953,N_1872);
nor U2516 (N_2516,N_1174,N_1841);
or U2517 (N_2517,N_1755,N_1900);
or U2518 (N_2518,N_1495,N_1141);
nor U2519 (N_2519,N_1827,N_1495);
nor U2520 (N_2520,N_1633,N_1618);
xnor U2521 (N_2521,N_1173,N_1249);
and U2522 (N_2522,N_1848,N_1483);
or U2523 (N_2523,N_1721,N_1599);
nor U2524 (N_2524,N_1648,N_1841);
nor U2525 (N_2525,N_1876,N_1313);
or U2526 (N_2526,N_1947,N_1496);
nor U2527 (N_2527,N_1655,N_1878);
nor U2528 (N_2528,N_1019,N_1633);
nor U2529 (N_2529,N_1136,N_1938);
nor U2530 (N_2530,N_1183,N_1136);
and U2531 (N_2531,N_1669,N_1208);
nand U2532 (N_2532,N_1714,N_1745);
nand U2533 (N_2533,N_1822,N_1989);
or U2534 (N_2534,N_1621,N_1675);
and U2535 (N_2535,N_1703,N_1224);
nand U2536 (N_2536,N_1025,N_1664);
or U2537 (N_2537,N_1971,N_1025);
and U2538 (N_2538,N_1761,N_1029);
nand U2539 (N_2539,N_1556,N_1527);
nand U2540 (N_2540,N_1660,N_1176);
nand U2541 (N_2541,N_1483,N_1594);
and U2542 (N_2542,N_1365,N_1299);
nor U2543 (N_2543,N_1848,N_1563);
or U2544 (N_2544,N_1831,N_1409);
and U2545 (N_2545,N_1537,N_1600);
nor U2546 (N_2546,N_1158,N_1030);
nor U2547 (N_2547,N_1106,N_1654);
or U2548 (N_2548,N_1986,N_1074);
nand U2549 (N_2549,N_1037,N_1073);
and U2550 (N_2550,N_1192,N_1017);
or U2551 (N_2551,N_1929,N_1160);
and U2552 (N_2552,N_1556,N_1203);
nor U2553 (N_2553,N_1287,N_1032);
nor U2554 (N_2554,N_1967,N_1720);
nor U2555 (N_2555,N_1196,N_1974);
nand U2556 (N_2556,N_1905,N_1792);
and U2557 (N_2557,N_1952,N_1626);
or U2558 (N_2558,N_1279,N_1477);
nor U2559 (N_2559,N_1029,N_1684);
nand U2560 (N_2560,N_1846,N_1380);
nand U2561 (N_2561,N_1952,N_1389);
and U2562 (N_2562,N_1302,N_1376);
nor U2563 (N_2563,N_1150,N_1421);
nand U2564 (N_2564,N_1681,N_1375);
nand U2565 (N_2565,N_1367,N_1017);
nor U2566 (N_2566,N_1902,N_1540);
and U2567 (N_2567,N_1350,N_1075);
and U2568 (N_2568,N_1121,N_1913);
nand U2569 (N_2569,N_1612,N_1428);
nand U2570 (N_2570,N_1287,N_1378);
and U2571 (N_2571,N_1185,N_1129);
nand U2572 (N_2572,N_1111,N_1774);
nor U2573 (N_2573,N_1061,N_1764);
and U2574 (N_2574,N_1615,N_1466);
nand U2575 (N_2575,N_1803,N_1561);
nor U2576 (N_2576,N_1499,N_1104);
nand U2577 (N_2577,N_1606,N_1373);
nor U2578 (N_2578,N_1016,N_1885);
or U2579 (N_2579,N_1088,N_1836);
or U2580 (N_2580,N_1010,N_1132);
nor U2581 (N_2581,N_1422,N_1972);
or U2582 (N_2582,N_1945,N_1248);
or U2583 (N_2583,N_1741,N_1052);
or U2584 (N_2584,N_1367,N_1365);
or U2585 (N_2585,N_1334,N_1682);
and U2586 (N_2586,N_1045,N_1085);
and U2587 (N_2587,N_1360,N_1263);
or U2588 (N_2588,N_1357,N_1621);
or U2589 (N_2589,N_1816,N_1987);
nor U2590 (N_2590,N_1963,N_1085);
nor U2591 (N_2591,N_1474,N_1486);
nand U2592 (N_2592,N_1934,N_1540);
nor U2593 (N_2593,N_1089,N_1228);
nor U2594 (N_2594,N_1384,N_1311);
nor U2595 (N_2595,N_1484,N_1678);
nand U2596 (N_2596,N_1410,N_1100);
and U2597 (N_2597,N_1445,N_1878);
nand U2598 (N_2598,N_1656,N_1265);
and U2599 (N_2599,N_1679,N_1320);
nand U2600 (N_2600,N_1447,N_1871);
or U2601 (N_2601,N_1773,N_1146);
nor U2602 (N_2602,N_1619,N_1108);
nor U2603 (N_2603,N_1809,N_1913);
or U2604 (N_2604,N_1615,N_1197);
and U2605 (N_2605,N_1722,N_1952);
and U2606 (N_2606,N_1565,N_1125);
or U2607 (N_2607,N_1178,N_1880);
and U2608 (N_2608,N_1895,N_1725);
and U2609 (N_2609,N_1861,N_1401);
nor U2610 (N_2610,N_1273,N_1079);
nand U2611 (N_2611,N_1535,N_1939);
or U2612 (N_2612,N_1382,N_1778);
or U2613 (N_2613,N_1899,N_1539);
nor U2614 (N_2614,N_1343,N_1853);
or U2615 (N_2615,N_1773,N_1744);
nor U2616 (N_2616,N_1337,N_1296);
nor U2617 (N_2617,N_1686,N_1835);
nand U2618 (N_2618,N_1818,N_1880);
or U2619 (N_2619,N_1147,N_1903);
nor U2620 (N_2620,N_1744,N_1790);
or U2621 (N_2621,N_1079,N_1509);
and U2622 (N_2622,N_1458,N_1844);
nor U2623 (N_2623,N_1225,N_1923);
and U2624 (N_2624,N_1111,N_1096);
nand U2625 (N_2625,N_1246,N_1721);
or U2626 (N_2626,N_1185,N_1602);
or U2627 (N_2627,N_1043,N_1750);
or U2628 (N_2628,N_1832,N_1428);
nor U2629 (N_2629,N_1084,N_1059);
and U2630 (N_2630,N_1234,N_1844);
or U2631 (N_2631,N_1721,N_1431);
or U2632 (N_2632,N_1132,N_1068);
nor U2633 (N_2633,N_1869,N_1876);
or U2634 (N_2634,N_1388,N_1827);
and U2635 (N_2635,N_1593,N_1697);
or U2636 (N_2636,N_1669,N_1223);
and U2637 (N_2637,N_1175,N_1768);
nand U2638 (N_2638,N_1483,N_1103);
nor U2639 (N_2639,N_1604,N_1204);
and U2640 (N_2640,N_1854,N_1270);
or U2641 (N_2641,N_1374,N_1085);
and U2642 (N_2642,N_1381,N_1691);
nand U2643 (N_2643,N_1956,N_1448);
nand U2644 (N_2644,N_1964,N_1314);
nor U2645 (N_2645,N_1534,N_1086);
nor U2646 (N_2646,N_1892,N_1308);
or U2647 (N_2647,N_1660,N_1443);
nand U2648 (N_2648,N_1981,N_1633);
or U2649 (N_2649,N_1121,N_1337);
nor U2650 (N_2650,N_1110,N_1020);
and U2651 (N_2651,N_1920,N_1048);
nand U2652 (N_2652,N_1255,N_1196);
xor U2653 (N_2653,N_1374,N_1287);
nor U2654 (N_2654,N_1281,N_1679);
nand U2655 (N_2655,N_1223,N_1784);
or U2656 (N_2656,N_1629,N_1392);
or U2657 (N_2657,N_1865,N_1556);
nor U2658 (N_2658,N_1731,N_1222);
or U2659 (N_2659,N_1497,N_1105);
nor U2660 (N_2660,N_1057,N_1989);
nand U2661 (N_2661,N_1820,N_1282);
nor U2662 (N_2662,N_1319,N_1055);
and U2663 (N_2663,N_1563,N_1131);
or U2664 (N_2664,N_1788,N_1268);
nand U2665 (N_2665,N_1062,N_1908);
nor U2666 (N_2666,N_1625,N_1374);
nor U2667 (N_2667,N_1908,N_1235);
or U2668 (N_2668,N_1287,N_1562);
and U2669 (N_2669,N_1258,N_1097);
nor U2670 (N_2670,N_1962,N_1443);
nand U2671 (N_2671,N_1393,N_1168);
and U2672 (N_2672,N_1495,N_1638);
or U2673 (N_2673,N_1705,N_1263);
nand U2674 (N_2674,N_1762,N_1708);
nand U2675 (N_2675,N_1745,N_1260);
or U2676 (N_2676,N_1477,N_1003);
nand U2677 (N_2677,N_1235,N_1265);
or U2678 (N_2678,N_1631,N_1128);
or U2679 (N_2679,N_1996,N_1432);
nor U2680 (N_2680,N_1475,N_1453);
nand U2681 (N_2681,N_1387,N_1027);
nand U2682 (N_2682,N_1768,N_1435);
nand U2683 (N_2683,N_1373,N_1492);
and U2684 (N_2684,N_1863,N_1406);
and U2685 (N_2685,N_1082,N_1160);
nand U2686 (N_2686,N_1760,N_1126);
and U2687 (N_2687,N_1044,N_1003);
nor U2688 (N_2688,N_1611,N_1935);
nor U2689 (N_2689,N_1513,N_1511);
or U2690 (N_2690,N_1499,N_1970);
and U2691 (N_2691,N_1296,N_1595);
and U2692 (N_2692,N_1741,N_1896);
nand U2693 (N_2693,N_1461,N_1569);
and U2694 (N_2694,N_1083,N_1077);
nor U2695 (N_2695,N_1622,N_1913);
and U2696 (N_2696,N_1182,N_1126);
nor U2697 (N_2697,N_1692,N_1385);
nor U2698 (N_2698,N_1659,N_1267);
and U2699 (N_2699,N_1059,N_1305);
or U2700 (N_2700,N_1332,N_1364);
and U2701 (N_2701,N_1583,N_1599);
and U2702 (N_2702,N_1058,N_1569);
nand U2703 (N_2703,N_1989,N_1128);
nor U2704 (N_2704,N_1353,N_1689);
and U2705 (N_2705,N_1444,N_1552);
nand U2706 (N_2706,N_1152,N_1405);
or U2707 (N_2707,N_1632,N_1092);
nand U2708 (N_2708,N_1447,N_1861);
nor U2709 (N_2709,N_1035,N_1995);
nor U2710 (N_2710,N_1381,N_1708);
nor U2711 (N_2711,N_1204,N_1893);
and U2712 (N_2712,N_1666,N_1688);
nor U2713 (N_2713,N_1628,N_1535);
nor U2714 (N_2714,N_1550,N_1128);
nand U2715 (N_2715,N_1520,N_1376);
and U2716 (N_2716,N_1024,N_1368);
or U2717 (N_2717,N_1066,N_1231);
nand U2718 (N_2718,N_1250,N_1082);
and U2719 (N_2719,N_1199,N_1827);
nand U2720 (N_2720,N_1046,N_1825);
and U2721 (N_2721,N_1896,N_1514);
nor U2722 (N_2722,N_1337,N_1248);
or U2723 (N_2723,N_1625,N_1515);
nand U2724 (N_2724,N_1181,N_1368);
nand U2725 (N_2725,N_1773,N_1743);
and U2726 (N_2726,N_1731,N_1943);
and U2727 (N_2727,N_1550,N_1181);
nand U2728 (N_2728,N_1268,N_1893);
or U2729 (N_2729,N_1391,N_1367);
nor U2730 (N_2730,N_1458,N_1609);
nor U2731 (N_2731,N_1960,N_1350);
or U2732 (N_2732,N_1129,N_1223);
or U2733 (N_2733,N_1529,N_1338);
or U2734 (N_2734,N_1214,N_1873);
or U2735 (N_2735,N_1067,N_1590);
nand U2736 (N_2736,N_1286,N_1374);
xor U2737 (N_2737,N_1225,N_1404);
or U2738 (N_2738,N_1525,N_1871);
nand U2739 (N_2739,N_1090,N_1165);
nand U2740 (N_2740,N_1311,N_1481);
and U2741 (N_2741,N_1498,N_1873);
nand U2742 (N_2742,N_1670,N_1553);
nand U2743 (N_2743,N_1835,N_1089);
nand U2744 (N_2744,N_1166,N_1376);
nor U2745 (N_2745,N_1895,N_1003);
nand U2746 (N_2746,N_1890,N_1093);
or U2747 (N_2747,N_1702,N_1257);
and U2748 (N_2748,N_1495,N_1728);
and U2749 (N_2749,N_1931,N_1914);
nor U2750 (N_2750,N_1409,N_1112);
nand U2751 (N_2751,N_1477,N_1854);
or U2752 (N_2752,N_1220,N_1099);
or U2753 (N_2753,N_1374,N_1438);
nand U2754 (N_2754,N_1889,N_1393);
nor U2755 (N_2755,N_1894,N_1069);
nor U2756 (N_2756,N_1336,N_1318);
or U2757 (N_2757,N_1960,N_1668);
or U2758 (N_2758,N_1287,N_1189);
nor U2759 (N_2759,N_1626,N_1216);
nor U2760 (N_2760,N_1560,N_1635);
nor U2761 (N_2761,N_1416,N_1195);
nor U2762 (N_2762,N_1160,N_1874);
nor U2763 (N_2763,N_1361,N_1912);
nor U2764 (N_2764,N_1928,N_1836);
and U2765 (N_2765,N_1388,N_1742);
and U2766 (N_2766,N_1811,N_1377);
and U2767 (N_2767,N_1136,N_1286);
nand U2768 (N_2768,N_1802,N_1021);
and U2769 (N_2769,N_1500,N_1478);
nand U2770 (N_2770,N_1482,N_1935);
xnor U2771 (N_2771,N_1594,N_1823);
and U2772 (N_2772,N_1675,N_1850);
nand U2773 (N_2773,N_1346,N_1776);
nor U2774 (N_2774,N_1038,N_1659);
nor U2775 (N_2775,N_1778,N_1186);
or U2776 (N_2776,N_1510,N_1599);
nand U2777 (N_2777,N_1378,N_1844);
or U2778 (N_2778,N_1192,N_1113);
nand U2779 (N_2779,N_1297,N_1972);
and U2780 (N_2780,N_1463,N_1688);
nor U2781 (N_2781,N_1456,N_1573);
nand U2782 (N_2782,N_1847,N_1724);
nand U2783 (N_2783,N_1395,N_1556);
nand U2784 (N_2784,N_1648,N_1472);
or U2785 (N_2785,N_1924,N_1758);
nand U2786 (N_2786,N_1654,N_1436);
nand U2787 (N_2787,N_1007,N_1439);
nor U2788 (N_2788,N_1224,N_1766);
nor U2789 (N_2789,N_1796,N_1998);
nand U2790 (N_2790,N_1176,N_1570);
and U2791 (N_2791,N_1466,N_1746);
nand U2792 (N_2792,N_1898,N_1155);
nand U2793 (N_2793,N_1039,N_1223);
nand U2794 (N_2794,N_1306,N_1494);
nand U2795 (N_2795,N_1815,N_1534);
or U2796 (N_2796,N_1293,N_1309);
nand U2797 (N_2797,N_1312,N_1755);
nor U2798 (N_2798,N_1402,N_1950);
nand U2799 (N_2799,N_1118,N_1150);
nor U2800 (N_2800,N_1003,N_1084);
or U2801 (N_2801,N_1914,N_1119);
nand U2802 (N_2802,N_1714,N_1120);
or U2803 (N_2803,N_1708,N_1757);
nand U2804 (N_2804,N_1101,N_1731);
nand U2805 (N_2805,N_1227,N_1460);
nand U2806 (N_2806,N_1441,N_1573);
nor U2807 (N_2807,N_1064,N_1693);
or U2808 (N_2808,N_1442,N_1303);
or U2809 (N_2809,N_1929,N_1197);
or U2810 (N_2810,N_1596,N_1103);
or U2811 (N_2811,N_1471,N_1541);
or U2812 (N_2812,N_1334,N_1988);
nor U2813 (N_2813,N_1680,N_1461);
nand U2814 (N_2814,N_1148,N_1048);
nor U2815 (N_2815,N_1814,N_1734);
nor U2816 (N_2816,N_1078,N_1290);
or U2817 (N_2817,N_1642,N_1994);
and U2818 (N_2818,N_1218,N_1276);
or U2819 (N_2819,N_1088,N_1399);
or U2820 (N_2820,N_1731,N_1261);
nand U2821 (N_2821,N_1423,N_1514);
or U2822 (N_2822,N_1972,N_1772);
nand U2823 (N_2823,N_1914,N_1421);
nand U2824 (N_2824,N_1503,N_1384);
nor U2825 (N_2825,N_1882,N_1668);
nor U2826 (N_2826,N_1693,N_1314);
and U2827 (N_2827,N_1847,N_1878);
nand U2828 (N_2828,N_1467,N_1661);
and U2829 (N_2829,N_1124,N_1256);
and U2830 (N_2830,N_1263,N_1508);
and U2831 (N_2831,N_1027,N_1059);
or U2832 (N_2832,N_1948,N_1856);
or U2833 (N_2833,N_1028,N_1003);
or U2834 (N_2834,N_1184,N_1165);
or U2835 (N_2835,N_1815,N_1820);
or U2836 (N_2836,N_1089,N_1887);
or U2837 (N_2837,N_1361,N_1702);
and U2838 (N_2838,N_1932,N_1167);
nand U2839 (N_2839,N_1094,N_1542);
nand U2840 (N_2840,N_1436,N_1062);
nand U2841 (N_2841,N_1930,N_1190);
or U2842 (N_2842,N_1066,N_1457);
or U2843 (N_2843,N_1086,N_1123);
and U2844 (N_2844,N_1918,N_1081);
and U2845 (N_2845,N_1957,N_1687);
nor U2846 (N_2846,N_1270,N_1866);
nand U2847 (N_2847,N_1611,N_1322);
and U2848 (N_2848,N_1302,N_1790);
nor U2849 (N_2849,N_1279,N_1256);
or U2850 (N_2850,N_1697,N_1208);
nand U2851 (N_2851,N_1129,N_1777);
or U2852 (N_2852,N_1795,N_1396);
nand U2853 (N_2853,N_1467,N_1984);
xor U2854 (N_2854,N_1124,N_1902);
nor U2855 (N_2855,N_1822,N_1969);
nand U2856 (N_2856,N_1465,N_1986);
nand U2857 (N_2857,N_1983,N_1278);
nor U2858 (N_2858,N_1932,N_1733);
and U2859 (N_2859,N_1374,N_1164);
nor U2860 (N_2860,N_1573,N_1900);
and U2861 (N_2861,N_1246,N_1353);
and U2862 (N_2862,N_1170,N_1725);
and U2863 (N_2863,N_1415,N_1016);
nor U2864 (N_2864,N_1460,N_1700);
nor U2865 (N_2865,N_1967,N_1638);
or U2866 (N_2866,N_1741,N_1735);
nor U2867 (N_2867,N_1866,N_1440);
and U2868 (N_2868,N_1321,N_1573);
and U2869 (N_2869,N_1043,N_1291);
and U2870 (N_2870,N_1073,N_1747);
and U2871 (N_2871,N_1324,N_1652);
nand U2872 (N_2872,N_1311,N_1933);
or U2873 (N_2873,N_1444,N_1689);
nand U2874 (N_2874,N_1531,N_1812);
nor U2875 (N_2875,N_1478,N_1641);
nand U2876 (N_2876,N_1220,N_1087);
and U2877 (N_2877,N_1780,N_1563);
and U2878 (N_2878,N_1767,N_1243);
nand U2879 (N_2879,N_1853,N_1156);
and U2880 (N_2880,N_1301,N_1189);
nor U2881 (N_2881,N_1704,N_1743);
nand U2882 (N_2882,N_1622,N_1523);
or U2883 (N_2883,N_1102,N_1058);
or U2884 (N_2884,N_1190,N_1489);
or U2885 (N_2885,N_1610,N_1631);
and U2886 (N_2886,N_1096,N_1064);
nand U2887 (N_2887,N_1154,N_1808);
or U2888 (N_2888,N_1121,N_1592);
nor U2889 (N_2889,N_1134,N_1661);
and U2890 (N_2890,N_1374,N_1822);
nor U2891 (N_2891,N_1859,N_1238);
nand U2892 (N_2892,N_1819,N_1425);
or U2893 (N_2893,N_1052,N_1131);
and U2894 (N_2894,N_1291,N_1531);
nor U2895 (N_2895,N_1144,N_1426);
or U2896 (N_2896,N_1769,N_1789);
nor U2897 (N_2897,N_1334,N_1206);
nand U2898 (N_2898,N_1077,N_1747);
and U2899 (N_2899,N_1139,N_1499);
or U2900 (N_2900,N_1409,N_1652);
or U2901 (N_2901,N_1235,N_1191);
or U2902 (N_2902,N_1009,N_1086);
nand U2903 (N_2903,N_1046,N_1988);
nor U2904 (N_2904,N_1448,N_1500);
and U2905 (N_2905,N_1465,N_1974);
nor U2906 (N_2906,N_1214,N_1001);
and U2907 (N_2907,N_1784,N_1281);
nand U2908 (N_2908,N_1189,N_1732);
nor U2909 (N_2909,N_1264,N_1936);
or U2910 (N_2910,N_1821,N_1127);
or U2911 (N_2911,N_1241,N_1226);
nand U2912 (N_2912,N_1382,N_1243);
nor U2913 (N_2913,N_1132,N_1452);
and U2914 (N_2914,N_1442,N_1978);
nor U2915 (N_2915,N_1244,N_1047);
nor U2916 (N_2916,N_1931,N_1064);
nor U2917 (N_2917,N_1984,N_1820);
nand U2918 (N_2918,N_1716,N_1199);
and U2919 (N_2919,N_1506,N_1225);
nor U2920 (N_2920,N_1242,N_1159);
and U2921 (N_2921,N_1100,N_1319);
nor U2922 (N_2922,N_1734,N_1892);
nand U2923 (N_2923,N_1367,N_1441);
nand U2924 (N_2924,N_1777,N_1915);
nand U2925 (N_2925,N_1067,N_1733);
and U2926 (N_2926,N_1975,N_1743);
nand U2927 (N_2927,N_1612,N_1125);
and U2928 (N_2928,N_1255,N_1964);
and U2929 (N_2929,N_1047,N_1027);
and U2930 (N_2930,N_1250,N_1021);
or U2931 (N_2931,N_1082,N_1401);
or U2932 (N_2932,N_1319,N_1202);
and U2933 (N_2933,N_1638,N_1863);
or U2934 (N_2934,N_1666,N_1929);
nand U2935 (N_2935,N_1515,N_1054);
and U2936 (N_2936,N_1788,N_1388);
nand U2937 (N_2937,N_1895,N_1438);
nand U2938 (N_2938,N_1574,N_1883);
nor U2939 (N_2939,N_1228,N_1052);
nor U2940 (N_2940,N_1966,N_1003);
and U2941 (N_2941,N_1719,N_1360);
and U2942 (N_2942,N_1101,N_1446);
nor U2943 (N_2943,N_1630,N_1522);
nor U2944 (N_2944,N_1658,N_1053);
nor U2945 (N_2945,N_1707,N_1612);
or U2946 (N_2946,N_1478,N_1240);
or U2947 (N_2947,N_1633,N_1968);
nor U2948 (N_2948,N_1644,N_1604);
nor U2949 (N_2949,N_1756,N_1914);
or U2950 (N_2950,N_1054,N_1889);
or U2951 (N_2951,N_1789,N_1553);
nor U2952 (N_2952,N_1927,N_1006);
or U2953 (N_2953,N_1796,N_1896);
and U2954 (N_2954,N_1909,N_1320);
or U2955 (N_2955,N_1870,N_1453);
or U2956 (N_2956,N_1788,N_1376);
nand U2957 (N_2957,N_1119,N_1135);
or U2958 (N_2958,N_1466,N_1126);
nor U2959 (N_2959,N_1749,N_1397);
and U2960 (N_2960,N_1951,N_1533);
or U2961 (N_2961,N_1380,N_1271);
or U2962 (N_2962,N_1724,N_1858);
or U2963 (N_2963,N_1691,N_1745);
nand U2964 (N_2964,N_1477,N_1412);
or U2965 (N_2965,N_1422,N_1075);
nor U2966 (N_2966,N_1530,N_1591);
or U2967 (N_2967,N_1689,N_1993);
nand U2968 (N_2968,N_1315,N_1999);
nand U2969 (N_2969,N_1663,N_1820);
or U2970 (N_2970,N_1271,N_1687);
and U2971 (N_2971,N_1425,N_1889);
or U2972 (N_2972,N_1531,N_1892);
nand U2973 (N_2973,N_1828,N_1798);
or U2974 (N_2974,N_1548,N_1726);
and U2975 (N_2975,N_1305,N_1774);
and U2976 (N_2976,N_1886,N_1577);
nor U2977 (N_2977,N_1524,N_1295);
and U2978 (N_2978,N_1609,N_1313);
and U2979 (N_2979,N_1800,N_1409);
or U2980 (N_2980,N_1744,N_1593);
nand U2981 (N_2981,N_1464,N_1906);
or U2982 (N_2982,N_1652,N_1242);
nor U2983 (N_2983,N_1806,N_1584);
nor U2984 (N_2984,N_1357,N_1615);
and U2985 (N_2985,N_1134,N_1500);
and U2986 (N_2986,N_1739,N_1245);
nand U2987 (N_2987,N_1633,N_1012);
nor U2988 (N_2988,N_1679,N_1858);
or U2989 (N_2989,N_1051,N_1908);
or U2990 (N_2990,N_1557,N_1266);
or U2991 (N_2991,N_1249,N_1370);
nor U2992 (N_2992,N_1007,N_1547);
nor U2993 (N_2993,N_1906,N_1101);
xnor U2994 (N_2994,N_1857,N_1676);
nand U2995 (N_2995,N_1313,N_1884);
or U2996 (N_2996,N_1406,N_1586);
nor U2997 (N_2997,N_1779,N_1521);
nor U2998 (N_2998,N_1145,N_1946);
or U2999 (N_2999,N_1104,N_1472);
or U3000 (N_3000,N_2236,N_2483);
nand U3001 (N_3001,N_2572,N_2391);
nor U3002 (N_3002,N_2747,N_2156);
or U3003 (N_3003,N_2459,N_2606);
nand U3004 (N_3004,N_2494,N_2290);
nand U3005 (N_3005,N_2099,N_2939);
or U3006 (N_3006,N_2071,N_2855);
or U3007 (N_3007,N_2949,N_2737);
nor U3008 (N_3008,N_2402,N_2348);
or U3009 (N_3009,N_2500,N_2049);
or U3010 (N_3010,N_2222,N_2374);
and U3011 (N_3011,N_2343,N_2937);
xor U3012 (N_3012,N_2132,N_2484);
or U3013 (N_3013,N_2018,N_2330);
nand U3014 (N_3014,N_2337,N_2151);
and U3015 (N_3015,N_2215,N_2858);
or U3016 (N_3016,N_2848,N_2158);
or U3017 (N_3017,N_2629,N_2845);
nand U3018 (N_3018,N_2295,N_2006);
or U3019 (N_3019,N_2147,N_2046);
and U3020 (N_3020,N_2639,N_2351);
nor U3021 (N_3021,N_2318,N_2405);
nand U3022 (N_3022,N_2204,N_2449);
nand U3023 (N_3023,N_2037,N_2661);
nand U3024 (N_3024,N_2008,N_2895);
or U3025 (N_3025,N_2186,N_2646);
nand U3026 (N_3026,N_2772,N_2864);
nand U3027 (N_3027,N_2160,N_2353);
nor U3028 (N_3028,N_2774,N_2728);
and U3029 (N_3029,N_2591,N_2656);
nand U3030 (N_3030,N_2423,N_2170);
nand U3031 (N_3031,N_2114,N_2061);
or U3032 (N_3032,N_2047,N_2091);
or U3033 (N_3033,N_2773,N_2513);
and U3034 (N_3034,N_2636,N_2843);
or U3035 (N_3035,N_2751,N_2805);
nor U3036 (N_3036,N_2291,N_2014);
nor U3037 (N_3037,N_2975,N_2896);
nor U3038 (N_3038,N_2744,N_2175);
nand U3039 (N_3039,N_2396,N_2732);
nor U3040 (N_3040,N_2064,N_2976);
and U3041 (N_3041,N_2922,N_2902);
nor U3042 (N_3042,N_2223,N_2561);
xor U3043 (N_3043,N_2971,N_2936);
nor U3044 (N_3044,N_2205,N_2134);
or U3045 (N_3045,N_2958,N_2955);
nand U3046 (N_3046,N_2954,N_2106);
nand U3047 (N_3047,N_2611,N_2225);
or U3048 (N_3048,N_2947,N_2441);
or U3049 (N_3049,N_2548,N_2682);
nor U3050 (N_3050,N_2228,N_2809);
nand U3051 (N_3051,N_2305,N_2480);
nand U3052 (N_3052,N_2662,N_2798);
or U3053 (N_3053,N_2694,N_2479);
or U3054 (N_3054,N_2509,N_2770);
and U3055 (N_3055,N_2393,N_2850);
nand U3056 (N_3056,N_2093,N_2900);
and U3057 (N_3057,N_2054,N_2825);
or U3058 (N_3058,N_2765,N_2553);
and U3059 (N_3059,N_2658,N_2621);
nor U3060 (N_3060,N_2407,N_2886);
nor U3061 (N_3061,N_2303,N_2516);
or U3062 (N_3062,N_2188,N_2543);
and U3063 (N_3063,N_2385,N_2574);
or U3064 (N_3064,N_2389,N_2628);
nand U3065 (N_3065,N_2721,N_2001);
xor U3066 (N_3066,N_2083,N_2795);
or U3067 (N_3067,N_2498,N_2078);
nor U3068 (N_3068,N_2255,N_2470);
and U3069 (N_3069,N_2388,N_2741);
and U3070 (N_3070,N_2802,N_2844);
or U3071 (N_3071,N_2398,N_2137);
nand U3072 (N_3072,N_2586,N_2101);
nor U3073 (N_3073,N_2050,N_2853);
and U3074 (N_3074,N_2691,N_2242);
and U3075 (N_3075,N_2571,N_2984);
or U3076 (N_3076,N_2076,N_2560);
nor U3077 (N_3077,N_2699,N_2635);
and U3078 (N_3078,N_2200,N_2593);
or U3079 (N_3079,N_2512,N_2127);
and U3080 (N_3080,N_2240,N_2720);
and U3081 (N_3081,N_2846,N_2447);
nand U3082 (N_3082,N_2820,N_2442);
nor U3083 (N_3083,N_2882,N_2644);
or U3084 (N_3084,N_2036,N_2022);
nor U3085 (N_3085,N_2126,N_2775);
nor U3086 (N_3086,N_2012,N_2670);
or U3087 (N_3087,N_2052,N_2196);
or U3088 (N_3088,N_2519,N_2929);
and U3089 (N_3089,N_2655,N_2739);
nor U3090 (N_3090,N_2950,N_2282);
nand U3091 (N_3091,N_2813,N_2254);
or U3092 (N_3092,N_2068,N_2179);
nor U3093 (N_3093,N_2811,N_2302);
or U3094 (N_3094,N_2030,N_2608);
nand U3095 (N_3095,N_2856,N_2368);
and U3096 (N_3096,N_2273,N_2003);
and U3097 (N_3097,N_2308,N_2214);
nor U3098 (N_3098,N_2503,N_2096);
nor U3099 (N_3099,N_2857,N_2476);
or U3100 (N_3100,N_2039,N_2812);
or U3101 (N_3101,N_2792,N_2007);
or U3102 (N_3102,N_2425,N_2314);
nor U3103 (N_3103,N_2582,N_2104);
and U3104 (N_3104,N_2903,N_2005);
nand U3105 (N_3105,N_2199,N_2926);
nor U3106 (N_3106,N_2729,N_2042);
and U3107 (N_3107,N_2438,N_2831);
nand U3108 (N_3108,N_2167,N_2779);
nand U3109 (N_3109,N_2111,N_2239);
nand U3110 (N_3110,N_2883,N_2326);
or U3111 (N_3111,N_2643,N_2235);
nand U3112 (N_3112,N_2311,N_2446);
and U3113 (N_3113,N_2803,N_2428);
and U3114 (N_3114,N_2490,N_2709);
nor U3115 (N_3115,N_2650,N_2202);
or U3116 (N_3116,N_2496,N_2766);
xnor U3117 (N_3117,N_2113,N_2991);
or U3118 (N_3118,N_2507,N_2310);
or U3119 (N_3119,N_2679,N_2377);
nand U3120 (N_3120,N_2115,N_2172);
and U3121 (N_3121,N_2725,N_2569);
nand U3122 (N_3122,N_2098,N_2365);
nand U3123 (N_3123,N_2387,N_2349);
nor U3124 (N_3124,N_2433,N_2704);
nor U3125 (N_3125,N_2993,N_2016);
or U3126 (N_3126,N_2434,N_2640);
or U3127 (N_3127,N_2027,N_2359);
nor U3128 (N_3128,N_2164,N_2087);
and U3129 (N_3129,N_2120,N_2514);
nor U3130 (N_3130,N_2762,N_2227);
nand U3131 (N_3131,N_2139,N_2965);
or U3132 (N_3132,N_2794,N_2689);
and U3133 (N_3133,N_2331,N_2505);
nor U3134 (N_3134,N_2998,N_2703);
nand U3135 (N_3135,N_2576,N_2315);
nand U3136 (N_3136,N_2573,N_2759);
or U3137 (N_3137,N_2581,N_2530);
nor U3138 (N_3138,N_2948,N_2231);
xnor U3139 (N_3139,N_2075,N_2243);
nand U3140 (N_3140,N_2609,N_2390);
nand U3141 (N_3141,N_2352,N_2072);
or U3142 (N_3142,N_2994,N_2714);
or U3143 (N_3143,N_2592,N_2383);
and U3144 (N_3144,N_2261,N_2230);
nand U3145 (N_3145,N_2600,N_2804);
and U3146 (N_3146,N_2757,N_2122);
nand U3147 (N_3147,N_2092,N_2019);
xnor U3148 (N_3148,N_2226,N_2817);
nor U3149 (N_3149,N_2945,N_2454);
nor U3150 (N_3150,N_2546,N_2081);
and U3151 (N_3151,N_2289,N_2191);
or U3152 (N_3152,N_2879,N_2545);
nor U3153 (N_3153,N_2304,N_2681);
nand U3154 (N_3154,N_2570,N_2781);
and U3155 (N_3155,N_2686,N_2131);
or U3156 (N_3156,N_2834,N_2916);
or U3157 (N_3157,N_2485,N_2914);
or U3158 (N_3158,N_2985,N_2822);
nand U3159 (N_3159,N_2403,N_2612);
and U3160 (N_3160,N_2642,N_2218);
nor U3161 (N_3161,N_2208,N_2323);
and U3162 (N_3162,N_2904,N_2869);
nor U3163 (N_3163,N_2118,N_2279);
and U3164 (N_3164,N_2453,N_2238);
and U3165 (N_3165,N_2198,N_2373);
nor U3166 (N_3166,N_2515,N_2034);
or U3167 (N_3167,N_2002,N_2893);
nor U3168 (N_3168,N_2938,N_2015);
and U3169 (N_3169,N_2429,N_2815);
nand U3170 (N_3170,N_2038,N_2163);
or U3171 (N_3171,N_2968,N_2927);
and U3172 (N_3172,N_2657,N_2378);
nand U3173 (N_3173,N_2959,N_2934);
or U3174 (N_3174,N_2149,N_2917);
nand U3175 (N_3175,N_2392,N_2241);
nand U3176 (N_3176,N_2767,N_2336);
and U3177 (N_3177,N_2253,N_2418);
and U3178 (N_3178,N_2312,N_2768);
and U3179 (N_3179,N_2731,N_2264);
nand U3180 (N_3180,N_2533,N_2990);
nand U3181 (N_3181,N_2043,N_2918);
nand U3182 (N_3182,N_2908,N_2055);
and U3183 (N_3183,N_2554,N_2652);
and U3184 (N_3184,N_2033,N_2482);
nor U3185 (N_3185,N_2082,N_2262);
or U3186 (N_3186,N_2342,N_2341);
or U3187 (N_3187,N_2563,N_2354);
nor U3188 (N_3188,N_2426,N_2596);
and U3189 (N_3189,N_2088,N_2232);
nor U3190 (N_3190,N_2784,N_2898);
or U3191 (N_3191,N_2880,N_2089);
nor U3192 (N_3192,N_2818,N_2502);
or U3193 (N_3193,N_2004,N_2417);
nor U3194 (N_3194,N_2444,N_2552);
or U3195 (N_3195,N_2165,N_2602);
or U3196 (N_3196,N_2169,N_2233);
and U3197 (N_3197,N_2601,N_2859);
nor U3198 (N_3198,N_2944,N_2736);
nor U3199 (N_3199,N_2931,N_2829);
or U3200 (N_3200,N_2685,N_2209);
or U3201 (N_3201,N_2084,N_2935);
nand U3202 (N_3202,N_2140,N_2473);
or U3203 (N_3203,N_2159,N_2840);
and U3204 (N_3204,N_2674,N_2603);
and U3205 (N_3205,N_2753,N_2746);
nor U3206 (N_3206,N_2266,N_2988);
nor U3207 (N_3207,N_2776,N_2257);
and U3208 (N_3208,N_2946,N_2216);
and U3209 (N_3209,N_2787,N_2666);
nand U3210 (N_3210,N_2983,N_2748);
nor U3211 (N_3211,N_2833,N_2771);
nor U3212 (N_3212,N_2123,N_2203);
or U3213 (N_3213,N_2211,N_2397);
and U3214 (N_3214,N_2356,N_2683);
nor U3215 (N_3215,N_2288,N_2070);
or U3216 (N_3216,N_2117,N_2987);
nand U3217 (N_3217,N_2977,N_2523);
nand U3218 (N_3218,N_2294,N_2852);
nor U3219 (N_3219,N_2420,N_2980);
and U3220 (N_3220,N_2119,N_2324);
nor U3221 (N_3221,N_2734,N_2828);
or U3222 (N_3222,N_2097,N_2017);
or U3223 (N_3223,N_2742,N_2783);
or U3224 (N_3224,N_2521,N_2372);
nand U3225 (N_3225,N_2141,N_2460);
or U3226 (N_3226,N_2210,N_2271);
nand U3227 (N_3227,N_2381,N_2816);
and U3228 (N_3228,N_2504,N_2891);
nand U3229 (N_3229,N_2901,N_2564);
or U3230 (N_3230,N_2491,N_2259);
or U3231 (N_3231,N_2942,N_2638);
or U3232 (N_3232,N_2073,N_2599);
nor U3233 (N_3233,N_2452,N_2872);
nor U3234 (N_3234,N_2249,N_2492);
nand U3235 (N_3235,N_2361,N_2427);
nand U3236 (N_3236,N_2386,N_2808);
and U3237 (N_3237,N_2675,N_2009);
nand U3238 (N_3238,N_2466,N_2108);
nand U3239 (N_3239,N_2693,N_2125);
and U3240 (N_3240,N_2468,N_2148);
nand U3241 (N_3241,N_2979,N_2966);
nand U3242 (N_3242,N_2566,N_2669);
or U3243 (N_3243,N_2345,N_2595);
or U3244 (N_3244,N_2796,N_2972);
nor U3245 (N_3245,N_2511,N_2974);
and U3246 (N_3246,N_2717,N_2517);
and U3247 (N_3247,N_2152,N_2031);
and U3248 (N_3248,N_2431,N_2486);
and U3249 (N_3249,N_2346,N_2416);
nor U3250 (N_3250,N_2045,N_2316);
nand U3251 (N_3251,N_2764,N_2634);
nor U3252 (N_3252,N_2873,N_2355);
or U3253 (N_3253,N_2472,N_2185);
nor U3254 (N_3254,N_2394,N_2688);
nand U3255 (N_3255,N_2411,N_2615);
and U3256 (N_3256,N_2889,N_2892);
or U3257 (N_3257,N_2105,N_2063);
or U3258 (N_3258,N_2969,N_2455);
and U3259 (N_3259,N_2298,N_2077);
nand U3260 (N_3260,N_2181,N_2430);
nand U3261 (N_3261,N_2506,N_2549);
or U3262 (N_3262,N_2328,N_2835);
and U3263 (N_3263,N_2032,N_2910);
and U3264 (N_3264,N_2184,N_2363);
or U3265 (N_3265,N_2439,N_2107);
or U3266 (N_3266,N_2534,N_2362);
nor U3267 (N_3267,N_2807,N_2888);
and U3268 (N_3268,N_2647,N_2863);
nor U3269 (N_3269,N_2544,N_2508);
nand U3270 (N_3270,N_2501,N_2617);
nor U3271 (N_3271,N_2244,N_2897);
nor U3272 (N_3272,N_2213,N_2598);
nor U3273 (N_3273,N_2450,N_2040);
nor U3274 (N_3274,N_2672,N_2786);
nand U3275 (N_3275,N_2827,N_2705);
and U3276 (N_3276,N_2868,N_2653);
nand U3277 (N_3277,N_2166,N_2219);
nor U3278 (N_3278,N_2707,N_2718);
nand U3279 (N_3279,N_2723,N_2422);
or U3280 (N_3280,N_2309,N_2269);
or U3281 (N_3281,N_2550,N_2369);
nor U3282 (N_3282,N_2195,N_2475);
or U3283 (N_3283,N_2671,N_2542);
nor U3284 (N_3284,N_2192,N_2906);
or U3285 (N_3285,N_2085,N_2632);
nand U3286 (N_3286,N_2722,N_2276);
or U3287 (N_3287,N_2605,N_2716);
and U3288 (N_3288,N_2162,N_2129);
nand U3289 (N_3289,N_2357,N_2687);
nor U3290 (N_3290,N_2410,N_2997);
nand U3291 (N_3291,N_2541,N_2680);
nand U3292 (N_3292,N_2135,N_2376);
or U3293 (N_3293,N_2058,N_2894);
nand U3294 (N_3294,N_2557,N_2727);
and U3295 (N_3295,N_2752,N_2281);
nor U3296 (N_3296,N_2293,N_2256);
nand U3297 (N_3297,N_2921,N_2823);
and U3298 (N_3298,N_2029,N_2594);
and U3299 (N_3299,N_2711,N_2079);
or U3300 (N_3300,N_2953,N_2778);
or U3301 (N_3301,N_2458,N_2437);
and U3302 (N_3302,N_2375,N_2613);
nand U3303 (N_3303,N_2995,N_2982);
or U3304 (N_3304,N_2440,N_2961);
nand U3305 (N_3305,N_2335,N_2793);
nand U3306 (N_3306,N_2319,N_2168);
and U3307 (N_3307,N_2654,N_2587);
nor U3308 (N_3308,N_2777,N_2155);
or U3309 (N_3309,N_2066,N_2957);
nor U3310 (N_3310,N_2763,N_2023);
nand U3311 (N_3311,N_2128,N_2297);
nand U3312 (N_3312,N_2649,N_2338);
and U3313 (N_3313,N_2415,N_2443);
or U3314 (N_3314,N_2641,N_2733);
nand U3315 (N_3315,N_2584,N_2663);
nor U3316 (N_3316,N_2830,N_2668);
nor U3317 (N_3317,N_2406,N_2146);
nor U3318 (N_3318,N_2445,N_2758);
or U3319 (N_3319,N_2788,N_2499);
or U3320 (N_3320,N_2915,N_2280);
nor U3321 (N_3321,N_2799,N_2876);
or U3322 (N_3322,N_2578,N_2189);
and U3323 (N_3323,N_2806,N_2604);
and U3324 (N_3324,N_2690,N_2234);
nand U3325 (N_3325,N_2952,N_2623);
nand U3326 (N_3326,N_2144,N_2960);
or U3327 (N_3327,N_2478,N_2327);
or U3328 (N_3328,N_2860,N_2967);
nand U3329 (N_3329,N_2469,N_2925);
nor U3330 (N_3330,N_2011,N_2350);
and U3331 (N_3331,N_2626,N_2756);
nand U3332 (N_3332,N_2260,N_2924);
and U3333 (N_3333,N_2618,N_2116);
and U3334 (N_3334,N_2754,N_2176);
or U3335 (N_3335,N_2780,N_2307);
and U3336 (N_3336,N_2251,N_2884);
or U3337 (N_3337,N_2174,N_2292);
nor U3338 (N_3338,N_2565,N_2451);
nand U3339 (N_3339,N_2143,N_2838);
and U3340 (N_3340,N_2999,N_2237);
and U3341 (N_3341,N_2692,N_2551);
nor U3342 (N_3342,N_2060,N_2836);
or U3343 (N_3343,N_2180,N_2110);
nand U3344 (N_3344,N_2627,N_2619);
or U3345 (N_3345,N_2024,N_2529);
nand U3346 (N_3346,N_2913,N_2713);
nand U3347 (N_3347,N_2660,N_2540);
nor U3348 (N_3348,N_2695,N_2667);
nor U3349 (N_3349,N_2332,N_2538);
nand U3350 (N_3350,N_2457,N_2630);
nor U3351 (N_3351,N_2648,N_2317);
or U3352 (N_3352,N_2263,N_2461);
and U3353 (N_3353,N_2875,N_2358);
and U3354 (N_3354,N_2197,N_2810);
nor U3355 (N_3355,N_2408,N_2526);
nand U3356 (N_3356,N_2992,N_2698);
or U3357 (N_3357,N_2826,N_2531);
or U3358 (N_3358,N_2854,N_2951);
nand U3359 (N_3359,N_2220,N_2080);
and U3360 (N_3360,N_2464,N_2432);
nand U3361 (N_3361,N_2659,N_2769);
and U3362 (N_3362,N_2905,N_2745);
xnor U3363 (N_3363,N_2981,N_2382);
xnor U3364 (N_3364,N_2035,N_2696);
nor U3365 (N_3365,N_2849,N_2726);
or U3366 (N_3366,N_2819,N_2537);
nor U3367 (N_3367,N_2735,N_2286);
or U3368 (N_3368,N_2932,N_2265);
nor U3369 (N_3369,N_2399,N_2724);
and U3370 (N_3370,N_2920,N_2178);
or U3371 (N_3371,N_2625,N_2814);
nand U3372 (N_3372,N_2371,N_2715);
nand U3373 (N_3373,N_2614,N_2585);
or U3374 (N_3374,N_2409,N_2130);
and U3375 (N_3375,N_2493,N_2067);
and U3376 (N_3376,N_2867,N_2899);
nand U3377 (N_3377,N_2964,N_2217);
nor U3378 (N_3378,N_2555,N_2851);
nor U3379 (N_3379,N_2048,N_2567);
and U3380 (N_3380,N_2284,N_2173);
nor U3381 (N_3381,N_2059,N_2102);
and U3382 (N_3382,N_2738,N_2919);
nand U3383 (N_3383,N_2142,N_2645);
or U3384 (N_3384,N_2866,N_2296);
or U3385 (N_3385,N_2673,N_2133);
xor U3386 (N_3386,N_2247,N_2488);
nor U3387 (N_3387,N_2283,N_2520);
nor U3388 (N_3388,N_2287,N_2909);
or U3389 (N_3389,N_2575,N_2597);
or U3390 (N_3390,N_2224,N_2299);
nand U3391 (N_3391,N_2069,N_2701);
nor U3392 (N_3392,N_2161,N_2360);
nor U3393 (N_3393,N_2145,N_2510);
and U3394 (N_3394,N_2865,N_2518);
and U3395 (N_3395,N_2183,N_2528);
or U3396 (N_3396,N_2911,N_2112);
nor U3397 (N_3397,N_2021,N_2051);
nand U3398 (N_3398,N_2633,N_2056);
nor U3399 (N_3399,N_2320,N_2755);
nor U3400 (N_3400,N_2963,N_2322);
nor U3401 (N_3401,N_2094,N_2885);
nand U3402 (N_3402,N_2252,N_2436);
or U3403 (N_3403,N_2871,N_2489);
nor U3404 (N_3404,N_2933,N_2086);
and U3405 (N_3405,N_2622,N_2325);
nor U3406 (N_3406,N_2138,N_2100);
nor U3407 (N_3407,N_2400,N_2041);
nand U3408 (N_3408,N_2404,N_2187);
and U3409 (N_3409,N_2495,N_2973);
nand U3410 (N_3410,N_2171,N_2559);
nor U3411 (N_3411,N_2471,N_2547);
and U3412 (N_3412,N_2678,N_2527);
and U3413 (N_3413,N_2229,N_2782);
and U3414 (N_3414,N_2025,N_2190);
nor U3415 (N_3415,N_2824,N_2607);
nor U3416 (N_3416,N_2923,N_2267);
nor U3417 (N_3417,N_2801,N_2334);
or U3418 (N_3418,N_2474,N_2201);
or U3419 (N_3419,N_2250,N_2702);
nand U3420 (N_3420,N_2384,N_2206);
nor U3421 (N_3421,N_2413,N_2862);
or U3422 (N_3422,N_2414,N_2740);
and U3423 (N_3423,N_2821,N_2577);
nand U3424 (N_3424,N_2562,N_2532);
nand U3425 (N_3425,N_2710,N_2467);
nand U3426 (N_3426,N_2785,N_2344);
and U3427 (N_3427,N_2347,N_2870);
nor U3428 (N_3428,N_2847,N_2340);
nand U3429 (N_3429,N_2380,N_2090);
and U3430 (N_3430,N_2610,N_2749);
and U3431 (N_3431,N_2277,N_2367);
and U3432 (N_3432,N_2637,N_2379);
or U3433 (N_3433,N_2278,N_2448);
and U3434 (N_3434,N_2074,N_2706);
or U3435 (N_3435,N_2333,N_2928);
nand U3436 (N_3436,N_2258,N_2841);
nand U3437 (N_3437,N_2028,N_2631);
or U3438 (N_3438,N_2525,N_2153);
or U3439 (N_3439,N_2121,N_2522);
or U3440 (N_3440,N_2000,N_2421);
and U3441 (N_3441,N_2588,N_2456);
nand U3442 (N_3442,N_2274,N_2065);
or U3443 (N_3443,N_2020,N_2095);
and U3444 (N_3444,N_2580,N_2497);
nand U3445 (N_3445,N_2760,N_2136);
and U3446 (N_3446,N_2481,N_2150);
nand U3447 (N_3447,N_2487,N_2370);
nand U3448 (N_3448,N_2881,N_2013);
and U3449 (N_3449,N_2986,N_2761);
and U3450 (N_3450,N_2890,N_2212);
nand U3451 (N_3451,N_2321,N_2535);
nor U3452 (N_3452,N_2193,N_2010);
or U3453 (N_3453,N_2941,N_2435);
xnor U3454 (N_3454,N_2246,N_2708);
nand U3455 (N_3455,N_2620,N_2996);
nand U3456 (N_3456,N_2877,N_2062);
nor U3457 (N_3457,N_2616,N_2624);
and U3458 (N_3458,N_2275,N_2664);
or U3459 (N_3459,N_2556,N_2750);
and U3460 (N_3460,N_2651,N_2157);
or U3461 (N_3461,N_2364,N_2697);
nor U3462 (N_3462,N_2300,N_2677);
and U3463 (N_3463,N_2874,N_2412);
or U3464 (N_3464,N_2989,N_2583);
nand U3465 (N_3465,N_2887,N_2221);
nor U3466 (N_3466,N_2800,N_2053);
or U3467 (N_3467,N_2424,N_2791);
or U3468 (N_3468,N_2956,N_2182);
or U3469 (N_3469,N_2339,N_2665);
nand U3470 (N_3470,N_2366,N_2943);
and U3471 (N_3471,N_2268,N_2306);
nand U3472 (N_3472,N_2568,N_2245);
nor U3473 (N_3473,N_2712,N_2272);
nand U3474 (N_3474,N_2207,N_2970);
nand U3475 (N_3475,N_2462,N_2797);
and U3476 (N_3476,N_2579,N_2194);
or U3477 (N_3477,N_2676,N_2684);
and U3478 (N_3478,N_2154,N_2329);
and U3479 (N_3479,N_2270,N_2177);
nand U3480 (N_3480,N_2842,N_2401);
and U3481 (N_3481,N_2477,N_2940);
and U3482 (N_3482,N_2700,N_2839);
nand U3483 (N_3483,N_2044,N_2743);
nand U3484 (N_3484,N_2790,N_2878);
nor U3485 (N_3485,N_2789,N_2719);
nor U3486 (N_3486,N_2026,N_2907);
nor U3487 (N_3487,N_2930,N_2109);
and U3488 (N_3488,N_2962,N_2539);
or U3489 (N_3489,N_2465,N_2589);
and U3490 (N_3490,N_2912,N_2248);
nor U3491 (N_3491,N_2463,N_2103);
or U3492 (N_3492,N_2730,N_2301);
nor U3493 (N_3493,N_2313,N_2832);
nand U3494 (N_3494,N_2536,N_2124);
nand U3495 (N_3495,N_2419,N_2590);
nor U3496 (N_3496,N_2057,N_2558);
nor U3497 (N_3497,N_2285,N_2978);
or U3498 (N_3498,N_2524,N_2861);
nand U3499 (N_3499,N_2837,N_2395);
nand U3500 (N_3500,N_2913,N_2937);
and U3501 (N_3501,N_2914,N_2210);
or U3502 (N_3502,N_2259,N_2014);
and U3503 (N_3503,N_2659,N_2111);
and U3504 (N_3504,N_2932,N_2972);
or U3505 (N_3505,N_2317,N_2600);
nor U3506 (N_3506,N_2977,N_2173);
nand U3507 (N_3507,N_2415,N_2120);
nor U3508 (N_3508,N_2776,N_2488);
nor U3509 (N_3509,N_2434,N_2500);
nand U3510 (N_3510,N_2649,N_2261);
nand U3511 (N_3511,N_2744,N_2829);
nor U3512 (N_3512,N_2882,N_2143);
and U3513 (N_3513,N_2194,N_2113);
and U3514 (N_3514,N_2244,N_2012);
and U3515 (N_3515,N_2235,N_2675);
nand U3516 (N_3516,N_2303,N_2590);
or U3517 (N_3517,N_2474,N_2758);
and U3518 (N_3518,N_2156,N_2961);
nand U3519 (N_3519,N_2743,N_2082);
nor U3520 (N_3520,N_2433,N_2671);
or U3521 (N_3521,N_2025,N_2405);
nor U3522 (N_3522,N_2088,N_2837);
nor U3523 (N_3523,N_2598,N_2610);
nor U3524 (N_3524,N_2707,N_2183);
nor U3525 (N_3525,N_2150,N_2086);
nor U3526 (N_3526,N_2375,N_2179);
nor U3527 (N_3527,N_2683,N_2817);
nor U3528 (N_3528,N_2953,N_2076);
nor U3529 (N_3529,N_2945,N_2992);
or U3530 (N_3530,N_2020,N_2172);
and U3531 (N_3531,N_2160,N_2920);
nor U3532 (N_3532,N_2012,N_2501);
nor U3533 (N_3533,N_2143,N_2960);
or U3534 (N_3534,N_2623,N_2616);
nand U3535 (N_3535,N_2728,N_2172);
or U3536 (N_3536,N_2714,N_2267);
nor U3537 (N_3537,N_2795,N_2741);
nand U3538 (N_3538,N_2724,N_2474);
nor U3539 (N_3539,N_2493,N_2854);
and U3540 (N_3540,N_2848,N_2747);
and U3541 (N_3541,N_2006,N_2217);
nand U3542 (N_3542,N_2756,N_2803);
nand U3543 (N_3543,N_2948,N_2731);
or U3544 (N_3544,N_2022,N_2924);
and U3545 (N_3545,N_2446,N_2223);
or U3546 (N_3546,N_2489,N_2585);
and U3547 (N_3547,N_2512,N_2743);
nor U3548 (N_3548,N_2652,N_2999);
nand U3549 (N_3549,N_2132,N_2060);
nand U3550 (N_3550,N_2536,N_2065);
nand U3551 (N_3551,N_2374,N_2549);
or U3552 (N_3552,N_2141,N_2665);
nor U3553 (N_3553,N_2744,N_2946);
and U3554 (N_3554,N_2070,N_2548);
or U3555 (N_3555,N_2574,N_2575);
and U3556 (N_3556,N_2710,N_2867);
nor U3557 (N_3557,N_2889,N_2962);
and U3558 (N_3558,N_2604,N_2404);
and U3559 (N_3559,N_2562,N_2612);
nand U3560 (N_3560,N_2378,N_2578);
and U3561 (N_3561,N_2302,N_2281);
nor U3562 (N_3562,N_2227,N_2020);
nand U3563 (N_3563,N_2202,N_2173);
nand U3564 (N_3564,N_2690,N_2000);
nand U3565 (N_3565,N_2131,N_2356);
or U3566 (N_3566,N_2082,N_2483);
nand U3567 (N_3567,N_2817,N_2156);
nand U3568 (N_3568,N_2330,N_2293);
and U3569 (N_3569,N_2222,N_2465);
nor U3570 (N_3570,N_2526,N_2574);
or U3571 (N_3571,N_2023,N_2580);
and U3572 (N_3572,N_2898,N_2633);
or U3573 (N_3573,N_2909,N_2915);
or U3574 (N_3574,N_2151,N_2223);
xor U3575 (N_3575,N_2543,N_2746);
nor U3576 (N_3576,N_2736,N_2103);
nand U3577 (N_3577,N_2860,N_2940);
nor U3578 (N_3578,N_2145,N_2983);
and U3579 (N_3579,N_2484,N_2240);
nand U3580 (N_3580,N_2637,N_2046);
nor U3581 (N_3581,N_2995,N_2169);
nand U3582 (N_3582,N_2823,N_2315);
or U3583 (N_3583,N_2323,N_2390);
or U3584 (N_3584,N_2912,N_2887);
and U3585 (N_3585,N_2966,N_2056);
xnor U3586 (N_3586,N_2053,N_2294);
and U3587 (N_3587,N_2147,N_2203);
nor U3588 (N_3588,N_2076,N_2720);
or U3589 (N_3589,N_2076,N_2613);
or U3590 (N_3590,N_2743,N_2478);
nor U3591 (N_3591,N_2911,N_2208);
nand U3592 (N_3592,N_2836,N_2860);
nor U3593 (N_3593,N_2582,N_2216);
xor U3594 (N_3594,N_2392,N_2022);
or U3595 (N_3595,N_2811,N_2270);
nand U3596 (N_3596,N_2019,N_2815);
or U3597 (N_3597,N_2646,N_2561);
nand U3598 (N_3598,N_2079,N_2436);
and U3599 (N_3599,N_2085,N_2922);
xnor U3600 (N_3600,N_2594,N_2743);
nor U3601 (N_3601,N_2258,N_2114);
or U3602 (N_3602,N_2163,N_2604);
nand U3603 (N_3603,N_2270,N_2762);
or U3604 (N_3604,N_2339,N_2097);
nand U3605 (N_3605,N_2630,N_2626);
and U3606 (N_3606,N_2346,N_2415);
nor U3607 (N_3607,N_2811,N_2136);
nor U3608 (N_3608,N_2057,N_2898);
nand U3609 (N_3609,N_2965,N_2632);
and U3610 (N_3610,N_2712,N_2943);
or U3611 (N_3611,N_2423,N_2578);
or U3612 (N_3612,N_2829,N_2836);
nor U3613 (N_3613,N_2832,N_2449);
nor U3614 (N_3614,N_2714,N_2599);
nor U3615 (N_3615,N_2219,N_2345);
and U3616 (N_3616,N_2148,N_2795);
and U3617 (N_3617,N_2138,N_2584);
or U3618 (N_3618,N_2014,N_2431);
nor U3619 (N_3619,N_2281,N_2015);
and U3620 (N_3620,N_2270,N_2347);
or U3621 (N_3621,N_2753,N_2097);
and U3622 (N_3622,N_2820,N_2008);
or U3623 (N_3623,N_2183,N_2817);
nand U3624 (N_3624,N_2830,N_2172);
nand U3625 (N_3625,N_2777,N_2701);
and U3626 (N_3626,N_2958,N_2889);
nor U3627 (N_3627,N_2622,N_2198);
nand U3628 (N_3628,N_2730,N_2723);
nor U3629 (N_3629,N_2928,N_2946);
or U3630 (N_3630,N_2804,N_2096);
nand U3631 (N_3631,N_2471,N_2731);
and U3632 (N_3632,N_2700,N_2330);
nor U3633 (N_3633,N_2430,N_2169);
nand U3634 (N_3634,N_2576,N_2352);
or U3635 (N_3635,N_2087,N_2358);
nor U3636 (N_3636,N_2899,N_2379);
nor U3637 (N_3637,N_2155,N_2393);
and U3638 (N_3638,N_2887,N_2350);
or U3639 (N_3639,N_2783,N_2195);
nor U3640 (N_3640,N_2487,N_2911);
nand U3641 (N_3641,N_2531,N_2053);
or U3642 (N_3642,N_2166,N_2546);
or U3643 (N_3643,N_2074,N_2143);
and U3644 (N_3644,N_2511,N_2369);
and U3645 (N_3645,N_2377,N_2043);
nor U3646 (N_3646,N_2634,N_2516);
nor U3647 (N_3647,N_2194,N_2777);
and U3648 (N_3648,N_2106,N_2140);
and U3649 (N_3649,N_2398,N_2803);
nand U3650 (N_3650,N_2915,N_2462);
or U3651 (N_3651,N_2148,N_2139);
nor U3652 (N_3652,N_2901,N_2761);
nand U3653 (N_3653,N_2605,N_2745);
or U3654 (N_3654,N_2015,N_2796);
or U3655 (N_3655,N_2890,N_2980);
or U3656 (N_3656,N_2778,N_2606);
nand U3657 (N_3657,N_2052,N_2123);
or U3658 (N_3658,N_2123,N_2226);
and U3659 (N_3659,N_2590,N_2416);
nand U3660 (N_3660,N_2191,N_2916);
nand U3661 (N_3661,N_2162,N_2283);
nand U3662 (N_3662,N_2784,N_2882);
or U3663 (N_3663,N_2018,N_2422);
and U3664 (N_3664,N_2664,N_2927);
and U3665 (N_3665,N_2312,N_2602);
xnor U3666 (N_3666,N_2487,N_2444);
nand U3667 (N_3667,N_2274,N_2569);
and U3668 (N_3668,N_2304,N_2291);
or U3669 (N_3669,N_2876,N_2625);
and U3670 (N_3670,N_2051,N_2795);
and U3671 (N_3671,N_2932,N_2868);
or U3672 (N_3672,N_2286,N_2697);
nor U3673 (N_3673,N_2528,N_2298);
and U3674 (N_3674,N_2780,N_2026);
nor U3675 (N_3675,N_2962,N_2608);
or U3676 (N_3676,N_2154,N_2404);
and U3677 (N_3677,N_2242,N_2854);
nand U3678 (N_3678,N_2336,N_2297);
nor U3679 (N_3679,N_2398,N_2840);
nand U3680 (N_3680,N_2830,N_2242);
or U3681 (N_3681,N_2156,N_2035);
or U3682 (N_3682,N_2499,N_2564);
or U3683 (N_3683,N_2396,N_2713);
and U3684 (N_3684,N_2436,N_2827);
or U3685 (N_3685,N_2574,N_2249);
nand U3686 (N_3686,N_2075,N_2900);
nor U3687 (N_3687,N_2321,N_2127);
and U3688 (N_3688,N_2825,N_2889);
nor U3689 (N_3689,N_2959,N_2660);
nand U3690 (N_3690,N_2316,N_2747);
or U3691 (N_3691,N_2214,N_2921);
and U3692 (N_3692,N_2818,N_2496);
nor U3693 (N_3693,N_2972,N_2904);
nor U3694 (N_3694,N_2448,N_2017);
and U3695 (N_3695,N_2416,N_2316);
or U3696 (N_3696,N_2532,N_2588);
and U3697 (N_3697,N_2887,N_2629);
or U3698 (N_3698,N_2748,N_2439);
nand U3699 (N_3699,N_2801,N_2043);
or U3700 (N_3700,N_2852,N_2819);
nor U3701 (N_3701,N_2855,N_2413);
nand U3702 (N_3702,N_2739,N_2714);
or U3703 (N_3703,N_2802,N_2519);
or U3704 (N_3704,N_2996,N_2863);
and U3705 (N_3705,N_2455,N_2231);
nand U3706 (N_3706,N_2876,N_2043);
or U3707 (N_3707,N_2244,N_2658);
or U3708 (N_3708,N_2227,N_2330);
nand U3709 (N_3709,N_2322,N_2000);
nor U3710 (N_3710,N_2110,N_2595);
and U3711 (N_3711,N_2742,N_2907);
or U3712 (N_3712,N_2149,N_2939);
nor U3713 (N_3713,N_2197,N_2256);
nand U3714 (N_3714,N_2402,N_2013);
nand U3715 (N_3715,N_2680,N_2761);
and U3716 (N_3716,N_2002,N_2734);
nand U3717 (N_3717,N_2677,N_2137);
nand U3718 (N_3718,N_2055,N_2335);
or U3719 (N_3719,N_2385,N_2686);
nor U3720 (N_3720,N_2940,N_2795);
or U3721 (N_3721,N_2316,N_2428);
nor U3722 (N_3722,N_2570,N_2697);
nand U3723 (N_3723,N_2454,N_2998);
and U3724 (N_3724,N_2584,N_2668);
nand U3725 (N_3725,N_2961,N_2283);
or U3726 (N_3726,N_2716,N_2161);
and U3727 (N_3727,N_2692,N_2200);
or U3728 (N_3728,N_2606,N_2919);
and U3729 (N_3729,N_2834,N_2449);
and U3730 (N_3730,N_2858,N_2416);
and U3731 (N_3731,N_2017,N_2123);
nand U3732 (N_3732,N_2573,N_2481);
or U3733 (N_3733,N_2076,N_2503);
nand U3734 (N_3734,N_2491,N_2539);
nor U3735 (N_3735,N_2466,N_2025);
and U3736 (N_3736,N_2496,N_2126);
or U3737 (N_3737,N_2261,N_2951);
nand U3738 (N_3738,N_2669,N_2705);
or U3739 (N_3739,N_2159,N_2954);
nand U3740 (N_3740,N_2595,N_2739);
and U3741 (N_3741,N_2787,N_2933);
nand U3742 (N_3742,N_2318,N_2033);
nand U3743 (N_3743,N_2779,N_2752);
nand U3744 (N_3744,N_2700,N_2531);
and U3745 (N_3745,N_2247,N_2828);
nand U3746 (N_3746,N_2264,N_2793);
and U3747 (N_3747,N_2613,N_2801);
and U3748 (N_3748,N_2197,N_2790);
and U3749 (N_3749,N_2824,N_2065);
and U3750 (N_3750,N_2509,N_2029);
or U3751 (N_3751,N_2158,N_2968);
or U3752 (N_3752,N_2724,N_2953);
or U3753 (N_3753,N_2646,N_2489);
and U3754 (N_3754,N_2404,N_2125);
nor U3755 (N_3755,N_2028,N_2085);
or U3756 (N_3756,N_2670,N_2694);
nand U3757 (N_3757,N_2135,N_2210);
or U3758 (N_3758,N_2335,N_2647);
or U3759 (N_3759,N_2845,N_2868);
or U3760 (N_3760,N_2051,N_2684);
nand U3761 (N_3761,N_2422,N_2575);
and U3762 (N_3762,N_2687,N_2141);
and U3763 (N_3763,N_2896,N_2618);
or U3764 (N_3764,N_2375,N_2670);
and U3765 (N_3765,N_2301,N_2396);
and U3766 (N_3766,N_2315,N_2177);
or U3767 (N_3767,N_2201,N_2903);
nand U3768 (N_3768,N_2407,N_2093);
and U3769 (N_3769,N_2557,N_2842);
and U3770 (N_3770,N_2999,N_2025);
and U3771 (N_3771,N_2839,N_2670);
nor U3772 (N_3772,N_2590,N_2598);
nand U3773 (N_3773,N_2042,N_2044);
or U3774 (N_3774,N_2723,N_2934);
or U3775 (N_3775,N_2244,N_2646);
nor U3776 (N_3776,N_2580,N_2505);
nand U3777 (N_3777,N_2109,N_2706);
and U3778 (N_3778,N_2760,N_2830);
nor U3779 (N_3779,N_2860,N_2717);
nand U3780 (N_3780,N_2199,N_2634);
nor U3781 (N_3781,N_2464,N_2140);
nand U3782 (N_3782,N_2796,N_2762);
and U3783 (N_3783,N_2491,N_2393);
and U3784 (N_3784,N_2279,N_2173);
nor U3785 (N_3785,N_2770,N_2736);
or U3786 (N_3786,N_2183,N_2966);
nor U3787 (N_3787,N_2165,N_2904);
and U3788 (N_3788,N_2374,N_2221);
nor U3789 (N_3789,N_2943,N_2743);
nand U3790 (N_3790,N_2838,N_2439);
nand U3791 (N_3791,N_2949,N_2440);
and U3792 (N_3792,N_2394,N_2567);
nand U3793 (N_3793,N_2363,N_2850);
and U3794 (N_3794,N_2273,N_2626);
and U3795 (N_3795,N_2818,N_2618);
nor U3796 (N_3796,N_2204,N_2220);
or U3797 (N_3797,N_2656,N_2426);
and U3798 (N_3798,N_2462,N_2773);
nor U3799 (N_3799,N_2165,N_2413);
nor U3800 (N_3800,N_2051,N_2233);
and U3801 (N_3801,N_2792,N_2461);
nor U3802 (N_3802,N_2588,N_2604);
nand U3803 (N_3803,N_2558,N_2328);
nand U3804 (N_3804,N_2323,N_2643);
nor U3805 (N_3805,N_2237,N_2371);
or U3806 (N_3806,N_2902,N_2687);
and U3807 (N_3807,N_2066,N_2711);
nor U3808 (N_3808,N_2683,N_2850);
and U3809 (N_3809,N_2223,N_2099);
nand U3810 (N_3810,N_2783,N_2068);
nor U3811 (N_3811,N_2325,N_2510);
nand U3812 (N_3812,N_2269,N_2416);
and U3813 (N_3813,N_2087,N_2684);
nand U3814 (N_3814,N_2518,N_2786);
or U3815 (N_3815,N_2119,N_2674);
and U3816 (N_3816,N_2458,N_2433);
nor U3817 (N_3817,N_2080,N_2300);
or U3818 (N_3818,N_2191,N_2109);
or U3819 (N_3819,N_2276,N_2950);
and U3820 (N_3820,N_2834,N_2627);
or U3821 (N_3821,N_2282,N_2092);
nor U3822 (N_3822,N_2137,N_2155);
and U3823 (N_3823,N_2323,N_2706);
or U3824 (N_3824,N_2525,N_2596);
nor U3825 (N_3825,N_2948,N_2162);
nor U3826 (N_3826,N_2487,N_2302);
or U3827 (N_3827,N_2293,N_2566);
and U3828 (N_3828,N_2489,N_2621);
or U3829 (N_3829,N_2597,N_2872);
or U3830 (N_3830,N_2386,N_2319);
nand U3831 (N_3831,N_2877,N_2190);
nor U3832 (N_3832,N_2082,N_2341);
and U3833 (N_3833,N_2842,N_2794);
nand U3834 (N_3834,N_2437,N_2172);
or U3835 (N_3835,N_2636,N_2236);
or U3836 (N_3836,N_2300,N_2291);
nor U3837 (N_3837,N_2455,N_2066);
and U3838 (N_3838,N_2016,N_2870);
or U3839 (N_3839,N_2230,N_2248);
nand U3840 (N_3840,N_2606,N_2900);
nor U3841 (N_3841,N_2367,N_2782);
or U3842 (N_3842,N_2104,N_2315);
nor U3843 (N_3843,N_2223,N_2313);
or U3844 (N_3844,N_2821,N_2675);
and U3845 (N_3845,N_2129,N_2036);
nor U3846 (N_3846,N_2391,N_2168);
or U3847 (N_3847,N_2867,N_2996);
and U3848 (N_3848,N_2750,N_2889);
or U3849 (N_3849,N_2829,N_2014);
and U3850 (N_3850,N_2465,N_2346);
or U3851 (N_3851,N_2590,N_2732);
nor U3852 (N_3852,N_2004,N_2132);
or U3853 (N_3853,N_2862,N_2778);
or U3854 (N_3854,N_2183,N_2998);
or U3855 (N_3855,N_2196,N_2493);
nand U3856 (N_3856,N_2837,N_2794);
and U3857 (N_3857,N_2711,N_2766);
or U3858 (N_3858,N_2357,N_2941);
or U3859 (N_3859,N_2923,N_2753);
and U3860 (N_3860,N_2820,N_2723);
nand U3861 (N_3861,N_2440,N_2652);
and U3862 (N_3862,N_2846,N_2825);
nand U3863 (N_3863,N_2139,N_2671);
or U3864 (N_3864,N_2937,N_2442);
nor U3865 (N_3865,N_2398,N_2434);
and U3866 (N_3866,N_2655,N_2462);
nor U3867 (N_3867,N_2510,N_2628);
nor U3868 (N_3868,N_2805,N_2634);
or U3869 (N_3869,N_2927,N_2871);
nand U3870 (N_3870,N_2563,N_2209);
and U3871 (N_3871,N_2643,N_2595);
or U3872 (N_3872,N_2858,N_2554);
nand U3873 (N_3873,N_2025,N_2541);
nor U3874 (N_3874,N_2345,N_2913);
and U3875 (N_3875,N_2791,N_2304);
and U3876 (N_3876,N_2223,N_2782);
and U3877 (N_3877,N_2079,N_2424);
xor U3878 (N_3878,N_2021,N_2938);
or U3879 (N_3879,N_2732,N_2243);
or U3880 (N_3880,N_2267,N_2206);
nand U3881 (N_3881,N_2747,N_2617);
and U3882 (N_3882,N_2045,N_2845);
or U3883 (N_3883,N_2551,N_2654);
or U3884 (N_3884,N_2113,N_2298);
and U3885 (N_3885,N_2991,N_2616);
or U3886 (N_3886,N_2213,N_2693);
nor U3887 (N_3887,N_2285,N_2363);
or U3888 (N_3888,N_2527,N_2627);
nand U3889 (N_3889,N_2348,N_2285);
nor U3890 (N_3890,N_2834,N_2825);
and U3891 (N_3891,N_2289,N_2629);
and U3892 (N_3892,N_2135,N_2527);
nor U3893 (N_3893,N_2553,N_2353);
nand U3894 (N_3894,N_2778,N_2612);
and U3895 (N_3895,N_2910,N_2047);
and U3896 (N_3896,N_2240,N_2849);
or U3897 (N_3897,N_2572,N_2157);
or U3898 (N_3898,N_2448,N_2354);
and U3899 (N_3899,N_2592,N_2805);
nand U3900 (N_3900,N_2680,N_2304);
and U3901 (N_3901,N_2299,N_2092);
nor U3902 (N_3902,N_2001,N_2532);
nor U3903 (N_3903,N_2718,N_2686);
and U3904 (N_3904,N_2975,N_2445);
xnor U3905 (N_3905,N_2024,N_2916);
and U3906 (N_3906,N_2199,N_2982);
nor U3907 (N_3907,N_2336,N_2519);
and U3908 (N_3908,N_2138,N_2161);
nand U3909 (N_3909,N_2519,N_2663);
nand U3910 (N_3910,N_2224,N_2676);
or U3911 (N_3911,N_2219,N_2098);
or U3912 (N_3912,N_2243,N_2367);
or U3913 (N_3913,N_2654,N_2087);
or U3914 (N_3914,N_2829,N_2184);
nand U3915 (N_3915,N_2154,N_2675);
or U3916 (N_3916,N_2409,N_2398);
and U3917 (N_3917,N_2810,N_2513);
or U3918 (N_3918,N_2592,N_2898);
nand U3919 (N_3919,N_2836,N_2325);
or U3920 (N_3920,N_2541,N_2359);
and U3921 (N_3921,N_2101,N_2059);
and U3922 (N_3922,N_2006,N_2753);
and U3923 (N_3923,N_2369,N_2903);
nor U3924 (N_3924,N_2616,N_2004);
and U3925 (N_3925,N_2454,N_2299);
nand U3926 (N_3926,N_2224,N_2292);
and U3927 (N_3927,N_2344,N_2106);
and U3928 (N_3928,N_2646,N_2730);
and U3929 (N_3929,N_2019,N_2630);
and U3930 (N_3930,N_2326,N_2603);
nor U3931 (N_3931,N_2896,N_2563);
nand U3932 (N_3932,N_2167,N_2557);
nand U3933 (N_3933,N_2653,N_2379);
nor U3934 (N_3934,N_2450,N_2995);
or U3935 (N_3935,N_2923,N_2958);
and U3936 (N_3936,N_2579,N_2859);
or U3937 (N_3937,N_2024,N_2216);
nand U3938 (N_3938,N_2392,N_2930);
and U3939 (N_3939,N_2063,N_2357);
and U3940 (N_3940,N_2503,N_2320);
nor U3941 (N_3941,N_2334,N_2950);
nand U3942 (N_3942,N_2806,N_2464);
nand U3943 (N_3943,N_2415,N_2075);
and U3944 (N_3944,N_2346,N_2002);
nor U3945 (N_3945,N_2734,N_2351);
nand U3946 (N_3946,N_2976,N_2668);
and U3947 (N_3947,N_2134,N_2533);
or U3948 (N_3948,N_2340,N_2438);
and U3949 (N_3949,N_2817,N_2977);
and U3950 (N_3950,N_2126,N_2836);
nor U3951 (N_3951,N_2661,N_2795);
or U3952 (N_3952,N_2205,N_2044);
nor U3953 (N_3953,N_2265,N_2257);
and U3954 (N_3954,N_2876,N_2649);
and U3955 (N_3955,N_2498,N_2227);
or U3956 (N_3956,N_2707,N_2396);
nand U3957 (N_3957,N_2225,N_2706);
nor U3958 (N_3958,N_2721,N_2073);
nor U3959 (N_3959,N_2939,N_2248);
nor U3960 (N_3960,N_2966,N_2693);
and U3961 (N_3961,N_2018,N_2509);
nor U3962 (N_3962,N_2713,N_2035);
nor U3963 (N_3963,N_2222,N_2044);
nand U3964 (N_3964,N_2757,N_2855);
nand U3965 (N_3965,N_2337,N_2755);
nand U3966 (N_3966,N_2746,N_2555);
or U3967 (N_3967,N_2812,N_2764);
and U3968 (N_3968,N_2513,N_2686);
and U3969 (N_3969,N_2591,N_2472);
or U3970 (N_3970,N_2464,N_2380);
and U3971 (N_3971,N_2110,N_2031);
or U3972 (N_3972,N_2867,N_2910);
nand U3973 (N_3973,N_2074,N_2484);
and U3974 (N_3974,N_2195,N_2016);
nand U3975 (N_3975,N_2007,N_2901);
or U3976 (N_3976,N_2134,N_2722);
or U3977 (N_3977,N_2444,N_2042);
and U3978 (N_3978,N_2930,N_2061);
or U3979 (N_3979,N_2671,N_2985);
or U3980 (N_3980,N_2087,N_2549);
and U3981 (N_3981,N_2192,N_2033);
or U3982 (N_3982,N_2329,N_2184);
and U3983 (N_3983,N_2255,N_2008);
nor U3984 (N_3984,N_2874,N_2687);
or U3985 (N_3985,N_2739,N_2339);
or U3986 (N_3986,N_2129,N_2742);
nor U3987 (N_3987,N_2415,N_2826);
and U3988 (N_3988,N_2828,N_2423);
or U3989 (N_3989,N_2224,N_2945);
nor U3990 (N_3990,N_2327,N_2723);
nand U3991 (N_3991,N_2093,N_2441);
and U3992 (N_3992,N_2959,N_2586);
nor U3993 (N_3993,N_2788,N_2580);
or U3994 (N_3994,N_2222,N_2198);
or U3995 (N_3995,N_2140,N_2637);
nor U3996 (N_3996,N_2573,N_2950);
nor U3997 (N_3997,N_2425,N_2051);
or U3998 (N_3998,N_2679,N_2379);
nand U3999 (N_3999,N_2465,N_2500);
or U4000 (N_4000,N_3312,N_3818);
nand U4001 (N_4001,N_3143,N_3166);
nor U4002 (N_4002,N_3007,N_3235);
or U4003 (N_4003,N_3656,N_3006);
and U4004 (N_4004,N_3853,N_3601);
nor U4005 (N_4005,N_3076,N_3699);
nand U4006 (N_4006,N_3282,N_3194);
nor U4007 (N_4007,N_3081,N_3281);
nor U4008 (N_4008,N_3942,N_3436);
or U4009 (N_4009,N_3617,N_3979);
nor U4010 (N_4010,N_3449,N_3239);
nand U4011 (N_4011,N_3990,N_3682);
or U4012 (N_4012,N_3987,N_3204);
nand U4013 (N_4013,N_3530,N_3623);
xnor U4014 (N_4014,N_3325,N_3876);
nor U4015 (N_4015,N_3859,N_3414);
or U4016 (N_4016,N_3430,N_3043);
nand U4017 (N_4017,N_3975,N_3273);
nor U4018 (N_4018,N_3776,N_3257);
nand U4019 (N_4019,N_3544,N_3680);
nor U4020 (N_4020,N_3778,N_3870);
nand U4021 (N_4021,N_3417,N_3574);
and U4022 (N_4022,N_3811,N_3802);
and U4023 (N_4023,N_3227,N_3265);
nor U4024 (N_4024,N_3666,N_3831);
or U4025 (N_4025,N_3063,N_3283);
nand U4026 (N_4026,N_3490,N_3170);
xor U4027 (N_4027,N_3279,N_3351);
nand U4028 (N_4028,N_3676,N_3982);
nand U4029 (N_4029,N_3340,N_3432);
or U4030 (N_4030,N_3499,N_3951);
nor U4031 (N_4031,N_3621,N_3613);
nand U4032 (N_4032,N_3952,N_3521);
and U4033 (N_4033,N_3764,N_3567);
nand U4034 (N_4034,N_3635,N_3415);
and U4035 (N_4035,N_3110,N_3927);
and U4036 (N_4036,N_3077,N_3503);
or U4037 (N_4037,N_3517,N_3010);
nor U4038 (N_4038,N_3736,N_3962);
nor U4039 (N_4039,N_3939,N_3577);
nand U4040 (N_4040,N_3959,N_3300);
nor U4041 (N_4041,N_3446,N_3406);
nand U4042 (N_4042,N_3518,N_3328);
and U4043 (N_4043,N_3657,N_3626);
nand U4044 (N_4044,N_3256,N_3700);
nand U4045 (N_4045,N_3379,N_3167);
nor U4046 (N_4046,N_3905,N_3153);
and U4047 (N_4047,N_3931,N_3899);
nor U4048 (N_4048,N_3375,N_3456);
xnor U4049 (N_4049,N_3228,N_3169);
nand U4050 (N_4050,N_3065,N_3485);
and U4051 (N_4051,N_3733,N_3610);
and U4052 (N_4052,N_3191,N_3690);
or U4053 (N_4053,N_3555,N_3286);
and U4054 (N_4054,N_3488,N_3923);
or U4055 (N_4055,N_3806,N_3426);
nand U4056 (N_4056,N_3599,N_3280);
or U4057 (N_4057,N_3024,N_3510);
and U4058 (N_4058,N_3096,N_3598);
xnor U4059 (N_4059,N_3374,N_3907);
or U4060 (N_4060,N_3856,N_3429);
nand U4061 (N_4061,N_3892,N_3726);
or U4062 (N_4062,N_3655,N_3968);
nor U4063 (N_4063,N_3121,N_3285);
nor U4064 (N_4064,N_3647,N_3674);
nand U4065 (N_4065,N_3612,N_3718);
or U4066 (N_4066,N_3304,N_3314);
or U4067 (N_4067,N_3734,N_3618);
or U4068 (N_4068,N_3398,N_3366);
nor U4069 (N_4069,N_3341,N_3537);
or U4070 (N_4070,N_3457,N_3898);
nand U4071 (N_4071,N_3493,N_3992);
nor U4072 (N_4072,N_3444,N_3837);
and U4073 (N_4073,N_3466,N_3478);
nand U4074 (N_4074,N_3134,N_3940);
nor U4075 (N_4075,N_3605,N_3335);
and U4076 (N_4076,N_3707,N_3452);
nor U4077 (N_4077,N_3247,N_3214);
or U4078 (N_4078,N_3423,N_3901);
nor U4079 (N_4079,N_3128,N_3721);
nand U4080 (N_4080,N_3402,N_3483);
nand U4081 (N_4081,N_3703,N_3439);
nor U4082 (N_4082,N_3342,N_3506);
and U4083 (N_4083,N_3048,N_3346);
nor U4084 (N_4084,N_3701,N_3221);
and U4085 (N_4085,N_3047,N_3269);
or U4086 (N_4086,N_3683,N_3288);
nor U4087 (N_4087,N_3516,N_3232);
nor U4088 (N_4088,N_3814,N_3509);
and U4089 (N_4089,N_3039,N_3447);
or U4090 (N_4090,N_3135,N_3477);
nor U4091 (N_4091,N_3332,N_3897);
nor U4092 (N_4092,N_3357,N_3889);
and U4093 (N_4093,N_3427,N_3860);
nand U4094 (N_4094,N_3428,N_3089);
nor U4095 (N_4095,N_3763,N_3264);
and U4096 (N_4096,N_3309,N_3155);
or U4097 (N_4097,N_3720,N_3461);
nor U4098 (N_4098,N_3099,N_3413);
nand U4099 (N_4099,N_3482,N_3162);
and U4100 (N_4100,N_3958,N_3592);
nor U4101 (N_4101,N_3520,N_3200);
nand U4102 (N_4102,N_3715,N_3971);
xor U4103 (N_4103,N_3476,N_3714);
and U4104 (N_4104,N_3513,N_3393);
and U4105 (N_4105,N_3753,N_3526);
nand U4106 (N_4106,N_3885,N_3215);
and U4107 (N_4107,N_3536,N_3179);
and U4108 (N_4108,N_3359,N_3389);
nand U4109 (N_4109,N_3563,N_3038);
and U4110 (N_4110,N_3486,N_3677);
and U4111 (N_4111,N_3706,N_3213);
nor U4112 (N_4112,N_3130,N_3921);
and U4113 (N_4113,N_3771,N_3104);
and U4114 (N_4114,N_3631,N_3229);
or U4115 (N_4115,N_3752,N_3412);
and U4116 (N_4116,N_3145,N_3098);
nand U4117 (N_4117,N_3558,N_3709);
nor U4118 (N_4118,N_3996,N_3069);
nand U4119 (N_4119,N_3688,N_3742);
xnor U4120 (N_4120,N_3887,N_3090);
and U4121 (N_4121,N_3930,N_3809);
xor U4122 (N_4122,N_3908,N_3535);
nand U4123 (N_4123,N_3122,N_3565);
or U4124 (N_4124,N_3739,N_3345);
or U4125 (N_4125,N_3593,N_3913);
nand U4126 (N_4126,N_3397,N_3826);
nor U4127 (N_4127,N_3133,N_3716);
and U4128 (N_4128,N_3851,N_3943);
nand U4129 (N_4129,N_3226,N_3804);
nor U4130 (N_4130,N_3137,N_3832);
nor U4131 (N_4131,N_3569,N_3311);
or U4132 (N_4132,N_3762,N_3953);
or U4133 (N_4133,N_3835,N_3556);
nand U4134 (N_4134,N_3016,N_3318);
or U4135 (N_4135,N_3453,N_3246);
nand U4136 (N_4136,N_3994,N_3534);
and U4137 (N_4137,N_3553,N_3479);
nor U4138 (N_4138,N_3508,N_3954);
or U4139 (N_4139,N_3021,N_3109);
nor U4140 (N_4140,N_3203,N_3541);
or U4141 (N_4141,N_3687,N_3017);
nor U4142 (N_4142,N_3545,N_3062);
or U4143 (N_4143,N_3050,N_3193);
and U4144 (N_4144,N_3582,N_3915);
nand U4145 (N_4145,N_3108,N_3333);
nor U4146 (N_4146,N_3585,N_3496);
and U4147 (N_4147,N_3140,N_3183);
or U4148 (N_4148,N_3362,N_3394);
or U4149 (N_4149,N_3723,N_3781);
xor U4150 (N_4150,N_3303,N_3425);
and U4151 (N_4151,N_3737,N_3157);
nor U4152 (N_4152,N_3652,N_3644);
and U4153 (N_4153,N_3040,N_3651);
nor U4154 (N_4154,N_3075,N_3861);
or U4155 (N_4155,N_3643,N_3295);
or U4156 (N_4156,N_3748,N_3348);
or U4157 (N_4157,N_3792,N_3009);
or U4158 (N_4158,N_3224,N_3926);
nand U4159 (N_4159,N_3165,N_3875);
nor U4160 (N_4160,N_3845,N_3049);
and U4161 (N_4161,N_3290,N_3163);
nor U4162 (N_4162,N_3025,N_3057);
or U4163 (N_4163,N_3985,N_3597);
or U4164 (N_4164,N_3828,N_3576);
nand U4165 (N_4165,N_3761,N_3800);
nor U4166 (N_4166,N_3659,N_3933);
and U4167 (N_4167,N_3275,N_3694);
nand U4168 (N_4168,N_3082,N_3139);
nand U4169 (N_4169,N_3253,N_3839);
and U4170 (N_4170,N_3579,N_3705);
or U4171 (N_4171,N_3936,N_3244);
nand U4172 (N_4172,N_3147,N_3507);
nor U4173 (N_4173,N_3815,N_3844);
or U4174 (N_4174,N_3031,N_3293);
or U4175 (N_4175,N_3186,N_3382);
nor U4176 (N_4176,N_3055,N_3354);
and U4177 (N_4177,N_3404,N_3578);
nand U4178 (N_4178,N_3307,N_3906);
nand U4179 (N_4179,N_3786,N_3796);
nor U4180 (N_4180,N_3973,N_3957);
nor U4181 (N_4181,N_3935,N_3401);
nand U4182 (N_4182,N_3243,N_3741);
nor U4183 (N_4183,N_3812,N_3465);
or U4184 (N_4184,N_3045,N_3271);
nor U4185 (N_4185,N_3724,N_3334);
and U4186 (N_4186,N_3918,N_3880);
or U4187 (N_4187,N_3471,N_3395);
or U4188 (N_4188,N_3441,N_3443);
and U4189 (N_4189,N_3036,N_3073);
or U4190 (N_4190,N_3777,N_3003);
and U4191 (N_4191,N_3500,N_3596);
or U4192 (N_4192,N_3738,N_3693);
or U4193 (N_4193,N_3299,N_3468);
or U4194 (N_4194,N_3667,N_3788);
and U4195 (N_4195,N_3824,N_3821);
nand U4196 (N_4196,N_3813,N_3410);
and U4197 (N_4197,N_3783,N_3525);
and U4198 (N_4198,N_3302,N_3042);
nor U4199 (N_4199,N_3174,N_3550);
nand U4200 (N_4200,N_3658,N_3202);
nand U4201 (N_4201,N_3494,N_3531);
and U4202 (N_4202,N_3629,N_3141);
nor U4203 (N_4203,N_3469,N_3171);
nor U4204 (N_4204,N_3053,N_3176);
xor U4205 (N_4205,N_3126,N_3969);
and U4206 (N_4206,N_3728,N_3983);
nor U4207 (N_4207,N_3888,N_3005);
nor U4208 (N_4208,N_3775,N_3230);
and U4209 (N_4209,N_3708,N_3250);
or U4210 (N_4210,N_3515,N_3416);
nand U4211 (N_4211,N_3313,N_3001);
nand U4212 (N_4212,N_3511,N_3127);
and U4213 (N_4213,N_3046,N_3350);
nor U4214 (N_4214,N_3320,N_3654);
nand U4215 (N_4215,N_3684,N_3864);
and U4216 (N_4216,N_3847,N_3527);
nand U4217 (N_4217,N_3902,N_3371);
and U4218 (N_4218,N_3240,N_3160);
or U4219 (N_4219,N_3301,N_3219);
nor U4220 (N_4220,N_3188,N_3893);
nand U4221 (N_4221,N_3172,N_3306);
nor U4222 (N_4222,N_3095,N_3867);
or U4223 (N_4223,N_3732,N_3825);
and U4224 (N_4224,N_3966,N_3549);
nand U4225 (N_4225,N_3884,N_3252);
and U4226 (N_4226,N_3435,N_3890);
or U4227 (N_4227,N_3497,N_3011);
nor U4228 (N_4228,N_3877,N_3255);
xor U4229 (N_4229,N_3418,N_3891);
or U4230 (N_4230,N_3795,N_3144);
and U4231 (N_4231,N_3114,N_3066);
or U4232 (N_4232,N_3873,N_3863);
or U4233 (N_4233,N_3759,N_3020);
or U4234 (N_4234,N_3937,N_3078);
and U4235 (N_4235,N_3030,N_3895);
and U4236 (N_4236,N_3989,N_3222);
nor U4237 (N_4237,N_3671,N_3013);
nand U4238 (N_4238,N_3780,N_3440);
or U4239 (N_4239,N_3624,N_3607);
nor U4240 (N_4240,N_3820,N_3142);
and U4241 (N_4241,N_3967,N_3561);
and U4242 (N_4242,N_3032,N_3974);
xor U4243 (N_4243,N_3087,N_3008);
nand U4244 (N_4244,N_3464,N_3241);
and U4245 (N_4245,N_3642,N_3697);
or U4246 (N_4246,N_3872,N_3437);
nor U4247 (N_4247,N_3882,N_3852);
nor U4248 (N_4248,N_3074,N_3970);
nor U4249 (N_4249,N_3562,N_3268);
or U4250 (N_4250,N_3522,N_3564);
and U4251 (N_4251,N_3196,N_3630);
nor U4252 (N_4252,N_3201,N_3731);
nor U4253 (N_4253,N_3619,N_3868);
and U4254 (N_4254,N_3858,N_3675);
nand U4255 (N_4255,N_3580,N_3287);
and U4256 (N_4256,N_3757,N_3627);
nand U4257 (N_4257,N_3997,N_3472);
nor U4258 (N_4258,N_3878,N_3770);
or U4259 (N_4259,N_3801,N_3584);
nor U4260 (N_4260,N_3051,N_3842);
nor U4261 (N_4261,N_3028,N_3259);
or U4262 (N_4262,N_3955,N_3586);
nand U4263 (N_4263,N_3692,N_3502);
nand U4264 (N_4264,N_3450,N_3662);
and U4265 (N_4265,N_3146,N_3310);
or U4266 (N_4266,N_3451,N_3729);
and U4267 (N_4267,N_3209,N_3023);
or U4268 (N_4268,N_3263,N_3571);
nand U4269 (N_4269,N_3071,N_3434);
nor U4270 (N_4270,N_3438,N_3976);
nor U4271 (N_4271,N_3588,N_3978);
nor U4272 (N_4272,N_3261,N_3600);
nand U4273 (N_4273,N_3717,N_3383);
nor U4274 (N_4274,N_3060,N_3105);
nor U4275 (N_4275,N_3192,N_3735);
nand U4276 (N_4276,N_3862,N_3914);
nor U4277 (N_4277,N_3322,N_3653);
nor U4278 (N_4278,N_3361,N_3101);
or U4279 (N_4279,N_3294,N_3808);
or U4280 (N_4280,N_3603,N_3223);
nand U4281 (N_4281,N_3743,N_3827);
nand U4282 (N_4282,N_3308,N_3187);
nor U4283 (N_4283,N_3484,N_3784);
nor U4284 (N_4284,N_3922,N_3681);
nor U4285 (N_4285,N_3180,N_3611);
nor U4286 (N_4286,N_3198,N_3014);
nand U4287 (N_4287,N_3691,N_3529);
and U4288 (N_4288,N_3524,N_3152);
nand U4289 (N_4289,N_3238,N_3356);
or U4290 (N_4290,N_3094,N_3422);
or U4291 (N_4291,N_3991,N_3092);
and U4292 (N_4292,N_3745,N_3834);
nor U4293 (N_4293,N_3963,N_3602);
or U4294 (N_4294,N_3072,N_3353);
nor U4295 (N_4295,N_3129,N_3758);
or U4296 (N_4296,N_3947,N_3945);
nand U4297 (N_4297,N_3722,N_3458);
nor U4298 (N_4298,N_3587,N_3316);
xnor U4299 (N_4299,N_3358,N_3512);
nor U4300 (N_4300,N_3977,N_3205);
nor U4301 (N_4301,N_3399,N_3924);
nor U4302 (N_4302,N_3760,N_3614);
or U4303 (N_4303,N_3993,N_3950);
or U4304 (N_4304,N_3782,N_3747);
nor U4305 (N_4305,N_3941,N_3857);
or U4306 (N_4306,N_3015,N_3843);
nand U4307 (N_4307,N_3551,N_3190);
or U4308 (N_4308,N_3481,N_3538);
or U4309 (N_4309,N_3236,N_3695);
and U4310 (N_4310,N_3920,N_3199);
nand U4311 (N_4311,N_3944,N_3177);
or U4312 (N_4312,N_3679,N_3124);
and U4313 (N_4313,N_3442,N_3298);
nor U4314 (N_4314,N_3474,N_3315);
or U4315 (N_4315,N_3058,N_3972);
and U4316 (N_4316,N_3523,N_3946);
nor U4317 (N_4317,N_3338,N_3672);
or U4318 (N_4318,N_3115,N_3823);
nand U4319 (N_4319,N_3665,N_3463);
nor U4320 (N_4320,N_3981,N_3668);
nand U4321 (N_4321,N_3473,N_3367);
nor U4322 (N_4322,N_3646,N_3276);
or U4323 (N_4323,N_3184,N_3208);
or U4324 (N_4324,N_3411,N_3297);
nor U4325 (N_4325,N_3216,N_3258);
and U4326 (N_4326,N_3111,N_3988);
and U4327 (N_4327,N_3871,N_3559);
or U4328 (N_4328,N_3620,N_3084);
xnor U4329 (N_4329,N_3138,N_3713);
and U4330 (N_4330,N_3164,N_3838);
nor U4331 (N_4331,N_3347,N_3197);
nor U4332 (N_4332,N_3547,N_3083);
and U4333 (N_4333,N_3103,N_3321);
nor U4334 (N_4334,N_3370,N_3686);
nor U4335 (N_4335,N_3131,N_3460);
nand U4336 (N_4336,N_3546,N_3896);
nand U4337 (N_4337,N_3033,N_3744);
nand U4338 (N_4338,N_3797,N_3448);
nand U4339 (N_4339,N_3363,N_3331);
nand U4340 (N_4340,N_3242,N_3625);
nand U4341 (N_4341,N_3634,N_3793);
or U4342 (N_4342,N_3381,N_3803);
or U4343 (N_4343,N_3022,N_3159);
or U4344 (N_4344,N_3749,N_3640);
nand U4345 (N_4345,N_3919,N_3120);
nand U4346 (N_4346,N_3552,N_3156);
or U4347 (N_4347,N_3097,N_3445);
nor U4348 (N_4348,N_3489,N_3339);
and U4349 (N_4349,N_3704,N_3670);
nor U4350 (N_4350,N_3249,N_3289);
or U4351 (N_4351,N_3475,N_3251);
or U4352 (N_4352,N_3344,N_3589);
xor U4353 (N_4353,N_3822,N_3830);
or U4354 (N_4354,N_3849,N_3696);
nand U4355 (N_4355,N_3396,N_3067);
nand U4356 (N_4356,N_3932,N_3819);
and U4357 (N_4357,N_3727,N_3305);
and U4358 (N_4358,N_3390,N_3376);
or U4359 (N_4359,N_3291,N_3254);
or U4360 (N_4360,N_3454,N_3116);
nand U4361 (N_4361,N_3807,N_3185);
or U4362 (N_4362,N_3234,N_3000);
or U4363 (N_4363,N_3424,N_3768);
nand U4364 (N_4364,N_3158,N_3773);
nor U4365 (N_4365,N_3319,N_3791);
or U4366 (N_4366,N_3591,N_3004);
nor U4367 (N_4367,N_3850,N_3034);
nand U4368 (N_4368,N_3664,N_3035);
nor U4369 (N_4369,N_3168,N_3514);
nor U4370 (N_4370,N_3278,N_3772);
nand U4371 (N_4371,N_3470,N_3150);
and U4372 (N_4372,N_3368,N_3372);
nand U4373 (N_4373,N_3790,N_3225);
and U4374 (N_4374,N_3149,N_3248);
or U4375 (N_4375,N_3879,N_3568);
nor U4376 (N_4376,N_3929,N_3154);
nor U4377 (N_4377,N_3495,N_3480);
and U4378 (N_4378,N_3903,N_3175);
and U4379 (N_4379,N_3702,N_3628);
and U4380 (N_4380,N_3900,N_3027);
or U4381 (N_4381,N_3491,N_3044);
nor U4382 (N_4382,N_3648,N_3638);
and U4383 (N_4383,N_3539,N_3641);
nand U4384 (N_4384,N_3649,N_3136);
nand U4385 (N_4385,N_3384,N_3961);
and U4386 (N_4386,N_3373,N_3938);
and U4387 (N_4387,N_3769,N_3056);
nand U4388 (N_4388,N_3329,N_3615);
nor U4389 (N_4389,N_3274,N_3632);
nand U4390 (N_4390,N_3387,N_3874);
nand U4391 (N_4391,N_3420,N_3779);
and U4392 (N_4392,N_3054,N_3365);
or U4393 (N_4393,N_3995,N_3391);
nand U4394 (N_4394,N_3840,N_3385);
and U4395 (N_4395,N_3841,N_3324);
and U4396 (N_4396,N_3816,N_3419);
nand U4397 (N_4397,N_3195,N_3220);
nand U4398 (N_4398,N_3799,N_3869);
nand U4399 (N_4399,N_3400,N_3118);
nor U4400 (N_4400,N_3848,N_3462);
nor U4401 (N_4401,N_3018,N_3916);
or U4402 (N_4402,N_3085,N_3836);
nor U4403 (N_4403,N_3829,N_3459);
nand U4404 (N_4404,N_3079,N_3178);
nor U4405 (N_4405,N_3548,N_3330);
nand U4406 (N_4406,N_3100,N_3106);
nor U4407 (N_4407,N_3504,N_3277);
nor U4408 (N_4408,N_3498,N_3751);
nor U4409 (N_4409,N_3364,N_3712);
or U4410 (N_4410,N_3960,N_3685);
and U4411 (N_4411,N_3673,N_3633);
nor U4412 (N_4412,N_3113,N_3403);
or U4413 (N_4413,N_3669,N_3233);
nor U4414 (N_4414,N_3528,N_3260);
nor U4415 (N_4415,N_3637,N_3698);
or U4416 (N_4416,N_3501,N_3774);
or U4417 (N_4417,N_3999,N_3928);
and U4418 (N_4418,N_3894,N_3262);
nor U4419 (N_4419,N_3678,N_3119);
nor U4420 (N_4420,N_3725,N_3029);
nand U4421 (N_4421,N_3026,N_3125);
or U4422 (N_4422,N_3608,N_3270);
or U4423 (N_4423,N_3855,N_3917);
and U4424 (N_4424,N_3467,N_3572);
nand U4425 (N_4425,N_3854,N_3212);
or U4426 (N_4426,N_3211,N_3217);
and U4427 (N_4427,N_3377,N_3355);
nor U4428 (N_4428,N_3881,N_3909);
or U4429 (N_4429,N_3161,N_3789);
nand U4430 (N_4430,N_3560,N_3292);
nor U4431 (N_4431,N_3590,N_3408);
or U4432 (N_4432,N_3616,N_3794);
or U4433 (N_4433,N_3112,N_3833);
nor U4434 (N_4434,N_3594,N_3540);
and U4435 (N_4435,N_3349,N_3817);
nor U4436 (N_4436,N_3189,N_3123);
nand U4437 (N_4437,N_3575,N_3934);
nand U4438 (N_4438,N_3070,N_3805);
nor U4439 (N_4439,N_3636,N_3661);
and U4440 (N_4440,N_3326,N_3785);
and U4441 (N_4441,N_3519,N_3998);
nand U4442 (N_4442,N_3392,N_3949);
or U4443 (N_4443,N_3787,N_3750);
nand U4444 (N_4444,N_3091,N_3767);
nor U4445 (N_4445,N_3019,N_3865);
nand U4446 (N_4446,N_3986,N_3730);
nor U4447 (N_4447,N_3904,N_3337);
or U4448 (N_4448,N_3284,N_3088);
nor U4449 (N_4449,N_3956,N_3570);
nand U4450 (N_4450,N_3052,N_3622);
and U4451 (N_4451,N_3581,N_3336);
nor U4452 (N_4452,N_3948,N_3645);
or U4453 (N_4453,N_3206,N_3405);
nor U4454 (N_4454,N_3925,N_3609);
nor U4455 (N_4455,N_3689,N_3231);
and U4456 (N_4456,N_3543,N_3719);
and U4457 (N_4457,N_3173,N_3086);
or U4458 (N_4458,N_3711,N_3352);
or U4459 (N_4459,N_3964,N_3754);
and U4460 (N_4460,N_3573,N_3041);
and U4461 (N_4461,N_3327,N_3554);
nor U4462 (N_4462,N_3037,N_3431);
nor U4463 (N_4463,N_3132,N_3980);
nand U4464 (N_4464,N_3912,N_3533);
and U4465 (N_4465,N_3505,N_3064);
nand U4466 (N_4466,N_3606,N_3487);
nand U4467 (N_4467,N_3557,N_3883);
nand U4468 (N_4468,N_3237,N_3059);
or U4469 (N_4469,N_3566,N_3660);
nand U4470 (N_4470,N_3421,N_3266);
nand U4471 (N_4471,N_3866,N_3107);
or U4472 (N_4472,N_3740,N_3746);
nand U4473 (N_4473,N_3360,N_3148);
or U4474 (N_4474,N_3207,N_3639);
or U4475 (N_4475,N_3218,N_3532);
nor U4476 (N_4476,N_3583,N_3117);
nor U4477 (N_4477,N_3407,N_3798);
or U4478 (N_4478,N_3409,N_3492);
nor U4479 (N_4479,N_3388,N_3984);
or U4480 (N_4480,N_3151,N_3245);
or U4481 (N_4481,N_3710,N_3296);
and U4482 (N_4482,N_3317,N_3210);
and U4483 (N_4483,N_3267,N_3756);
or U4484 (N_4484,N_3102,N_3846);
and U4485 (N_4485,N_3093,N_3433);
nor U4486 (N_4486,N_3386,N_3002);
nand U4487 (N_4487,N_3343,N_3181);
nand U4488 (N_4488,N_3380,N_3810);
and U4489 (N_4489,N_3604,N_3272);
nand U4490 (N_4490,N_3455,N_3378);
nor U4491 (N_4491,N_3910,N_3650);
nand U4492 (N_4492,N_3766,N_3663);
nand U4493 (N_4493,N_3765,N_3182);
nand U4494 (N_4494,N_3068,N_3542);
or U4495 (N_4495,N_3323,N_3886);
nand U4496 (N_4496,N_3911,N_3012);
or U4497 (N_4497,N_3595,N_3061);
nor U4498 (N_4498,N_3755,N_3965);
or U4499 (N_4499,N_3369,N_3080);
or U4500 (N_4500,N_3313,N_3422);
and U4501 (N_4501,N_3740,N_3818);
and U4502 (N_4502,N_3241,N_3647);
nor U4503 (N_4503,N_3921,N_3759);
nand U4504 (N_4504,N_3133,N_3967);
nor U4505 (N_4505,N_3147,N_3688);
or U4506 (N_4506,N_3965,N_3826);
nand U4507 (N_4507,N_3583,N_3749);
nor U4508 (N_4508,N_3789,N_3481);
nor U4509 (N_4509,N_3722,N_3120);
nand U4510 (N_4510,N_3537,N_3096);
or U4511 (N_4511,N_3673,N_3398);
and U4512 (N_4512,N_3134,N_3335);
or U4513 (N_4513,N_3698,N_3483);
or U4514 (N_4514,N_3643,N_3812);
nor U4515 (N_4515,N_3711,N_3443);
nor U4516 (N_4516,N_3148,N_3189);
or U4517 (N_4517,N_3438,N_3882);
nor U4518 (N_4518,N_3170,N_3699);
nor U4519 (N_4519,N_3718,N_3717);
nor U4520 (N_4520,N_3434,N_3519);
and U4521 (N_4521,N_3798,N_3680);
and U4522 (N_4522,N_3196,N_3444);
nand U4523 (N_4523,N_3417,N_3030);
and U4524 (N_4524,N_3186,N_3384);
and U4525 (N_4525,N_3934,N_3843);
nor U4526 (N_4526,N_3769,N_3286);
nor U4527 (N_4527,N_3245,N_3907);
nand U4528 (N_4528,N_3370,N_3817);
and U4529 (N_4529,N_3917,N_3621);
nor U4530 (N_4530,N_3283,N_3815);
or U4531 (N_4531,N_3427,N_3781);
or U4532 (N_4532,N_3837,N_3808);
and U4533 (N_4533,N_3245,N_3408);
and U4534 (N_4534,N_3646,N_3385);
nand U4535 (N_4535,N_3966,N_3928);
nor U4536 (N_4536,N_3055,N_3237);
or U4537 (N_4537,N_3111,N_3419);
nor U4538 (N_4538,N_3214,N_3982);
xnor U4539 (N_4539,N_3657,N_3095);
and U4540 (N_4540,N_3202,N_3085);
xnor U4541 (N_4541,N_3583,N_3290);
and U4542 (N_4542,N_3866,N_3236);
or U4543 (N_4543,N_3839,N_3127);
nor U4544 (N_4544,N_3145,N_3281);
and U4545 (N_4545,N_3274,N_3044);
nand U4546 (N_4546,N_3241,N_3339);
and U4547 (N_4547,N_3400,N_3286);
and U4548 (N_4548,N_3629,N_3846);
nand U4549 (N_4549,N_3167,N_3405);
nor U4550 (N_4550,N_3136,N_3615);
nand U4551 (N_4551,N_3853,N_3345);
nor U4552 (N_4552,N_3021,N_3096);
nand U4553 (N_4553,N_3033,N_3463);
or U4554 (N_4554,N_3830,N_3389);
nor U4555 (N_4555,N_3932,N_3454);
nand U4556 (N_4556,N_3533,N_3113);
or U4557 (N_4557,N_3446,N_3390);
or U4558 (N_4558,N_3521,N_3311);
or U4559 (N_4559,N_3299,N_3591);
nor U4560 (N_4560,N_3810,N_3005);
or U4561 (N_4561,N_3990,N_3785);
nand U4562 (N_4562,N_3894,N_3308);
or U4563 (N_4563,N_3883,N_3947);
nand U4564 (N_4564,N_3943,N_3155);
nand U4565 (N_4565,N_3677,N_3334);
nand U4566 (N_4566,N_3210,N_3892);
nand U4567 (N_4567,N_3215,N_3935);
nand U4568 (N_4568,N_3497,N_3121);
nand U4569 (N_4569,N_3615,N_3100);
and U4570 (N_4570,N_3004,N_3344);
nor U4571 (N_4571,N_3950,N_3315);
nor U4572 (N_4572,N_3530,N_3121);
xnor U4573 (N_4573,N_3666,N_3577);
or U4574 (N_4574,N_3771,N_3277);
nand U4575 (N_4575,N_3964,N_3844);
nor U4576 (N_4576,N_3315,N_3488);
nor U4577 (N_4577,N_3362,N_3087);
nor U4578 (N_4578,N_3796,N_3221);
or U4579 (N_4579,N_3461,N_3146);
nand U4580 (N_4580,N_3597,N_3528);
nand U4581 (N_4581,N_3788,N_3025);
or U4582 (N_4582,N_3590,N_3009);
nand U4583 (N_4583,N_3956,N_3698);
nand U4584 (N_4584,N_3871,N_3827);
nand U4585 (N_4585,N_3328,N_3326);
and U4586 (N_4586,N_3573,N_3578);
nor U4587 (N_4587,N_3300,N_3839);
nor U4588 (N_4588,N_3634,N_3737);
or U4589 (N_4589,N_3858,N_3911);
nor U4590 (N_4590,N_3172,N_3565);
nor U4591 (N_4591,N_3380,N_3066);
nand U4592 (N_4592,N_3142,N_3548);
nor U4593 (N_4593,N_3686,N_3325);
nor U4594 (N_4594,N_3043,N_3958);
nand U4595 (N_4595,N_3271,N_3264);
or U4596 (N_4596,N_3145,N_3336);
and U4597 (N_4597,N_3974,N_3838);
nand U4598 (N_4598,N_3359,N_3973);
nand U4599 (N_4599,N_3627,N_3012);
and U4600 (N_4600,N_3062,N_3377);
nand U4601 (N_4601,N_3421,N_3050);
nor U4602 (N_4602,N_3929,N_3771);
and U4603 (N_4603,N_3707,N_3229);
and U4604 (N_4604,N_3039,N_3035);
nor U4605 (N_4605,N_3195,N_3576);
xor U4606 (N_4606,N_3452,N_3658);
nand U4607 (N_4607,N_3384,N_3795);
and U4608 (N_4608,N_3105,N_3204);
or U4609 (N_4609,N_3128,N_3935);
or U4610 (N_4610,N_3633,N_3049);
or U4611 (N_4611,N_3526,N_3107);
and U4612 (N_4612,N_3124,N_3224);
nand U4613 (N_4613,N_3740,N_3947);
nand U4614 (N_4614,N_3613,N_3585);
nor U4615 (N_4615,N_3905,N_3993);
and U4616 (N_4616,N_3281,N_3950);
and U4617 (N_4617,N_3272,N_3730);
or U4618 (N_4618,N_3217,N_3226);
and U4619 (N_4619,N_3398,N_3778);
nand U4620 (N_4620,N_3297,N_3967);
and U4621 (N_4621,N_3290,N_3384);
and U4622 (N_4622,N_3313,N_3692);
or U4623 (N_4623,N_3933,N_3543);
nand U4624 (N_4624,N_3268,N_3342);
nor U4625 (N_4625,N_3262,N_3727);
nand U4626 (N_4626,N_3139,N_3309);
or U4627 (N_4627,N_3986,N_3135);
nand U4628 (N_4628,N_3336,N_3415);
and U4629 (N_4629,N_3356,N_3760);
nor U4630 (N_4630,N_3944,N_3851);
and U4631 (N_4631,N_3846,N_3071);
nand U4632 (N_4632,N_3853,N_3966);
or U4633 (N_4633,N_3260,N_3317);
and U4634 (N_4634,N_3148,N_3854);
nor U4635 (N_4635,N_3410,N_3843);
nand U4636 (N_4636,N_3091,N_3756);
and U4637 (N_4637,N_3067,N_3746);
nand U4638 (N_4638,N_3648,N_3472);
nand U4639 (N_4639,N_3778,N_3843);
nor U4640 (N_4640,N_3306,N_3844);
xor U4641 (N_4641,N_3864,N_3328);
nor U4642 (N_4642,N_3528,N_3844);
nor U4643 (N_4643,N_3939,N_3807);
and U4644 (N_4644,N_3833,N_3066);
and U4645 (N_4645,N_3496,N_3178);
or U4646 (N_4646,N_3444,N_3764);
nor U4647 (N_4647,N_3226,N_3908);
or U4648 (N_4648,N_3422,N_3142);
or U4649 (N_4649,N_3663,N_3939);
nand U4650 (N_4650,N_3188,N_3684);
or U4651 (N_4651,N_3666,N_3429);
nor U4652 (N_4652,N_3528,N_3590);
and U4653 (N_4653,N_3757,N_3318);
nand U4654 (N_4654,N_3338,N_3968);
nor U4655 (N_4655,N_3599,N_3272);
nor U4656 (N_4656,N_3909,N_3574);
and U4657 (N_4657,N_3653,N_3461);
and U4658 (N_4658,N_3087,N_3218);
nand U4659 (N_4659,N_3464,N_3510);
nand U4660 (N_4660,N_3505,N_3625);
and U4661 (N_4661,N_3367,N_3415);
or U4662 (N_4662,N_3739,N_3521);
and U4663 (N_4663,N_3403,N_3880);
and U4664 (N_4664,N_3776,N_3474);
nor U4665 (N_4665,N_3830,N_3670);
and U4666 (N_4666,N_3421,N_3871);
or U4667 (N_4667,N_3944,N_3382);
nand U4668 (N_4668,N_3183,N_3814);
or U4669 (N_4669,N_3524,N_3824);
and U4670 (N_4670,N_3254,N_3385);
and U4671 (N_4671,N_3018,N_3275);
or U4672 (N_4672,N_3255,N_3637);
xnor U4673 (N_4673,N_3309,N_3057);
nor U4674 (N_4674,N_3354,N_3700);
nand U4675 (N_4675,N_3848,N_3282);
nand U4676 (N_4676,N_3134,N_3653);
nand U4677 (N_4677,N_3477,N_3963);
and U4678 (N_4678,N_3154,N_3104);
nor U4679 (N_4679,N_3200,N_3493);
nor U4680 (N_4680,N_3827,N_3255);
nor U4681 (N_4681,N_3186,N_3334);
nand U4682 (N_4682,N_3678,N_3652);
and U4683 (N_4683,N_3936,N_3793);
or U4684 (N_4684,N_3479,N_3053);
nand U4685 (N_4685,N_3307,N_3493);
nor U4686 (N_4686,N_3628,N_3366);
nor U4687 (N_4687,N_3790,N_3059);
nor U4688 (N_4688,N_3246,N_3276);
and U4689 (N_4689,N_3780,N_3993);
and U4690 (N_4690,N_3103,N_3457);
nand U4691 (N_4691,N_3783,N_3741);
and U4692 (N_4692,N_3627,N_3842);
nor U4693 (N_4693,N_3112,N_3749);
and U4694 (N_4694,N_3694,N_3440);
and U4695 (N_4695,N_3805,N_3829);
nand U4696 (N_4696,N_3097,N_3323);
nand U4697 (N_4697,N_3897,N_3350);
nor U4698 (N_4698,N_3613,N_3574);
or U4699 (N_4699,N_3178,N_3643);
or U4700 (N_4700,N_3160,N_3813);
nand U4701 (N_4701,N_3251,N_3845);
xnor U4702 (N_4702,N_3736,N_3684);
nor U4703 (N_4703,N_3834,N_3450);
and U4704 (N_4704,N_3253,N_3805);
nor U4705 (N_4705,N_3334,N_3630);
or U4706 (N_4706,N_3320,N_3002);
nand U4707 (N_4707,N_3019,N_3597);
or U4708 (N_4708,N_3761,N_3773);
or U4709 (N_4709,N_3780,N_3039);
nor U4710 (N_4710,N_3723,N_3121);
and U4711 (N_4711,N_3846,N_3178);
nand U4712 (N_4712,N_3889,N_3444);
or U4713 (N_4713,N_3614,N_3156);
or U4714 (N_4714,N_3747,N_3841);
nand U4715 (N_4715,N_3783,N_3638);
or U4716 (N_4716,N_3485,N_3408);
or U4717 (N_4717,N_3147,N_3176);
nand U4718 (N_4718,N_3419,N_3402);
and U4719 (N_4719,N_3656,N_3861);
nor U4720 (N_4720,N_3512,N_3965);
nand U4721 (N_4721,N_3977,N_3182);
nand U4722 (N_4722,N_3471,N_3826);
nand U4723 (N_4723,N_3807,N_3685);
and U4724 (N_4724,N_3684,N_3679);
or U4725 (N_4725,N_3958,N_3593);
nand U4726 (N_4726,N_3570,N_3924);
and U4727 (N_4727,N_3740,N_3082);
nand U4728 (N_4728,N_3508,N_3461);
nand U4729 (N_4729,N_3163,N_3701);
and U4730 (N_4730,N_3804,N_3999);
nor U4731 (N_4731,N_3065,N_3287);
or U4732 (N_4732,N_3058,N_3579);
or U4733 (N_4733,N_3586,N_3053);
or U4734 (N_4734,N_3184,N_3315);
nor U4735 (N_4735,N_3027,N_3743);
and U4736 (N_4736,N_3851,N_3272);
or U4737 (N_4737,N_3941,N_3711);
nor U4738 (N_4738,N_3170,N_3619);
nand U4739 (N_4739,N_3968,N_3706);
or U4740 (N_4740,N_3241,N_3856);
nand U4741 (N_4741,N_3360,N_3916);
or U4742 (N_4742,N_3582,N_3306);
or U4743 (N_4743,N_3309,N_3566);
and U4744 (N_4744,N_3487,N_3769);
nor U4745 (N_4745,N_3950,N_3971);
nand U4746 (N_4746,N_3951,N_3669);
nand U4747 (N_4747,N_3523,N_3983);
or U4748 (N_4748,N_3383,N_3099);
nor U4749 (N_4749,N_3190,N_3884);
nor U4750 (N_4750,N_3615,N_3819);
xor U4751 (N_4751,N_3353,N_3330);
or U4752 (N_4752,N_3702,N_3137);
and U4753 (N_4753,N_3118,N_3969);
or U4754 (N_4754,N_3830,N_3578);
nand U4755 (N_4755,N_3984,N_3126);
or U4756 (N_4756,N_3638,N_3434);
or U4757 (N_4757,N_3977,N_3836);
and U4758 (N_4758,N_3572,N_3823);
nor U4759 (N_4759,N_3911,N_3100);
nand U4760 (N_4760,N_3788,N_3716);
nor U4761 (N_4761,N_3216,N_3632);
nand U4762 (N_4762,N_3868,N_3212);
nor U4763 (N_4763,N_3428,N_3174);
and U4764 (N_4764,N_3021,N_3501);
nor U4765 (N_4765,N_3485,N_3444);
and U4766 (N_4766,N_3983,N_3941);
nand U4767 (N_4767,N_3983,N_3093);
or U4768 (N_4768,N_3529,N_3006);
nor U4769 (N_4769,N_3355,N_3120);
or U4770 (N_4770,N_3520,N_3300);
or U4771 (N_4771,N_3204,N_3613);
nand U4772 (N_4772,N_3738,N_3328);
nor U4773 (N_4773,N_3225,N_3835);
and U4774 (N_4774,N_3787,N_3697);
and U4775 (N_4775,N_3802,N_3198);
or U4776 (N_4776,N_3347,N_3784);
and U4777 (N_4777,N_3182,N_3749);
and U4778 (N_4778,N_3060,N_3155);
nor U4779 (N_4779,N_3536,N_3290);
and U4780 (N_4780,N_3097,N_3871);
nor U4781 (N_4781,N_3556,N_3758);
and U4782 (N_4782,N_3487,N_3829);
nor U4783 (N_4783,N_3701,N_3195);
or U4784 (N_4784,N_3121,N_3890);
or U4785 (N_4785,N_3808,N_3072);
nand U4786 (N_4786,N_3885,N_3073);
or U4787 (N_4787,N_3585,N_3436);
nand U4788 (N_4788,N_3450,N_3543);
and U4789 (N_4789,N_3380,N_3729);
or U4790 (N_4790,N_3782,N_3848);
and U4791 (N_4791,N_3231,N_3425);
nand U4792 (N_4792,N_3960,N_3814);
and U4793 (N_4793,N_3729,N_3819);
nor U4794 (N_4794,N_3947,N_3291);
or U4795 (N_4795,N_3820,N_3015);
nand U4796 (N_4796,N_3824,N_3816);
nand U4797 (N_4797,N_3500,N_3358);
nor U4798 (N_4798,N_3954,N_3495);
and U4799 (N_4799,N_3849,N_3340);
or U4800 (N_4800,N_3340,N_3258);
nand U4801 (N_4801,N_3933,N_3257);
or U4802 (N_4802,N_3196,N_3684);
nand U4803 (N_4803,N_3431,N_3022);
or U4804 (N_4804,N_3502,N_3101);
nor U4805 (N_4805,N_3118,N_3632);
and U4806 (N_4806,N_3727,N_3090);
or U4807 (N_4807,N_3954,N_3633);
nor U4808 (N_4808,N_3447,N_3312);
xor U4809 (N_4809,N_3598,N_3841);
nor U4810 (N_4810,N_3807,N_3942);
and U4811 (N_4811,N_3359,N_3210);
nand U4812 (N_4812,N_3551,N_3120);
nor U4813 (N_4813,N_3887,N_3376);
or U4814 (N_4814,N_3317,N_3681);
xor U4815 (N_4815,N_3990,N_3675);
or U4816 (N_4816,N_3740,N_3484);
and U4817 (N_4817,N_3718,N_3196);
or U4818 (N_4818,N_3268,N_3247);
and U4819 (N_4819,N_3911,N_3366);
nor U4820 (N_4820,N_3970,N_3716);
and U4821 (N_4821,N_3257,N_3747);
or U4822 (N_4822,N_3794,N_3182);
and U4823 (N_4823,N_3438,N_3835);
or U4824 (N_4824,N_3711,N_3669);
nor U4825 (N_4825,N_3969,N_3035);
and U4826 (N_4826,N_3965,N_3053);
nor U4827 (N_4827,N_3825,N_3787);
and U4828 (N_4828,N_3633,N_3004);
nand U4829 (N_4829,N_3603,N_3861);
xor U4830 (N_4830,N_3469,N_3359);
nor U4831 (N_4831,N_3586,N_3959);
and U4832 (N_4832,N_3582,N_3561);
nor U4833 (N_4833,N_3608,N_3470);
nor U4834 (N_4834,N_3651,N_3098);
nand U4835 (N_4835,N_3704,N_3536);
nand U4836 (N_4836,N_3892,N_3621);
nor U4837 (N_4837,N_3142,N_3245);
nor U4838 (N_4838,N_3546,N_3498);
nand U4839 (N_4839,N_3261,N_3192);
nand U4840 (N_4840,N_3689,N_3886);
and U4841 (N_4841,N_3506,N_3712);
nor U4842 (N_4842,N_3059,N_3883);
nor U4843 (N_4843,N_3512,N_3010);
nand U4844 (N_4844,N_3362,N_3003);
xnor U4845 (N_4845,N_3969,N_3984);
and U4846 (N_4846,N_3177,N_3404);
nor U4847 (N_4847,N_3514,N_3797);
nor U4848 (N_4848,N_3301,N_3343);
and U4849 (N_4849,N_3161,N_3930);
nand U4850 (N_4850,N_3030,N_3248);
and U4851 (N_4851,N_3379,N_3277);
or U4852 (N_4852,N_3949,N_3547);
and U4853 (N_4853,N_3035,N_3151);
nor U4854 (N_4854,N_3475,N_3347);
or U4855 (N_4855,N_3461,N_3411);
nand U4856 (N_4856,N_3738,N_3464);
and U4857 (N_4857,N_3351,N_3611);
or U4858 (N_4858,N_3270,N_3495);
nor U4859 (N_4859,N_3017,N_3237);
nand U4860 (N_4860,N_3733,N_3553);
nor U4861 (N_4861,N_3839,N_3864);
or U4862 (N_4862,N_3760,N_3209);
and U4863 (N_4863,N_3512,N_3259);
xor U4864 (N_4864,N_3019,N_3294);
nor U4865 (N_4865,N_3445,N_3053);
or U4866 (N_4866,N_3848,N_3523);
and U4867 (N_4867,N_3912,N_3416);
nand U4868 (N_4868,N_3390,N_3035);
nor U4869 (N_4869,N_3172,N_3011);
and U4870 (N_4870,N_3965,N_3819);
or U4871 (N_4871,N_3252,N_3044);
or U4872 (N_4872,N_3611,N_3589);
nor U4873 (N_4873,N_3687,N_3581);
nand U4874 (N_4874,N_3498,N_3384);
or U4875 (N_4875,N_3863,N_3704);
nor U4876 (N_4876,N_3953,N_3806);
nor U4877 (N_4877,N_3667,N_3506);
or U4878 (N_4878,N_3823,N_3320);
xor U4879 (N_4879,N_3854,N_3286);
nand U4880 (N_4880,N_3131,N_3037);
nor U4881 (N_4881,N_3750,N_3857);
nand U4882 (N_4882,N_3451,N_3189);
and U4883 (N_4883,N_3097,N_3591);
and U4884 (N_4884,N_3640,N_3068);
and U4885 (N_4885,N_3714,N_3173);
nor U4886 (N_4886,N_3898,N_3592);
nor U4887 (N_4887,N_3440,N_3176);
nand U4888 (N_4888,N_3247,N_3001);
nand U4889 (N_4889,N_3652,N_3508);
nand U4890 (N_4890,N_3995,N_3684);
nor U4891 (N_4891,N_3186,N_3896);
or U4892 (N_4892,N_3978,N_3315);
nor U4893 (N_4893,N_3411,N_3190);
nor U4894 (N_4894,N_3158,N_3405);
nand U4895 (N_4895,N_3329,N_3840);
nand U4896 (N_4896,N_3504,N_3970);
or U4897 (N_4897,N_3282,N_3070);
nand U4898 (N_4898,N_3953,N_3236);
nor U4899 (N_4899,N_3041,N_3293);
or U4900 (N_4900,N_3083,N_3495);
nor U4901 (N_4901,N_3301,N_3155);
and U4902 (N_4902,N_3567,N_3245);
or U4903 (N_4903,N_3102,N_3384);
or U4904 (N_4904,N_3548,N_3641);
nor U4905 (N_4905,N_3375,N_3426);
nor U4906 (N_4906,N_3769,N_3205);
or U4907 (N_4907,N_3564,N_3450);
nor U4908 (N_4908,N_3179,N_3315);
or U4909 (N_4909,N_3432,N_3572);
nand U4910 (N_4910,N_3246,N_3233);
nand U4911 (N_4911,N_3435,N_3320);
or U4912 (N_4912,N_3023,N_3494);
nand U4913 (N_4913,N_3291,N_3596);
and U4914 (N_4914,N_3978,N_3894);
xnor U4915 (N_4915,N_3027,N_3423);
and U4916 (N_4916,N_3658,N_3666);
and U4917 (N_4917,N_3563,N_3336);
nor U4918 (N_4918,N_3592,N_3963);
xnor U4919 (N_4919,N_3394,N_3088);
and U4920 (N_4920,N_3274,N_3351);
and U4921 (N_4921,N_3815,N_3911);
nand U4922 (N_4922,N_3603,N_3014);
nor U4923 (N_4923,N_3662,N_3726);
or U4924 (N_4924,N_3657,N_3218);
or U4925 (N_4925,N_3295,N_3624);
nor U4926 (N_4926,N_3964,N_3643);
nor U4927 (N_4927,N_3260,N_3712);
nor U4928 (N_4928,N_3057,N_3427);
nand U4929 (N_4929,N_3371,N_3501);
nand U4930 (N_4930,N_3284,N_3082);
nor U4931 (N_4931,N_3280,N_3396);
xor U4932 (N_4932,N_3014,N_3380);
xnor U4933 (N_4933,N_3940,N_3664);
and U4934 (N_4934,N_3761,N_3181);
or U4935 (N_4935,N_3102,N_3086);
nand U4936 (N_4936,N_3650,N_3821);
or U4937 (N_4937,N_3902,N_3805);
or U4938 (N_4938,N_3700,N_3154);
or U4939 (N_4939,N_3919,N_3627);
and U4940 (N_4940,N_3350,N_3290);
nor U4941 (N_4941,N_3576,N_3229);
nor U4942 (N_4942,N_3345,N_3002);
nor U4943 (N_4943,N_3013,N_3066);
or U4944 (N_4944,N_3747,N_3405);
or U4945 (N_4945,N_3515,N_3372);
and U4946 (N_4946,N_3352,N_3477);
nand U4947 (N_4947,N_3751,N_3625);
nand U4948 (N_4948,N_3992,N_3954);
or U4949 (N_4949,N_3777,N_3914);
nand U4950 (N_4950,N_3213,N_3036);
nand U4951 (N_4951,N_3635,N_3590);
and U4952 (N_4952,N_3402,N_3092);
and U4953 (N_4953,N_3838,N_3147);
and U4954 (N_4954,N_3395,N_3461);
or U4955 (N_4955,N_3262,N_3712);
nor U4956 (N_4956,N_3846,N_3247);
or U4957 (N_4957,N_3691,N_3624);
nand U4958 (N_4958,N_3071,N_3321);
and U4959 (N_4959,N_3116,N_3051);
nor U4960 (N_4960,N_3577,N_3532);
and U4961 (N_4961,N_3240,N_3962);
and U4962 (N_4962,N_3949,N_3722);
nor U4963 (N_4963,N_3267,N_3115);
and U4964 (N_4964,N_3972,N_3609);
nor U4965 (N_4965,N_3512,N_3394);
and U4966 (N_4966,N_3653,N_3167);
or U4967 (N_4967,N_3315,N_3136);
nand U4968 (N_4968,N_3657,N_3395);
and U4969 (N_4969,N_3252,N_3628);
or U4970 (N_4970,N_3087,N_3136);
or U4971 (N_4971,N_3811,N_3402);
or U4972 (N_4972,N_3810,N_3469);
nor U4973 (N_4973,N_3969,N_3663);
and U4974 (N_4974,N_3093,N_3617);
nand U4975 (N_4975,N_3468,N_3861);
or U4976 (N_4976,N_3480,N_3719);
nor U4977 (N_4977,N_3182,N_3118);
and U4978 (N_4978,N_3951,N_3110);
nand U4979 (N_4979,N_3803,N_3249);
or U4980 (N_4980,N_3179,N_3978);
nor U4981 (N_4981,N_3090,N_3384);
nor U4982 (N_4982,N_3375,N_3293);
or U4983 (N_4983,N_3519,N_3168);
and U4984 (N_4984,N_3802,N_3864);
and U4985 (N_4985,N_3510,N_3993);
or U4986 (N_4986,N_3354,N_3747);
or U4987 (N_4987,N_3525,N_3199);
or U4988 (N_4988,N_3019,N_3913);
and U4989 (N_4989,N_3014,N_3539);
and U4990 (N_4990,N_3888,N_3588);
or U4991 (N_4991,N_3173,N_3205);
nand U4992 (N_4992,N_3344,N_3643);
nand U4993 (N_4993,N_3016,N_3382);
nor U4994 (N_4994,N_3544,N_3990);
or U4995 (N_4995,N_3219,N_3222);
nand U4996 (N_4996,N_3362,N_3702);
and U4997 (N_4997,N_3140,N_3415);
and U4998 (N_4998,N_3510,N_3631);
nor U4999 (N_4999,N_3098,N_3707);
nand UO_0 (O_0,N_4590,N_4087);
and UO_1 (O_1,N_4318,N_4122);
nor UO_2 (O_2,N_4094,N_4718);
nor UO_3 (O_3,N_4507,N_4526);
nand UO_4 (O_4,N_4705,N_4444);
nand UO_5 (O_5,N_4785,N_4216);
nor UO_6 (O_6,N_4648,N_4263);
and UO_7 (O_7,N_4544,N_4312);
or UO_8 (O_8,N_4661,N_4083);
or UO_9 (O_9,N_4587,N_4824);
and UO_10 (O_10,N_4163,N_4267);
or UO_11 (O_11,N_4652,N_4669);
and UO_12 (O_12,N_4126,N_4425);
nor UO_13 (O_13,N_4496,N_4070);
nand UO_14 (O_14,N_4963,N_4048);
nor UO_15 (O_15,N_4497,N_4096);
nand UO_16 (O_16,N_4665,N_4819);
nor UO_17 (O_17,N_4671,N_4513);
or UO_18 (O_18,N_4381,N_4942);
or UO_19 (O_19,N_4626,N_4064);
nand UO_20 (O_20,N_4879,N_4723);
and UO_21 (O_21,N_4435,N_4757);
or UO_22 (O_22,N_4749,N_4128);
or UO_23 (O_23,N_4609,N_4328);
nor UO_24 (O_24,N_4232,N_4235);
nand UO_25 (O_25,N_4599,N_4870);
nor UO_26 (O_26,N_4647,N_4485);
nor UO_27 (O_27,N_4811,N_4564);
nor UO_28 (O_28,N_4180,N_4281);
nor UO_29 (O_29,N_4023,N_4234);
nor UO_30 (O_30,N_4270,N_4617);
or UO_31 (O_31,N_4585,N_4890);
or UO_32 (O_32,N_4997,N_4199);
nor UO_33 (O_33,N_4251,N_4744);
nand UO_34 (O_34,N_4539,N_4129);
and UO_35 (O_35,N_4324,N_4220);
nor UO_36 (O_36,N_4548,N_4771);
nor UO_37 (O_37,N_4923,N_4189);
nor UO_38 (O_38,N_4510,N_4957);
and UO_39 (O_39,N_4115,N_4020);
nand UO_40 (O_40,N_4568,N_4569);
nor UO_41 (O_41,N_4368,N_4708);
or UO_42 (O_42,N_4334,N_4344);
nand UO_43 (O_43,N_4442,N_4243);
or UO_44 (O_44,N_4441,N_4773);
or UO_45 (O_45,N_4546,N_4833);
nand UO_46 (O_46,N_4698,N_4340);
and UO_47 (O_47,N_4950,N_4909);
nand UO_48 (O_48,N_4006,N_4753);
nand UO_49 (O_49,N_4802,N_4371);
nor UO_50 (O_50,N_4296,N_4223);
and UO_51 (O_51,N_4641,N_4466);
nor UO_52 (O_52,N_4953,N_4619);
or UO_53 (O_53,N_4213,N_4822);
and UO_54 (O_54,N_4460,N_4552);
and UO_55 (O_55,N_4016,N_4628);
nand UO_56 (O_56,N_4856,N_4151);
nor UO_57 (O_57,N_4149,N_4433);
nand UO_58 (O_58,N_4256,N_4388);
or UO_59 (O_59,N_4706,N_4712);
nor UO_60 (O_60,N_4028,N_4204);
and UO_61 (O_61,N_4398,N_4376);
and UO_62 (O_62,N_4470,N_4039);
and UO_63 (O_63,N_4105,N_4673);
and UO_64 (O_64,N_4404,N_4634);
and UO_65 (O_65,N_4022,N_4306);
nor UO_66 (O_66,N_4101,N_4035);
nor UO_67 (O_67,N_4534,N_4735);
or UO_68 (O_68,N_4644,N_4616);
or UO_69 (O_69,N_4522,N_4409);
nand UO_70 (O_70,N_4517,N_4882);
nand UO_71 (O_71,N_4295,N_4717);
nor UO_72 (O_72,N_4104,N_4147);
and UO_73 (O_73,N_4554,N_4214);
or UO_74 (O_74,N_4203,N_4314);
xnor UO_75 (O_75,N_4872,N_4157);
nor UO_76 (O_76,N_4095,N_4166);
or UO_77 (O_77,N_4715,N_4403);
or UO_78 (O_78,N_4264,N_4218);
nor UO_79 (O_79,N_4037,N_4484);
nor UO_80 (O_80,N_4479,N_4412);
and UO_81 (O_81,N_4471,N_4797);
nand UO_82 (O_82,N_4816,N_4250);
or UO_83 (O_83,N_4138,N_4261);
nand UO_84 (O_84,N_4451,N_4922);
and UO_85 (O_85,N_4191,N_4003);
nand UO_86 (O_86,N_4254,N_4495);
nand UO_87 (O_87,N_4774,N_4065);
or UO_88 (O_88,N_4044,N_4960);
and UO_89 (O_89,N_4134,N_4415);
or UO_90 (O_90,N_4366,N_4174);
nand UO_91 (O_91,N_4472,N_4826);
or UO_92 (O_92,N_4042,N_4280);
and UO_93 (O_93,N_4084,N_4370);
or UO_94 (O_94,N_4931,N_4165);
nor UO_95 (O_95,N_4493,N_4756);
and UO_96 (O_96,N_4211,N_4766);
and UO_97 (O_97,N_4878,N_4730);
or UO_98 (O_98,N_4574,N_4528);
nor UO_99 (O_99,N_4969,N_4373);
nand UO_100 (O_100,N_4810,N_4563);
or UO_101 (O_101,N_4352,N_4248);
nor UO_102 (O_102,N_4697,N_4937);
nor UO_103 (O_103,N_4456,N_4760);
or UO_104 (O_104,N_4518,N_4386);
and UO_105 (O_105,N_4406,N_4947);
or UO_106 (O_106,N_4259,N_4168);
or UO_107 (O_107,N_4612,N_4202);
nor UO_108 (O_108,N_4500,N_4868);
nand UO_109 (O_109,N_4419,N_4242);
and UO_110 (O_110,N_4776,N_4193);
or UO_111 (O_111,N_4136,N_4855);
and UO_112 (O_112,N_4764,N_4655);
or UO_113 (O_113,N_4965,N_4973);
xnor UO_114 (O_114,N_4778,N_4289);
and UO_115 (O_115,N_4883,N_4450);
xor UO_116 (O_116,N_4643,N_4888);
and UO_117 (O_117,N_4558,N_4996);
nor UO_118 (O_118,N_4750,N_4173);
nor UO_119 (O_119,N_4029,N_4565);
nor UO_120 (O_120,N_4262,N_4567);
and UO_121 (O_121,N_4972,N_4967);
and UO_122 (O_122,N_4047,N_4310);
nor UO_123 (O_123,N_4278,N_4678);
nor UO_124 (O_124,N_4355,N_4977);
nor UO_125 (O_125,N_4089,N_4463);
xor UO_126 (O_126,N_4672,N_4536);
and UO_127 (O_127,N_4781,N_4311);
and UO_128 (O_128,N_4841,N_4422);
nand UO_129 (O_129,N_4072,N_4688);
nor UO_130 (O_130,N_4566,N_4508);
nand UO_131 (O_131,N_4139,N_4579);
and UO_132 (O_132,N_4102,N_4374);
nand UO_133 (O_133,N_4452,N_4176);
and UO_134 (O_134,N_4219,N_4863);
nor UO_135 (O_135,N_4867,N_4217);
and UO_136 (O_136,N_4358,N_4144);
nand UO_137 (O_137,N_4142,N_4835);
or UO_138 (O_138,N_4125,N_4813);
and UO_139 (O_139,N_4015,N_4086);
nor UO_140 (O_140,N_4754,N_4237);
nand UO_141 (O_141,N_4746,N_4146);
and UO_142 (O_142,N_4864,N_4762);
nand UO_143 (O_143,N_4545,N_4710);
nor UO_144 (O_144,N_4247,N_4091);
and UO_145 (O_145,N_4831,N_4081);
or UO_146 (O_146,N_4745,N_4114);
or UO_147 (O_147,N_4828,N_4761);
or UO_148 (O_148,N_4962,N_4130);
and UO_149 (O_149,N_4474,N_4755);
nand UO_150 (O_150,N_4881,N_4783);
nand UO_151 (O_151,N_4946,N_4309);
or UO_152 (O_152,N_4702,N_4951);
nor UO_153 (O_153,N_4359,N_4181);
and UO_154 (O_154,N_4523,N_4955);
or UO_155 (O_155,N_4971,N_4431);
nand UO_156 (O_156,N_4468,N_4054);
or UO_157 (O_157,N_4695,N_4600);
nor UO_158 (O_158,N_4687,N_4194);
nor UO_159 (O_159,N_4793,N_4696);
and UO_160 (O_160,N_4562,N_4332);
or UO_161 (O_161,N_4052,N_4758);
nor UO_162 (O_162,N_4529,N_4492);
nand UO_163 (O_163,N_4230,N_4759);
and UO_164 (O_164,N_4722,N_4935);
and UO_165 (O_165,N_4055,N_4159);
nand UO_166 (O_166,N_4618,N_4869);
or UO_167 (O_167,N_4423,N_4814);
or UO_168 (O_168,N_4555,N_4538);
nand UO_169 (O_169,N_4459,N_4741);
nor UO_170 (O_170,N_4524,N_4288);
nand UO_171 (O_171,N_4928,N_4823);
and UO_172 (O_172,N_4827,N_4681);
nand UO_173 (O_173,N_4691,N_4933);
and UO_174 (O_174,N_4862,N_4448);
nand UO_175 (O_175,N_4876,N_4998);
and UO_176 (O_176,N_4121,N_4337);
or UO_177 (O_177,N_4910,N_4905);
nor UO_178 (O_178,N_4417,N_4748);
and UO_179 (O_179,N_4784,N_4238);
or UO_180 (O_180,N_4786,N_4620);
nand UO_181 (O_181,N_4155,N_4763);
and UO_182 (O_182,N_4791,N_4990);
nand UO_183 (O_183,N_4919,N_4901);
and UO_184 (O_184,N_4063,N_4794);
nand UO_185 (O_185,N_4740,N_4920);
and UO_186 (O_186,N_4719,N_4663);
or UO_187 (O_187,N_4943,N_4026);
or UO_188 (O_188,N_4603,N_4009);
nand UO_189 (O_189,N_4858,N_4336);
xnor UO_190 (O_190,N_4326,N_4212);
xnor UO_191 (O_191,N_4668,N_4884);
nor UO_192 (O_192,N_4577,N_4354);
nand UO_193 (O_193,N_4111,N_4184);
nand UO_194 (O_194,N_4300,N_4349);
or UO_195 (O_195,N_4724,N_4198);
nor UO_196 (O_196,N_4050,N_4098);
and UO_197 (O_197,N_4911,N_4610);
or UO_198 (O_198,N_4525,N_4886);
or UO_199 (O_199,N_4488,N_4926);
nor UO_200 (O_200,N_4509,N_4632);
or UO_201 (O_201,N_4046,N_4221);
and UO_202 (O_202,N_4611,N_4821);
or UO_203 (O_203,N_4934,N_4938);
and UO_204 (O_204,N_4018,N_4080);
and UO_205 (O_205,N_4043,N_4475);
nor UO_206 (O_206,N_4253,N_4290);
nand UO_207 (O_207,N_4330,N_4578);
or UO_208 (O_208,N_4768,N_4806);
nand UO_209 (O_209,N_4427,N_4847);
nor UO_210 (O_210,N_4584,N_4927);
and UO_211 (O_211,N_4553,N_4818);
nand UO_212 (O_212,N_4769,N_4512);
xor UO_213 (O_213,N_4473,N_4375);
and UO_214 (O_214,N_4976,N_4670);
and UO_215 (O_215,N_4342,N_4851);
nor UO_216 (O_216,N_4292,N_4979);
and UO_217 (O_217,N_4701,N_4800);
or UO_218 (O_218,N_4772,N_4642);
nand UO_219 (O_219,N_4224,N_4408);
nor UO_220 (O_220,N_4649,N_4143);
and UO_221 (O_221,N_4315,N_4645);
nand UO_222 (O_222,N_4160,N_4978);
nand UO_223 (O_223,N_4653,N_4726);
nand UO_224 (O_224,N_4593,N_4830);
xnor UO_225 (O_225,N_4657,N_4988);
and UO_226 (O_226,N_4405,N_4437);
and UO_227 (O_227,N_4171,N_4550);
and UO_228 (O_228,N_4258,N_4245);
and UO_229 (O_229,N_4930,N_4120);
nor UO_230 (O_230,N_4123,N_4000);
and UO_231 (O_231,N_4209,N_4924);
nor UO_232 (O_232,N_4327,N_4736);
nand UO_233 (O_233,N_4317,N_4394);
and UO_234 (O_234,N_4693,N_4387);
nand UO_235 (O_235,N_4066,N_4414);
and UO_236 (O_236,N_4325,N_4302);
or UO_237 (O_237,N_4287,N_4981);
or UO_238 (O_238,N_4164,N_4313);
nor UO_239 (O_239,N_4921,N_4458);
nor UO_240 (O_240,N_4865,N_4056);
nor UO_241 (O_241,N_4737,N_4454);
nor UO_242 (O_242,N_4154,N_4162);
or UO_243 (O_243,N_4900,N_4656);
nand UO_244 (O_244,N_4440,N_4179);
or UO_245 (O_245,N_4389,N_4156);
and UO_246 (O_246,N_4276,N_4476);
nand UO_247 (O_247,N_4361,N_4449);
or UO_248 (O_248,N_4241,N_4541);
nand UO_249 (O_249,N_4227,N_4137);
nor UO_250 (O_250,N_4983,N_4535);
or UO_251 (O_251,N_4426,N_4236);
or UO_252 (O_252,N_4752,N_4885);
or UO_253 (O_253,N_4622,N_4266);
or UO_254 (O_254,N_4030,N_4540);
nand UO_255 (O_255,N_4436,N_4838);
or UO_256 (O_256,N_4895,N_4438);
nand UO_257 (O_257,N_4231,N_4131);
and UO_258 (O_258,N_4798,N_4075);
nand UO_259 (O_259,N_4684,N_4896);
and UO_260 (O_260,N_4952,N_4447);
nor UO_261 (O_261,N_4260,N_4514);
and UO_262 (O_262,N_4112,N_4853);
or UO_263 (O_263,N_4385,N_4024);
or UO_264 (O_264,N_4861,N_4742);
nand UO_265 (O_265,N_4032,N_4058);
nor UO_266 (O_266,N_4738,N_4487);
nor UO_267 (O_267,N_4646,N_4792);
and UO_268 (O_268,N_4453,N_4304);
or UO_269 (O_269,N_4348,N_4041);
nor UO_270 (O_270,N_4530,N_4989);
and UO_271 (O_271,N_4852,N_4999);
nand UO_272 (O_272,N_4443,N_4694);
nor UO_273 (O_273,N_4378,N_4092);
and UO_274 (O_274,N_4418,N_4906);
xor UO_275 (O_275,N_4707,N_4511);
and UO_276 (O_276,N_4339,N_4229);
or UO_277 (O_277,N_4416,N_4076);
and UO_278 (O_278,N_4107,N_4897);
nor UO_279 (O_279,N_4836,N_4891);
and UO_280 (O_280,N_4547,N_4172);
and UO_281 (O_281,N_4588,N_4936);
nor UO_282 (O_282,N_4581,N_4071);
nand UO_283 (O_283,N_4843,N_4045);
and UO_284 (O_284,N_4170,N_4877);
nor UO_285 (O_285,N_4274,N_4255);
or UO_286 (O_286,N_4365,N_4807);
nand UO_287 (O_287,N_4805,N_4594);
nor UO_288 (O_288,N_4341,N_4721);
and UO_289 (O_289,N_4595,N_4297);
and UO_290 (O_290,N_4363,N_4008);
xnor UO_291 (O_291,N_4636,N_4889);
or UO_292 (O_292,N_4161,N_4467);
nor UO_293 (O_293,N_4014,N_4145);
or UO_294 (O_294,N_4974,N_4675);
nor UO_295 (O_295,N_4908,N_4874);
and UO_296 (O_296,N_4503,N_4432);
and UO_297 (O_297,N_4049,N_4502);
or UO_298 (O_298,N_4573,N_4233);
and UO_299 (O_299,N_4457,N_4228);
nor UO_300 (O_300,N_4469,N_4100);
or UO_301 (O_301,N_4153,N_4239);
nand UO_302 (O_302,N_4845,N_4362);
nor UO_303 (O_303,N_4499,N_4069);
nand UO_304 (O_304,N_4871,N_4659);
nor UO_305 (O_305,N_4623,N_4531);
or UO_306 (O_306,N_4521,N_4789);
or UO_307 (O_307,N_4350,N_4141);
nand UO_308 (O_308,N_4703,N_4731);
nor UO_309 (O_309,N_4682,N_4478);
nand UO_310 (O_310,N_4837,N_4391);
and UO_311 (O_311,N_4068,N_4367);
and UO_312 (O_312,N_4504,N_4323);
or UO_313 (O_313,N_4483,N_4597);
nor UO_314 (O_314,N_4025,N_4053);
and UO_315 (O_315,N_4074,N_4799);
nor UO_316 (O_316,N_4013,N_4903);
or UO_317 (O_317,N_4273,N_4848);
or UO_318 (O_318,N_4866,N_4062);
nand UO_319 (O_319,N_4803,N_4372);
nor UO_320 (O_320,N_4265,N_4021);
or UO_321 (O_321,N_4667,N_4185);
nor UO_322 (O_322,N_4307,N_4462);
nor UO_323 (O_323,N_4177,N_4034);
nor UO_324 (O_324,N_4152,N_4140);
and UO_325 (O_325,N_4956,N_4169);
and UO_326 (O_326,N_4093,N_4482);
nor UO_327 (O_327,N_4994,N_4894);
and UO_328 (O_328,N_4892,N_4082);
and UO_329 (O_329,N_4904,N_4777);
nand UO_330 (O_330,N_4700,N_4246);
and UO_331 (O_331,N_4480,N_4380);
or UO_332 (O_332,N_4625,N_4196);
nand UO_333 (O_333,N_4902,N_4301);
nor UO_334 (O_334,N_4351,N_4917);
nor UO_335 (O_335,N_4490,N_4109);
nand UO_336 (O_336,N_4711,N_4127);
nand UO_337 (O_337,N_4991,N_4148);
or UO_338 (O_338,N_4549,N_4608);
or UO_339 (O_339,N_4004,N_4486);
nor UO_340 (O_340,N_4225,N_4880);
nand UO_341 (O_341,N_4941,N_4743);
or UO_342 (O_342,N_4303,N_4446);
nor UO_343 (O_343,N_4775,N_4286);
nor UO_344 (O_344,N_4801,N_4932);
or UO_345 (O_345,N_4051,N_4489);
and UO_346 (O_346,N_4812,N_4244);
and UO_347 (O_347,N_4704,N_4277);
or UO_348 (O_348,N_4788,N_4804);
or UO_349 (O_349,N_4968,N_4491);
and UO_350 (O_350,N_4560,N_4377);
and UO_351 (O_351,N_4424,N_4322);
and UO_352 (O_352,N_4410,N_4970);
nor UO_353 (O_353,N_4846,N_4108);
or UO_354 (O_354,N_4699,N_4685);
and UO_355 (O_355,N_4556,N_4501);
and UO_356 (O_356,N_4571,N_4929);
or UO_357 (O_357,N_4282,N_4561);
and UO_358 (O_358,N_4898,N_4734);
nand UO_359 (O_359,N_4240,N_4596);
and UO_360 (O_360,N_4002,N_4073);
nor UO_361 (O_361,N_4820,N_4815);
nor UO_362 (O_362,N_4033,N_4012);
or UO_363 (O_363,N_4321,N_4739);
or UO_364 (O_364,N_4716,N_4592);
nand UO_365 (O_365,N_4605,N_4893);
and UO_366 (O_366,N_4559,N_4421);
nand UO_367 (O_367,N_4019,N_4333);
nand UO_368 (O_368,N_4631,N_4477);
and UO_369 (O_369,N_4939,N_4078);
or UO_370 (O_370,N_4132,N_4949);
and UO_371 (O_371,N_4975,N_4602);
nor UO_372 (O_372,N_4011,N_4017);
or UO_373 (O_373,N_4606,N_4343);
or UO_374 (O_374,N_4966,N_4840);
or UO_375 (O_375,N_4948,N_4283);
nand UO_376 (O_376,N_4298,N_4787);
and UO_377 (O_377,N_4654,N_4099);
nand UO_378 (O_378,N_4925,N_4215);
nand UO_379 (O_379,N_4633,N_4319);
or UO_380 (O_380,N_4899,N_4364);
nand UO_381 (O_381,N_4958,N_4186);
or UO_382 (O_382,N_4085,N_4875);
nor UO_383 (O_383,N_4158,N_4533);
nor UO_384 (O_384,N_4790,N_4175);
nand UO_385 (O_385,N_4506,N_4519);
or UO_386 (O_386,N_4945,N_4940);
nor UO_387 (O_387,N_4293,N_4059);
nand UO_388 (O_388,N_4356,N_4207);
or UO_389 (O_389,N_4360,N_4944);
and UO_390 (O_390,N_4110,N_4150);
nor UO_391 (O_391,N_4713,N_4679);
or UO_392 (O_392,N_4188,N_4401);
nor UO_393 (O_393,N_4434,N_4913);
and UO_394 (O_394,N_4411,N_4627);
nor UO_395 (O_395,N_4331,N_4873);
nand UO_396 (O_396,N_4964,N_4727);
nor UO_397 (O_397,N_4635,N_4183);
or UO_398 (O_398,N_4257,N_4226);
or UO_399 (O_399,N_4720,N_4249);
nor UO_400 (O_400,N_4190,N_4346);
and UO_401 (O_401,N_4572,N_4182);
or UO_402 (O_402,N_4779,N_4393);
nor UO_403 (O_403,N_4379,N_4658);
nand UO_404 (O_404,N_4464,N_4335);
nor UO_405 (O_405,N_4116,N_4993);
or UO_406 (O_406,N_4689,N_4557);
nor UO_407 (O_407,N_4113,N_4369);
nand UO_408 (O_408,N_4576,N_4601);
and UO_409 (O_409,N_4982,N_4516);
xnor UO_410 (O_410,N_4780,N_4860);
nand UO_411 (O_411,N_4268,N_4201);
nand UO_412 (O_412,N_4725,N_4854);
and UO_413 (O_413,N_4118,N_4347);
and UO_414 (O_414,N_4455,N_4206);
nor UO_415 (O_415,N_4650,N_4542);
and UO_416 (O_416,N_4208,N_4527);
nand UO_417 (O_417,N_4660,N_4001);
or UO_418 (O_418,N_4915,N_4392);
nor UO_419 (O_419,N_4850,N_4995);
and UO_420 (O_420,N_4680,N_4195);
nand UO_421 (O_421,N_4271,N_4692);
or UO_422 (O_422,N_4395,N_4187);
nor UO_423 (O_423,N_4613,N_4674);
or UO_424 (O_424,N_4305,N_4839);
nand UO_425 (O_425,N_4400,N_4420);
and UO_426 (O_426,N_4589,N_4269);
nand UO_427 (O_427,N_4402,N_4106);
or UO_428 (O_428,N_4604,N_4097);
nor UO_429 (O_429,N_4200,N_4959);
nor UO_430 (O_430,N_4686,N_4357);
or UO_431 (O_431,N_4825,N_4210);
nor UO_432 (O_432,N_4690,N_4067);
nand UO_433 (O_433,N_4980,N_4407);
and UO_434 (O_434,N_4077,N_4834);
nand UO_435 (O_435,N_4445,N_4010);
and UO_436 (O_436,N_4651,N_4551);
nand UO_437 (O_437,N_4570,N_4677);
xnor UO_438 (O_438,N_4676,N_4197);
or UO_439 (O_439,N_4316,N_4383);
nor UO_440 (O_440,N_4709,N_4284);
nor UO_441 (O_441,N_4808,N_4320);
or UO_442 (O_442,N_4252,N_4986);
nor UO_443 (O_443,N_4057,N_4732);
and UO_444 (O_444,N_4461,N_4914);
nor UO_445 (O_445,N_4345,N_4857);
and UO_446 (O_446,N_4912,N_4505);
or UO_447 (O_447,N_4961,N_4765);
or UO_448 (O_448,N_4222,N_4782);
nor UO_449 (O_449,N_4624,N_4714);
or UO_450 (O_450,N_4829,N_4543);
nor UO_451 (O_451,N_4844,N_4916);
and UO_452 (O_452,N_4399,N_4575);
nor UO_453 (O_453,N_4767,N_4353);
nand UO_454 (O_454,N_4481,N_4582);
nor UO_455 (O_455,N_4520,N_4729);
nor UO_456 (O_456,N_4272,N_4494);
nor UO_457 (O_457,N_4907,N_4683);
and UO_458 (O_458,N_4954,N_4498);
or UO_459 (O_459,N_4817,N_4036);
or UO_460 (O_460,N_4428,N_4887);
nor UO_461 (O_461,N_4397,N_4291);
nand UO_462 (O_462,N_4580,N_4384);
nand UO_463 (O_463,N_4088,N_4279);
and UO_464 (O_464,N_4664,N_4809);
or UO_465 (O_465,N_4733,N_4728);
nor UO_466 (O_466,N_4178,N_4040);
nand UO_467 (O_467,N_4133,N_4796);
and UO_468 (O_468,N_4638,N_4751);
or UO_469 (O_469,N_4308,N_4090);
nand UO_470 (O_470,N_4640,N_4537);
and UO_471 (O_471,N_4770,N_4666);
nand UO_472 (O_472,N_4614,N_4135);
and UO_473 (O_473,N_4031,N_4607);
and UO_474 (O_474,N_4598,N_4117);
or UO_475 (O_475,N_4167,N_4103);
and UO_476 (O_476,N_4465,N_4591);
and UO_477 (O_477,N_4061,N_4987);
xnor UO_478 (O_478,N_4439,N_4027);
or UO_479 (O_479,N_4795,N_4299);
and UO_480 (O_480,N_4038,N_4382);
or UO_481 (O_481,N_4390,N_4842);
xnor UO_482 (O_482,N_4007,N_4621);
or UO_483 (O_483,N_4985,N_4747);
nand UO_484 (O_484,N_4413,N_4662);
nand UO_485 (O_485,N_4629,N_4294);
nor UO_486 (O_486,N_4119,N_4586);
or UO_487 (O_487,N_4285,N_4515);
nand UO_488 (O_488,N_4984,N_4992);
nand UO_489 (O_489,N_4124,N_4849);
or UO_490 (O_490,N_4630,N_4583);
nand UO_491 (O_491,N_4329,N_4832);
nand UO_492 (O_492,N_4079,N_4918);
and UO_493 (O_493,N_4615,N_4060);
nor UO_494 (O_494,N_4396,N_4192);
nor UO_495 (O_495,N_4338,N_4005);
nand UO_496 (O_496,N_4639,N_4430);
or UO_497 (O_497,N_4859,N_4205);
nor UO_498 (O_498,N_4637,N_4429);
or UO_499 (O_499,N_4532,N_4275);
and UO_500 (O_500,N_4564,N_4928);
nand UO_501 (O_501,N_4552,N_4491);
nor UO_502 (O_502,N_4739,N_4626);
nor UO_503 (O_503,N_4161,N_4259);
and UO_504 (O_504,N_4496,N_4179);
or UO_505 (O_505,N_4463,N_4027);
nor UO_506 (O_506,N_4131,N_4326);
and UO_507 (O_507,N_4128,N_4245);
nor UO_508 (O_508,N_4094,N_4858);
and UO_509 (O_509,N_4745,N_4597);
and UO_510 (O_510,N_4199,N_4655);
nand UO_511 (O_511,N_4612,N_4986);
and UO_512 (O_512,N_4952,N_4912);
and UO_513 (O_513,N_4352,N_4389);
or UO_514 (O_514,N_4434,N_4715);
nor UO_515 (O_515,N_4573,N_4705);
nand UO_516 (O_516,N_4967,N_4021);
and UO_517 (O_517,N_4624,N_4324);
nand UO_518 (O_518,N_4451,N_4135);
nor UO_519 (O_519,N_4644,N_4362);
and UO_520 (O_520,N_4287,N_4232);
and UO_521 (O_521,N_4724,N_4789);
nor UO_522 (O_522,N_4406,N_4178);
nand UO_523 (O_523,N_4102,N_4914);
nor UO_524 (O_524,N_4203,N_4371);
nand UO_525 (O_525,N_4985,N_4424);
nand UO_526 (O_526,N_4602,N_4655);
nand UO_527 (O_527,N_4320,N_4442);
nand UO_528 (O_528,N_4279,N_4608);
or UO_529 (O_529,N_4085,N_4152);
nor UO_530 (O_530,N_4443,N_4782);
nand UO_531 (O_531,N_4757,N_4446);
nor UO_532 (O_532,N_4734,N_4994);
nor UO_533 (O_533,N_4262,N_4287);
nand UO_534 (O_534,N_4364,N_4144);
nor UO_535 (O_535,N_4773,N_4711);
or UO_536 (O_536,N_4731,N_4724);
or UO_537 (O_537,N_4527,N_4936);
and UO_538 (O_538,N_4911,N_4030);
and UO_539 (O_539,N_4922,N_4880);
or UO_540 (O_540,N_4974,N_4321);
and UO_541 (O_541,N_4275,N_4099);
nand UO_542 (O_542,N_4365,N_4055);
or UO_543 (O_543,N_4462,N_4735);
nand UO_544 (O_544,N_4789,N_4482);
or UO_545 (O_545,N_4819,N_4722);
and UO_546 (O_546,N_4868,N_4188);
and UO_547 (O_547,N_4817,N_4355);
or UO_548 (O_548,N_4179,N_4626);
nand UO_549 (O_549,N_4239,N_4869);
nor UO_550 (O_550,N_4776,N_4989);
nand UO_551 (O_551,N_4299,N_4925);
or UO_552 (O_552,N_4199,N_4789);
nor UO_553 (O_553,N_4620,N_4832);
or UO_554 (O_554,N_4422,N_4612);
nor UO_555 (O_555,N_4282,N_4903);
nor UO_556 (O_556,N_4061,N_4690);
and UO_557 (O_557,N_4231,N_4858);
nand UO_558 (O_558,N_4013,N_4099);
nor UO_559 (O_559,N_4600,N_4070);
or UO_560 (O_560,N_4284,N_4584);
nor UO_561 (O_561,N_4233,N_4975);
nand UO_562 (O_562,N_4735,N_4085);
nor UO_563 (O_563,N_4552,N_4961);
nand UO_564 (O_564,N_4458,N_4692);
and UO_565 (O_565,N_4871,N_4996);
nor UO_566 (O_566,N_4684,N_4970);
nand UO_567 (O_567,N_4555,N_4127);
and UO_568 (O_568,N_4278,N_4646);
and UO_569 (O_569,N_4294,N_4540);
and UO_570 (O_570,N_4563,N_4227);
nand UO_571 (O_571,N_4012,N_4556);
nand UO_572 (O_572,N_4627,N_4912);
nor UO_573 (O_573,N_4345,N_4882);
and UO_574 (O_574,N_4589,N_4925);
or UO_575 (O_575,N_4451,N_4019);
and UO_576 (O_576,N_4731,N_4638);
nand UO_577 (O_577,N_4149,N_4631);
and UO_578 (O_578,N_4774,N_4011);
and UO_579 (O_579,N_4856,N_4012);
or UO_580 (O_580,N_4721,N_4479);
and UO_581 (O_581,N_4548,N_4814);
nor UO_582 (O_582,N_4328,N_4364);
nor UO_583 (O_583,N_4051,N_4242);
and UO_584 (O_584,N_4267,N_4166);
nand UO_585 (O_585,N_4001,N_4208);
nor UO_586 (O_586,N_4084,N_4315);
or UO_587 (O_587,N_4234,N_4646);
or UO_588 (O_588,N_4453,N_4365);
nand UO_589 (O_589,N_4103,N_4349);
or UO_590 (O_590,N_4970,N_4157);
nor UO_591 (O_591,N_4768,N_4486);
nand UO_592 (O_592,N_4212,N_4050);
or UO_593 (O_593,N_4913,N_4397);
or UO_594 (O_594,N_4370,N_4355);
nor UO_595 (O_595,N_4158,N_4787);
nand UO_596 (O_596,N_4437,N_4852);
nor UO_597 (O_597,N_4044,N_4314);
or UO_598 (O_598,N_4376,N_4202);
nor UO_599 (O_599,N_4962,N_4518);
nor UO_600 (O_600,N_4347,N_4548);
nand UO_601 (O_601,N_4886,N_4142);
nor UO_602 (O_602,N_4293,N_4886);
or UO_603 (O_603,N_4683,N_4806);
nor UO_604 (O_604,N_4087,N_4776);
nor UO_605 (O_605,N_4158,N_4989);
or UO_606 (O_606,N_4998,N_4350);
xnor UO_607 (O_607,N_4062,N_4602);
nor UO_608 (O_608,N_4858,N_4689);
or UO_609 (O_609,N_4338,N_4678);
or UO_610 (O_610,N_4450,N_4436);
nor UO_611 (O_611,N_4748,N_4815);
nand UO_612 (O_612,N_4742,N_4102);
nor UO_613 (O_613,N_4690,N_4027);
nor UO_614 (O_614,N_4298,N_4193);
or UO_615 (O_615,N_4581,N_4128);
nor UO_616 (O_616,N_4278,N_4595);
and UO_617 (O_617,N_4143,N_4365);
nand UO_618 (O_618,N_4736,N_4722);
and UO_619 (O_619,N_4173,N_4080);
or UO_620 (O_620,N_4883,N_4181);
nor UO_621 (O_621,N_4775,N_4030);
and UO_622 (O_622,N_4200,N_4775);
or UO_623 (O_623,N_4808,N_4711);
or UO_624 (O_624,N_4493,N_4239);
nor UO_625 (O_625,N_4979,N_4854);
and UO_626 (O_626,N_4044,N_4717);
nor UO_627 (O_627,N_4409,N_4474);
or UO_628 (O_628,N_4526,N_4545);
nor UO_629 (O_629,N_4705,N_4748);
nand UO_630 (O_630,N_4764,N_4772);
nand UO_631 (O_631,N_4184,N_4965);
or UO_632 (O_632,N_4483,N_4570);
and UO_633 (O_633,N_4907,N_4856);
nor UO_634 (O_634,N_4213,N_4372);
nor UO_635 (O_635,N_4294,N_4256);
or UO_636 (O_636,N_4008,N_4596);
nand UO_637 (O_637,N_4654,N_4197);
or UO_638 (O_638,N_4704,N_4491);
nand UO_639 (O_639,N_4824,N_4773);
nand UO_640 (O_640,N_4847,N_4124);
nand UO_641 (O_641,N_4960,N_4836);
nand UO_642 (O_642,N_4170,N_4270);
or UO_643 (O_643,N_4833,N_4871);
nand UO_644 (O_644,N_4589,N_4683);
or UO_645 (O_645,N_4583,N_4744);
nand UO_646 (O_646,N_4634,N_4621);
or UO_647 (O_647,N_4049,N_4828);
nor UO_648 (O_648,N_4880,N_4989);
and UO_649 (O_649,N_4596,N_4937);
and UO_650 (O_650,N_4272,N_4937);
nand UO_651 (O_651,N_4898,N_4700);
and UO_652 (O_652,N_4993,N_4065);
nor UO_653 (O_653,N_4564,N_4225);
and UO_654 (O_654,N_4273,N_4138);
nand UO_655 (O_655,N_4234,N_4926);
or UO_656 (O_656,N_4410,N_4901);
and UO_657 (O_657,N_4309,N_4924);
nor UO_658 (O_658,N_4572,N_4835);
or UO_659 (O_659,N_4527,N_4913);
nand UO_660 (O_660,N_4809,N_4339);
nand UO_661 (O_661,N_4813,N_4286);
or UO_662 (O_662,N_4783,N_4855);
nor UO_663 (O_663,N_4122,N_4123);
and UO_664 (O_664,N_4350,N_4752);
nor UO_665 (O_665,N_4966,N_4668);
and UO_666 (O_666,N_4008,N_4904);
nand UO_667 (O_667,N_4672,N_4775);
or UO_668 (O_668,N_4185,N_4585);
or UO_669 (O_669,N_4104,N_4667);
nor UO_670 (O_670,N_4136,N_4651);
and UO_671 (O_671,N_4861,N_4867);
and UO_672 (O_672,N_4915,N_4455);
nor UO_673 (O_673,N_4768,N_4159);
nor UO_674 (O_674,N_4095,N_4521);
or UO_675 (O_675,N_4083,N_4193);
and UO_676 (O_676,N_4541,N_4494);
nor UO_677 (O_677,N_4677,N_4449);
or UO_678 (O_678,N_4492,N_4356);
and UO_679 (O_679,N_4284,N_4231);
or UO_680 (O_680,N_4531,N_4353);
nor UO_681 (O_681,N_4199,N_4227);
xor UO_682 (O_682,N_4190,N_4284);
or UO_683 (O_683,N_4190,N_4669);
nor UO_684 (O_684,N_4255,N_4848);
nand UO_685 (O_685,N_4406,N_4119);
or UO_686 (O_686,N_4936,N_4410);
and UO_687 (O_687,N_4195,N_4843);
nand UO_688 (O_688,N_4106,N_4364);
nand UO_689 (O_689,N_4475,N_4272);
nor UO_690 (O_690,N_4283,N_4217);
and UO_691 (O_691,N_4054,N_4057);
nor UO_692 (O_692,N_4654,N_4408);
or UO_693 (O_693,N_4636,N_4475);
nor UO_694 (O_694,N_4718,N_4636);
or UO_695 (O_695,N_4235,N_4539);
or UO_696 (O_696,N_4633,N_4814);
or UO_697 (O_697,N_4067,N_4190);
nand UO_698 (O_698,N_4908,N_4397);
nand UO_699 (O_699,N_4108,N_4326);
nor UO_700 (O_700,N_4342,N_4747);
nand UO_701 (O_701,N_4558,N_4343);
or UO_702 (O_702,N_4476,N_4256);
nor UO_703 (O_703,N_4099,N_4192);
and UO_704 (O_704,N_4389,N_4144);
and UO_705 (O_705,N_4528,N_4094);
and UO_706 (O_706,N_4066,N_4043);
and UO_707 (O_707,N_4976,N_4475);
nand UO_708 (O_708,N_4486,N_4297);
and UO_709 (O_709,N_4203,N_4535);
and UO_710 (O_710,N_4005,N_4436);
nor UO_711 (O_711,N_4922,N_4001);
and UO_712 (O_712,N_4749,N_4995);
or UO_713 (O_713,N_4540,N_4229);
or UO_714 (O_714,N_4101,N_4427);
xor UO_715 (O_715,N_4187,N_4258);
and UO_716 (O_716,N_4095,N_4111);
nor UO_717 (O_717,N_4931,N_4297);
nand UO_718 (O_718,N_4841,N_4011);
nand UO_719 (O_719,N_4332,N_4707);
or UO_720 (O_720,N_4508,N_4296);
or UO_721 (O_721,N_4600,N_4583);
nor UO_722 (O_722,N_4005,N_4579);
and UO_723 (O_723,N_4640,N_4452);
or UO_724 (O_724,N_4564,N_4043);
nand UO_725 (O_725,N_4323,N_4753);
nor UO_726 (O_726,N_4451,N_4549);
nor UO_727 (O_727,N_4589,N_4919);
xor UO_728 (O_728,N_4735,N_4066);
nor UO_729 (O_729,N_4339,N_4606);
or UO_730 (O_730,N_4376,N_4578);
nor UO_731 (O_731,N_4348,N_4589);
or UO_732 (O_732,N_4580,N_4694);
and UO_733 (O_733,N_4080,N_4954);
nor UO_734 (O_734,N_4133,N_4116);
nand UO_735 (O_735,N_4225,N_4318);
or UO_736 (O_736,N_4818,N_4432);
nor UO_737 (O_737,N_4252,N_4853);
nor UO_738 (O_738,N_4788,N_4559);
nand UO_739 (O_739,N_4982,N_4041);
or UO_740 (O_740,N_4047,N_4665);
or UO_741 (O_741,N_4583,N_4275);
and UO_742 (O_742,N_4329,N_4531);
and UO_743 (O_743,N_4541,N_4584);
and UO_744 (O_744,N_4958,N_4733);
nor UO_745 (O_745,N_4442,N_4435);
nand UO_746 (O_746,N_4945,N_4540);
or UO_747 (O_747,N_4158,N_4477);
and UO_748 (O_748,N_4496,N_4004);
nand UO_749 (O_749,N_4508,N_4353);
and UO_750 (O_750,N_4233,N_4881);
nor UO_751 (O_751,N_4554,N_4728);
or UO_752 (O_752,N_4983,N_4229);
nor UO_753 (O_753,N_4648,N_4713);
xor UO_754 (O_754,N_4786,N_4217);
and UO_755 (O_755,N_4814,N_4550);
and UO_756 (O_756,N_4079,N_4495);
and UO_757 (O_757,N_4394,N_4383);
and UO_758 (O_758,N_4415,N_4214);
or UO_759 (O_759,N_4658,N_4333);
or UO_760 (O_760,N_4675,N_4356);
nand UO_761 (O_761,N_4651,N_4401);
and UO_762 (O_762,N_4868,N_4674);
nor UO_763 (O_763,N_4996,N_4530);
or UO_764 (O_764,N_4677,N_4813);
nand UO_765 (O_765,N_4259,N_4217);
nand UO_766 (O_766,N_4698,N_4556);
nand UO_767 (O_767,N_4554,N_4718);
nor UO_768 (O_768,N_4675,N_4079);
and UO_769 (O_769,N_4664,N_4553);
nand UO_770 (O_770,N_4559,N_4675);
nand UO_771 (O_771,N_4579,N_4479);
and UO_772 (O_772,N_4394,N_4963);
nand UO_773 (O_773,N_4428,N_4455);
and UO_774 (O_774,N_4061,N_4578);
and UO_775 (O_775,N_4076,N_4185);
nor UO_776 (O_776,N_4855,N_4278);
or UO_777 (O_777,N_4477,N_4331);
nor UO_778 (O_778,N_4853,N_4516);
and UO_779 (O_779,N_4084,N_4882);
or UO_780 (O_780,N_4064,N_4068);
nand UO_781 (O_781,N_4974,N_4016);
or UO_782 (O_782,N_4937,N_4961);
and UO_783 (O_783,N_4480,N_4913);
nand UO_784 (O_784,N_4804,N_4406);
nand UO_785 (O_785,N_4220,N_4219);
nor UO_786 (O_786,N_4170,N_4774);
nor UO_787 (O_787,N_4258,N_4280);
or UO_788 (O_788,N_4069,N_4868);
nor UO_789 (O_789,N_4335,N_4847);
nor UO_790 (O_790,N_4207,N_4492);
nor UO_791 (O_791,N_4496,N_4538);
nand UO_792 (O_792,N_4729,N_4790);
or UO_793 (O_793,N_4625,N_4786);
nand UO_794 (O_794,N_4834,N_4205);
nor UO_795 (O_795,N_4056,N_4377);
nand UO_796 (O_796,N_4879,N_4812);
nor UO_797 (O_797,N_4050,N_4329);
nor UO_798 (O_798,N_4698,N_4768);
xnor UO_799 (O_799,N_4413,N_4267);
and UO_800 (O_800,N_4953,N_4948);
nor UO_801 (O_801,N_4512,N_4203);
or UO_802 (O_802,N_4094,N_4785);
nor UO_803 (O_803,N_4387,N_4702);
nor UO_804 (O_804,N_4132,N_4989);
and UO_805 (O_805,N_4862,N_4261);
and UO_806 (O_806,N_4570,N_4562);
nand UO_807 (O_807,N_4832,N_4210);
or UO_808 (O_808,N_4600,N_4316);
or UO_809 (O_809,N_4289,N_4404);
and UO_810 (O_810,N_4819,N_4061);
and UO_811 (O_811,N_4173,N_4442);
nand UO_812 (O_812,N_4188,N_4514);
or UO_813 (O_813,N_4388,N_4646);
nand UO_814 (O_814,N_4454,N_4835);
or UO_815 (O_815,N_4852,N_4925);
and UO_816 (O_816,N_4516,N_4986);
nor UO_817 (O_817,N_4310,N_4542);
nor UO_818 (O_818,N_4265,N_4737);
and UO_819 (O_819,N_4313,N_4206);
nor UO_820 (O_820,N_4222,N_4306);
and UO_821 (O_821,N_4779,N_4751);
nor UO_822 (O_822,N_4401,N_4572);
or UO_823 (O_823,N_4345,N_4778);
nand UO_824 (O_824,N_4301,N_4640);
xnor UO_825 (O_825,N_4945,N_4771);
nand UO_826 (O_826,N_4409,N_4482);
and UO_827 (O_827,N_4946,N_4484);
nor UO_828 (O_828,N_4657,N_4639);
nor UO_829 (O_829,N_4794,N_4842);
nor UO_830 (O_830,N_4585,N_4341);
or UO_831 (O_831,N_4626,N_4078);
and UO_832 (O_832,N_4800,N_4863);
nand UO_833 (O_833,N_4411,N_4744);
nand UO_834 (O_834,N_4144,N_4397);
nand UO_835 (O_835,N_4537,N_4481);
nor UO_836 (O_836,N_4185,N_4306);
nand UO_837 (O_837,N_4586,N_4524);
nand UO_838 (O_838,N_4666,N_4320);
nand UO_839 (O_839,N_4996,N_4094);
nand UO_840 (O_840,N_4627,N_4677);
nand UO_841 (O_841,N_4748,N_4036);
nand UO_842 (O_842,N_4412,N_4804);
nand UO_843 (O_843,N_4219,N_4312);
and UO_844 (O_844,N_4037,N_4007);
or UO_845 (O_845,N_4676,N_4229);
nand UO_846 (O_846,N_4335,N_4307);
or UO_847 (O_847,N_4671,N_4824);
nor UO_848 (O_848,N_4761,N_4472);
nand UO_849 (O_849,N_4328,N_4389);
and UO_850 (O_850,N_4140,N_4260);
nor UO_851 (O_851,N_4967,N_4324);
nor UO_852 (O_852,N_4729,N_4484);
nor UO_853 (O_853,N_4395,N_4358);
and UO_854 (O_854,N_4142,N_4277);
nor UO_855 (O_855,N_4398,N_4391);
nor UO_856 (O_856,N_4486,N_4376);
or UO_857 (O_857,N_4753,N_4820);
nor UO_858 (O_858,N_4758,N_4538);
nand UO_859 (O_859,N_4761,N_4393);
or UO_860 (O_860,N_4395,N_4881);
and UO_861 (O_861,N_4301,N_4627);
nand UO_862 (O_862,N_4149,N_4731);
nor UO_863 (O_863,N_4222,N_4165);
nor UO_864 (O_864,N_4225,N_4140);
nor UO_865 (O_865,N_4272,N_4761);
nand UO_866 (O_866,N_4343,N_4227);
nor UO_867 (O_867,N_4240,N_4327);
nand UO_868 (O_868,N_4197,N_4032);
or UO_869 (O_869,N_4669,N_4497);
and UO_870 (O_870,N_4026,N_4651);
and UO_871 (O_871,N_4467,N_4735);
nand UO_872 (O_872,N_4076,N_4271);
nor UO_873 (O_873,N_4714,N_4800);
or UO_874 (O_874,N_4912,N_4899);
nand UO_875 (O_875,N_4159,N_4916);
or UO_876 (O_876,N_4336,N_4053);
or UO_877 (O_877,N_4206,N_4597);
and UO_878 (O_878,N_4283,N_4907);
or UO_879 (O_879,N_4842,N_4125);
or UO_880 (O_880,N_4387,N_4040);
or UO_881 (O_881,N_4153,N_4855);
and UO_882 (O_882,N_4283,N_4744);
nand UO_883 (O_883,N_4972,N_4502);
and UO_884 (O_884,N_4867,N_4167);
nor UO_885 (O_885,N_4247,N_4566);
nand UO_886 (O_886,N_4365,N_4115);
nor UO_887 (O_887,N_4290,N_4906);
nand UO_888 (O_888,N_4657,N_4838);
nor UO_889 (O_889,N_4732,N_4157);
and UO_890 (O_890,N_4756,N_4829);
nand UO_891 (O_891,N_4023,N_4220);
or UO_892 (O_892,N_4291,N_4271);
nor UO_893 (O_893,N_4164,N_4120);
nand UO_894 (O_894,N_4021,N_4224);
nand UO_895 (O_895,N_4606,N_4432);
nor UO_896 (O_896,N_4040,N_4112);
nor UO_897 (O_897,N_4389,N_4047);
or UO_898 (O_898,N_4215,N_4700);
nor UO_899 (O_899,N_4630,N_4313);
or UO_900 (O_900,N_4276,N_4111);
and UO_901 (O_901,N_4862,N_4983);
nor UO_902 (O_902,N_4256,N_4931);
nand UO_903 (O_903,N_4479,N_4627);
or UO_904 (O_904,N_4956,N_4717);
nand UO_905 (O_905,N_4810,N_4428);
nor UO_906 (O_906,N_4844,N_4792);
or UO_907 (O_907,N_4802,N_4954);
nand UO_908 (O_908,N_4159,N_4329);
nor UO_909 (O_909,N_4036,N_4077);
nand UO_910 (O_910,N_4649,N_4667);
nand UO_911 (O_911,N_4149,N_4909);
and UO_912 (O_912,N_4729,N_4606);
or UO_913 (O_913,N_4450,N_4913);
nand UO_914 (O_914,N_4010,N_4516);
or UO_915 (O_915,N_4911,N_4348);
or UO_916 (O_916,N_4091,N_4980);
or UO_917 (O_917,N_4918,N_4146);
or UO_918 (O_918,N_4029,N_4698);
nand UO_919 (O_919,N_4944,N_4055);
nand UO_920 (O_920,N_4916,N_4332);
or UO_921 (O_921,N_4510,N_4459);
and UO_922 (O_922,N_4855,N_4919);
or UO_923 (O_923,N_4256,N_4833);
nor UO_924 (O_924,N_4322,N_4525);
and UO_925 (O_925,N_4468,N_4573);
nand UO_926 (O_926,N_4379,N_4759);
nand UO_927 (O_927,N_4772,N_4312);
or UO_928 (O_928,N_4263,N_4442);
nand UO_929 (O_929,N_4294,N_4870);
nand UO_930 (O_930,N_4388,N_4400);
or UO_931 (O_931,N_4490,N_4592);
or UO_932 (O_932,N_4485,N_4378);
nor UO_933 (O_933,N_4817,N_4283);
nand UO_934 (O_934,N_4553,N_4642);
or UO_935 (O_935,N_4899,N_4751);
or UO_936 (O_936,N_4034,N_4161);
or UO_937 (O_937,N_4534,N_4731);
nor UO_938 (O_938,N_4540,N_4601);
nor UO_939 (O_939,N_4216,N_4888);
or UO_940 (O_940,N_4471,N_4282);
or UO_941 (O_941,N_4194,N_4259);
nor UO_942 (O_942,N_4032,N_4409);
nand UO_943 (O_943,N_4173,N_4586);
nor UO_944 (O_944,N_4690,N_4857);
and UO_945 (O_945,N_4910,N_4338);
nor UO_946 (O_946,N_4650,N_4113);
nand UO_947 (O_947,N_4130,N_4085);
nor UO_948 (O_948,N_4812,N_4483);
or UO_949 (O_949,N_4129,N_4184);
and UO_950 (O_950,N_4170,N_4857);
nor UO_951 (O_951,N_4676,N_4245);
and UO_952 (O_952,N_4321,N_4093);
nand UO_953 (O_953,N_4471,N_4614);
or UO_954 (O_954,N_4588,N_4537);
and UO_955 (O_955,N_4293,N_4600);
or UO_956 (O_956,N_4002,N_4534);
nand UO_957 (O_957,N_4437,N_4177);
nand UO_958 (O_958,N_4610,N_4768);
and UO_959 (O_959,N_4339,N_4981);
and UO_960 (O_960,N_4813,N_4425);
nand UO_961 (O_961,N_4592,N_4059);
or UO_962 (O_962,N_4901,N_4669);
or UO_963 (O_963,N_4625,N_4604);
and UO_964 (O_964,N_4792,N_4917);
nand UO_965 (O_965,N_4176,N_4355);
and UO_966 (O_966,N_4412,N_4236);
nor UO_967 (O_967,N_4643,N_4868);
nor UO_968 (O_968,N_4946,N_4146);
and UO_969 (O_969,N_4669,N_4712);
nand UO_970 (O_970,N_4721,N_4922);
and UO_971 (O_971,N_4360,N_4167);
and UO_972 (O_972,N_4872,N_4916);
nor UO_973 (O_973,N_4601,N_4412);
and UO_974 (O_974,N_4829,N_4908);
or UO_975 (O_975,N_4356,N_4831);
and UO_976 (O_976,N_4623,N_4986);
nand UO_977 (O_977,N_4937,N_4174);
or UO_978 (O_978,N_4466,N_4133);
nor UO_979 (O_979,N_4567,N_4992);
or UO_980 (O_980,N_4884,N_4741);
nor UO_981 (O_981,N_4714,N_4822);
or UO_982 (O_982,N_4823,N_4044);
nor UO_983 (O_983,N_4534,N_4170);
or UO_984 (O_984,N_4276,N_4326);
nand UO_985 (O_985,N_4978,N_4179);
xor UO_986 (O_986,N_4626,N_4741);
nor UO_987 (O_987,N_4777,N_4092);
nand UO_988 (O_988,N_4136,N_4042);
nand UO_989 (O_989,N_4402,N_4934);
or UO_990 (O_990,N_4065,N_4570);
or UO_991 (O_991,N_4826,N_4454);
nand UO_992 (O_992,N_4020,N_4122);
nand UO_993 (O_993,N_4095,N_4858);
nand UO_994 (O_994,N_4898,N_4991);
nor UO_995 (O_995,N_4432,N_4587);
nand UO_996 (O_996,N_4430,N_4634);
nand UO_997 (O_997,N_4990,N_4057);
nor UO_998 (O_998,N_4429,N_4522);
nand UO_999 (O_999,N_4763,N_4902);
endmodule